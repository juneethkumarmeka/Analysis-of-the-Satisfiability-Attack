module basic_1000_10000_1500_5_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_667,In_981);
nand U1 (N_1,In_230,In_715);
nand U2 (N_2,In_85,In_849);
and U3 (N_3,In_990,In_30);
and U4 (N_4,In_743,In_323);
nand U5 (N_5,In_569,In_185);
or U6 (N_6,In_695,In_589);
nand U7 (N_7,In_196,In_79);
nor U8 (N_8,In_699,In_255);
nor U9 (N_9,In_174,In_385);
or U10 (N_10,In_438,In_409);
nor U11 (N_11,In_198,In_908);
or U12 (N_12,In_959,In_77);
or U13 (N_13,In_577,In_962);
and U14 (N_14,In_756,In_413);
nor U15 (N_15,In_456,In_750);
and U16 (N_16,In_712,In_175);
nor U17 (N_17,In_860,In_274);
or U18 (N_18,In_247,In_843);
and U19 (N_19,In_298,In_925);
and U20 (N_20,In_285,In_625);
or U21 (N_21,In_958,In_53);
or U22 (N_22,In_565,In_499);
and U23 (N_23,In_273,In_143);
nor U24 (N_24,In_523,In_878);
nand U25 (N_25,In_311,In_360);
or U26 (N_26,In_21,In_113);
xnor U27 (N_27,In_633,In_339);
and U28 (N_28,In_834,In_295);
or U29 (N_29,In_294,In_514);
nor U30 (N_30,In_162,In_946);
xor U31 (N_31,In_232,In_706);
or U32 (N_32,In_60,In_349);
nor U33 (N_33,In_257,In_328);
nand U34 (N_34,In_39,In_128);
or U35 (N_35,In_37,In_653);
and U36 (N_36,In_307,In_893);
or U37 (N_37,In_837,In_703);
nand U38 (N_38,In_270,In_416);
and U39 (N_39,In_898,In_389);
and U40 (N_40,In_354,In_731);
and U41 (N_41,In_634,In_467);
or U42 (N_42,In_482,In_497);
or U43 (N_43,In_192,In_194);
nor U44 (N_44,In_377,In_637);
nand U45 (N_45,In_992,In_963);
xor U46 (N_46,In_444,In_197);
and U47 (N_47,In_741,In_333);
nor U48 (N_48,In_331,In_662);
or U49 (N_49,In_205,In_478);
or U50 (N_50,In_261,In_29);
and U51 (N_51,In_819,In_529);
or U52 (N_52,In_110,In_248);
nor U53 (N_53,In_423,In_442);
or U54 (N_54,In_351,In_820);
nor U55 (N_55,In_508,In_635);
nor U56 (N_56,In_595,In_810);
nor U57 (N_57,In_338,In_334);
nand U58 (N_58,In_817,In_164);
nor U59 (N_59,In_66,In_484);
and U60 (N_60,In_507,In_462);
and U61 (N_61,In_322,In_666);
and U62 (N_62,In_96,In_249);
nor U63 (N_63,In_694,In_808);
nand U64 (N_64,In_888,In_774);
or U65 (N_65,In_346,In_884);
and U66 (N_66,In_614,In_915);
and U67 (N_67,In_557,In_121);
or U68 (N_68,In_234,In_564);
or U69 (N_69,In_101,In_81);
and U70 (N_70,In_350,In_572);
nand U71 (N_71,In_278,In_387);
nor U72 (N_72,In_277,In_450);
and U73 (N_73,In_840,In_437);
nand U74 (N_74,In_826,In_760);
or U75 (N_75,In_594,In_811);
nor U76 (N_76,In_347,In_996);
and U77 (N_77,In_567,In_618);
and U78 (N_78,In_142,In_670);
and U79 (N_79,In_525,In_610);
or U80 (N_80,In_861,In_199);
or U81 (N_81,In_698,In_7);
and U82 (N_82,In_493,In_70);
nand U83 (N_83,In_830,In_624);
or U84 (N_84,In_486,In_693);
or U85 (N_85,In_873,In_987);
nand U86 (N_86,In_537,In_552);
nor U87 (N_87,In_373,In_630);
nand U88 (N_88,In_988,In_803);
nand U89 (N_89,In_161,In_882);
or U90 (N_90,In_593,In_296);
or U91 (N_91,In_616,In_768);
xor U92 (N_92,In_118,In_747);
and U93 (N_93,In_558,In_742);
nor U94 (N_94,In_217,In_713);
nor U95 (N_95,In_83,In_880);
and U96 (N_96,In_879,In_405);
nand U97 (N_97,In_325,In_802);
nor U98 (N_98,In_584,In_272);
and U99 (N_99,In_87,In_263);
or U100 (N_100,In_541,In_718);
and U101 (N_101,In_986,In_288);
nand U102 (N_102,In_180,In_611);
nand U103 (N_103,In_209,In_74);
or U104 (N_104,In_907,In_33);
nor U105 (N_105,In_201,In_800);
or U106 (N_106,In_782,In_429);
or U107 (N_107,In_448,In_492);
nand U108 (N_108,In_835,In_92);
and U109 (N_109,In_48,In_677);
nor U110 (N_110,In_227,In_571);
or U111 (N_111,In_443,In_968);
or U112 (N_112,In_606,In_554);
or U113 (N_113,In_17,In_721);
or U114 (N_114,In_723,In_392);
and U115 (N_115,In_141,In_560);
or U116 (N_116,In_176,In_178);
xnor U117 (N_117,In_870,In_816);
or U118 (N_118,In_159,In_902);
nand U119 (N_119,In_645,In_765);
and U120 (N_120,In_852,In_379);
and U121 (N_121,In_526,In_867);
and U122 (N_122,In_924,In_366);
and U123 (N_123,In_961,In_146);
or U124 (N_124,In_476,In_642);
or U125 (N_125,In_682,In_651);
or U126 (N_126,In_626,In_211);
and U127 (N_127,In_983,In_853);
and U128 (N_128,In_381,In_166);
nor U129 (N_129,In_190,In_275);
or U130 (N_130,In_568,In_937);
nor U131 (N_131,In_388,In_623);
and U132 (N_132,In_220,In_652);
or U133 (N_133,In_581,In_431);
nor U134 (N_134,In_369,In_675);
and U135 (N_135,In_324,In_397);
nor U136 (N_136,In_244,In_754);
and U137 (N_137,In_5,In_40);
nor U138 (N_138,In_63,In_761);
and U139 (N_139,In_399,In_579);
nor U140 (N_140,In_485,In_510);
or U141 (N_141,In_72,In_701);
or U142 (N_142,In_470,In_258);
and U143 (N_143,In_503,In_518);
or U144 (N_144,In_749,In_965);
nand U145 (N_145,In_789,In_213);
nand U146 (N_146,In_231,In_43);
and U147 (N_147,In_999,In_191);
nor U148 (N_148,In_780,In_791);
nor U149 (N_149,In_805,In_422);
nor U150 (N_150,In_597,In_868);
and U151 (N_151,In_301,In_950);
or U152 (N_152,In_342,In_382);
nand U153 (N_153,In_664,In_866);
nand U154 (N_154,In_535,In_32);
or U155 (N_155,In_297,In_692);
or U156 (N_156,In_974,In_858);
nand U157 (N_157,In_984,In_864);
nor U158 (N_158,In_465,In_973);
and U159 (N_159,In_219,In_62);
nor U160 (N_160,In_851,In_772);
nand U161 (N_161,In_951,In_299);
nand U162 (N_162,In_886,In_436);
and U163 (N_163,In_73,In_994);
or U164 (N_164,In_336,In_726);
and U165 (N_165,In_940,In_26);
nor U166 (N_166,In_80,In_939);
nand U167 (N_167,In_620,In_942);
and U168 (N_168,In_287,In_315);
or U169 (N_169,In_343,In_909);
and U170 (N_170,In_419,In_463);
xor U171 (N_171,In_49,In_490);
or U172 (N_172,In_345,In_599);
nor U173 (N_173,In_639,In_11);
xor U174 (N_174,In_376,In_1);
nand U175 (N_175,In_250,In_914);
nor U176 (N_176,In_441,In_547);
and U177 (N_177,In_41,In_31);
nand U178 (N_178,In_900,In_913);
nand U179 (N_179,In_582,In_67);
and U180 (N_180,In_794,In_472);
nor U181 (N_181,In_223,In_979);
nand U182 (N_182,In_293,In_970);
and U183 (N_183,In_955,In_519);
nor U184 (N_184,In_781,In_663);
and U185 (N_185,In_407,In_842);
nor U186 (N_186,In_414,In_18);
or U187 (N_187,In_938,In_545);
nor U188 (N_188,In_302,In_303);
and U189 (N_189,In_788,In_520);
nor U190 (N_190,In_468,In_759);
nor U191 (N_191,In_475,In_348);
nand U192 (N_192,In_932,In_544);
nand U193 (N_193,In_35,In_575);
nor U194 (N_194,In_200,In_286);
or U195 (N_195,In_276,In_55);
and U196 (N_196,In_615,In_269);
or U197 (N_197,In_776,In_352);
or U198 (N_198,In_592,In_69);
nand U199 (N_199,In_638,In_154);
and U200 (N_200,In_832,In_733);
or U201 (N_201,In_739,In_995);
or U202 (N_202,In_107,In_921);
or U203 (N_203,In_453,In_136);
nor U204 (N_204,In_402,In_583);
or U205 (N_205,In_56,In_580);
nand U206 (N_206,In_513,In_869);
nor U207 (N_207,In_871,In_167);
nand U208 (N_208,In_910,In_237);
and U209 (N_209,In_536,In_729);
or U210 (N_210,In_145,In_736);
and U211 (N_211,In_551,In_256);
nor U212 (N_212,In_326,In_114);
or U213 (N_213,In_889,In_44);
or U214 (N_214,In_173,In_783);
and U215 (N_215,In_341,In_367);
nor U216 (N_216,In_291,In_848);
and U217 (N_217,In_312,In_38);
nand U218 (N_218,In_822,In_762);
nor U219 (N_219,In_813,In_152);
and U220 (N_220,In_596,In_430);
nor U221 (N_221,In_403,In_51);
or U222 (N_222,In_933,In_737);
xor U223 (N_223,In_374,In_59);
or U224 (N_224,In_412,In_978);
and U225 (N_225,In_836,In_155);
nand U226 (N_226,In_240,In_236);
nand U227 (N_227,In_10,In_673);
and U228 (N_228,In_93,In_515);
or U229 (N_229,In_941,In_829);
nand U230 (N_230,In_847,In_918);
or U231 (N_231,In_282,In_24);
nand U232 (N_232,In_559,In_50);
nand U233 (N_233,In_183,In_763);
and U234 (N_234,In_604,In_27);
nand U235 (N_235,In_831,In_576);
nand U236 (N_236,In_119,In_420);
or U237 (N_237,In_516,In_90);
nand U238 (N_238,In_455,In_268);
and U239 (N_239,In_945,In_289);
nor U240 (N_240,In_855,In_976);
or U241 (N_241,In_149,In_753);
and U242 (N_242,In_658,In_578);
or U243 (N_243,In_496,In_757);
or U244 (N_244,In_716,In_137);
nand U245 (N_245,In_679,In_151);
or U246 (N_246,In_944,In_766);
nand U247 (N_247,In_993,In_125);
nand U248 (N_248,In_158,In_202);
and U249 (N_249,In_501,In_449);
or U250 (N_250,In_329,In_517);
nor U251 (N_251,In_702,In_483);
and U252 (N_252,In_171,In_566);
nand U253 (N_253,In_375,In_491);
nand U254 (N_254,In_896,In_435);
nor U255 (N_255,In_498,In_253);
and U256 (N_256,In_647,In_359);
or U257 (N_257,In_424,In_916);
nor U258 (N_258,In_265,In_827);
nand U259 (N_259,In_758,In_587);
or U260 (N_260,In_4,In_505);
and U261 (N_261,In_147,In_14);
or U262 (N_262,In_953,In_935);
or U263 (N_263,In_428,In_215);
or U264 (N_264,In_744,In_458);
nor U265 (N_265,In_184,In_46);
and U266 (N_266,In_506,In_94);
nand U267 (N_267,In_260,In_862);
and U268 (N_268,In_923,In_335);
nand U269 (N_269,In_665,In_370);
and U270 (N_270,In_64,In_75);
nor U271 (N_271,In_193,In_327);
or U272 (N_272,In_457,In_977);
nor U273 (N_273,In_310,In_971);
nor U274 (N_274,In_674,In_714);
or U275 (N_275,In_875,In_401);
nand U276 (N_276,In_99,In_306);
and U277 (N_277,In_332,In_393);
nand U278 (N_278,In_903,In_115);
nand U279 (N_279,In_495,In_607);
nor U280 (N_280,In_13,In_704);
or U281 (N_281,In_686,In_12);
nor U282 (N_282,In_127,In_446);
nor U283 (N_283,In_730,In_23);
nand U284 (N_284,In_105,In_109);
and U285 (N_285,In_169,In_655);
and U286 (N_286,In_504,In_168);
nor U287 (N_287,In_644,In_464);
nor U288 (N_288,In_522,In_111);
and U289 (N_289,In_793,In_206);
nand U290 (N_290,In_710,In_372);
nand U291 (N_291,In_725,In_640);
and U292 (N_292,In_216,In_627);
or U293 (N_293,In_434,In_313);
and U294 (N_294,In_52,In_553);
or U295 (N_295,In_735,In_844);
and U296 (N_296,In_812,In_588);
or U297 (N_297,In_724,In_130);
nand U298 (N_298,In_132,In_691);
nor U299 (N_299,In_678,In_418);
or U300 (N_300,In_391,In_58);
nor U301 (N_301,In_380,In_309);
xnor U302 (N_302,In_960,In_972);
and U303 (N_303,In_204,In_809);
nor U304 (N_304,In_885,In_748);
and U305 (N_305,In_316,In_660);
or U306 (N_306,In_779,In_148);
and U307 (N_307,In_531,In_195);
xor U308 (N_308,In_887,In_815);
nor U309 (N_309,In_512,In_487);
and U310 (N_310,In_86,In_989);
or U311 (N_311,In_943,In_680);
nand U312 (N_312,In_912,In_591);
and U313 (N_313,In_841,In_9);
nand U314 (N_314,In_489,In_421);
nor U315 (N_315,In_262,In_36);
and U316 (N_316,In_68,In_689);
xnor U317 (N_317,In_612,In_411);
or U318 (N_318,In_460,In_823);
nor U319 (N_319,In_337,In_6);
nand U320 (N_320,In_524,In_8);
and U321 (N_321,In_969,In_0);
nor U322 (N_322,In_106,In_947);
and U323 (N_323,In_755,In_991);
nor U324 (N_324,In_967,In_771);
nor U325 (N_325,In_922,In_292);
and U326 (N_326,In_573,In_561);
and U327 (N_327,In_927,In_356);
and U328 (N_328,In_112,In_471);
nand U329 (N_329,In_585,In_532);
and U330 (N_330,In_267,In_534);
or U331 (N_331,In_636,In_318);
or U332 (N_332,In_628,In_229);
and U333 (N_333,In_165,In_91);
nor U334 (N_334,In_459,In_857);
or U335 (N_335,In_617,In_764);
nor U336 (N_336,In_222,In_926);
or U337 (N_337,In_980,In_494);
nor U338 (N_338,In_905,In_65);
nor U339 (N_339,In_806,In_892);
nor U340 (N_340,In_872,In_440);
nor U341 (N_341,In_542,In_308);
or U342 (N_342,In_883,In_384);
nor U343 (N_343,In_648,In_140);
or U344 (N_344,In_321,In_15);
nand U345 (N_345,In_839,In_603);
nand U346 (N_346,In_952,In_368);
and U347 (N_347,In_371,In_283);
and U348 (N_348,In_622,In_188);
nand U349 (N_349,In_717,In_97);
nand U350 (N_350,In_804,In_856);
or U351 (N_351,In_708,In_221);
nor U352 (N_352,In_461,In_84);
nand U353 (N_353,In_172,In_562);
or U354 (N_354,In_353,In_543);
and U355 (N_355,In_386,In_527);
or U356 (N_356,In_271,In_357);
or U357 (N_357,In_317,In_957);
and U358 (N_358,In_116,In_745);
nor U359 (N_359,In_122,In_254);
xor U360 (N_360,In_891,In_71);
xor U361 (N_361,In_711,In_734);
or U362 (N_362,In_574,In_383);
or U363 (N_363,In_452,In_709);
nand U364 (N_364,In_242,In_123);
and U365 (N_365,In_245,In_19);
nor U366 (N_366,In_966,In_683);
or U367 (N_367,In_395,In_931);
nor U368 (N_368,In_47,In_330);
or U369 (N_369,In_466,In_934);
and U370 (N_370,In_88,In_904);
and U371 (N_371,In_187,In_656);
nand U372 (N_372,In_144,In_563);
and U373 (N_373,In_228,In_134);
nand U374 (N_374,In_865,In_845);
and U375 (N_375,In_259,In_801);
nor U376 (N_376,In_246,In_138);
nor U377 (N_377,In_225,In_182);
or U378 (N_378,In_833,In_157);
nand U379 (N_379,In_920,In_825);
nor U380 (N_380,In_850,In_433);
nor U381 (N_381,In_394,In_181);
nand U382 (N_382,In_751,In_133);
or U383 (N_383,In_929,In_954);
nor U384 (N_384,In_672,In_45);
or U385 (N_385,In_160,In_224);
or U386 (N_386,In_778,In_319);
nand U387 (N_387,In_266,In_378);
or U388 (N_388,In_488,In_632);
xnor U389 (N_389,In_814,In_669);
nand U390 (N_390,In_117,In_208);
nand U391 (N_391,In_156,In_641);
nand U392 (N_392,In_894,In_451);
and U393 (N_393,In_828,In_602);
or U394 (N_394,In_767,In_807);
and U395 (N_395,In_415,In_340);
nand U396 (N_396,In_539,In_700);
or U397 (N_397,In_659,In_676);
nand U398 (N_398,In_124,In_671);
or U399 (N_399,In_792,In_426);
nand U400 (N_400,In_629,In_846);
and U401 (N_401,In_521,In_363);
or U402 (N_402,In_773,In_280);
nor U403 (N_403,In_42,In_480);
or U404 (N_404,In_473,In_2);
nor U405 (N_405,In_688,In_207);
nor U406 (N_406,In_170,In_684);
and U407 (N_407,In_390,In_243);
and U408 (N_408,In_153,In_481);
or U409 (N_409,In_78,In_404);
or U410 (N_410,In_601,In_281);
or U411 (N_411,In_685,In_985);
and U412 (N_412,In_727,In_936);
and U413 (N_413,In_752,In_108);
nor U414 (N_414,In_570,In_235);
nor U415 (N_415,In_82,In_997);
and U416 (N_416,In_203,In_777);
or U417 (N_417,In_163,In_613);
nand U418 (N_418,In_439,In_362);
nand U419 (N_419,In_54,In_241);
or U420 (N_420,In_746,In_212);
or U421 (N_421,In_975,In_590);
or U422 (N_422,In_150,In_930);
or U423 (N_423,In_264,In_720);
or U424 (N_424,In_608,In_398);
nand U425 (N_425,In_854,In_214);
nand U426 (N_426,In_728,In_251);
nor U427 (N_427,In_890,In_548);
xnor U428 (N_428,In_824,In_477);
nor U429 (N_429,In_690,In_28);
or U430 (N_430,In_22,In_897);
nor U431 (N_431,In_775,In_252);
nand U432 (N_432,In_540,In_98);
nand U433 (N_433,In_131,In_300);
and U434 (N_434,In_135,In_314);
or U435 (N_435,In_838,In_210);
or U436 (N_436,In_998,In_445);
or U437 (N_437,In_454,In_320);
nor U438 (N_438,In_406,In_425);
and U439 (N_439,In_928,In_738);
nor U440 (N_440,In_821,In_586);
and U441 (N_441,In_538,In_770);
and U442 (N_442,In_722,In_239);
nor U443 (N_443,In_396,In_917);
nand U444 (N_444,In_732,In_57);
nand U445 (N_445,In_102,In_189);
xor U446 (N_446,In_16,In_500);
nor U447 (N_447,In_631,In_61);
nand U448 (N_448,In_179,In_95);
or U449 (N_449,In_34,In_740);
and U450 (N_450,In_797,In_355);
nand U451 (N_451,In_661,In_956);
nor U452 (N_452,In_304,In_233);
nor U453 (N_453,In_100,In_609);
nor U454 (N_454,In_364,In_859);
and U455 (N_455,In_874,In_818);
nand U456 (N_456,In_528,In_697);
and U457 (N_457,In_226,In_305);
nand U458 (N_458,In_408,In_795);
or U459 (N_459,In_687,In_901);
and U460 (N_460,In_598,In_344);
and U461 (N_461,In_719,In_139);
or U462 (N_462,In_427,In_643);
nor U463 (N_463,In_863,In_705);
nand U464 (N_464,In_696,In_410);
nand U465 (N_465,In_479,In_769);
and U466 (N_466,In_964,In_949);
nor U467 (N_467,In_786,In_546);
xor U468 (N_468,In_502,In_533);
nor U469 (N_469,In_982,In_785);
nand U470 (N_470,In_365,In_877);
or U471 (N_471,In_619,In_654);
or U472 (N_472,In_798,In_400);
nor U473 (N_473,In_549,In_279);
or U474 (N_474,In_881,In_530);
or U475 (N_475,In_657,In_89);
or U476 (N_476,In_876,In_895);
nor U477 (N_477,In_668,In_447);
nand U478 (N_478,In_238,In_784);
and U479 (N_479,In_432,In_948);
or U480 (N_480,In_555,In_76);
nand U481 (N_481,In_600,In_919);
and U482 (N_482,In_25,In_218);
or U483 (N_483,In_20,In_284);
and U484 (N_484,In_509,In_126);
nor U485 (N_485,In_474,In_186);
and U486 (N_486,In_796,In_104);
or U487 (N_487,In_646,In_129);
nor U488 (N_488,In_361,In_649);
nand U489 (N_489,In_799,In_3);
and U490 (N_490,In_177,In_790);
and U491 (N_491,In_707,In_103);
or U492 (N_492,In_417,In_120);
xor U493 (N_493,In_469,In_621);
or U494 (N_494,In_911,In_605);
nor U495 (N_495,In_787,In_358);
nand U496 (N_496,In_681,In_650);
or U497 (N_497,In_290,In_511);
nor U498 (N_498,In_899,In_556);
nor U499 (N_499,In_550,In_906);
and U500 (N_500,In_108,In_874);
and U501 (N_501,In_245,In_318);
nor U502 (N_502,In_917,In_549);
or U503 (N_503,In_43,In_157);
and U504 (N_504,In_422,In_91);
or U505 (N_505,In_840,In_112);
nand U506 (N_506,In_588,In_226);
or U507 (N_507,In_878,In_620);
or U508 (N_508,In_93,In_690);
and U509 (N_509,In_981,In_150);
and U510 (N_510,In_450,In_599);
nor U511 (N_511,In_681,In_830);
nor U512 (N_512,In_303,In_544);
nor U513 (N_513,In_325,In_240);
or U514 (N_514,In_14,In_906);
and U515 (N_515,In_130,In_934);
and U516 (N_516,In_447,In_242);
or U517 (N_517,In_905,In_698);
or U518 (N_518,In_515,In_798);
nand U519 (N_519,In_677,In_59);
nor U520 (N_520,In_840,In_226);
nor U521 (N_521,In_141,In_380);
and U522 (N_522,In_624,In_458);
nand U523 (N_523,In_337,In_93);
and U524 (N_524,In_101,In_564);
nor U525 (N_525,In_119,In_647);
and U526 (N_526,In_225,In_412);
or U527 (N_527,In_958,In_892);
and U528 (N_528,In_618,In_150);
and U529 (N_529,In_881,In_358);
and U530 (N_530,In_215,In_423);
nand U531 (N_531,In_897,In_799);
xnor U532 (N_532,In_992,In_160);
xnor U533 (N_533,In_431,In_362);
and U534 (N_534,In_672,In_538);
and U535 (N_535,In_903,In_121);
nand U536 (N_536,In_81,In_209);
nor U537 (N_537,In_426,In_731);
or U538 (N_538,In_53,In_63);
nand U539 (N_539,In_750,In_220);
or U540 (N_540,In_254,In_127);
nor U541 (N_541,In_255,In_882);
or U542 (N_542,In_772,In_253);
nor U543 (N_543,In_121,In_366);
and U544 (N_544,In_762,In_182);
xnor U545 (N_545,In_163,In_154);
and U546 (N_546,In_61,In_151);
and U547 (N_547,In_75,In_183);
and U548 (N_548,In_914,In_600);
nor U549 (N_549,In_554,In_429);
xor U550 (N_550,In_418,In_180);
nor U551 (N_551,In_548,In_673);
and U552 (N_552,In_851,In_927);
and U553 (N_553,In_597,In_968);
nand U554 (N_554,In_578,In_903);
and U555 (N_555,In_238,In_484);
nor U556 (N_556,In_26,In_135);
and U557 (N_557,In_204,In_387);
nand U558 (N_558,In_905,In_128);
nand U559 (N_559,In_720,In_746);
nand U560 (N_560,In_838,In_590);
and U561 (N_561,In_153,In_183);
nand U562 (N_562,In_566,In_658);
nand U563 (N_563,In_563,In_968);
nor U564 (N_564,In_687,In_103);
nor U565 (N_565,In_972,In_767);
nor U566 (N_566,In_962,In_824);
and U567 (N_567,In_927,In_894);
xnor U568 (N_568,In_475,In_176);
or U569 (N_569,In_542,In_102);
and U570 (N_570,In_697,In_257);
xor U571 (N_571,In_316,In_616);
nor U572 (N_572,In_987,In_973);
and U573 (N_573,In_678,In_819);
and U574 (N_574,In_307,In_18);
xor U575 (N_575,In_974,In_573);
nand U576 (N_576,In_339,In_648);
and U577 (N_577,In_219,In_17);
nor U578 (N_578,In_145,In_839);
nor U579 (N_579,In_695,In_577);
nand U580 (N_580,In_279,In_410);
nor U581 (N_581,In_227,In_164);
or U582 (N_582,In_998,In_503);
nor U583 (N_583,In_441,In_193);
nand U584 (N_584,In_550,In_24);
nor U585 (N_585,In_954,In_458);
nand U586 (N_586,In_139,In_837);
nand U587 (N_587,In_911,In_362);
nor U588 (N_588,In_317,In_391);
nor U589 (N_589,In_807,In_389);
and U590 (N_590,In_39,In_684);
nand U591 (N_591,In_57,In_825);
or U592 (N_592,In_792,In_47);
or U593 (N_593,In_225,In_757);
or U594 (N_594,In_566,In_77);
nand U595 (N_595,In_471,In_710);
nor U596 (N_596,In_935,In_813);
or U597 (N_597,In_479,In_185);
nor U598 (N_598,In_111,In_371);
nor U599 (N_599,In_143,In_133);
and U600 (N_600,In_943,In_389);
or U601 (N_601,In_735,In_665);
nand U602 (N_602,In_34,In_119);
nand U603 (N_603,In_308,In_392);
nor U604 (N_604,In_461,In_292);
nor U605 (N_605,In_131,In_46);
nor U606 (N_606,In_667,In_370);
nor U607 (N_607,In_659,In_181);
or U608 (N_608,In_996,In_213);
nor U609 (N_609,In_131,In_261);
nor U610 (N_610,In_862,In_76);
nand U611 (N_611,In_279,In_239);
and U612 (N_612,In_23,In_895);
nand U613 (N_613,In_748,In_389);
nand U614 (N_614,In_941,In_574);
or U615 (N_615,In_723,In_214);
nand U616 (N_616,In_629,In_258);
nor U617 (N_617,In_677,In_941);
nor U618 (N_618,In_845,In_742);
or U619 (N_619,In_232,In_568);
or U620 (N_620,In_946,In_852);
and U621 (N_621,In_15,In_827);
and U622 (N_622,In_219,In_814);
nand U623 (N_623,In_515,In_164);
nand U624 (N_624,In_265,In_78);
xor U625 (N_625,In_254,In_772);
nand U626 (N_626,In_968,In_734);
and U627 (N_627,In_723,In_324);
nand U628 (N_628,In_208,In_488);
nand U629 (N_629,In_874,In_506);
or U630 (N_630,In_168,In_441);
nor U631 (N_631,In_571,In_239);
nor U632 (N_632,In_853,In_474);
or U633 (N_633,In_412,In_545);
and U634 (N_634,In_747,In_863);
and U635 (N_635,In_34,In_434);
nand U636 (N_636,In_19,In_994);
xor U637 (N_637,In_820,In_684);
nor U638 (N_638,In_325,In_244);
nand U639 (N_639,In_494,In_839);
and U640 (N_640,In_164,In_183);
and U641 (N_641,In_873,In_588);
nand U642 (N_642,In_843,In_397);
nor U643 (N_643,In_667,In_453);
nand U644 (N_644,In_645,In_223);
nand U645 (N_645,In_818,In_61);
nor U646 (N_646,In_809,In_616);
nand U647 (N_647,In_928,In_71);
nand U648 (N_648,In_882,In_130);
nand U649 (N_649,In_843,In_151);
nand U650 (N_650,In_941,In_631);
nand U651 (N_651,In_456,In_164);
or U652 (N_652,In_212,In_529);
nand U653 (N_653,In_909,In_870);
nand U654 (N_654,In_234,In_801);
nor U655 (N_655,In_854,In_198);
nand U656 (N_656,In_964,In_937);
nand U657 (N_657,In_392,In_748);
nor U658 (N_658,In_718,In_528);
nand U659 (N_659,In_490,In_479);
nand U660 (N_660,In_408,In_973);
and U661 (N_661,In_927,In_410);
or U662 (N_662,In_642,In_412);
nand U663 (N_663,In_613,In_269);
and U664 (N_664,In_577,In_388);
and U665 (N_665,In_588,In_558);
and U666 (N_666,In_706,In_570);
or U667 (N_667,In_553,In_838);
xnor U668 (N_668,In_313,In_795);
or U669 (N_669,In_497,In_843);
nor U670 (N_670,In_175,In_453);
or U671 (N_671,In_243,In_80);
xor U672 (N_672,In_498,In_949);
nand U673 (N_673,In_826,In_230);
or U674 (N_674,In_581,In_775);
and U675 (N_675,In_902,In_885);
and U676 (N_676,In_149,In_835);
or U677 (N_677,In_666,In_427);
and U678 (N_678,In_3,In_590);
or U679 (N_679,In_786,In_533);
xnor U680 (N_680,In_142,In_563);
or U681 (N_681,In_689,In_279);
and U682 (N_682,In_805,In_494);
or U683 (N_683,In_619,In_412);
nor U684 (N_684,In_507,In_198);
nand U685 (N_685,In_338,In_11);
nand U686 (N_686,In_700,In_706);
and U687 (N_687,In_540,In_977);
nand U688 (N_688,In_34,In_818);
nor U689 (N_689,In_28,In_541);
nand U690 (N_690,In_880,In_978);
nand U691 (N_691,In_318,In_601);
nand U692 (N_692,In_214,In_104);
and U693 (N_693,In_841,In_627);
nor U694 (N_694,In_508,In_72);
and U695 (N_695,In_830,In_984);
nor U696 (N_696,In_995,In_737);
and U697 (N_697,In_909,In_335);
nor U698 (N_698,In_304,In_248);
and U699 (N_699,In_598,In_270);
xnor U700 (N_700,In_135,In_184);
nand U701 (N_701,In_371,In_515);
nor U702 (N_702,In_268,In_251);
nor U703 (N_703,In_607,In_767);
nor U704 (N_704,In_117,In_742);
or U705 (N_705,In_28,In_89);
nor U706 (N_706,In_728,In_888);
nor U707 (N_707,In_181,In_168);
and U708 (N_708,In_448,In_653);
nor U709 (N_709,In_158,In_38);
or U710 (N_710,In_832,In_663);
nor U711 (N_711,In_105,In_467);
or U712 (N_712,In_235,In_263);
and U713 (N_713,In_776,In_484);
or U714 (N_714,In_753,In_266);
or U715 (N_715,In_806,In_620);
or U716 (N_716,In_636,In_406);
or U717 (N_717,In_13,In_161);
or U718 (N_718,In_984,In_820);
or U719 (N_719,In_651,In_831);
and U720 (N_720,In_624,In_916);
and U721 (N_721,In_485,In_19);
or U722 (N_722,In_749,In_747);
or U723 (N_723,In_430,In_138);
nand U724 (N_724,In_914,In_920);
and U725 (N_725,In_856,In_267);
nor U726 (N_726,In_695,In_793);
nand U727 (N_727,In_574,In_650);
nand U728 (N_728,In_43,In_194);
nand U729 (N_729,In_325,In_456);
nand U730 (N_730,In_638,In_528);
or U731 (N_731,In_292,In_351);
and U732 (N_732,In_813,In_402);
nor U733 (N_733,In_101,In_710);
nor U734 (N_734,In_346,In_294);
nor U735 (N_735,In_246,In_385);
nand U736 (N_736,In_958,In_559);
or U737 (N_737,In_73,In_887);
or U738 (N_738,In_950,In_633);
xor U739 (N_739,In_183,In_102);
nand U740 (N_740,In_230,In_688);
nand U741 (N_741,In_834,In_568);
or U742 (N_742,In_239,In_181);
and U743 (N_743,In_113,In_165);
and U744 (N_744,In_330,In_704);
and U745 (N_745,In_69,In_752);
or U746 (N_746,In_529,In_857);
or U747 (N_747,In_881,In_953);
or U748 (N_748,In_686,In_77);
and U749 (N_749,In_386,In_547);
xor U750 (N_750,In_148,In_543);
or U751 (N_751,In_790,In_198);
or U752 (N_752,In_155,In_954);
nor U753 (N_753,In_574,In_541);
or U754 (N_754,In_368,In_220);
nor U755 (N_755,In_420,In_792);
and U756 (N_756,In_812,In_387);
and U757 (N_757,In_108,In_436);
nand U758 (N_758,In_523,In_587);
xor U759 (N_759,In_301,In_497);
and U760 (N_760,In_576,In_821);
or U761 (N_761,In_186,In_198);
or U762 (N_762,In_128,In_361);
nand U763 (N_763,In_33,In_45);
nand U764 (N_764,In_107,In_123);
nand U765 (N_765,In_236,In_937);
and U766 (N_766,In_901,In_361);
nand U767 (N_767,In_625,In_922);
or U768 (N_768,In_5,In_222);
and U769 (N_769,In_203,In_858);
and U770 (N_770,In_276,In_204);
and U771 (N_771,In_343,In_799);
nand U772 (N_772,In_769,In_30);
nor U773 (N_773,In_870,In_193);
nor U774 (N_774,In_820,In_437);
nand U775 (N_775,In_287,In_278);
and U776 (N_776,In_90,In_647);
or U777 (N_777,In_577,In_231);
nor U778 (N_778,In_494,In_45);
and U779 (N_779,In_412,In_990);
nand U780 (N_780,In_78,In_399);
nor U781 (N_781,In_64,In_708);
or U782 (N_782,In_412,In_631);
nor U783 (N_783,In_551,In_264);
and U784 (N_784,In_978,In_552);
nand U785 (N_785,In_569,In_58);
and U786 (N_786,In_237,In_146);
nor U787 (N_787,In_554,In_490);
or U788 (N_788,In_490,In_422);
and U789 (N_789,In_56,In_793);
and U790 (N_790,In_838,In_623);
and U791 (N_791,In_862,In_218);
nor U792 (N_792,In_848,In_354);
xor U793 (N_793,In_802,In_519);
or U794 (N_794,In_931,In_280);
nor U795 (N_795,In_772,In_297);
nor U796 (N_796,In_729,In_572);
nor U797 (N_797,In_890,In_544);
nor U798 (N_798,In_596,In_234);
nor U799 (N_799,In_889,In_337);
and U800 (N_800,In_116,In_506);
nor U801 (N_801,In_643,In_784);
or U802 (N_802,In_39,In_191);
or U803 (N_803,In_17,In_403);
or U804 (N_804,In_402,In_906);
or U805 (N_805,In_58,In_258);
and U806 (N_806,In_227,In_588);
and U807 (N_807,In_193,In_688);
nor U808 (N_808,In_859,In_304);
and U809 (N_809,In_599,In_558);
nand U810 (N_810,In_458,In_857);
nor U811 (N_811,In_487,In_343);
nand U812 (N_812,In_631,In_188);
and U813 (N_813,In_393,In_303);
or U814 (N_814,In_65,In_807);
nand U815 (N_815,In_480,In_640);
nand U816 (N_816,In_391,In_686);
nor U817 (N_817,In_976,In_856);
and U818 (N_818,In_630,In_260);
nand U819 (N_819,In_440,In_569);
nor U820 (N_820,In_828,In_487);
xor U821 (N_821,In_360,In_795);
and U822 (N_822,In_854,In_425);
nor U823 (N_823,In_562,In_421);
and U824 (N_824,In_699,In_446);
nand U825 (N_825,In_369,In_819);
and U826 (N_826,In_825,In_531);
nor U827 (N_827,In_70,In_227);
nor U828 (N_828,In_17,In_958);
and U829 (N_829,In_348,In_901);
and U830 (N_830,In_465,In_417);
nand U831 (N_831,In_813,In_923);
nand U832 (N_832,In_952,In_278);
and U833 (N_833,In_63,In_468);
nor U834 (N_834,In_871,In_792);
and U835 (N_835,In_555,In_959);
and U836 (N_836,In_76,In_27);
nand U837 (N_837,In_364,In_190);
nand U838 (N_838,In_376,In_500);
nor U839 (N_839,In_586,In_771);
nand U840 (N_840,In_801,In_800);
nand U841 (N_841,In_712,In_469);
nand U842 (N_842,In_987,In_26);
nand U843 (N_843,In_870,In_207);
nor U844 (N_844,In_740,In_426);
nand U845 (N_845,In_607,In_806);
nor U846 (N_846,In_408,In_548);
nor U847 (N_847,In_580,In_908);
nand U848 (N_848,In_40,In_642);
nor U849 (N_849,In_585,In_464);
or U850 (N_850,In_467,In_183);
nand U851 (N_851,In_114,In_86);
and U852 (N_852,In_61,In_73);
nand U853 (N_853,In_498,In_802);
and U854 (N_854,In_812,In_638);
nand U855 (N_855,In_415,In_857);
nand U856 (N_856,In_83,In_983);
or U857 (N_857,In_613,In_596);
or U858 (N_858,In_364,In_973);
nand U859 (N_859,In_671,In_395);
and U860 (N_860,In_231,In_238);
and U861 (N_861,In_616,In_47);
nor U862 (N_862,In_312,In_675);
nand U863 (N_863,In_648,In_546);
or U864 (N_864,In_960,In_929);
and U865 (N_865,In_143,In_0);
or U866 (N_866,In_574,In_739);
or U867 (N_867,In_764,In_469);
or U868 (N_868,In_627,In_416);
and U869 (N_869,In_903,In_880);
nand U870 (N_870,In_505,In_599);
nor U871 (N_871,In_977,In_359);
nor U872 (N_872,In_472,In_5);
nand U873 (N_873,In_764,In_780);
or U874 (N_874,In_355,In_506);
or U875 (N_875,In_296,In_416);
nor U876 (N_876,In_247,In_34);
or U877 (N_877,In_360,In_985);
or U878 (N_878,In_255,In_47);
nor U879 (N_879,In_613,In_512);
nor U880 (N_880,In_165,In_615);
nand U881 (N_881,In_150,In_192);
nand U882 (N_882,In_169,In_400);
and U883 (N_883,In_716,In_23);
nand U884 (N_884,In_976,In_967);
xnor U885 (N_885,In_810,In_829);
and U886 (N_886,In_242,In_361);
nand U887 (N_887,In_680,In_69);
xor U888 (N_888,In_433,In_393);
xnor U889 (N_889,In_744,In_28);
or U890 (N_890,In_217,In_82);
and U891 (N_891,In_450,In_511);
nor U892 (N_892,In_135,In_885);
nand U893 (N_893,In_613,In_843);
or U894 (N_894,In_152,In_664);
nand U895 (N_895,In_785,In_117);
nor U896 (N_896,In_794,In_11);
nor U897 (N_897,In_294,In_639);
nor U898 (N_898,In_84,In_708);
nand U899 (N_899,In_686,In_259);
and U900 (N_900,In_611,In_330);
or U901 (N_901,In_235,In_917);
nor U902 (N_902,In_895,In_589);
nor U903 (N_903,In_378,In_291);
nand U904 (N_904,In_518,In_414);
nor U905 (N_905,In_948,In_852);
and U906 (N_906,In_999,In_520);
nor U907 (N_907,In_147,In_121);
and U908 (N_908,In_325,In_307);
nor U909 (N_909,In_703,In_622);
nor U910 (N_910,In_467,In_476);
nor U911 (N_911,In_98,In_50);
xnor U912 (N_912,In_96,In_596);
or U913 (N_913,In_666,In_901);
nor U914 (N_914,In_79,In_113);
and U915 (N_915,In_665,In_432);
nor U916 (N_916,In_851,In_963);
and U917 (N_917,In_683,In_162);
and U918 (N_918,In_497,In_173);
nor U919 (N_919,In_673,In_555);
or U920 (N_920,In_320,In_48);
nor U921 (N_921,In_78,In_863);
nor U922 (N_922,In_161,In_396);
nand U923 (N_923,In_852,In_252);
and U924 (N_924,In_804,In_632);
or U925 (N_925,In_649,In_562);
and U926 (N_926,In_349,In_812);
nor U927 (N_927,In_248,In_616);
nor U928 (N_928,In_329,In_393);
nor U929 (N_929,In_459,In_130);
nor U930 (N_930,In_758,In_804);
or U931 (N_931,In_550,In_991);
nor U932 (N_932,In_45,In_132);
or U933 (N_933,In_306,In_64);
or U934 (N_934,In_993,In_105);
nand U935 (N_935,In_257,In_816);
nor U936 (N_936,In_526,In_456);
or U937 (N_937,In_930,In_641);
and U938 (N_938,In_833,In_761);
nand U939 (N_939,In_569,In_107);
nor U940 (N_940,In_304,In_589);
nor U941 (N_941,In_693,In_482);
nor U942 (N_942,In_438,In_40);
nor U943 (N_943,In_793,In_781);
nor U944 (N_944,In_270,In_591);
and U945 (N_945,In_305,In_431);
nand U946 (N_946,In_230,In_21);
and U947 (N_947,In_35,In_174);
and U948 (N_948,In_951,In_427);
and U949 (N_949,In_764,In_553);
xnor U950 (N_950,In_253,In_569);
nor U951 (N_951,In_307,In_834);
nor U952 (N_952,In_796,In_157);
nand U953 (N_953,In_680,In_93);
nor U954 (N_954,In_413,In_55);
nand U955 (N_955,In_320,In_139);
and U956 (N_956,In_916,In_556);
nand U957 (N_957,In_65,In_598);
or U958 (N_958,In_927,In_533);
nand U959 (N_959,In_529,In_570);
nor U960 (N_960,In_878,In_315);
nand U961 (N_961,In_92,In_900);
and U962 (N_962,In_221,In_29);
nand U963 (N_963,In_711,In_811);
nand U964 (N_964,In_161,In_832);
nor U965 (N_965,In_757,In_673);
nor U966 (N_966,In_191,In_631);
nand U967 (N_967,In_121,In_717);
nor U968 (N_968,In_92,In_937);
xnor U969 (N_969,In_213,In_954);
nand U970 (N_970,In_980,In_295);
nand U971 (N_971,In_972,In_195);
nand U972 (N_972,In_608,In_549);
or U973 (N_973,In_468,In_890);
and U974 (N_974,In_693,In_452);
nor U975 (N_975,In_379,In_288);
nand U976 (N_976,In_919,In_909);
or U977 (N_977,In_361,In_794);
nand U978 (N_978,In_964,In_129);
nor U979 (N_979,In_94,In_96);
nand U980 (N_980,In_559,In_396);
or U981 (N_981,In_164,In_285);
nor U982 (N_982,In_560,In_863);
nor U983 (N_983,In_746,In_240);
nor U984 (N_984,In_124,In_270);
or U985 (N_985,In_977,In_614);
nor U986 (N_986,In_64,In_679);
or U987 (N_987,In_564,In_227);
nor U988 (N_988,In_383,In_316);
or U989 (N_989,In_257,In_108);
nor U990 (N_990,In_202,In_801);
nor U991 (N_991,In_366,In_14);
xnor U992 (N_992,In_258,In_526);
nor U993 (N_993,In_607,In_405);
or U994 (N_994,In_535,In_12);
and U995 (N_995,In_693,In_768);
and U996 (N_996,In_895,In_773);
nor U997 (N_997,In_660,In_800);
nor U998 (N_998,In_699,In_120);
nand U999 (N_999,In_796,In_736);
nand U1000 (N_1000,In_86,In_793);
or U1001 (N_1001,In_28,In_452);
or U1002 (N_1002,In_759,In_361);
or U1003 (N_1003,In_822,In_317);
or U1004 (N_1004,In_803,In_579);
nor U1005 (N_1005,In_524,In_1);
or U1006 (N_1006,In_765,In_161);
nor U1007 (N_1007,In_907,In_296);
or U1008 (N_1008,In_387,In_311);
nand U1009 (N_1009,In_274,In_65);
or U1010 (N_1010,In_320,In_42);
or U1011 (N_1011,In_184,In_638);
and U1012 (N_1012,In_170,In_644);
nand U1013 (N_1013,In_840,In_906);
and U1014 (N_1014,In_537,In_582);
nand U1015 (N_1015,In_585,In_66);
nor U1016 (N_1016,In_942,In_250);
and U1017 (N_1017,In_608,In_81);
nor U1018 (N_1018,In_743,In_700);
nor U1019 (N_1019,In_98,In_9);
and U1020 (N_1020,In_5,In_896);
or U1021 (N_1021,In_197,In_228);
nand U1022 (N_1022,In_88,In_724);
or U1023 (N_1023,In_23,In_382);
nor U1024 (N_1024,In_564,In_526);
and U1025 (N_1025,In_724,In_919);
and U1026 (N_1026,In_711,In_72);
nor U1027 (N_1027,In_616,In_258);
nor U1028 (N_1028,In_914,In_627);
nor U1029 (N_1029,In_77,In_929);
nand U1030 (N_1030,In_182,In_444);
or U1031 (N_1031,In_4,In_386);
nand U1032 (N_1032,In_36,In_659);
nand U1033 (N_1033,In_642,In_58);
or U1034 (N_1034,In_646,In_729);
nor U1035 (N_1035,In_976,In_862);
or U1036 (N_1036,In_472,In_111);
nand U1037 (N_1037,In_990,In_390);
and U1038 (N_1038,In_20,In_489);
nor U1039 (N_1039,In_166,In_870);
nand U1040 (N_1040,In_300,In_359);
or U1041 (N_1041,In_691,In_4);
nand U1042 (N_1042,In_835,In_834);
nor U1043 (N_1043,In_739,In_861);
and U1044 (N_1044,In_66,In_939);
nand U1045 (N_1045,In_532,In_961);
nand U1046 (N_1046,In_496,In_371);
nand U1047 (N_1047,In_56,In_414);
nor U1048 (N_1048,In_403,In_586);
nand U1049 (N_1049,In_520,In_36);
and U1050 (N_1050,In_825,In_628);
nor U1051 (N_1051,In_206,In_110);
and U1052 (N_1052,In_542,In_968);
or U1053 (N_1053,In_727,In_169);
nor U1054 (N_1054,In_629,In_954);
nand U1055 (N_1055,In_940,In_802);
nand U1056 (N_1056,In_125,In_605);
nor U1057 (N_1057,In_698,In_81);
or U1058 (N_1058,In_616,In_525);
and U1059 (N_1059,In_464,In_43);
nor U1060 (N_1060,In_861,In_412);
xor U1061 (N_1061,In_977,In_559);
or U1062 (N_1062,In_320,In_861);
nor U1063 (N_1063,In_397,In_46);
xnor U1064 (N_1064,In_814,In_712);
or U1065 (N_1065,In_695,In_492);
or U1066 (N_1066,In_873,In_730);
xor U1067 (N_1067,In_170,In_924);
nand U1068 (N_1068,In_996,In_547);
nor U1069 (N_1069,In_884,In_659);
nor U1070 (N_1070,In_737,In_289);
or U1071 (N_1071,In_99,In_704);
nor U1072 (N_1072,In_125,In_104);
xor U1073 (N_1073,In_772,In_416);
nor U1074 (N_1074,In_478,In_166);
and U1075 (N_1075,In_21,In_513);
and U1076 (N_1076,In_783,In_233);
nand U1077 (N_1077,In_560,In_328);
or U1078 (N_1078,In_249,In_778);
nand U1079 (N_1079,In_199,In_939);
or U1080 (N_1080,In_803,In_830);
or U1081 (N_1081,In_287,In_617);
or U1082 (N_1082,In_290,In_345);
xnor U1083 (N_1083,In_755,In_51);
or U1084 (N_1084,In_714,In_727);
or U1085 (N_1085,In_990,In_649);
nand U1086 (N_1086,In_996,In_450);
xor U1087 (N_1087,In_458,In_310);
and U1088 (N_1088,In_154,In_27);
nand U1089 (N_1089,In_111,In_660);
nor U1090 (N_1090,In_32,In_307);
or U1091 (N_1091,In_264,In_681);
or U1092 (N_1092,In_618,In_50);
nand U1093 (N_1093,In_894,In_377);
or U1094 (N_1094,In_763,In_456);
nand U1095 (N_1095,In_485,In_402);
or U1096 (N_1096,In_347,In_57);
nor U1097 (N_1097,In_879,In_196);
or U1098 (N_1098,In_167,In_805);
nor U1099 (N_1099,In_643,In_173);
nor U1100 (N_1100,In_91,In_378);
nor U1101 (N_1101,In_894,In_658);
nor U1102 (N_1102,In_678,In_720);
and U1103 (N_1103,In_769,In_104);
and U1104 (N_1104,In_464,In_19);
nor U1105 (N_1105,In_390,In_105);
and U1106 (N_1106,In_41,In_384);
and U1107 (N_1107,In_958,In_460);
and U1108 (N_1108,In_634,In_495);
and U1109 (N_1109,In_447,In_752);
nand U1110 (N_1110,In_518,In_46);
or U1111 (N_1111,In_684,In_124);
nor U1112 (N_1112,In_118,In_221);
nand U1113 (N_1113,In_215,In_603);
nand U1114 (N_1114,In_484,In_370);
xor U1115 (N_1115,In_330,In_96);
and U1116 (N_1116,In_442,In_518);
nand U1117 (N_1117,In_739,In_388);
nand U1118 (N_1118,In_567,In_96);
nand U1119 (N_1119,In_894,In_725);
nand U1120 (N_1120,In_859,In_316);
nand U1121 (N_1121,In_933,In_375);
or U1122 (N_1122,In_157,In_727);
nor U1123 (N_1123,In_903,In_646);
nand U1124 (N_1124,In_297,In_599);
or U1125 (N_1125,In_514,In_111);
and U1126 (N_1126,In_691,In_701);
and U1127 (N_1127,In_232,In_98);
or U1128 (N_1128,In_747,In_956);
xor U1129 (N_1129,In_202,In_591);
nand U1130 (N_1130,In_363,In_630);
nor U1131 (N_1131,In_897,In_777);
and U1132 (N_1132,In_745,In_533);
or U1133 (N_1133,In_634,In_146);
nand U1134 (N_1134,In_746,In_81);
and U1135 (N_1135,In_713,In_635);
nand U1136 (N_1136,In_668,In_479);
and U1137 (N_1137,In_472,In_85);
nor U1138 (N_1138,In_840,In_803);
nor U1139 (N_1139,In_593,In_568);
nor U1140 (N_1140,In_516,In_627);
nor U1141 (N_1141,In_699,In_380);
and U1142 (N_1142,In_844,In_228);
nor U1143 (N_1143,In_579,In_650);
and U1144 (N_1144,In_160,In_215);
and U1145 (N_1145,In_442,In_144);
nor U1146 (N_1146,In_732,In_930);
or U1147 (N_1147,In_222,In_26);
nand U1148 (N_1148,In_930,In_196);
nor U1149 (N_1149,In_362,In_246);
or U1150 (N_1150,In_597,In_404);
nand U1151 (N_1151,In_171,In_369);
nand U1152 (N_1152,In_97,In_224);
nor U1153 (N_1153,In_568,In_714);
nor U1154 (N_1154,In_702,In_611);
and U1155 (N_1155,In_746,In_988);
and U1156 (N_1156,In_629,In_744);
or U1157 (N_1157,In_615,In_176);
and U1158 (N_1158,In_232,In_827);
and U1159 (N_1159,In_272,In_671);
or U1160 (N_1160,In_906,In_565);
or U1161 (N_1161,In_443,In_232);
nand U1162 (N_1162,In_905,In_145);
and U1163 (N_1163,In_281,In_673);
nor U1164 (N_1164,In_130,In_428);
or U1165 (N_1165,In_703,In_594);
or U1166 (N_1166,In_411,In_942);
or U1167 (N_1167,In_9,In_411);
and U1168 (N_1168,In_309,In_438);
or U1169 (N_1169,In_166,In_620);
or U1170 (N_1170,In_52,In_101);
nand U1171 (N_1171,In_911,In_314);
or U1172 (N_1172,In_21,In_61);
nand U1173 (N_1173,In_799,In_217);
xor U1174 (N_1174,In_506,In_185);
nand U1175 (N_1175,In_189,In_50);
or U1176 (N_1176,In_657,In_440);
nor U1177 (N_1177,In_748,In_340);
or U1178 (N_1178,In_363,In_904);
nor U1179 (N_1179,In_763,In_853);
and U1180 (N_1180,In_119,In_423);
nor U1181 (N_1181,In_1,In_763);
and U1182 (N_1182,In_363,In_413);
and U1183 (N_1183,In_131,In_213);
or U1184 (N_1184,In_274,In_875);
nor U1185 (N_1185,In_34,In_561);
nand U1186 (N_1186,In_686,In_646);
or U1187 (N_1187,In_501,In_483);
nor U1188 (N_1188,In_316,In_432);
nand U1189 (N_1189,In_492,In_837);
nor U1190 (N_1190,In_827,In_40);
nor U1191 (N_1191,In_184,In_672);
nor U1192 (N_1192,In_83,In_93);
nor U1193 (N_1193,In_546,In_195);
or U1194 (N_1194,In_77,In_740);
or U1195 (N_1195,In_698,In_574);
nand U1196 (N_1196,In_588,In_537);
nor U1197 (N_1197,In_809,In_638);
nor U1198 (N_1198,In_271,In_422);
and U1199 (N_1199,In_150,In_393);
or U1200 (N_1200,In_988,In_451);
or U1201 (N_1201,In_653,In_87);
nand U1202 (N_1202,In_485,In_158);
or U1203 (N_1203,In_184,In_213);
and U1204 (N_1204,In_324,In_823);
nand U1205 (N_1205,In_185,In_668);
and U1206 (N_1206,In_79,In_850);
or U1207 (N_1207,In_923,In_46);
nor U1208 (N_1208,In_342,In_950);
and U1209 (N_1209,In_886,In_545);
nand U1210 (N_1210,In_657,In_875);
nor U1211 (N_1211,In_206,In_428);
or U1212 (N_1212,In_863,In_925);
and U1213 (N_1213,In_382,In_2);
and U1214 (N_1214,In_333,In_375);
or U1215 (N_1215,In_514,In_528);
nand U1216 (N_1216,In_855,In_937);
or U1217 (N_1217,In_473,In_370);
or U1218 (N_1218,In_625,In_879);
xnor U1219 (N_1219,In_389,In_877);
nor U1220 (N_1220,In_407,In_501);
nor U1221 (N_1221,In_117,In_524);
nor U1222 (N_1222,In_832,In_290);
or U1223 (N_1223,In_674,In_534);
or U1224 (N_1224,In_454,In_240);
and U1225 (N_1225,In_673,In_899);
xnor U1226 (N_1226,In_914,In_971);
nor U1227 (N_1227,In_986,In_361);
nand U1228 (N_1228,In_559,In_435);
or U1229 (N_1229,In_678,In_821);
and U1230 (N_1230,In_572,In_565);
nor U1231 (N_1231,In_161,In_896);
and U1232 (N_1232,In_169,In_562);
and U1233 (N_1233,In_948,In_865);
or U1234 (N_1234,In_427,In_302);
or U1235 (N_1235,In_455,In_697);
nand U1236 (N_1236,In_358,In_594);
or U1237 (N_1237,In_690,In_49);
or U1238 (N_1238,In_7,In_406);
and U1239 (N_1239,In_51,In_266);
or U1240 (N_1240,In_191,In_141);
and U1241 (N_1241,In_346,In_577);
and U1242 (N_1242,In_536,In_545);
or U1243 (N_1243,In_188,In_843);
or U1244 (N_1244,In_499,In_540);
and U1245 (N_1245,In_859,In_37);
nand U1246 (N_1246,In_618,In_172);
nand U1247 (N_1247,In_491,In_307);
nand U1248 (N_1248,In_77,In_825);
and U1249 (N_1249,In_159,In_25);
nor U1250 (N_1250,In_583,In_236);
nor U1251 (N_1251,In_806,In_255);
and U1252 (N_1252,In_428,In_510);
and U1253 (N_1253,In_416,In_363);
nand U1254 (N_1254,In_8,In_969);
nor U1255 (N_1255,In_649,In_348);
and U1256 (N_1256,In_984,In_565);
nor U1257 (N_1257,In_547,In_594);
nand U1258 (N_1258,In_572,In_487);
nor U1259 (N_1259,In_735,In_227);
or U1260 (N_1260,In_970,In_621);
or U1261 (N_1261,In_514,In_952);
nor U1262 (N_1262,In_21,In_580);
and U1263 (N_1263,In_805,In_561);
nor U1264 (N_1264,In_889,In_901);
nor U1265 (N_1265,In_516,In_164);
nand U1266 (N_1266,In_488,In_923);
nand U1267 (N_1267,In_399,In_534);
or U1268 (N_1268,In_905,In_239);
or U1269 (N_1269,In_253,In_535);
and U1270 (N_1270,In_294,In_305);
nor U1271 (N_1271,In_856,In_405);
or U1272 (N_1272,In_614,In_684);
and U1273 (N_1273,In_830,In_918);
or U1274 (N_1274,In_912,In_939);
nand U1275 (N_1275,In_609,In_735);
and U1276 (N_1276,In_180,In_782);
nor U1277 (N_1277,In_808,In_216);
nand U1278 (N_1278,In_255,In_802);
and U1279 (N_1279,In_158,In_374);
and U1280 (N_1280,In_557,In_2);
nor U1281 (N_1281,In_718,In_311);
xor U1282 (N_1282,In_193,In_648);
or U1283 (N_1283,In_783,In_487);
and U1284 (N_1284,In_582,In_274);
nand U1285 (N_1285,In_819,In_558);
or U1286 (N_1286,In_454,In_641);
nor U1287 (N_1287,In_63,In_921);
and U1288 (N_1288,In_858,In_824);
nand U1289 (N_1289,In_462,In_802);
nand U1290 (N_1290,In_235,In_312);
nand U1291 (N_1291,In_909,In_166);
and U1292 (N_1292,In_734,In_843);
or U1293 (N_1293,In_160,In_716);
nand U1294 (N_1294,In_333,In_833);
nor U1295 (N_1295,In_161,In_511);
and U1296 (N_1296,In_423,In_979);
nor U1297 (N_1297,In_780,In_896);
or U1298 (N_1298,In_437,In_253);
or U1299 (N_1299,In_214,In_944);
and U1300 (N_1300,In_955,In_160);
or U1301 (N_1301,In_314,In_515);
or U1302 (N_1302,In_229,In_627);
and U1303 (N_1303,In_588,In_185);
or U1304 (N_1304,In_260,In_147);
and U1305 (N_1305,In_286,In_75);
or U1306 (N_1306,In_357,In_664);
nor U1307 (N_1307,In_395,In_43);
nor U1308 (N_1308,In_794,In_832);
and U1309 (N_1309,In_861,In_938);
or U1310 (N_1310,In_339,In_112);
or U1311 (N_1311,In_824,In_584);
nand U1312 (N_1312,In_13,In_223);
nand U1313 (N_1313,In_597,In_807);
nor U1314 (N_1314,In_289,In_861);
or U1315 (N_1315,In_806,In_15);
nor U1316 (N_1316,In_843,In_367);
nand U1317 (N_1317,In_426,In_393);
and U1318 (N_1318,In_211,In_793);
nor U1319 (N_1319,In_3,In_911);
and U1320 (N_1320,In_943,In_234);
nor U1321 (N_1321,In_31,In_346);
nand U1322 (N_1322,In_981,In_178);
nor U1323 (N_1323,In_790,In_192);
or U1324 (N_1324,In_309,In_677);
nor U1325 (N_1325,In_512,In_688);
and U1326 (N_1326,In_473,In_94);
or U1327 (N_1327,In_537,In_379);
or U1328 (N_1328,In_963,In_75);
or U1329 (N_1329,In_324,In_195);
nor U1330 (N_1330,In_891,In_468);
nand U1331 (N_1331,In_986,In_147);
and U1332 (N_1332,In_264,In_522);
xor U1333 (N_1333,In_525,In_209);
nor U1334 (N_1334,In_534,In_775);
or U1335 (N_1335,In_228,In_798);
and U1336 (N_1336,In_532,In_682);
xnor U1337 (N_1337,In_796,In_90);
and U1338 (N_1338,In_502,In_86);
or U1339 (N_1339,In_608,In_222);
or U1340 (N_1340,In_7,In_595);
nand U1341 (N_1341,In_974,In_579);
nand U1342 (N_1342,In_126,In_739);
or U1343 (N_1343,In_912,In_52);
nor U1344 (N_1344,In_499,In_484);
and U1345 (N_1345,In_903,In_186);
or U1346 (N_1346,In_465,In_618);
xor U1347 (N_1347,In_837,In_352);
nand U1348 (N_1348,In_687,In_558);
nand U1349 (N_1349,In_623,In_409);
nand U1350 (N_1350,In_760,In_549);
and U1351 (N_1351,In_755,In_191);
nand U1352 (N_1352,In_168,In_637);
nand U1353 (N_1353,In_939,In_54);
and U1354 (N_1354,In_433,In_627);
nand U1355 (N_1355,In_331,In_115);
nor U1356 (N_1356,In_94,In_649);
nor U1357 (N_1357,In_711,In_336);
nor U1358 (N_1358,In_267,In_183);
nor U1359 (N_1359,In_188,In_185);
and U1360 (N_1360,In_19,In_519);
or U1361 (N_1361,In_123,In_39);
nand U1362 (N_1362,In_507,In_512);
or U1363 (N_1363,In_323,In_161);
nand U1364 (N_1364,In_860,In_522);
nand U1365 (N_1365,In_914,In_639);
nor U1366 (N_1366,In_10,In_698);
nor U1367 (N_1367,In_741,In_905);
nor U1368 (N_1368,In_170,In_917);
and U1369 (N_1369,In_872,In_898);
or U1370 (N_1370,In_546,In_622);
or U1371 (N_1371,In_282,In_536);
nand U1372 (N_1372,In_310,In_960);
nor U1373 (N_1373,In_686,In_933);
or U1374 (N_1374,In_392,In_842);
or U1375 (N_1375,In_66,In_436);
xnor U1376 (N_1376,In_274,In_930);
and U1377 (N_1377,In_869,In_3);
or U1378 (N_1378,In_523,In_697);
and U1379 (N_1379,In_623,In_593);
nor U1380 (N_1380,In_582,In_503);
nor U1381 (N_1381,In_986,In_82);
nand U1382 (N_1382,In_244,In_281);
and U1383 (N_1383,In_654,In_357);
nor U1384 (N_1384,In_972,In_741);
or U1385 (N_1385,In_945,In_234);
nand U1386 (N_1386,In_478,In_391);
nor U1387 (N_1387,In_772,In_634);
nand U1388 (N_1388,In_829,In_102);
nor U1389 (N_1389,In_719,In_624);
or U1390 (N_1390,In_328,In_188);
nor U1391 (N_1391,In_145,In_518);
nor U1392 (N_1392,In_219,In_223);
or U1393 (N_1393,In_69,In_561);
nor U1394 (N_1394,In_75,In_782);
or U1395 (N_1395,In_555,In_941);
or U1396 (N_1396,In_465,In_197);
and U1397 (N_1397,In_501,In_892);
nand U1398 (N_1398,In_772,In_428);
nor U1399 (N_1399,In_983,In_187);
nand U1400 (N_1400,In_554,In_302);
or U1401 (N_1401,In_794,In_211);
and U1402 (N_1402,In_518,In_372);
nand U1403 (N_1403,In_365,In_355);
or U1404 (N_1404,In_441,In_979);
nor U1405 (N_1405,In_979,In_765);
or U1406 (N_1406,In_255,In_831);
or U1407 (N_1407,In_721,In_764);
nand U1408 (N_1408,In_947,In_644);
nor U1409 (N_1409,In_81,In_230);
and U1410 (N_1410,In_408,In_898);
or U1411 (N_1411,In_449,In_502);
nand U1412 (N_1412,In_104,In_448);
nand U1413 (N_1413,In_300,In_866);
nand U1414 (N_1414,In_835,In_26);
nor U1415 (N_1415,In_955,In_716);
nor U1416 (N_1416,In_963,In_926);
xnor U1417 (N_1417,In_724,In_496);
nand U1418 (N_1418,In_227,In_515);
and U1419 (N_1419,In_827,In_737);
nand U1420 (N_1420,In_77,In_778);
or U1421 (N_1421,In_437,In_224);
or U1422 (N_1422,In_144,In_520);
and U1423 (N_1423,In_604,In_57);
or U1424 (N_1424,In_687,In_328);
or U1425 (N_1425,In_954,In_373);
nor U1426 (N_1426,In_864,In_204);
nand U1427 (N_1427,In_735,In_61);
nand U1428 (N_1428,In_576,In_877);
nor U1429 (N_1429,In_457,In_21);
or U1430 (N_1430,In_344,In_215);
nand U1431 (N_1431,In_66,In_241);
nand U1432 (N_1432,In_293,In_11);
nand U1433 (N_1433,In_167,In_236);
nand U1434 (N_1434,In_348,In_660);
or U1435 (N_1435,In_705,In_364);
or U1436 (N_1436,In_922,In_138);
and U1437 (N_1437,In_521,In_585);
nor U1438 (N_1438,In_261,In_855);
or U1439 (N_1439,In_76,In_684);
or U1440 (N_1440,In_563,In_271);
nand U1441 (N_1441,In_108,In_144);
nor U1442 (N_1442,In_965,In_557);
nor U1443 (N_1443,In_660,In_990);
nand U1444 (N_1444,In_698,In_18);
or U1445 (N_1445,In_525,In_271);
nor U1446 (N_1446,In_3,In_401);
nor U1447 (N_1447,In_666,In_162);
or U1448 (N_1448,In_14,In_234);
nor U1449 (N_1449,In_428,In_386);
and U1450 (N_1450,In_268,In_982);
nor U1451 (N_1451,In_261,In_63);
nor U1452 (N_1452,In_9,In_179);
nand U1453 (N_1453,In_947,In_225);
nor U1454 (N_1454,In_348,In_793);
xor U1455 (N_1455,In_900,In_274);
nor U1456 (N_1456,In_420,In_328);
and U1457 (N_1457,In_942,In_65);
nor U1458 (N_1458,In_73,In_386);
or U1459 (N_1459,In_10,In_325);
and U1460 (N_1460,In_569,In_994);
nor U1461 (N_1461,In_495,In_288);
or U1462 (N_1462,In_173,In_635);
or U1463 (N_1463,In_773,In_819);
and U1464 (N_1464,In_978,In_739);
xor U1465 (N_1465,In_658,In_338);
nand U1466 (N_1466,In_503,In_639);
nand U1467 (N_1467,In_742,In_813);
or U1468 (N_1468,In_676,In_47);
nor U1469 (N_1469,In_311,In_217);
and U1470 (N_1470,In_263,In_822);
nor U1471 (N_1471,In_426,In_368);
nand U1472 (N_1472,In_403,In_604);
and U1473 (N_1473,In_643,In_933);
or U1474 (N_1474,In_579,In_998);
or U1475 (N_1475,In_364,In_481);
or U1476 (N_1476,In_530,In_459);
nor U1477 (N_1477,In_444,In_726);
and U1478 (N_1478,In_339,In_88);
nor U1479 (N_1479,In_975,In_683);
or U1480 (N_1480,In_932,In_531);
or U1481 (N_1481,In_935,In_740);
nor U1482 (N_1482,In_588,In_772);
nand U1483 (N_1483,In_576,In_531);
nor U1484 (N_1484,In_585,In_792);
and U1485 (N_1485,In_968,In_334);
nand U1486 (N_1486,In_848,In_47);
nor U1487 (N_1487,In_940,In_621);
and U1488 (N_1488,In_193,In_366);
and U1489 (N_1489,In_270,In_48);
nand U1490 (N_1490,In_130,In_875);
and U1491 (N_1491,In_191,In_337);
nor U1492 (N_1492,In_510,In_253);
nor U1493 (N_1493,In_590,In_103);
nor U1494 (N_1494,In_389,In_202);
or U1495 (N_1495,In_716,In_647);
or U1496 (N_1496,In_30,In_831);
nand U1497 (N_1497,In_786,In_345);
and U1498 (N_1498,In_666,In_881);
nor U1499 (N_1499,In_379,In_831);
or U1500 (N_1500,In_998,In_53);
or U1501 (N_1501,In_346,In_114);
or U1502 (N_1502,In_984,In_236);
nand U1503 (N_1503,In_502,In_104);
or U1504 (N_1504,In_405,In_965);
nor U1505 (N_1505,In_215,In_38);
nor U1506 (N_1506,In_764,In_533);
or U1507 (N_1507,In_632,In_356);
nor U1508 (N_1508,In_689,In_906);
xnor U1509 (N_1509,In_643,In_554);
nand U1510 (N_1510,In_750,In_395);
nor U1511 (N_1511,In_185,In_367);
nor U1512 (N_1512,In_71,In_936);
nand U1513 (N_1513,In_759,In_470);
and U1514 (N_1514,In_454,In_157);
and U1515 (N_1515,In_639,In_255);
and U1516 (N_1516,In_333,In_170);
and U1517 (N_1517,In_219,In_474);
nor U1518 (N_1518,In_229,In_586);
or U1519 (N_1519,In_355,In_620);
or U1520 (N_1520,In_324,In_392);
nor U1521 (N_1521,In_116,In_119);
and U1522 (N_1522,In_483,In_147);
nand U1523 (N_1523,In_684,In_357);
xor U1524 (N_1524,In_179,In_850);
or U1525 (N_1525,In_627,In_616);
nor U1526 (N_1526,In_573,In_431);
nor U1527 (N_1527,In_484,In_227);
nand U1528 (N_1528,In_540,In_734);
nand U1529 (N_1529,In_707,In_702);
and U1530 (N_1530,In_877,In_357);
nand U1531 (N_1531,In_359,In_880);
and U1532 (N_1532,In_921,In_156);
nand U1533 (N_1533,In_812,In_483);
nor U1534 (N_1534,In_136,In_829);
or U1535 (N_1535,In_252,In_854);
nand U1536 (N_1536,In_504,In_777);
or U1537 (N_1537,In_736,In_705);
nor U1538 (N_1538,In_815,In_261);
nor U1539 (N_1539,In_775,In_976);
nor U1540 (N_1540,In_531,In_957);
nand U1541 (N_1541,In_682,In_351);
nand U1542 (N_1542,In_177,In_483);
nand U1543 (N_1543,In_913,In_613);
nor U1544 (N_1544,In_638,In_71);
and U1545 (N_1545,In_16,In_984);
or U1546 (N_1546,In_641,In_986);
nor U1547 (N_1547,In_458,In_39);
or U1548 (N_1548,In_396,In_358);
nand U1549 (N_1549,In_972,In_185);
nand U1550 (N_1550,In_793,In_648);
and U1551 (N_1551,In_963,In_958);
or U1552 (N_1552,In_401,In_296);
nor U1553 (N_1553,In_872,In_687);
nand U1554 (N_1554,In_813,In_110);
nor U1555 (N_1555,In_155,In_135);
xor U1556 (N_1556,In_311,In_91);
or U1557 (N_1557,In_214,In_673);
or U1558 (N_1558,In_733,In_803);
nand U1559 (N_1559,In_34,In_67);
and U1560 (N_1560,In_898,In_244);
nand U1561 (N_1561,In_743,In_222);
or U1562 (N_1562,In_137,In_507);
or U1563 (N_1563,In_861,In_407);
nor U1564 (N_1564,In_44,In_172);
nor U1565 (N_1565,In_346,In_613);
nor U1566 (N_1566,In_159,In_526);
or U1567 (N_1567,In_329,In_939);
or U1568 (N_1568,In_37,In_159);
and U1569 (N_1569,In_590,In_725);
and U1570 (N_1570,In_176,In_38);
and U1571 (N_1571,In_763,In_589);
nor U1572 (N_1572,In_323,In_81);
nor U1573 (N_1573,In_644,In_741);
or U1574 (N_1574,In_105,In_885);
nor U1575 (N_1575,In_465,In_579);
or U1576 (N_1576,In_908,In_95);
nand U1577 (N_1577,In_927,In_766);
nor U1578 (N_1578,In_404,In_623);
nand U1579 (N_1579,In_730,In_542);
nand U1580 (N_1580,In_55,In_336);
xor U1581 (N_1581,In_437,In_267);
nand U1582 (N_1582,In_52,In_273);
nor U1583 (N_1583,In_517,In_377);
and U1584 (N_1584,In_382,In_810);
nand U1585 (N_1585,In_27,In_449);
nand U1586 (N_1586,In_837,In_483);
and U1587 (N_1587,In_97,In_455);
xor U1588 (N_1588,In_213,In_798);
nand U1589 (N_1589,In_972,In_107);
and U1590 (N_1590,In_108,In_168);
or U1591 (N_1591,In_446,In_825);
and U1592 (N_1592,In_338,In_588);
and U1593 (N_1593,In_950,In_845);
nand U1594 (N_1594,In_735,In_194);
or U1595 (N_1595,In_722,In_882);
and U1596 (N_1596,In_261,In_343);
nor U1597 (N_1597,In_326,In_216);
and U1598 (N_1598,In_528,In_319);
nor U1599 (N_1599,In_476,In_215);
nor U1600 (N_1600,In_534,In_246);
and U1601 (N_1601,In_825,In_468);
nand U1602 (N_1602,In_15,In_241);
nand U1603 (N_1603,In_613,In_267);
and U1604 (N_1604,In_353,In_64);
nand U1605 (N_1605,In_265,In_609);
and U1606 (N_1606,In_761,In_815);
or U1607 (N_1607,In_834,In_806);
nand U1608 (N_1608,In_315,In_752);
or U1609 (N_1609,In_162,In_792);
or U1610 (N_1610,In_259,In_562);
nor U1611 (N_1611,In_436,In_540);
and U1612 (N_1612,In_35,In_775);
nor U1613 (N_1613,In_572,In_533);
nand U1614 (N_1614,In_629,In_375);
nand U1615 (N_1615,In_656,In_229);
nand U1616 (N_1616,In_507,In_668);
nor U1617 (N_1617,In_374,In_737);
and U1618 (N_1618,In_357,In_442);
or U1619 (N_1619,In_100,In_264);
nand U1620 (N_1620,In_32,In_93);
nand U1621 (N_1621,In_73,In_423);
and U1622 (N_1622,In_931,In_264);
and U1623 (N_1623,In_930,In_775);
nand U1624 (N_1624,In_420,In_578);
or U1625 (N_1625,In_641,In_169);
or U1626 (N_1626,In_974,In_39);
and U1627 (N_1627,In_35,In_34);
and U1628 (N_1628,In_154,In_33);
or U1629 (N_1629,In_571,In_167);
or U1630 (N_1630,In_168,In_995);
or U1631 (N_1631,In_623,In_136);
nand U1632 (N_1632,In_659,In_595);
or U1633 (N_1633,In_83,In_595);
and U1634 (N_1634,In_274,In_100);
and U1635 (N_1635,In_394,In_706);
or U1636 (N_1636,In_319,In_536);
nand U1637 (N_1637,In_501,In_925);
or U1638 (N_1638,In_668,In_372);
nor U1639 (N_1639,In_694,In_515);
nor U1640 (N_1640,In_738,In_764);
and U1641 (N_1641,In_700,In_75);
and U1642 (N_1642,In_720,In_132);
nand U1643 (N_1643,In_728,In_329);
and U1644 (N_1644,In_90,In_781);
nor U1645 (N_1645,In_121,In_573);
or U1646 (N_1646,In_757,In_456);
nor U1647 (N_1647,In_935,In_429);
xor U1648 (N_1648,In_49,In_759);
nor U1649 (N_1649,In_242,In_645);
and U1650 (N_1650,In_705,In_320);
or U1651 (N_1651,In_180,In_692);
nand U1652 (N_1652,In_948,In_784);
or U1653 (N_1653,In_599,In_462);
nand U1654 (N_1654,In_229,In_730);
or U1655 (N_1655,In_93,In_853);
nand U1656 (N_1656,In_163,In_21);
or U1657 (N_1657,In_977,In_561);
or U1658 (N_1658,In_164,In_924);
and U1659 (N_1659,In_799,In_871);
nor U1660 (N_1660,In_726,In_216);
or U1661 (N_1661,In_571,In_879);
or U1662 (N_1662,In_69,In_684);
and U1663 (N_1663,In_43,In_753);
nand U1664 (N_1664,In_175,In_914);
and U1665 (N_1665,In_191,In_947);
or U1666 (N_1666,In_912,In_482);
nand U1667 (N_1667,In_201,In_673);
and U1668 (N_1668,In_325,In_811);
or U1669 (N_1669,In_915,In_178);
or U1670 (N_1670,In_331,In_661);
nor U1671 (N_1671,In_485,In_464);
and U1672 (N_1672,In_627,In_889);
nand U1673 (N_1673,In_267,In_679);
nand U1674 (N_1674,In_837,In_219);
nor U1675 (N_1675,In_347,In_359);
or U1676 (N_1676,In_301,In_310);
nor U1677 (N_1677,In_977,In_923);
nand U1678 (N_1678,In_758,In_145);
and U1679 (N_1679,In_561,In_943);
or U1680 (N_1680,In_685,In_553);
and U1681 (N_1681,In_199,In_317);
nand U1682 (N_1682,In_451,In_871);
nor U1683 (N_1683,In_726,In_21);
nand U1684 (N_1684,In_170,In_60);
and U1685 (N_1685,In_312,In_500);
nand U1686 (N_1686,In_912,In_381);
or U1687 (N_1687,In_289,In_650);
nand U1688 (N_1688,In_271,In_863);
nand U1689 (N_1689,In_925,In_602);
xor U1690 (N_1690,In_316,In_318);
xnor U1691 (N_1691,In_452,In_787);
and U1692 (N_1692,In_171,In_348);
and U1693 (N_1693,In_84,In_129);
nand U1694 (N_1694,In_496,In_156);
nor U1695 (N_1695,In_445,In_85);
or U1696 (N_1696,In_409,In_761);
xnor U1697 (N_1697,In_135,In_95);
and U1698 (N_1698,In_11,In_708);
nor U1699 (N_1699,In_178,In_448);
and U1700 (N_1700,In_306,In_33);
nand U1701 (N_1701,In_378,In_492);
or U1702 (N_1702,In_56,In_977);
and U1703 (N_1703,In_749,In_12);
nand U1704 (N_1704,In_778,In_967);
nor U1705 (N_1705,In_497,In_839);
nor U1706 (N_1706,In_397,In_65);
nand U1707 (N_1707,In_833,In_224);
nand U1708 (N_1708,In_626,In_746);
nand U1709 (N_1709,In_750,In_553);
nand U1710 (N_1710,In_846,In_686);
nor U1711 (N_1711,In_236,In_902);
and U1712 (N_1712,In_769,In_950);
or U1713 (N_1713,In_115,In_13);
or U1714 (N_1714,In_913,In_621);
and U1715 (N_1715,In_511,In_999);
nor U1716 (N_1716,In_459,In_434);
or U1717 (N_1717,In_540,In_547);
nor U1718 (N_1718,In_926,In_499);
nand U1719 (N_1719,In_23,In_486);
nor U1720 (N_1720,In_332,In_189);
nor U1721 (N_1721,In_935,In_796);
xor U1722 (N_1722,In_875,In_146);
nand U1723 (N_1723,In_97,In_750);
xor U1724 (N_1724,In_267,In_181);
nand U1725 (N_1725,In_123,In_978);
nand U1726 (N_1726,In_439,In_93);
and U1727 (N_1727,In_680,In_770);
and U1728 (N_1728,In_964,In_182);
and U1729 (N_1729,In_427,In_66);
nor U1730 (N_1730,In_601,In_109);
nor U1731 (N_1731,In_977,In_157);
or U1732 (N_1732,In_395,In_776);
nor U1733 (N_1733,In_991,In_198);
nand U1734 (N_1734,In_70,In_347);
or U1735 (N_1735,In_136,In_338);
nor U1736 (N_1736,In_683,In_183);
and U1737 (N_1737,In_990,In_994);
and U1738 (N_1738,In_253,In_164);
and U1739 (N_1739,In_224,In_623);
or U1740 (N_1740,In_567,In_459);
or U1741 (N_1741,In_601,In_406);
or U1742 (N_1742,In_852,In_772);
or U1743 (N_1743,In_361,In_913);
nor U1744 (N_1744,In_541,In_941);
nor U1745 (N_1745,In_174,In_925);
nor U1746 (N_1746,In_850,In_189);
nand U1747 (N_1747,In_557,In_555);
and U1748 (N_1748,In_219,In_207);
nor U1749 (N_1749,In_596,In_83);
or U1750 (N_1750,In_902,In_255);
nor U1751 (N_1751,In_569,In_395);
or U1752 (N_1752,In_225,In_453);
or U1753 (N_1753,In_300,In_641);
nand U1754 (N_1754,In_815,In_764);
nand U1755 (N_1755,In_506,In_8);
or U1756 (N_1756,In_506,In_632);
nand U1757 (N_1757,In_595,In_319);
or U1758 (N_1758,In_713,In_625);
nor U1759 (N_1759,In_984,In_829);
or U1760 (N_1760,In_38,In_638);
nand U1761 (N_1761,In_323,In_888);
and U1762 (N_1762,In_191,In_64);
nand U1763 (N_1763,In_475,In_493);
nand U1764 (N_1764,In_724,In_222);
and U1765 (N_1765,In_226,In_614);
nand U1766 (N_1766,In_656,In_31);
and U1767 (N_1767,In_971,In_384);
and U1768 (N_1768,In_575,In_320);
nand U1769 (N_1769,In_484,In_431);
nand U1770 (N_1770,In_173,In_521);
or U1771 (N_1771,In_215,In_985);
nand U1772 (N_1772,In_903,In_871);
nor U1773 (N_1773,In_309,In_553);
nand U1774 (N_1774,In_36,In_614);
nand U1775 (N_1775,In_647,In_159);
nor U1776 (N_1776,In_139,In_437);
nor U1777 (N_1777,In_547,In_596);
nand U1778 (N_1778,In_334,In_896);
nor U1779 (N_1779,In_802,In_374);
and U1780 (N_1780,In_799,In_44);
or U1781 (N_1781,In_21,In_247);
or U1782 (N_1782,In_866,In_39);
nand U1783 (N_1783,In_559,In_430);
xor U1784 (N_1784,In_676,In_256);
and U1785 (N_1785,In_525,In_624);
or U1786 (N_1786,In_15,In_147);
nand U1787 (N_1787,In_707,In_521);
or U1788 (N_1788,In_126,In_292);
nand U1789 (N_1789,In_380,In_715);
xnor U1790 (N_1790,In_695,In_961);
nor U1791 (N_1791,In_400,In_273);
or U1792 (N_1792,In_949,In_714);
or U1793 (N_1793,In_3,In_602);
and U1794 (N_1794,In_536,In_996);
or U1795 (N_1795,In_149,In_622);
and U1796 (N_1796,In_508,In_207);
nand U1797 (N_1797,In_816,In_830);
and U1798 (N_1798,In_407,In_931);
or U1799 (N_1799,In_291,In_51);
nor U1800 (N_1800,In_206,In_318);
or U1801 (N_1801,In_27,In_547);
or U1802 (N_1802,In_328,In_94);
and U1803 (N_1803,In_449,In_109);
xor U1804 (N_1804,In_155,In_117);
nand U1805 (N_1805,In_642,In_26);
nand U1806 (N_1806,In_725,In_51);
nor U1807 (N_1807,In_815,In_421);
or U1808 (N_1808,In_941,In_727);
nor U1809 (N_1809,In_790,In_401);
and U1810 (N_1810,In_127,In_139);
and U1811 (N_1811,In_445,In_71);
nand U1812 (N_1812,In_349,In_559);
nand U1813 (N_1813,In_717,In_62);
and U1814 (N_1814,In_798,In_721);
and U1815 (N_1815,In_214,In_336);
or U1816 (N_1816,In_835,In_165);
nand U1817 (N_1817,In_118,In_776);
nor U1818 (N_1818,In_257,In_919);
or U1819 (N_1819,In_349,In_293);
nor U1820 (N_1820,In_403,In_205);
nor U1821 (N_1821,In_887,In_798);
nor U1822 (N_1822,In_609,In_832);
nand U1823 (N_1823,In_612,In_349);
nand U1824 (N_1824,In_835,In_380);
or U1825 (N_1825,In_897,In_102);
and U1826 (N_1826,In_916,In_775);
or U1827 (N_1827,In_994,In_954);
nand U1828 (N_1828,In_25,In_9);
nor U1829 (N_1829,In_279,In_214);
nor U1830 (N_1830,In_52,In_927);
nand U1831 (N_1831,In_153,In_367);
xnor U1832 (N_1832,In_466,In_842);
nor U1833 (N_1833,In_636,In_740);
and U1834 (N_1834,In_413,In_211);
nor U1835 (N_1835,In_948,In_715);
or U1836 (N_1836,In_338,In_510);
and U1837 (N_1837,In_466,In_614);
nand U1838 (N_1838,In_911,In_111);
nor U1839 (N_1839,In_554,In_777);
nor U1840 (N_1840,In_296,In_867);
and U1841 (N_1841,In_822,In_505);
nand U1842 (N_1842,In_23,In_305);
and U1843 (N_1843,In_14,In_621);
nand U1844 (N_1844,In_247,In_188);
nand U1845 (N_1845,In_115,In_644);
and U1846 (N_1846,In_274,In_644);
nand U1847 (N_1847,In_171,In_355);
or U1848 (N_1848,In_289,In_667);
nand U1849 (N_1849,In_938,In_871);
and U1850 (N_1850,In_481,In_945);
or U1851 (N_1851,In_51,In_855);
nand U1852 (N_1852,In_189,In_924);
and U1853 (N_1853,In_359,In_909);
nand U1854 (N_1854,In_144,In_196);
nor U1855 (N_1855,In_921,In_252);
nor U1856 (N_1856,In_126,In_560);
or U1857 (N_1857,In_535,In_161);
and U1858 (N_1858,In_310,In_657);
nand U1859 (N_1859,In_55,In_25);
and U1860 (N_1860,In_762,In_474);
nor U1861 (N_1861,In_339,In_19);
or U1862 (N_1862,In_992,In_497);
nand U1863 (N_1863,In_458,In_887);
nor U1864 (N_1864,In_282,In_232);
nand U1865 (N_1865,In_757,In_7);
or U1866 (N_1866,In_179,In_386);
or U1867 (N_1867,In_940,In_741);
nor U1868 (N_1868,In_216,In_507);
nor U1869 (N_1869,In_50,In_314);
and U1870 (N_1870,In_896,In_255);
nand U1871 (N_1871,In_493,In_830);
nand U1872 (N_1872,In_808,In_384);
nand U1873 (N_1873,In_882,In_533);
nand U1874 (N_1874,In_54,In_683);
and U1875 (N_1875,In_967,In_556);
nand U1876 (N_1876,In_465,In_905);
nand U1877 (N_1877,In_582,In_753);
or U1878 (N_1878,In_33,In_992);
nor U1879 (N_1879,In_661,In_35);
or U1880 (N_1880,In_434,In_646);
or U1881 (N_1881,In_584,In_952);
nor U1882 (N_1882,In_596,In_8);
and U1883 (N_1883,In_846,In_467);
and U1884 (N_1884,In_719,In_697);
or U1885 (N_1885,In_76,In_408);
and U1886 (N_1886,In_405,In_360);
nor U1887 (N_1887,In_460,In_93);
or U1888 (N_1888,In_526,In_425);
and U1889 (N_1889,In_934,In_394);
and U1890 (N_1890,In_220,In_445);
xor U1891 (N_1891,In_3,In_436);
or U1892 (N_1892,In_738,In_654);
and U1893 (N_1893,In_601,In_861);
xor U1894 (N_1894,In_191,In_407);
or U1895 (N_1895,In_189,In_835);
or U1896 (N_1896,In_177,In_799);
or U1897 (N_1897,In_995,In_449);
and U1898 (N_1898,In_901,In_639);
or U1899 (N_1899,In_94,In_828);
nor U1900 (N_1900,In_991,In_566);
nor U1901 (N_1901,In_591,In_663);
nand U1902 (N_1902,In_833,In_564);
or U1903 (N_1903,In_132,In_795);
nor U1904 (N_1904,In_914,In_77);
nor U1905 (N_1905,In_434,In_133);
nor U1906 (N_1906,In_584,In_10);
and U1907 (N_1907,In_66,In_559);
nor U1908 (N_1908,In_604,In_49);
and U1909 (N_1909,In_784,In_201);
nor U1910 (N_1910,In_933,In_237);
nor U1911 (N_1911,In_489,In_256);
or U1912 (N_1912,In_446,In_553);
and U1913 (N_1913,In_650,In_619);
nor U1914 (N_1914,In_846,In_65);
or U1915 (N_1915,In_170,In_950);
and U1916 (N_1916,In_17,In_921);
and U1917 (N_1917,In_389,In_141);
nor U1918 (N_1918,In_881,In_356);
or U1919 (N_1919,In_459,In_645);
and U1920 (N_1920,In_958,In_508);
and U1921 (N_1921,In_854,In_903);
nor U1922 (N_1922,In_339,In_486);
nor U1923 (N_1923,In_440,In_737);
and U1924 (N_1924,In_937,In_492);
nand U1925 (N_1925,In_908,In_998);
and U1926 (N_1926,In_775,In_885);
nor U1927 (N_1927,In_841,In_932);
nor U1928 (N_1928,In_143,In_770);
or U1929 (N_1929,In_607,In_438);
nand U1930 (N_1930,In_561,In_800);
nand U1931 (N_1931,In_132,In_808);
xnor U1932 (N_1932,In_625,In_988);
and U1933 (N_1933,In_492,In_359);
or U1934 (N_1934,In_297,In_647);
or U1935 (N_1935,In_582,In_429);
and U1936 (N_1936,In_389,In_432);
nor U1937 (N_1937,In_968,In_319);
nand U1938 (N_1938,In_735,In_329);
nand U1939 (N_1939,In_379,In_947);
nand U1940 (N_1940,In_287,In_753);
or U1941 (N_1941,In_706,In_867);
and U1942 (N_1942,In_342,In_865);
nor U1943 (N_1943,In_718,In_214);
and U1944 (N_1944,In_296,In_945);
or U1945 (N_1945,In_824,In_753);
nor U1946 (N_1946,In_632,In_210);
nand U1947 (N_1947,In_283,In_252);
and U1948 (N_1948,In_666,In_869);
and U1949 (N_1949,In_46,In_760);
xnor U1950 (N_1950,In_443,In_349);
nand U1951 (N_1951,In_307,In_405);
and U1952 (N_1952,In_265,In_770);
or U1953 (N_1953,In_750,In_519);
nand U1954 (N_1954,In_309,In_397);
or U1955 (N_1955,In_344,In_736);
and U1956 (N_1956,In_148,In_824);
or U1957 (N_1957,In_989,In_412);
or U1958 (N_1958,In_736,In_490);
and U1959 (N_1959,In_557,In_530);
or U1960 (N_1960,In_376,In_225);
nor U1961 (N_1961,In_333,In_466);
nand U1962 (N_1962,In_250,In_780);
or U1963 (N_1963,In_508,In_652);
or U1964 (N_1964,In_984,In_720);
and U1965 (N_1965,In_754,In_492);
or U1966 (N_1966,In_236,In_894);
or U1967 (N_1967,In_665,In_29);
xor U1968 (N_1968,In_620,In_107);
nor U1969 (N_1969,In_206,In_643);
or U1970 (N_1970,In_718,In_133);
nor U1971 (N_1971,In_832,In_568);
or U1972 (N_1972,In_979,In_316);
or U1973 (N_1973,In_699,In_137);
and U1974 (N_1974,In_781,In_945);
nor U1975 (N_1975,In_41,In_871);
xor U1976 (N_1976,In_506,In_884);
nor U1977 (N_1977,In_532,In_500);
and U1978 (N_1978,In_30,In_723);
nor U1979 (N_1979,In_657,In_400);
or U1980 (N_1980,In_546,In_6);
nor U1981 (N_1981,In_663,In_482);
nand U1982 (N_1982,In_605,In_816);
and U1983 (N_1983,In_493,In_735);
xor U1984 (N_1984,In_600,In_324);
or U1985 (N_1985,In_632,In_63);
and U1986 (N_1986,In_234,In_175);
and U1987 (N_1987,In_560,In_944);
nand U1988 (N_1988,In_756,In_559);
nor U1989 (N_1989,In_829,In_163);
nor U1990 (N_1990,In_643,In_862);
or U1991 (N_1991,In_789,In_963);
or U1992 (N_1992,In_355,In_917);
and U1993 (N_1993,In_977,In_818);
nor U1994 (N_1994,In_283,In_626);
nand U1995 (N_1995,In_334,In_709);
nor U1996 (N_1996,In_166,In_927);
or U1997 (N_1997,In_622,In_247);
nand U1998 (N_1998,In_136,In_632);
nor U1999 (N_1999,In_229,In_809);
or U2000 (N_2000,N_879,N_442);
and U2001 (N_2001,N_1772,N_1261);
and U2002 (N_2002,N_1244,N_1659);
nor U2003 (N_2003,N_440,N_1307);
and U2004 (N_2004,N_983,N_805);
nand U2005 (N_2005,N_1057,N_353);
nand U2006 (N_2006,N_808,N_558);
and U2007 (N_2007,N_1375,N_1703);
xor U2008 (N_2008,N_295,N_10);
or U2009 (N_2009,N_119,N_886);
xor U2010 (N_2010,N_1252,N_1129);
nor U2011 (N_2011,N_1683,N_1037);
nor U2012 (N_2012,N_1367,N_1473);
nand U2013 (N_2013,N_1648,N_1004);
nand U2014 (N_2014,N_1290,N_1634);
or U2015 (N_2015,N_817,N_202);
nand U2016 (N_2016,N_1480,N_1530);
nand U2017 (N_2017,N_1064,N_449);
or U2018 (N_2018,N_168,N_1883);
or U2019 (N_2019,N_1087,N_261);
nor U2020 (N_2020,N_1785,N_1669);
or U2021 (N_2021,N_1327,N_1361);
xnor U2022 (N_2022,N_660,N_350);
nor U2023 (N_2023,N_782,N_634);
nand U2024 (N_2024,N_1387,N_315);
nand U2025 (N_2025,N_1423,N_1276);
nand U2026 (N_2026,N_146,N_7);
or U2027 (N_2027,N_1242,N_1750);
nor U2028 (N_2028,N_1233,N_1201);
or U2029 (N_2029,N_151,N_655);
and U2030 (N_2030,N_990,N_1408);
nand U2031 (N_2031,N_99,N_1968);
nand U2032 (N_2032,N_1902,N_316);
xor U2033 (N_2033,N_55,N_1250);
nand U2034 (N_2034,N_845,N_587);
and U2035 (N_2035,N_1954,N_737);
nor U2036 (N_2036,N_1826,N_632);
nand U2037 (N_2037,N_1690,N_87);
or U2038 (N_2038,N_452,N_1300);
nand U2039 (N_2039,N_1786,N_1085);
and U2040 (N_2040,N_1237,N_1781);
xnor U2041 (N_2041,N_1102,N_358);
and U2042 (N_2042,N_1165,N_616);
nor U2043 (N_2043,N_1831,N_161);
xor U2044 (N_2044,N_1534,N_1488);
and U2045 (N_2045,N_968,N_481);
and U2046 (N_2046,N_508,N_1892);
nor U2047 (N_2047,N_1662,N_1827);
or U2048 (N_2048,N_1868,N_33);
or U2049 (N_2049,N_412,N_1302);
and U2050 (N_2050,N_606,N_1305);
or U2051 (N_2051,N_838,N_901);
and U2052 (N_2052,N_665,N_1493);
and U2053 (N_2053,N_563,N_494);
nor U2054 (N_2054,N_1414,N_919);
nor U2055 (N_2055,N_1281,N_1208);
and U2056 (N_2056,N_1068,N_43);
nand U2057 (N_2057,N_195,N_1819);
or U2058 (N_2058,N_975,N_1602);
nor U2059 (N_2059,N_1841,N_944);
and U2060 (N_2060,N_1579,N_222);
or U2061 (N_2061,N_1097,N_1298);
and U2062 (N_2062,N_911,N_989);
nand U2063 (N_2063,N_1961,N_884);
nand U2064 (N_2064,N_1607,N_1294);
or U2065 (N_2065,N_1500,N_1823);
nand U2066 (N_2066,N_755,N_1432);
or U2067 (N_2067,N_1222,N_1855);
and U2068 (N_2068,N_1181,N_1696);
nor U2069 (N_2069,N_874,N_757);
and U2070 (N_2070,N_1199,N_468);
or U2071 (N_2071,N_285,N_1107);
nand U2072 (N_2072,N_601,N_1470);
nor U2073 (N_2073,N_1877,N_882);
nor U2074 (N_2074,N_383,N_1232);
or U2075 (N_2075,N_1725,N_1874);
and U2076 (N_2076,N_1542,N_305);
nor U2077 (N_2077,N_312,N_600);
or U2078 (N_2078,N_1718,N_594);
or U2079 (N_2079,N_98,N_188);
nor U2080 (N_2080,N_1840,N_1914);
or U2081 (N_2081,N_1507,N_623);
nor U2082 (N_2082,N_1635,N_1506);
xor U2083 (N_2083,N_740,N_1957);
or U2084 (N_2084,N_267,N_1582);
xor U2085 (N_2085,N_434,N_1809);
and U2086 (N_2086,N_724,N_60);
nor U2087 (N_2087,N_889,N_448);
nand U2088 (N_2088,N_1550,N_59);
and U2089 (N_2089,N_1235,N_1857);
and U2090 (N_2090,N_1538,N_1131);
or U2091 (N_2091,N_186,N_556);
and U2092 (N_2092,N_1436,N_226);
and U2093 (N_2093,N_795,N_1933);
nor U2094 (N_2094,N_1697,N_1929);
and U2095 (N_2095,N_1734,N_970);
or U2096 (N_2096,N_1454,N_44);
or U2097 (N_2097,N_1067,N_609);
nor U2098 (N_2098,N_368,N_986);
or U2099 (N_2099,N_235,N_612);
nand U2100 (N_2100,N_359,N_1562);
xor U2101 (N_2101,N_334,N_598);
and U2102 (N_2102,N_565,N_1600);
and U2103 (N_2103,N_1611,N_1701);
and U2104 (N_2104,N_1640,N_735);
and U2105 (N_2105,N_908,N_1969);
nand U2106 (N_2106,N_1006,N_890);
or U2107 (N_2107,N_1518,N_993);
nand U2108 (N_2108,N_197,N_876);
nand U2109 (N_2109,N_391,N_1134);
or U2110 (N_2110,N_995,N_144);
nand U2111 (N_2111,N_933,N_1282);
nand U2112 (N_2112,N_1873,N_713);
nor U2113 (N_2113,N_1391,N_388);
or U2114 (N_2114,N_1452,N_1625);
nor U2115 (N_2115,N_1073,N_716);
or U2116 (N_2116,N_1137,N_281);
or U2117 (N_2117,N_291,N_1706);
nor U2118 (N_2118,N_164,N_1974);
and U2119 (N_2119,N_252,N_469);
or U2120 (N_2120,N_303,N_1565);
nand U2121 (N_2121,N_187,N_20);
nand U2122 (N_2122,N_1918,N_1403);
nand U2123 (N_2123,N_1395,N_1077);
nand U2124 (N_2124,N_1450,N_1657);
nor U2125 (N_2125,N_318,N_1908);
and U2126 (N_2126,N_321,N_1462);
nor U2127 (N_2127,N_400,N_1025);
or U2128 (N_2128,N_210,N_117);
and U2129 (N_2129,N_324,N_75);
or U2130 (N_2130,N_384,N_552);
or U2131 (N_2131,N_1845,N_1140);
nor U2132 (N_2132,N_1901,N_1663);
and U2133 (N_2133,N_779,N_823);
and U2134 (N_2134,N_822,N_1529);
nor U2135 (N_2135,N_1489,N_910);
nor U2136 (N_2136,N_483,N_1641);
nand U2137 (N_2137,N_814,N_714);
nor U2138 (N_2138,N_1653,N_277);
nand U2139 (N_2139,N_873,N_1378);
and U2140 (N_2140,N_288,N_208);
nor U2141 (N_2141,N_668,N_1637);
nor U2142 (N_2142,N_1574,N_30);
or U2143 (N_2143,N_663,N_1977);
nor U2144 (N_2144,N_1339,N_806);
nand U2145 (N_2145,N_500,N_1859);
and U2146 (N_2146,N_535,N_1570);
nor U2147 (N_2147,N_1944,N_298);
and U2148 (N_2148,N_1495,N_1413);
or U2149 (N_2149,N_1265,N_1689);
and U2150 (N_2150,N_920,N_1490);
nand U2151 (N_2151,N_342,N_1712);
or U2152 (N_2152,N_1054,N_102);
or U2153 (N_2153,N_1870,N_122);
nand U2154 (N_2154,N_1956,N_1161);
nor U2155 (N_2155,N_923,N_752);
and U2156 (N_2156,N_193,N_465);
nor U2157 (N_2157,N_1854,N_1921);
or U2158 (N_2158,N_644,N_1084);
nor U2159 (N_2159,N_1224,N_491);
xnor U2160 (N_2160,N_649,N_1311);
and U2161 (N_2161,N_216,N_477);
and U2162 (N_2162,N_503,N_871);
and U2163 (N_2163,N_1952,N_1062);
nor U2164 (N_2164,N_774,N_1850);
and U2165 (N_2165,N_223,N_237);
nor U2166 (N_2166,N_541,N_775);
nand U2167 (N_2167,N_1978,N_1434);
nor U2168 (N_2168,N_1342,N_1775);
and U2169 (N_2169,N_666,N_1492);
nor U2170 (N_2170,N_1789,N_271);
nand U2171 (N_2171,N_626,N_1959);
nand U2172 (N_2172,N_238,N_249);
nor U2173 (N_2173,N_683,N_1899);
and U2174 (N_2174,N_524,N_1360);
or U2175 (N_2175,N_702,N_693);
nand U2176 (N_2176,N_1114,N_520);
and U2177 (N_2177,N_568,N_1098);
and U2178 (N_2178,N_1086,N_1658);
nand U2179 (N_2179,N_1048,N_1905);
or U2180 (N_2180,N_1404,N_425);
nand U2181 (N_2181,N_1504,N_1453);
nor U2182 (N_2182,N_1082,N_464);
nand U2183 (N_2183,N_977,N_341);
and U2184 (N_2184,N_573,N_641);
nand U2185 (N_2185,N_1843,N_739);
or U2186 (N_2186,N_569,N_1966);
or U2187 (N_2187,N_1245,N_894);
and U2188 (N_2188,N_527,N_1428);
nand U2189 (N_2189,N_893,N_1477);
nand U2190 (N_2190,N_505,N_1295);
nor U2191 (N_2191,N_332,N_785);
and U2192 (N_2192,N_559,N_1766);
nand U2193 (N_2193,N_1036,N_1458);
nor U2194 (N_2194,N_1430,N_1771);
and U2195 (N_2195,N_1846,N_1306);
nor U2196 (N_2196,N_380,N_972);
nand U2197 (N_2197,N_320,N_750);
nor U2198 (N_2198,N_366,N_1011);
nor U2199 (N_2199,N_1881,N_1100);
nand U2200 (N_2200,N_1805,N_141);
or U2201 (N_2201,N_1088,N_1885);
nand U2202 (N_2202,N_708,N_1108);
and U2203 (N_2203,N_936,N_546);
nand U2204 (N_2204,N_185,N_432);
and U2205 (N_2205,N_1419,N_11);
or U2206 (N_2206,N_1746,N_218);
nor U2207 (N_2207,N_1728,N_511);
and U2208 (N_2208,N_645,N_611);
nand U2209 (N_2209,N_470,N_175);
and U2210 (N_2210,N_1382,N_1155);
nor U2211 (N_2211,N_262,N_180);
or U2212 (N_2212,N_1168,N_1896);
or U2213 (N_2213,N_1886,N_610);
and U2214 (N_2214,N_1947,N_1118);
xor U2215 (N_2215,N_1444,N_162);
and U2216 (N_2216,N_1070,N_1851);
nor U2217 (N_2217,N_217,N_1953);
nand U2218 (N_2218,N_1499,N_314);
or U2219 (N_2219,N_1937,N_1629);
and U2220 (N_2220,N_1756,N_71);
and U2221 (N_2221,N_1922,N_918);
and U2222 (N_2222,N_653,N_331);
or U2223 (N_2223,N_333,N_1743);
or U2224 (N_2224,N_1995,N_128);
nand U2225 (N_2225,N_1111,N_373);
or U2226 (N_2226,N_209,N_517);
nand U2227 (N_2227,N_1214,N_1691);
xor U2228 (N_2228,N_694,N_733);
and U2229 (N_2229,N_112,N_86);
or U2230 (N_2230,N_1943,N_1511);
and U2231 (N_2231,N_1080,N_1520);
and U2232 (N_2232,N_1643,N_952);
or U2233 (N_2233,N_1106,N_229);
nand U2234 (N_2234,N_958,N_545);
and U2235 (N_2235,N_1400,N_1536);
or U2236 (N_2236,N_1175,N_1987);
nor U2237 (N_2237,N_156,N_971);
nand U2238 (N_2238,N_844,N_927);
and U2239 (N_2239,N_1702,N_864);
or U2240 (N_2240,N_1186,N_444);
and U2241 (N_2241,N_953,N_709);
nor U2242 (N_2242,N_407,N_435);
nand U2243 (N_2243,N_999,N_1861);
nor U2244 (N_2244,N_1219,N_969);
nand U2245 (N_2245,N_1171,N_1626);
xor U2246 (N_2246,N_681,N_509);
and U2247 (N_2247,N_1029,N_121);
and U2248 (N_2248,N_1173,N_1748);
nor U2249 (N_2249,N_863,N_386);
nand U2250 (N_2250,N_1674,N_943);
nand U2251 (N_2251,N_1397,N_1704);
and U2252 (N_2252,N_613,N_361);
and U2253 (N_2253,N_337,N_1486);
nor U2254 (N_2254,N_1303,N_1251);
nand U2255 (N_2255,N_1150,N_1983);
or U2256 (N_2256,N_1313,N_1194);
nor U2257 (N_2257,N_1469,N_74);
or U2258 (N_2258,N_1263,N_1038);
nand U2259 (N_2259,N_1013,N_1225);
nand U2260 (N_2260,N_1865,N_457);
and U2261 (N_2261,N_415,N_1061);
or U2262 (N_2262,N_934,N_370);
and U2263 (N_2263,N_791,N_1793);
or U2264 (N_2264,N_1271,N_1571);
or U2265 (N_2265,N_532,N_973);
nand U2266 (N_2266,N_1727,N_1291);
nor U2267 (N_2267,N_323,N_475);
nand U2268 (N_2268,N_1457,N_73);
xor U2269 (N_2269,N_652,N_513);
or U2270 (N_2270,N_297,N_1623);
xor U2271 (N_2271,N_1380,N_45);
nor U2272 (N_2272,N_1695,N_181);
or U2273 (N_2273,N_1445,N_1849);
nand U2274 (N_2274,N_1894,N_47);
and U2275 (N_2275,N_78,N_280);
nor U2276 (N_2276,N_1461,N_1063);
and U2277 (N_2277,N_1289,N_1754);
nand U2278 (N_2278,N_1374,N_287);
or U2279 (N_2279,N_917,N_1167);
nor U2280 (N_2280,N_1708,N_766);
and U2281 (N_2281,N_1796,N_325);
nand U2282 (N_2282,N_1744,N_89);
nand U2283 (N_2283,N_1151,N_234);
or U2284 (N_2284,N_753,N_1363);
or U2285 (N_2285,N_1483,N_802);
nand U2286 (N_2286,N_1532,N_1973);
nor U2287 (N_2287,N_270,N_302);
or U2288 (N_2288,N_1343,N_566);
and U2289 (N_2289,N_996,N_1810);
and U2290 (N_2290,N_604,N_640);
or U2291 (N_2291,N_607,N_26);
nand U2292 (N_2292,N_1561,N_810);
nand U2293 (N_2293,N_1964,N_834);
nand U2294 (N_2294,N_393,N_854);
or U2295 (N_2295,N_1677,N_1915);
and U2296 (N_2296,N_682,N_439);
and U2297 (N_2297,N_1527,N_436);
and U2298 (N_2298,N_576,N_1284);
nor U2299 (N_2299,N_205,N_1656);
or U2300 (N_2300,N_1350,N_1553);
and U2301 (N_2301,N_1911,N_1045);
or U2302 (N_2302,N_1847,N_1985);
xnor U2303 (N_2303,N_233,N_1309);
nand U2304 (N_2304,N_446,N_340);
and U2305 (N_2305,N_1965,N_1531);
or U2306 (N_2306,N_347,N_585);
and U2307 (N_2307,N_855,N_451);
nand U2308 (N_2308,N_1021,N_1948);
and U2309 (N_2309,N_1633,N_322);
and U2310 (N_2310,N_723,N_21);
nor U2311 (N_2311,N_497,N_25);
nor U2312 (N_2312,N_1514,N_504);
or U2313 (N_2313,N_1930,N_1613);
nor U2314 (N_2314,N_2,N_1838);
nand U2315 (N_2315,N_1588,N_176);
nor U2316 (N_2316,N_1928,N_720);
and U2317 (N_2317,N_1320,N_792);
or U2318 (N_2318,N_284,N_41);
or U2319 (N_2319,N_1729,N_414);
and U2320 (N_2320,N_1076,N_27);
nand U2321 (N_2321,N_247,N_93);
nor U2322 (N_2322,N_1997,N_1834);
and U2323 (N_2323,N_754,N_165);
nand U2324 (N_2324,N_1142,N_1906);
nor U2325 (N_2325,N_289,N_1630);
xor U2326 (N_2326,N_1693,N_955);
nor U2327 (N_2327,N_8,N_1485);
nand U2328 (N_2328,N_1425,N_215);
or U2329 (N_2329,N_839,N_430);
nand U2330 (N_2330,N_240,N_15);
nor U2331 (N_2331,N_1524,N_1249);
nor U2332 (N_2332,N_1700,N_658);
or U2333 (N_2333,N_1256,N_523);
nand U2334 (N_2334,N_1345,N_1898);
or U2335 (N_2335,N_484,N_327);
nor U2336 (N_2336,N_206,N_1152);
and U2337 (N_2337,N_1684,N_1405);
and U2338 (N_2338,N_1768,N_892);
and U2339 (N_2339,N_1083,N_1047);
or U2340 (N_2340,N_1717,N_132);
or U2341 (N_2341,N_19,N_741);
and U2342 (N_2342,N_813,N_821);
nand U2343 (N_2343,N_251,N_1238);
and U2344 (N_2344,N_677,N_1639);
nand U2345 (N_2345,N_670,N_116);
or U2346 (N_2346,N_804,N_914);
nand U2347 (N_2347,N_620,N_1722);
or U2348 (N_2348,N_931,N_1971);
nor U2349 (N_2349,N_945,N_129);
or U2350 (N_2350,N_152,N_963);
nor U2351 (N_2351,N_1191,N_883);
and U2352 (N_2352,N_1248,N_932);
nand U2353 (N_2353,N_136,N_109);
or U2354 (N_2354,N_1897,N_1940);
and U2355 (N_2355,N_1075,N_1113);
or U2356 (N_2356,N_476,N_940);
or U2357 (N_2357,N_157,N_888);
or U2358 (N_2358,N_1660,N_1705);
or U2359 (N_2359,N_70,N_900);
or U2360 (N_2360,N_335,N_1369);
nand U2361 (N_2361,N_184,N_1742);
nor U2362 (N_2362,N_1162,N_1891);
or U2363 (N_2363,N_4,N_1655);
or U2364 (N_2364,N_339,N_1330);
nand U2365 (N_2365,N_1907,N_1931);
nor U2366 (N_2366,N_1719,N_575);
and U2367 (N_2367,N_651,N_1523);
nor U2368 (N_2368,N_837,N_273);
nor U2369 (N_2369,N_125,N_1159);
nand U2370 (N_2370,N_1539,N_1678);
or U2371 (N_2371,N_507,N_867);
nand U2372 (N_2372,N_1817,N_979);
and U2373 (N_2373,N_1502,N_12);
nor U2374 (N_2374,N_1610,N_46);
and U2375 (N_2375,N_657,N_219);
and U2376 (N_2376,N_345,N_1308);
nand U2377 (N_2377,N_1143,N_732);
and U2378 (N_2378,N_1226,N_1352);
nand U2379 (N_2379,N_1122,N_1286);
nand U2380 (N_2380,N_1460,N_395);
nor U2381 (N_2381,N_362,N_530);
and U2382 (N_2382,N_959,N_643);
and U2383 (N_2383,N_1144,N_1044);
nor U2384 (N_2384,N_53,N_1581);
or U2385 (N_2385,N_572,N_593);
or U2386 (N_2386,N_376,N_521);
or U2387 (N_2387,N_294,N_695);
or U2388 (N_2388,N_1732,N_1560);
nor U2389 (N_2389,N_381,N_661);
nor U2390 (N_2390,N_1337,N_897);
or U2391 (N_2391,N_629,N_143);
nor U2392 (N_2392,N_1266,N_394);
or U2393 (N_2393,N_1407,N_293);
and U2394 (N_2394,N_150,N_269);
nor U2395 (N_2395,N_1145,N_1779);
nor U2396 (N_2396,N_997,N_126);
or U2397 (N_2397,N_904,N_1736);
and U2398 (N_2398,N_499,N_1148);
or U2399 (N_2399,N_1218,N_1815);
xnor U2400 (N_2400,N_1014,N_1333);
nor U2401 (N_2401,N_369,N_1384);
and U2402 (N_2402,N_1751,N_236);
or U2403 (N_2403,N_194,N_1784);
and U2404 (N_2404,N_304,N_1467);
nand U2405 (N_2405,N_1525,N_1652);
nand U2406 (N_2406,N_1355,N_385);
or U2407 (N_2407,N_1254,N_1449);
nor U2408 (N_2408,N_1945,N_104);
and U2409 (N_2409,N_1946,N_1517);
nand U2410 (N_2410,N_1758,N_313);
nor U2411 (N_2411,N_76,N_1814);
nor U2412 (N_2412,N_765,N_836);
and U2413 (N_2413,N_718,N_841);
xor U2414 (N_2414,N_988,N_1875);
or U2415 (N_2415,N_950,N_801);
nor U2416 (N_2416,N_1034,N_248);
and U2417 (N_2417,N_1665,N_1128);
nand U2418 (N_2418,N_1341,N_760);
and U2419 (N_2419,N_1362,N_691);
and U2420 (N_2420,N_1509,N_510);
nand U2421 (N_2421,N_231,N_537);
and U2422 (N_2422,N_747,N_909);
nor U2423 (N_2423,N_769,N_1205);
or U2424 (N_2424,N_416,N_992);
or U2425 (N_2425,N_1429,N_1278);
nor U2426 (N_2426,N_492,N_590);
or U2427 (N_2427,N_1269,N_1554);
nand U2428 (N_2428,N_1903,N_1319);
and U2429 (N_2429,N_1867,N_1206);
nor U2430 (N_2430,N_748,N_1839);
nand U2431 (N_2431,N_1545,N_1670);
nor U2432 (N_2432,N_1210,N_1878);
and U2433 (N_2433,N_707,N_1900);
nor U2434 (N_2434,N_1544,N_1889);
or U2435 (N_2435,N_533,N_946);
nand U2436 (N_2436,N_820,N_204);
and U2437 (N_2437,N_1636,N_851);
and U2438 (N_2438,N_478,N_1005);
nand U2439 (N_2439,N_1476,N_1566);
nand U2440 (N_2440,N_1353,N_466);
nand U2441 (N_2441,N_1316,N_1055);
nand U2442 (N_2442,N_420,N_255);
or U2443 (N_2443,N_110,N_1919);
or U2444 (N_2444,N_232,N_1427);
and U2445 (N_2445,N_1912,N_1935);
nand U2446 (N_2446,N_712,N_1770);
or U2447 (N_2447,N_227,N_1576);
and U2448 (N_2448,N_1526,N_1608);
and U2449 (N_2449,N_1280,N_1039);
or U2450 (N_2450,N_37,N_1074);
and U2451 (N_2451,N_698,N_472);
nand U2452 (N_2452,N_697,N_1923);
and U2453 (N_2453,N_1651,N_1595);
nor U2454 (N_2454,N_1887,N_1698);
nand U2455 (N_2455,N_423,N_1563);
or U2456 (N_2456,N_1050,N_846);
and U2457 (N_2457,N_1567,N_408);
or U2458 (N_2458,N_656,N_300);
nand U2459 (N_2459,N_1220,N_1422);
and U2460 (N_2460,N_551,N_998);
nor U2461 (N_2461,N_865,N_816);
nand U2462 (N_2462,N_1125,N_1791);
nand U2463 (N_2463,N_957,N_1515);
and U2464 (N_2464,N_967,N_1749);
and U2465 (N_2465,N_1549,N_1926);
nor U2466 (N_2466,N_1924,N_1325);
nand U2467 (N_2467,N_9,N_1568);
and U2468 (N_2468,N_1464,N_1864);
nor U2469 (N_2469,N_1163,N_1501);
xor U2470 (N_2470,N_727,N_1802);
nand U2471 (N_2471,N_1951,N_1274);
nor U2472 (N_2472,N_699,N_583);
nand U2473 (N_2473,N_543,N_1109);
and U2474 (N_2474,N_1988,N_127);
or U2475 (N_2475,N_428,N_878);
nor U2476 (N_2476,N_1466,N_274);
or U2477 (N_2477,N_1331,N_1120);
nor U2478 (N_2478,N_1135,N_1176);
and U2479 (N_2479,N_1241,N_994);
nand U2480 (N_2480,N_1016,N_1752);
and U2481 (N_2481,N_1836,N_1158);
nor U2482 (N_2482,N_456,N_1592);
nand U2483 (N_2483,N_818,N_1835);
and U2484 (N_2484,N_106,N_591);
and U2485 (N_2485,N_895,N_1593);
or U2486 (N_2486,N_554,N_1);
nand U2487 (N_2487,N_605,N_1202);
or U2488 (N_2488,N_137,N_692);
and U2489 (N_2489,N_1223,N_352);
nand U2490 (N_2490,N_498,N_413);
or U2491 (N_2491,N_1389,N_1012);
or U2492 (N_2492,N_1322,N_172);
nor U2493 (N_2493,N_1156,N_1820);
and U2494 (N_2494,N_159,N_987);
or U2495 (N_2495,N_1015,N_948);
or U2496 (N_2496,N_1417,N_1621);
nor U2497 (N_2497,N_1687,N_101);
and U2498 (N_2498,N_1679,N_730);
or U2499 (N_2499,N_1713,N_406);
xor U2500 (N_2500,N_1354,N_522);
nand U2501 (N_2501,N_147,N_860);
nand U2502 (N_2502,N_113,N_1324);
nand U2503 (N_2503,N_1431,N_1247);
nor U2504 (N_2504,N_256,N_1059);
nand U2505 (N_2505,N_555,N_1439);
or U2506 (N_2506,N_1958,N_1105);
and U2507 (N_2507,N_1979,N_1848);
and U2508 (N_2508,N_438,N_1573);
nor U2509 (N_2509,N_1590,N_64);
nand U2510 (N_2510,N_1963,N_48);
nor U2511 (N_2511,N_96,N_130);
or U2512 (N_2512,N_578,N_1797);
or U2513 (N_2513,N_1009,N_124);
nand U2514 (N_2514,N_696,N_858);
nand U2515 (N_2515,N_1688,N_1127);
nor U2516 (N_2516,N_1557,N_1780);
or U2517 (N_2517,N_662,N_58);
and U2518 (N_2518,N_1627,N_1583);
and U2519 (N_2519,N_1215,N_461);
nor U2520 (N_2520,N_283,N_1297);
and U2521 (N_2521,N_907,N_560);
nor U2522 (N_2522,N_1346,N_614);
and U2523 (N_2523,N_1496,N_1760);
nand U2524 (N_2524,N_1270,N_1481);
or U2525 (N_2525,N_597,N_744);
nor U2526 (N_2526,N_835,N_1090);
and U2527 (N_2527,N_639,N_1993);
nor U2528 (N_2528,N_1253,N_584);
or U2529 (N_2529,N_706,N_377);
or U2530 (N_2530,N_767,N_349);
nor U2531 (N_2531,N_803,N_763);
or U2532 (N_2532,N_853,N_738);
nand U2533 (N_2533,N_1671,N_196);
and U2534 (N_2534,N_398,N_419);
or U2535 (N_2535,N_1852,N_978);
or U2536 (N_2536,N_1709,N_100);
or U2537 (N_2537,N_704,N_1335);
nor U2538 (N_2538,N_1095,N_1195);
and U2539 (N_2539,N_965,N_726);
and U2540 (N_2540,N_1720,N_825);
nor U2541 (N_2541,N_1739,N_843);
nor U2542 (N_2542,N_711,N_1018);
and U2543 (N_2543,N_1412,N_228);
and U2544 (N_2544,N_540,N_1196);
and U2545 (N_2545,N_1383,N_23);
or U2546 (N_2546,N_81,N_1535);
nand U2547 (N_2547,N_1990,N_885);
nor U2548 (N_2548,N_896,N_974);
and U2549 (N_2549,N_1081,N_749);
nand U2550 (N_2550,N_1310,N_947);
and U2551 (N_2551,N_625,N_1371);
or U2552 (N_2552,N_1673,N_463);
nor U2553 (N_2553,N_149,N_1394);
and U2554 (N_2554,N_759,N_1858);
nand U2555 (N_2555,N_829,N_746);
and U2556 (N_2556,N_1487,N_1910);
nor U2557 (N_2557,N_1031,N_1141);
nand U2558 (N_2558,N_371,N_1606);
and U2559 (N_2559,N_1686,N_1312);
nor U2560 (N_2560,N_1904,N_1615);
or U2561 (N_2561,N_688,N_1041);
or U2562 (N_2562,N_1317,N_778);
nand U2563 (N_2563,N_1149,N_246);
nor U2564 (N_2564,N_770,N_1628);
or U2565 (N_2565,N_1596,N_462);
nand U2566 (N_2566,N_1551,N_1415);
and U2567 (N_2567,N_1154,N_984);
nand U2568 (N_2568,N_916,N_1216);
nor U2569 (N_2569,N_221,N_1209);
or U2570 (N_2570,N_684,N_1685);
nor U2571 (N_2571,N_243,N_1980);
nor U2572 (N_2572,N_1160,N_260);
and U2573 (N_2573,N_1733,N_1584);
nand U2574 (N_2574,N_177,N_115);
or U2575 (N_2575,N_1277,N_581);
or U2576 (N_2576,N_1349,N_1392);
nand U2577 (N_2577,N_482,N_1645);
nand U2578 (N_2578,N_225,N_1649);
nor U2579 (N_2579,N_1177,N_780);
nand U2580 (N_2580,N_241,N_1440);
nor U2581 (N_2581,N_1273,N_1200);
nand U2582 (N_2582,N_564,N_1552);
nand U2583 (N_2583,N_1666,N_824);
and U2584 (N_2584,N_1447,N_579);
or U2585 (N_2585,N_553,N_768);
nor U2586 (N_2586,N_1829,N_1315);
nand U2587 (N_2587,N_515,N_133);
nor U2588 (N_2588,N_148,N_1385);
nand U2589 (N_2589,N_1738,N_372);
nor U2590 (N_2590,N_731,N_736);
or U2591 (N_2591,N_453,N_57);
nand U2592 (N_2592,N_1019,N_636);
nor U2593 (N_2593,N_1654,N_1246);
nand U2594 (N_2594,N_311,N_72);
and U2595 (N_2595,N_1586,N_455);
and U2596 (N_2596,N_811,N_534);
or U2597 (N_2597,N_1787,N_1301);
nand U2598 (N_2598,N_798,N_467);
and U2599 (N_2599,N_1724,N_1730);
nand U2600 (N_2600,N_1917,N_1259);
and U2601 (N_2601,N_276,N_1116);
nand U2602 (N_2602,N_1424,N_1103);
or U2603 (N_2603,N_63,N_925);
or U2604 (N_2604,N_1999,N_1996);
nor U2605 (N_2605,N_574,N_542);
nor U2606 (N_2606,N_1185,N_794);
nand U2607 (N_2607,N_422,N_50);
or U2608 (N_2608,N_1650,N_90);
nor U2609 (N_2609,N_789,N_728);
nand U2610 (N_2610,N_1773,N_1555);
nand U2611 (N_2611,N_1540,N_1368);
and U2612 (N_2612,N_809,N_1828);
or U2613 (N_2613,N_877,N_1882);
xnor U2614 (N_2614,N_268,N_915);
nand U2615 (N_2615,N_756,N_717);
and U2616 (N_2616,N_207,N_1842);
nand U2617 (N_2617,N_1052,N_1792);
or U2618 (N_2618,N_646,N_582);
nand U2619 (N_2619,N_1747,N_906);
nor U2620 (N_2620,N_870,N_351);
nor U2621 (N_2621,N_40,N_1762);
nor U2622 (N_2622,N_1765,N_1644);
nor U2623 (N_2623,N_966,N_1420);
and U2624 (N_2624,N_153,N_536);
nor U2625 (N_2625,N_111,N_1876);
nand U2626 (N_2626,N_426,N_550);
and U2627 (N_2627,N_1459,N_396);
nor U2628 (N_2628,N_1955,N_1624);
and U2629 (N_2629,N_571,N_348);
nor U2630 (N_2630,N_265,N_145);
or U2631 (N_2631,N_495,N_1399);
or U2632 (N_2632,N_705,N_244);
nand U2633 (N_2633,N_826,N_797);
or U2634 (N_2634,N_1465,N_266);
or U2635 (N_2635,N_1564,N_1472);
nor U2636 (N_2636,N_679,N_454);
and U2637 (N_2637,N_1268,N_627);
nor U2638 (N_2638,N_1871,N_715);
nor U2639 (N_2639,N_1416,N_1373);
nor U2640 (N_2640,N_799,N_1856);
nand U2641 (N_2641,N_1410,N_344);
nand U2642 (N_2642,N_92,N_788);
nor U2643 (N_2643,N_34,N_1409);
or U2644 (N_2644,N_848,N_171);
or U2645 (N_2645,N_1288,N_1264);
and U2646 (N_2646,N_781,N_1916);
nand U2647 (N_2647,N_319,N_1604);
nor U2648 (N_2648,N_424,N_673);
nor U2649 (N_2649,N_928,N_1456);
nor U2650 (N_2650,N_123,N_1110);
nand U2651 (N_2651,N_832,N_1455);
nand U2652 (N_2652,N_935,N_301);
nand U2653 (N_2653,N_642,N_1710);
nand U2654 (N_2654,N_1351,N_903);
nand U2655 (N_2655,N_382,N_1283);
nand U2656 (N_2656,N_635,N_964);
and U2657 (N_2657,N_1920,N_1975);
and U2658 (N_2658,N_962,N_404);
nor U2659 (N_2659,N_1808,N_847);
or U2660 (N_2660,N_842,N_1795);
nand U2661 (N_2661,N_139,N_902);
or U2662 (N_2662,N_296,N_1777);
or U2663 (N_2663,N_680,N_190);
nand U2664 (N_2664,N_1811,N_1764);
and U2665 (N_2665,N_279,N_1179);
and U2666 (N_2666,N_1078,N_1418);
xor U2667 (N_2667,N_1197,N_1441);
xnor U2668 (N_2668,N_743,N_529);
and U2669 (N_2669,N_561,N_787);
nand U2670 (N_2670,N_450,N_1631);
and U2671 (N_2671,N_1478,N_1800);
nand U2672 (N_2672,N_1471,N_722);
nand U2673 (N_2673,N_1740,N_6);
xor U2674 (N_2674,N_1184,N_1058);
or U2675 (N_2675,N_976,N_721);
and U2676 (N_2676,N_1715,N_1296);
and U2677 (N_2677,N_399,N_687);
and U2678 (N_2678,N_592,N_674);
or U2679 (N_2679,N_1597,N_538);
nor U2680 (N_2680,N_479,N_624);
and U2681 (N_2681,N_734,N_108);
or U2682 (N_2682,N_1601,N_1032);
nand U2683 (N_2683,N_608,N_856);
nor U2684 (N_2684,N_1401,N_880);
nor U2685 (N_2685,N_1694,N_310);
and U2686 (N_2686,N_308,N_82);
and U2687 (N_2687,N_1869,N_1612);
nor U2688 (N_2688,N_650,N_1002);
or U2689 (N_2689,N_771,N_857);
nor U2690 (N_2690,N_1243,N_1323);
and U2691 (N_2691,N_776,N_441);
or U2692 (N_2692,N_68,N_1262);
xnor U2693 (N_2693,N_596,N_1236);
and U2694 (N_2694,N_1794,N_392);
or U2695 (N_2695,N_360,N_189);
nand U2696 (N_2696,N_66,N_1825);
and U2697 (N_2697,N_1126,N_622);
or U2698 (N_2698,N_1783,N_199);
and U2699 (N_2699,N_1609,N_619);
or U2700 (N_2700,N_80,N_926);
nor U2701 (N_2701,N_1421,N_899);
nor U2702 (N_2702,N_1170,N_35);
and U2703 (N_2703,N_166,N_1172);
and U2704 (N_2704,N_1146,N_1909);
and U2705 (N_2705,N_212,N_405);
and U2706 (N_2706,N_1379,N_1620);
nor U2707 (N_2707,N_1051,N_1027);
nor U2708 (N_2708,N_812,N_1402);
nand U2709 (N_2709,N_1913,N_637);
nand U2710 (N_2710,N_1007,N_155);
nand U2711 (N_2711,N_1589,N_548);
and U2712 (N_2712,N_1451,N_1211);
nand U2713 (N_2713,N_1065,N_1366);
nand U2714 (N_2714,N_866,N_1121);
or U2715 (N_2715,N_615,N_1321);
and U2716 (N_2716,N_1813,N_1484);
and U2717 (N_2717,N_621,N_1723);
and U2718 (N_2718,N_1056,N_1443);
and U2719 (N_2719,N_514,N_1279);
and U2720 (N_2720,N_905,N_1498);
nand U2721 (N_2721,N_1183,N_1803);
or U2722 (N_2722,N_648,N_1049);
nand U2723 (N_2723,N_32,N_411);
nand U2724 (N_2724,N_1326,N_375);
nor U2725 (N_2725,N_254,N_1942);
and U2726 (N_2726,N_1711,N_140);
and U2727 (N_2727,N_51,N_1984);
nand U2728 (N_2728,N_1231,N_800);
or U2729 (N_2729,N_1119,N_135);
nor U2730 (N_2730,N_954,N_887);
nor U2731 (N_2731,N_39,N_1101);
and U2732 (N_2732,N_577,N_869);
nand U2733 (N_2733,N_183,N_881);
nand U2734 (N_2734,N_1731,N_91);
and U2735 (N_2735,N_329,N_570);
nand U2736 (N_2736,N_24,N_1994);
and U2737 (N_2737,N_777,N_1962);
and U2738 (N_2738,N_114,N_1448);
nand U2739 (N_2739,N_1681,N_496);
and U2740 (N_2740,N_1822,N_486);
nor U2741 (N_2741,N_338,N_1895);
or U2742 (N_2742,N_387,N_88);
nand U2743 (N_2743,N_1862,N_1755);
and U2744 (N_2744,N_1187,N_374);
or U2745 (N_2745,N_942,N_1598);
nor U2746 (N_2746,N_427,N_242);
or U2747 (N_2747,N_1941,N_429);
nor U2748 (N_2748,N_1257,N_528);
nor U2749 (N_2749,N_690,N_1040);
nor U2750 (N_2750,N_418,N_1821);
or U2751 (N_2751,N_1138,N_859);
nand U2752 (N_2752,N_961,N_42);
or U2753 (N_2753,N_1830,N_1991);
or U2754 (N_2754,N_1198,N_1788);
and U2755 (N_2755,N_257,N_1519);
or U2756 (N_2756,N_1547,N_1938);
or U2757 (N_2757,N_1837,N_258);
nand U2758 (N_2758,N_160,N_54);
and U2759 (N_2759,N_1692,N_1166);
xnor U2760 (N_2760,N_460,N_891);
or U2761 (N_2761,N_1426,N_1411);
nor U2762 (N_2762,N_1949,N_1661);
xnor U2763 (N_2763,N_170,N_796);
or U2764 (N_2764,N_1406,N_1763);
nand U2765 (N_2765,N_1503,N_417);
nor U2766 (N_2766,N_230,N_1981);
nand U2767 (N_2767,N_356,N_1505);
or U2768 (N_2768,N_1304,N_62);
and U2769 (N_2769,N_930,N_1591);
xnor U2770 (N_2770,N_549,N_1559);
nand U2771 (N_2771,N_1193,N_1932);
nand U2772 (N_2772,N_1619,N_1347);
or U2773 (N_2773,N_742,N_493);
and U2774 (N_2774,N_328,N_1386);
nand U2775 (N_2775,N_1178,N_14);
and U2776 (N_2776,N_758,N_1132);
nand U2777 (N_2777,N_163,N_833);
nand U2778 (N_2778,N_1516,N_1863);
and U2779 (N_2779,N_107,N_173);
and U2780 (N_2780,N_676,N_1494);
xnor U2781 (N_2781,N_61,N_647);
or U2782 (N_2782,N_1759,N_773);
nor U2783 (N_2783,N_5,N_52);
nand U2784 (N_2784,N_307,N_1992);
nor U2785 (N_2785,N_786,N_1396);
and U2786 (N_2786,N_421,N_409);
nor U2787 (N_2787,N_1541,N_1099);
and U2788 (N_2788,N_1798,N_1675);
and U2789 (N_2789,N_603,N_1676);
and U2790 (N_2790,N_518,N_437);
or U2791 (N_2791,N_1260,N_336);
nor U2792 (N_2792,N_1543,N_745);
nor U2793 (N_2793,N_1577,N_1844);
nand U2794 (N_2794,N_667,N_588);
or U2795 (N_2795,N_1388,N_250);
xnor U2796 (N_2796,N_402,N_292);
nor U2797 (N_2797,N_1468,N_1491);
or U2798 (N_2798,N_1934,N_317);
nor U2799 (N_2799,N_28,N_77);
or U2800 (N_2800,N_1575,N_343);
nand U2801 (N_2801,N_580,N_1348);
or U2802 (N_2802,N_1188,N_367);
and U2803 (N_2803,N_410,N_1446);
and U2804 (N_2804,N_913,N_1790);
and U2805 (N_2805,N_473,N_431);
nor U2806 (N_2806,N_1603,N_1605);
and U2807 (N_2807,N_1042,N_1580);
nand U2808 (N_2808,N_868,N_1510);
and U2809 (N_2809,N_1482,N_1950);
or U2810 (N_2810,N_1275,N_526);
xor U2811 (N_2811,N_1053,N_1816);
and U2812 (N_2812,N_1680,N_263);
nor U2813 (N_2813,N_1230,N_38);
nor U2814 (N_2814,N_1497,N_264);
and U2815 (N_2815,N_1853,N_1046);
nand U2816 (N_2816,N_16,N_275);
nand U2817 (N_2817,N_363,N_1026);
and U2818 (N_2818,N_1672,N_103);
nor U2819 (N_2819,N_1761,N_1336);
or U2820 (N_2820,N_761,N_1998);
nand U2821 (N_2821,N_1558,N_599);
and U2822 (N_2822,N_949,N_191);
and U2823 (N_2823,N_1769,N_725);
or U2824 (N_2824,N_1217,N_389);
and U2825 (N_2825,N_617,N_638);
nand U2826 (N_2826,N_762,N_1647);
nand U2827 (N_2827,N_1017,N_1599);
or U2828 (N_2828,N_547,N_1028);
nand U2829 (N_2829,N_1001,N_1617);
xor U2830 (N_2830,N_1438,N_793);
nand U2831 (N_2831,N_253,N_445);
and U2832 (N_2832,N_1147,N_79);
or U2833 (N_2833,N_95,N_1035);
nand U2834 (N_2834,N_403,N_1884);
nand U2835 (N_2835,N_29,N_557);
nand U2836 (N_2836,N_1569,N_67);
or U2837 (N_2837,N_1292,N_1936);
nand U2838 (N_2838,N_378,N_586);
xnor U2839 (N_2839,N_1043,N_474);
and U2840 (N_2840,N_539,N_1091);
nand U2841 (N_2841,N_531,N_1123);
nor U2842 (N_2842,N_1318,N_220);
xor U2843 (N_2843,N_443,N_595);
and U2844 (N_2844,N_1329,N_1089);
nor U2845 (N_2845,N_169,N_669);
and U2846 (N_2846,N_1726,N_1357);
nand U2847 (N_2847,N_1365,N_1513);
and U2848 (N_2848,N_1376,N_1239);
nor U2849 (N_2849,N_357,N_991);
nor U2850 (N_2850,N_602,N_488);
and U2851 (N_2851,N_1521,N_85);
nor U2852 (N_2852,N_1735,N_506);
or U2853 (N_2853,N_245,N_516);
nand U2854 (N_2854,N_201,N_354);
and U2855 (N_2855,N_1377,N_1638);
and U2856 (N_2856,N_1548,N_1030);
and U2857 (N_2857,N_1124,N_751);
or U2858 (N_2858,N_480,N_562);
nand U2859 (N_2859,N_1104,N_1344);
or U2860 (N_2860,N_1893,N_1287);
nor U2861 (N_2861,N_1982,N_1437);
and U2862 (N_2862,N_1182,N_1618);
or U2863 (N_2863,N_729,N_1860);
and U2864 (N_2864,N_1572,N_1340);
nand U2865 (N_2865,N_364,N_1880);
and U2866 (N_2866,N_1442,N_1293);
and U2867 (N_2867,N_22,N_18);
nand U2868 (N_2868,N_1115,N_815);
nor U2869 (N_2869,N_512,N_1000);
and U2870 (N_2870,N_1578,N_1925);
xnor U2871 (N_2871,N_1024,N_1986);
nand U2872 (N_2872,N_211,N_1334);
or U2873 (N_2873,N_1066,N_1370);
and U2874 (N_2874,N_1757,N_390);
nor U2875 (N_2875,N_1240,N_689);
nor U2876 (N_2876,N_1632,N_299);
or U2877 (N_2877,N_1338,N_939);
nand U2878 (N_2878,N_1801,N_1096);
nand U2879 (N_2879,N_1189,N_179);
and U2880 (N_2880,N_628,N_401);
nand U2881 (N_2881,N_1682,N_982);
nand U2882 (N_2882,N_1398,N_1364);
and U2883 (N_2883,N_633,N_1463);
nor U2884 (N_2884,N_1153,N_49);
and U2885 (N_2885,N_1976,N_849);
or U2886 (N_2886,N_1927,N_664);
nor U2887 (N_2887,N_1699,N_525);
and U2888 (N_2888,N_142,N_1522);
nor U2889 (N_2889,N_956,N_1022);
nand U2890 (N_2890,N_286,N_1475);
and U2891 (N_2891,N_1234,N_198);
nand U2892 (N_2892,N_1190,N_174);
and U2893 (N_2893,N_1782,N_1285);
nor U2894 (N_2894,N_1667,N_960);
or U2895 (N_2895,N_1512,N_1668);
and U2896 (N_2896,N_1192,N_589);
nand U2897 (N_2897,N_1372,N_1072);
nor U2898 (N_2898,N_912,N_1060);
nand U2899 (N_2899,N_875,N_1832);
nand U2900 (N_2900,N_1093,N_83);
nand U2901 (N_2901,N_1010,N_65);
or U2902 (N_2902,N_490,N_1537);
nor U2903 (N_2903,N_489,N_772);
nand U2904 (N_2904,N_1799,N_1164);
or U2905 (N_2905,N_397,N_981);
and U2906 (N_2906,N_1229,N_1356);
nand U2907 (N_2907,N_1435,N_501);
nor U2908 (N_2908,N_1133,N_84);
or U2909 (N_2909,N_1741,N_830);
nand U2910 (N_2910,N_807,N_784);
nor U2911 (N_2911,N_618,N_929);
nand U2912 (N_2912,N_272,N_1776);
and U2913 (N_2913,N_1174,N_1614);
nand U2914 (N_2914,N_1778,N_922);
nor U2915 (N_2915,N_898,N_938);
and U2916 (N_2916,N_519,N_1328);
or U2917 (N_2917,N_56,N_365);
and U2918 (N_2918,N_1008,N_703);
or U2919 (N_2919,N_1267,N_213);
nand U2920 (N_2920,N_1721,N_1818);
xor U2921 (N_2921,N_1888,N_1033);
nor U2922 (N_2922,N_1960,N_306);
or U2923 (N_2923,N_1255,N_1433);
nor U2924 (N_2924,N_1767,N_1332);
or U2925 (N_2925,N_69,N_831);
and U2926 (N_2926,N_192,N_1139);
nand U2927 (N_2927,N_1939,N_924);
nor U2928 (N_2928,N_282,N_1812);
and U2929 (N_2929,N_1616,N_654);
and U2930 (N_2930,N_937,N_1180);
nor U2931 (N_2931,N_675,N_154);
or U2932 (N_2932,N_1528,N_1117);
nor U2933 (N_2933,N_861,N_182);
or U2934 (N_2934,N_1556,N_1587);
or U2935 (N_2935,N_214,N_1071);
nor U2936 (N_2936,N_502,N_259);
nand U2937 (N_2937,N_764,N_167);
nor U2938 (N_2938,N_1664,N_134);
nor U2939 (N_2939,N_1359,N_278);
nand U2940 (N_2940,N_200,N_1646);
and U2941 (N_2941,N_980,N_31);
and U2942 (N_2942,N_1737,N_862);
nand U2943 (N_2943,N_1479,N_346);
nand U2944 (N_2944,N_97,N_1474);
and U2945 (N_2945,N_355,N_1227);
or U2946 (N_2946,N_485,N_118);
or U2947 (N_2947,N_1258,N_1136);
nor U2948 (N_2948,N_1228,N_1642);
nand U2949 (N_2949,N_1069,N_544);
nor U2950 (N_2950,N_790,N_1972);
nor U2951 (N_2951,N_36,N_828);
nor U2952 (N_2952,N_326,N_1594);
or U2953 (N_2953,N_105,N_1714);
and U2954 (N_2954,N_1221,N_685);
and U2955 (N_2955,N_783,N_827);
nand U2956 (N_2956,N_631,N_1774);
nand U2957 (N_2957,N_1358,N_1003);
and U2958 (N_2958,N_120,N_178);
nand U2959 (N_2959,N_433,N_951);
or U2960 (N_2960,N_1314,N_630);
nor U2961 (N_2961,N_1020,N_1753);
nand U2962 (N_2962,N_819,N_678);
nand U2963 (N_2963,N_700,N_1707);
nor U2964 (N_2964,N_239,N_158);
nor U2965 (N_2965,N_1546,N_0);
nor U2966 (N_2966,N_330,N_1833);
nor U2967 (N_2967,N_458,N_719);
or U2968 (N_2968,N_985,N_1130);
and U2969 (N_2969,N_1213,N_686);
and U2970 (N_2970,N_1890,N_941);
nor U2971 (N_2971,N_1804,N_840);
nand U2972 (N_2972,N_203,N_701);
or U2973 (N_2973,N_471,N_459);
nor U2974 (N_2974,N_224,N_1390);
nor U2975 (N_2975,N_1824,N_1381);
or U2976 (N_2976,N_131,N_1092);
and U2977 (N_2977,N_1169,N_1533);
and U2978 (N_2978,N_17,N_379);
or U2979 (N_2979,N_659,N_1272);
nand U2980 (N_2980,N_1023,N_1585);
nand U2981 (N_2981,N_447,N_1970);
or U2982 (N_2982,N_1212,N_1622);
or U2983 (N_2983,N_1112,N_1967);
nor U2984 (N_2984,N_3,N_13);
nand U2985 (N_2985,N_1716,N_1508);
and U2986 (N_2986,N_1207,N_921);
or U2987 (N_2987,N_671,N_852);
nand U2988 (N_2988,N_1807,N_872);
and U2989 (N_2989,N_1872,N_1094);
or U2990 (N_2990,N_850,N_1806);
nor U2991 (N_2991,N_138,N_290);
and U2992 (N_2992,N_1866,N_1393);
nand U2993 (N_2993,N_309,N_487);
and U2994 (N_2994,N_672,N_567);
nor U2995 (N_2995,N_1879,N_710);
and U2996 (N_2996,N_1299,N_94);
or U2997 (N_2997,N_1157,N_1204);
nand U2998 (N_2998,N_1989,N_1745);
nor U2999 (N_2999,N_1079,N_1203);
nand U3000 (N_3000,N_600,N_11);
and U3001 (N_3001,N_1822,N_1612);
or U3002 (N_3002,N_830,N_931);
and U3003 (N_3003,N_702,N_1938);
nand U3004 (N_3004,N_1293,N_580);
xnor U3005 (N_3005,N_525,N_148);
and U3006 (N_3006,N_948,N_1229);
or U3007 (N_3007,N_152,N_1174);
nor U3008 (N_3008,N_399,N_1573);
or U3009 (N_3009,N_1620,N_100);
nor U3010 (N_3010,N_630,N_788);
nor U3011 (N_3011,N_102,N_940);
nor U3012 (N_3012,N_1722,N_1159);
and U3013 (N_3013,N_486,N_1652);
nor U3014 (N_3014,N_204,N_948);
or U3015 (N_3015,N_823,N_1240);
and U3016 (N_3016,N_699,N_1215);
nor U3017 (N_3017,N_929,N_1874);
and U3018 (N_3018,N_1694,N_636);
and U3019 (N_3019,N_296,N_1601);
nand U3020 (N_3020,N_110,N_28);
or U3021 (N_3021,N_1281,N_862);
nor U3022 (N_3022,N_1813,N_1350);
and U3023 (N_3023,N_1693,N_1354);
or U3024 (N_3024,N_1314,N_1002);
nor U3025 (N_3025,N_728,N_1007);
or U3026 (N_3026,N_26,N_1978);
nand U3027 (N_3027,N_1809,N_567);
nand U3028 (N_3028,N_71,N_19);
and U3029 (N_3029,N_1312,N_487);
or U3030 (N_3030,N_1311,N_321);
and U3031 (N_3031,N_37,N_1193);
nor U3032 (N_3032,N_52,N_964);
and U3033 (N_3033,N_1627,N_1452);
or U3034 (N_3034,N_1156,N_917);
nor U3035 (N_3035,N_1501,N_1776);
or U3036 (N_3036,N_889,N_743);
or U3037 (N_3037,N_75,N_1853);
nand U3038 (N_3038,N_1296,N_1963);
nand U3039 (N_3039,N_1133,N_1609);
and U3040 (N_3040,N_1192,N_1285);
nor U3041 (N_3041,N_712,N_1124);
or U3042 (N_3042,N_731,N_922);
nor U3043 (N_3043,N_817,N_0);
or U3044 (N_3044,N_703,N_1056);
or U3045 (N_3045,N_604,N_1730);
nand U3046 (N_3046,N_161,N_721);
nand U3047 (N_3047,N_1816,N_253);
nand U3048 (N_3048,N_1502,N_64);
xnor U3049 (N_3049,N_265,N_284);
or U3050 (N_3050,N_677,N_256);
nand U3051 (N_3051,N_1250,N_108);
nand U3052 (N_3052,N_1049,N_962);
nand U3053 (N_3053,N_1413,N_1365);
and U3054 (N_3054,N_1052,N_99);
and U3055 (N_3055,N_1069,N_1049);
or U3056 (N_3056,N_134,N_453);
nand U3057 (N_3057,N_1671,N_1924);
nor U3058 (N_3058,N_428,N_168);
nor U3059 (N_3059,N_550,N_1152);
nor U3060 (N_3060,N_704,N_700);
or U3061 (N_3061,N_211,N_1069);
xor U3062 (N_3062,N_689,N_88);
nand U3063 (N_3063,N_552,N_1039);
nor U3064 (N_3064,N_421,N_1330);
nor U3065 (N_3065,N_242,N_1403);
nand U3066 (N_3066,N_644,N_1610);
xor U3067 (N_3067,N_1749,N_843);
and U3068 (N_3068,N_1704,N_133);
nor U3069 (N_3069,N_902,N_853);
nand U3070 (N_3070,N_220,N_1690);
or U3071 (N_3071,N_306,N_720);
nor U3072 (N_3072,N_594,N_657);
or U3073 (N_3073,N_1825,N_483);
nor U3074 (N_3074,N_1140,N_411);
nor U3075 (N_3075,N_1835,N_556);
or U3076 (N_3076,N_513,N_869);
and U3077 (N_3077,N_172,N_828);
and U3078 (N_3078,N_1848,N_1825);
nand U3079 (N_3079,N_1198,N_275);
nor U3080 (N_3080,N_1926,N_1302);
and U3081 (N_3081,N_1221,N_847);
nor U3082 (N_3082,N_894,N_1894);
nor U3083 (N_3083,N_694,N_1671);
and U3084 (N_3084,N_187,N_145);
or U3085 (N_3085,N_1378,N_1976);
or U3086 (N_3086,N_1357,N_677);
or U3087 (N_3087,N_1936,N_147);
or U3088 (N_3088,N_1556,N_1852);
nand U3089 (N_3089,N_1453,N_499);
or U3090 (N_3090,N_1021,N_1581);
and U3091 (N_3091,N_886,N_1355);
or U3092 (N_3092,N_1758,N_1320);
and U3093 (N_3093,N_1510,N_757);
nand U3094 (N_3094,N_1721,N_176);
nor U3095 (N_3095,N_1603,N_1704);
nor U3096 (N_3096,N_1582,N_1060);
nand U3097 (N_3097,N_220,N_1754);
or U3098 (N_3098,N_470,N_1353);
nand U3099 (N_3099,N_889,N_1708);
nor U3100 (N_3100,N_972,N_114);
nand U3101 (N_3101,N_377,N_1004);
nand U3102 (N_3102,N_784,N_1163);
nor U3103 (N_3103,N_1930,N_63);
nand U3104 (N_3104,N_21,N_1920);
nor U3105 (N_3105,N_1977,N_1601);
nor U3106 (N_3106,N_1561,N_1034);
and U3107 (N_3107,N_519,N_652);
xnor U3108 (N_3108,N_715,N_744);
nor U3109 (N_3109,N_843,N_1571);
and U3110 (N_3110,N_665,N_992);
and U3111 (N_3111,N_480,N_1071);
nand U3112 (N_3112,N_925,N_311);
nor U3113 (N_3113,N_991,N_1750);
or U3114 (N_3114,N_1377,N_585);
or U3115 (N_3115,N_1328,N_1746);
nor U3116 (N_3116,N_619,N_110);
nor U3117 (N_3117,N_1438,N_1255);
nor U3118 (N_3118,N_1487,N_1028);
and U3119 (N_3119,N_1763,N_1012);
nor U3120 (N_3120,N_1799,N_1722);
and U3121 (N_3121,N_772,N_310);
xor U3122 (N_3122,N_982,N_944);
nand U3123 (N_3123,N_1126,N_1344);
nor U3124 (N_3124,N_1692,N_155);
nand U3125 (N_3125,N_1906,N_1302);
xnor U3126 (N_3126,N_163,N_14);
xor U3127 (N_3127,N_1693,N_28);
nor U3128 (N_3128,N_647,N_1484);
or U3129 (N_3129,N_1912,N_1800);
or U3130 (N_3130,N_777,N_1468);
nor U3131 (N_3131,N_1431,N_1417);
and U3132 (N_3132,N_1411,N_1549);
nor U3133 (N_3133,N_1182,N_1120);
and U3134 (N_3134,N_1527,N_605);
or U3135 (N_3135,N_1084,N_72);
nor U3136 (N_3136,N_146,N_116);
nor U3137 (N_3137,N_1222,N_1277);
or U3138 (N_3138,N_736,N_1901);
nand U3139 (N_3139,N_1756,N_873);
or U3140 (N_3140,N_200,N_769);
or U3141 (N_3141,N_1168,N_452);
or U3142 (N_3142,N_131,N_1073);
or U3143 (N_3143,N_1030,N_1212);
nand U3144 (N_3144,N_955,N_1871);
nand U3145 (N_3145,N_848,N_823);
nor U3146 (N_3146,N_1723,N_1098);
nand U3147 (N_3147,N_1064,N_947);
or U3148 (N_3148,N_579,N_479);
or U3149 (N_3149,N_1497,N_1664);
nand U3150 (N_3150,N_1181,N_1070);
nand U3151 (N_3151,N_1886,N_687);
or U3152 (N_3152,N_301,N_1172);
nand U3153 (N_3153,N_1183,N_1014);
nand U3154 (N_3154,N_1123,N_765);
and U3155 (N_3155,N_1060,N_1296);
nand U3156 (N_3156,N_1286,N_789);
and U3157 (N_3157,N_1504,N_1448);
nor U3158 (N_3158,N_908,N_1279);
or U3159 (N_3159,N_252,N_919);
nor U3160 (N_3160,N_1696,N_1112);
and U3161 (N_3161,N_612,N_594);
nand U3162 (N_3162,N_70,N_780);
nand U3163 (N_3163,N_1329,N_438);
or U3164 (N_3164,N_1733,N_160);
nor U3165 (N_3165,N_521,N_254);
and U3166 (N_3166,N_1053,N_1638);
nor U3167 (N_3167,N_1339,N_1443);
and U3168 (N_3168,N_456,N_1066);
nor U3169 (N_3169,N_1402,N_309);
or U3170 (N_3170,N_301,N_1550);
nand U3171 (N_3171,N_266,N_1277);
or U3172 (N_3172,N_1702,N_881);
and U3173 (N_3173,N_452,N_980);
nand U3174 (N_3174,N_250,N_1507);
and U3175 (N_3175,N_907,N_124);
nor U3176 (N_3176,N_135,N_929);
nor U3177 (N_3177,N_400,N_1480);
nand U3178 (N_3178,N_17,N_1948);
and U3179 (N_3179,N_366,N_398);
or U3180 (N_3180,N_105,N_576);
or U3181 (N_3181,N_546,N_59);
or U3182 (N_3182,N_573,N_1047);
xnor U3183 (N_3183,N_838,N_316);
nor U3184 (N_3184,N_1424,N_1433);
nand U3185 (N_3185,N_1283,N_66);
or U3186 (N_3186,N_322,N_374);
nor U3187 (N_3187,N_110,N_1806);
and U3188 (N_3188,N_393,N_110);
or U3189 (N_3189,N_606,N_1796);
nor U3190 (N_3190,N_1061,N_1625);
or U3191 (N_3191,N_1548,N_1141);
or U3192 (N_3192,N_1941,N_361);
nand U3193 (N_3193,N_1906,N_1595);
nor U3194 (N_3194,N_796,N_1077);
nand U3195 (N_3195,N_609,N_1342);
nor U3196 (N_3196,N_996,N_515);
nor U3197 (N_3197,N_955,N_977);
nor U3198 (N_3198,N_95,N_281);
nor U3199 (N_3199,N_99,N_1152);
and U3200 (N_3200,N_1443,N_191);
nand U3201 (N_3201,N_1281,N_237);
or U3202 (N_3202,N_1338,N_352);
and U3203 (N_3203,N_652,N_1174);
or U3204 (N_3204,N_1229,N_1044);
nor U3205 (N_3205,N_1089,N_1726);
nand U3206 (N_3206,N_1750,N_1779);
or U3207 (N_3207,N_749,N_966);
nand U3208 (N_3208,N_1353,N_1280);
or U3209 (N_3209,N_1626,N_1888);
and U3210 (N_3210,N_1472,N_848);
and U3211 (N_3211,N_452,N_323);
and U3212 (N_3212,N_775,N_912);
nand U3213 (N_3213,N_304,N_1395);
or U3214 (N_3214,N_703,N_1444);
and U3215 (N_3215,N_444,N_1679);
nor U3216 (N_3216,N_500,N_1188);
or U3217 (N_3217,N_275,N_1680);
nand U3218 (N_3218,N_1888,N_189);
nand U3219 (N_3219,N_961,N_657);
and U3220 (N_3220,N_1324,N_1747);
and U3221 (N_3221,N_679,N_1396);
or U3222 (N_3222,N_1039,N_896);
nand U3223 (N_3223,N_738,N_1869);
and U3224 (N_3224,N_674,N_1490);
and U3225 (N_3225,N_1647,N_721);
and U3226 (N_3226,N_1050,N_303);
and U3227 (N_3227,N_1501,N_1262);
xor U3228 (N_3228,N_90,N_957);
nand U3229 (N_3229,N_1160,N_1608);
nor U3230 (N_3230,N_1057,N_150);
nor U3231 (N_3231,N_375,N_1831);
nand U3232 (N_3232,N_551,N_1763);
and U3233 (N_3233,N_355,N_82);
nand U3234 (N_3234,N_224,N_1496);
nor U3235 (N_3235,N_618,N_1268);
nor U3236 (N_3236,N_1555,N_1455);
or U3237 (N_3237,N_1870,N_1743);
nand U3238 (N_3238,N_1381,N_450);
nor U3239 (N_3239,N_1006,N_381);
or U3240 (N_3240,N_968,N_1487);
and U3241 (N_3241,N_149,N_1643);
or U3242 (N_3242,N_723,N_639);
nor U3243 (N_3243,N_437,N_379);
or U3244 (N_3244,N_1477,N_247);
xor U3245 (N_3245,N_1531,N_293);
nand U3246 (N_3246,N_1434,N_1771);
nand U3247 (N_3247,N_1369,N_478);
and U3248 (N_3248,N_1972,N_1268);
nor U3249 (N_3249,N_195,N_168);
nor U3250 (N_3250,N_1614,N_1128);
and U3251 (N_3251,N_123,N_1665);
and U3252 (N_3252,N_1497,N_1012);
nor U3253 (N_3253,N_1739,N_115);
nor U3254 (N_3254,N_1959,N_889);
nand U3255 (N_3255,N_1564,N_943);
xor U3256 (N_3256,N_440,N_221);
nand U3257 (N_3257,N_356,N_375);
and U3258 (N_3258,N_1349,N_1955);
nand U3259 (N_3259,N_1424,N_1881);
nor U3260 (N_3260,N_161,N_1250);
nand U3261 (N_3261,N_1572,N_524);
nor U3262 (N_3262,N_636,N_46);
and U3263 (N_3263,N_319,N_363);
or U3264 (N_3264,N_935,N_1860);
or U3265 (N_3265,N_1945,N_1135);
nor U3266 (N_3266,N_985,N_1755);
or U3267 (N_3267,N_1862,N_453);
nand U3268 (N_3268,N_857,N_144);
and U3269 (N_3269,N_910,N_1107);
nor U3270 (N_3270,N_279,N_658);
and U3271 (N_3271,N_1791,N_444);
nor U3272 (N_3272,N_514,N_1896);
or U3273 (N_3273,N_624,N_1432);
nand U3274 (N_3274,N_135,N_1499);
and U3275 (N_3275,N_1779,N_632);
nand U3276 (N_3276,N_400,N_1332);
nand U3277 (N_3277,N_1765,N_1084);
and U3278 (N_3278,N_430,N_282);
nor U3279 (N_3279,N_699,N_695);
nor U3280 (N_3280,N_451,N_644);
nor U3281 (N_3281,N_1083,N_1805);
nor U3282 (N_3282,N_660,N_1546);
nand U3283 (N_3283,N_1523,N_388);
nand U3284 (N_3284,N_1602,N_1298);
or U3285 (N_3285,N_583,N_1144);
nand U3286 (N_3286,N_635,N_1471);
or U3287 (N_3287,N_634,N_640);
or U3288 (N_3288,N_1797,N_1850);
and U3289 (N_3289,N_1049,N_1401);
or U3290 (N_3290,N_723,N_615);
nor U3291 (N_3291,N_1466,N_68);
nand U3292 (N_3292,N_1638,N_66);
or U3293 (N_3293,N_85,N_235);
or U3294 (N_3294,N_1474,N_314);
or U3295 (N_3295,N_1930,N_688);
and U3296 (N_3296,N_778,N_236);
and U3297 (N_3297,N_62,N_1748);
nand U3298 (N_3298,N_371,N_1047);
nand U3299 (N_3299,N_775,N_881);
or U3300 (N_3300,N_1154,N_1086);
nand U3301 (N_3301,N_1427,N_462);
and U3302 (N_3302,N_1316,N_564);
nand U3303 (N_3303,N_706,N_1647);
nand U3304 (N_3304,N_1795,N_848);
nand U3305 (N_3305,N_813,N_236);
nand U3306 (N_3306,N_484,N_1187);
nor U3307 (N_3307,N_232,N_1276);
nor U3308 (N_3308,N_934,N_1330);
nor U3309 (N_3309,N_1622,N_348);
nor U3310 (N_3310,N_287,N_283);
and U3311 (N_3311,N_1223,N_1816);
nor U3312 (N_3312,N_735,N_461);
or U3313 (N_3313,N_155,N_726);
xnor U3314 (N_3314,N_70,N_893);
and U3315 (N_3315,N_1686,N_1148);
and U3316 (N_3316,N_1800,N_301);
and U3317 (N_3317,N_1904,N_864);
or U3318 (N_3318,N_1283,N_24);
or U3319 (N_3319,N_1538,N_1533);
or U3320 (N_3320,N_563,N_1536);
or U3321 (N_3321,N_770,N_1599);
and U3322 (N_3322,N_50,N_409);
and U3323 (N_3323,N_14,N_1508);
nand U3324 (N_3324,N_455,N_1313);
or U3325 (N_3325,N_750,N_1206);
or U3326 (N_3326,N_1490,N_209);
or U3327 (N_3327,N_1424,N_1698);
nor U3328 (N_3328,N_1158,N_1763);
nand U3329 (N_3329,N_905,N_925);
nand U3330 (N_3330,N_552,N_307);
nand U3331 (N_3331,N_1375,N_308);
xor U3332 (N_3332,N_1251,N_26);
and U3333 (N_3333,N_406,N_1478);
nor U3334 (N_3334,N_190,N_425);
and U3335 (N_3335,N_1894,N_229);
and U3336 (N_3336,N_1392,N_335);
or U3337 (N_3337,N_1716,N_1695);
nand U3338 (N_3338,N_463,N_1026);
nor U3339 (N_3339,N_1185,N_1865);
and U3340 (N_3340,N_266,N_1664);
and U3341 (N_3341,N_609,N_502);
xor U3342 (N_3342,N_1883,N_1624);
xnor U3343 (N_3343,N_313,N_1432);
or U3344 (N_3344,N_1169,N_936);
nor U3345 (N_3345,N_935,N_1869);
or U3346 (N_3346,N_429,N_1184);
or U3347 (N_3347,N_1042,N_385);
nor U3348 (N_3348,N_1560,N_62);
or U3349 (N_3349,N_619,N_411);
or U3350 (N_3350,N_1367,N_995);
nor U3351 (N_3351,N_1855,N_522);
nand U3352 (N_3352,N_295,N_721);
and U3353 (N_3353,N_383,N_35);
or U3354 (N_3354,N_1889,N_1921);
and U3355 (N_3355,N_559,N_252);
or U3356 (N_3356,N_1462,N_1185);
and U3357 (N_3357,N_1012,N_899);
nor U3358 (N_3358,N_851,N_998);
and U3359 (N_3359,N_104,N_143);
nand U3360 (N_3360,N_1403,N_1738);
nand U3361 (N_3361,N_1870,N_195);
nand U3362 (N_3362,N_1753,N_69);
or U3363 (N_3363,N_487,N_1569);
or U3364 (N_3364,N_1626,N_1450);
nor U3365 (N_3365,N_817,N_1290);
nor U3366 (N_3366,N_1888,N_1902);
nor U3367 (N_3367,N_1897,N_1969);
nor U3368 (N_3368,N_1048,N_1200);
or U3369 (N_3369,N_413,N_1507);
and U3370 (N_3370,N_515,N_109);
nor U3371 (N_3371,N_878,N_236);
or U3372 (N_3372,N_1991,N_1116);
and U3373 (N_3373,N_1461,N_1923);
nand U3374 (N_3374,N_715,N_1353);
nor U3375 (N_3375,N_1053,N_1015);
or U3376 (N_3376,N_1739,N_1344);
nand U3377 (N_3377,N_1079,N_41);
or U3378 (N_3378,N_1060,N_194);
nand U3379 (N_3379,N_219,N_1928);
nor U3380 (N_3380,N_1312,N_356);
nand U3381 (N_3381,N_642,N_708);
or U3382 (N_3382,N_1462,N_938);
nand U3383 (N_3383,N_749,N_1231);
and U3384 (N_3384,N_787,N_173);
or U3385 (N_3385,N_1945,N_1809);
or U3386 (N_3386,N_1061,N_1270);
nand U3387 (N_3387,N_887,N_41);
nor U3388 (N_3388,N_997,N_608);
nand U3389 (N_3389,N_823,N_1963);
or U3390 (N_3390,N_1899,N_811);
and U3391 (N_3391,N_1649,N_489);
nand U3392 (N_3392,N_374,N_330);
nor U3393 (N_3393,N_1423,N_1315);
or U3394 (N_3394,N_1642,N_587);
nand U3395 (N_3395,N_1841,N_1890);
and U3396 (N_3396,N_1021,N_351);
or U3397 (N_3397,N_1655,N_155);
and U3398 (N_3398,N_970,N_1245);
and U3399 (N_3399,N_1096,N_1237);
or U3400 (N_3400,N_1969,N_948);
nor U3401 (N_3401,N_452,N_1879);
nand U3402 (N_3402,N_1855,N_1377);
nand U3403 (N_3403,N_1449,N_1993);
nor U3404 (N_3404,N_1356,N_1706);
nor U3405 (N_3405,N_1054,N_1102);
and U3406 (N_3406,N_290,N_817);
and U3407 (N_3407,N_77,N_378);
and U3408 (N_3408,N_1298,N_1965);
nor U3409 (N_3409,N_1822,N_324);
or U3410 (N_3410,N_1937,N_564);
and U3411 (N_3411,N_1276,N_4);
and U3412 (N_3412,N_1324,N_1521);
xor U3413 (N_3413,N_567,N_1444);
nand U3414 (N_3414,N_581,N_369);
xnor U3415 (N_3415,N_1914,N_943);
and U3416 (N_3416,N_452,N_206);
and U3417 (N_3417,N_840,N_45);
and U3418 (N_3418,N_679,N_411);
or U3419 (N_3419,N_1108,N_68);
and U3420 (N_3420,N_16,N_875);
and U3421 (N_3421,N_575,N_917);
nand U3422 (N_3422,N_923,N_755);
nand U3423 (N_3423,N_1655,N_1289);
nand U3424 (N_3424,N_334,N_1126);
xnor U3425 (N_3425,N_703,N_918);
nor U3426 (N_3426,N_562,N_238);
nand U3427 (N_3427,N_1771,N_1394);
nor U3428 (N_3428,N_667,N_1074);
nor U3429 (N_3429,N_544,N_864);
or U3430 (N_3430,N_544,N_733);
nor U3431 (N_3431,N_1843,N_826);
nor U3432 (N_3432,N_713,N_625);
or U3433 (N_3433,N_1787,N_297);
nand U3434 (N_3434,N_1594,N_1283);
nand U3435 (N_3435,N_1314,N_98);
and U3436 (N_3436,N_942,N_440);
and U3437 (N_3437,N_1395,N_1937);
nor U3438 (N_3438,N_71,N_611);
nand U3439 (N_3439,N_1745,N_1227);
and U3440 (N_3440,N_1582,N_454);
and U3441 (N_3441,N_566,N_14);
or U3442 (N_3442,N_444,N_1035);
and U3443 (N_3443,N_137,N_739);
nand U3444 (N_3444,N_701,N_1181);
and U3445 (N_3445,N_1338,N_1509);
nor U3446 (N_3446,N_26,N_1855);
nand U3447 (N_3447,N_272,N_127);
nor U3448 (N_3448,N_186,N_264);
and U3449 (N_3449,N_1170,N_727);
or U3450 (N_3450,N_1485,N_547);
or U3451 (N_3451,N_1728,N_71);
or U3452 (N_3452,N_1799,N_528);
and U3453 (N_3453,N_1953,N_1582);
or U3454 (N_3454,N_838,N_1921);
or U3455 (N_3455,N_495,N_383);
or U3456 (N_3456,N_833,N_726);
or U3457 (N_3457,N_1920,N_1852);
or U3458 (N_3458,N_1233,N_1445);
or U3459 (N_3459,N_1388,N_87);
or U3460 (N_3460,N_704,N_973);
or U3461 (N_3461,N_263,N_1253);
or U3462 (N_3462,N_1862,N_1029);
nor U3463 (N_3463,N_543,N_47);
and U3464 (N_3464,N_1508,N_672);
or U3465 (N_3465,N_279,N_666);
nand U3466 (N_3466,N_1015,N_1513);
and U3467 (N_3467,N_1562,N_1746);
or U3468 (N_3468,N_1997,N_1245);
and U3469 (N_3469,N_281,N_1045);
nor U3470 (N_3470,N_310,N_432);
or U3471 (N_3471,N_1049,N_1245);
or U3472 (N_3472,N_1338,N_1228);
and U3473 (N_3473,N_290,N_1246);
and U3474 (N_3474,N_1149,N_1535);
or U3475 (N_3475,N_516,N_74);
nand U3476 (N_3476,N_1648,N_978);
nand U3477 (N_3477,N_958,N_131);
and U3478 (N_3478,N_1791,N_971);
nand U3479 (N_3479,N_1625,N_263);
or U3480 (N_3480,N_204,N_525);
nand U3481 (N_3481,N_1926,N_1555);
or U3482 (N_3482,N_1827,N_1661);
nor U3483 (N_3483,N_916,N_1196);
nor U3484 (N_3484,N_1046,N_1512);
and U3485 (N_3485,N_1436,N_659);
and U3486 (N_3486,N_1902,N_987);
and U3487 (N_3487,N_1682,N_152);
and U3488 (N_3488,N_426,N_1635);
or U3489 (N_3489,N_568,N_875);
and U3490 (N_3490,N_1339,N_1584);
or U3491 (N_3491,N_889,N_363);
or U3492 (N_3492,N_394,N_1607);
or U3493 (N_3493,N_45,N_1437);
xnor U3494 (N_3494,N_52,N_1346);
nor U3495 (N_3495,N_1311,N_1249);
nand U3496 (N_3496,N_1473,N_1233);
or U3497 (N_3497,N_420,N_1715);
and U3498 (N_3498,N_1575,N_1379);
and U3499 (N_3499,N_229,N_1308);
nor U3500 (N_3500,N_1577,N_1973);
and U3501 (N_3501,N_1781,N_1286);
xor U3502 (N_3502,N_958,N_1426);
nor U3503 (N_3503,N_1110,N_1816);
nor U3504 (N_3504,N_355,N_170);
or U3505 (N_3505,N_969,N_549);
and U3506 (N_3506,N_536,N_1276);
nor U3507 (N_3507,N_768,N_1932);
and U3508 (N_3508,N_981,N_1541);
and U3509 (N_3509,N_1398,N_1671);
nor U3510 (N_3510,N_1756,N_607);
nand U3511 (N_3511,N_248,N_42);
or U3512 (N_3512,N_570,N_1911);
nand U3513 (N_3513,N_999,N_859);
and U3514 (N_3514,N_1916,N_1343);
nand U3515 (N_3515,N_924,N_74);
nand U3516 (N_3516,N_1338,N_858);
xnor U3517 (N_3517,N_1480,N_1094);
nor U3518 (N_3518,N_1452,N_584);
nand U3519 (N_3519,N_188,N_1341);
and U3520 (N_3520,N_763,N_1308);
and U3521 (N_3521,N_1301,N_1586);
or U3522 (N_3522,N_727,N_1292);
nor U3523 (N_3523,N_136,N_1521);
and U3524 (N_3524,N_1097,N_1010);
and U3525 (N_3525,N_789,N_1288);
nand U3526 (N_3526,N_899,N_136);
or U3527 (N_3527,N_576,N_399);
or U3528 (N_3528,N_1485,N_893);
and U3529 (N_3529,N_887,N_1675);
or U3530 (N_3530,N_492,N_1228);
or U3531 (N_3531,N_1090,N_1936);
nand U3532 (N_3532,N_365,N_885);
or U3533 (N_3533,N_149,N_1733);
nor U3534 (N_3534,N_321,N_1097);
or U3535 (N_3535,N_1356,N_1159);
nand U3536 (N_3536,N_749,N_1466);
nor U3537 (N_3537,N_1766,N_1881);
nor U3538 (N_3538,N_1977,N_1267);
and U3539 (N_3539,N_1283,N_1817);
nor U3540 (N_3540,N_277,N_1986);
nor U3541 (N_3541,N_1635,N_1576);
nor U3542 (N_3542,N_766,N_889);
nand U3543 (N_3543,N_1658,N_749);
and U3544 (N_3544,N_1014,N_1908);
nor U3545 (N_3545,N_1658,N_1995);
and U3546 (N_3546,N_1983,N_263);
nand U3547 (N_3547,N_1478,N_1497);
nand U3548 (N_3548,N_1425,N_903);
or U3549 (N_3549,N_853,N_1602);
and U3550 (N_3550,N_1868,N_1146);
nand U3551 (N_3551,N_36,N_1501);
or U3552 (N_3552,N_1349,N_414);
and U3553 (N_3553,N_496,N_1853);
nor U3554 (N_3554,N_1159,N_1508);
or U3555 (N_3555,N_85,N_635);
and U3556 (N_3556,N_1021,N_1114);
or U3557 (N_3557,N_1802,N_1960);
and U3558 (N_3558,N_1209,N_1221);
or U3559 (N_3559,N_148,N_920);
nor U3560 (N_3560,N_547,N_1868);
and U3561 (N_3561,N_362,N_1959);
and U3562 (N_3562,N_1476,N_499);
or U3563 (N_3563,N_1351,N_1989);
nor U3564 (N_3564,N_393,N_35);
nand U3565 (N_3565,N_472,N_1387);
nor U3566 (N_3566,N_1641,N_1413);
nor U3567 (N_3567,N_943,N_288);
and U3568 (N_3568,N_672,N_1639);
nor U3569 (N_3569,N_1233,N_777);
or U3570 (N_3570,N_703,N_761);
xor U3571 (N_3571,N_600,N_188);
or U3572 (N_3572,N_781,N_1428);
xnor U3573 (N_3573,N_1837,N_1506);
nor U3574 (N_3574,N_1103,N_912);
nand U3575 (N_3575,N_1756,N_1607);
and U3576 (N_3576,N_1204,N_275);
and U3577 (N_3577,N_1444,N_1344);
and U3578 (N_3578,N_1817,N_1289);
or U3579 (N_3579,N_71,N_819);
nor U3580 (N_3580,N_1990,N_479);
nand U3581 (N_3581,N_996,N_960);
nand U3582 (N_3582,N_108,N_174);
nor U3583 (N_3583,N_1530,N_1503);
and U3584 (N_3584,N_1398,N_1681);
nand U3585 (N_3585,N_1942,N_981);
or U3586 (N_3586,N_744,N_1665);
nand U3587 (N_3587,N_45,N_442);
nand U3588 (N_3588,N_505,N_1161);
nor U3589 (N_3589,N_1320,N_577);
nor U3590 (N_3590,N_865,N_270);
and U3591 (N_3591,N_1209,N_1019);
nand U3592 (N_3592,N_999,N_1317);
and U3593 (N_3593,N_634,N_627);
nand U3594 (N_3594,N_103,N_825);
nand U3595 (N_3595,N_165,N_1044);
nor U3596 (N_3596,N_1576,N_687);
or U3597 (N_3597,N_1643,N_1020);
nor U3598 (N_3598,N_1060,N_87);
and U3599 (N_3599,N_76,N_401);
nand U3600 (N_3600,N_421,N_1424);
and U3601 (N_3601,N_1018,N_729);
and U3602 (N_3602,N_138,N_498);
or U3603 (N_3603,N_957,N_1767);
or U3604 (N_3604,N_1191,N_1112);
or U3605 (N_3605,N_1542,N_1422);
nor U3606 (N_3606,N_536,N_65);
nand U3607 (N_3607,N_1716,N_1284);
nand U3608 (N_3608,N_56,N_1913);
or U3609 (N_3609,N_1177,N_1042);
and U3610 (N_3610,N_1274,N_1315);
nor U3611 (N_3611,N_735,N_1008);
nand U3612 (N_3612,N_448,N_1951);
nand U3613 (N_3613,N_406,N_622);
nand U3614 (N_3614,N_740,N_5);
nor U3615 (N_3615,N_1299,N_1976);
nor U3616 (N_3616,N_1563,N_360);
and U3617 (N_3617,N_1767,N_1080);
and U3618 (N_3618,N_1322,N_49);
or U3619 (N_3619,N_1899,N_1260);
xor U3620 (N_3620,N_1243,N_953);
or U3621 (N_3621,N_277,N_1154);
or U3622 (N_3622,N_1926,N_403);
nand U3623 (N_3623,N_1219,N_1367);
and U3624 (N_3624,N_1092,N_354);
and U3625 (N_3625,N_1993,N_1592);
nor U3626 (N_3626,N_1506,N_1849);
or U3627 (N_3627,N_792,N_1107);
and U3628 (N_3628,N_1421,N_1119);
nand U3629 (N_3629,N_836,N_241);
xnor U3630 (N_3630,N_1933,N_813);
or U3631 (N_3631,N_1487,N_194);
nand U3632 (N_3632,N_1937,N_719);
nor U3633 (N_3633,N_150,N_972);
nand U3634 (N_3634,N_133,N_335);
nor U3635 (N_3635,N_1637,N_488);
and U3636 (N_3636,N_40,N_746);
nand U3637 (N_3637,N_85,N_813);
or U3638 (N_3638,N_1691,N_210);
nor U3639 (N_3639,N_328,N_1526);
and U3640 (N_3640,N_318,N_1267);
nand U3641 (N_3641,N_598,N_1107);
nand U3642 (N_3642,N_680,N_1347);
and U3643 (N_3643,N_1445,N_340);
or U3644 (N_3644,N_1883,N_1687);
or U3645 (N_3645,N_813,N_865);
or U3646 (N_3646,N_1604,N_186);
nor U3647 (N_3647,N_1006,N_1122);
nor U3648 (N_3648,N_676,N_1907);
nand U3649 (N_3649,N_623,N_1405);
nand U3650 (N_3650,N_1734,N_1097);
or U3651 (N_3651,N_1512,N_1959);
or U3652 (N_3652,N_227,N_367);
nand U3653 (N_3653,N_1485,N_952);
and U3654 (N_3654,N_414,N_1463);
nand U3655 (N_3655,N_40,N_1479);
nor U3656 (N_3656,N_518,N_1515);
and U3657 (N_3657,N_1433,N_426);
or U3658 (N_3658,N_634,N_1989);
nand U3659 (N_3659,N_550,N_1334);
nand U3660 (N_3660,N_1940,N_442);
nand U3661 (N_3661,N_1159,N_1349);
nor U3662 (N_3662,N_1918,N_1185);
nor U3663 (N_3663,N_757,N_1069);
and U3664 (N_3664,N_1655,N_766);
and U3665 (N_3665,N_1848,N_1322);
nand U3666 (N_3666,N_1988,N_1932);
nor U3667 (N_3667,N_1333,N_1778);
nand U3668 (N_3668,N_1055,N_1269);
nor U3669 (N_3669,N_1506,N_416);
or U3670 (N_3670,N_1943,N_39);
nor U3671 (N_3671,N_436,N_1724);
or U3672 (N_3672,N_1077,N_1792);
nand U3673 (N_3673,N_1980,N_567);
nand U3674 (N_3674,N_1089,N_1238);
or U3675 (N_3675,N_1755,N_1038);
nor U3676 (N_3676,N_767,N_68);
or U3677 (N_3677,N_1095,N_1334);
nor U3678 (N_3678,N_1865,N_596);
nor U3679 (N_3679,N_102,N_1076);
or U3680 (N_3680,N_1459,N_1969);
nor U3681 (N_3681,N_1832,N_971);
or U3682 (N_3682,N_509,N_1241);
nor U3683 (N_3683,N_182,N_1966);
or U3684 (N_3684,N_1602,N_299);
or U3685 (N_3685,N_1467,N_1509);
or U3686 (N_3686,N_616,N_673);
nor U3687 (N_3687,N_1297,N_158);
nor U3688 (N_3688,N_1472,N_1735);
or U3689 (N_3689,N_771,N_359);
nand U3690 (N_3690,N_24,N_1498);
nor U3691 (N_3691,N_833,N_1150);
nor U3692 (N_3692,N_507,N_905);
and U3693 (N_3693,N_1420,N_421);
nand U3694 (N_3694,N_1861,N_1034);
and U3695 (N_3695,N_1999,N_969);
and U3696 (N_3696,N_405,N_452);
nor U3697 (N_3697,N_1441,N_666);
or U3698 (N_3698,N_515,N_1529);
and U3699 (N_3699,N_963,N_1956);
nand U3700 (N_3700,N_1595,N_1578);
nand U3701 (N_3701,N_1072,N_1520);
or U3702 (N_3702,N_1697,N_1238);
nor U3703 (N_3703,N_1219,N_799);
nand U3704 (N_3704,N_633,N_121);
nand U3705 (N_3705,N_1726,N_1816);
or U3706 (N_3706,N_569,N_1363);
nor U3707 (N_3707,N_524,N_1931);
nand U3708 (N_3708,N_609,N_770);
nand U3709 (N_3709,N_1908,N_1665);
or U3710 (N_3710,N_1987,N_1951);
and U3711 (N_3711,N_214,N_721);
nor U3712 (N_3712,N_1349,N_1747);
nor U3713 (N_3713,N_1813,N_775);
nor U3714 (N_3714,N_1250,N_1299);
xor U3715 (N_3715,N_1677,N_1889);
nand U3716 (N_3716,N_358,N_562);
or U3717 (N_3717,N_1177,N_451);
and U3718 (N_3718,N_336,N_1276);
nand U3719 (N_3719,N_4,N_698);
nor U3720 (N_3720,N_1627,N_436);
xor U3721 (N_3721,N_1689,N_1398);
and U3722 (N_3722,N_685,N_896);
nor U3723 (N_3723,N_1513,N_965);
or U3724 (N_3724,N_819,N_731);
or U3725 (N_3725,N_1031,N_963);
or U3726 (N_3726,N_1408,N_311);
or U3727 (N_3727,N_1669,N_1921);
nand U3728 (N_3728,N_1160,N_1703);
nor U3729 (N_3729,N_1022,N_1541);
and U3730 (N_3730,N_1167,N_1455);
nand U3731 (N_3731,N_938,N_457);
or U3732 (N_3732,N_1327,N_1348);
or U3733 (N_3733,N_1218,N_499);
and U3734 (N_3734,N_653,N_156);
nor U3735 (N_3735,N_315,N_516);
or U3736 (N_3736,N_388,N_1866);
and U3737 (N_3737,N_1452,N_1261);
or U3738 (N_3738,N_1008,N_1580);
nand U3739 (N_3739,N_1554,N_1958);
and U3740 (N_3740,N_1103,N_429);
or U3741 (N_3741,N_198,N_399);
nand U3742 (N_3742,N_1300,N_1680);
or U3743 (N_3743,N_1230,N_52);
and U3744 (N_3744,N_790,N_1386);
or U3745 (N_3745,N_218,N_1410);
and U3746 (N_3746,N_999,N_1470);
or U3747 (N_3747,N_546,N_1436);
and U3748 (N_3748,N_705,N_905);
nor U3749 (N_3749,N_1267,N_1372);
nand U3750 (N_3750,N_142,N_779);
or U3751 (N_3751,N_1293,N_1857);
or U3752 (N_3752,N_1874,N_1933);
and U3753 (N_3753,N_346,N_1596);
nand U3754 (N_3754,N_1284,N_655);
nand U3755 (N_3755,N_983,N_773);
or U3756 (N_3756,N_640,N_1002);
and U3757 (N_3757,N_85,N_1293);
and U3758 (N_3758,N_1622,N_1612);
nand U3759 (N_3759,N_1194,N_959);
nand U3760 (N_3760,N_586,N_1207);
nor U3761 (N_3761,N_1868,N_947);
or U3762 (N_3762,N_1061,N_1344);
or U3763 (N_3763,N_78,N_194);
nand U3764 (N_3764,N_375,N_1913);
nor U3765 (N_3765,N_1042,N_275);
or U3766 (N_3766,N_222,N_323);
nand U3767 (N_3767,N_1271,N_1509);
or U3768 (N_3768,N_86,N_781);
or U3769 (N_3769,N_19,N_1154);
nand U3770 (N_3770,N_306,N_506);
or U3771 (N_3771,N_1180,N_797);
or U3772 (N_3772,N_553,N_1207);
and U3773 (N_3773,N_16,N_1004);
and U3774 (N_3774,N_899,N_80);
nor U3775 (N_3775,N_1191,N_388);
nand U3776 (N_3776,N_411,N_461);
nand U3777 (N_3777,N_1608,N_13);
nand U3778 (N_3778,N_88,N_837);
or U3779 (N_3779,N_674,N_992);
nand U3780 (N_3780,N_235,N_1678);
nor U3781 (N_3781,N_1391,N_1685);
or U3782 (N_3782,N_1082,N_1734);
nor U3783 (N_3783,N_1492,N_338);
or U3784 (N_3784,N_611,N_1448);
nor U3785 (N_3785,N_1839,N_783);
nor U3786 (N_3786,N_1184,N_1204);
or U3787 (N_3787,N_1529,N_1368);
nor U3788 (N_3788,N_462,N_1431);
or U3789 (N_3789,N_1240,N_306);
and U3790 (N_3790,N_1071,N_1583);
and U3791 (N_3791,N_839,N_1058);
and U3792 (N_3792,N_1601,N_1492);
nor U3793 (N_3793,N_1664,N_1342);
and U3794 (N_3794,N_508,N_1817);
nor U3795 (N_3795,N_578,N_105);
nor U3796 (N_3796,N_90,N_428);
nor U3797 (N_3797,N_285,N_1537);
xnor U3798 (N_3798,N_995,N_1000);
and U3799 (N_3799,N_911,N_933);
nand U3800 (N_3800,N_1294,N_62);
nor U3801 (N_3801,N_768,N_1073);
nor U3802 (N_3802,N_148,N_448);
nand U3803 (N_3803,N_1977,N_408);
nand U3804 (N_3804,N_1555,N_1256);
or U3805 (N_3805,N_1388,N_320);
or U3806 (N_3806,N_584,N_1897);
nor U3807 (N_3807,N_660,N_1540);
and U3808 (N_3808,N_1901,N_1426);
and U3809 (N_3809,N_760,N_1967);
or U3810 (N_3810,N_1214,N_1602);
nor U3811 (N_3811,N_1800,N_1359);
xnor U3812 (N_3812,N_1020,N_608);
nand U3813 (N_3813,N_438,N_1116);
nor U3814 (N_3814,N_1089,N_1302);
and U3815 (N_3815,N_211,N_126);
nand U3816 (N_3816,N_1878,N_1561);
nor U3817 (N_3817,N_161,N_1111);
nor U3818 (N_3818,N_1076,N_676);
xnor U3819 (N_3819,N_671,N_1798);
and U3820 (N_3820,N_107,N_1852);
nor U3821 (N_3821,N_319,N_1234);
and U3822 (N_3822,N_975,N_698);
or U3823 (N_3823,N_1015,N_1820);
nor U3824 (N_3824,N_143,N_648);
nor U3825 (N_3825,N_988,N_1785);
nor U3826 (N_3826,N_636,N_1693);
nand U3827 (N_3827,N_1878,N_1028);
nor U3828 (N_3828,N_44,N_1168);
and U3829 (N_3829,N_51,N_1204);
or U3830 (N_3830,N_13,N_1088);
nor U3831 (N_3831,N_528,N_651);
nand U3832 (N_3832,N_1688,N_540);
xnor U3833 (N_3833,N_654,N_1135);
or U3834 (N_3834,N_694,N_767);
nor U3835 (N_3835,N_79,N_1465);
nand U3836 (N_3836,N_1372,N_552);
nor U3837 (N_3837,N_1182,N_1052);
nor U3838 (N_3838,N_1741,N_204);
nor U3839 (N_3839,N_1811,N_1974);
and U3840 (N_3840,N_1253,N_1061);
nor U3841 (N_3841,N_553,N_563);
nor U3842 (N_3842,N_104,N_903);
and U3843 (N_3843,N_1981,N_1471);
nand U3844 (N_3844,N_1880,N_1551);
or U3845 (N_3845,N_115,N_1437);
nand U3846 (N_3846,N_1492,N_1712);
and U3847 (N_3847,N_1025,N_1106);
or U3848 (N_3848,N_943,N_1843);
nor U3849 (N_3849,N_1897,N_976);
or U3850 (N_3850,N_944,N_932);
or U3851 (N_3851,N_1462,N_1874);
and U3852 (N_3852,N_431,N_36);
nand U3853 (N_3853,N_1649,N_1690);
or U3854 (N_3854,N_879,N_378);
nand U3855 (N_3855,N_1438,N_234);
and U3856 (N_3856,N_1310,N_1786);
nand U3857 (N_3857,N_1188,N_1063);
xnor U3858 (N_3858,N_163,N_1347);
or U3859 (N_3859,N_1690,N_1468);
nand U3860 (N_3860,N_1758,N_1192);
and U3861 (N_3861,N_1117,N_1501);
nor U3862 (N_3862,N_1793,N_445);
xor U3863 (N_3863,N_1180,N_1457);
and U3864 (N_3864,N_1050,N_1161);
and U3865 (N_3865,N_806,N_178);
or U3866 (N_3866,N_329,N_883);
nand U3867 (N_3867,N_1795,N_1629);
and U3868 (N_3868,N_361,N_1532);
nor U3869 (N_3869,N_1044,N_1280);
and U3870 (N_3870,N_107,N_1616);
or U3871 (N_3871,N_1124,N_1673);
xnor U3872 (N_3872,N_1371,N_1410);
and U3873 (N_3873,N_120,N_1856);
or U3874 (N_3874,N_418,N_1169);
or U3875 (N_3875,N_1969,N_507);
or U3876 (N_3876,N_432,N_954);
and U3877 (N_3877,N_919,N_1237);
or U3878 (N_3878,N_798,N_1218);
nand U3879 (N_3879,N_1807,N_500);
nand U3880 (N_3880,N_1479,N_1611);
and U3881 (N_3881,N_1929,N_1805);
or U3882 (N_3882,N_55,N_488);
nor U3883 (N_3883,N_1669,N_109);
or U3884 (N_3884,N_1648,N_1147);
nand U3885 (N_3885,N_1806,N_1247);
nand U3886 (N_3886,N_1050,N_1252);
or U3887 (N_3887,N_40,N_1622);
nor U3888 (N_3888,N_679,N_1042);
or U3889 (N_3889,N_1112,N_1600);
xor U3890 (N_3890,N_1585,N_126);
xor U3891 (N_3891,N_149,N_789);
nand U3892 (N_3892,N_706,N_805);
nand U3893 (N_3893,N_1928,N_1417);
nor U3894 (N_3894,N_1535,N_1709);
and U3895 (N_3895,N_140,N_1007);
and U3896 (N_3896,N_1678,N_165);
or U3897 (N_3897,N_940,N_843);
or U3898 (N_3898,N_1296,N_1671);
nor U3899 (N_3899,N_814,N_881);
nand U3900 (N_3900,N_1163,N_1568);
or U3901 (N_3901,N_1374,N_936);
nand U3902 (N_3902,N_593,N_563);
and U3903 (N_3903,N_1058,N_940);
nand U3904 (N_3904,N_1296,N_1046);
xnor U3905 (N_3905,N_75,N_1630);
or U3906 (N_3906,N_775,N_181);
and U3907 (N_3907,N_578,N_736);
nand U3908 (N_3908,N_1630,N_29);
or U3909 (N_3909,N_926,N_1879);
and U3910 (N_3910,N_1112,N_1548);
and U3911 (N_3911,N_622,N_299);
nand U3912 (N_3912,N_560,N_1474);
or U3913 (N_3913,N_1246,N_1206);
nor U3914 (N_3914,N_541,N_1911);
nand U3915 (N_3915,N_1562,N_1524);
and U3916 (N_3916,N_1105,N_1455);
or U3917 (N_3917,N_615,N_388);
nand U3918 (N_3918,N_1594,N_964);
and U3919 (N_3919,N_1645,N_532);
and U3920 (N_3920,N_1887,N_999);
nor U3921 (N_3921,N_801,N_1729);
and U3922 (N_3922,N_1395,N_1980);
nand U3923 (N_3923,N_1953,N_162);
nor U3924 (N_3924,N_1032,N_634);
nor U3925 (N_3925,N_95,N_1024);
nor U3926 (N_3926,N_1335,N_166);
nor U3927 (N_3927,N_369,N_428);
and U3928 (N_3928,N_1510,N_1165);
nand U3929 (N_3929,N_594,N_243);
nor U3930 (N_3930,N_1887,N_165);
and U3931 (N_3931,N_704,N_1454);
nand U3932 (N_3932,N_1985,N_165);
and U3933 (N_3933,N_1121,N_1882);
or U3934 (N_3934,N_229,N_899);
nor U3935 (N_3935,N_1520,N_1260);
and U3936 (N_3936,N_1410,N_966);
nor U3937 (N_3937,N_471,N_1165);
or U3938 (N_3938,N_1535,N_242);
and U3939 (N_3939,N_309,N_923);
and U3940 (N_3940,N_1057,N_920);
nand U3941 (N_3941,N_863,N_1483);
nand U3942 (N_3942,N_1060,N_388);
and U3943 (N_3943,N_265,N_69);
nand U3944 (N_3944,N_1666,N_598);
nor U3945 (N_3945,N_975,N_816);
or U3946 (N_3946,N_380,N_692);
or U3947 (N_3947,N_258,N_362);
or U3948 (N_3948,N_986,N_1738);
or U3949 (N_3949,N_1147,N_1612);
and U3950 (N_3950,N_1433,N_1136);
nor U3951 (N_3951,N_1392,N_996);
nand U3952 (N_3952,N_420,N_980);
nor U3953 (N_3953,N_765,N_1169);
nor U3954 (N_3954,N_1707,N_672);
nor U3955 (N_3955,N_812,N_1030);
nand U3956 (N_3956,N_1733,N_302);
or U3957 (N_3957,N_999,N_1618);
nand U3958 (N_3958,N_1859,N_932);
nor U3959 (N_3959,N_1595,N_68);
and U3960 (N_3960,N_1840,N_681);
and U3961 (N_3961,N_322,N_1783);
nor U3962 (N_3962,N_403,N_1006);
nand U3963 (N_3963,N_1885,N_1096);
nand U3964 (N_3964,N_272,N_1342);
nand U3965 (N_3965,N_704,N_1052);
nor U3966 (N_3966,N_1981,N_248);
nand U3967 (N_3967,N_1497,N_686);
nand U3968 (N_3968,N_1522,N_1665);
xor U3969 (N_3969,N_485,N_1418);
nor U3970 (N_3970,N_921,N_376);
nand U3971 (N_3971,N_326,N_1287);
xor U3972 (N_3972,N_11,N_438);
nor U3973 (N_3973,N_852,N_1661);
nor U3974 (N_3974,N_1059,N_357);
nor U3975 (N_3975,N_833,N_979);
nand U3976 (N_3976,N_466,N_463);
or U3977 (N_3977,N_572,N_1170);
and U3978 (N_3978,N_967,N_530);
nand U3979 (N_3979,N_668,N_1609);
nor U3980 (N_3980,N_547,N_1744);
nor U3981 (N_3981,N_1947,N_1047);
nand U3982 (N_3982,N_641,N_561);
or U3983 (N_3983,N_216,N_1967);
and U3984 (N_3984,N_412,N_1962);
or U3985 (N_3985,N_670,N_1691);
nor U3986 (N_3986,N_1969,N_1362);
nor U3987 (N_3987,N_1826,N_505);
or U3988 (N_3988,N_567,N_39);
nor U3989 (N_3989,N_1361,N_984);
nor U3990 (N_3990,N_743,N_612);
and U3991 (N_3991,N_1502,N_989);
or U3992 (N_3992,N_1618,N_1438);
nand U3993 (N_3993,N_177,N_202);
and U3994 (N_3994,N_1488,N_373);
and U3995 (N_3995,N_1841,N_1833);
nor U3996 (N_3996,N_992,N_791);
nand U3997 (N_3997,N_1033,N_1078);
and U3998 (N_3998,N_1645,N_1962);
nand U3999 (N_3999,N_1978,N_1384);
or U4000 (N_4000,N_3079,N_3908);
and U4001 (N_4001,N_2618,N_2073);
and U4002 (N_4002,N_3081,N_3287);
nand U4003 (N_4003,N_2343,N_2958);
or U4004 (N_4004,N_2535,N_2558);
and U4005 (N_4005,N_3049,N_3887);
or U4006 (N_4006,N_2701,N_2715);
or U4007 (N_4007,N_2931,N_3331);
nand U4008 (N_4008,N_2988,N_2703);
nor U4009 (N_4009,N_2069,N_3947);
nor U4010 (N_4010,N_3562,N_3102);
and U4011 (N_4011,N_2990,N_3439);
or U4012 (N_4012,N_2731,N_2268);
nand U4013 (N_4013,N_3504,N_3796);
or U4014 (N_4014,N_2012,N_2240);
nor U4015 (N_4015,N_3836,N_2885);
and U4016 (N_4016,N_3561,N_2400);
nand U4017 (N_4017,N_2808,N_3142);
or U4018 (N_4018,N_3986,N_3804);
nor U4019 (N_4019,N_3031,N_3851);
nand U4020 (N_4020,N_2824,N_2258);
nand U4021 (N_4021,N_3445,N_3355);
and U4022 (N_4022,N_3095,N_3353);
nand U4023 (N_4023,N_2660,N_3199);
nand U4024 (N_4024,N_3954,N_2003);
nor U4025 (N_4025,N_3437,N_3792);
and U4026 (N_4026,N_3741,N_2373);
or U4027 (N_4027,N_3289,N_3164);
nand U4028 (N_4028,N_3111,N_3458);
and U4029 (N_4029,N_2076,N_2880);
nor U4030 (N_4030,N_3131,N_2491);
nand U4031 (N_4031,N_2560,N_3980);
or U4032 (N_4032,N_3361,N_2181);
nand U4033 (N_4033,N_3548,N_2661);
or U4034 (N_4034,N_2394,N_2792);
or U4035 (N_4035,N_3175,N_2937);
and U4036 (N_4036,N_2709,N_2192);
and U4037 (N_4037,N_3197,N_2779);
and U4038 (N_4038,N_2545,N_2755);
nand U4039 (N_4039,N_2455,N_2876);
or U4040 (N_4040,N_3498,N_3028);
or U4041 (N_4041,N_3221,N_2909);
and U4042 (N_4042,N_3256,N_3043);
and U4043 (N_4043,N_2927,N_3674);
and U4044 (N_4044,N_2780,N_3528);
nand U4045 (N_4045,N_3687,N_2199);
and U4046 (N_4046,N_2286,N_2162);
and U4047 (N_4047,N_2859,N_2460);
or U4048 (N_4048,N_3708,N_2631);
or U4049 (N_4049,N_3113,N_2402);
and U4050 (N_4050,N_2443,N_2719);
or U4051 (N_4051,N_3655,N_3753);
nand U4052 (N_4052,N_2478,N_3509);
nor U4053 (N_4053,N_2208,N_2765);
nor U4054 (N_4054,N_3271,N_2772);
and U4055 (N_4055,N_2431,N_2338);
and U4056 (N_4056,N_2810,N_2092);
nand U4057 (N_4057,N_3858,N_3592);
or U4058 (N_4058,N_2263,N_3122);
nand U4059 (N_4059,N_3441,N_3936);
nand U4060 (N_4060,N_2839,N_2607);
or U4061 (N_4061,N_2399,N_2131);
and U4062 (N_4062,N_3946,N_3025);
nand U4063 (N_4063,N_2959,N_3745);
or U4064 (N_4064,N_2116,N_3988);
nand U4065 (N_4065,N_3731,N_3672);
nand U4066 (N_4066,N_3564,N_2220);
nand U4067 (N_4067,N_2643,N_3097);
nor U4068 (N_4068,N_2337,N_3448);
nand U4069 (N_4069,N_3965,N_3715);
nand U4070 (N_4070,N_3922,N_2027);
nand U4071 (N_4071,N_2700,N_3570);
and U4072 (N_4072,N_2509,N_3832);
nor U4073 (N_4073,N_3538,N_3984);
nand U4074 (N_4074,N_3841,N_2356);
and U4075 (N_4075,N_2318,N_3608);
nand U4076 (N_4076,N_3363,N_3651);
nand U4077 (N_4077,N_3647,N_3485);
and U4078 (N_4078,N_3955,N_3360);
nor U4079 (N_4079,N_3285,N_3830);
nor U4080 (N_4080,N_2842,N_3295);
and U4081 (N_4081,N_3044,N_3154);
nand U4082 (N_4082,N_3174,N_2969);
or U4083 (N_4083,N_2712,N_3502);
and U4084 (N_4084,N_3557,N_2355);
nor U4085 (N_4085,N_2065,N_2050);
and U4086 (N_4086,N_3698,N_3755);
nand U4087 (N_4087,N_2456,N_2393);
and U4088 (N_4088,N_2507,N_2853);
nand U4089 (N_4089,N_3457,N_3738);
or U4090 (N_4090,N_3168,N_3928);
nor U4091 (N_4091,N_3637,N_3501);
nor U4092 (N_4092,N_3177,N_2999);
nand U4093 (N_4093,N_2469,N_2597);
or U4094 (N_4094,N_2036,N_2042);
nor U4095 (N_4095,N_2976,N_2943);
nor U4096 (N_4096,N_3091,N_3218);
and U4097 (N_4097,N_2482,N_2571);
nand U4098 (N_4098,N_3616,N_3325);
nor U4099 (N_4099,N_2276,N_3904);
nor U4100 (N_4100,N_2289,N_3159);
and U4101 (N_4101,N_2517,N_2905);
and U4102 (N_4102,N_3801,N_2840);
nor U4103 (N_4103,N_2487,N_2161);
nand U4104 (N_4104,N_3640,N_3911);
or U4105 (N_4105,N_2021,N_3932);
and U4106 (N_4106,N_2279,N_2492);
and U4107 (N_4107,N_2655,N_3278);
or U4108 (N_4108,N_3949,N_3701);
nand U4109 (N_4109,N_3549,N_3683);
nor U4110 (N_4110,N_2067,N_2864);
nand U4111 (N_4111,N_3491,N_3248);
or U4112 (N_4112,N_2372,N_3938);
nand U4113 (N_4113,N_2854,N_3891);
and U4114 (N_4114,N_2266,N_3976);
nand U4115 (N_4115,N_3873,N_3306);
or U4116 (N_4116,N_2615,N_3893);
nand U4117 (N_4117,N_2424,N_3080);
nand U4118 (N_4118,N_2973,N_3811);
nor U4119 (N_4119,N_2056,N_2923);
nor U4120 (N_4120,N_3395,N_3497);
or U4121 (N_4121,N_2101,N_3193);
and U4122 (N_4122,N_2107,N_3371);
nor U4123 (N_4123,N_2757,N_3983);
nor U4124 (N_4124,N_2419,N_2401);
nor U4125 (N_4125,N_3297,N_3269);
nand U4126 (N_4126,N_2771,N_3446);
and U4127 (N_4127,N_2446,N_3188);
or U4128 (N_4128,N_2426,N_3462);
or U4129 (N_4129,N_3684,N_3558);
or U4130 (N_4130,N_2762,N_3885);
nand U4131 (N_4131,N_2459,N_3664);
or U4132 (N_4132,N_2415,N_3789);
or U4133 (N_4133,N_2883,N_2573);
and U4134 (N_4134,N_2196,N_2519);
nor U4135 (N_4135,N_3861,N_3522);
or U4136 (N_4136,N_3597,N_3894);
nor U4137 (N_4137,N_2233,N_2601);
or U4138 (N_4138,N_3317,N_2895);
nor U4139 (N_4139,N_3078,N_2984);
and U4140 (N_4140,N_3240,N_3077);
nand U4141 (N_4141,N_3896,N_2906);
nand U4142 (N_4142,N_3607,N_3048);
or U4143 (N_4143,N_3052,N_3614);
nor U4144 (N_4144,N_3042,N_2530);
and U4145 (N_4145,N_2499,N_2423);
or U4146 (N_4146,N_3427,N_3732);
or U4147 (N_4147,N_2805,N_2201);
nor U4148 (N_4148,N_3493,N_3393);
or U4149 (N_4149,N_3369,N_2114);
and U4150 (N_4150,N_2480,N_2777);
nor U4151 (N_4151,N_3797,N_2711);
nor U4152 (N_4152,N_2246,N_3807);
or U4153 (N_4153,N_2879,N_3082);
or U4154 (N_4154,N_2011,N_2468);
nor U4155 (N_4155,N_2139,N_3694);
and U4156 (N_4156,N_3827,N_3200);
or U4157 (N_4157,N_3585,N_2595);
nand U4158 (N_4158,N_3442,N_3423);
or U4159 (N_4159,N_2591,N_2288);
or U4160 (N_4160,N_2685,N_2942);
nor U4161 (N_4161,N_3160,N_3249);
nor U4162 (N_4162,N_2664,N_2054);
or U4163 (N_4163,N_3888,N_3757);
nand U4164 (N_4164,N_2062,N_2292);
and U4165 (N_4165,N_3957,N_3103);
nor U4166 (N_4166,N_2638,N_2120);
nor U4167 (N_4167,N_2458,N_3410);
nor U4168 (N_4168,N_3776,N_2881);
xor U4169 (N_4169,N_2869,N_2911);
nand U4170 (N_4170,N_2163,N_2970);
nor U4171 (N_4171,N_2518,N_2158);
nor U4172 (N_4172,N_3405,N_3967);
nor U4173 (N_4173,N_3587,N_3128);
and U4174 (N_4174,N_3610,N_3606);
nor U4175 (N_4175,N_3316,N_3034);
and U4176 (N_4176,N_2537,N_2612);
nor U4177 (N_4177,N_3966,N_3087);
or U4178 (N_4178,N_3161,N_3951);
and U4179 (N_4179,N_3670,N_3959);
nor U4180 (N_4180,N_3436,N_3336);
nand U4181 (N_4181,N_2955,N_2602);
nor U4182 (N_4182,N_3320,N_3675);
nor U4183 (N_4183,N_2294,N_3473);
and U4184 (N_4184,N_3870,N_3009);
xor U4185 (N_4185,N_3308,N_2362);
nor U4186 (N_4186,N_3378,N_2115);
nor U4187 (N_4187,N_2714,N_2781);
and U4188 (N_4188,N_2211,N_3004);
and U4189 (N_4189,N_2407,N_3781);
nand U4190 (N_4190,N_2678,N_3150);
nand U4191 (N_4191,N_2982,N_2849);
nor U4192 (N_4192,N_2872,N_3429);
nor U4193 (N_4193,N_2369,N_2374);
and U4194 (N_4194,N_3345,N_2658);
nand U4195 (N_4195,N_3581,N_3808);
nand U4196 (N_4196,N_3513,N_3389);
or U4197 (N_4197,N_2704,N_2531);
nor U4198 (N_4198,N_2441,N_2740);
or U4199 (N_4199,N_3507,N_3318);
and U4200 (N_4200,N_3902,N_2185);
nor U4201 (N_4201,N_3440,N_2527);
nand U4202 (N_4202,N_2662,N_2699);
and U4203 (N_4203,N_2555,N_3580);
nor U4204 (N_4204,N_2690,N_2089);
nand U4205 (N_4205,N_3997,N_3703);
nand U4206 (N_4206,N_2835,N_3905);
nand U4207 (N_4207,N_3254,N_2551);
and U4208 (N_4208,N_2766,N_3677);
and U4209 (N_4209,N_2317,N_2322);
or U4210 (N_4210,N_2514,N_3415);
nor U4211 (N_4211,N_3018,N_3426);
or U4212 (N_4212,N_2748,N_3601);
or U4213 (N_4213,N_3815,N_2633);
and U4214 (N_4214,N_2086,N_2308);
nand U4215 (N_4215,N_3104,N_3969);
or U4216 (N_4216,N_3996,N_3892);
nand U4217 (N_4217,N_3045,N_2617);
and U4218 (N_4218,N_3234,N_3418);
and U4219 (N_4219,N_3213,N_3192);
nor U4220 (N_4220,N_3619,N_3981);
and U4221 (N_4221,N_3973,N_2910);
or U4222 (N_4222,N_2032,N_2410);
xnor U4223 (N_4223,N_2102,N_3481);
or U4224 (N_4224,N_3076,N_3229);
nor U4225 (N_4225,N_2698,N_3276);
and U4226 (N_4226,N_2972,N_2465);
or U4227 (N_4227,N_2243,N_2717);
nor U4228 (N_4228,N_2341,N_3722);
or U4229 (N_4229,N_3833,N_2417);
and U4230 (N_4230,N_2437,N_2668);
nor U4231 (N_4231,N_2019,N_2304);
and U4232 (N_4232,N_2146,N_2098);
nand U4233 (N_4233,N_2467,N_2386);
xor U4234 (N_4234,N_3994,N_3382);
or U4235 (N_4235,N_2406,N_2368);
and U4236 (N_4236,N_2033,N_3322);
or U4237 (N_4237,N_3280,N_2600);
and U4238 (N_4238,N_2091,N_2111);
nand U4239 (N_4239,N_2037,N_3086);
or U4240 (N_4240,N_2747,N_2015);
or U4241 (N_4241,N_3525,N_3559);
or U4242 (N_4242,N_2838,N_2819);
nor U4243 (N_4243,N_3059,N_3073);
nor U4244 (N_4244,N_2347,N_2309);
and U4245 (N_4245,N_2521,N_2626);
and U4246 (N_4246,N_2544,N_3186);
nor U4247 (N_4247,N_3147,N_3995);
and U4248 (N_4248,N_2630,N_3825);
or U4249 (N_4249,N_2414,N_3682);
and U4250 (N_4250,N_2803,N_3214);
nor U4251 (N_4251,N_3014,N_3339);
nor U4252 (N_4252,N_3107,N_3477);
and U4253 (N_4253,N_2759,N_2339);
or U4254 (N_4254,N_2344,N_3390);
or U4255 (N_4255,N_2857,N_2109);
nand U4256 (N_4256,N_2252,N_2946);
nand U4257 (N_4257,N_3692,N_2147);
or U4258 (N_4258,N_2776,N_2725);
and U4259 (N_4259,N_2950,N_3895);
or U4260 (N_4260,N_3913,N_3835);
or U4261 (N_4261,N_2398,N_3281);
nor U4262 (N_4262,N_3829,N_2121);
and U4263 (N_4263,N_2085,N_3183);
nand U4264 (N_4264,N_2488,N_3296);
nand U4265 (N_4265,N_2496,N_3544);
and U4266 (N_4266,N_2082,N_2242);
nor U4267 (N_4267,N_2649,N_2815);
and U4268 (N_4268,N_3621,N_2583);
or U4269 (N_4269,N_3000,N_2951);
or U4270 (N_4270,N_2094,N_2651);
nand U4271 (N_4271,N_3632,N_2957);
and U4272 (N_4272,N_3706,N_2045);
nand U4273 (N_4273,N_3482,N_3774);
nor U4274 (N_4274,N_2793,N_2845);
nor U4275 (N_4275,N_3739,N_3541);
nand U4276 (N_4276,N_2886,N_3085);
nand U4277 (N_4277,N_2014,N_3487);
or U4278 (N_4278,N_3535,N_3618);
nor U4279 (N_4279,N_2647,N_3024);
and U4280 (N_4280,N_2035,N_3579);
or U4281 (N_4281,N_3720,N_3596);
or U4282 (N_4282,N_2827,N_3734);
and U4283 (N_4283,N_3121,N_2063);
nand U4284 (N_4284,N_3617,N_3189);
xnor U4285 (N_4285,N_2817,N_3124);
or U4286 (N_4286,N_3822,N_2635);
nor U4287 (N_4287,N_2164,N_2058);
and U4288 (N_4288,N_2599,N_2787);
or U4289 (N_4289,N_3421,N_3689);
or U4290 (N_4290,N_2898,N_3236);
or U4291 (N_4291,N_3464,N_3201);
nor U4292 (N_4292,N_2742,N_3003);
and U4293 (N_4293,N_2479,N_2202);
nand U4294 (N_4294,N_3066,N_2687);
and U4295 (N_4295,N_3093,N_2737);
nand U4296 (N_4296,N_3479,N_2379);
nor U4297 (N_4297,N_3212,N_3869);
and U4298 (N_4298,N_3132,N_2924);
nor U4299 (N_4299,N_3726,N_3404);
nor U4300 (N_4300,N_2302,N_3241);
and U4301 (N_4301,N_2157,N_2052);
or U4302 (N_4302,N_2475,N_3071);
or U4303 (N_4303,N_3293,N_2088);
nand U4304 (N_4304,N_2296,N_2893);
nand U4305 (N_4305,N_2580,N_3046);
nor U4306 (N_4306,N_3784,N_3709);
or U4307 (N_4307,N_3862,N_3927);
or U4308 (N_4308,N_3785,N_3488);
and U4309 (N_4309,N_2642,N_3347);
and U4310 (N_4310,N_2295,N_3163);
or U4311 (N_4311,N_3842,N_2452);
and U4312 (N_4312,N_3406,N_2108);
nor U4313 (N_4313,N_2112,N_3217);
nand U4314 (N_4314,N_2697,N_2176);
and U4315 (N_4315,N_3717,N_3411);
or U4316 (N_4316,N_2044,N_3206);
nand U4317 (N_4317,N_3403,N_2450);
and U4318 (N_4318,N_3070,N_3391);
nand U4319 (N_4319,N_3162,N_2980);
nand U4320 (N_4320,N_3349,N_3257);
nor U4321 (N_4321,N_3056,N_3736);
and U4322 (N_4322,N_3484,N_2659);
nor U4323 (N_4323,N_3678,N_2129);
and U4324 (N_4324,N_3941,N_3286);
nand U4325 (N_4325,N_2562,N_2669);
and U4326 (N_4326,N_3247,N_2038);
nor U4327 (N_4327,N_2511,N_3323);
nand U4328 (N_4328,N_2281,N_3845);
nand U4329 (N_4329,N_3699,N_2320);
and U4330 (N_4330,N_2938,N_2075);
nor U4331 (N_4331,N_3151,N_3718);
nor U4332 (N_4332,N_2917,N_2209);
nor U4333 (N_4333,N_3230,N_3510);
or U4334 (N_4334,N_3875,N_3496);
nand U4335 (N_4335,N_3114,N_3645);
nand U4336 (N_4336,N_2170,N_3723);
nand U4337 (N_4337,N_3775,N_3083);
nand U4338 (N_4338,N_2123,N_2148);
or U4339 (N_4339,N_3026,N_3622);
nand U4340 (N_4340,N_2614,N_3139);
and U4341 (N_4341,N_2609,N_3642);
nand U4342 (N_4342,N_3176,N_3555);
nor U4343 (N_4343,N_3072,N_3765);
or U4344 (N_4344,N_2553,N_3790);
nor U4345 (N_4345,N_2724,N_3989);
nand U4346 (N_4346,N_3294,N_2439);
or U4347 (N_4347,N_2383,N_3846);
and U4348 (N_4348,N_3279,N_3005);
nor U4349 (N_4349,N_3237,N_3847);
and U4350 (N_4350,N_3676,N_2730);
and U4351 (N_4351,N_2168,N_3474);
or U4352 (N_4352,N_3324,N_2770);
nand U4353 (N_4353,N_2000,N_3761);
or U4354 (N_4354,N_2169,N_3542);
nor U4355 (N_4355,N_2047,N_2542);
or U4356 (N_4356,N_3916,N_3179);
and U4357 (N_4357,N_2870,N_2582);
and U4358 (N_4358,N_3012,N_3215);
xor U4359 (N_4359,N_2673,N_2213);
or U4360 (N_4360,N_2871,N_2941);
xnor U4361 (N_4361,N_3724,N_2693);
nor U4362 (N_4362,N_2641,N_2193);
and U4363 (N_4363,N_2746,N_2505);
or U4364 (N_4364,N_2016,N_2675);
and U4365 (N_4365,N_3744,N_2851);
nand U4366 (N_4366,N_2897,N_3780);
xor U4367 (N_4367,N_2652,N_3854);
and U4368 (N_4368,N_3534,N_3291);
nand U4369 (N_4369,N_2506,N_2986);
nand U4370 (N_4370,N_2855,N_2150);
or U4371 (N_4371,N_3639,N_2022);
or U4372 (N_4372,N_2928,N_3490);
nor U4373 (N_4373,N_3313,N_3547);
or U4374 (N_4374,N_2274,N_3660);
and U4375 (N_4375,N_2814,N_3187);
nand U4376 (N_4376,N_3629,N_2397);
nor U4377 (N_4377,N_2490,N_3918);
nor U4378 (N_4378,N_2875,N_2282);
or U4379 (N_4379,N_2723,N_3173);
nand U4380 (N_4380,N_2624,N_3565);
nand U4381 (N_4381,N_3962,N_2945);
and U4382 (N_4382,N_2061,N_2336);
and U4383 (N_4383,N_2884,N_3728);
or U4384 (N_4384,N_3799,N_2570);
and U4385 (N_4385,N_2964,N_2829);
or U4386 (N_4386,N_3567,N_3330);
and U4387 (N_4387,N_3144,N_2918);
nand U4388 (N_4388,N_3233,N_2285);
nor U4389 (N_4389,N_3275,N_2900);
or U4390 (N_4390,N_2733,N_3588);
or U4391 (N_4391,N_2447,N_2370);
and U4392 (N_4392,N_3392,N_2914);
or U4393 (N_4393,N_2313,N_2667);
and U4394 (N_4394,N_2682,N_2833);
nor U4395 (N_4395,N_3613,N_2994);
nand U4396 (N_4396,N_3524,N_2843);
nor U4397 (N_4397,N_2761,N_2299);
and U4398 (N_4398,N_2497,N_2745);
nand U4399 (N_4399,N_2563,N_2874);
or U4400 (N_4400,N_3563,N_3716);
nand U4401 (N_4401,N_2913,N_2798);
or U4402 (N_4402,N_3855,N_2696);
and U4403 (N_4403,N_2809,N_3120);
or U4404 (N_4404,N_3770,N_3149);
nand U4405 (N_4405,N_3352,N_2405);
nor U4406 (N_4406,N_3374,N_2348);
and U4407 (N_4407,N_3036,N_2221);
and U4408 (N_4408,N_2436,N_2576);
and U4409 (N_4409,N_3050,N_2239);
and U4410 (N_4410,N_3864,N_3809);
and U4411 (N_4411,N_3400,N_3993);
and U4412 (N_4412,N_2858,N_2182);
and U4413 (N_4413,N_2837,N_3520);
nand U4414 (N_4414,N_3117,N_2671);
or U4415 (N_4415,N_3863,N_2411);
nor U4416 (N_4416,N_2903,N_2095);
and U4417 (N_4417,N_2180,N_2550);
nor U4418 (N_4418,N_2194,N_2464);
or U4419 (N_4419,N_3839,N_3730);
nor U4420 (N_4420,N_3387,N_3551);
nor U4421 (N_4421,N_2760,N_3469);
nand U4422 (N_4422,N_2080,N_3310);
or U4423 (N_4423,N_2778,N_2218);
nand U4424 (N_4424,N_3992,N_2451);
nor U4425 (N_4425,N_3417,N_2782);
or U4426 (N_4426,N_3968,N_2680);
xor U4427 (N_4427,N_3511,N_3106);
nand U4428 (N_4428,N_2862,N_3466);
nand U4429 (N_4429,N_3679,N_2967);
and U4430 (N_4430,N_3057,N_3595);
xor U4431 (N_4431,N_3216,N_3714);
nand U4432 (N_4432,N_3243,N_3032);
nand U4433 (N_4433,N_2473,N_3690);
nor U4434 (N_4434,N_2387,N_2919);
nor U4435 (N_4435,N_2672,N_2818);
or U4436 (N_4436,N_2526,N_2297);
or U4437 (N_4437,N_2977,N_3455);
nor U4438 (N_4438,N_3878,N_2841);
or U4439 (N_4439,N_3628,N_3630);
or U4440 (N_4440,N_3859,N_3460);
nand U4441 (N_4441,N_2822,N_3831);
and U4442 (N_4442,N_2418,N_2828);
or U4443 (N_4443,N_3654,N_3897);
nor U4444 (N_4444,N_3794,N_2223);
and U4445 (N_4445,N_2028,N_2229);
nand U4446 (N_4446,N_3386,N_3136);
or U4447 (N_4447,N_2084,N_3681);
nand U4448 (N_4448,N_3523,N_2254);
or U4449 (N_4449,N_2785,N_3376);
and U4450 (N_4450,N_2413,N_3643);
or U4451 (N_4451,N_2603,N_3612);
or U4452 (N_4452,N_3971,N_3866);
nand U4453 (N_4453,N_3519,N_3424);
xnor U4454 (N_4454,N_2001,N_2224);
nand U4455 (N_4455,N_2427,N_3633);
nor U4456 (N_4456,N_3700,N_3798);
nor U4457 (N_4457,N_2449,N_2342);
xor U4458 (N_4458,N_2325,N_3646);
nor U4459 (N_4459,N_3449,N_2915);
or U4460 (N_4460,N_2357,N_3963);
nand U4461 (N_4461,N_3625,N_2593);
nor U4462 (N_4462,N_3506,N_3209);
and U4463 (N_4463,N_3751,N_2093);
nor U4464 (N_4464,N_2264,N_3975);
xnor U4465 (N_4465,N_2152,N_2728);
xor U4466 (N_4466,N_3047,N_2645);
or U4467 (N_4467,N_2825,N_3574);
xor U4468 (N_4468,N_2960,N_3252);
or U4469 (N_4469,N_2259,N_3244);
or U4470 (N_4470,N_3985,N_3270);
and U4471 (N_4471,N_2899,N_3958);
and U4472 (N_4472,N_2486,N_2996);
nor U4473 (N_4473,N_3433,N_2269);
xnor U4474 (N_4474,N_2908,N_3268);
or U4475 (N_4475,N_3431,N_2271);
nand U4476 (N_4476,N_2234,N_3334);
and U4477 (N_4477,N_2217,N_3088);
or U4478 (N_4478,N_3029,N_2978);
and U4479 (N_4479,N_3346,N_2632);
and U4480 (N_4480,N_2018,N_3169);
nand U4481 (N_4481,N_3550,N_2261);
and U4482 (N_4482,N_3274,N_2256);
nand U4483 (N_4483,N_2278,N_3521);
or U4484 (N_4484,N_3364,N_2377);
or U4485 (N_4485,N_3990,N_3857);
nand U4486 (N_4486,N_3263,N_2691);
and U4487 (N_4487,N_2504,N_3022);
or U4488 (N_4488,N_3397,N_3589);
nor U4489 (N_4489,N_3053,N_3101);
or U4490 (N_4490,N_3450,N_2113);
or U4491 (N_4491,N_2625,N_2547);
or U4492 (N_4492,N_3710,N_2183);
nor U4493 (N_4493,N_2998,N_3537);
nand U4494 (N_4494,N_3152,N_3351);
or U4495 (N_4495,N_3428,N_3035);
or U4496 (N_4496,N_3593,N_3368);
and U4497 (N_4497,N_3196,N_3590);
nand U4498 (N_4498,N_2366,N_3327);
and U4499 (N_4499,N_3008,N_3090);
nor U4500 (N_4500,N_3365,N_3583);
and U4501 (N_4501,N_2442,N_2608);
nor U4502 (N_4502,N_3702,N_3020);
or U4503 (N_4503,N_2440,N_2686);
nand U4504 (N_4504,N_3923,N_3220);
and U4505 (N_4505,N_3019,N_2865);
nand U4506 (N_4506,N_2137,N_2351);
nand U4507 (N_4507,N_3470,N_2749);
and U4508 (N_4508,N_2557,N_2890);
nor U4509 (N_4509,N_2363,N_2713);
or U4510 (N_4510,N_3153,N_3649);
nand U4511 (N_4511,N_3309,N_2750);
nand U4512 (N_4512,N_2319,N_3972);
or U4513 (N_4513,N_3225,N_3594);
and U4514 (N_4514,N_3366,N_2953);
nand U4515 (N_4515,N_3609,N_3974);
xor U4516 (N_4516,N_3027,N_2581);
and U4517 (N_4517,N_3231,N_3903);
nor U4518 (N_4518,N_2244,N_2207);
or U4519 (N_4519,N_2333,N_2284);
and U4520 (N_4520,N_3582,N_3166);
nor U4521 (N_4521,N_3385,N_2706);
and U4522 (N_4522,N_2813,N_3791);
and U4523 (N_4523,N_2797,N_3850);
nand U4524 (N_4524,N_3573,N_2189);
nor U4525 (N_4525,N_2820,N_2247);
and U4526 (N_4526,N_2435,N_2710);
nor U4527 (N_4527,N_3661,N_3194);
and U4528 (N_4528,N_2589,N_3514);
nor U4529 (N_4529,N_3991,N_2151);
xnor U4530 (N_4530,N_3930,N_3806);
or U4531 (N_4531,N_3624,N_3853);
nand U4532 (N_4532,N_2334,N_2756);
and U4533 (N_4533,N_2734,N_2907);
nand U4534 (N_4534,N_3223,N_2445);
nor U4535 (N_4535,N_3098,N_2026);
nand U4536 (N_4536,N_3826,N_2305);
or U4537 (N_4537,N_3326,N_3062);
nand U4538 (N_4538,N_2006,N_3171);
and U4539 (N_4539,N_2323,N_3865);
nand U4540 (N_4540,N_3074,N_3148);
or U4541 (N_4541,N_2744,N_3486);
and U4542 (N_4542,N_2009,N_2390);
nor U4543 (N_4543,N_3760,N_2057);
and U4544 (N_4544,N_2948,N_3222);
nand U4545 (N_4545,N_2471,N_3133);
or U4546 (N_4546,N_3603,N_2572);
nand U4547 (N_4547,N_3729,N_2536);
nand U4548 (N_4548,N_2380,N_2741);
or U4549 (N_4549,N_2789,N_2767);
or U4550 (N_4550,N_2392,N_3977);
and U4551 (N_4551,N_2764,N_2352);
nor U4552 (N_4552,N_3685,N_2421);
or U4553 (N_4553,N_2922,N_3879);
nand U4554 (N_4554,N_2606,N_3359);
or U4555 (N_4555,N_3172,N_3416);
nand U4556 (N_4556,N_3251,N_2204);
nand U4557 (N_4557,N_3953,N_3238);
or U4558 (N_4558,N_3123,N_2214);
or U4559 (N_4559,N_3413,N_2823);
nor U4560 (N_4560,N_2171,N_3657);
nor U4561 (N_4561,N_2552,N_2694);
nor U4562 (N_4562,N_3711,N_2375);
nor U4563 (N_4563,N_3401,N_2203);
xnor U4564 (N_4564,N_2916,N_3265);
nor U4565 (N_4565,N_3627,N_3586);
nor U4566 (N_4566,N_3912,N_3210);
and U4567 (N_4567,N_2125,N_3882);
nor U4568 (N_4568,N_2079,N_3979);
nand U4569 (N_4569,N_3435,N_3602);
nor U4570 (N_4570,N_2901,N_3503);
nor U4571 (N_4571,N_3051,N_3680);
nor U4572 (N_4572,N_2934,N_3157);
nand U4573 (N_4573,N_2408,N_2270);
or U4574 (N_4574,N_2388,N_2077);
and U4575 (N_4575,N_2083,N_2328);
or U4576 (N_4576,N_2238,N_3362);
nor U4577 (N_4577,N_3707,N_3467);
nor U4578 (N_4578,N_3058,N_2307);
nand U4579 (N_4579,N_3611,N_2160);
nand U4580 (N_4580,N_3735,N_2359);
nand U4581 (N_4581,N_2060,N_2995);
or U4582 (N_4582,N_2025,N_2949);
or U4583 (N_4583,N_3793,N_2689);
nand U4584 (N_4584,N_2989,N_3170);
nor U4585 (N_4585,N_3060,N_3552);
or U4586 (N_4586,N_3096,N_3877);
nand U4587 (N_4587,N_2007,N_2024);
nand U4588 (N_4588,N_3067,N_2844);
xor U4589 (N_4589,N_3112,N_2997);
or U4590 (N_4590,N_2412,N_2739);
and U4591 (N_4591,N_2726,N_2971);
or U4592 (N_4592,N_3227,N_2130);
nor U4593 (N_4593,N_3636,N_3890);
nor U4594 (N_4594,N_3653,N_3505);
nand U4595 (N_4595,N_2605,N_2821);
nor U4596 (N_4596,N_2364,N_2041);
and U4597 (N_4597,N_3752,N_2522);
nor U4598 (N_4598,N_3940,N_2290);
nand U4599 (N_4599,N_3964,N_3099);
nand U4600 (N_4600,N_2866,N_2523);
nand U4601 (N_4601,N_2665,N_2312);
nand U4602 (N_4602,N_2005,N_3756);
or U4603 (N_4603,N_3658,N_3224);
nor U4604 (N_4604,N_3768,N_3178);
nand U4605 (N_4605,N_2097,N_3394);
nor U4606 (N_4606,N_2251,N_2987);
nor U4607 (N_4607,N_2738,N_2087);
or U4608 (N_4608,N_2034,N_3805);
nand U4609 (N_4609,N_2262,N_2186);
nor U4610 (N_4610,N_3130,N_3041);
and U4611 (N_4611,N_3033,N_2768);
or U4612 (N_4612,N_2935,N_3412);
nand U4613 (N_4613,N_2769,N_3343);
or U4614 (N_4614,N_2513,N_3463);
and U4615 (N_4615,N_2975,N_3970);
nor U4616 (N_4616,N_2167,N_2330);
nor U4617 (N_4617,N_3228,N_2887);
and U4618 (N_4618,N_3821,N_2117);
nor U4619 (N_4619,N_3942,N_2684);
and U4620 (N_4620,N_3571,N_3377);
or U4621 (N_4621,N_3615,N_3315);
or U4622 (N_4622,N_2483,N_3771);
and U4623 (N_4623,N_2064,N_3591);
and U4624 (N_4624,N_2554,N_3697);
or U4625 (N_4625,N_2461,N_2140);
nand U4626 (N_4626,N_3749,N_3190);
or U4627 (N_4627,N_3471,N_3673);
nor U4628 (N_4628,N_3817,N_3358);
or U4629 (N_4629,N_2735,N_3526);
or U4630 (N_4630,N_3898,N_3907);
nor U4631 (N_4631,N_2345,N_3909);
or U4632 (N_4632,N_2260,N_3813);
or U4633 (N_4633,N_2968,N_2830);
or U4634 (N_4634,N_2628,N_3527);
or U4635 (N_4635,N_3876,N_2031);
nor U4636 (N_4636,N_2850,N_2882);
or U4637 (N_4637,N_3667,N_2620);
and U4638 (N_4638,N_2929,N_3290);
and U4639 (N_4639,N_2873,N_2543);
xnor U4640 (N_4640,N_2799,N_2613);
xnor U4641 (N_4641,N_2800,N_2273);
or U4642 (N_4642,N_3758,N_2053);
nand U4643 (N_4643,N_3388,N_3540);
and U4644 (N_4644,N_2637,N_2758);
nor U4645 (N_4645,N_3476,N_2718);
nand U4646 (N_4646,N_2867,N_3191);
xnor U4647 (N_4647,N_2653,N_2559);
nand U4648 (N_4648,N_2072,N_3712);
nand U4649 (N_4649,N_2049,N_3235);
or U4650 (N_4650,N_3219,N_3883);
nand U4651 (N_4651,N_3348,N_2891);
xor U4652 (N_4652,N_3860,N_3328);
nand U4653 (N_4653,N_2051,N_2763);
nor U4654 (N_4654,N_2640,N_3828);
or U4655 (N_4655,N_3508,N_3226);
xnor U4656 (N_4656,N_2836,N_3370);
nor U4657 (N_4657,N_3100,N_2683);
or U4658 (N_4658,N_3115,N_2020);
or U4659 (N_4659,N_2122,N_3084);
or U4660 (N_4660,N_3465,N_2592);
nand U4661 (N_4661,N_2248,N_2629);
nor U4662 (N_4662,N_2433,N_3788);
nor U4663 (N_4663,N_2099,N_2892);
and U4664 (N_4664,N_2743,N_2070);
or U4665 (N_4665,N_3432,N_2291);
and U4666 (N_4666,N_2524,N_2991);
or U4667 (N_4667,N_2802,N_2241);
or U4668 (N_4668,N_2481,N_3094);
or U4669 (N_4669,N_3599,N_2226);
nor U4670 (N_4670,N_2878,N_3844);
nor U4671 (N_4671,N_3943,N_3648);
nor U4672 (N_4672,N_3998,N_3232);
nor U4673 (N_4673,N_2979,N_3638);
nand U4674 (N_4674,N_3631,N_3329);
or U4675 (N_4675,N_2232,N_2110);
nand U4676 (N_4676,N_3626,N_3303);
and U4677 (N_4677,N_3773,N_3665);
and U4678 (N_4678,N_2752,N_2143);
xor U4679 (N_4679,N_2727,N_3447);
and U4680 (N_4680,N_2255,N_2237);
nor U4681 (N_4681,N_3007,N_3553);
or U4682 (N_4682,N_3783,N_2587);
or U4683 (N_4683,N_3407,N_2932);
and U4684 (N_4684,N_2846,N_2416);
nand U4685 (N_4685,N_2267,N_3874);
nand U4686 (N_4686,N_3604,N_2944);
xnor U4687 (N_4687,N_2327,N_2376);
or U4688 (N_4688,N_3489,N_2566);
or U4689 (N_4689,N_3198,N_3443);
and U4690 (N_4690,N_2773,N_3284);
or U4691 (N_4691,N_2353,N_3367);
and U4692 (N_4692,N_2634,N_2705);
nand U4693 (N_4693,N_2275,N_2155);
or U4694 (N_4694,N_3292,N_2230);
or U4695 (N_4695,N_2154,N_3620);
xor U4696 (N_4696,N_3332,N_3341);
nand U4697 (N_4697,N_2993,N_2500);
and U4698 (N_4698,N_3695,N_3924);
or U4699 (N_4699,N_3314,N_3748);
and U4700 (N_4700,N_2470,N_3372);
and U4701 (N_4701,N_3444,N_2179);
nand U4702 (N_4702,N_3021,N_3641);
or U4703 (N_4703,N_3516,N_3158);
or U4704 (N_4704,N_3384,N_3434);
nand U4705 (N_4705,N_2391,N_2774);
or U4706 (N_4706,N_3092,N_3944);
nand U4707 (N_4707,N_3623,N_2540);
or U4708 (N_4708,N_3422,N_2753);
and U4709 (N_4709,N_2736,N_3945);
nand U4710 (N_4710,N_2852,N_3272);
nand U4711 (N_4711,N_2961,N_3333);
and U4712 (N_4712,N_2508,N_3451);
nor U4713 (N_4713,N_3305,N_2963);
or U4714 (N_4714,N_2503,N_2729);
nand U4715 (N_4715,N_3258,N_2231);
nor U4716 (N_4716,N_2751,N_3311);
nor U4717 (N_4717,N_3956,N_2303);
or U4718 (N_4718,N_3635,N_3302);
or U4719 (N_4719,N_3545,N_3001);
nor U4720 (N_4720,N_3802,N_3438);
nand U4721 (N_4721,N_3764,N_3242);
or U4722 (N_4722,N_3299,N_2175);
and U4723 (N_4723,N_3145,N_2434);
nor U4724 (N_4724,N_2832,N_3480);
or U4725 (N_4725,N_2623,N_2293);
or U4726 (N_4726,N_3662,N_3886);
xor U4727 (N_4727,N_3575,N_2806);
or U4728 (N_4728,N_2564,N_3778);
nor U4729 (N_4729,N_2444,N_3906);
xnor U4730 (N_4730,N_3782,N_2191);
nand U4731 (N_4731,N_3307,N_2974);
nand U4732 (N_4732,N_2621,N_2956);
or U4733 (N_4733,N_2432,N_3843);
and U4734 (N_4734,N_2801,N_3396);
nor U4735 (N_4735,N_2834,N_3691);
or U4736 (N_4736,N_3512,N_3253);
nand U4737 (N_4737,N_3634,N_2596);
or U4738 (N_4738,N_3135,N_3536);
nor U4739 (N_4739,N_3260,N_3931);
nand U4740 (N_4740,N_2716,N_3156);
xnor U4741 (N_4741,N_2378,N_2796);
and U4742 (N_4742,N_3246,N_2586);
nor U4743 (N_4743,N_2495,N_2775);
nand U4744 (N_4744,N_3705,N_2816);
and U4745 (N_4745,N_2422,N_2066);
or U4746 (N_4746,N_3203,N_3065);
or U4747 (N_4747,N_3713,N_2489);
nor U4748 (N_4748,N_2132,N_3182);
nor U4749 (N_4749,N_2794,N_3023);
or U4750 (N_4750,N_2396,N_3787);
or U4751 (N_4751,N_2791,N_3999);
nor U4752 (N_4752,N_2529,N_3185);
and U4753 (N_4753,N_2280,N_3109);
nand U4754 (N_4754,N_3578,N_2074);
nor U4755 (N_4755,N_3075,N_3650);
and U4756 (N_4756,N_3814,N_2936);
nand U4757 (N_4757,N_3719,N_3452);
nor U4758 (N_4758,N_2205,N_2860);
nor U4759 (N_4759,N_3011,N_3952);
nand U4760 (N_4760,N_2350,N_2732);
and U4761 (N_4761,N_2636,N_3848);
and U4762 (N_4762,N_3577,N_2585);
or U4763 (N_4763,N_3211,N_3600);
nor U4764 (N_4764,N_2611,N_3354);
or U4765 (N_4765,N_3483,N_2863);
nor U4766 (N_4766,N_2720,N_3747);
nand U4767 (N_4767,N_3155,N_2287);
or U4768 (N_4768,N_3127,N_3824);
nor U4769 (N_4769,N_2992,N_3960);
and U4770 (N_4770,N_2314,N_2043);
nor U4771 (N_4771,N_2466,N_2940);
or U4772 (N_4772,N_2198,N_2485);
nand U4773 (N_4773,N_3871,N_2174);
nand U4774 (N_4774,N_3380,N_2474);
nor U4775 (N_4775,N_3129,N_3381);
nand U4776 (N_4776,N_2650,N_2676);
nand U4777 (N_4777,N_3054,N_3357);
nor U4778 (N_4778,N_2933,N_2361);
or U4779 (N_4779,N_2215,N_3414);
nor U4780 (N_4780,N_2448,N_2688);
nand U4781 (N_4781,N_2100,N_3688);
and U4782 (N_4782,N_2298,N_3978);
nor U4783 (N_4783,N_2172,N_2354);
or U4784 (N_4784,N_3666,N_2498);
or U4785 (N_4785,N_2788,N_3934);
or U4786 (N_4786,N_3468,N_3379);
nor U4787 (N_4787,N_2081,N_2128);
nand U4788 (N_4788,N_2888,N_2861);
or U4789 (N_4789,N_3566,N_3030);
nand U4790 (N_4790,N_2590,N_3935);
xnor U4791 (N_4791,N_2463,N_3277);
nand U4792 (N_4792,N_2385,N_3917);
nand U4793 (N_4793,N_3420,N_3013);
or U4794 (N_4794,N_3803,N_2538);
nor U4795 (N_4795,N_3063,N_2939);
nand U4796 (N_4796,N_3543,N_2124);
or U4797 (N_4797,N_3759,N_2331);
and U4798 (N_4798,N_2721,N_3560);
nand U4799 (N_4799,N_3425,N_3880);
and U4800 (N_4800,N_3002,N_3742);
nor U4801 (N_4801,N_2604,N_2654);
nor U4802 (N_4802,N_3398,N_2666);
nand U4803 (N_4803,N_3663,N_3725);
xnor U4804 (N_4804,N_2657,N_2227);
nor U4805 (N_4805,N_2681,N_2301);
nor U4806 (N_4806,N_2178,N_3914);
and U4807 (N_4807,N_3852,N_2384);
or U4808 (N_4808,N_3750,N_2588);
nor U4809 (N_4809,N_3652,N_2187);
and U4810 (N_4810,N_2454,N_3454);
and U4811 (N_4811,N_2340,N_3165);
or U4812 (N_4812,N_2677,N_2030);
nand U4813 (N_4813,N_2277,N_2786);
and U4814 (N_4814,N_2925,N_2197);
or U4815 (N_4815,N_3915,N_3068);
and U4816 (N_4816,N_3539,N_2539);
xnor U4817 (N_4817,N_3119,N_2920);
nand U4818 (N_4818,N_3300,N_2166);
nor U4819 (N_4819,N_3267,N_2804);
or U4820 (N_4820,N_2145,N_2040);
nand U4821 (N_4821,N_3763,N_3383);
nor U4822 (N_4822,N_3772,N_2225);
or U4823 (N_4823,N_3430,N_2472);
nor U4824 (N_4824,N_3146,N_3402);
and U4825 (N_4825,N_2068,N_3301);
and U4826 (N_4826,N_3069,N_2133);
and U4827 (N_4827,N_3919,N_3338);
nand U4828 (N_4828,N_3015,N_3016);
nand U4829 (N_4829,N_3459,N_3335);
nand U4830 (N_4830,N_2245,N_3929);
and U4831 (N_4831,N_2568,N_3818);
and U4832 (N_4832,N_2627,N_2646);
and U4833 (N_4833,N_2575,N_3529);
or U4834 (N_4834,N_3321,N_3881);
nor U4835 (N_4835,N_3342,N_3181);
and U4836 (N_4836,N_2159,N_3948);
nor U4837 (N_4837,N_2104,N_2754);
nor U4838 (N_4838,N_2210,N_2722);
or U4839 (N_4839,N_3939,N_2371);
nor U4840 (N_4840,N_3184,N_2702);
nand U4841 (N_4841,N_3116,N_2329);
nand U4842 (N_4842,N_3475,N_3546);
or U4843 (N_4843,N_2541,N_3554);
nand U4844 (N_4844,N_2250,N_3532);
xnor U4845 (N_4845,N_2430,N_2177);
nand U4846 (N_4846,N_3568,N_3849);
nand U4847 (N_4847,N_3118,N_3762);
nor U4848 (N_4848,N_3061,N_2556);
nor U4849 (N_4849,N_2090,N_2184);
nor U4850 (N_4850,N_2708,N_2300);
or U4851 (N_4851,N_3264,N_3834);
and U4852 (N_4852,N_2515,N_3933);
nor U4853 (N_4853,N_2574,N_2010);
nand U4854 (N_4854,N_3298,N_3656);
nor U4855 (N_4855,N_3356,N_3499);
or U4856 (N_4856,N_2425,N_2648);
and U4857 (N_4857,N_3108,N_2584);
and U4858 (N_4858,N_3375,N_3531);
and U4859 (N_4859,N_2306,N_2457);
and U4860 (N_4860,N_2981,N_2952);
or U4861 (N_4861,N_3572,N_3921);
and U4862 (N_4862,N_3038,N_2257);
xnor U4863 (N_4863,N_2048,N_2856);
nand U4864 (N_4864,N_3900,N_3786);
and U4865 (N_4865,N_2533,N_3961);
nand U4866 (N_4866,N_3704,N_2947);
or U4867 (N_4867,N_2494,N_2656);
and U4868 (N_4868,N_2848,N_2316);
nand U4869 (N_4869,N_2409,N_3576);
nor U4870 (N_4870,N_2265,N_2404);
and U4871 (N_4871,N_2311,N_2059);
nor U4872 (N_4872,N_3659,N_3250);
or U4873 (N_4873,N_3868,N_3304);
xnor U4874 (N_4874,N_2896,N_2216);
nor U4875 (N_4875,N_2367,N_2462);
nand U4876 (N_4876,N_2071,N_2096);
and U4877 (N_4877,N_3205,N_3453);
and U4878 (N_4878,N_3584,N_2190);
and U4879 (N_4879,N_2528,N_2594);
nand U4880 (N_4880,N_2105,N_3820);
xor U4881 (N_4881,N_3125,N_3556);
nor U4882 (N_4882,N_3837,N_3239);
and U4883 (N_4883,N_3105,N_3273);
nor U4884 (N_4884,N_3180,N_2004);
or U4885 (N_4885,N_2039,N_2200);
and U4886 (N_4886,N_2135,N_2395);
nand U4887 (N_4887,N_3569,N_3779);
nand U4888 (N_4888,N_2692,N_3461);
nand U4889 (N_4889,N_2141,N_2807);
or U4890 (N_4890,N_3530,N_2548);
or U4891 (N_4891,N_2428,N_3017);
nand U4892 (N_4892,N_3899,N_3671);
nand U4893 (N_4893,N_3767,N_3810);
nand U4894 (N_4894,N_2579,N_3533);
or U4895 (N_4895,N_3350,N_3733);
nor U4896 (N_4896,N_2679,N_2532);
or U4897 (N_4897,N_2310,N_3064);
nand U4898 (N_4898,N_2283,N_3202);
and U4899 (N_4899,N_2644,N_3693);
and U4900 (N_4900,N_2639,N_3872);
or U4901 (N_4901,N_2324,N_3696);
or U4902 (N_4902,N_3754,N_2966);
and U4903 (N_4903,N_2326,N_2349);
nand U4904 (N_4904,N_2783,N_3037);
and U4905 (N_4905,N_2078,N_3337);
and U4906 (N_4906,N_3456,N_2403);
or U4907 (N_4907,N_3686,N_2965);
nor U4908 (N_4908,N_3478,N_2103);
and U4909 (N_4909,N_2222,N_3500);
nor U4910 (N_4910,N_2930,N_2008);
and U4911 (N_4911,N_3167,N_3419);
nor U4912 (N_4912,N_2954,N_3766);
xnor U4913 (N_4913,N_2153,N_2889);
xor U4914 (N_4914,N_3373,N_2868);
nor U4915 (N_4915,N_3920,N_3266);
or U4916 (N_4916,N_2811,N_2249);
nand U4917 (N_4917,N_2546,N_3769);
and U4918 (N_4918,N_3143,N_2561);
and U4919 (N_4919,N_3819,N_3743);
nor U4920 (N_4920,N_3137,N_2520);
nor U4921 (N_4921,N_2195,N_3039);
xnor U4922 (N_4922,N_2577,N_3283);
and U4923 (N_4923,N_3494,N_3089);
or U4924 (N_4924,N_2926,N_3950);
and U4925 (N_4925,N_3282,N_2565);
and U4926 (N_4926,N_2235,N_3598);
xnor U4927 (N_4927,N_3010,N_2501);
or U4928 (N_4928,N_2477,N_2173);
and U4929 (N_4929,N_3195,N_2236);
and U4930 (N_4930,N_2127,N_2212);
and U4931 (N_4931,N_2619,N_2985);
and U4932 (N_4932,N_3208,N_2118);
or U4933 (N_4933,N_3668,N_3737);
or U4934 (N_4934,N_3207,N_3746);
or U4935 (N_4935,N_3138,N_2962);
nand U4936 (N_4936,N_3040,N_3006);
xor U4937 (N_4937,N_3472,N_3901);
and U4938 (N_4938,N_3926,N_2420);
and U4939 (N_4939,N_2134,N_2610);
nor U4940 (N_4940,N_3399,N_3937);
and U4941 (N_4941,N_3838,N_2315);
nand U4942 (N_4942,N_2156,N_2438);
nor U4943 (N_4943,N_3605,N_3727);
or U4944 (N_4944,N_2877,N_2790);
nand U4945 (N_4945,N_2831,N_2902);
nand U4946 (N_4946,N_2138,N_3910);
and U4947 (N_4947,N_3777,N_2046);
nand U4948 (N_4948,N_2136,N_3812);
or U4949 (N_4949,N_2534,N_2429);
xor U4950 (N_4950,N_2784,N_3518);
xnor U4951 (N_4951,N_2013,N_2567);
nand U4952 (N_4952,N_2360,N_3262);
or U4953 (N_4953,N_2106,N_3204);
and U4954 (N_4954,N_2253,N_3889);
nor U4955 (N_4955,N_2598,N_2622);
nand U4956 (N_4956,N_2382,N_2453);
nand U4957 (N_4957,N_2029,N_2493);
xnor U4958 (N_4958,N_3925,N_2707);
nor U4959 (N_4959,N_3126,N_3823);
or U4960 (N_4960,N_2381,N_2358);
or U4961 (N_4961,N_3261,N_2219);
and U4962 (N_4962,N_2023,N_3515);
nand U4963 (N_4963,N_3055,N_2119);
or U4964 (N_4964,N_3408,N_2055);
nand U4965 (N_4965,N_2228,N_2549);
or U4966 (N_4966,N_3721,N_3344);
nor U4967 (N_4967,N_2335,N_2002);
or U4968 (N_4968,N_3245,N_2695);
nor U4969 (N_4969,N_2525,N_2144);
nand U4970 (N_4970,N_2912,N_2795);
and U4971 (N_4971,N_3255,N_3795);
nand U4972 (N_4972,N_2512,N_2321);
nor U4973 (N_4973,N_3495,N_3987);
xnor U4974 (N_4974,N_3259,N_2812);
nor U4975 (N_4975,N_2569,N_2142);
and U4976 (N_4976,N_3492,N_2663);
nand U4977 (N_4977,N_2149,N_2332);
or U4978 (N_4978,N_2510,N_2921);
nand U4979 (N_4979,N_2578,N_3884);
xor U4980 (N_4980,N_3340,N_2847);
nor U4981 (N_4981,N_2502,N_3141);
and U4982 (N_4982,N_2188,N_3867);
and U4983 (N_4983,N_2206,N_3134);
and U4984 (N_4984,N_3517,N_2272);
xnor U4985 (N_4985,N_2365,N_3840);
nor U4986 (N_4986,N_2904,N_3856);
nand U4987 (N_4987,N_2346,N_3312);
nor U4988 (N_4988,N_3740,N_3800);
nand U4989 (N_4989,N_2476,N_2826);
nor U4990 (N_4990,N_3110,N_3288);
nand U4991 (N_4991,N_2674,N_2616);
nor U4992 (N_4992,N_2484,N_3140);
and U4993 (N_4993,N_2389,N_3982);
nand U4994 (N_4994,N_3319,N_3669);
and U4995 (N_4995,N_2017,N_2894);
nor U4996 (N_4996,N_2165,N_2126);
nand U4997 (N_4997,N_2983,N_2670);
nor U4998 (N_4998,N_3816,N_3644);
nor U4999 (N_4999,N_2516,N_3409);
nand U5000 (N_5000,N_3646,N_3247);
nor U5001 (N_5001,N_2143,N_2553);
nand U5002 (N_5002,N_3829,N_3670);
and U5003 (N_5003,N_2735,N_2305);
nand U5004 (N_5004,N_2391,N_3478);
nand U5005 (N_5005,N_2242,N_2877);
nor U5006 (N_5006,N_3589,N_3952);
xor U5007 (N_5007,N_3439,N_3591);
nand U5008 (N_5008,N_2448,N_2332);
nand U5009 (N_5009,N_2027,N_3052);
and U5010 (N_5010,N_3388,N_3933);
nor U5011 (N_5011,N_3412,N_2344);
nand U5012 (N_5012,N_3368,N_2191);
nand U5013 (N_5013,N_2011,N_3118);
nor U5014 (N_5014,N_2016,N_3633);
nand U5015 (N_5015,N_2529,N_2242);
and U5016 (N_5016,N_3996,N_2447);
nand U5017 (N_5017,N_2088,N_3812);
and U5018 (N_5018,N_3472,N_3260);
nor U5019 (N_5019,N_2333,N_3444);
nor U5020 (N_5020,N_2748,N_3954);
nor U5021 (N_5021,N_2023,N_2611);
and U5022 (N_5022,N_2943,N_2130);
nor U5023 (N_5023,N_3036,N_2153);
xnor U5024 (N_5024,N_2759,N_3323);
or U5025 (N_5025,N_2977,N_2526);
nor U5026 (N_5026,N_2210,N_2211);
and U5027 (N_5027,N_2822,N_2096);
or U5028 (N_5028,N_3971,N_3203);
and U5029 (N_5029,N_3362,N_3063);
nor U5030 (N_5030,N_3466,N_3688);
nor U5031 (N_5031,N_2196,N_3702);
or U5032 (N_5032,N_2971,N_3753);
and U5033 (N_5033,N_2694,N_2735);
and U5034 (N_5034,N_3060,N_3840);
nand U5035 (N_5035,N_2019,N_2721);
nand U5036 (N_5036,N_3340,N_2494);
and U5037 (N_5037,N_2927,N_2682);
nand U5038 (N_5038,N_3717,N_3023);
or U5039 (N_5039,N_3384,N_2211);
and U5040 (N_5040,N_2153,N_2789);
or U5041 (N_5041,N_3146,N_3092);
and U5042 (N_5042,N_3552,N_3348);
and U5043 (N_5043,N_3444,N_2733);
nor U5044 (N_5044,N_3152,N_2868);
and U5045 (N_5045,N_2691,N_3676);
or U5046 (N_5046,N_3992,N_3597);
and U5047 (N_5047,N_3830,N_3491);
nand U5048 (N_5048,N_3659,N_3928);
nand U5049 (N_5049,N_2698,N_2192);
nor U5050 (N_5050,N_3067,N_3930);
xor U5051 (N_5051,N_3923,N_3081);
or U5052 (N_5052,N_2702,N_3434);
nand U5053 (N_5053,N_2983,N_3783);
nor U5054 (N_5054,N_2414,N_3840);
nor U5055 (N_5055,N_3342,N_2888);
or U5056 (N_5056,N_3964,N_2699);
nor U5057 (N_5057,N_2360,N_2163);
xor U5058 (N_5058,N_2533,N_2021);
nor U5059 (N_5059,N_2965,N_2731);
or U5060 (N_5060,N_2682,N_3130);
or U5061 (N_5061,N_3245,N_2241);
nor U5062 (N_5062,N_2921,N_3893);
nor U5063 (N_5063,N_2195,N_2358);
and U5064 (N_5064,N_3423,N_2368);
or U5065 (N_5065,N_2923,N_3787);
nor U5066 (N_5066,N_2427,N_3169);
nand U5067 (N_5067,N_2355,N_3956);
nand U5068 (N_5068,N_2223,N_3052);
nand U5069 (N_5069,N_2566,N_3230);
and U5070 (N_5070,N_3365,N_2062);
or U5071 (N_5071,N_2180,N_2349);
xor U5072 (N_5072,N_2687,N_2808);
or U5073 (N_5073,N_2560,N_3936);
or U5074 (N_5074,N_3174,N_2894);
nor U5075 (N_5075,N_3379,N_3251);
and U5076 (N_5076,N_3419,N_2586);
and U5077 (N_5077,N_3579,N_3661);
or U5078 (N_5078,N_2553,N_2230);
and U5079 (N_5079,N_3530,N_3305);
xnor U5080 (N_5080,N_3402,N_3130);
or U5081 (N_5081,N_2071,N_2120);
and U5082 (N_5082,N_2575,N_2716);
nor U5083 (N_5083,N_2866,N_3482);
and U5084 (N_5084,N_2851,N_2333);
or U5085 (N_5085,N_3138,N_2746);
nand U5086 (N_5086,N_2037,N_2631);
or U5087 (N_5087,N_2115,N_2099);
xor U5088 (N_5088,N_2806,N_3262);
xor U5089 (N_5089,N_2489,N_3810);
nand U5090 (N_5090,N_3873,N_2744);
nand U5091 (N_5091,N_2161,N_2375);
xnor U5092 (N_5092,N_3235,N_3044);
xnor U5093 (N_5093,N_2038,N_2515);
nor U5094 (N_5094,N_2334,N_2732);
nor U5095 (N_5095,N_2169,N_3526);
nand U5096 (N_5096,N_3393,N_2440);
or U5097 (N_5097,N_3895,N_2260);
nor U5098 (N_5098,N_3472,N_3481);
xnor U5099 (N_5099,N_2862,N_3362);
and U5100 (N_5100,N_2611,N_2348);
and U5101 (N_5101,N_2102,N_3874);
or U5102 (N_5102,N_3887,N_2432);
or U5103 (N_5103,N_3589,N_3548);
nand U5104 (N_5104,N_2795,N_3775);
xor U5105 (N_5105,N_3123,N_3124);
nand U5106 (N_5106,N_3223,N_2525);
and U5107 (N_5107,N_2337,N_3143);
or U5108 (N_5108,N_3892,N_2955);
or U5109 (N_5109,N_2716,N_3753);
or U5110 (N_5110,N_3157,N_3925);
and U5111 (N_5111,N_3227,N_2361);
nand U5112 (N_5112,N_2787,N_3046);
and U5113 (N_5113,N_3407,N_2310);
or U5114 (N_5114,N_2195,N_3662);
nand U5115 (N_5115,N_3410,N_3250);
nand U5116 (N_5116,N_3813,N_3842);
nand U5117 (N_5117,N_2861,N_3334);
or U5118 (N_5118,N_2148,N_3613);
nand U5119 (N_5119,N_2598,N_2710);
or U5120 (N_5120,N_3685,N_3211);
nor U5121 (N_5121,N_3942,N_3717);
and U5122 (N_5122,N_3647,N_3315);
nor U5123 (N_5123,N_3795,N_3352);
or U5124 (N_5124,N_3707,N_2346);
nor U5125 (N_5125,N_3786,N_3488);
nor U5126 (N_5126,N_2388,N_2770);
and U5127 (N_5127,N_2266,N_2949);
nor U5128 (N_5128,N_2103,N_2448);
nand U5129 (N_5129,N_3220,N_3517);
or U5130 (N_5130,N_2607,N_3343);
or U5131 (N_5131,N_3262,N_3169);
xor U5132 (N_5132,N_2699,N_3925);
nor U5133 (N_5133,N_2673,N_3724);
xor U5134 (N_5134,N_2394,N_2143);
or U5135 (N_5135,N_2757,N_2386);
nor U5136 (N_5136,N_2095,N_2776);
or U5137 (N_5137,N_3412,N_2976);
or U5138 (N_5138,N_3977,N_3120);
or U5139 (N_5139,N_3841,N_3699);
nor U5140 (N_5140,N_2428,N_3825);
nand U5141 (N_5141,N_3761,N_3328);
nor U5142 (N_5142,N_2646,N_2490);
xor U5143 (N_5143,N_3663,N_2984);
or U5144 (N_5144,N_3097,N_2832);
or U5145 (N_5145,N_2096,N_3322);
xor U5146 (N_5146,N_3331,N_2583);
or U5147 (N_5147,N_3218,N_3053);
nand U5148 (N_5148,N_2820,N_3566);
and U5149 (N_5149,N_2667,N_2203);
or U5150 (N_5150,N_3461,N_3200);
and U5151 (N_5151,N_2803,N_2216);
or U5152 (N_5152,N_2824,N_3769);
nor U5153 (N_5153,N_3269,N_2778);
nand U5154 (N_5154,N_2186,N_2605);
nor U5155 (N_5155,N_2714,N_3476);
nor U5156 (N_5156,N_2619,N_3998);
nand U5157 (N_5157,N_3037,N_2003);
nand U5158 (N_5158,N_3175,N_2483);
and U5159 (N_5159,N_2786,N_3212);
and U5160 (N_5160,N_3949,N_2280);
and U5161 (N_5161,N_3015,N_3584);
and U5162 (N_5162,N_3968,N_2528);
or U5163 (N_5163,N_2210,N_2122);
xnor U5164 (N_5164,N_2990,N_3074);
nand U5165 (N_5165,N_2572,N_3643);
and U5166 (N_5166,N_3256,N_2250);
or U5167 (N_5167,N_2358,N_2953);
or U5168 (N_5168,N_2315,N_3846);
or U5169 (N_5169,N_2577,N_3042);
or U5170 (N_5170,N_3010,N_3125);
nand U5171 (N_5171,N_2888,N_3888);
or U5172 (N_5172,N_3385,N_2565);
and U5173 (N_5173,N_3036,N_2849);
nand U5174 (N_5174,N_3357,N_3384);
or U5175 (N_5175,N_3614,N_3076);
and U5176 (N_5176,N_3230,N_2390);
or U5177 (N_5177,N_2570,N_2166);
or U5178 (N_5178,N_3179,N_3701);
nand U5179 (N_5179,N_2375,N_3988);
or U5180 (N_5180,N_2755,N_2737);
or U5181 (N_5181,N_2911,N_2922);
or U5182 (N_5182,N_2118,N_2693);
nand U5183 (N_5183,N_3285,N_2188);
nor U5184 (N_5184,N_2900,N_3403);
and U5185 (N_5185,N_2571,N_2518);
and U5186 (N_5186,N_2122,N_3746);
xnor U5187 (N_5187,N_3785,N_2914);
xor U5188 (N_5188,N_2630,N_2221);
nand U5189 (N_5189,N_2785,N_2568);
and U5190 (N_5190,N_3964,N_2147);
or U5191 (N_5191,N_2031,N_3864);
nor U5192 (N_5192,N_3356,N_3892);
xor U5193 (N_5193,N_3163,N_2715);
or U5194 (N_5194,N_2864,N_3000);
nor U5195 (N_5195,N_2690,N_3497);
nand U5196 (N_5196,N_2107,N_2795);
nand U5197 (N_5197,N_3551,N_3650);
nor U5198 (N_5198,N_2465,N_2179);
nand U5199 (N_5199,N_3388,N_3459);
nand U5200 (N_5200,N_2035,N_2418);
or U5201 (N_5201,N_3347,N_2224);
or U5202 (N_5202,N_3582,N_3469);
or U5203 (N_5203,N_2519,N_3246);
and U5204 (N_5204,N_3178,N_2977);
nor U5205 (N_5205,N_2535,N_3430);
nand U5206 (N_5206,N_2850,N_2507);
nand U5207 (N_5207,N_3763,N_2465);
nand U5208 (N_5208,N_2712,N_3784);
and U5209 (N_5209,N_2078,N_3226);
or U5210 (N_5210,N_3075,N_2780);
and U5211 (N_5211,N_3209,N_2911);
nor U5212 (N_5212,N_2996,N_3511);
nand U5213 (N_5213,N_2652,N_2895);
or U5214 (N_5214,N_3875,N_2315);
or U5215 (N_5215,N_2920,N_3538);
and U5216 (N_5216,N_2663,N_3752);
nand U5217 (N_5217,N_2800,N_2266);
nor U5218 (N_5218,N_3647,N_2787);
or U5219 (N_5219,N_3567,N_2746);
xor U5220 (N_5220,N_3891,N_2766);
or U5221 (N_5221,N_2671,N_3733);
nand U5222 (N_5222,N_2826,N_3306);
nor U5223 (N_5223,N_3497,N_3743);
xnor U5224 (N_5224,N_3093,N_2028);
nand U5225 (N_5225,N_2355,N_2333);
nor U5226 (N_5226,N_2761,N_2160);
or U5227 (N_5227,N_3568,N_3064);
and U5228 (N_5228,N_3154,N_3546);
and U5229 (N_5229,N_2143,N_3491);
nand U5230 (N_5230,N_2056,N_3970);
nor U5231 (N_5231,N_2827,N_3513);
or U5232 (N_5232,N_3199,N_2038);
nor U5233 (N_5233,N_3449,N_3169);
nand U5234 (N_5234,N_2496,N_3418);
nand U5235 (N_5235,N_2014,N_3812);
and U5236 (N_5236,N_3228,N_2625);
or U5237 (N_5237,N_3918,N_2041);
nor U5238 (N_5238,N_2193,N_2226);
nor U5239 (N_5239,N_3542,N_3896);
nor U5240 (N_5240,N_3108,N_3983);
nor U5241 (N_5241,N_2888,N_3887);
or U5242 (N_5242,N_3525,N_3051);
or U5243 (N_5243,N_3955,N_3413);
and U5244 (N_5244,N_3586,N_3739);
or U5245 (N_5245,N_3408,N_3572);
nor U5246 (N_5246,N_2710,N_2750);
xnor U5247 (N_5247,N_3232,N_2576);
and U5248 (N_5248,N_2203,N_3690);
and U5249 (N_5249,N_2334,N_2966);
nor U5250 (N_5250,N_3390,N_3784);
nor U5251 (N_5251,N_2879,N_2077);
and U5252 (N_5252,N_2722,N_2730);
nand U5253 (N_5253,N_3386,N_3791);
nor U5254 (N_5254,N_2069,N_3713);
nand U5255 (N_5255,N_3401,N_3812);
and U5256 (N_5256,N_2293,N_3602);
nor U5257 (N_5257,N_2418,N_2320);
or U5258 (N_5258,N_2410,N_3757);
nand U5259 (N_5259,N_3791,N_3422);
and U5260 (N_5260,N_2802,N_3712);
or U5261 (N_5261,N_2636,N_3259);
nand U5262 (N_5262,N_2801,N_2409);
nand U5263 (N_5263,N_2530,N_2082);
nand U5264 (N_5264,N_2512,N_2848);
nand U5265 (N_5265,N_2833,N_2131);
nor U5266 (N_5266,N_2777,N_3162);
nand U5267 (N_5267,N_3743,N_2288);
or U5268 (N_5268,N_2218,N_3141);
nor U5269 (N_5269,N_2902,N_3957);
and U5270 (N_5270,N_2752,N_3145);
and U5271 (N_5271,N_2012,N_2615);
nand U5272 (N_5272,N_3579,N_3670);
and U5273 (N_5273,N_3444,N_2409);
nand U5274 (N_5274,N_2377,N_3342);
and U5275 (N_5275,N_3923,N_2765);
nand U5276 (N_5276,N_2719,N_3172);
nand U5277 (N_5277,N_2175,N_2665);
nand U5278 (N_5278,N_2791,N_2172);
nand U5279 (N_5279,N_2226,N_3958);
nor U5280 (N_5280,N_2378,N_2312);
nand U5281 (N_5281,N_3133,N_3271);
or U5282 (N_5282,N_2869,N_3997);
nor U5283 (N_5283,N_2729,N_2938);
or U5284 (N_5284,N_2508,N_2791);
nand U5285 (N_5285,N_3640,N_3176);
or U5286 (N_5286,N_3081,N_2238);
and U5287 (N_5287,N_3822,N_2794);
nor U5288 (N_5288,N_3492,N_2224);
nor U5289 (N_5289,N_3505,N_2852);
or U5290 (N_5290,N_3040,N_2159);
nand U5291 (N_5291,N_2187,N_3781);
nand U5292 (N_5292,N_2468,N_2114);
nor U5293 (N_5293,N_2341,N_3052);
nand U5294 (N_5294,N_3929,N_2734);
and U5295 (N_5295,N_3080,N_3879);
or U5296 (N_5296,N_3431,N_2265);
nand U5297 (N_5297,N_2050,N_3232);
nand U5298 (N_5298,N_2188,N_3433);
or U5299 (N_5299,N_2290,N_2212);
and U5300 (N_5300,N_2844,N_2722);
nand U5301 (N_5301,N_2946,N_3174);
nand U5302 (N_5302,N_3969,N_2514);
nand U5303 (N_5303,N_3685,N_2400);
or U5304 (N_5304,N_3918,N_3861);
and U5305 (N_5305,N_2111,N_2898);
or U5306 (N_5306,N_2365,N_3029);
nor U5307 (N_5307,N_3061,N_3967);
nor U5308 (N_5308,N_3800,N_2214);
nor U5309 (N_5309,N_2087,N_3330);
nand U5310 (N_5310,N_2791,N_2161);
and U5311 (N_5311,N_2095,N_3043);
and U5312 (N_5312,N_2472,N_2147);
or U5313 (N_5313,N_2780,N_2451);
and U5314 (N_5314,N_2671,N_3751);
or U5315 (N_5315,N_2369,N_2928);
and U5316 (N_5316,N_3251,N_3470);
and U5317 (N_5317,N_2332,N_2682);
nand U5318 (N_5318,N_3217,N_3700);
nor U5319 (N_5319,N_3795,N_2255);
nor U5320 (N_5320,N_2988,N_2087);
nand U5321 (N_5321,N_2062,N_2050);
or U5322 (N_5322,N_3283,N_3017);
or U5323 (N_5323,N_3519,N_3896);
or U5324 (N_5324,N_2473,N_3183);
nand U5325 (N_5325,N_2395,N_3255);
nand U5326 (N_5326,N_2752,N_2387);
nor U5327 (N_5327,N_2796,N_3899);
and U5328 (N_5328,N_2927,N_2000);
and U5329 (N_5329,N_3845,N_2188);
nand U5330 (N_5330,N_2836,N_3663);
nor U5331 (N_5331,N_3893,N_2841);
or U5332 (N_5332,N_3652,N_2757);
and U5333 (N_5333,N_3477,N_2685);
xnor U5334 (N_5334,N_2254,N_2573);
nor U5335 (N_5335,N_3468,N_2159);
or U5336 (N_5336,N_2127,N_3679);
nand U5337 (N_5337,N_2330,N_2174);
nor U5338 (N_5338,N_3903,N_2438);
and U5339 (N_5339,N_3558,N_2277);
or U5340 (N_5340,N_2794,N_2964);
nor U5341 (N_5341,N_3033,N_2312);
and U5342 (N_5342,N_2395,N_2321);
or U5343 (N_5343,N_2574,N_3752);
nand U5344 (N_5344,N_2690,N_2895);
nand U5345 (N_5345,N_2616,N_3425);
or U5346 (N_5346,N_2608,N_2613);
nor U5347 (N_5347,N_2895,N_2965);
nor U5348 (N_5348,N_3187,N_3499);
nand U5349 (N_5349,N_2589,N_3590);
and U5350 (N_5350,N_3183,N_2210);
nand U5351 (N_5351,N_3435,N_3758);
or U5352 (N_5352,N_2702,N_3951);
or U5353 (N_5353,N_2090,N_2215);
nand U5354 (N_5354,N_3234,N_3615);
xnor U5355 (N_5355,N_2415,N_2421);
or U5356 (N_5356,N_3119,N_3768);
nand U5357 (N_5357,N_2866,N_3827);
nand U5358 (N_5358,N_3260,N_3694);
nor U5359 (N_5359,N_2553,N_2192);
and U5360 (N_5360,N_3401,N_2111);
nor U5361 (N_5361,N_2925,N_2098);
and U5362 (N_5362,N_3826,N_2236);
or U5363 (N_5363,N_2059,N_3479);
nor U5364 (N_5364,N_3799,N_3754);
or U5365 (N_5365,N_3436,N_2568);
nor U5366 (N_5366,N_3029,N_3913);
nand U5367 (N_5367,N_2108,N_2675);
nor U5368 (N_5368,N_3206,N_3800);
nand U5369 (N_5369,N_3100,N_3187);
nand U5370 (N_5370,N_2638,N_3745);
and U5371 (N_5371,N_3873,N_2292);
and U5372 (N_5372,N_3581,N_3313);
or U5373 (N_5373,N_2393,N_2240);
or U5374 (N_5374,N_2244,N_3617);
nand U5375 (N_5375,N_2622,N_2633);
nor U5376 (N_5376,N_2830,N_3988);
nor U5377 (N_5377,N_2919,N_3272);
nand U5378 (N_5378,N_2515,N_3571);
or U5379 (N_5379,N_2672,N_3756);
and U5380 (N_5380,N_3684,N_2666);
nand U5381 (N_5381,N_3273,N_2104);
nand U5382 (N_5382,N_2660,N_2246);
nand U5383 (N_5383,N_3553,N_3475);
nand U5384 (N_5384,N_2272,N_2912);
nand U5385 (N_5385,N_3943,N_2851);
nor U5386 (N_5386,N_2012,N_2164);
nand U5387 (N_5387,N_2949,N_3737);
nor U5388 (N_5388,N_3473,N_3450);
nor U5389 (N_5389,N_2125,N_3293);
and U5390 (N_5390,N_3561,N_2345);
xnor U5391 (N_5391,N_3728,N_2283);
nand U5392 (N_5392,N_3135,N_2603);
nor U5393 (N_5393,N_2225,N_2075);
nand U5394 (N_5394,N_3529,N_3605);
nand U5395 (N_5395,N_2517,N_3068);
or U5396 (N_5396,N_2385,N_3751);
nor U5397 (N_5397,N_3367,N_2128);
or U5398 (N_5398,N_2452,N_2828);
and U5399 (N_5399,N_3577,N_3069);
nor U5400 (N_5400,N_2027,N_3700);
nand U5401 (N_5401,N_2989,N_2888);
and U5402 (N_5402,N_2616,N_3639);
nand U5403 (N_5403,N_3266,N_2000);
nand U5404 (N_5404,N_3581,N_2832);
nor U5405 (N_5405,N_3826,N_3868);
nand U5406 (N_5406,N_3954,N_2760);
and U5407 (N_5407,N_3596,N_2976);
nor U5408 (N_5408,N_3055,N_2279);
nor U5409 (N_5409,N_2543,N_2288);
xor U5410 (N_5410,N_2589,N_3658);
and U5411 (N_5411,N_3185,N_3566);
nor U5412 (N_5412,N_3679,N_2292);
nor U5413 (N_5413,N_2184,N_2557);
nor U5414 (N_5414,N_2710,N_3296);
and U5415 (N_5415,N_2091,N_3127);
or U5416 (N_5416,N_3681,N_2994);
and U5417 (N_5417,N_2039,N_2762);
or U5418 (N_5418,N_2994,N_3585);
or U5419 (N_5419,N_3175,N_3255);
nand U5420 (N_5420,N_2005,N_3294);
nor U5421 (N_5421,N_2958,N_2138);
and U5422 (N_5422,N_3860,N_3200);
and U5423 (N_5423,N_3376,N_2994);
nor U5424 (N_5424,N_2590,N_3654);
nor U5425 (N_5425,N_3327,N_2123);
nand U5426 (N_5426,N_2579,N_3264);
and U5427 (N_5427,N_2465,N_3826);
nor U5428 (N_5428,N_3015,N_2912);
nor U5429 (N_5429,N_3513,N_2487);
or U5430 (N_5430,N_3085,N_2246);
nand U5431 (N_5431,N_2475,N_2064);
and U5432 (N_5432,N_2958,N_3120);
nand U5433 (N_5433,N_2480,N_3508);
nor U5434 (N_5434,N_2389,N_2782);
or U5435 (N_5435,N_3317,N_3337);
and U5436 (N_5436,N_2582,N_3238);
and U5437 (N_5437,N_2999,N_2797);
nand U5438 (N_5438,N_2706,N_3155);
nor U5439 (N_5439,N_3617,N_2434);
or U5440 (N_5440,N_3507,N_2625);
nor U5441 (N_5441,N_3666,N_3499);
or U5442 (N_5442,N_3189,N_3005);
nand U5443 (N_5443,N_3848,N_3045);
and U5444 (N_5444,N_2840,N_3699);
nor U5445 (N_5445,N_2299,N_2091);
or U5446 (N_5446,N_3168,N_2661);
and U5447 (N_5447,N_2407,N_2161);
or U5448 (N_5448,N_2058,N_2471);
nor U5449 (N_5449,N_2224,N_3416);
or U5450 (N_5450,N_3776,N_3832);
nand U5451 (N_5451,N_3612,N_2903);
or U5452 (N_5452,N_2717,N_2914);
nand U5453 (N_5453,N_3325,N_3524);
nor U5454 (N_5454,N_2925,N_2832);
and U5455 (N_5455,N_2568,N_2266);
nand U5456 (N_5456,N_3819,N_3301);
or U5457 (N_5457,N_3938,N_2582);
xnor U5458 (N_5458,N_2699,N_2421);
or U5459 (N_5459,N_2166,N_3413);
and U5460 (N_5460,N_3297,N_2062);
nand U5461 (N_5461,N_2238,N_3141);
or U5462 (N_5462,N_2106,N_2818);
nor U5463 (N_5463,N_2476,N_2624);
or U5464 (N_5464,N_3642,N_3907);
or U5465 (N_5465,N_3226,N_2971);
nand U5466 (N_5466,N_3165,N_2752);
or U5467 (N_5467,N_2372,N_2614);
xor U5468 (N_5468,N_2535,N_2387);
and U5469 (N_5469,N_3551,N_3972);
and U5470 (N_5470,N_3632,N_2938);
and U5471 (N_5471,N_2387,N_3860);
and U5472 (N_5472,N_3948,N_3098);
and U5473 (N_5473,N_3503,N_3083);
nand U5474 (N_5474,N_2762,N_3447);
nor U5475 (N_5475,N_2558,N_3636);
nor U5476 (N_5476,N_2104,N_2290);
and U5477 (N_5477,N_3247,N_2152);
or U5478 (N_5478,N_3802,N_3903);
nand U5479 (N_5479,N_2717,N_2405);
and U5480 (N_5480,N_3285,N_3029);
and U5481 (N_5481,N_2780,N_3668);
nor U5482 (N_5482,N_2357,N_2871);
nand U5483 (N_5483,N_3205,N_3904);
and U5484 (N_5484,N_3391,N_3056);
nand U5485 (N_5485,N_2448,N_2218);
and U5486 (N_5486,N_3808,N_2964);
nand U5487 (N_5487,N_2249,N_2111);
nor U5488 (N_5488,N_2348,N_2716);
nor U5489 (N_5489,N_2945,N_2121);
nor U5490 (N_5490,N_2561,N_2363);
and U5491 (N_5491,N_3128,N_3641);
nand U5492 (N_5492,N_3882,N_2500);
and U5493 (N_5493,N_3328,N_2091);
and U5494 (N_5494,N_3532,N_3651);
or U5495 (N_5495,N_3925,N_2519);
and U5496 (N_5496,N_3105,N_2837);
nand U5497 (N_5497,N_3255,N_3596);
nand U5498 (N_5498,N_2386,N_3144);
nor U5499 (N_5499,N_2240,N_3760);
and U5500 (N_5500,N_2172,N_2860);
nor U5501 (N_5501,N_2837,N_3868);
and U5502 (N_5502,N_3679,N_3700);
nor U5503 (N_5503,N_3567,N_2589);
nor U5504 (N_5504,N_2088,N_3807);
or U5505 (N_5505,N_2605,N_2736);
nand U5506 (N_5506,N_2867,N_3905);
nand U5507 (N_5507,N_2388,N_2263);
or U5508 (N_5508,N_2451,N_2343);
and U5509 (N_5509,N_3363,N_2530);
nand U5510 (N_5510,N_3384,N_3854);
nor U5511 (N_5511,N_2568,N_2451);
nor U5512 (N_5512,N_2805,N_2125);
and U5513 (N_5513,N_2306,N_2550);
or U5514 (N_5514,N_3224,N_2253);
nor U5515 (N_5515,N_3719,N_3751);
or U5516 (N_5516,N_3377,N_3306);
or U5517 (N_5517,N_3159,N_3876);
nand U5518 (N_5518,N_3204,N_2588);
nor U5519 (N_5519,N_2791,N_3801);
nand U5520 (N_5520,N_2470,N_2117);
nand U5521 (N_5521,N_2491,N_2534);
nand U5522 (N_5522,N_2548,N_2911);
nand U5523 (N_5523,N_3137,N_2875);
nor U5524 (N_5524,N_2220,N_2673);
or U5525 (N_5525,N_3584,N_2669);
nand U5526 (N_5526,N_3949,N_2187);
or U5527 (N_5527,N_3497,N_3705);
or U5528 (N_5528,N_3942,N_3457);
and U5529 (N_5529,N_2571,N_3820);
or U5530 (N_5530,N_3668,N_3568);
nand U5531 (N_5531,N_3115,N_2910);
nor U5532 (N_5532,N_3991,N_2897);
and U5533 (N_5533,N_2872,N_3371);
and U5534 (N_5534,N_2924,N_2019);
nor U5535 (N_5535,N_3362,N_3014);
nand U5536 (N_5536,N_2364,N_2071);
or U5537 (N_5537,N_3165,N_2431);
nor U5538 (N_5538,N_2075,N_3398);
nor U5539 (N_5539,N_3601,N_3389);
nor U5540 (N_5540,N_3119,N_2023);
nand U5541 (N_5541,N_3875,N_2443);
nor U5542 (N_5542,N_3501,N_2898);
nand U5543 (N_5543,N_2648,N_3972);
nor U5544 (N_5544,N_2794,N_3853);
or U5545 (N_5545,N_2646,N_3141);
nor U5546 (N_5546,N_3910,N_2107);
and U5547 (N_5547,N_3411,N_2815);
or U5548 (N_5548,N_3506,N_3486);
nand U5549 (N_5549,N_2103,N_2811);
or U5550 (N_5550,N_2907,N_2189);
nor U5551 (N_5551,N_2317,N_3675);
or U5552 (N_5552,N_3030,N_2911);
or U5553 (N_5553,N_2674,N_3503);
and U5554 (N_5554,N_3015,N_2044);
or U5555 (N_5555,N_3598,N_3413);
nor U5556 (N_5556,N_2053,N_2669);
nand U5557 (N_5557,N_3196,N_3108);
xor U5558 (N_5558,N_3808,N_2821);
nor U5559 (N_5559,N_2074,N_3877);
or U5560 (N_5560,N_3753,N_3121);
and U5561 (N_5561,N_3305,N_3836);
nand U5562 (N_5562,N_3663,N_2777);
or U5563 (N_5563,N_3544,N_2948);
nand U5564 (N_5564,N_3840,N_2976);
nor U5565 (N_5565,N_2101,N_3022);
nor U5566 (N_5566,N_3279,N_2023);
and U5567 (N_5567,N_3693,N_2475);
nand U5568 (N_5568,N_3754,N_3309);
nor U5569 (N_5569,N_3109,N_2958);
or U5570 (N_5570,N_3800,N_2907);
nand U5571 (N_5571,N_2609,N_3199);
and U5572 (N_5572,N_2420,N_2780);
and U5573 (N_5573,N_2776,N_3224);
or U5574 (N_5574,N_3600,N_3667);
and U5575 (N_5575,N_2829,N_2696);
nor U5576 (N_5576,N_2050,N_2211);
nor U5577 (N_5577,N_3292,N_2527);
xnor U5578 (N_5578,N_3731,N_2083);
nor U5579 (N_5579,N_2734,N_3123);
and U5580 (N_5580,N_3403,N_3531);
or U5581 (N_5581,N_3188,N_2872);
nand U5582 (N_5582,N_2261,N_3392);
nand U5583 (N_5583,N_2343,N_3491);
or U5584 (N_5584,N_2011,N_3854);
nand U5585 (N_5585,N_2800,N_3353);
nor U5586 (N_5586,N_3475,N_3059);
and U5587 (N_5587,N_3368,N_3579);
nor U5588 (N_5588,N_2105,N_2061);
and U5589 (N_5589,N_3606,N_3209);
nand U5590 (N_5590,N_2327,N_3250);
nand U5591 (N_5591,N_2552,N_2626);
or U5592 (N_5592,N_2740,N_2082);
nand U5593 (N_5593,N_2811,N_3675);
or U5594 (N_5594,N_3115,N_2348);
nand U5595 (N_5595,N_3378,N_3842);
nor U5596 (N_5596,N_3343,N_3920);
and U5597 (N_5597,N_2924,N_2242);
and U5598 (N_5598,N_3699,N_3145);
or U5599 (N_5599,N_3622,N_3022);
and U5600 (N_5600,N_3286,N_2805);
nand U5601 (N_5601,N_3464,N_2694);
and U5602 (N_5602,N_3253,N_2520);
or U5603 (N_5603,N_3954,N_2654);
or U5604 (N_5604,N_2690,N_2814);
nand U5605 (N_5605,N_3229,N_2130);
or U5606 (N_5606,N_3557,N_3702);
xor U5607 (N_5607,N_2382,N_3596);
or U5608 (N_5608,N_3280,N_2131);
or U5609 (N_5609,N_3016,N_3641);
nand U5610 (N_5610,N_3666,N_2724);
nand U5611 (N_5611,N_3255,N_3852);
nand U5612 (N_5612,N_2134,N_3425);
nor U5613 (N_5613,N_3822,N_2341);
nor U5614 (N_5614,N_3865,N_3546);
nor U5615 (N_5615,N_3143,N_2902);
nand U5616 (N_5616,N_3496,N_2782);
nor U5617 (N_5617,N_2922,N_3375);
or U5618 (N_5618,N_3107,N_3554);
and U5619 (N_5619,N_3278,N_2454);
and U5620 (N_5620,N_2748,N_2040);
or U5621 (N_5621,N_3656,N_3033);
nand U5622 (N_5622,N_2418,N_3594);
and U5623 (N_5623,N_2945,N_2333);
nor U5624 (N_5624,N_2653,N_3670);
or U5625 (N_5625,N_3499,N_2001);
nor U5626 (N_5626,N_3777,N_3692);
nor U5627 (N_5627,N_3083,N_3072);
nor U5628 (N_5628,N_2071,N_3310);
or U5629 (N_5629,N_3638,N_3500);
nor U5630 (N_5630,N_2128,N_2352);
or U5631 (N_5631,N_2658,N_3556);
nor U5632 (N_5632,N_2244,N_2830);
and U5633 (N_5633,N_3864,N_3605);
or U5634 (N_5634,N_3810,N_2479);
and U5635 (N_5635,N_3508,N_3945);
and U5636 (N_5636,N_3086,N_3438);
nor U5637 (N_5637,N_2513,N_2156);
nor U5638 (N_5638,N_3673,N_2715);
nor U5639 (N_5639,N_3274,N_3440);
nand U5640 (N_5640,N_3420,N_3060);
and U5641 (N_5641,N_3912,N_3703);
and U5642 (N_5642,N_3882,N_2393);
or U5643 (N_5643,N_2231,N_2804);
and U5644 (N_5644,N_3022,N_3112);
nand U5645 (N_5645,N_3014,N_3222);
nand U5646 (N_5646,N_3885,N_2988);
nor U5647 (N_5647,N_3693,N_2159);
or U5648 (N_5648,N_3808,N_3451);
and U5649 (N_5649,N_3318,N_3577);
or U5650 (N_5650,N_3416,N_2722);
or U5651 (N_5651,N_3206,N_2714);
or U5652 (N_5652,N_2515,N_2681);
and U5653 (N_5653,N_2915,N_3690);
and U5654 (N_5654,N_3242,N_2795);
or U5655 (N_5655,N_3960,N_2598);
or U5656 (N_5656,N_3875,N_2611);
and U5657 (N_5657,N_3183,N_3074);
and U5658 (N_5658,N_2429,N_2886);
nand U5659 (N_5659,N_3070,N_2801);
or U5660 (N_5660,N_3819,N_3414);
nor U5661 (N_5661,N_2503,N_3897);
and U5662 (N_5662,N_3389,N_2464);
nor U5663 (N_5663,N_2819,N_2162);
or U5664 (N_5664,N_3946,N_3754);
xor U5665 (N_5665,N_2447,N_2106);
nor U5666 (N_5666,N_3799,N_2374);
and U5667 (N_5667,N_2081,N_2582);
and U5668 (N_5668,N_3015,N_2814);
nor U5669 (N_5669,N_3510,N_2578);
nand U5670 (N_5670,N_3951,N_2191);
nor U5671 (N_5671,N_3639,N_3567);
and U5672 (N_5672,N_3257,N_2014);
nor U5673 (N_5673,N_3486,N_3154);
nor U5674 (N_5674,N_3613,N_3509);
nand U5675 (N_5675,N_2416,N_3615);
nand U5676 (N_5676,N_2837,N_3164);
xor U5677 (N_5677,N_3201,N_2168);
nor U5678 (N_5678,N_3612,N_3454);
nand U5679 (N_5679,N_2896,N_3960);
nor U5680 (N_5680,N_3126,N_2005);
nor U5681 (N_5681,N_2618,N_3473);
nor U5682 (N_5682,N_3544,N_3422);
nand U5683 (N_5683,N_2737,N_3038);
nand U5684 (N_5684,N_3620,N_2325);
nand U5685 (N_5685,N_3498,N_2881);
and U5686 (N_5686,N_3158,N_3310);
nor U5687 (N_5687,N_2529,N_3477);
nor U5688 (N_5688,N_3740,N_3801);
nand U5689 (N_5689,N_2665,N_2644);
or U5690 (N_5690,N_3843,N_3150);
nor U5691 (N_5691,N_2057,N_3715);
xnor U5692 (N_5692,N_3990,N_3007);
nor U5693 (N_5693,N_2895,N_3628);
nand U5694 (N_5694,N_3480,N_2616);
nor U5695 (N_5695,N_2181,N_2043);
and U5696 (N_5696,N_2811,N_3083);
nand U5697 (N_5697,N_2794,N_3426);
xor U5698 (N_5698,N_2474,N_2118);
nor U5699 (N_5699,N_2435,N_2580);
or U5700 (N_5700,N_2897,N_3898);
and U5701 (N_5701,N_3131,N_3561);
and U5702 (N_5702,N_2523,N_3847);
and U5703 (N_5703,N_3378,N_2879);
or U5704 (N_5704,N_3977,N_3606);
nand U5705 (N_5705,N_2556,N_3133);
or U5706 (N_5706,N_2973,N_3405);
nor U5707 (N_5707,N_3287,N_2419);
nor U5708 (N_5708,N_2866,N_3781);
nor U5709 (N_5709,N_3193,N_3619);
nor U5710 (N_5710,N_2232,N_2355);
nand U5711 (N_5711,N_3717,N_3498);
nor U5712 (N_5712,N_3469,N_2975);
or U5713 (N_5713,N_3768,N_2905);
and U5714 (N_5714,N_3918,N_3125);
nor U5715 (N_5715,N_3724,N_3749);
or U5716 (N_5716,N_2275,N_3976);
and U5717 (N_5717,N_2729,N_3505);
nor U5718 (N_5718,N_3224,N_3573);
and U5719 (N_5719,N_3446,N_3942);
or U5720 (N_5720,N_3544,N_2411);
or U5721 (N_5721,N_3073,N_3033);
nor U5722 (N_5722,N_2090,N_2579);
or U5723 (N_5723,N_3584,N_2076);
or U5724 (N_5724,N_2405,N_3932);
nand U5725 (N_5725,N_3639,N_3254);
nand U5726 (N_5726,N_3658,N_2196);
nand U5727 (N_5727,N_2142,N_2723);
nor U5728 (N_5728,N_3616,N_3846);
nand U5729 (N_5729,N_3730,N_3505);
and U5730 (N_5730,N_3680,N_2092);
nand U5731 (N_5731,N_3686,N_3161);
nor U5732 (N_5732,N_3540,N_2027);
nand U5733 (N_5733,N_3685,N_2740);
nor U5734 (N_5734,N_3664,N_3002);
or U5735 (N_5735,N_3473,N_3098);
nor U5736 (N_5736,N_2728,N_2206);
nor U5737 (N_5737,N_3380,N_2780);
and U5738 (N_5738,N_2780,N_2187);
and U5739 (N_5739,N_2747,N_3210);
or U5740 (N_5740,N_3751,N_2861);
nand U5741 (N_5741,N_3433,N_3986);
or U5742 (N_5742,N_3404,N_2145);
and U5743 (N_5743,N_2053,N_2620);
or U5744 (N_5744,N_3975,N_3326);
and U5745 (N_5745,N_3972,N_3668);
or U5746 (N_5746,N_3789,N_2736);
or U5747 (N_5747,N_2703,N_2456);
nor U5748 (N_5748,N_2702,N_2427);
and U5749 (N_5749,N_2098,N_2732);
nor U5750 (N_5750,N_3496,N_3101);
and U5751 (N_5751,N_3631,N_2309);
nand U5752 (N_5752,N_2606,N_2834);
and U5753 (N_5753,N_2377,N_2189);
or U5754 (N_5754,N_2286,N_2122);
nand U5755 (N_5755,N_2143,N_3463);
and U5756 (N_5756,N_3471,N_2787);
xor U5757 (N_5757,N_2973,N_2942);
or U5758 (N_5758,N_3927,N_2342);
nor U5759 (N_5759,N_2917,N_2105);
nor U5760 (N_5760,N_3644,N_3886);
nand U5761 (N_5761,N_3844,N_3102);
nand U5762 (N_5762,N_3506,N_2860);
and U5763 (N_5763,N_2118,N_3450);
and U5764 (N_5764,N_3611,N_2299);
nor U5765 (N_5765,N_2686,N_3374);
nand U5766 (N_5766,N_2452,N_3804);
or U5767 (N_5767,N_3158,N_3708);
or U5768 (N_5768,N_3000,N_3189);
and U5769 (N_5769,N_2108,N_3237);
nor U5770 (N_5770,N_2477,N_3717);
or U5771 (N_5771,N_3058,N_3962);
and U5772 (N_5772,N_2929,N_2981);
nand U5773 (N_5773,N_2589,N_2904);
nand U5774 (N_5774,N_3613,N_2300);
nand U5775 (N_5775,N_3975,N_2221);
and U5776 (N_5776,N_2314,N_2551);
and U5777 (N_5777,N_3584,N_3122);
and U5778 (N_5778,N_3159,N_2637);
and U5779 (N_5779,N_3250,N_2963);
or U5780 (N_5780,N_3714,N_2802);
or U5781 (N_5781,N_2648,N_3843);
nand U5782 (N_5782,N_2818,N_3726);
and U5783 (N_5783,N_3871,N_2169);
nor U5784 (N_5784,N_2768,N_2528);
nor U5785 (N_5785,N_2787,N_2240);
xnor U5786 (N_5786,N_3470,N_2147);
nand U5787 (N_5787,N_3077,N_3139);
and U5788 (N_5788,N_2756,N_2267);
nand U5789 (N_5789,N_2584,N_3973);
or U5790 (N_5790,N_3419,N_3767);
or U5791 (N_5791,N_3496,N_3680);
and U5792 (N_5792,N_2755,N_3652);
or U5793 (N_5793,N_3794,N_2518);
and U5794 (N_5794,N_2832,N_2738);
nor U5795 (N_5795,N_3400,N_2974);
nand U5796 (N_5796,N_2271,N_2339);
nor U5797 (N_5797,N_2386,N_3379);
and U5798 (N_5798,N_3260,N_3085);
nand U5799 (N_5799,N_3273,N_3752);
nand U5800 (N_5800,N_3783,N_2146);
or U5801 (N_5801,N_2271,N_3735);
and U5802 (N_5802,N_2479,N_3573);
nand U5803 (N_5803,N_2925,N_2368);
or U5804 (N_5804,N_2718,N_3581);
nor U5805 (N_5805,N_3117,N_3659);
nand U5806 (N_5806,N_2226,N_2501);
nand U5807 (N_5807,N_2529,N_2078);
or U5808 (N_5808,N_3713,N_3828);
nand U5809 (N_5809,N_3081,N_3312);
and U5810 (N_5810,N_3028,N_2612);
and U5811 (N_5811,N_3730,N_3573);
nand U5812 (N_5812,N_2699,N_2268);
nor U5813 (N_5813,N_2503,N_3565);
nand U5814 (N_5814,N_2966,N_3269);
or U5815 (N_5815,N_3480,N_3661);
or U5816 (N_5816,N_3073,N_3195);
and U5817 (N_5817,N_2268,N_2715);
and U5818 (N_5818,N_3127,N_3437);
and U5819 (N_5819,N_2043,N_3555);
and U5820 (N_5820,N_2819,N_3376);
nor U5821 (N_5821,N_2353,N_2254);
nand U5822 (N_5822,N_2769,N_2127);
xor U5823 (N_5823,N_2038,N_3338);
and U5824 (N_5824,N_2303,N_2712);
xnor U5825 (N_5825,N_3069,N_2287);
and U5826 (N_5826,N_2509,N_3932);
nand U5827 (N_5827,N_3734,N_2903);
nor U5828 (N_5828,N_3864,N_3611);
nor U5829 (N_5829,N_3899,N_2312);
or U5830 (N_5830,N_3555,N_3026);
nor U5831 (N_5831,N_2949,N_2428);
or U5832 (N_5832,N_2702,N_3227);
and U5833 (N_5833,N_3939,N_3853);
or U5834 (N_5834,N_2408,N_2388);
nor U5835 (N_5835,N_3723,N_2890);
or U5836 (N_5836,N_3988,N_2920);
nand U5837 (N_5837,N_3061,N_2559);
nand U5838 (N_5838,N_3518,N_2269);
nor U5839 (N_5839,N_2890,N_3629);
and U5840 (N_5840,N_3621,N_2853);
nand U5841 (N_5841,N_2178,N_3523);
nor U5842 (N_5842,N_2001,N_3669);
nand U5843 (N_5843,N_2844,N_3735);
nor U5844 (N_5844,N_2783,N_2053);
and U5845 (N_5845,N_2755,N_3272);
or U5846 (N_5846,N_3195,N_2281);
and U5847 (N_5847,N_3290,N_2861);
xor U5848 (N_5848,N_2850,N_3873);
and U5849 (N_5849,N_2293,N_2441);
nor U5850 (N_5850,N_3849,N_2348);
or U5851 (N_5851,N_2441,N_3657);
nand U5852 (N_5852,N_3789,N_3937);
nor U5853 (N_5853,N_2844,N_2390);
nand U5854 (N_5854,N_3088,N_2127);
nor U5855 (N_5855,N_2894,N_2829);
nand U5856 (N_5856,N_3130,N_2426);
or U5857 (N_5857,N_2991,N_3763);
or U5858 (N_5858,N_3977,N_2923);
nand U5859 (N_5859,N_2816,N_3921);
and U5860 (N_5860,N_3386,N_2138);
nor U5861 (N_5861,N_3347,N_3191);
or U5862 (N_5862,N_2488,N_2046);
and U5863 (N_5863,N_3965,N_2293);
or U5864 (N_5864,N_2019,N_2710);
or U5865 (N_5865,N_3854,N_3437);
or U5866 (N_5866,N_3247,N_3264);
nand U5867 (N_5867,N_3240,N_2943);
nand U5868 (N_5868,N_2168,N_2939);
and U5869 (N_5869,N_3975,N_3715);
and U5870 (N_5870,N_2199,N_2604);
nor U5871 (N_5871,N_3773,N_3569);
nand U5872 (N_5872,N_3532,N_3472);
and U5873 (N_5873,N_3778,N_2713);
or U5874 (N_5874,N_3810,N_3461);
and U5875 (N_5875,N_3208,N_2288);
nor U5876 (N_5876,N_2150,N_3555);
and U5877 (N_5877,N_2782,N_3883);
nor U5878 (N_5878,N_3616,N_3561);
nor U5879 (N_5879,N_3742,N_3589);
and U5880 (N_5880,N_3105,N_3336);
nand U5881 (N_5881,N_2925,N_2699);
or U5882 (N_5882,N_2479,N_3410);
and U5883 (N_5883,N_3310,N_2185);
nor U5884 (N_5884,N_2334,N_3135);
nand U5885 (N_5885,N_2993,N_3740);
or U5886 (N_5886,N_2010,N_2054);
nand U5887 (N_5887,N_3241,N_3806);
nor U5888 (N_5888,N_2384,N_2273);
and U5889 (N_5889,N_2339,N_3821);
or U5890 (N_5890,N_2727,N_2353);
and U5891 (N_5891,N_2953,N_2077);
nand U5892 (N_5892,N_3427,N_3880);
nand U5893 (N_5893,N_2677,N_2542);
nand U5894 (N_5894,N_3160,N_3673);
nand U5895 (N_5895,N_3193,N_2610);
or U5896 (N_5896,N_3939,N_3242);
or U5897 (N_5897,N_2755,N_3445);
and U5898 (N_5898,N_2218,N_2941);
nand U5899 (N_5899,N_3209,N_3641);
nor U5900 (N_5900,N_2575,N_2226);
and U5901 (N_5901,N_2998,N_2238);
and U5902 (N_5902,N_3542,N_2683);
and U5903 (N_5903,N_3225,N_3117);
nor U5904 (N_5904,N_2366,N_3821);
nor U5905 (N_5905,N_3995,N_2450);
and U5906 (N_5906,N_2888,N_2920);
and U5907 (N_5907,N_3081,N_3308);
xnor U5908 (N_5908,N_2896,N_2563);
or U5909 (N_5909,N_3812,N_3389);
nor U5910 (N_5910,N_2681,N_3518);
or U5911 (N_5911,N_3670,N_3694);
nand U5912 (N_5912,N_3010,N_2030);
xor U5913 (N_5913,N_2140,N_3752);
or U5914 (N_5914,N_2384,N_2904);
or U5915 (N_5915,N_3798,N_3934);
nand U5916 (N_5916,N_2287,N_2714);
nor U5917 (N_5917,N_2822,N_3248);
and U5918 (N_5918,N_2911,N_2829);
nor U5919 (N_5919,N_3005,N_2673);
or U5920 (N_5920,N_3199,N_2266);
and U5921 (N_5921,N_2547,N_2465);
xnor U5922 (N_5922,N_2155,N_2259);
or U5923 (N_5923,N_3844,N_3388);
nand U5924 (N_5924,N_3233,N_2628);
and U5925 (N_5925,N_3410,N_3201);
and U5926 (N_5926,N_3470,N_3654);
nor U5927 (N_5927,N_2515,N_2093);
and U5928 (N_5928,N_2418,N_3295);
or U5929 (N_5929,N_3252,N_2784);
nor U5930 (N_5930,N_2300,N_3147);
and U5931 (N_5931,N_3054,N_3329);
or U5932 (N_5932,N_3057,N_2173);
nand U5933 (N_5933,N_3316,N_3247);
nor U5934 (N_5934,N_2893,N_3111);
nor U5935 (N_5935,N_2341,N_2637);
and U5936 (N_5936,N_2471,N_3004);
and U5937 (N_5937,N_3856,N_3130);
and U5938 (N_5938,N_3708,N_2180);
nand U5939 (N_5939,N_2148,N_3983);
nor U5940 (N_5940,N_2148,N_3661);
or U5941 (N_5941,N_2991,N_2506);
or U5942 (N_5942,N_3452,N_3639);
and U5943 (N_5943,N_2677,N_2779);
nand U5944 (N_5944,N_3171,N_3054);
and U5945 (N_5945,N_3607,N_2119);
nand U5946 (N_5946,N_3594,N_3884);
or U5947 (N_5947,N_2658,N_3227);
nor U5948 (N_5948,N_3372,N_2018);
nor U5949 (N_5949,N_2310,N_2736);
or U5950 (N_5950,N_2414,N_2007);
or U5951 (N_5951,N_2630,N_3150);
nor U5952 (N_5952,N_3170,N_3132);
and U5953 (N_5953,N_3394,N_3673);
nor U5954 (N_5954,N_2910,N_2102);
or U5955 (N_5955,N_2988,N_2411);
xor U5956 (N_5956,N_2248,N_2485);
and U5957 (N_5957,N_3130,N_2180);
nand U5958 (N_5958,N_2246,N_2171);
nand U5959 (N_5959,N_2323,N_2173);
or U5960 (N_5960,N_2500,N_3468);
or U5961 (N_5961,N_2919,N_3745);
nor U5962 (N_5962,N_3362,N_2506);
nand U5963 (N_5963,N_3929,N_2524);
or U5964 (N_5964,N_2768,N_2739);
nor U5965 (N_5965,N_2745,N_2110);
nor U5966 (N_5966,N_3471,N_2092);
or U5967 (N_5967,N_2084,N_3659);
nor U5968 (N_5968,N_2632,N_2924);
nor U5969 (N_5969,N_2732,N_2791);
nor U5970 (N_5970,N_3050,N_2865);
and U5971 (N_5971,N_3020,N_2685);
nor U5972 (N_5972,N_2037,N_3198);
nand U5973 (N_5973,N_2358,N_2736);
nor U5974 (N_5974,N_3775,N_2918);
nand U5975 (N_5975,N_3669,N_3965);
and U5976 (N_5976,N_3040,N_3480);
nand U5977 (N_5977,N_2224,N_3265);
xnor U5978 (N_5978,N_3160,N_2888);
nor U5979 (N_5979,N_2590,N_2464);
nand U5980 (N_5980,N_3874,N_2163);
or U5981 (N_5981,N_3982,N_3935);
nor U5982 (N_5982,N_2879,N_3846);
or U5983 (N_5983,N_3313,N_2081);
nand U5984 (N_5984,N_2639,N_2338);
and U5985 (N_5985,N_3353,N_3669);
or U5986 (N_5986,N_3104,N_2710);
nor U5987 (N_5987,N_2579,N_3559);
nand U5988 (N_5988,N_2205,N_2579);
and U5989 (N_5989,N_2827,N_3888);
or U5990 (N_5990,N_2029,N_3542);
nand U5991 (N_5991,N_2477,N_2029);
nor U5992 (N_5992,N_3803,N_3774);
or U5993 (N_5993,N_3405,N_3362);
nor U5994 (N_5994,N_2138,N_2803);
nand U5995 (N_5995,N_3343,N_3412);
or U5996 (N_5996,N_3218,N_3280);
and U5997 (N_5997,N_3137,N_2332);
and U5998 (N_5998,N_2912,N_2648);
or U5999 (N_5999,N_2135,N_3218);
nor U6000 (N_6000,N_5337,N_5914);
or U6001 (N_6001,N_4465,N_5974);
nor U6002 (N_6002,N_4380,N_4159);
nand U6003 (N_6003,N_5441,N_4880);
nor U6004 (N_6004,N_4117,N_5215);
nor U6005 (N_6005,N_5066,N_4344);
nand U6006 (N_6006,N_4251,N_4663);
and U6007 (N_6007,N_4543,N_4078);
or U6008 (N_6008,N_4626,N_4444);
or U6009 (N_6009,N_4792,N_4167);
nand U6010 (N_6010,N_5932,N_4305);
nand U6011 (N_6011,N_4328,N_5274);
nand U6012 (N_6012,N_4490,N_5519);
or U6013 (N_6013,N_4058,N_5963);
nand U6014 (N_6014,N_4367,N_5820);
nand U6015 (N_6015,N_5291,N_5767);
nor U6016 (N_6016,N_5443,N_4314);
or U6017 (N_6017,N_5709,N_4243);
and U6018 (N_6018,N_4487,N_4226);
and U6019 (N_6019,N_4933,N_5080);
nor U6020 (N_6020,N_5206,N_4410);
or U6021 (N_6021,N_4787,N_4870);
nor U6022 (N_6022,N_4469,N_5877);
nor U6023 (N_6023,N_4640,N_5711);
and U6024 (N_6024,N_4704,N_5892);
nand U6025 (N_6025,N_5158,N_5193);
nor U6026 (N_6026,N_5115,N_4241);
or U6027 (N_6027,N_4895,N_4178);
and U6028 (N_6028,N_4074,N_5937);
or U6029 (N_6029,N_5393,N_4807);
or U6030 (N_6030,N_5414,N_5145);
or U6031 (N_6031,N_4882,N_4146);
or U6032 (N_6032,N_4100,N_5675);
or U6033 (N_6033,N_4655,N_4789);
nand U6034 (N_6034,N_5303,N_4841);
or U6035 (N_6035,N_5517,N_5059);
or U6036 (N_6036,N_4397,N_5299);
and U6037 (N_6037,N_4061,N_4160);
nor U6038 (N_6038,N_5972,N_5791);
or U6039 (N_6039,N_4554,N_4216);
nand U6040 (N_6040,N_5968,N_4550);
or U6041 (N_6041,N_5072,N_4921);
and U6042 (N_6042,N_5379,N_5246);
nand U6043 (N_6043,N_5812,N_5620);
nand U6044 (N_6044,N_4953,N_4233);
nand U6045 (N_6045,N_4671,N_4264);
nor U6046 (N_6046,N_4588,N_5221);
nand U6047 (N_6047,N_4327,N_5686);
or U6048 (N_6048,N_4986,N_4449);
nor U6049 (N_6049,N_4248,N_5452);
or U6050 (N_6050,N_5341,N_5903);
or U6051 (N_6051,N_5887,N_5752);
and U6052 (N_6052,N_5876,N_5084);
and U6053 (N_6053,N_4832,N_4702);
nand U6054 (N_6054,N_4125,N_5495);
nand U6055 (N_6055,N_5964,N_5200);
nand U6056 (N_6056,N_4130,N_4309);
xnor U6057 (N_6057,N_5902,N_4811);
nand U6058 (N_6058,N_4959,N_4416);
nor U6059 (N_6059,N_4362,N_4040);
nor U6060 (N_6060,N_4334,N_4985);
and U6061 (N_6061,N_4276,N_4786);
nor U6062 (N_6062,N_5491,N_4637);
nor U6063 (N_6063,N_5535,N_4573);
and U6064 (N_6064,N_4038,N_5021);
and U6065 (N_6065,N_4854,N_5800);
and U6066 (N_6066,N_4105,N_4129);
and U6067 (N_6067,N_5760,N_4437);
nor U6068 (N_6068,N_4068,N_5797);
nand U6069 (N_6069,N_4945,N_5631);
and U6070 (N_6070,N_4548,N_4127);
nor U6071 (N_6071,N_5566,N_5543);
xor U6072 (N_6072,N_4358,N_5060);
nand U6073 (N_6073,N_5858,N_4732);
or U6074 (N_6074,N_4725,N_5473);
nand U6075 (N_6075,N_5068,N_5598);
or U6076 (N_6076,N_5014,N_4631);
nor U6077 (N_6077,N_4915,N_4360);
nand U6078 (N_6078,N_4684,N_5548);
and U6079 (N_6079,N_4996,N_5195);
nor U6080 (N_6080,N_5478,N_4477);
nand U6081 (N_6081,N_5981,N_4612);
nor U6082 (N_6082,N_5666,N_4376);
and U6083 (N_6083,N_5328,N_4292);
nand U6084 (N_6084,N_5449,N_4135);
nor U6085 (N_6085,N_5415,N_5198);
and U6086 (N_6086,N_4995,N_5496);
nor U6087 (N_6087,N_5288,N_5143);
or U6088 (N_6088,N_4253,N_5657);
or U6089 (N_6089,N_5971,N_5308);
and U6090 (N_6090,N_4373,N_4116);
nor U6091 (N_6091,N_5107,N_4949);
or U6092 (N_6092,N_5833,N_5326);
nand U6093 (N_6093,N_4443,N_5640);
nand U6094 (N_6094,N_4692,N_5925);
or U6095 (N_6095,N_4955,N_4194);
nand U6096 (N_6096,N_5584,N_4330);
nor U6097 (N_6097,N_4186,N_5644);
and U6098 (N_6098,N_5431,N_5210);
nand U6099 (N_6099,N_4516,N_5660);
and U6100 (N_6100,N_4095,N_5184);
and U6101 (N_6101,N_4374,N_4859);
or U6102 (N_6102,N_5875,N_4559);
or U6103 (N_6103,N_5942,N_4576);
nand U6104 (N_6104,N_4746,N_4418);
nor U6105 (N_6105,N_4413,N_4150);
nand U6106 (N_6106,N_4674,N_4969);
nor U6107 (N_6107,N_4153,N_4780);
nor U6108 (N_6108,N_5838,N_5081);
nand U6109 (N_6109,N_5088,N_4467);
xnor U6110 (N_6110,N_4500,N_5306);
nand U6111 (N_6111,N_4273,N_4521);
and U6112 (N_6112,N_4258,N_4365);
nor U6113 (N_6113,N_5146,N_5841);
nor U6114 (N_6114,N_4428,N_5343);
or U6115 (N_6115,N_5224,N_5798);
nor U6116 (N_6116,N_4102,N_5777);
and U6117 (N_6117,N_5094,N_4662);
nand U6118 (N_6118,N_5695,N_4765);
and U6119 (N_6119,N_5279,N_5975);
nand U6120 (N_6120,N_4885,N_5626);
or U6121 (N_6121,N_5842,N_5715);
nand U6122 (N_6122,N_5860,N_5751);
nor U6123 (N_6123,N_4349,N_4904);
nand U6124 (N_6124,N_4999,N_4733);
or U6125 (N_6125,N_4658,N_4383);
nand U6126 (N_6126,N_4705,N_5119);
nor U6127 (N_6127,N_4110,N_5104);
nor U6128 (N_6128,N_5289,N_4438);
and U6129 (N_6129,N_4647,N_4024);
nand U6130 (N_6130,N_5102,N_5037);
nand U6131 (N_6131,N_4246,N_5216);
nor U6132 (N_6132,N_4666,N_5499);
and U6133 (N_6133,N_5966,N_4983);
nand U6134 (N_6134,N_5240,N_4862);
and U6135 (N_6135,N_4526,N_5806);
or U6136 (N_6136,N_5559,N_4575);
or U6137 (N_6137,N_5136,N_4389);
or U6138 (N_6138,N_4336,N_5978);
nand U6139 (N_6139,N_4615,N_4403);
nor U6140 (N_6140,N_5128,N_5827);
and U6141 (N_6141,N_5673,N_4254);
nor U6142 (N_6142,N_5888,N_5911);
nor U6143 (N_6143,N_4475,N_5690);
nand U6144 (N_6144,N_4053,N_5948);
and U6145 (N_6145,N_5542,N_5993);
and U6146 (N_6146,N_4242,N_5696);
or U6147 (N_6147,N_5560,N_5900);
nor U6148 (N_6148,N_4103,N_5167);
and U6149 (N_6149,N_4407,N_5395);
and U6150 (N_6150,N_5041,N_4990);
and U6151 (N_6151,N_4463,N_4071);
and U6152 (N_6152,N_4917,N_5718);
or U6153 (N_6153,N_4998,N_5509);
or U6154 (N_6154,N_4506,N_4422);
nor U6155 (N_6155,N_4051,N_5223);
nor U6156 (N_6156,N_5386,N_4865);
nor U6157 (N_6157,N_4343,N_4960);
nor U6158 (N_6158,N_4080,N_5671);
nand U6159 (N_6159,N_4141,N_5672);
and U6160 (N_6160,N_5537,N_4440);
nor U6161 (N_6161,N_5321,N_5346);
or U6162 (N_6162,N_4517,N_4082);
or U6163 (N_6163,N_5831,N_4022);
nor U6164 (N_6164,N_4479,N_5073);
and U6165 (N_6165,N_4085,N_4262);
and U6166 (N_6166,N_5748,N_4011);
nand U6167 (N_6167,N_5263,N_4333);
or U6168 (N_6168,N_5460,N_5528);
nand U6169 (N_6169,N_5042,N_4583);
nand U6170 (N_6170,N_5416,N_4472);
nor U6171 (N_6171,N_4866,N_4451);
nor U6172 (N_6172,N_4412,N_5407);
and U6173 (N_6173,N_5179,N_4355);
nor U6174 (N_6174,N_4297,N_4822);
nand U6175 (N_6175,N_4363,N_5356);
xnor U6176 (N_6176,N_4873,N_5025);
and U6177 (N_6177,N_5728,N_5749);
or U6178 (N_6178,N_4687,N_5765);
nor U6179 (N_6179,N_5141,N_4607);
xor U6180 (N_6180,N_4527,N_4834);
or U6181 (N_6181,N_5684,N_5522);
and U6182 (N_6182,N_4280,N_5430);
and U6183 (N_6183,N_4329,N_5648);
nand U6184 (N_6184,N_5761,N_5110);
nand U6185 (N_6185,N_5867,N_5924);
nand U6186 (N_6186,N_5811,N_5227);
or U6187 (N_6187,N_5050,N_4567);
or U6188 (N_6188,N_4016,N_5608);
nand U6189 (N_6189,N_4419,N_5864);
and U6190 (N_6190,N_4402,N_4689);
xnor U6191 (N_6191,N_4197,N_4592);
nor U6192 (N_6192,N_4934,N_5387);
xor U6193 (N_6193,N_4525,N_5455);
and U6194 (N_6194,N_5744,N_4657);
and U6195 (N_6195,N_4207,N_5795);
nor U6196 (N_6196,N_4686,N_5471);
or U6197 (N_6197,N_4529,N_5355);
nor U6198 (N_6198,N_4505,N_5302);
nand U6199 (N_6199,N_4200,N_5470);
nor U6200 (N_6200,N_5890,N_4668);
nor U6201 (N_6201,N_4177,N_4111);
and U6202 (N_6202,N_5220,N_5380);
nand U6203 (N_6203,N_4726,N_4813);
nand U6204 (N_6204,N_5627,N_4137);
nand U6205 (N_6205,N_5362,N_5276);
nand U6206 (N_6206,N_5917,N_5861);
and U6207 (N_6207,N_5889,N_5687);
or U6208 (N_6208,N_4988,N_4743);
nand U6209 (N_6209,N_5821,N_5769);
nor U6210 (N_6210,N_4709,N_4259);
nand U6211 (N_6211,N_5004,N_4325);
nand U6212 (N_6212,N_4954,N_5638);
nand U6213 (N_6213,N_4348,N_5207);
nand U6214 (N_6214,N_4599,N_4989);
or U6215 (N_6215,N_4893,N_4978);
nand U6216 (N_6216,N_5152,N_5348);
and U6217 (N_6217,N_5586,N_4131);
nor U6218 (N_6218,N_4369,N_5707);
or U6219 (N_6219,N_5316,N_5610);
or U6220 (N_6220,N_4508,N_4232);
or U6221 (N_6221,N_4690,N_4790);
and U6222 (N_6222,N_5052,N_4044);
nor U6223 (N_6223,N_4315,N_4851);
nand U6224 (N_6224,N_4468,N_4648);
and U6225 (N_6225,N_5336,N_5815);
nor U6226 (N_6226,N_5197,N_5730);
or U6227 (N_6227,N_5534,N_5540);
nor U6228 (N_6228,N_4126,N_5565);
xnor U6229 (N_6229,N_5661,N_4208);
or U6230 (N_6230,N_5603,N_4268);
and U6231 (N_6231,N_5219,N_4619);
and U6232 (N_6232,N_4287,N_5365);
nand U6233 (N_6233,N_4547,N_4481);
and U6234 (N_6234,N_5309,N_5401);
nor U6235 (N_6235,N_5421,N_5249);
or U6236 (N_6236,N_5307,N_5419);
xor U6237 (N_6237,N_4542,N_4156);
and U6238 (N_6238,N_4981,N_4749);
nand U6239 (N_6239,N_5771,N_5413);
or U6240 (N_6240,N_4238,N_4830);
and U6241 (N_6241,N_5217,N_4182);
nand U6242 (N_6242,N_5970,N_5774);
nand U6243 (N_6243,N_5539,N_4015);
and U6244 (N_6244,N_5446,N_4947);
nor U6245 (N_6245,N_4083,N_5149);
and U6246 (N_6246,N_4964,N_4997);
nand U6247 (N_6247,N_5254,N_4215);
nand U6248 (N_6248,N_5040,N_4871);
and U6249 (N_6249,N_4639,N_4203);
xnor U6250 (N_6250,N_4828,N_4884);
xnor U6251 (N_6251,N_4499,N_5766);
nand U6252 (N_6252,N_4535,N_4014);
and U6253 (N_6253,N_4918,N_4942);
nand U6254 (N_6254,N_4594,N_4544);
nand U6255 (N_6255,N_4638,N_4236);
nor U6256 (N_6256,N_4426,N_5936);
nor U6257 (N_6257,N_5454,N_5371);
nor U6258 (N_6258,N_5778,N_5015);
and U6259 (N_6259,N_4758,N_4553);
nand U6260 (N_6260,N_4844,N_5133);
and U6261 (N_6261,N_5743,N_5712);
and U6262 (N_6262,N_4204,N_4518);
or U6263 (N_6263,N_5609,N_4541);
or U6264 (N_6264,N_5654,N_5893);
and U6265 (N_6265,N_5783,N_4935);
and U6266 (N_6266,N_4555,N_4166);
nor U6267 (N_6267,N_4134,N_5301);
or U6268 (N_6268,N_4461,N_4042);
and U6269 (N_6269,N_5445,N_5029);
nor U6270 (N_6270,N_4067,N_5868);
and U6271 (N_6271,N_5720,N_5422);
and U6272 (N_6272,N_4019,N_5637);
nand U6273 (N_6273,N_5991,N_5009);
and U6274 (N_6274,N_5725,N_5006);
or U6275 (N_6275,N_5226,N_5116);
and U6276 (N_6276,N_4906,N_5030);
or U6277 (N_6277,N_5855,N_5679);
nor U6278 (N_6278,N_5161,N_5634);
nor U6279 (N_6279,N_5469,N_5142);
or U6280 (N_6280,N_4411,N_5733);
or U6281 (N_6281,N_5947,N_5112);
nand U6282 (N_6282,N_4266,N_4063);
or U6283 (N_6283,N_4275,N_4578);
or U6284 (N_6284,N_4534,N_5448);
or U6285 (N_6285,N_5385,N_5324);
and U6286 (N_6286,N_4605,N_4353);
nand U6287 (N_6287,N_5781,N_4730);
or U6288 (N_6288,N_4055,N_5245);
nand U6289 (N_6289,N_5992,N_4609);
and U6290 (N_6290,N_5989,N_4625);
or U6291 (N_6291,N_5588,N_4825);
or U6292 (N_6292,N_4218,N_4887);
nand U6293 (N_6293,N_4342,N_5320);
and U6294 (N_6294,N_4504,N_5344);
nor U6295 (N_6295,N_5429,N_5949);
nor U6296 (N_6296,N_4277,N_4048);
or U6297 (N_6297,N_4294,N_5463);
nor U6298 (N_6298,N_5375,N_4591);
or U6299 (N_6299,N_4614,N_4433);
nand U6300 (N_6300,N_4711,N_4486);
nor U6301 (N_6301,N_4975,N_4772);
nor U6302 (N_6302,N_5294,N_5525);
or U6303 (N_6303,N_5390,N_4029);
or U6304 (N_6304,N_4770,N_4084);
or U6305 (N_6305,N_4323,N_5601);
nand U6306 (N_6306,N_5689,N_4184);
nand U6307 (N_6307,N_4435,N_5782);
nor U6308 (N_6308,N_5898,N_4718);
nand U6309 (N_6309,N_4032,N_5959);
or U6310 (N_6310,N_4919,N_5808);
and U6311 (N_6311,N_4809,N_5359);
and U6312 (N_6312,N_5201,N_5374);
or U6313 (N_6313,N_5138,N_5378);
and U6314 (N_6314,N_5427,N_5552);
nand U6315 (N_6315,N_4179,N_5182);
and U6316 (N_6316,N_4923,N_4282);
nor U6317 (N_6317,N_5700,N_5651);
or U6318 (N_6318,N_4391,N_4524);
nand U6319 (N_6319,N_4863,N_4723);
or U6320 (N_6320,N_5794,N_5181);
nor U6321 (N_6321,N_5439,N_4217);
nor U6322 (N_6322,N_4028,N_5281);
and U6323 (N_6323,N_5754,N_4027);
nor U6324 (N_6324,N_5273,N_5531);
nor U6325 (N_6325,N_5434,N_4821);
or U6326 (N_6326,N_5101,N_5545);
nand U6327 (N_6327,N_4109,N_5590);
and U6328 (N_6328,N_5114,N_5096);
nor U6329 (N_6329,N_4375,N_4528);
nor U6330 (N_6330,N_4677,N_4898);
nor U6331 (N_6331,N_5367,N_5252);
and U6332 (N_6332,N_4581,N_5646);
or U6333 (N_6333,N_4453,N_5406);
and U6334 (N_6334,N_4768,N_5502);
xnor U6335 (N_6335,N_5053,N_4227);
xor U6336 (N_6336,N_5484,N_5597);
or U6337 (N_6337,N_4783,N_4318);
nor U6338 (N_6338,N_5412,N_5802);
or U6339 (N_6339,N_4002,N_4800);
or U6340 (N_6340,N_5553,N_4021);
or U6341 (N_6341,N_5810,N_5488);
nand U6342 (N_6342,N_4742,N_5756);
nor U6343 (N_6343,N_5804,N_5705);
and U6344 (N_6344,N_5726,N_4874);
or U6345 (N_6345,N_5587,N_5938);
nor U6346 (N_6346,N_5879,N_4447);
xnor U6347 (N_6347,N_4691,N_5943);
and U6348 (N_6348,N_5571,N_5173);
and U6349 (N_6349,N_4875,N_5438);
nand U6350 (N_6350,N_5662,N_5747);
and U6351 (N_6351,N_5475,N_5830);
or U6352 (N_6352,N_5961,N_5490);
and U6353 (N_6353,N_5514,N_5614);
nor U6354 (N_6354,N_5247,N_5214);
and U6355 (N_6355,N_4206,N_5000);
or U6356 (N_6356,N_4271,N_4423);
nand U6357 (N_6357,N_4406,N_5319);
or U6358 (N_6358,N_4722,N_5127);
xnor U6359 (N_6359,N_5596,N_4124);
or U6360 (N_6360,N_5391,N_5740);
and U6361 (N_6361,N_4198,N_4039);
nand U6362 (N_6362,N_4812,N_4927);
nor U6363 (N_6363,N_5061,N_5134);
nand U6364 (N_6364,N_5347,N_5039);
and U6365 (N_6365,N_5916,N_5853);
nor U6366 (N_6366,N_5624,N_4710);
nand U6367 (N_6367,N_5501,N_5880);
nand U6368 (N_6368,N_4636,N_5846);
and U6369 (N_6369,N_4698,N_4034);
and U6370 (N_6370,N_5186,N_5950);
nor U6371 (N_6371,N_4739,N_5919);
and U6372 (N_6372,N_4755,N_5757);
nand U6373 (N_6373,N_4572,N_5418);
nand U6374 (N_6374,N_4260,N_4191);
nor U6375 (N_6375,N_4714,N_5529);
nand U6376 (N_6376,N_4774,N_5459);
xnor U6377 (N_6377,N_4304,N_4628);
nand U6378 (N_6378,N_5232,N_4172);
nor U6379 (N_6379,N_4672,N_4688);
and U6380 (N_6380,N_4026,N_4401);
and U6381 (N_6381,N_4400,N_4269);
nor U6382 (N_6382,N_4209,N_5283);
or U6383 (N_6383,N_4897,N_5054);
nand U6384 (N_6384,N_4478,N_5047);
or U6385 (N_6385,N_4890,N_4202);
and U6386 (N_6386,N_5140,N_5954);
and U6387 (N_6387,N_4760,N_4793);
or U6388 (N_6388,N_5241,N_5826);
nor U6389 (N_6389,N_5476,N_5716);
nor U6390 (N_6390,N_5650,N_5489);
or U6391 (N_6391,N_4138,N_4624);
xnor U6392 (N_6392,N_5659,N_5485);
nand U6393 (N_6393,N_5480,N_4660);
and U6394 (N_6394,N_5417,N_4498);
or U6395 (N_6395,N_4052,N_5334);
and U6396 (N_6396,N_4370,N_5062);
and U6397 (N_6397,N_4415,N_4932);
or U6398 (N_6398,N_5844,N_4128);
nand U6399 (N_6399,N_4247,N_5033);
nand U6400 (N_6400,N_5595,N_5031);
or U6401 (N_6401,N_5298,N_4149);
or U6402 (N_6402,N_4551,N_4993);
and U6403 (N_6403,N_4359,N_5594);
xor U6404 (N_6404,N_4377,N_5960);
nor U6405 (N_6405,N_5670,N_5100);
and U6406 (N_6406,N_4840,N_4905);
xnor U6407 (N_6407,N_5639,N_5296);
nor U6408 (N_6408,N_5456,N_5847);
or U6409 (N_6409,N_4940,N_5776);
and U6410 (N_6410,N_4701,N_5300);
or U6411 (N_6411,N_5792,N_5250);
and U6412 (N_6412,N_5849,N_5945);
and U6413 (N_6413,N_4916,N_4261);
and U6414 (N_6414,N_4798,N_5225);
nand U6415 (N_6415,N_5388,N_5891);
nor U6416 (N_6416,N_5222,N_4424);
and U6417 (N_6417,N_5951,N_4968);
or U6418 (N_6418,N_5151,N_4912);
nand U6419 (N_6419,N_5667,N_4777);
nor U6420 (N_6420,N_4913,N_5233);
and U6421 (N_6421,N_4480,N_5965);
and U6422 (N_6422,N_5618,N_4741);
or U6423 (N_6423,N_4627,N_5315);
nor U6424 (N_6424,N_4381,N_5866);
or U6425 (N_6425,N_4914,N_5688);
and U6426 (N_6426,N_4221,N_5286);
and U6427 (N_6427,N_4069,N_4823);
or U6428 (N_6428,N_4971,N_4496);
and U6429 (N_6429,N_5275,N_5038);
nor U6430 (N_6430,N_5918,N_5404);
or U6431 (N_6431,N_4861,N_5836);
or U6432 (N_6432,N_4845,N_4006);
or U6433 (N_6433,N_4899,N_5996);
nor U6434 (N_6434,N_4796,N_4173);
or U6435 (N_6435,N_4119,N_5630);
nor U6436 (N_6436,N_5024,N_4574);
or U6437 (N_6437,N_4556,N_5230);
nor U6438 (N_6438,N_5423,N_4031);
and U6439 (N_6439,N_5086,N_4509);
nor U6440 (N_6440,N_4511,N_4560);
and U6441 (N_6441,N_5051,N_5763);
nor U6442 (N_6442,N_4601,N_5332);
or U6443 (N_6443,N_4060,N_4858);
and U6444 (N_6444,N_5779,N_5585);
nand U6445 (N_6445,N_4970,N_5611);
or U6446 (N_6446,N_4492,N_4267);
nand U6447 (N_6447,N_5424,N_4099);
and U6448 (N_6448,N_4810,N_5358);
or U6449 (N_6449,N_4645,N_5708);
nor U6450 (N_6450,N_5056,N_5635);
or U6451 (N_6451,N_4434,N_5739);
nor U6452 (N_6452,N_5479,N_4962);
nand U6453 (N_6453,N_5510,N_4944);
nand U6454 (N_6454,N_5257,N_5238);
or U6455 (N_6455,N_4293,N_5530);
nor U6456 (N_6456,N_4966,N_4713);
nor U6457 (N_6457,N_5462,N_4168);
nor U6458 (N_6458,N_4386,N_5856);
nand U6459 (N_6459,N_5305,N_4093);
and U6460 (N_6460,N_4096,N_4075);
and U6461 (N_6461,N_4864,N_5255);
and U6462 (N_6462,N_4231,N_4421);
or U6463 (N_6463,N_4171,N_4092);
nand U6464 (N_6464,N_5381,N_4345);
nand U6465 (N_6465,N_4902,N_5269);
or U6466 (N_6466,N_5985,N_4808);
or U6467 (N_6467,N_4473,N_4888);
nand U6468 (N_6468,N_5885,N_5389);
nand U6469 (N_6469,N_4900,N_5126);
nand U6470 (N_6470,N_5568,N_5704);
nand U6471 (N_6471,N_4488,N_5472);
nand U6472 (N_6472,N_4289,N_5411);
nor U6473 (N_6473,N_5825,N_5894);
or U6474 (N_6474,N_5262,N_4081);
and U6475 (N_6475,N_4321,N_5976);
and U6476 (N_6476,N_5027,N_4489);
nor U6477 (N_6477,N_4680,N_4540);
and U6478 (N_6478,N_5314,N_5664);
nor U6479 (N_6479,N_5373,N_4673);
nand U6480 (N_6480,N_5713,N_5135);
nand U6481 (N_6481,N_4169,N_4459);
and U6482 (N_6482,N_4234,N_4351);
or U6483 (N_6483,N_5617,N_4963);
nand U6484 (N_6484,N_5939,N_4512);
or U6485 (N_6485,N_4728,N_5155);
and U6486 (N_6486,N_4946,N_4339);
nor U6487 (N_6487,N_5979,N_5005);
and U6488 (N_6488,N_4311,N_5863);
or U6489 (N_6489,N_5615,N_4757);
xnor U6490 (N_6490,N_5816,N_5737);
nand U6491 (N_6491,N_4815,N_4967);
or U6492 (N_6492,N_5677,N_5619);
nand U6493 (N_6493,N_5928,N_5492);
nor U6494 (N_6494,N_4062,N_5998);
nor U6495 (N_6495,N_5335,N_5461);
nand U6496 (N_6496,N_4632,N_4335);
nor U6497 (N_6497,N_5208,N_4883);
and U6498 (N_6498,N_5370,N_5962);
nor U6499 (N_6499,N_5987,N_4445);
xnor U6500 (N_6500,N_5398,N_4452);
nor U6501 (N_6501,N_5655,N_4826);
nor U6502 (N_6502,N_4154,N_5645);
or U6503 (N_6503,N_4427,N_5809);
or U6504 (N_6504,N_4901,N_5194);
or U6505 (N_6505,N_5676,N_5997);
or U6506 (N_6506,N_4641,N_5032);
or U6507 (N_6507,N_5106,N_5253);
and U6508 (N_6508,N_5043,N_5357);
and U6509 (N_6509,N_5526,N_4991);
or U6510 (N_6510,N_4079,N_4608);
nor U6511 (N_6511,N_4066,N_4337);
nor U6512 (N_6512,N_4889,N_5131);
nor U6513 (N_6513,N_5921,N_5506);
and U6514 (N_6514,N_5329,N_5327);
nor U6515 (N_6515,N_5019,N_4903);
or U6516 (N_6516,N_4302,N_4176);
and U6517 (N_6517,N_5768,N_5498);
or U6518 (N_6518,N_5244,N_4519);
xnor U6519 (N_6519,N_5160,N_4721);
nor U6520 (N_6520,N_5159,N_5504);
and U6521 (N_6521,N_4561,N_4417);
nand U6522 (N_6522,N_4307,N_5697);
nor U6523 (N_6523,N_4892,N_4513);
or U6524 (N_6524,N_4552,N_4706);
nor U6525 (N_6525,N_4533,N_4773);
nor U6526 (N_6526,N_5403,N_5701);
nor U6527 (N_6527,N_4976,N_5234);
nor U6528 (N_6528,N_4121,N_5563);
and U6529 (N_6529,N_4364,N_5691);
or U6530 (N_6530,N_5909,N_4497);
nor U6531 (N_6531,N_4462,N_4908);
nand U6532 (N_6532,N_4057,N_4522);
nor U6533 (N_6533,N_5538,N_4797);
and U6534 (N_6534,N_5188,N_5266);
nand U6535 (N_6535,N_5083,N_4244);
and U6536 (N_6536,N_4012,N_4939);
or U6537 (N_6537,N_5272,N_4784);
nand U6538 (N_6538,N_4170,N_4211);
and U6539 (N_6539,N_4008,N_5067);
or U6540 (N_6540,N_4087,N_4485);
nor U6541 (N_6541,N_4623,N_5085);
or U6542 (N_6542,N_5518,N_5466);
nand U6543 (N_6543,N_5507,N_4001);
nand U6544 (N_6544,N_4779,N_4388);
and U6545 (N_6545,N_4201,N_4751);
nor U6546 (N_6546,N_4643,N_5770);
nor U6547 (N_6547,N_4164,N_5762);
or U6548 (N_6548,N_4752,N_4196);
and U6549 (N_6549,N_5310,N_4886);
nor U6550 (N_6550,N_4539,N_5178);
and U6551 (N_6551,N_5541,N_5555);
nor U6552 (N_6552,N_4795,N_5564);
and U6553 (N_6553,N_5036,N_5579);
nor U6554 (N_6554,N_5270,N_5722);
or U6555 (N_6555,N_4018,N_5817);
or U6556 (N_6556,N_5350,N_4157);
and U6557 (N_6557,N_4466,N_5828);
and U6558 (N_6558,N_4306,N_4676);
nand U6559 (N_6559,N_4464,N_5191);
nor U6560 (N_6560,N_5785,N_4118);
xnor U6561 (N_6561,N_5967,N_4470);
nor U6562 (N_6562,N_4838,N_4973);
or U6563 (N_6563,N_4237,N_4911);
nand U6564 (N_6564,N_4065,N_4298);
and U6565 (N_6565,N_4707,N_5527);
and U6566 (N_6566,N_5665,N_5913);
nand U6567 (N_6567,N_5034,N_4501);
and U6568 (N_6568,N_4474,N_5091);
and U6569 (N_6569,N_5818,N_5486);
or U6570 (N_6570,N_5409,N_4799);
nand U6571 (N_6571,N_4776,N_4394);
nor U6572 (N_6572,N_5859,N_5772);
and U6573 (N_6573,N_5986,N_5905);
nand U6574 (N_6574,N_5105,N_4090);
nand U6575 (N_6575,N_4432,N_4740);
and U6576 (N_6576,N_5277,N_5805);
nor U6577 (N_6577,N_4876,N_4143);
nor U6578 (N_6578,N_4291,N_5397);
and U6579 (N_6579,N_5574,N_4948);
and U6580 (N_6580,N_5192,N_4046);
nor U6581 (N_6581,N_4634,N_4181);
nand U6582 (N_6582,N_5994,N_4735);
or U6583 (N_6583,N_5011,N_4086);
and U6584 (N_6584,N_5578,N_4571);
nor U6585 (N_6585,N_4929,N_5046);
nand U6586 (N_6586,N_5714,N_5330);
nand U6587 (N_6587,N_4112,N_4041);
nand U6588 (N_6588,N_5154,N_5840);
or U6589 (N_6589,N_5633,N_5901);
nand U6590 (N_6590,N_5515,N_5139);
nand U6591 (N_6591,N_5103,N_5613);
nand U6592 (N_6592,N_4974,N_5570);
nor U6593 (N_6593,N_5957,N_5843);
nor U6594 (N_6594,N_5099,N_5318);
and U6595 (N_6595,N_5983,N_5487);
nand U6596 (N_6596,N_4162,N_5002);
or U6597 (N_6597,N_5256,N_4195);
or U6598 (N_6598,N_5512,N_4439);
nor U6599 (N_6599,N_5732,N_5477);
nand U6600 (N_6600,N_4460,N_4324);
or U6601 (N_6601,N_5750,N_4951);
nand U6602 (N_6602,N_5583,N_5264);
and U6603 (N_6603,N_4515,N_4286);
nor U6604 (N_6604,N_4621,N_5384);
nand U6605 (N_6605,N_4108,N_5311);
nand U6606 (N_6606,N_5211,N_4274);
nor U6607 (N_6607,N_4303,N_4101);
and U6608 (N_6608,N_4009,N_5121);
or U6609 (N_6609,N_5372,N_5605);
and U6610 (N_6610,N_5464,N_4650);
nand U6611 (N_6611,N_5278,N_5440);
or U6612 (N_6612,N_4759,N_5973);
or U6613 (N_6613,N_4430,N_4514);
nor U6614 (N_6614,N_5721,N_5910);
or U6615 (N_6615,N_4604,N_5010);
nand U6616 (N_6616,N_5093,N_4867);
xor U6617 (N_6617,N_4545,N_5628);
and U6618 (N_6618,N_4133,N_4602);
and U6619 (N_6619,N_5551,N_5205);
and U6620 (N_6620,N_4503,N_4132);
nand U6621 (N_6621,N_4665,N_4222);
nand U6622 (N_6622,N_5361,N_4331);
and U6623 (N_6623,N_5228,N_5426);
nand U6624 (N_6624,N_4618,N_4754);
nand U6625 (N_6625,N_5544,N_5642);
or U6626 (N_6626,N_4843,N_4279);
nand U6627 (N_6627,N_5394,N_4586);
nor U6628 (N_6628,N_5111,N_5458);
nand U6629 (N_6629,N_5874,N_5352);
or U6630 (N_6630,N_5511,N_4229);
or U6631 (N_6631,N_4729,N_4272);
nor U6632 (N_6632,N_5457,N_4425);
and U6633 (N_6633,N_5287,N_5016);
xor U6634 (N_6634,N_5952,N_5731);
nand U6635 (N_6635,N_5048,N_5203);
or U6636 (N_6636,N_4617,N_5786);
and U6637 (N_6637,N_4804,N_5168);
or U6638 (N_6638,N_5706,N_5213);
and U6639 (N_6639,N_5304,N_5282);
nand U6640 (N_6640,N_4629,N_4536);
nand U6641 (N_6641,N_4635,N_5402);
nand U6642 (N_6642,N_5789,N_4442);
and U6643 (N_6643,N_5710,N_5170);
or U6644 (N_6644,N_5632,N_5399);
or U6645 (N_6645,N_4979,N_4398);
nor U6646 (N_6646,N_4020,N_5123);
or U6647 (N_6647,N_4188,N_4767);
nor U6648 (N_6648,N_5087,N_5819);
nand U6649 (N_6649,N_4163,N_4669);
nor U6650 (N_6650,N_5500,N_4992);
or U6651 (N_6651,N_5044,N_5338);
nand U6652 (N_6652,N_5738,N_4956);
nor U6653 (N_6653,N_5420,N_5163);
nand U6654 (N_6654,N_4580,N_4659);
nor U6655 (N_6655,N_5450,N_5915);
or U6656 (N_6656,N_4393,N_5408);
and U6657 (N_6657,N_5796,N_4649);
nand U6658 (N_6658,N_5118,N_5018);
or U6659 (N_6659,N_5995,N_5070);
nor U6660 (N_6660,N_5636,N_5023);
nand U6661 (N_6661,N_5871,N_4013);
nor U6662 (N_6662,N_4354,N_4685);
or U6663 (N_6663,N_5508,N_4283);
xor U6664 (N_6664,N_5685,N_5239);
or U6665 (N_6665,N_5857,N_5396);
and U6666 (N_6666,N_5323,N_4748);
nor U6667 (N_6667,N_5977,N_4762);
or U6668 (N_6668,N_4869,N_5683);
nand U6669 (N_6669,N_4152,N_5742);
or U6670 (N_6670,N_4147,N_5561);
nand U6671 (N_6671,N_5055,N_4520);
nand U6672 (N_6672,N_5592,N_5243);
nor U6673 (N_6673,N_4842,N_4371);
nand U6674 (N_6674,N_5652,N_4054);
xor U6675 (N_6675,N_4214,N_5602);
or U6676 (N_6676,N_5342,N_5280);
or U6677 (N_6677,N_4630,N_4980);
nand U6678 (N_6678,N_5929,N_4313);
or U6679 (N_6679,N_5190,N_4037);
nor U6680 (N_6680,N_5573,N_5884);
nand U6681 (N_6681,N_4745,N_5907);
xor U6682 (N_6682,N_4409,N_5172);
and U6683 (N_6683,N_5242,N_5908);
nor U6684 (N_6684,N_5678,N_4436);
nor U6685 (N_6685,N_5313,N_5124);
or U6686 (N_6686,N_4482,N_4562);
nor U6687 (N_6687,N_5787,N_5556);
nand U6688 (N_6688,N_4523,N_5493);
nor U6689 (N_6689,N_5435,N_5656);
or U6690 (N_6690,N_4610,N_5265);
nor U6691 (N_6691,N_5870,N_4926);
nor U6692 (N_6692,N_4734,N_4265);
nand U6693 (N_6693,N_4356,N_4879);
and U6694 (N_6694,N_4531,N_4644);
xnor U6695 (N_6695,N_4600,N_4835);
nand U6696 (N_6696,N_4881,N_4778);
and U6697 (N_6697,N_4756,N_4719);
nor U6698 (N_6698,N_4420,N_4652);
nand U6699 (N_6699,N_5897,N_4431);
nand U6700 (N_6700,N_5883,N_5185);
nor U6701 (N_6701,N_5108,N_4005);
or U6702 (N_6702,N_5183,N_4458);
and U6703 (N_6703,N_5784,N_4396);
nand U6704 (N_6704,N_4763,N_4372);
and U6705 (N_6705,N_4557,N_5658);
nor U6706 (N_6706,N_4616,N_5505);
or U6707 (N_6707,N_5850,N_4750);
nor U6708 (N_6708,N_5591,N_5392);
or U6709 (N_6709,N_4284,N_4484);
nor U6710 (N_6710,N_4175,N_4382);
nor U6711 (N_6711,N_5383,N_4192);
and U6712 (N_6712,N_4322,N_5122);
nor U6713 (N_6713,N_4049,N_4378);
and U6714 (N_6714,N_4700,N_5483);
or U6715 (N_6715,N_4045,N_5984);
nor U6716 (N_6716,N_4151,N_5790);
or U6717 (N_6717,N_4877,N_4136);
xor U6718 (N_6718,N_4301,N_4696);
nand U6719 (N_6719,N_5369,N_5523);
nand U6720 (N_6720,N_5474,N_5865);
nand U6721 (N_6721,N_5807,N_5581);
nor U6722 (N_6722,N_4144,N_5363);
nor U6723 (N_6723,N_5063,N_5166);
nor U6724 (N_6724,N_4025,N_5717);
nand U6725 (N_6725,N_5137,N_4724);
xor U6726 (N_6726,N_5199,N_5261);
nand U6727 (N_6727,N_5360,N_5698);
or U6728 (N_6728,N_5425,N_4727);
nand U6729 (N_6729,N_4836,N_5600);
nor U6730 (N_6730,N_5775,N_4390);
xor U6731 (N_6731,N_4399,N_5467);
or U6732 (N_6732,N_4316,N_5494);
or U6733 (N_6733,N_5881,N_4860);
or U6734 (N_6734,N_5940,N_5832);
nor U6735 (N_6735,N_5196,N_4113);
and U6736 (N_6736,N_4070,N_4582);
or U6737 (N_6737,N_4653,N_4088);
or U6738 (N_6738,N_5267,N_4185);
nor U6739 (N_6739,N_4347,N_4747);
nand U6740 (N_6740,N_4801,N_4853);
and U6741 (N_6741,N_4252,N_4549);
nor U6742 (N_6742,N_5169,N_5547);
or U6743 (N_6743,N_4285,N_5290);
nor U6744 (N_6744,N_5616,N_4454);
nand U6745 (N_6745,N_4073,N_5734);
xor U6746 (N_6746,N_4190,N_4577);
and U6747 (N_6747,N_4114,N_5681);
nor U6748 (N_6748,N_5647,N_5896);
nand U6749 (N_6749,N_4493,N_4532);
and U6750 (N_6750,N_5575,N_4139);
and U6751 (N_6751,N_4288,N_4829);
nand U6752 (N_6752,N_4537,N_4350);
or U6753 (N_6753,N_5532,N_5990);
nand U6754 (N_6754,N_5562,N_5218);
nor U6755 (N_6755,N_4384,N_4846);
xnor U6756 (N_6756,N_5235,N_4731);
or U6757 (N_6757,N_4738,N_5453);
nand U6758 (N_6758,N_4670,N_5284);
nor U6759 (N_6759,N_5157,N_4456);
or U6760 (N_6760,N_5941,N_4681);
nor U6761 (N_6761,N_5935,N_4675);
or U6762 (N_6762,N_5669,N_4230);
xor U6763 (N_6763,N_5366,N_5869);
or U6764 (N_6764,N_5922,N_4744);
or U6765 (N_6765,N_5988,N_4245);
and U6766 (N_6766,N_5125,N_5674);
xnor U6767 (N_6767,N_5295,N_4546);
nor U6768 (N_6768,N_4165,N_5074);
or U6769 (N_6769,N_4965,N_4256);
and U6770 (N_6770,N_5297,N_4868);
nand U6771 (N_6771,N_5451,N_4094);
nand U6772 (N_6772,N_4140,N_5175);
or U6773 (N_6773,N_5607,N_4716);
nand U6774 (N_6774,N_4593,N_4507);
nand U6775 (N_6775,N_4097,N_4189);
and U6776 (N_6776,N_5623,N_4235);
and U6777 (N_6777,N_5699,N_4831);
nand U6778 (N_6778,N_4596,N_5931);
nand U6779 (N_6779,N_4446,N_4766);
and U6780 (N_6780,N_4872,N_5723);
nor U6781 (N_6781,N_5322,N_5165);
and U6782 (N_6782,N_4106,N_5852);
and U6783 (N_6783,N_4368,N_4646);
or U6784 (N_6784,N_4047,N_5410);
or U6785 (N_6785,N_4000,N_4925);
or U6786 (N_6786,N_5621,N_5694);
nand U6787 (N_6787,N_4952,N_4310);
or U6788 (N_6788,N_4148,N_4319);
xor U6789 (N_6789,N_5773,N_5934);
nand U6790 (N_6790,N_4161,N_4352);
nand U6791 (N_6791,N_4661,N_5333);
or U6792 (N_6792,N_4010,N_5933);
nor U6793 (N_6793,N_5129,N_5209);
nor U6794 (N_6794,N_5813,N_5873);
or U6795 (N_6795,N_5204,N_4107);
nand U6796 (N_6796,N_5682,N_4930);
and U6797 (N_6797,N_5753,N_4036);
and U6798 (N_6798,N_4558,N_5376);
and U6799 (N_6799,N_5824,N_4255);
nand U6800 (N_6800,N_4761,N_5001);
and U6801 (N_6801,N_5641,N_4708);
or U6802 (N_6802,N_4852,N_4341);
nor U6803 (N_6803,N_4982,N_5331);
xor U6804 (N_6804,N_5113,N_5022);
and U6805 (N_6805,N_4408,N_5400);
nand U6806 (N_6806,N_5148,N_4299);
and U6807 (N_6807,N_5872,N_5153);
nand U6808 (N_6808,N_5882,N_5920);
nor U6809 (N_6809,N_5076,N_4187);
or U6810 (N_6810,N_4769,N_5312);
and U6811 (N_6811,N_5851,N_4338);
nor U6812 (N_6812,N_4223,N_4891);
or U6813 (N_6813,N_5546,N_5339);
nor U6814 (N_6814,N_4295,N_4312);
xor U6815 (N_6815,N_4936,N_5405);
nor U6816 (N_6816,N_4606,N_4366);
or U6817 (N_6817,N_5663,N_5822);
nor U6818 (N_6818,N_4603,N_4395);
and U6819 (N_6819,N_4405,N_4450);
nand U6820 (N_6820,N_5437,N_4785);
and U6821 (N_6821,N_5079,N_5064);
and U6822 (N_6822,N_4894,N_5735);
and U6823 (N_6823,N_4183,N_5071);
and U6824 (N_6824,N_4579,N_4346);
nor U6825 (N_6825,N_4098,N_5622);
nor U6826 (N_6826,N_4240,N_5187);
or U6827 (N_6827,N_4030,N_4228);
nor U6828 (N_6828,N_5433,N_4817);
and U6829 (N_6829,N_5729,N_5746);
xor U6830 (N_6830,N_4943,N_5759);
and U6831 (N_6831,N_4794,N_5436);
nand U6832 (N_6832,N_5171,N_5285);
nor U6833 (N_6833,N_4569,N_5980);
xor U6834 (N_6834,N_5069,N_4589);
and U6835 (N_6835,N_4017,N_4448);
and U6836 (N_6836,N_4145,N_5927);
and U6837 (N_6837,N_5839,N_5444);
or U6838 (N_6838,N_5912,N_5268);
nor U6839 (N_6839,N_5823,N_5745);
or U6840 (N_6840,N_4224,N_5364);
or U6841 (N_6841,N_4239,N_4839);
or U6842 (N_6842,N_5593,N_4715);
nor U6843 (N_6843,N_5468,N_5567);
or U6844 (N_6844,N_5020,N_4379);
and U6845 (N_6845,N_5130,N_5349);
and U6846 (N_6846,N_5829,N_5764);
and U6847 (N_6847,N_5572,N_5599);
and U6848 (N_6848,N_4004,N_5117);
nor U6849 (N_6849,N_4225,N_4984);
and U6850 (N_6850,N_4595,N_4429);
and U6851 (N_6851,N_4142,N_5814);
or U6852 (N_6852,N_4664,N_5432);
nor U6853 (N_6853,N_4819,N_4056);
and U6854 (N_6854,N_4667,N_4300);
and U6855 (N_6855,N_5089,N_5793);
nor U6856 (N_6856,N_4281,N_4695);
and U6857 (N_6857,N_5082,N_4697);
nor U6858 (N_6858,N_4495,N_4855);
nand U6859 (N_6859,N_4788,N_4909);
nor U6860 (N_6860,N_5899,N_5906);
or U6861 (N_6861,N_5692,N_5132);
nor U6862 (N_6862,N_4568,N_4633);
or U6863 (N_6863,N_5576,N_4457);
nor U6864 (N_6864,N_4824,N_4972);
or U6865 (N_6865,N_5354,N_4494);
nand U6866 (N_6866,N_4931,N_5558);
and U6867 (N_6867,N_4802,N_5837);
or U6868 (N_6868,N_4720,N_5248);
and U6869 (N_6869,N_5077,N_5788);
or U6870 (N_6870,N_4924,N_5351);
nand U6871 (N_6871,N_5162,N_5164);
or U6872 (N_6872,N_4850,N_5144);
or U6873 (N_6873,N_4848,N_4174);
and U6874 (N_6874,N_5258,N_4679);
or U6875 (N_6875,N_5862,N_5629);
or U6876 (N_6876,N_4598,N_5180);
nand U6877 (N_6877,N_5895,N_4896);
nand U6878 (N_6878,N_4387,N_4035);
xor U6879 (N_6879,N_4023,N_4249);
and U6880 (N_6880,N_4805,N_5702);
and U6881 (N_6881,N_4317,N_4033);
nor U6882 (N_6882,N_4120,N_5606);
or U6883 (N_6883,N_4320,N_4611);
and U6884 (N_6884,N_4340,N_5382);
and U6885 (N_6885,N_4977,N_5803);
and U6886 (N_6886,N_5758,N_4613);
or U6887 (N_6887,N_4922,N_5447);
and U6888 (N_6888,N_4566,N_4849);
nor U6889 (N_6889,N_5680,N_5442);
xnor U6890 (N_6890,N_5589,N_4104);
or U6891 (N_6891,N_5693,N_5090);
or U6892 (N_6892,N_5058,N_5801);
nor U6893 (N_6893,N_4219,N_5926);
nand U6894 (N_6894,N_4538,N_4007);
nand U6895 (N_6895,N_5848,N_4332);
xor U6896 (N_6896,N_5095,N_4597);
and U6897 (N_6897,N_4483,N_5007);
nor U6898 (N_6898,N_4158,N_5098);
nor U6899 (N_6899,N_5497,N_5353);
nand U6900 (N_6900,N_5727,N_5878);
nand U6901 (N_6901,N_4585,N_5008);
nand U6902 (N_6902,N_5465,N_4803);
nand U6903 (N_6903,N_5045,N_5953);
or U6904 (N_6904,N_5513,N_4622);
or U6905 (N_6905,N_4064,N_5003);
or U6906 (N_6906,N_4180,N_5147);
and U6907 (N_6907,N_4651,N_5969);
nor U6908 (N_6908,N_4220,N_5325);
and U6909 (N_6909,N_5643,N_4958);
and U6910 (N_6910,N_4570,N_4775);
nor U6911 (N_6911,N_4957,N_4003);
or U6912 (N_6912,N_5345,N_5503);
nor U6913 (N_6913,N_4050,N_4642);
or U6914 (N_6914,N_5834,N_5017);
nor U6915 (N_6915,N_4199,N_4827);
and U6916 (N_6916,N_4736,N_4205);
or U6917 (N_6917,N_5292,N_5012);
and U6918 (N_6918,N_4278,N_4587);
and U6919 (N_6919,N_5231,N_4326);
nor U6920 (N_6920,N_5886,N_4806);
and U6921 (N_6921,N_4987,N_5156);
nand U6922 (N_6922,N_4920,N_5923);
nor U6923 (N_6923,N_5799,N_4043);
and U6924 (N_6924,N_5854,N_5482);
xor U6925 (N_6925,N_5189,N_4530);
nor U6926 (N_6926,N_4814,N_5612);
nor U6927 (N_6927,N_5577,N_4584);
nor U6928 (N_6928,N_4290,N_4122);
or U6929 (N_6929,N_4683,N_5999);
and U6930 (N_6930,N_5057,N_5521);
nand U6931 (N_6931,N_4656,N_4076);
and U6932 (N_6932,N_4961,N_5481);
nand U6933 (N_6933,N_4563,N_5653);
or U6934 (N_6934,N_5956,N_5150);
or U6935 (N_6935,N_5944,N_5251);
or U6936 (N_6936,N_5340,N_4155);
and U6937 (N_6937,N_4994,N_5202);
and U6938 (N_6938,N_4491,N_4212);
nand U6939 (N_6939,N_5075,N_4941);
nand U6940 (N_6940,N_4357,N_5719);
or U6941 (N_6941,N_5035,N_5293);
nor U6942 (N_6942,N_5741,N_5260);
nor U6943 (N_6943,N_5557,N_4213);
or U6944 (N_6944,N_5026,N_5904);
nor U6945 (N_6945,N_5780,N_5930);
nand U6946 (N_6946,N_4703,N_5845);
or U6947 (N_6947,N_5550,N_5271);
xnor U6948 (N_6948,N_4392,N_4502);
and U6949 (N_6949,N_4308,N_5625);
or U6950 (N_6950,N_4072,N_4385);
or U6951 (N_6951,N_5955,N_5703);
or U6952 (N_6952,N_4878,N_4699);
nand U6953 (N_6953,N_5092,N_4123);
or U6954 (N_6954,N_5013,N_4833);
and U6955 (N_6955,N_4781,N_4856);
or U6956 (N_6956,N_5049,N_5524);
nor U6957 (N_6957,N_5428,N_4455);
nand U6958 (N_6958,N_5946,N_4510);
nor U6959 (N_6959,N_4115,N_5604);
nand U6960 (N_6960,N_4263,N_4782);
nand U6961 (N_6961,N_5582,N_4820);
nor U6962 (N_6962,N_4441,N_4737);
nor U6963 (N_6963,N_4361,N_4678);
and U6964 (N_6964,N_5368,N_5212);
and U6965 (N_6965,N_5078,N_5229);
or U6966 (N_6966,N_5982,N_5120);
or U6967 (N_6967,N_4950,N_5649);
or U6968 (N_6968,N_5736,N_4764);
or U6969 (N_6969,N_4816,N_4910);
xor U6970 (N_6970,N_5533,N_4771);
nand U6971 (N_6971,N_4296,N_4257);
nor U6972 (N_6972,N_5097,N_5536);
nor U6973 (N_6973,N_5580,N_5174);
nand U6974 (N_6974,N_5668,N_5554);
nor U6975 (N_6975,N_5549,N_4791);
nand U6976 (N_6976,N_5176,N_4565);
nand U6977 (N_6977,N_4476,N_4682);
and U6978 (N_6978,N_5569,N_4937);
nor U6979 (N_6979,N_4938,N_4620);
nor U6980 (N_6980,N_5177,N_4404);
and U6981 (N_6981,N_4847,N_5028);
and U6982 (N_6982,N_5516,N_4928);
nor U6983 (N_6983,N_5724,N_5237);
nand U6984 (N_6984,N_5377,N_4414);
nor U6985 (N_6985,N_4250,N_4270);
or U6986 (N_6986,N_4753,N_4564);
nand U6987 (N_6987,N_4693,N_5958);
nor U6988 (N_6988,N_5520,N_4712);
or U6989 (N_6989,N_4059,N_5065);
xor U6990 (N_6990,N_4818,N_4717);
or U6991 (N_6991,N_5236,N_5317);
nand U6992 (N_6992,N_4907,N_4590);
nor U6993 (N_6993,N_5835,N_4694);
or U6994 (N_6994,N_4091,N_4654);
nand U6995 (N_6995,N_4077,N_4210);
nor U6996 (N_6996,N_5109,N_4471);
nor U6997 (N_6997,N_4089,N_4837);
nand U6998 (N_6998,N_5755,N_4193);
nor U6999 (N_6999,N_5259,N_4857);
nor U7000 (N_7000,N_4542,N_5860);
and U7001 (N_7001,N_5036,N_5659);
or U7002 (N_7002,N_5730,N_4347);
nor U7003 (N_7003,N_5265,N_4872);
or U7004 (N_7004,N_5837,N_4671);
nor U7005 (N_7005,N_5149,N_5029);
nor U7006 (N_7006,N_5581,N_4614);
or U7007 (N_7007,N_4871,N_5669);
nand U7008 (N_7008,N_4354,N_4716);
and U7009 (N_7009,N_5607,N_4016);
nand U7010 (N_7010,N_4826,N_4151);
and U7011 (N_7011,N_4518,N_4833);
or U7012 (N_7012,N_5535,N_5523);
nand U7013 (N_7013,N_5786,N_4359);
and U7014 (N_7014,N_4954,N_4168);
and U7015 (N_7015,N_5734,N_5554);
or U7016 (N_7016,N_4360,N_5551);
or U7017 (N_7017,N_5156,N_4289);
nand U7018 (N_7018,N_5022,N_4114);
nor U7019 (N_7019,N_5193,N_5982);
or U7020 (N_7020,N_5586,N_4346);
and U7021 (N_7021,N_5034,N_5772);
or U7022 (N_7022,N_5255,N_4948);
nor U7023 (N_7023,N_4054,N_5717);
nand U7024 (N_7024,N_4859,N_4566);
and U7025 (N_7025,N_4120,N_4851);
nand U7026 (N_7026,N_5472,N_4853);
nor U7027 (N_7027,N_4352,N_4857);
and U7028 (N_7028,N_4367,N_5492);
nor U7029 (N_7029,N_4552,N_5032);
or U7030 (N_7030,N_5148,N_5447);
and U7031 (N_7031,N_5691,N_5822);
or U7032 (N_7032,N_4011,N_5953);
nor U7033 (N_7033,N_4759,N_4998);
and U7034 (N_7034,N_4818,N_5774);
nor U7035 (N_7035,N_5282,N_4137);
nand U7036 (N_7036,N_5213,N_4891);
nor U7037 (N_7037,N_4417,N_4304);
nor U7038 (N_7038,N_4754,N_5293);
or U7039 (N_7039,N_5131,N_5560);
or U7040 (N_7040,N_4821,N_4436);
nor U7041 (N_7041,N_5982,N_4370);
or U7042 (N_7042,N_5327,N_5132);
or U7043 (N_7043,N_5336,N_4395);
xor U7044 (N_7044,N_5104,N_4534);
nor U7045 (N_7045,N_5770,N_4942);
or U7046 (N_7046,N_4679,N_4114);
nor U7047 (N_7047,N_4067,N_4242);
and U7048 (N_7048,N_5174,N_5900);
or U7049 (N_7049,N_5798,N_4520);
nor U7050 (N_7050,N_5904,N_5223);
nor U7051 (N_7051,N_4703,N_5075);
nand U7052 (N_7052,N_5616,N_5311);
or U7053 (N_7053,N_4458,N_4229);
or U7054 (N_7054,N_5989,N_4538);
or U7055 (N_7055,N_5524,N_4569);
nor U7056 (N_7056,N_4206,N_5372);
nand U7057 (N_7057,N_4278,N_4193);
nand U7058 (N_7058,N_5972,N_5278);
or U7059 (N_7059,N_5819,N_4699);
or U7060 (N_7060,N_5133,N_5974);
nor U7061 (N_7061,N_5476,N_5004);
nor U7062 (N_7062,N_4502,N_4010);
nand U7063 (N_7063,N_4617,N_5873);
and U7064 (N_7064,N_5601,N_4322);
nor U7065 (N_7065,N_4504,N_4387);
and U7066 (N_7066,N_5029,N_5242);
and U7067 (N_7067,N_5047,N_5056);
and U7068 (N_7068,N_4447,N_4575);
and U7069 (N_7069,N_5564,N_4133);
and U7070 (N_7070,N_5753,N_4096);
and U7071 (N_7071,N_5680,N_5877);
nor U7072 (N_7072,N_5229,N_5084);
nand U7073 (N_7073,N_4084,N_5910);
nand U7074 (N_7074,N_5386,N_5714);
and U7075 (N_7075,N_4428,N_4156);
xnor U7076 (N_7076,N_5082,N_4838);
nand U7077 (N_7077,N_5707,N_5087);
or U7078 (N_7078,N_4899,N_5494);
nand U7079 (N_7079,N_5252,N_4332);
nor U7080 (N_7080,N_5159,N_5088);
or U7081 (N_7081,N_4114,N_4699);
and U7082 (N_7082,N_5851,N_4474);
nand U7083 (N_7083,N_5868,N_4052);
or U7084 (N_7084,N_5303,N_4379);
nand U7085 (N_7085,N_5955,N_5023);
xor U7086 (N_7086,N_5088,N_4759);
nor U7087 (N_7087,N_4666,N_4824);
or U7088 (N_7088,N_4779,N_5381);
or U7089 (N_7089,N_5122,N_5737);
nor U7090 (N_7090,N_5920,N_4572);
nor U7091 (N_7091,N_4530,N_4532);
nor U7092 (N_7092,N_4690,N_5065);
nand U7093 (N_7093,N_5547,N_4369);
nand U7094 (N_7094,N_4960,N_5993);
or U7095 (N_7095,N_5195,N_4258);
and U7096 (N_7096,N_5929,N_4286);
or U7097 (N_7097,N_5369,N_4357);
and U7098 (N_7098,N_5135,N_4922);
nand U7099 (N_7099,N_5529,N_4916);
and U7100 (N_7100,N_4283,N_4428);
or U7101 (N_7101,N_4388,N_4191);
xnor U7102 (N_7102,N_4270,N_5760);
nand U7103 (N_7103,N_5312,N_5582);
and U7104 (N_7104,N_4839,N_4632);
and U7105 (N_7105,N_5457,N_4718);
nand U7106 (N_7106,N_5233,N_4084);
nand U7107 (N_7107,N_5624,N_4038);
nor U7108 (N_7108,N_5441,N_4951);
nor U7109 (N_7109,N_5044,N_5586);
nand U7110 (N_7110,N_5602,N_5620);
nand U7111 (N_7111,N_5227,N_5460);
nor U7112 (N_7112,N_5721,N_4695);
nor U7113 (N_7113,N_4317,N_4809);
nor U7114 (N_7114,N_5174,N_4319);
and U7115 (N_7115,N_4424,N_5415);
or U7116 (N_7116,N_5507,N_5252);
nand U7117 (N_7117,N_5507,N_5980);
and U7118 (N_7118,N_4869,N_4432);
or U7119 (N_7119,N_4830,N_4338);
nand U7120 (N_7120,N_4559,N_4937);
nor U7121 (N_7121,N_4803,N_4331);
and U7122 (N_7122,N_5203,N_5305);
or U7123 (N_7123,N_4246,N_4686);
nor U7124 (N_7124,N_4998,N_5484);
and U7125 (N_7125,N_4041,N_5172);
nor U7126 (N_7126,N_4786,N_4156);
or U7127 (N_7127,N_4292,N_4464);
nand U7128 (N_7128,N_4461,N_5819);
nor U7129 (N_7129,N_4040,N_5633);
and U7130 (N_7130,N_5856,N_4913);
and U7131 (N_7131,N_4535,N_5668);
nor U7132 (N_7132,N_4176,N_5853);
or U7133 (N_7133,N_4817,N_4535);
and U7134 (N_7134,N_5130,N_5764);
nand U7135 (N_7135,N_4554,N_5849);
or U7136 (N_7136,N_4470,N_4317);
or U7137 (N_7137,N_5750,N_5385);
nand U7138 (N_7138,N_4143,N_4287);
nor U7139 (N_7139,N_5211,N_5461);
or U7140 (N_7140,N_5053,N_5830);
nand U7141 (N_7141,N_4212,N_4650);
nand U7142 (N_7142,N_4025,N_4453);
and U7143 (N_7143,N_4873,N_4428);
or U7144 (N_7144,N_4603,N_4621);
nand U7145 (N_7145,N_4807,N_4274);
nand U7146 (N_7146,N_4954,N_5062);
nand U7147 (N_7147,N_4789,N_5733);
nand U7148 (N_7148,N_4310,N_5288);
nor U7149 (N_7149,N_5712,N_4488);
nand U7150 (N_7150,N_5583,N_5017);
nand U7151 (N_7151,N_4523,N_5705);
nor U7152 (N_7152,N_5546,N_4728);
nor U7153 (N_7153,N_4314,N_4438);
nand U7154 (N_7154,N_4260,N_4223);
xnor U7155 (N_7155,N_4948,N_5040);
nor U7156 (N_7156,N_4781,N_5675);
nor U7157 (N_7157,N_4578,N_5243);
and U7158 (N_7158,N_5358,N_4036);
or U7159 (N_7159,N_5231,N_4232);
nand U7160 (N_7160,N_5817,N_4900);
nor U7161 (N_7161,N_4800,N_4345);
and U7162 (N_7162,N_4483,N_4540);
and U7163 (N_7163,N_5935,N_5473);
or U7164 (N_7164,N_5096,N_4947);
nand U7165 (N_7165,N_4032,N_5318);
and U7166 (N_7166,N_4485,N_4670);
nor U7167 (N_7167,N_5794,N_5360);
nand U7168 (N_7168,N_5899,N_4941);
and U7169 (N_7169,N_5999,N_4953);
nand U7170 (N_7170,N_4792,N_5553);
nor U7171 (N_7171,N_4245,N_4447);
nand U7172 (N_7172,N_5825,N_4527);
or U7173 (N_7173,N_4911,N_5532);
and U7174 (N_7174,N_4168,N_5541);
nand U7175 (N_7175,N_5400,N_4463);
nor U7176 (N_7176,N_5911,N_4280);
nor U7177 (N_7177,N_4555,N_4220);
and U7178 (N_7178,N_5621,N_5296);
or U7179 (N_7179,N_4891,N_5567);
nor U7180 (N_7180,N_5303,N_4313);
and U7181 (N_7181,N_4737,N_5689);
nor U7182 (N_7182,N_4914,N_4673);
and U7183 (N_7183,N_5886,N_5997);
nor U7184 (N_7184,N_4109,N_4977);
and U7185 (N_7185,N_5798,N_4975);
and U7186 (N_7186,N_5863,N_4114);
or U7187 (N_7187,N_5590,N_4866);
nand U7188 (N_7188,N_5988,N_4803);
nor U7189 (N_7189,N_5731,N_5798);
and U7190 (N_7190,N_5604,N_5433);
nand U7191 (N_7191,N_5614,N_5704);
or U7192 (N_7192,N_5753,N_4199);
or U7193 (N_7193,N_5841,N_4889);
nor U7194 (N_7194,N_4137,N_5359);
nor U7195 (N_7195,N_5984,N_5998);
and U7196 (N_7196,N_5085,N_4270);
nor U7197 (N_7197,N_5221,N_4029);
and U7198 (N_7198,N_5665,N_4995);
nor U7199 (N_7199,N_5063,N_4207);
or U7200 (N_7200,N_5210,N_4471);
nor U7201 (N_7201,N_4555,N_5319);
and U7202 (N_7202,N_5416,N_5593);
and U7203 (N_7203,N_4955,N_5161);
xnor U7204 (N_7204,N_4959,N_4236);
nor U7205 (N_7205,N_5298,N_5009);
nor U7206 (N_7206,N_4682,N_5246);
or U7207 (N_7207,N_4405,N_4878);
nor U7208 (N_7208,N_4573,N_5732);
or U7209 (N_7209,N_4388,N_5698);
or U7210 (N_7210,N_5955,N_5941);
nand U7211 (N_7211,N_5250,N_4522);
or U7212 (N_7212,N_4799,N_4609);
nor U7213 (N_7213,N_4082,N_5713);
nand U7214 (N_7214,N_4094,N_5767);
or U7215 (N_7215,N_4738,N_5333);
or U7216 (N_7216,N_5400,N_4718);
or U7217 (N_7217,N_5800,N_4648);
or U7218 (N_7218,N_5056,N_5644);
nor U7219 (N_7219,N_5858,N_5097);
and U7220 (N_7220,N_4892,N_5189);
nor U7221 (N_7221,N_5538,N_5416);
or U7222 (N_7222,N_5060,N_5659);
or U7223 (N_7223,N_5144,N_5540);
nor U7224 (N_7224,N_5233,N_5072);
and U7225 (N_7225,N_5685,N_4700);
xnor U7226 (N_7226,N_4318,N_5655);
nand U7227 (N_7227,N_5069,N_5750);
nand U7228 (N_7228,N_4822,N_4882);
nor U7229 (N_7229,N_4356,N_4268);
or U7230 (N_7230,N_4028,N_4763);
nand U7231 (N_7231,N_5104,N_4028);
or U7232 (N_7232,N_5948,N_5003);
and U7233 (N_7233,N_4378,N_5080);
nor U7234 (N_7234,N_5723,N_5799);
or U7235 (N_7235,N_4877,N_5333);
or U7236 (N_7236,N_5986,N_4766);
nor U7237 (N_7237,N_4444,N_5249);
or U7238 (N_7238,N_4038,N_5739);
or U7239 (N_7239,N_4655,N_4380);
nand U7240 (N_7240,N_5462,N_5571);
nand U7241 (N_7241,N_4290,N_4857);
nand U7242 (N_7242,N_4946,N_4604);
and U7243 (N_7243,N_5123,N_5450);
or U7244 (N_7244,N_5154,N_4282);
nor U7245 (N_7245,N_4721,N_5826);
nor U7246 (N_7246,N_4840,N_4209);
and U7247 (N_7247,N_5639,N_4694);
and U7248 (N_7248,N_4680,N_4285);
nand U7249 (N_7249,N_4984,N_4917);
nand U7250 (N_7250,N_5742,N_5870);
or U7251 (N_7251,N_5708,N_4460);
nand U7252 (N_7252,N_4491,N_5501);
nor U7253 (N_7253,N_4198,N_5670);
nor U7254 (N_7254,N_4449,N_4401);
and U7255 (N_7255,N_4516,N_4062);
or U7256 (N_7256,N_5707,N_5900);
nand U7257 (N_7257,N_5481,N_5433);
or U7258 (N_7258,N_4926,N_4149);
nand U7259 (N_7259,N_5454,N_5075);
or U7260 (N_7260,N_5305,N_4786);
nand U7261 (N_7261,N_5224,N_5124);
and U7262 (N_7262,N_5436,N_4371);
nor U7263 (N_7263,N_5125,N_5943);
or U7264 (N_7264,N_5620,N_4802);
nor U7265 (N_7265,N_4466,N_4144);
nor U7266 (N_7266,N_5907,N_5529);
and U7267 (N_7267,N_5125,N_4801);
and U7268 (N_7268,N_4487,N_5839);
and U7269 (N_7269,N_4998,N_5424);
nand U7270 (N_7270,N_4010,N_5687);
xnor U7271 (N_7271,N_5999,N_4131);
xor U7272 (N_7272,N_4711,N_4903);
nor U7273 (N_7273,N_4168,N_5674);
or U7274 (N_7274,N_5522,N_4869);
or U7275 (N_7275,N_4256,N_5723);
or U7276 (N_7276,N_4390,N_5615);
nand U7277 (N_7277,N_4198,N_4315);
nand U7278 (N_7278,N_5953,N_5368);
nand U7279 (N_7279,N_5768,N_5077);
nor U7280 (N_7280,N_4121,N_5410);
nand U7281 (N_7281,N_5780,N_5570);
and U7282 (N_7282,N_4893,N_4208);
and U7283 (N_7283,N_4025,N_5989);
nand U7284 (N_7284,N_5351,N_4420);
or U7285 (N_7285,N_4429,N_5257);
and U7286 (N_7286,N_4641,N_4170);
and U7287 (N_7287,N_4197,N_5639);
nor U7288 (N_7288,N_4436,N_4666);
nand U7289 (N_7289,N_4782,N_4869);
or U7290 (N_7290,N_5087,N_4791);
nor U7291 (N_7291,N_4582,N_5525);
and U7292 (N_7292,N_4011,N_5107);
nor U7293 (N_7293,N_5902,N_5812);
nor U7294 (N_7294,N_4636,N_5505);
nor U7295 (N_7295,N_4619,N_4029);
or U7296 (N_7296,N_4604,N_5863);
nand U7297 (N_7297,N_4820,N_5954);
and U7298 (N_7298,N_4994,N_4371);
or U7299 (N_7299,N_5085,N_5956);
nand U7300 (N_7300,N_5144,N_5272);
and U7301 (N_7301,N_5690,N_5872);
and U7302 (N_7302,N_4612,N_4469);
or U7303 (N_7303,N_4239,N_4278);
or U7304 (N_7304,N_5347,N_4034);
nand U7305 (N_7305,N_5799,N_5853);
or U7306 (N_7306,N_5050,N_4072);
or U7307 (N_7307,N_5175,N_4970);
or U7308 (N_7308,N_4750,N_5992);
and U7309 (N_7309,N_5768,N_5050);
or U7310 (N_7310,N_5185,N_4489);
nor U7311 (N_7311,N_4782,N_4653);
and U7312 (N_7312,N_4706,N_4918);
nand U7313 (N_7313,N_5463,N_4890);
nand U7314 (N_7314,N_5255,N_4179);
or U7315 (N_7315,N_4366,N_4368);
and U7316 (N_7316,N_4233,N_4353);
and U7317 (N_7317,N_4264,N_4304);
or U7318 (N_7318,N_4751,N_5052);
and U7319 (N_7319,N_4128,N_5409);
or U7320 (N_7320,N_4824,N_4336);
nand U7321 (N_7321,N_4530,N_4222);
nand U7322 (N_7322,N_4033,N_5750);
nor U7323 (N_7323,N_4923,N_4145);
and U7324 (N_7324,N_4229,N_4144);
nor U7325 (N_7325,N_5462,N_5782);
or U7326 (N_7326,N_4780,N_5569);
or U7327 (N_7327,N_5569,N_5329);
and U7328 (N_7328,N_4581,N_5090);
or U7329 (N_7329,N_4228,N_4539);
nor U7330 (N_7330,N_5200,N_4829);
nor U7331 (N_7331,N_5357,N_5630);
and U7332 (N_7332,N_5346,N_5728);
nand U7333 (N_7333,N_4370,N_4121);
or U7334 (N_7334,N_4437,N_4663);
and U7335 (N_7335,N_4631,N_5102);
and U7336 (N_7336,N_4649,N_4019);
nor U7337 (N_7337,N_5840,N_5196);
xor U7338 (N_7338,N_5304,N_5414);
nand U7339 (N_7339,N_4108,N_4918);
nand U7340 (N_7340,N_4475,N_5281);
nand U7341 (N_7341,N_4612,N_4934);
and U7342 (N_7342,N_5002,N_5181);
or U7343 (N_7343,N_5675,N_5508);
and U7344 (N_7344,N_4719,N_5162);
nand U7345 (N_7345,N_4320,N_5070);
nand U7346 (N_7346,N_5936,N_4094);
and U7347 (N_7347,N_5449,N_5314);
nor U7348 (N_7348,N_4741,N_4955);
nor U7349 (N_7349,N_5208,N_5319);
nand U7350 (N_7350,N_4435,N_5045);
and U7351 (N_7351,N_5191,N_5480);
nor U7352 (N_7352,N_4918,N_5205);
and U7353 (N_7353,N_4022,N_5111);
and U7354 (N_7354,N_4214,N_5497);
xor U7355 (N_7355,N_4648,N_5719);
or U7356 (N_7356,N_4244,N_5355);
nand U7357 (N_7357,N_5208,N_5267);
and U7358 (N_7358,N_4182,N_5043);
nand U7359 (N_7359,N_4422,N_4380);
nor U7360 (N_7360,N_4230,N_4120);
and U7361 (N_7361,N_4106,N_4104);
or U7362 (N_7362,N_5689,N_4070);
nand U7363 (N_7363,N_4212,N_4293);
nand U7364 (N_7364,N_5303,N_4734);
nand U7365 (N_7365,N_5534,N_4804);
or U7366 (N_7366,N_5291,N_5456);
nor U7367 (N_7367,N_5126,N_4424);
and U7368 (N_7368,N_5656,N_5282);
nor U7369 (N_7369,N_4146,N_4513);
nand U7370 (N_7370,N_5118,N_5612);
or U7371 (N_7371,N_5378,N_5555);
nor U7372 (N_7372,N_4539,N_5539);
or U7373 (N_7373,N_4420,N_4448);
nand U7374 (N_7374,N_4034,N_5972);
xor U7375 (N_7375,N_4927,N_5387);
nand U7376 (N_7376,N_5638,N_4743);
nor U7377 (N_7377,N_4968,N_4113);
nand U7378 (N_7378,N_4029,N_5474);
and U7379 (N_7379,N_5087,N_4275);
nand U7380 (N_7380,N_5956,N_5399);
nand U7381 (N_7381,N_4805,N_4872);
nor U7382 (N_7382,N_5466,N_4498);
nor U7383 (N_7383,N_4763,N_5256);
and U7384 (N_7384,N_5627,N_5216);
or U7385 (N_7385,N_4651,N_4096);
or U7386 (N_7386,N_5110,N_5345);
nand U7387 (N_7387,N_5381,N_5246);
or U7388 (N_7388,N_5647,N_4443);
nand U7389 (N_7389,N_4128,N_4184);
and U7390 (N_7390,N_5729,N_4046);
and U7391 (N_7391,N_4105,N_5653);
nand U7392 (N_7392,N_4263,N_4726);
nor U7393 (N_7393,N_5166,N_5195);
and U7394 (N_7394,N_5456,N_5866);
nand U7395 (N_7395,N_5879,N_5474);
or U7396 (N_7396,N_4480,N_4508);
nor U7397 (N_7397,N_5575,N_4420);
nand U7398 (N_7398,N_4153,N_5415);
nor U7399 (N_7399,N_4917,N_5484);
nor U7400 (N_7400,N_5084,N_5331);
nand U7401 (N_7401,N_4238,N_4039);
and U7402 (N_7402,N_5043,N_5898);
nor U7403 (N_7403,N_4795,N_5421);
or U7404 (N_7404,N_5082,N_5222);
nor U7405 (N_7405,N_5823,N_5310);
nand U7406 (N_7406,N_4291,N_4310);
or U7407 (N_7407,N_5350,N_5061);
and U7408 (N_7408,N_5418,N_5106);
and U7409 (N_7409,N_5583,N_5330);
nand U7410 (N_7410,N_4520,N_4150);
nand U7411 (N_7411,N_4877,N_4437);
and U7412 (N_7412,N_5746,N_4145);
nor U7413 (N_7413,N_4329,N_5408);
or U7414 (N_7414,N_5172,N_5532);
xor U7415 (N_7415,N_4638,N_4873);
or U7416 (N_7416,N_5000,N_4469);
or U7417 (N_7417,N_5750,N_4446);
nand U7418 (N_7418,N_4717,N_4366);
or U7419 (N_7419,N_5151,N_5687);
nor U7420 (N_7420,N_4119,N_4712);
and U7421 (N_7421,N_5135,N_4463);
and U7422 (N_7422,N_4558,N_5284);
or U7423 (N_7423,N_5789,N_4700);
nor U7424 (N_7424,N_5674,N_5273);
nor U7425 (N_7425,N_5321,N_5581);
and U7426 (N_7426,N_4215,N_4893);
nor U7427 (N_7427,N_4085,N_4324);
nand U7428 (N_7428,N_4898,N_5273);
xor U7429 (N_7429,N_4455,N_5980);
nand U7430 (N_7430,N_4617,N_5121);
or U7431 (N_7431,N_4354,N_5314);
nor U7432 (N_7432,N_4505,N_5689);
and U7433 (N_7433,N_4843,N_4832);
nor U7434 (N_7434,N_5565,N_5276);
or U7435 (N_7435,N_4682,N_5213);
and U7436 (N_7436,N_4149,N_5741);
or U7437 (N_7437,N_4927,N_4058);
or U7438 (N_7438,N_4682,N_5270);
nor U7439 (N_7439,N_5614,N_4893);
or U7440 (N_7440,N_5425,N_5062);
xnor U7441 (N_7441,N_4885,N_5200);
or U7442 (N_7442,N_4923,N_4705);
or U7443 (N_7443,N_4159,N_4838);
and U7444 (N_7444,N_4968,N_5675);
nand U7445 (N_7445,N_5573,N_4958);
and U7446 (N_7446,N_5470,N_4079);
and U7447 (N_7447,N_4056,N_5919);
or U7448 (N_7448,N_5320,N_4155);
and U7449 (N_7449,N_5801,N_4781);
nor U7450 (N_7450,N_5864,N_5930);
and U7451 (N_7451,N_4095,N_5683);
nand U7452 (N_7452,N_5750,N_5569);
nand U7453 (N_7453,N_4019,N_4313);
nor U7454 (N_7454,N_5510,N_5956);
nand U7455 (N_7455,N_5952,N_4950);
nand U7456 (N_7456,N_5148,N_4234);
or U7457 (N_7457,N_5501,N_5650);
nand U7458 (N_7458,N_4543,N_5892);
and U7459 (N_7459,N_5658,N_5872);
nand U7460 (N_7460,N_4431,N_5508);
and U7461 (N_7461,N_4689,N_5865);
nor U7462 (N_7462,N_5343,N_4156);
xnor U7463 (N_7463,N_5923,N_5580);
or U7464 (N_7464,N_5371,N_5658);
or U7465 (N_7465,N_5089,N_5490);
nand U7466 (N_7466,N_5369,N_4064);
nand U7467 (N_7467,N_4583,N_4525);
nor U7468 (N_7468,N_4742,N_5306);
nand U7469 (N_7469,N_4028,N_5760);
or U7470 (N_7470,N_4010,N_4324);
nand U7471 (N_7471,N_5063,N_4131);
nor U7472 (N_7472,N_5298,N_4935);
nand U7473 (N_7473,N_4386,N_4579);
or U7474 (N_7474,N_5427,N_4134);
nand U7475 (N_7475,N_5493,N_4458);
and U7476 (N_7476,N_4874,N_4280);
nor U7477 (N_7477,N_4267,N_5723);
or U7478 (N_7478,N_4172,N_5639);
nand U7479 (N_7479,N_4897,N_4800);
and U7480 (N_7480,N_4294,N_4396);
and U7481 (N_7481,N_4047,N_4490);
nand U7482 (N_7482,N_5776,N_5327);
nor U7483 (N_7483,N_4454,N_5225);
or U7484 (N_7484,N_5289,N_4972);
and U7485 (N_7485,N_4722,N_4561);
and U7486 (N_7486,N_5339,N_4008);
and U7487 (N_7487,N_4359,N_4629);
or U7488 (N_7488,N_4261,N_4738);
nor U7489 (N_7489,N_5374,N_5403);
or U7490 (N_7490,N_5343,N_5387);
and U7491 (N_7491,N_5877,N_4414);
nand U7492 (N_7492,N_4872,N_5963);
nor U7493 (N_7493,N_4130,N_5156);
and U7494 (N_7494,N_5978,N_4455);
and U7495 (N_7495,N_5421,N_4950);
nor U7496 (N_7496,N_5087,N_5046);
or U7497 (N_7497,N_4484,N_4247);
and U7498 (N_7498,N_5387,N_4509);
and U7499 (N_7499,N_4467,N_4209);
nand U7500 (N_7500,N_4428,N_4180);
or U7501 (N_7501,N_4882,N_5683);
xnor U7502 (N_7502,N_5711,N_5900);
nand U7503 (N_7503,N_5687,N_5943);
and U7504 (N_7504,N_4282,N_4541);
and U7505 (N_7505,N_4400,N_5214);
xnor U7506 (N_7506,N_4073,N_5844);
and U7507 (N_7507,N_5697,N_4428);
or U7508 (N_7508,N_4513,N_5877);
and U7509 (N_7509,N_5436,N_4000);
nand U7510 (N_7510,N_5915,N_5369);
or U7511 (N_7511,N_4403,N_4519);
or U7512 (N_7512,N_5618,N_4340);
nor U7513 (N_7513,N_5168,N_5087);
and U7514 (N_7514,N_4443,N_4619);
nand U7515 (N_7515,N_4470,N_4159);
or U7516 (N_7516,N_5409,N_5784);
nand U7517 (N_7517,N_4317,N_4406);
or U7518 (N_7518,N_4288,N_5662);
and U7519 (N_7519,N_4931,N_4343);
or U7520 (N_7520,N_4684,N_5927);
or U7521 (N_7521,N_4207,N_4875);
or U7522 (N_7522,N_4517,N_4574);
or U7523 (N_7523,N_5643,N_5327);
and U7524 (N_7524,N_4652,N_4016);
nor U7525 (N_7525,N_5728,N_4023);
nand U7526 (N_7526,N_4142,N_5481);
or U7527 (N_7527,N_4668,N_5137);
or U7528 (N_7528,N_5785,N_5942);
nand U7529 (N_7529,N_4286,N_4992);
nand U7530 (N_7530,N_4018,N_5966);
or U7531 (N_7531,N_5503,N_4998);
nor U7532 (N_7532,N_5705,N_4153);
or U7533 (N_7533,N_5410,N_5646);
nand U7534 (N_7534,N_5620,N_4047);
xor U7535 (N_7535,N_5142,N_5217);
nor U7536 (N_7536,N_5259,N_4417);
or U7537 (N_7537,N_4060,N_5948);
nand U7538 (N_7538,N_5540,N_5809);
and U7539 (N_7539,N_4390,N_4744);
and U7540 (N_7540,N_4002,N_4069);
xnor U7541 (N_7541,N_4128,N_5120);
and U7542 (N_7542,N_5891,N_5824);
or U7543 (N_7543,N_4318,N_4681);
nor U7544 (N_7544,N_5507,N_4814);
and U7545 (N_7545,N_4871,N_4333);
or U7546 (N_7546,N_4196,N_4383);
nor U7547 (N_7547,N_4561,N_4541);
nand U7548 (N_7548,N_5520,N_4128);
nor U7549 (N_7549,N_5750,N_5460);
and U7550 (N_7550,N_4096,N_5530);
and U7551 (N_7551,N_5106,N_4962);
nor U7552 (N_7552,N_4908,N_4421);
or U7553 (N_7553,N_4638,N_4686);
and U7554 (N_7554,N_5403,N_5417);
nand U7555 (N_7555,N_5924,N_4127);
and U7556 (N_7556,N_4784,N_4113);
nand U7557 (N_7557,N_4668,N_4242);
nand U7558 (N_7558,N_5066,N_4054);
and U7559 (N_7559,N_5260,N_5825);
nor U7560 (N_7560,N_4687,N_5744);
nor U7561 (N_7561,N_5019,N_5913);
and U7562 (N_7562,N_5057,N_5787);
nor U7563 (N_7563,N_4857,N_5441);
or U7564 (N_7564,N_4567,N_4476);
or U7565 (N_7565,N_4426,N_5629);
nor U7566 (N_7566,N_5504,N_4865);
nand U7567 (N_7567,N_5802,N_5967);
nand U7568 (N_7568,N_4103,N_4533);
or U7569 (N_7569,N_5022,N_4333);
and U7570 (N_7570,N_5236,N_4269);
and U7571 (N_7571,N_4536,N_4154);
nand U7572 (N_7572,N_4772,N_4498);
and U7573 (N_7573,N_5570,N_5943);
nand U7574 (N_7574,N_5107,N_4897);
nor U7575 (N_7575,N_4097,N_4228);
nand U7576 (N_7576,N_4192,N_5693);
nor U7577 (N_7577,N_5600,N_4200);
and U7578 (N_7578,N_5413,N_4581);
and U7579 (N_7579,N_4217,N_5632);
and U7580 (N_7580,N_4156,N_5857);
nand U7581 (N_7581,N_5898,N_5842);
nor U7582 (N_7582,N_4428,N_5123);
nor U7583 (N_7583,N_5819,N_4412);
nand U7584 (N_7584,N_4700,N_5588);
or U7585 (N_7585,N_5047,N_5399);
nand U7586 (N_7586,N_4446,N_4311);
nor U7587 (N_7587,N_4760,N_5714);
nor U7588 (N_7588,N_4038,N_4183);
nor U7589 (N_7589,N_4617,N_5970);
nor U7590 (N_7590,N_5772,N_4477);
and U7591 (N_7591,N_4031,N_5825);
and U7592 (N_7592,N_4837,N_4928);
nand U7593 (N_7593,N_4579,N_5553);
or U7594 (N_7594,N_4627,N_5902);
nor U7595 (N_7595,N_5761,N_5308);
nor U7596 (N_7596,N_4388,N_5956);
and U7597 (N_7597,N_4175,N_4925);
or U7598 (N_7598,N_5584,N_5783);
nand U7599 (N_7599,N_4871,N_4659);
or U7600 (N_7600,N_5113,N_5544);
or U7601 (N_7601,N_4041,N_4463);
nor U7602 (N_7602,N_5842,N_5139);
nor U7603 (N_7603,N_4227,N_5604);
nand U7604 (N_7604,N_4906,N_5203);
nand U7605 (N_7605,N_4901,N_4534);
and U7606 (N_7606,N_5222,N_4979);
nand U7607 (N_7607,N_5676,N_5405);
or U7608 (N_7608,N_4819,N_4172);
nand U7609 (N_7609,N_5247,N_4952);
or U7610 (N_7610,N_5343,N_5258);
or U7611 (N_7611,N_4571,N_4755);
or U7612 (N_7612,N_4056,N_5509);
or U7613 (N_7613,N_5956,N_4464);
and U7614 (N_7614,N_5732,N_5284);
nor U7615 (N_7615,N_5647,N_5562);
nand U7616 (N_7616,N_5676,N_4878);
and U7617 (N_7617,N_5716,N_4073);
and U7618 (N_7618,N_4650,N_5124);
and U7619 (N_7619,N_4430,N_5671);
nand U7620 (N_7620,N_5340,N_4491);
and U7621 (N_7621,N_5972,N_4480);
nand U7622 (N_7622,N_4990,N_5349);
and U7623 (N_7623,N_5067,N_5756);
and U7624 (N_7624,N_5624,N_4184);
or U7625 (N_7625,N_4580,N_5047);
nand U7626 (N_7626,N_5901,N_5361);
and U7627 (N_7627,N_4432,N_4500);
nand U7628 (N_7628,N_4017,N_4525);
nand U7629 (N_7629,N_4080,N_4936);
and U7630 (N_7630,N_5200,N_4236);
nor U7631 (N_7631,N_4931,N_5697);
nand U7632 (N_7632,N_4328,N_4343);
xor U7633 (N_7633,N_5219,N_5111);
and U7634 (N_7634,N_5503,N_4310);
nor U7635 (N_7635,N_5699,N_5029);
or U7636 (N_7636,N_4833,N_5828);
and U7637 (N_7637,N_5554,N_5324);
or U7638 (N_7638,N_4427,N_5525);
or U7639 (N_7639,N_5219,N_4977);
or U7640 (N_7640,N_5314,N_4696);
and U7641 (N_7641,N_4240,N_5768);
or U7642 (N_7642,N_4332,N_5297);
and U7643 (N_7643,N_5145,N_4136);
or U7644 (N_7644,N_5234,N_4804);
nor U7645 (N_7645,N_4463,N_4771);
or U7646 (N_7646,N_5065,N_4636);
nand U7647 (N_7647,N_4800,N_5421);
or U7648 (N_7648,N_4107,N_5431);
nor U7649 (N_7649,N_4162,N_4308);
or U7650 (N_7650,N_5188,N_5319);
or U7651 (N_7651,N_4863,N_5640);
and U7652 (N_7652,N_5151,N_4141);
and U7653 (N_7653,N_4012,N_5632);
xor U7654 (N_7654,N_4159,N_4077);
and U7655 (N_7655,N_4043,N_4637);
nor U7656 (N_7656,N_4064,N_4275);
or U7657 (N_7657,N_4573,N_5835);
and U7658 (N_7658,N_5985,N_4379);
and U7659 (N_7659,N_4742,N_5151);
nand U7660 (N_7660,N_4470,N_5223);
nand U7661 (N_7661,N_4150,N_5172);
and U7662 (N_7662,N_5479,N_5592);
and U7663 (N_7663,N_4656,N_5595);
and U7664 (N_7664,N_5380,N_5489);
nor U7665 (N_7665,N_5148,N_5503);
and U7666 (N_7666,N_5371,N_5076);
nor U7667 (N_7667,N_5626,N_4698);
and U7668 (N_7668,N_5107,N_5532);
nand U7669 (N_7669,N_5507,N_4711);
and U7670 (N_7670,N_4543,N_5338);
and U7671 (N_7671,N_4411,N_5592);
or U7672 (N_7672,N_5455,N_4580);
and U7673 (N_7673,N_5558,N_5165);
nand U7674 (N_7674,N_5952,N_4854);
nor U7675 (N_7675,N_4201,N_4228);
nor U7676 (N_7676,N_4727,N_5055);
nor U7677 (N_7677,N_4049,N_4624);
or U7678 (N_7678,N_4539,N_4400);
and U7679 (N_7679,N_4481,N_4574);
and U7680 (N_7680,N_5336,N_4292);
nand U7681 (N_7681,N_5031,N_5785);
nand U7682 (N_7682,N_4391,N_4343);
and U7683 (N_7683,N_5568,N_4056);
nand U7684 (N_7684,N_4721,N_4813);
nand U7685 (N_7685,N_4823,N_4339);
or U7686 (N_7686,N_5077,N_4177);
nor U7687 (N_7687,N_4268,N_5233);
nor U7688 (N_7688,N_5600,N_5537);
or U7689 (N_7689,N_4946,N_5331);
nor U7690 (N_7690,N_5487,N_5328);
or U7691 (N_7691,N_5488,N_5481);
or U7692 (N_7692,N_5243,N_5289);
and U7693 (N_7693,N_4738,N_4307);
and U7694 (N_7694,N_5487,N_4505);
or U7695 (N_7695,N_4503,N_4588);
nor U7696 (N_7696,N_4250,N_5170);
and U7697 (N_7697,N_4664,N_5529);
nor U7698 (N_7698,N_5428,N_5197);
nor U7699 (N_7699,N_4756,N_5654);
nor U7700 (N_7700,N_5589,N_4556);
and U7701 (N_7701,N_4255,N_4481);
and U7702 (N_7702,N_4375,N_4390);
nor U7703 (N_7703,N_5886,N_5079);
and U7704 (N_7704,N_5567,N_5548);
and U7705 (N_7705,N_5179,N_4448);
nand U7706 (N_7706,N_4405,N_5347);
nand U7707 (N_7707,N_5914,N_4640);
nor U7708 (N_7708,N_4157,N_4852);
nor U7709 (N_7709,N_5300,N_4668);
or U7710 (N_7710,N_4485,N_5137);
nand U7711 (N_7711,N_5186,N_5641);
nand U7712 (N_7712,N_4352,N_4268);
nand U7713 (N_7713,N_4991,N_5185);
nor U7714 (N_7714,N_5591,N_4379);
or U7715 (N_7715,N_5038,N_4098);
and U7716 (N_7716,N_4929,N_4445);
nor U7717 (N_7717,N_4123,N_4878);
or U7718 (N_7718,N_5399,N_4897);
and U7719 (N_7719,N_5847,N_5608);
and U7720 (N_7720,N_5592,N_5623);
nand U7721 (N_7721,N_4170,N_4744);
and U7722 (N_7722,N_4433,N_4362);
or U7723 (N_7723,N_5321,N_5361);
nor U7724 (N_7724,N_4898,N_5058);
nand U7725 (N_7725,N_4306,N_5374);
or U7726 (N_7726,N_4753,N_5639);
nand U7727 (N_7727,N_5603,N_5532);
nand U7728 (N_7728,N_4335,N_4887);
nor U7729 (N_7729,N_4731,N_5676);
and U7730 (N_7730,N_4846,N_4745);
nor U7731 (N_7731,N_4064,N_4173);
nor U7732 (N_7732,N_4644,N_5440);
and U7733 (N_7733,N_5655,N_5373);
and U7734 (N_7734,N_5876,N_4675);
or U7735 (N_7735,N_5440,N_5685);
nand U7736 (N_7736,N_5659,N_4655);
or U7737 (N_7737,N_5592,N_5869);
nor U7738 (N_7738,N_4106,N_4888);
or U7739 (N_7739,N_4422,N_5575);
or U7740 (N_7740,N_5858,N_5297);
nand U7741 (N_7741,N_4075,N_4127);
nand U7742 (N_7742,N_4682,N_5193);
and U7743 (N_7743,N_4819,N_4243);
or U7744 (N_7744,N_5390,N_4598);
nor U7745 (N_7745,N_4205,N_5873);
nand U7746 (N_7746,N_5214,N_4988);
nor U7747 (N_7747,N_5084,N_4397);
or U7748 (N_7748,N_5860,N_5934);
and U7749 (N_7749,N_5992,N_5416);
or U7750 (N_7750,N_5919,N_5528);
or U7751 (N_7751,N_4053,N_5179);
and U7752 (N_7752,N_4954,N_4072);
nand U7753 (N_7753,N_4464,N_5886);
nand U7754 (N_7754,N_5674,N_5951);
or U7755 (N_7755,N_4856,N_5293);
and U7756 (N_7756,N_5384,N_5160);
or U7757 (N_7757,N_5585,N_4095);
or U7758 (N_7758,N_4295,N_5517);
nor U7759 (N_7759,N_5746,N_5768);
nand U7760 (N_7760,N_5747,N_5247);
nor U7761 (N_7761,N_5754,N_5942);
nand U7762 (N_7762,N_4285,N_4693);
nand U7763 (N_7763,N_5159,N_5956);
nand U7764 (N_7764,N_4399,N_4897);
or U7765 (N_7765,N_4410,N_5536);
nand U7766 (N_7766,N_5239,N_4633);
or U7767 (N_7767,N_5109,N_4428);
nor U7768 (N_7768,N_4780,N_5107);
and U7769 (N_7769,N_5140,N_4465);
or U7770 (N_7770,N_5408,N_4729);
or U7771 (N_7771,N_5783,N_5149);
nand U7772 (N_7772,N_5786,N_4645);
and U7773 (N_7773,N_5734,N_5331);
and U7774 (N_7774,N_5561,N_5724);
xnor U7775 (N_7775,N_5393,N_5723);
nor U7776 (N_7776,N_4034,N_5537);
nor U7777 (N_7777,N_5509,N_5499);
and U7778 (N_7778,N_5463,N_4838);
xnor U7779 (N_7779,N_4989,N_4897);
nor U7780 (N_7780,N_4261,N_4418);
nand U7781 (N_7781,N_5802,N_4652);
xor U7782 (N_7782,N_5145,N_4989);
nand U7783 (N_7783,N_4941,N_4218);
or U7784 (N_7784,N_5245,N_5526);
or U7785 (N_7785,N_5780,N_5174);
and U7786 (N_7786,N_4987,N_4179);
nand U7787 (N_7787,N_4609,N_5015);
and U7788 (N_7788,N_4580,N_4113);
and U7789 (N_7789,N_5753,N_5867);
or U7790 (N_7790,N_4289,N_4727);
or U7791 (N_7791,N_5464,N_5986);
and U7792 (N_7792,N_5368,N_5829);
nand U7793 (N_7793,N_4714,N_5527);
and U7794 (N_7794,N_4484,N_4108);
and U7795 (N_7795,N_4778,N_4571);
nor U7796 (N_7796,N_4115,N_4950);
nand U7797 (N_7797,N_5275,N_4482);
or U7798 (N_7798,N_5250,N_5894);
nor U7799 (N_7799,N_4018,N_5636);
and U7800 (N_7800,N_4240,N_4612);
or U7801 (N_7801,N_5547,N_5571);
nand U7802 (N_7802,N_5201,N_4091);
nand U7803 (N_7803,N_4362,N_4650);
and U7804 (N_7804,N_4027,N_4666);
nor U7805 (N_7805,N_4358,N_5673);
and U7806 (N_7806,N_4762,N_5932);
and U7807 (N_7807,N_5886,N_4776);
and U7808 (N_7808,N_4997,N_4276);
nand U7809 (N_7809,N_5526,N_5355);
and U7810 (N_7810,N_5847,N_4329);
or U7811 (N_7811,N_5494,N_4972);
nor U7812 (N_7812,N_4780,N_5053);
nor U7813 (N_7813,N_4908,N_5019);
nor U7814 (N_7814,N_4931,N_5626);
nor U7815 (N_7815,N_5613,N_5844);
or U7816 (N_7816,N_5714,N_4753);
or U7817 (N_7817,N_5205,N_4243);
nand U7818 (N_7818,N_5414,N_4112);
nand U7819 (N_7819,N_4934,N_5125);
nand U7820 (N_7820,N_4841,N_5106);
or U7821 (N_7821,N_4151,N_4571);
nand U7822 (N_7822,N_5336,N_4563);
nor U7823 (N_7823,N_5043,N_5155);
nand U7824 (N_7824,N_4785,N_5491);
and U7825 (N_7825,N_4790,N_4176);
nand U7826 (N_7826,N_4004,N_5159);
and U7827 (N_7827,N_4162,N_4820);
nand U7828 (N_7828,N_4143,N_4092);
nor U7829 (N_7829,N_4456,N_5036);
xor U7830 (N_7830,N_4422,N_5907);
nor U7831 (N_7831,N_4133,N_5723);
or U7832 (N_7832,N_5561,N_4449);
nor U7833 (N_7833,N_4082,N_5163);
nor U7834 (N_7834,N_4378,N_5671);
and U7835 (N_7835,N_5334,N_5252);
nor U7836 (N_7836,N_4271,N_4925);
or U7837 (N_7837,N_5777,N_4888);
and U7838 (N_7838,N_4691,N_5094);
nor U7839 (N_7839,N_4476,N_4989);
nand U7840 (N_7840,N_4195,N_5806);
and U7841 (N_7841,N_5367,N_5528);
nand U7842 (N_7842,N_4328,N_4351);
nor U7843 (N_7843,N_5352,N_4421);
nand U7844 (N_7844,N_4209,N_4038);
nand U7845 (N_7845,N_4315,N_5836);
or U7846 (N_7846,N_5989,N_5240);
and U7847 (N_7847,N_5650,N_4725);
and U7848 (N_7848,N_5088,N_5373);
or U7849 (N_7849,N_4102,N_4609);
nand U7850 (N_7850,N_5868,N_5192);
or U7851 (N_7851,N_5092,N_4038);
and U7852 (N_7852,N_4179,N_4891);
nor U7853 (N_7853,N_5378,N_4041);
nor U7854 (N_7854,N_4552,N_5362);
and U7855 (N_7855,N_5982,N_4026);
nor U7856 (N_7856,N_4219,N_4961);
nand U7857 (N_7857,N_5287,N_4640);
nor U7858 (N_7858,N_4253,N_5910);
nand U7859 (N_7859,N_5921,N_4195);
and U7860 (N_7860,N_4298,N_5913);
nor U7861 (N_7861,N_5624,N_4272);
nand U7862 (N_7862,N_4231,N_5348);
nor U7863 (N_7863,N_5501,N_5498);
nand U7864 (N_7864,N_5769,N_4865);
nand U7865 (N_7865,N_4423,N_4106);
or U7866 (N_7866,N_5549,N_4844);
and U7867 (N_7867,N_5880,N_5346);
and U7868 (N_7868,N_4317,N_5141);
and U7869 (N_7869,N_5323,N_5298);
and U7870 (N_7870,N_4149,N_5903);
or U7871 (N_7871,N_4333,N_4525);
or U7872 (N_7872,N_4717,N_4608);
and U7873 (N_7873,N_5934,N_5046);
nor U7874 (N_7874,N_4953,N_4310);
nand U7875 (N_7875,N_4051,N_5199);
and U7876 (N_7876,N_5959,N_5427);
nand U7877 (N_7877,N_5189,N_4555);
xor U7878 (N_7878,N_4201,N_4249);
nand U7879 (N_7879,N_4353,N_4947);
or U7880 (N_7880,N_5674,N_5300);
and U7881 (N_7881,N_4506,N_4125);
and U7882 (N_7882,N_4331,N_4829);
or U7883 (N_7883,N_5506,N_5181);
nand U7884 (N_7884,N_4277,N_5206);
nor U7885 (N_7885,N_4714,N_5883);
and U7886 (N_7886,N_4835,N_4848);
or U7887 (N_7887,N_5951,N_4858);
or U7888 (N_7888,N_5698,N_5681);
nand U7889 (N_7889,N_4577,N_5337);
and U7890 (N_7890,N_5902,N_5112);
nand U7891 (N_7891,N_4070,N_4000);
or U7892 (N_7892,N_4910,N_5867);
nor U7893 (N_7893,N_4130,N_4067);
and U7894 (N_7894,N_4959,N_5289);
or U7895 (N_7895,N_5529,N_4074);
nor U7896 (N_7896,N_5609,N_4390);
or U7897 (N_7897,N_4380,N_5519);
nand U7898 (N_7898,N_4878,N_5510);
nor U7899 (N_7899,N_4005,N_5189);
nand U7900 (N_7900,N_5487,N_5263);
nand U7901 (N_7901,N_5519,N_4357);
or U7902 (N_7902,N_4850,N_4294);
nand U7903 (N_7903,N_5921,N_5994);
and U7904 (N_7904,N_4300,N_4292);
nand U7905 (N_7905,N_5994,N_4785);
nor U7906 (N_7906,N_5282,N_5764);
nor U7907 (N_7907,N_4306,N_5180);
nand U7908 (N_7908,N_5424,N_4440);
and U7909 (N_7909,N_4951,N_4066);
nand U7910 (N_7910,N_4006,N_4572);
nor U7911 (N_7911,N_5581,N_5313);
nand U7912 (N_7912,N_5920,N_4740);
nand U7913 (N_7913,N_4064,N_4279);
nand U7914 (N_7914,N_5258,N_5028);
nand U7915 (N_7915,N_5861,N_5289);
and U7916 (N_7916,N_4281,N_4311);
nor U7917 (N_7917,N_5391,N_5562);
nand U7918 (N_7918,N_4192,N_4336);
nor U7919 (N_7919,N_5879,N_4774);
nand U7920 (N_7920,N_4822,N_4440);
nor U7921 (N_7921,N_4994,N_4367);
and U7922 (N_7922,N_4552,N_4141);
or U7923 (N_7923,N_5978,N_5599);
or U7924 (N_7924,N_5533,N_4169);
and U7925 (N_7925,N_5052,N_5129);
and U7926 (N_7926,N_5017,N_5882);
or U7927 (N_7927,N_4525,N_4109);
nand U7928 (N_7928,N_5850,N_4718);
or U7929 (N_7929,N_5757,N_5245);
nand U7930 (N_7930,N_4427,N_4123);
nand U7931 (N_7931,N_5367,N_5447);
nand U7932 (N_7932,N_5453,N_5520);
and U7933 (N_7933,N_4264,N_4145);
or U7934 (N_7934,N_4651,N_4401);
nor U7935 (N_7935,N_5944,N_5061);
and U7936 (N_7936,N_4275,N_4955);
and U7937 (N_7937,N_4159,N_4416);
and U7938 (N_7938,N_5820,N_4733);
or U7939 (N_7939,N_4927,N_4832);
nor U7940 (N_7940,N_5248,N_4005);
nand U7941 (N_7941,N_5894,N_4634);
nor U7942 (N_7942,N_5303,N_4941);
and U7943 (N_7943,N_5751,N_4362);
or U7944 (N_7944,N_4037,N_4640);
or U7945 (N_7945,N_5519,N_5806);
nor U7946 (N_7946,N_4297,N_4871);
and U7947 (N_7947,N_5239,N_5496);
nand U7948 (N_7948,N_5700,N_5696);
xnor U7949 (N_7949,N_4539,N_5215);
and U7950 (N_7950,N_5721,N_4013);
and U7951 (N_7951,N_4322,N_5793);
nor U7952 (N_7952,N_4069,N_5473);
and U7953 (N_7953,N_4249,N_4665);
nand U7954 (N_7954,N_4500,N_4023);
nand U7955 (N_7955,N_5304,N_4286);
nand U7956 (N_7956,N_5532,N_4555);
nand U7957 (N_7957,N_4651,N_4518);
nor U7958 (N_7958,N_4180,N_5126);
nand U7959 (N_7959,N_4607,N_5511);
nand U7960 (N_7960,N_4068,N_4387);
nor U7961 (N_7961,N_4480,N_4780);
and U7962 (N_7962,N_4647,N_4727);
nand U7963 (N_7963,N_5734,N_4184);
nand U7964 (N_7964,N_4452,N_4842);
and U7965 (N_7965,N_4333,N_4310);
and U7966 (N_7966,N_4233,N_4226);
nand U7967 (N_7967,N_4209,N_5742);
nand U7968 (N_7968,N_5248,N_4446);
or U7969 (N_7969,N_4814,N_4576);
and U7970 (N_7970,N_5762,N_5877);
and U7971 (N_7971,N_5957,N_4275);
nor U7972 (N_7972,N_4511,N_5999);
and U7973 (N_7973,N_4618,N_5116);
or U7974 (N_7974,N_5598,N_5074);
nand U7975 (N_7975,N_4673,N_5700);
and U7976 (N_7976,N_5557,N_4472);
and U7977 (N_7977,N_5058,N_5533);
and U7978 (N_7978,N_4810,N_4909);
nor U7979 (N_7979,N_5175,N_4573);
nor U7980 (N_7980,N_4464,N_4196);
or U7981 (N_7981,N_4002,N_4212);
or U7982 (N_7982,N_4528,N_4774);
xor U7983 (N_7983,N_5737,N_4860);
nand U7984 (N_7984,N_5265,N_4196);
and U7985 (N_7985,N_5603,N_4218);
nor U7986 (N_7986,N_4597,N_4992);
nand U7987 (N_7987,N_5331,N_4698);
nor U7988 (N_7988,N_5349,N_4420);
or U7989 (N_7989,N_5056,N_5901);
or U7990 (N_7990,N_5833,N_5652);
and U7991 (N_7991,N_5310,N_5664);
nand U7992 (N_7992,N_5804,N_5631);
and U7993 (N_7993,N_5363,N_4597);
or U7994 (N_7994,N_4039,N_4746);
and U7995 (N_7995,N_5642,N_4578);
nor U7996 (N_7996,N_4290,N_4728);
nor U7997 (N_7997,N_4933,N_5004);
or U7998 (N_7998,N_4157,N_5949);
and U7999 (N_7999,N_5005,N_4034);
nand U8000 (N_8000,N_7278,N_7810);
or U8001 (N_8001,N_6756,N_6576);
and U8002 (N_8002,N_6708,N_7713);
nand U8003 (N_8003,N_7426,N_6110);
nand U8004 (N_8004,N_6017,N_7799);
nand U8005 (N_8005,N_6952,N_7884);
and U8006 (N_8006,N_6285,N_7023);
or U8007 (N_8007,N_7806,N_6601);
and U8008 (N_8008,N_7195,N_6899);
and U8009 (N_8009,N_7314,N_7999);
and U8010 (N_8010,N_6956,N_6637);
nand U8011 (N_8011,N_6325,N_7991);
nand U8012 (N_8012,N_6830,N_6297);
nand U8013 (N_8013,N_6492,N_6578);
nand U8014 (N_8014,N_6726,N_7769);
nor U8015 (N_8015,N_6875,N_6214);
nor U8016 (N_8016,N_6998,N_6567);
or U8017 (N_8017,N_6200,N_6937);
and U8018 (N_8018,N_7581,N_7365);
or U8019 (N_8019,N_6840,N_6183);
or U8020 (N_8020,N_6903,N_7311);
nand U8021 (N_8021,N_6659,N_7431);
nand U8022 (N_8022,N_7688,N_7227);
or U8023 (N_8023,N_6364,N_7905);
xor U8024 (N_8024,N_6662,N_6494);
and U8025 (N_8025,N_6457,N_6163);
nor U8026 (N_8026,N_6877,N_7368);
xor U8027 (N_8027,N_6044,N_7469);
nand U8028 (N_8028,N_7893,N_6219);
nand U8029 (N_8029,N_7734,N_6078);
or U8030 (N_8030,N_6604,N_6119);
nor U8031 (N_8031,N_6700,N_7952);
or U8032 (N_8032,N_6283,N_7402);
nand U8033 (N_8033,N_6995,N_7282);
and U8034 (N_8034,N_7434,N_7464);
and U8035 (N_8035,N_7582,N_6780);
and U8036 (N_8036,N_7101,N_7720);
or U8037 (N_8037,N_7624,N_7946);
nor U8038 (N_8038,N_7290,N_7319);
nand U8039 (N_8039,N_6256,N_6721);
nor U8040 (N_8040,N_7505,N_6893);
or U8041 (N_8041,N_6684,N_6201);
nor U8042 (N_8042,N_7940,N_6921);
nand U8043 (N_8043,N_6501,N_6738);
or U8044 (N_8044,N_6591,N_6057);
or U8045 (N_8045,N_7007,N_6098);
and U8046 (N_8046,N_7403,N_6733);
nor U8047 (N_8047,N_7951,N_6159);
or U8048 (N_8048,N_6557,N_7941);
or U8049 (N_8049,N_6913,N_6933);
and U8050 (N_8050,N_7437,N_6254);
nor U8051 (N_8051,N_6841,N_6025);
nand U8052 (N_8052,N_7604,N_6021);
and U8053 (N_8053,N_7832,N_6340);
nand U8054 (N_8054,N_6130,N_7718);
or U8055 (N_8055,N_7309,N_6945);
or U8056 (N_8056,N_7163,N_6376);
nand U8057 (N_8057,N_7261,N_7771);
and U8058 (N_8058,N_7514,N_7153);
nor U8059 (N_8059,N_6408,N_7038);
nor U8060 (N_8060,N_6487,N_7009);
nand U8061 (N_8061,N_7215,N_7056);
nor U8062 (N_8062,N_6486,N_6282);
nand U8063 (N_8063,N_7093,N_7399);
and U8064 (N_8064,N_7149,N_7691);
nand U8065 (N_8065,N_6851,N_7800);
and U8066 (N_8066,N_6301,N_7229);
or U8067 (N_8067,N_6572,N_7871);
or U8068 (N_8068,N_6004,N_7166);
and U8069 (N_8069,N_6338,N_6895);
or U8070 (N_8070,N_6414,N_7144);
nand U8071 (N_8071,N_6737,N_7914);
nor U8072 (N_8072,N_6232,N_6676);
xnor U8073 (N_8073,N_6208,N_7306);
xnor U8074 (N_8074,N_7156,N_7566);
and U8075 (N_8075,N_6885,N_6826);
and U8076 (N_8076,N_6073,N_7934);
and U8077 (N_8077,N_6174,N_6905);
nand U8078 (N_8078,N_6904,N_6093);
or U8079 (N_8079,N_7356,N_6609);
and U8080 (N_8080,N_7367,N_6361);
nor U8081 (N_8081,N_7214,N_6446);
or U8082 (N_8082,N_7213,N_7533);
or U8083 (N_8083,N_6689,N_7335);
xnor U8084 (N_8084,N_7128,N_7879);
and U8085 (N_8085,N_7021,N_6982);
nand U8086 (N_8086,N_7135,N_7867);
and U8087 (N_8087,N_7292,N_6357);
nand U8088 (N_8088,N_7191,N_7202);
nor U8089 (N_8089,N_6918,N_7726);
nor U8090 (N_8090,N_7005,N_7266);
or U8091 (N_8091,N_7289,N_6648);
nand U8092 (N_8092,N_6991,N_7661);
and U8093 (N_8093,N_7658,N_7171);
and U8094 (N_8094,N_7079,N_6311);
nor U8095 (N_8095,N_6561,N_7666);
nor U8096 (N_8096,N_7897,N_6139);
and U8097 (N_8097,N_6362,N_7383);
nor U8098 (N_8098,N_6327,N_6673);
nor U8099 (N_8099,N_7498,N_7528);
nand U8100 (N_8100,N_6951,N_6696);
and U8101 (N_8101,N_6013,N_7092);
nor U8102 (N_8102,N_6041,N_7150);
or U8103 (N_8103,N_7842,N_7558);
or U8104 (N_8104,N_6805,N_7424);
or U8105 (N_8105,N_7578,N_7555);
nor U8106 (N_8106,N_7542,N_7413);
and U8107 (N_8107,N_7042,N_7181);
nor U8108 (N_8108,N_6321,N_7735);
or U8109 (N_8109,N_6770,N_7915);
xor U8110 (N_8110,N_6251,N_6079);
and U8111 (N_8111,N_7129,N_7053);
and U8112 (N_8112,N_7747,N_6072);
xnor U8113 (N_8113,N_6702,N_6538);
nor U8114 (N_8114,N_7669,N_6331);
or U8115 (N_8115,N_6483,N_7583);
or U8116 (N_8116,N_7158,N_7540);
or U8117 (N_8117,N_7616,N_6114);
nor U8118 (N_8118,N_7858,N_6391);
and U8119 (N_8119,N_6445,N_6644);
nor U8120 (N_8120,N_7516,N_7972);
and U8121 (N_8121,N_6916,N_7241);
and U8122 (N_8122,N_6766,N_7379);
and U8123 (N_8123,N_6817,N_7201);
nor U8124 (N_8124,N_7378,N_6108);
nand U8125 (N_8125,N_6687,N_6085);
nand U8126 (N_8126,N_7850,N_7955);
xnor U8127 (N_8127,N_6531,N_7126);
nor U8128 (N_8128,N_7255,N_7866);
nor U8129 (N_8129,N_6479,N_7446);
or U8130 (N_8130,N_7428,N_7878);
nor U8131 (N_8131,N_6053,N_7170);
nand U8132 (N_8132,N_7945,N_7554);
and U8133 (N_8133,N_7980,N_6943);
and U8134 (N_8134,N_6564,N_6158);
and U8135 (N_8135,N_7630,N_7580);
nand U8136 (N_8136,N_7244,N_7108);
nand U8137 (N_8137,N_6475,N_6808);
nor U8138 (N_8138,N_6882,N_6366);
nand U8139 (N_8139,N_6404,N_7541);
or U8140 (N_8140,N_6096,N_7325);
or U8141 (N_8141,N_6860,N_6758);
nor U8142 (N_8142,N_7793,N_7707);
nand U8143 (N_8143,N_6101,N_6190);
nor U8144 (N_8144,N_6415,N_7614);
or U8145 (N_8145,N_7141,N_7621);
and U8146 (N_8146,N_7326,N_6107);
nand U8147 (N_8147,N_7176,N_6465);
nand U8148 (N_8148,N_7697,N_7327);
or U8149 (N_8149,N_6188,N_7748);
or U8150 (N_8150,N_6223,N_6925);
nand U8151 (N_8151,N_6424,N_6771);
and U8152 (N_8152,N_7281,N_7853);
nor U8153 (N_8153,N_7313,N_7859);
nand U8154 (N_8154,N_7174,N_6761);
and U8155 (N_8155,N_7466,N_7393);
and U8156 (N_8156,N_7162,N_6339);
or U8157 (N_8157,N_6897,N_6596);
nor U8158 (N_8158,N_7308,N_6051);
or U8159 (N_8159,N_6599,N_6398);
nor U8160 (N_8160,N_6290,N_7118);
nor U8161 (N_8161,N_6575,N_6355);
nand U8162 (N_8162,N_7324,N_7104);
and U8163 (N_8163,N_6996,N_7245);
nor U8164 (N_8164,N_7569,N_7496);
nand U8165 (N_8165,N_7950,N_6498);
or U8166 (N_8166,N_7510,N_6109);
and U8167 (N_8167,N_6205,N_7018);
and U8168 (N_8168,N_6542,N_6461);
nor U8169 (N_8169,N_6224,N_6410);
xor U8170 (N_8170,N_6554,N_6822);
and U8171 (N_8171,N_6789,N_7632);
nand U8172 (N_8172,N_6328,N_7686);
or U8173 (N_8173,N_7740,N_6622);
and U8174 (N_8174,N_7277,N_6820);
nand U8175 (N_8175,N_7762,N_6587);
nand U8176 (N_8176,N_6309,N_6510);
nor U8177 (N_8177,N_6611,N_6835);
nand U8178 (N_8178,N_7962,N_7231);
xor U8179 (N_8179,N_7210,N_7273);
nor U8180 (N_8180,N_6195,N_6135);
and U8181 (N_8181,N_6832,N_7029);
and U8182 (N_8182,N_6682,N_7722);
and U8183 (N_8183,N_7636,N_6812);
and U8184 (N_8184,N_7060,N_7909);
nor U8185 (N_8185,N_7240,N_7727);
nand U8186 (N_8186,N_7550,N_6803);
nor U8187 (N_8187,N_7845,N_7435);
and U8188 (N_8188,N_7836,N_7396);
nor U8189 (N_8189,N_6735,N_7796);
nor U8190 (N_8190,N_6128,N_6022);
and U8191 (N_8191,N_7209,N_6981);
and U8192 (N_8192,N_6744,N_6975);
nand U8193 (N_8193,N_7138,N_6873);
or U8194 (N_8194,N_6102,N_6928);
or U8195 (N_8195,N_6675,N_7679);
nand U8196 (N_8196,N_6731,N_6047);
nor U8197 (N_8197,N_6762,N_7175);
or U8198 (N_8198,N_6798,N_7594);
and U8199 (N_8199,N_6718,N_6111);
or U8200 (N_8200,N_6967,N_7360);
nand U8201 (N_8201,N_6577,N_6674);
nand U8202 (N_8202,N_6693,N_7638);
and U8203 (N_8203,N_6631,N_6661);
and U8204 (N_8204,N_7287,N_6294);
and U8205 (N_8205,N_6570,N_6957);
or U8206 (N_8206,N_6252,N_6768);
nor U8207 (N_8207,N_6056,N_7130);
or U8208 (N_8208,N_6389,N_6630);
and U8209 (N_8209,N_7812,N_7818);
or U8210 (N_8210,N_6026,N_7398);
and U8211 (N_8211,N_6437,N_7072);
or U8212 (N_8212,N_7565,N_6330);
or U8213 (N_8213,N_6009,N_6239);
and U8214 (N_8214,N_6582,N_7530);
or U8215 (N_8215,N_6070,N_7220);
or U8216 (N_8216,N_6260,N_7139);
nand U8217 (N_8217,N_6180,N_7539);
or U8218 (N_8218,N_7095,N_7027);
nand U8219 (N_8219,N_7837,N_6350);
or U8220 (N_8220,N_6263,N_6528);
or U8221 (N_8221,N_7329,N_7640);
xnor U8222 (N_8222,N_7067,N_7116);
nor U8223 (N_8223,N_7825,N_7193);
or U8224 (N_8224,N_7113,N_6862);
and U8225 (N_8225,N_6354,N_6062);
and U8226 (N_8226,N_6192,N_7830);
and U8227 (N_8227,N_6767,N_7167);
nand U8228 (N_8228,N_7251,N_6865);
and U8229 (N_8229,N_7804,N_7271);
nor U8230 (N_8230,N_6211,N_6716);
and U8231 (N_8231,N_7136,N_7062);
and U8232 (N_8232,N_7462,N_7559);
nor U8233 (N_8233,N_6137,N_7807);
nor U8234 (N_8234,N_7047,N_7409);
nand U8235 (N_8235,N_6132,N_6908);
nor U8236 (N_8236,N_6887,N_6169);
and U8237 (N_8237,N_6750,N_6651);
and U8238 (N_8238,N_7288,N_6199);
and U8239 (N_8239,N_6417,N_7381);
or U8240 (N_8240,N_7698,N_7711);
or U8241 (N_8241,N_6255,N_7928);
and U8242 (N_8242,N_7607,N_6319);
nand U8243 (N_8243,N_6955,N_6462);
nor U8244 (N_8244,N_6593,N_7217);
and U8245 (N_8245,N_7664,N_7448);
nand U8246 (N_8246,N_7099,N_7506);
nor U8247 (N_8247,N_7598,N_6763);
or U8248 (N_8248,N_6329,N_6068);
nand U8249 (N_8249,N_7875,N_6580);
nor U8250 (N_8250,N_7061,N_6827);
and U8251 (N_8251,N_7743,N_7610);
nand U8252 (N_8252,N_7387,N_7082);
xor U8253 (N_8253,N_7772,N_6291);
or U8254 (N_8254,N_7423,N_7293);
and U8255 (N_8255,N_7562,N_7179);
nand U8256 (N_8256,N_7258,N_7328);
and U8257 (N_8257,N_6464,N_6246);
or U8258 (N_8258,N_6317,N_6560);
nor U8259 (N_8259,N_7133,N_6143);
nor U8260 (N_8260,N_7421,N_7246);
nand U8261 (N_8261,N_6390,N_7297);
xor U8262 (N_8262,N_7775,N_6506);
and U8263 (N_8263,N_6909,N_6295);
or U8264 (N_8264,N_7729,N_6603);
nand U8265 (N_8265,N_7236,N_6965);
nor U8266 (N_8266,N_7585,N_7809);
or U8267 (N_8267,N_7696,N_7532);
nand U8268 (N_8268,N_6852,N_6743);
and U8269 (N_8269,N_6799,N_6449);
and U8270 (N_8270,N_7186,N_6663);
and U8271 (N_8271,N_7519,N_6615);
nor U8272 (N_8272,N_6012,N_6490);
or U8273 (N_8273,N_6772,N_7194);
or U8274 (N_8274,N_7184,N_7567);
and U8275 (N_8275,N_6606,N_6588);
xnor U8276 (N_8276,N_6720,N_7545);
nor U8277 (N_8277,N_6058,N_6729);
and U8278 (N_8278,N_6162,N_6517);
and U8279 (N_8279,N_6476,N_7798);
or U8280 (N_8280,N_7451,N_7637);
or U8281 (N_8281,N_6455,N_7511);
and U8282 (N_8282,N_7020,N_6927);
nor U8283 (N_8283,N_6237,N_6172);
nand U8284 (N_8284,N_6342,N_7350);
or U8285 (N_8285,N_6828,N_6002);
nand U8286 (N_8286,N_7472,N_6382);
or U8287 (N_8287,N_7257,N_7123);
nand U8288 (N_8288,N_6848,N_7146);
and U8289 (N_8289,N_7786,N_7781);
nand U8290 (N_8290,N_7702,N_6221);
and U8291 (N_8291,N_7477,N_7492);
xnor U8292 (N_8292,N_7197,N_7612);
or U8293 (N_8293,N_6052,N_7015);
nor U8294 (N_8294,N_6837,N_7407);
and U8295 (N_8295,N_6749,N_7317);
nor U8296 (N_8296,N_6050,N_6715);
and U8297 (N_8297,N_6233,N_7342);
nand U8298 (N_8298,N_6960,N_6323);
nand U8299 (N_8299,N_7508,N_7779);
and U8300 (N_8300,N_7000,N_6258);
and U8301 (N_8301,N_7745,N_7183);
nand U8302 (N_8302,N_6787,N_6495);
and U8303 (N_8303,N_7004,N_6493);
and U8304 (N_8304,N_6405,N_6378);
and U8305 (N_8305,N_6847,N_7377);
nand U8306 (N_8306,N_7022,N_6469);
and U8307 (N_8307,N_7303,N_7064);
or U8308 (N_8308,N_6272,N_7642);
nand U8309 (N_8309,N_7764,N_6213);
and U8310 (N_8310,N_7976,N_6800);
nor U8311 (N_8311,N_6625,N_7674);
nand U8312 (N_8312,N_6833,N_7959);
or U8313 (N_8313,N_7097,N_6748);
nand U8314 (N_8314,N_7650,N_6641);
nor U8315 (N_8315,N_7280,N_7537);
nor U8316 (N_8316,N_7947,N_6719);
nor U8317 (N_8317,N_7593,N_7552);
xor U8318 (N_8318,N_6029,N_6594);
or U8319 (N_8319,N_7907,N_7370);
nand U8320 (N_8320,N_6428,N_7331);
nand U8321 (N_8321,N_6392,N_7982);
or U8322 (N_8322,N_7137,N_6341);
nand U8323 (N_8323,N_6986,N_6745);
or U8324 (N_8324,N_7861,N_7937);
or U8325 (N_8325,N_6416,N_6193);
and U8326 (N_8326,N_7336,N_7468);
nor U8327 (N_8327,N_6123,N_7078);
and U8328 (N_8328,N_6683,N_7668);
or U8329 (N_8329,N_7717,N_6535);
and U8330 (N_8330,N_6558,N_6880);
nor U8331 (N_8331,N_7429,N_6092);
or U8332 (N_8332,N_7045,N_6970);
and U8333 (N_8333,N_7320,N_6972);
nor U8334 (N_8334,N_7284,N_6046);
or U8335 (N_8335,N_7458,N_7778);
and U8336 (N_8336,N_7672,N_7164);
or U8337 (N_8337,N_7339,N_7646);
nand U8338 (N_8338,N_7418,N_6326);
and U8339 (N_8339,N_6187,N_6536);
nand U8340 (N_8340,N_6774,N_6360);
and U8341 (N_8341,N_7939,N_6838);
nor U8342 (N_8342,N_7821,N_6896);
nor U8343 (N_8343,N_6949,N_6654);
nand U8344 (N_8344,N_6706,N_6509);
or U8345 (N_8345,N_7459,N_7933);
or U8346 (N_8346,N_7752,N_7110);
or U8347 (N_8347,N_7076,N_6579);
and U8348 (N_8348,N_7894,N_6430);
nand U8349 (N_8349,N_6829,N_6612);
or U8350 (N_8350,N_6931,N_7994);
or U8351 (N_8351,N_7322,N_6194);
and U8352 (N_8352,N_6842,N_6600);
or U8353 (N_8353,N_7008,N_7016);
nand U8354 (N_8354,N_6695,N_7815);
or U8355 (N_8355,N_7344,N_7475);
nand U8356 (N_8356,N_7746,N_7188);
or U8357 (N_8357,N_7724,N_6060);
nand U8358 (N_8358,N_7456,N_7989);
nor U8359 (N_8359,N_6134,N_6018);
or U8360 (N_8360,N_7906,N_6007);
nor U8361 (N_8361,N_6574,N_6668);
nor U8362 (N_8362,N_7613,N_6334);
nor U8363 (N_8363,N_6653,N_7685);
xor U8364 (N_8364,N_6534,N_6488);
nor U8365 (N_8365,N_7924,N_7046);
and U8366 (N_8366,N_6278,N_7927);
xnor U8367 (N_8367,N_6503,N_7543);
nand U8368 (N_8368,N_7026,N_6215);
xnor U8369 (N_8369,N_7970,N_6973);
nand U8370 (N_8370,N_7119,N_7675);
nor U8371 (N_8371,N_6915,N_7680);
and U8372 (N_8372,N_7601,N_6597);
or U8373 (N_8373,N_7503,N_7974);
nor U8374 (N_8374,N_7958,N_6399);
nand U8375 (N_8375,N_7071,N_7736);
or U8376 (N_8376,N_7971,N_6627);
or U8377 (N_8377,N_6177,N_7829);
nand U8378 (N_8378,N_7080,N_6642);
nand U8379 (N_8379,N_7651,N_6439);
or U8380 (N_8380,N_6598,N_7997);
nor U8381 (N_8381,N_6836,N_6831);
and U8382 (N_8382,N_6377,N_6934);
or U8383 (N_8383,N_7791,N_7547);
and U8384 (N_8384,N_7883,N_7460);
nand U8385 (N_8385,N_6333,N_6170);
nor U8386 (N_8386,N_7349,N_7086);
or U8387 (N_8387,N_7232,N_7911);
or U8388 (N_8388,N_7480,N_7501);
nand U8389 (N_8389,N_7731,N_7641);
or U8390 (N_8390,N_6383,N_7443);
or U8391 (N_8391,N_6989,N_6442);
or U8392 (N_8392,N_6089,N_6126);
nand U8393 (N_8393,N_7877,N_6940);
or U8394 (N_8394,N_6878,N_7903);
xor U8395 (N_8395,N_7839,N_7068);
nor U8396 (N_8396,N_6898,N_7003);
nor U8397 (N_8397,N_6456,N_6454);
nand U8398 (N_8398,N_7857,N_6262);
or U8399 (N_8399,N_6470,N_6306);
nor U8400 (N_8400,N_6784,N_7645);
nand U8401 (N_8401,N_7270,N_7759);
and U8402 (N_8402,N_6403,N_7301);
or U8403 (N_8403,N_6008,N_7814);
and U8404 (N_8404,N_7089,N_6125);
nand U8405 (N_8405,N_6752,N_6429);
nand U8406 (N_8406,N_6261,N_6724);
and U8407 (N_8407,N_7114,N_6930);
nor U8408 (N_8408,N_6434,N_7028);
nand U8409 (N_8409,N_7831,N_6807);
nand U8410 (N_8410,N_7353,N_6138);
or U8411 (N_8411,N_6063,N_6853);
or U8412 (N_8412,N_7719,N_7216);
nand U8413 (N_8413,N_7105,N_6691);
or U8414 (N_8414,N_6303,N_6347);
and U8415 (N_8415,N_6395,N_6529);
nand U8416 (N_8416,N_7985,N_7094);
nor U8417 (N_8417,N_6349,N_7152);
or U8418 (N_8418,N_7364,N_7900);
nand U8419 (N_8419,N_6153,N_6049);
nand U8420 (N_8420,N_6891,N_7908);
xnor U8421 (N_8421,N_6298,N_6149);
nand U8422 (N_8422,N_6267,N_6811);
and U8423 (N_8423,N_6121,N_6791);
nor U8424 (N_8424,N_6924,N_7250);
and U8425 (N_8425,N_6947,N_6452);
xor U8426 (N_8426,N_6167,N_6795);
and U8427 (N_8427,N_7820,N_6458);
or U8428 (N_8428,N_6938,N_7557);
or U8429 (N_8429,N_6148,N_7238);
nor U8430 (N_8430,N_7230,N_6796);
nand U8431 (N_8431,N_7892,N_6276);
and U8432 (N_8432,N_6315,N_6459);
or U8433 (N_8433,N_6202,N_7912);
or U8434 (N_8434,N_7487,N_6868);
nand U8435 (N_8435,N_6804,N_7750);
and U8436 (N_8436,N_7534,N_7654);
or U8437 (N_8437,N_7995,N_7587);
nor U8438 (N_8438,N_6385,N_7561);
or U8439 (N_8439,N_6307,N_6590);
nand U8440 (N_8440,N_6335,N_7031);
or U8441 (N_8441,N_7710,N_7371);
or U8442 (N_8442,N_7784,N_6238);
nor U8443 (N_8443,N_6546,N_6027);
or U8444 (N_8444,N_6605,N_6508);
and U8445 (N_8445,N_7253,N_7758);
nand U8446 (N_8446,N_7037,N_6589);
nand U8447 (N_8447,N_6806,N_6001);
nand U8448 (N_8448,N_7010,N_6220);
and U8449 (N_8449,N_7148,N_7474);
and U8450 (N_8450,N_7954,N_6480);
nor U8451 (N_8451,N_6065,N_6874);
nor U8452 (N_8452,N_7112,N_6423);
and U8453 (N_8453,N_6608,N_7657);
and U8454 (N_8454,N_7676,N_6157);
nor U8455 (N_8455,N_6179,N_6419);
or U8456 (N_8456,N_7611,N_7478);
and U8457 (N_8457,N_7918,N_7990);
and U8458 (N_8458,N_6173,N_6502);
nor U8459 (N_8459,N_7048,N_6969);
or U8460 (N_8460,N_7033,N_6435);
or U8461 (N_8461,N_6086,N_6993);
or U8462 (N_8462,N_7692,N_6024);
and U8463 (N_8463,N_7960,N_7828);
nor U8464 (N_8464,N_6369,N_7441);
or U8465 (N_8465,N_7237,N_6664);
and U8466 (N_8466,N_6394,N_6697);
xor U8467 (N_8467,N_7819,N_6643);
nor U8468 (N_8468,N_7140,N_7966);
or U8469 (N_8469,N_7880,N_7036);
nor U8470 (N_8470,N_7969,N_6393);
and U8471 (N_8471,N_7520,N_7011);
nor U8472 (N_8472,N_6257,N_6210);
or U8473 (N_8473,N_6900,N_6067);
or U8474 (N_8474,N_6779,N_7864);
and U8475 (N_8475,N_6866,N_7233);
nand U8476 (N_8476,N_6019,N_7121);
nand U8477 (N_8477,N_7763,N_6974);
nand U8478 (N_8478,N_7283,N_6929);
and U8479 (N_8479,N_7524,N_7790);
nand U8480 (N_8480,N_6048,N_6274);
or U8481 (N_8481,N_7494,N_6966);
nor U8482 (N_8482,N_7049,N_6620);
nand U8483 (N_8483,N_6857,N_6551);
and U8484 (N_8484,N_6614,N_6727);
and U8485 (N_8485,N_7863,N_6760);
nor U8486 (N_8486,N_7373,N_7816);
or U8487 (N_8487,N_7629,N_6322);
or U8488 (N_8488,N_6421,N_6015);
nor U8489 (N_8489,N_6562,N_7573);
and U8490 (N_8490,N_7538,N_7512);
nand U8491 (N_8491,N_6935,N_6523);
nand U8492 (N_8492,N_7107,N_6164);
nor U8493 (N_8493,N_6759,N_6939);
nand U8494 (N_8494,N_6075,N_6638);
and U8495 (N_8495,N_7507,N_7703);
nand U8496 (N_8496,N_6856,N_7142);
or U8497 (N_8497,N_7394,N_7930);
and U8498 (N_8498,N_6226,N_6628);
and U8499 (N_8499,N_7635,N_6030);
or U8500 (N_8500,N_7332,N_7334);
and U8501 (N_8501,N_6242,N_6616);
or U8502 (N_8502,N_7262,N_7526);
nand U8503 (N_8503,N_6773,N_6346);
and U8504 (N_8504,N_7973,N_6370);
nand U8505 (N_8505,N_6879,N_7715);
nand U8506 (N_8506,N_7868,N_6527);
nor U8507 (N_8507,N_7678,N_6834);
nand U8508 (N_8508,N_7206,N_6932);
or U8509 (N_8509,N_6521,N_7885);
or U8510 (N_8510,N_6318,N_7926);
nand U8511 (N_8511,N_6553,N_6185);
xor U8512 (N_8512,N_7014,N_7913);
nor U8513 (N_8513,N_6769,N_7333);
nor U8514 (N_8514,N_7157,N_6356);
nand U8515 (N_8515,N_7275,N_7730);
nor U8516 (N_8516,N_7035,N_7584);
nor U8517 (N_8517,N_6755,N_6288);
or U8518 (N_8518,N_7476,N_7961);
nand U8519 (N_8519,N_7102,N_7165);
nand U8520 (N_8520,N_7874,N_6189);
and U8521 (N_8521,N_6544,N_7767);
and U8522 (N_8522,N_6447,N_7628);
or U8523 (N_8523,N_7935,N_6031);
or U8524 (N_8524,N_6507,N_7789);
and U8525 (N_8525,N_6782,N_7127);
nand U8526 (N_8526,N_7700,N_7298);
nor U8527 (N_8527,N_6373,N_7286);
nor U8528 (N_8528,N_7527,N_7777);
nor U8529 (N_8529,N_7560,N_7670);
nor U8530 (N_8530,N_7663,N_7756);
and U8531 (N_8531,N_6964,N_7485);
and U8532 (N_8532,N_6374,N_7454);
or U8533 (N_8533,N_7643,N_6402);
nor U8534 (N_8534,N_7160,N_7708);
and U8535 (N_8535,N_6548,N_7354);
and U8536 (N_8536,N_7504,N_7404);
or U8537 (N_8537,N_7438,N_6978);
nand U8538 (N_8538,N_6984,N_6387);
or U8539 (N_8539,N_6692,N_6225);
nor U8540 (N_8540,N_6640,N_6586);
and U8541 (N_8541,N_6305,N_6751);
or U8542 (N_8542,N_7579,N_7944);
or U8543 (N_8543,N_6992,N_6112);
nor U8544 (N_8544,N_6368,N_7050);
nor U8545 (N_8545,N_7088,N_6854);
or U8546 (N_8546,N_7482,N_7264);
and U8547 (N_8547,N_7405,N_6746);
nand U8548 (N_8548,N_7662,N_7359);
or U8549 (N_8549,N_7998,N_7340);
nor U8550 (N_8550,N_6976,N_6504);
and U8551 (N_8551,N_6103,N_6858);
and U8552 (N_8552,N_6003,N_6105);
nand U8553 (N_8553,N_6730,N_6710);
nand U8554 (N_8554,N_7797,N_6825);
nor U8555 (N_8555,N_7925,N_7013);
nor U8556 (N_8556,N_7401,N_6212);
and U8557 (N_8557,N_7223,N_6296);
nor U8558 (N_8558,N_7801,N_6181);
and U8559 (N_8559,N_6665,N_7147);
or U8560 (N_8560,N_7436,N_6792);
and U8561 (N_8561,N_7346,N_6634);
nor U8562 (N_8562,N_7198,N_6118);
nor U8563 (N_8563,N_6091,N_7988);
nand U8564 (N_8564,N_7041,N_6635);
nor U8565 (N_8565,N_6717,N_6151);
or U8566 (N_8566,N_6082,N_6160);
and U8567 (N_8567,N_7384,N_7936);
nor U8568 (N_8568,N_7633,N_6699);
nor U8569 (N_8569,N_7721,N_6516);
and U8570 (N_8570,N_7606,N_6244);
and U8571 (N_8571,N_7430,N_7285);
nand U8572 (N_8572,N_6639,N_6106);
nor U8573 (N_8573,N_6043,N_6270);
and U8574 (N_8574,N_6400,N_7655);
or U8575 (N_8575,N_6453,N_7956);
and U8576 (N_8576,N_7098,N_6191);
nand U8577 (N_8577,N_7575,N_7742);
nor U8578 (N_8578,N_6491,N_7051);
nor U8579 (N_8579,N_6293,N_6712);
and U8580 (N_8580,N_6292,N_7932);
nand U8581 (N_8581,N_6505,N_6077);
nor U8582 (N_8582,N_6816,N_7996);
and U8583 (N_8583,N_6351,N_6520);
and U8584 (N_8584,N_7363,N_6788);
and U8585 (N_8585,N_6636,N_6556);
nand U8586 (N_8586,N_7766,N_6809);
nor U8587 (N_8587,N_6519,N_6433);
and U8588 (N_8588,N_6006,N_6413);
nor U8589 (N_8589,N_7185,N_6154);
and U8590 (N_8590,N_6268,N_7862);
nor U8591 (N_8591,N_6472,N_7701);
or U8592 (N_8592,N_6083,N_7084);
or U8593 (N_8593,N_6645,N_7315);
and U8594 (N_8594,N_7599,N_7077);
nand U8595 (N_8595,N_7929,N_6563);
nand U8596 (N_8596,N_6777,N_7983);
nand U8597 (N_8597,N_7856,N_6273);
or U8598 (N_8598,N_7902,N_6038);
nor U8599 (N_8599,N_7822,N_7548);
or U8600 (N_8600,N_6530,N_7882);
and U8601 (N_8601,N_6451,N_7397);
nor U8602 (N_8602,N_6647,N_6814);
nor U8603 (N_8603,N_7588,N_7390);
or U8604 (N_8604,N_6216,N_6045);
and U8605 (N_8605,N_7639,N_6420);
or U8606 (N_8606,N_7473,N_7461);
nand U8607 (N_8607,N_6725,N_6485);
xor U8608 (N_8608,N_7891,N_7723);
nor U8609 (N_8609,N_6818,N_7433);
nor U8610 (N_8610,N_7805,N_6705);
and U8611 (N_8611,N_6672,N_7132);
and U8612 (N_8612,N_6740,N_7602);
or U8613 (N_8613,N_7844,N_7375);
or U8614 (N_8614,N_7212,N_7024);
or U8615 (N_8615,N_7949,N_6821);
nand U8616 (N_8616,N_7551,N_6790);
and U8617 (N_8617,N_7341,N_7109);
nor U8618 (N_8618,N_6894,N_7416);
nor U8619 (N_8619,N_7852,N_7310);
and U8620 (N_8620,N_6890,N_6384);
nor U8621 (N_8621,N_6876,N_6610);
and U8622 (N_8622,N_7699,N_6097);
nor U8623 (N_8623,N_6707,N_6566);
nand U8624 (N_8624,N_6100,N_6926);
nor U8625 (N_8625,N_7385,N_6243);
nand U8626 (N_8626,N_6136,N_6670);
nor U8627 (N_8627,N_7690,N_7753);
nor U8628 (N_8628,N_6036,N_6482);
and U8629 (N_8629,N_7802,N_7774);
or U8630 (N_8630,N_6289,N_7168);
or U8631 (N_8631,N_7841,N_7975);
nand U8632 (N_8632,N_6371,N_7369);
nand U8633 (N_8633,N_6765,N_6000);
or U8634 (N_8634,N_6117,N_6997);
nand U8635 (N_8635,N_6113,N_7840);
or U8636 (N_8636,N_7235,N_7833);
nor U8637 (N_8637,N_7773,N_6316);
nand U8638 (N_8638,N_7824,N_7192);
or U8639 (N_8639,N_7876,N_6165);
nor U8640 (N_8640,N_7873,N_7305);
and U8641 (N_8641,N_6253,N_7667);
or U8642 (N_8642,N_7953,N_7169);
nor U8643 (N_8643,N_6230,N_6671);
or U8644 (N_8644,N_6352,N_7291);
or U8645 (N_8645,N_7860,N_6069);
xor U8646 (N_8646,N_7531,N_7019);
and U8647 (N_8647,N_7795,N_7296);
xor U8648 (N_8648,N_7739,N_6679);
nor U8649 (N_8649,N_6688,N_6802);
nand U8650 (N_8650,N_6308,N_7408);
nand U8651 (N_8651,N_6304,N_7222);
and U8652 (N_8652,N_7155,N_6889);
nor U8653 (N_8653,N_6146,N_7673);
or U8654 (N_8654,N_6460,N_7916);
nand U8655 (N_8655,N_6178,N_6287);
and U8656 (N_8656,N_6312,N_6764);
nor U8657 (N_8657,N_6626,N_6388);
nand U8658 (N_8658,N_7295,N_7922);
or U8659 (N_8659,N_6427,N_7665);
or U8660 (N_8660,N_6020,N_7190);
nor U8661 (N_8661,N_6059,N_7017);
and U8662 (N_8662,N_6005,N_6206);
nor U8663 (N_8663,N_6090,N_7964);
or U8664 (N_8664,N_7254,N_6265);
nor U8665 (N_8665,N_6156,N_7709);
nor U8666 (N_8666,N_7811,N_6014);
and U8667 (N_8667,N_6793,N_7770);
or U8668 (N_8668,N_7267,N_7869);
or U8669 (N_8669,N_6204,N_6203);
or U8670 (N_8670,N_7615,N_6471);
nor U8671 (N_8671,N_6526,N_6088);
and U8672 (N_8672,N_6431,N_6076);
nor U8673 (N_8673,N_7063,N_6127);
nor U8674 (N_8674,N_7452,N_7749);
and U8675 (N_8675,N_6074,N_6613);
and U8676 (N_8676,N_6397,N_7732);
or U8677 (N_8677,N_6284,N_6621);
or U8678 (N_8678,N_7917,N_7259);
or U8679 (N_8679,N_6228,N_7358);
nor U8680 (N_8680,N_7410,N_7890);
and U8681 (N_8681,N_7817,N_6552);
or U8682 (N_8682,N_7870,N_6942);
nand U8683 (N_8683,N_7090,N_7488);
nor U8684 (N_8684,N_7608,N_7942);
or U8685 (N_8685,N_6467,N_7943);
nor U8686 (N_8686,N_7075,N_7263);
nand U8687 (N_8687,N_6741,N_7012);
nor U8688 (N_8688,N_6489,N_6595);
nand U8689 (N_8689,N_6686,N_7714);
or U8690 (N_8690,N_7835,N_7304);
and U8691 (N_8691,N_7484,N_7388);
nand U8692 (N_8692,N_6532,N_6694);
or U8693 (N_8693,N_6855,N_6240);
nand U8694 (N_8694,N_6064,N_6649);
nor U8695 (N_8695,N_7001,N_7272);
and U8696 (N_8696,N_6099,N_7243);
or U8697 (N_8697,N_6537,N_6236);
nor U8698 (N_8698,N_6959,N_7415);
nand U8699 (N_8699,N_6742,N_6184);
xor U8700 (N_8700,N_7556,N_6839);
or U8701 (N_8701,N_6144,N_7276);
nor U8702 (N_8702,N_6629,N_7294);
nand U8703 (N_8703,N_7855,N_7728);
nor U8704 (N_8704,N_7920,N_6463);
nor U8705 (N_8705,N_6175,N_6150);
and U8706 (N_8706,N_7553,N_6728);
nand U8707 (N_8707,N_7957,N_6299);
and U8708 (N_8708,N_6279,N_7386);
nand U8709 (N_8709,N_6946,N_7647);
or U8710 (N_8710,N_6155,N_7025);
or U8711 (N_8711,N_6619,N_7725);
nor U8712 (N_8712,N_7631,N_7895);
nand U8713 (N_8713,N_6669,N_6300);
and U8714 (N_8714,N_6685,N_7269);
or U8715 (N_8715,N_6901,N_6426);
nor U8716 (N_8716,N_7159,N_6034);
nand U8717 (N_8717,N_6678,N_7380);
or U8718 (N_8718,N_7299,N_7603);
nand U8719 (N_8719,N_6133,N_7338);
and U8720 (N_8720,N_6518,N_6500);
and U8721 (N_8721,N_7151,N_6286);
nor U8722 (N_8722,N_6910,N_6660);
nor U8723 (N_8723,N_7187,N_6313);
nand U8724 (N_8724,N_7843,N_7252);
nand U8725 (N_8725,N_6124,N_7854);
or U8726 (N_8726,N_6142,N_6365);
and U8727 (N_8727,N_7361,N_6698);
or U8728 (N_8728,N_7522,N_6736);
nand U8729 (N_8729,N_6441,N_6473);
nand U8730 (N_8730,N_7529,N_6152);
or U8731 (N_8731,N_7712,N_6171);
or U8732 (N_8732,N_7977,N_6690);
nor U8733 (N_8733,N_7355,N_7923);
and U8734 (N_8734,N_6953,N_7218);
nand U8735 (N_8735,N_6140,N_7006);
or U8736 (N_8736,N_7260,N_7279);
nand U8737 (N_8737,N_7986,N_7043);
xor U8738 (N_8738,N_6958,N_6432);
xor U8739 (N_8739,N_7649,N_6514);
nor U8740 (N_8740,N_7465,N_7741);
nor U8741 (N_8741,N_6066,N_7948);
or U8742 (N_8742,N_6565,N_7173);
nand U8743 (N_8743,N_7576,N_7330);
nand U8744 (N_8744,N_7391,N_7652);
and U8745 (N_8745,N_6477,N_6320);
or U8746 (N_8746,N_6919,N_7609);
or U8747 (N_8747,N_6734,N_7605);
nand U8748 (N_8748,N_7744,N_7889);
nor U8749 (N_8749,N_6511,N_6864);
nand U8750 (N_8750,N_7660,N_7463);
nor U8751 (N_8751,N_7992,N_7827);
nand U8752 (N_8752,N_7788,N_6042);
and U8753 (N_8753,N_6302,N_6568);
or U8754 (N_8754,N_7886,N_6207);
or U8755 (N_8755,N_6372,N_6120);
or U8756 (N_8756,N_7372,N_7776);
or U8757 (N_8757,N_6781,N_7622);
nor U8758 (N_8758,N_6650,N_7671);
and U8759 (N_8759,N_6581,N_6623);
nor U8760 (N_8760,N_7106,N_7568);
nand U8761 (N_8761,N_6166,N_6711);
or U8762 (N_8762,N_6961,N_6886);
and U8763 (N_8763,N_7577,N_6844);
nor U8764 (N_8764,N_7425,N_7030);
or U8765 (N_8765,N_6954,N_7794);
nor U8766 (N_8766,N_7199,N_6658);
or U8767 (N_8767,N_6499,N_6539);
and U8768 (N_8768,N_6227,N_6337);
or U8769 (N_8769,N_7204,N_6797);
and U8770 (N_8770,N_7525,N_6823);
and U8771 (N_8771,N_6450,N_6248);
or U8772 (N_8772,N_7931,N_7447);
and U8773 (N_8773,N_6944,N_7901);
or U8774 (N_8774,N_7682,N_7470);
nor U8775 (N_8775,N_6776,N_6081);
or U8776 (N_8776,N_6161,N_7838);
and U8777 (N_8777,N_7172,N_6550);
nor U8778 (N_8778,N_7120,N_7442);
nand U8779 (N_8779,N_6028,N_7693);
and U8780 (N_8780,N_6681,N_7357);
nor U8781 (N_8781,N_7392,N_7792);
or U8782 (N_8782,N_6411,N_7034);
nor U8783 (N_8783,N_6657,N_6229);
nand U8784 (N_8784,N_7189,N_7145);
and U8785 (N_8785,N_6314,N_7716);
nand U8786 (N_8786,N_6988,N_6412);
and U8787 (N_8787,N_6245,N_6701);
nand U8788 (N_8788,N_7872,N_7226);
or U8789 (N_8789,N_6861,N_6406);
or U8790 (N_8790,N_7052,N_6094);
or U8791 (N_8791,N_7596,N_7938);
nor U8792 (N_8792,N_6775,N_7834);
and U8793 (N_8793,N_7705,N_6122);
and U8794 (N_8794,N_6407,N_7704);
nor U8795 (N_8795,N_6888,N_6754);
nand U8796 (N_8796,N_7445,N_7362);
nand U8797 (N_8797,N_7249,N_7455);
or U8798 (N_8798,N_6655,N_7733);
or U8799 (N_8799,N_7486,N_7302);
nand U8800 (N_8800,N_7083,N_6218);
or U8801 (N_8801,N_7124,N_6061);
nor U8802 (N_8802,N_6914,N_7312);
and U8803 (N_8803,N_7131,N_7826);
and U8804 (N_8804,N_7471,N_7919);
nand U8805 (N_8805,N_6241,N_6484);
nor U8806 (N_8806,N_7489,N_6824);
and U8807 (N_8807,N_7419,N_7499);
nor U8808 (N_8808,N_6055,N_6963);
nand U8809 (N_8809,N_7590,N_6231);
xor U8810 (N_8810,N_6444,N_7518);
nand U8811 (N_8811,N_7754,N_7427);
and U8812 (N_8812,N_7626,N_7205);
nand U8813 (N_8813,N_6785,N_7178);
nand U8814 (N_8814,N_7968,N_7808);
nor U8815 (N_8815,N_6709,N_7439);
and U8816 (N_8816,N_7683,N_7694);
nand U8817 (N_8817,N_6379,N_6522);
xor U8818 (N_8818,N_6443,N_7627);
or U8819 (N_8819,N_7787,N_6666);
or U8820 (N_8820,N_6994,N_7888);
nor U8821 (N_8821,N_6813,N_6999);
and U8822 (N_8822,N_7002,N_7400);
or U8823 (N_8823,N_7343,N_7366);
nor U8824 (N_8824,N_6543,N_6819);
nand U8825 (N_8825,N_7406,N_7846);
nand U8826 (N_8826,N_7563,N_6084);
nand U8827 (N_8827,N_7644,N_6541);
nor U8828 (N_8828,N_6474,N_6182);
nor U8829 (N_8829,N_6859,N_6032);
and U8830 (N_8830,N_6515,N_6980);
or U8831 (N_8831,N_6129,N_7963);
nor U8832 (N_8832,N_6147,N_7921);
and U8833 (N_8833,N_6235,N_6652);
nand U8834 (N_8834,N_7345,N_6936);
nor U8835 (N_8835,N_7783,N_7479);
nand U8836 (N_8836,N_6332,N_7450);
nor U8837 (N_8837,N_7659,N_6656);
nor U8838 (N_8838,N_7074,N_7481);
nand U8839 (N_8839,N_7617,N_7417);
nor U8840 (N_8840,N_6850,N_6892);
nor U8841 (N_8841,N_6023,N_6884);
and U8842 (N_8842,N_6396,N_7813);
and U8843 (N_8843,N_6145,N_6436);
and U8844 (N_8844,N_6040,N_6448);
and U8845 (N_8845,N_7851,N_7904);
xnor U8846 (N_8846,N_6985,N_6358);
xnor U8847 (N_8847,N_6095,N_7592);
nor U8848 (N_8848,N_6367,N_6275);
nor U8849 (N_8849,N_6525,N_7307);
and U8850 (N_8850,N_7881,N_6667);
or U8851 (N_8851,N_7656,N_7200);
nor U8852 (N_8852,N_6902,N_6714);
or U8853 (N_8853,N_6478,N_7318);
and U8854 (N_8854,N_7572,N_6440);
nor U8855 (N_8855,N_6979,N_7065);
nor U8856 (N_8856,N_6249,N_7081);
nand U8857 (N_8857,N_7987,N_7493);
xnor U8858 (N_8858,N_6723,N_7681);
nand U8859 (N_8859,N_6176,N_6863);
and U8860 (N_8860,N_6540,N_7111);
nor U8861 (N_8861,N_7896,N_7422);
nor U8862 (N_8862,N_7502,N_7347);
nor U8863 (N_8863,N_6584,N_7096);
and U8864 (N_8864,N_7695,N_7161);
or U8865 (N_8865,N_6186,N_6912);
nor U8866 (N_8866,N_7595,N_7760);
or U8867 (N_8867,N_7115,N_6425);
nor U8868 (N_8868,N_6917,N_6569);
nand U8869 (N_8869,N_6983,N_7444);
xnor U8870 (N_8870,N_6054,N_6646);
or U8871 (N_8871,N_6545,N_6222);
nand U8872 (N_8872,N_7196,N_6116);
nor U8873 (N_8873,N_7453,N_6533);
xnor U8874 (N_8874,N_7411,N_7981);
or U8875 (N_8875,N_6677,N_7965);
nor U8876 (N_8876,N_6713,N_7085);
nor U8877 (N_8877,N_6266,N_7521);
or U8878 (N_8878,N_7549,N_7591);
nand U8879 (N_8879,N_7500,N_6922);
nor U8880 (N_8880,N_6033,N_6496);
and U8881 (N_8881,N_7382,N_7490);
nand U8882 (N_8882,N_6375,N_6869);
or U8883 (N_8883,N_6923,N_7618);
or U8884 (N_8884,N_7757,N_7570);
and U8885 (N_8885,N_7689,N_6438);
or U8886 (N_8886,N_7070,N_6381);
nand U8887 (N_8887,N_7544,N_6871);
nand U8888 (N_8888,N_7597,N_7910);
and U8889 (N_8889,N_6722,N_7653);
and U8890 (N_8890,N_7803,N_6217);
or U8891 (N_8891,N_6920,N_6348);
and U8892 (N_8892,N_7040,N_7337);
or U8893 (N_8893,N_6757,N_7323);
or U8894 (N_8894,N_6845,N_6115);
nor U8895 (N_8895,N_6011,N_7066);
or U8896 (N_8896,N_6786,N_6234);
or U8897 (N_8897,N_6624,N_7091);
and U8898 (N_8898,N_7457,N_7586);
and U8899 (N_8899,N_7300,N_6962);
nor U8900 (N_8900,N_7449,N_6418);
nand U8901 (N_8901,N_6409,N_7073);
nand U8902 (N_8902,N_7117,N_7899);
and U8903 (N_8903,N_6324,N_7256);
nand U8904 (N_8904,N_7044,N_6209);
nor U8905 (N_8905,N_7177,N_6585);
or U8906 (N_8906,N_6197,N_6607);
or U8907 (N_8907,N_6753,N_7316);
nand U8908 (N_8908,N_7059,N_6353);
nor U8909 (N_8909,N_6633,N_6883);
nor U8910 (N_8910,N_6571,N_7967);
nand U8911 (N_8911,N_6987,N_6843);
xor U8912 (N_8912,N_6271,N_7057);
nand U8913 (N_8913,N_7887,N_7823);
nor U8914 (N_8914,N_6363,N_7623);
nand U8915 (N_8915,N_7412,N_7574);
nor U8916 (N_8916,N_6131,N_7495);
or U8917 (N_8917,N_7154,N_6977);
and U8918 (N_8918,N_6336,N_6259);
nand U8919 (N_8919,N_7523,N_6950);
nand U8920 (N_8920,N_7180,N_7979);
and U8921 (N_8921,N_7619,N_6632);
or U8922 (N_8922,N_6141,N_6386);
and U8923 (N_8923,N_7589,N_7497);
and U8924 (N_8924,N_6783,N_6990);
nor U8925 (N_8925,N_7706,N_6846);
nor U8926 (N_8926,N_6680,N_7467);
nor U8927 (N_8927,N_6794,N_7224);
nand U8928 (N_8928,N_7513,N_7755);
nand U8929 (N_8929,N_7535,N_6547);
or U8930 (N_8930,N_6466,N_7242);
nor U8931 (N_8931,N_7782,N_6602);
nor U8932 (N_8932,N_7208,N_6468);
or U8933 (N_8933,N_7225,N_6401);
and U8934 (N_8934,N_6104,N_7536);
nand U8935 (N_8935,N_7234,N_7564);
and U8936 (N_8936,N_7374,N_6849);
and U8937 (N_8937,N_6269,N_7055);
or U8938 (N_8938,N_7737,N_6815);
nand U8939 (N_8939,N_7847,N_6583);
or U8940 (N_8940,N_6497,N_7483);
or U8941 (N_8941,N_6555,N_7898);
nor U8942 (N_8942,N_7440,N_6280);
and U8943 (N_8943,N_6481,N_6867);
nor U8944 (N_8944,N_7620,N_7058);
or U8945 (N_8945,N_7221,N_7039);
nand U8946 (N_8946,N_6080,N_7143);
and U8947 (N_8947,N_7432,N_7054);
nor U8948 (N_8948,N_7268,N_6035);
nand U8949 (N_8949,N_7122,N_6513);
nand U8950 (N_8950,N_7248,N_6592);
or U8951 (N_8951,N_6422,N_6911);
nor U8952 (N_8952,N_6948,N_7352);
or U8953 (N_8953,N_6196,N_7219);
and U8954 (N_8954,N_6872,N_6037);
nand U8955 (N_8955,N_7517,N_7600);
or U8956 (N_8956,N_6380,N_6906);
nand U8957 (N_8957,N_6703,N_6281);
nand U8958 (N_8958,N_6732,N_6617);
nand U8959 (N_8959,N_6039,N_7069);
nor U8960 (N_8960,N_6739,N_7207);
nand U8961 (N_8961,N_7780,N_7849);
nor U8962 (N_8962,N_7414,N_6010);
nand U8963 (N_8963,N_6778,N_7087);
and U8964 (N_8964,N_7571,N_6247);
nand U8965 (N_8965,N_7677,N_7203);
or U8966 (N_8966,N_6907,N_6801);
and U8967 (N_8967,N_7376,N_7239);
nor U8968 (N_8968,N_6310,N_7348);
nand U8969 (N_8969,N_6618,N_6087);
and U8970 (N_8970,N_7228,N_6512);
nand U8971 (N_8971,N_6524,N_7134);
nor U8972 (N_8972,N_7321,N_7684);
and U8973 (N_8973,N_7182,N_7103);
and U8974 (N_8974,N_7625,N_7768);
and U8975 (N_8975,N_7351,N_7211);
or U8976 (N_8976,N_7546,N_6264);
or U8977 (N_8977,N_7984,N_6344);
nand U8978 (N_8978,N_7761,N_6747);
nor U8979 (N_8979,N_6250,N_7247);
nand U8980 (N_8980,N_6359,N_7265);
and U8981 (N_8981,N_7420,N_7491);
nor U8982 (N_8982,N_7634,N_6704);
or U8983 (N_8983,N_7395,N_7785);
and U8984 (N_8984,N_6277,N_6559);
nand U8985 (N_8985,N_6198,N_7100);
nor U8986 (N_8986,N_6870,N_7865);
nand U8987 (N_8987,N_6549,N_6941);
nand U8988 (N_8988,N_7274,N_6971);
and U8989 (N_8989,N_7978,N_7648);
and U8990 (N_8990,N_7993,N_7687);
and U8991 (N_8991,N_6168,N_6343);
or U8992 (N_8992,N_6968,N_6881);
and U8993 (N_8993,N_7032,N_7515);
nor U8994 (N_8994,N_7509,N_6345);
nand U8995 (N_8995,N_6071,N_6573);
nor U8996 (N_8996,N_7389,N_7125);
and U8997 (N_8997,N_7848,N_7738);
and U8998 (N_8998,N_6016,N_6810);
nand U8999 (N_8999,N_7765,N_7751);
and U9000 (N_9000,N_6476,N_6676);
nor U9001 (N_9001,N_7189,N_6946);
nand U9002 (N_9002,N_6011,N_7087);
or U9003 (N_9003,N_7840,N_6194);
nand U9004 (N_9004,N_6315,N_7207);
or U9005 (N_9005,N_7941,N_6541);
and U9006 (N_9006,N_6693,N_6731);
or U9007 (N_9007,N_6573,N_6633);
or U9008 (N_9008,N_7759,N_7903);
nand U9009 (N_9009,N_7297,N_7468);
nor U9010 (N_9010,N_7824,N_7419);
and U9011 (N_9011,N_7252,N_7749);
nor U9012 (N_9012,N_7375,N_6080);
nand U9013 (N_9013,N_6387,N_7016);
and U9014 (N_9014,N_6795,N_7848);
nor U9015 (N_9015,N_7937,N_6287);
and U9016 (N_9016,N_6114,N_6597);
and U9017 (N_9017,N_6307,N_7637);
nand U9018 (N_9018,N_6327,N_6104);
or U9019 (N_9019,N_6852,N_6233);
and U9020 (N_9020,N_7634,N_7395);
or U9021 (N_9021,N_7143,N_6945);
and U9022 (N_9022,N_7441,N_6374);
or U9023 (N_9023,N_6297,N_6998);
or U9024 (N_9024,N_7274,N_6263);
or U9025 (N_9025,N_6819,N_6761);
or U9026 (N_9026,N_7462,N_7639);
and U9027 (N_9027,N_6138,N_7320);
and U9028 (N_9028,N_7950,N_6536);
nor U9029 (N_9029,N_7627,N_6863);
nor U9030 (N_9030,N_7839,N_7962);
nor U9031 (N_9031,N_6877,N_6766);
and U9032 (N_9032,N_7711,N_6032);
or U9033 (N_9033,N_6329,N_7693);
nand U9034 (N_9034,N_7454,N_7921);
nand U9035 (N_9035,N_7892,N_7370);
and U9036 (N_9036,N_7516,N_6694);
or U9037 (N_9037,N_6964,N_6106);
nor U9038 (N_9038,N_6856,N_7607);
xor U9039 (N_9039,N_6936,N_6439);
or U9040 (N_9040,N_7767,N_6065);
nor U9041 (N_9041,N_6139,N_7145);
or U9042 (N_9042,N_6552,N_7932);
nand U9043 (N_9043,N_6626,N_7424);
and U9044 (N_9044,N_7192,N_6482);
nand U9045 (N_9045,N_6298,N_6235);
nand U9046 (N_9046,N_7231,N_6370);
and U9047 (N_9047,N_6186,N_6852);
nor U9048 (N_9048,N_7060,N_7849);
and U9049 (N_9049,N_7921,N_6401);
or U9050 (N_9050,N_6056,N_6499);
nor U9051 (N_9051,N_6763,N_7417);
nand U9052 (N_9052,N_6337,N_7991);
nand U9053 (N_9053,N_6264,N_6103);
nand U9054 (N_9054,N_6424,N_6229);
nand U9055 (N_9055,N_7041,N_6616);
nor U9056 (N_9056,N_7371,N_6646);
nand U9057 (N_9057,N_6062,N_6400);
nand U9058 (N_9058,N_6578,N_7223);
or U9059 (N_9059,N_6309,N_6012);
nor U9060 (N_9060,N_6273,N_7226);
or U9061 (N_9061,N_7648,N_6519);
nor U9062 (N_9062,N_6892,N_6480);
or U9063 (N_9063,N_6117,N_7645);
nor U9064 (N_9064,N_7005,N_6125);
nor U9065 (N_9065,N_6848,N_6650);
and U9066 (N_9066,N_7645,N_6239);
or U9067 (N_9067,N_6075,N_6820);
nand U9068 (N_9068,N_7352,N_6158);
xor U9069 (N_9069,N_6287,N_7846);
and U9070 (N_9070,N_6283,N_6157);
nor U9071 (N_9071,N_6858,N_7309);
nand U9072 (N_9072,N_6964,N_6684);
and U9073 (N_9073,N_7876,N_6731);
nand U9074 (N_9074,N_6710,N_7433);
and U9075 (N_9075,N_6694,N_6776);
or U9076 (N_9076,N_7587,N_6380);
nor U9077 (N_9077,N_6756,N_6377);
nand U9078 (N_9078,N_6557,N_7119);
or U9079 (N_9079,N_7487,N_7912);
nor U9080 (N_9080,N_6964,N_6037);
nor U9081 (N_9081,N_7779,N_6004);
or U9082 (N_9082,N_7630,N_7644);
or U9083 (N_9083,N_7754,N_6682);
nor U9084 (N_9084,N_7664,N_6990);
nor U9085 (N_9085,N_6431,N_6340);
xor U9086 (N_9086,N_6905,N_6307);
nor U9087 (N_9087,N_7682,N_7172);
and U9088 (N_9088,N_6314,N_6586);
and U9089 (N_9089,N_6581,N_7501);
and U9090 (N_9090,N_6144,N_6734);
and U9091 (N_9091,N_6266,N_7554);
nor U9092 (N_9092,N_6245,N_6188);
or U9093 (N_9093,N_6993,N_6352);
xor U9094 (N_9094,N_7988,N_7105);
nor U9095 (N_9095,N_7701,N_6648);
nand U9096 (N_9096,N_6528,N_6682);
or U9097 (N_9097,N_6915,N_6859);
and U9098 (N_9098,N_6081,N_6950);
or U9099 (N_9099,N_6798,N_7101);
nor U9100 (N_9100,N_7939,N_6779);
and U9101 (N_9101,N_6404,N_6788);
and U9102 (N_9102,N_7952,N_6555);
nand U9103 (N_9103,N_7824,N_7316);
and U9104 (N_9104,N_6639,N_6763);
and U9105 (N_9105,N_7518,N_7514);
nand U9106 (N_9106,N_7832,N_6577);
and U9107 (N_9107,N_7929,N_7289);
and U9108 (N_9108,N_6045,N_7509);
or U9109 (N_9109,N_7250,N_6053);
or U9110 (N_9110,N_7145,N_7879);
nor U9111 (N_9111,N_6884,N_7971);
nor U9112 (N_9112,N_7126,N_7016);
nand U9113 (N_9113,N_7046,N_7705);
xor U9114 (N_9114,N_7147,N_7890);
nor U9115 (N_9115,N_6167,N_6260);
nor U9116 (N_9116,N_7928,N_6037);
or U9117 (N_9117,N_7177,N_7583);
or U9118 (N_9118,N_7154,N_6605);
and U9119 (N_9119,N_6675,N_6415);
or U9120 (N_9120,N_7557,N_6878);
and U9121 (N_9121,N_7950,N_7642);
or U9122 (N_9122,N_7313,N_7831);
and U9123 (N_9123,N_6146,N_6916);
nor U9124 (N_9124,N_7863,N_6008);
and U9125 (N_9125,N_7302,N_6536);
nand U9126 (N_9126,N_7374,N_7987);
and U9127 (N_9127,N_6894,N_7953);
or U9128 (N_9128,N_6644,N_6629);
or U9129 (N_9129,N_6471,N_6760);
nand U9130 (N_9130,N_6298,N_6116);
xor U9131 (N_9131,N_7300,N_7273);
xor U9132 (N_9132,N_7115,N_6762);
or U9133 (N_9133,N_6258,N_7264);
nand U9134 (N_9134,N_6682,N_7081);
nor U9135 (N_9135,N_7523,N_7008);
or U9136 (N_9136,N_6794,N_6137);
or U9137 (N_9137,N_7056,N_7248);
nand U9138 (N_9138,N_6174,N_7212);
or U9139 (N_9139,N_6844,N_6323);
nor U9140 (N_9140,N_6261,N_7567);
nor U9141 (N_9141,N_7954,N_7133);
and U9142 (N_9142,N_7894,N_7390);
or U9143 (N_9143,N_7695,N_7910);
nand U9144 (N_9144,N_7898,N_7390);
nand U9145 (N_9145,N_7157,N_7421);
and U9146 (N_9146,N_7148,N_7398);
nor U9147 (N_9147,N_7989,N_7106);
nor U9148 (N_9148,N_6155,N_7428);
or U9149 (N_9149,N_6567,N_6510);
nor U9150 (N_9150,N_6245,N_7167);
nand U9151 (N_9151,N_6307,N_7407);
nor U9152 (N_9152,N_7144,N_7332);
nand U9153 (N_9153,N_6095,N_7641);
nor U9154 (N_9154,N_6163,N_6729);
nor U9155 (N_9155,N_7837,N_7156);
or U9156 (N_9156,N_7882,N_6457);
nand U9157 (N_9157,N_6160,N_6361);
and U9158 (N_9158,N_6659,N_6842);
nand U9159 (N_9159,N_6248,N_6278);
or U9160 (N_9160,N_7682,N_6191);
and U9161 (N_9161,N_7564,N_7820);
nor U9162 (N_9162,N_6821,N_6842);
nor U9163 (N_9163,N_7487,N_6585);
nor U9164 (N_9164,N_6843,N_6253);
nor U9165 (N_9165,N_7638,N_6490);
nor U9166 (N_9166,N_6929,N_6936);
nand U9167 (N_9167,N_7016,N_6273);
or U9168 (N_9168,N_6516,N_7535);
and U9169 (N_9169,N_6918,N_7901);
nand U9170 (N_9170,N_7701,N_7294);
or U9171 (N_9171,N_6894,N_6726);
nor U9172 (N_9172,N_6293,N_7540);
xnor U9173 (N_9173,N_6850,N_6246);
nor U9174 (N_9174,N_7077,N_7668);
or U9175 (N_9175,N_6947,N_6523);
nand U9176 (N_9176,N_7041,N_6739);
and U9177 (N_9177,N_7332,N_6405);
nor U9178 (N_9178,N_7604,N_7252);
or U9179 (N_9179,N_7807,N_6313);
nor U9180 (N_9180,N_7033,N_7208);
and U9181 (N_9181,N_6076,N_7159);
nand U9182 (N_9182,N_7997,N_7839);
and U9183 (N_9183,N_7529,N_6587);
nor U9184 (N_9184,N_6766,N_6909);
nand U9185 (N_9185,N_7405,N_7578);
nor U9186 (N_9186,N_7371,N_6738);
nand U9187 (N_9187,N_6851,N_7933);
nor U9188 (N_9188,N_7558,N_6973);
or U9189 (N_9189,N_7586,N_7949);
nor U9190 (N_9190,N_7796,N_7299);
and U9191 (N_9191,N_7925,N_7100);
or U9192 (N_9192,N_7893,N_6126);
nor U9193 (N_9193,N_6971,N_6223);
nand U9194 (N_9194,N_6767,N_6807);
nor U9195 (N_9195,N_7867,N_7713);
nor U9196 (N_9196,N_7731,N_6926);
or U9197 (N_9197,N_6222,N_7830);
and U9198 (N_9198,N_7803,N_7722);
nor U9199 (N_9199,N_7170,N_6048);
nand U9200 (N_9200,N_6007,N_7328);
nand U9201 (N_9201,N_7841,N_7871);
or U9202 (N_9202,N_7172,N_7081);
or U9203 (N_9203,N_7991,N_6290);
nand U9204 (N_9204,N_7474,N_7740);
nor U9205 (N_9205,N_7906,N_7610);
nand U9206 (N_9206,N_6618,N_6002);
nor U9207 (N_9207,N_7229,N_6572);
or U9208 (N_9208,N_7155,N_7592);
xnor U9209 (N_9209,N_7164,N_6653);
nand U9210 (N_9210,N_6455,N_7883);
nor U9211 (N_9211,N_6101,N_7628);
or U9212 (N_9212,N_6216,N_7964);
and U9213 (N_9213,N_6482,N_7865);
or U9214 (N_9214,N_6078,N_7500);
nor U9215 (N_9215,N_6173,N_7107);
nor U9216 (N_9216,N_6905,N_6613);
or U9217 (N_9217,N_7626,N_6283);
nand U9218 (N_9218,N_6731,N_7679);
and U9219 (N_9219,N_6266,N_6594);
or U9220 (N_9220,N_6063,N_7158);
nand U9221 (N_9221,N_7868,N_7348);
or U9222 (N_9222,N_6584,N_7935);
and U9223 (N_9223,N_6188,N_6552);
nand U9224 (N_9224,N_7931,N_7137);
and U9225 (N_9225,N_7110,N_7568);
nor U9226 (N_9226,N_7339,N_6136);
nor U9227 (N_9227,N_6362,N_7650);
or U9228 (N_9228,N_7167,N_6471);
nand U9229 (N_9229,N_6200,N_6564);
nor U9230 (N_9230,N_7679,N_6348);
and U9231 (N_9231,N_6075,N_6724);
and U9232 (N_9232,N_6537,N_6626);
and U9233 (N_9233,N_7736,N_7638);
and U9234 (N_9234,N_7140,N_6637);
and U9235 (N_9235,N_7970,N_6498);
nand U9236 (N_9236,N_7083,N_7696);
or U9237 (N_9237,N_6803,N_7822);
or U9238 (N_9238,N_7880,N_6392);
nand U9239 (N_9239,N_7216,N_6425);
xor U9240 (N_9240,N_7481,N_7312);
or U9241 (N_9241,N_7813,N_7594);
nand U9242 (N_9242,N_7502,N_7891);
nor U9243 (N_9243,N_7440,N_6237);
and U9244 (N_9244,N_6816,N_7686);
or U9245 (N_9245,N_6343,N_6371);
and U9246 (N_9246,N_7167,N_7355);
xnor U9247 (N_9247,N_7002,N_6021);
or U9248 (N_9248,N_6858,N_6143);
nor U9249 (N_9249,N_7645,N_6084);
nor U9250 (N_9250,N_7763,N_6189);
xnor U9251 (N_9251,N_6564,N_6532);
or U9252 (N_9252,N_7822,N_7996);
nand U9253 (N_9253,N_7994,N_6744);
nand U9254 (N_9254,N_7348,N_6417);
or U9255 (N_9255,N_7355,N_7252);
nand U9256 (N_9256,N_6708,N_6014);
nand U9257 (N_9257,N_7495,N_7271);
and U9258 (N_9258,N_6567,N_7717);
nand U9259 (N_9259,N_7947,N_7481);
or U9260 (N_9260,N_7449,N_7838);
nand U9261 (N_9261,N_6397,N_6512);
nor U9262 (N_9262,N_7229,N_6193);
nand U9263 (N_9263,N_7144,N_7237);
nand U9264 (N_9264,N_6768,N_7350);
nor U9265 (N_9265,N_6874,N_7121);
nor U9266 (N_9266,N_7517,N_6695);
and U9267 (N_9267,N_6682,N_6466);
nand U9268 (N_9268,N_7752,N_7318);
or U9269 (N_9269,N_7644,N_6714);
or U9270 (N_9270,N_6909,N_7825);
nor U9271 (N_9271,N_7225,N_6235);
or U9272 (N_9272,N_6418,N_6541);
and U9273 (N_9273,N_7315,N_6398);
and U9274 (N_9274,N_7026,N_7301);
and U9275 (N_9275,N_7077,N_6105);
and U9276 (N_9276,N_6751,N_7087);
nor U9277 (N_9277,N_6497,N_6832);
nor U9278 (N_9278,N_7567,N_6816);
nor U9279 (N_9279,N_6537,N_6817);
and U9280 (N_9280,N_7487,N_6687);
nor U9281 (N_9281,N_7291,N_6755);
or U9282 (N_9282,N_7512,N_7135);
nand U9283 (N_9283,N_6209,N_6728);
xor U9284 (N_9284,N_7580,N_7624);
nand U9285 (N_9285,N_7513,N_7464);
nor U9286 (N_9286,N_6215,N_7323);
nor U9287 (N_9287,N_7403,N_7827);
nand U9288 (N_9288,N_7244,N_6910);
nor U9289 (N_9289,N_6164,N_7097);
nand U9290 (N_9290,N_7992,N_6697);
or U9291 (N_9291,N_6552,N_6702);
and U9292 (N_9292,N_6724,N_6004);
nand U9293 (N_9293,N_6448,N_7012);
nor U9294 (N_9294,N_7985,N_6066);
or U9295 (N_9295,N_7312,N_6546);
nor U9296 (N_9296,N_6188,N_7032);
or U9297 (N_9297,N_7443,N_7064);
and U9298 (N_9298,N_6542,N_6072);
or U9299 (N_9299,N_7031,N_7482);
nand U9300 (N_9300,N_6591,N_7702);
or U9301 (N_9301,N_7155,N_7404);
or U9302 (N_9302,N_7987,N_7114);
or U9303 (N_9303,N_7741,N_6621);
and U9304 (N_9304,N_6568,N_6373);
nand U9305 (N_9305,N_7161,N_6210);
nor U9306 (N_9306,N_7200,N_6371);
or U9307 (N_9307,N_7175,N_6319);
and U9308 (N_9308,N_7074,N_6927);
xor U9309 (N_9309,N_7048,N_6558);
or U9310 (N_9310,N_6779,N_6500);
and U9311 (N_9311,N_7166,N_7933);
nor U9312 (N_9312,N_7415,N_7193);
nor U9313 (N_9313,N_6796,N_6557);
and U9314 (N_9314,N_6908,N_7563);
or U9315 (N_9315,N_6250,N_7595);
or U9316 (N_9316,N_7068,N_6613);
nor U9317 (N_9317,N_6166,N_6370);
nor U9318 (N_9318,N_7585,N_7022);
nand U9319 (N_9319,N_7414,N_7568);
nor U9320 (N_9320,N_6123,N_7124);
or U9321 (N_9321,N_7162,N_7491);
or U9322 (N_9322,N_6192,N_6441);
nand U9323 (N_9323,N_6250,N_6520);
nand U9324 (N_9324,N_6034,N_7052);
nand U9325 (N_9325,N_6606,N_7024);
nand U9326 (N_9326,N_7165,N_6754);
or U9327 (N_9327,N_6864,N_6551);
nor U9328 (N_9328,N_6894,N_6584);
and U9329 (N_9329,N_6916,N_7516);
or U9330 (N_9330,N_6090,N_7349);
and U9331 (N_9331,N_7871,N_7316);
and U9332 (N_9332,N_6771,N_6186);
or U9333 (N_9333,N_7785,N_7510);
and U9334 (N_9334,N_7913,N_6981);
and U9335 (N_9335,N_6562,N_7128);
nand U9336 (N_9336,N_7563,N_6730);
nor U9337 (N_9337,N_7784,N_7903);
nor U9338 (N_9338,N_7038,N_6393);
nor U9339 (N_9339,N_6216,N_7318);
nand U9340 (N_9340,N_6585,N_7843);
or U9341 (N_9341,N_7383,N_7918);
and U9342 (N_9342,N_6962,N_6761);
nor U9343 (N_9343,N_6479,N_6544);
nor U9344 (N_9344,N_6419,N_6459);
and U9345 (N_9345,N_7069,N_6994);
and U9346 (N_9346,N_7289,N_7778);
and U9347 (N_9347,N_6853,N_7729);
nand U9348 (N_9348,N_6378,N_6106);
nor U9349 (N_9349,N_6561,N_6245);
or U9350 (N_9350,N_6923,N_6486);
nor U9351 (N_9351,N_6441,N_7820);
and U9352 (N_9352,N_7215,N_7784);
and U9353 (N_9353,N_7338,N_7895);
nand U9354 (N_9354,N_6241,N_6054);
nor U9355 (N_9355,N_7325,N_7915);
nor U9356 (N_9356,N_6690,N_6548);
nand U9357 (N_9357,N_6710,N_6058);
nor U9358 (N_9358,N_6390,N_6238);
and U9359 (N_9359,N_7322,N_6106);
nor U9360 (N_9360,N_7937,N_7834);
and U9361 (N_9361,N_6102,N_7878);
nor U9362 (N_9362,N_6878,N_7299);
or U9363 (N_9363,N_7574,N_7550);
or U9364 (N_9364,N_7987,N_7310);
nor U9365 (N_9365,N_7219,N_6190);
and U9366 (N_9366,N_6006,N_6845);
nand U9367 (N_9367,N_6308,N_6248);
or U9368 (N_9368,N_6031,N_7137);
or U9369 (N_9369,N_7789,N_6287);
nand U9370 (N_9370,N_7704,N_6955);
nand U9371 (N_9371,N_7143,N_6861);
or U9372 (N_9372,N_6885,N_6150);
or U9373 (N_9373,N_6779,N_6073);
or U9374 (N_9374,N_7719,N_7396);
or U9375 (N_9375,N_7786,N_6890);
and U9376 (N_9376,N_6805,N_7208);
nor U9377 (N_9377,N_6661,N_6008);
or U9378 (N_9378,N_7808,N_6741);
nand U9379 (N_9379,N_6950,N_7748);
and U9380 (N_9380,N_6479,N_6692);
nand U9381 (N_9381,N_7058,N_6143);
nor U9382 (N_9382,N_6721,N_6493);
nand U9383 (N_9383,N_7469,N_7389);
and U9384 (N_9384,N_7429,N_7956);
or U9385 (N_9385,N_7442,N_7536);
and U9386 (N_9386,N_7777,N_7259);
or U9387 (N_9387,N_6366,N_7661);
nand U9388 (N_9388,N_6295,N_6468);
nand U9389 (N_9389,N_6785,N_6248);
nand U9390 (N_9390,N_6851,N_7236);
and U9391 (N_9391,N_7638,N_7762);
nand U9392 (N_9392,N_7179,N_6455);
and U9393 (N_9393,N_7917,N_7165);
or U9394 (N_9394,N_6493,N_7910);
nor U9395 (N_9395,N_6391,N_7126);
and U9396 (N_9396,N_6908,N_6012);
nand U9397 (N_9397,N_6398,N_7891);
or U9398 (N_9398,N_7053,N_6185);
or U9399 (N_9399,N_7218,N_6500);
nand U9400 (N_9400,N_7030,N_6336);
xnor U9401 (N_9401,N_7460,N_7610);
nand U9402 (N_9402,N_7761,N_7734);
nor U9403 (N_9403,N_6520,N_7725);
nand U9404 (N_9404,N_7362,N_7093);
and U9405 (N_9405,N_7542,N_7735);
nor U9406 (N_9406,N_7180,N_6834);
or U9407 (N_9407,N_6027,N_7101);
or U9408 (N_9408,N_7755,N_6165);
nand U9409 (N_9409,N_7298,N_6684);
and U9410 (N_9410,N_7330,N_6452);
nor U9411 (N_9411,N_6602,N_6003);
and U9412 (N_9412,N_7471,N_7101);
nor U9413 (N_9413,N_7433,N_6070);
xor U9414 (N_9414,N_7911,N_6844);
or U9415 (N_9415,N_6975,N_6884);
or U9416 (N_9416,N_7264,N_6104);
nand U9417 (N_9417,N_6214,N_6269);
or U9418 (N_9418,N_7195,N_6005);
or U9419 (N_9419,N_6529,N_6313);
or U9420 (N_9420,N_6559,N_7799);
and U9421 (N_9421,N_6218,N_7134);
xor U9422 (N_9422,N_7368,N_6257);
nand U9423 (N_9423,N_7968,N_6624);
and U9424 (N_9424,N_6031,N_7299);
nor U9425 (N_9425,N_6856,N_7887);
or U9426 (N_9426,N_6921,N_6952);
and U9427 (N_9427,N_7209,N_6036);
nor U9428 (N_9428,N_7617,N_7419);
and U9429 (N_9429,N_6457,N_6361);
or U9430 (N_9430,N_7364,N_7045);
or U9431 (N_9431,N_6696,N_6641);
nor U9432 (N_9432,N_6779,N_6829);
or U9433 (N_9433,N_7858,N_6979);
nand U9434 (N_9434,N_7395,N_6279);
nor U9435 (N_9435,N_7778,N_7321);
nor U9436 (N_9436,N_6447,N_6938);
and U9437 (N_9437,N_7580,N_6013);
nand U9438 (N_9438,N_7241,N_7047);
nor U9439 (N_9439,N_7515,N_6623);
or U9440 (N_9440,N_7700,N_6825);
nand U9441 (N_9441,N_7718,N_7584);
nand U9442 (N_9442,N_6698,N_6094);
or U9443 (N_9443,N_6657,N_6970);
nor U9444 (N_9444,N_6263,N_7009);
or U9445 (N_9445,N_7386,N_6476);
nor U9446 (N_9446,N_6538,N_6006);
nand U9447 (N_9447,N_6343,N_7466);
nor U9448 (N_9448,N_6605,N_6033);
nor U9449 (N_9449,N_6614,N_6680);
and U9450 (N_9450,N_7556,N_7577);
or U9451 (N_9451,N_7852,N_7549);
or U9452 (N_9452,N_6570,N_6731);
and U9453 (N_9453,N_7533,N_6180);
and U9454 (N_9454,N_6346,N_7489);
and U9455 (N_9455,N_7517,N_6230);
nor U9456 (N_9456,N_6196,N_6136);
nor U9457 (N_9457,N_7743,N_6323);
or U9458 (N_9458,N_7875,N_7045);
or U9459 (N_9459,N_6693,N_7402);
xnor U9460 (N_9460,N_6039,N_6878);
and U9461 (N_9461,N_7358,N_7252);
and U9462 (N_9462,N_7189,N_6343);
or U9463 (N_9463,N_7733,N_7161);
or U9464 (N_9464,N_7663,N_7192);
nor U9465 (N_9465,N_7834,N_6991);
nand U9466 (N_9466,N_7897,N_6117);
or U9467 (N_9467,N_7518,N_7516);
nor U9468 (N_9468,N_7960,N_7629);
or U9469 (N_9469,N_6578,N_7796);
nand U9470 (N_9470,N_6960,N_7645);
nand U9471 (N_9471,N_7898,N_6259);
nand U9472 (N_9472,N_7372,N_6187);
nand U9473 (N_9473,N_6648,N_6514);
or U9474 (N_9474,N_7431,N_7329);
nand U9475 (N_9475,N_6687,N_7859);
and U9476 (N_9476,N_7421,N_6862);
nor U9477 (N_9477,N_7452,N_6055);
and U9478 (N_9478,N_6635,N_7512);
or U9479 (N_9479,N_7224,N_7005);
or U9480 (N_9480,N_6055,N_7489);
and U9481 (N_9481,N_7420,N_7848);
or U9482 (N_9482,N_6038,N_7268);
nor U9483 (N_9483,N_7731,N_7819);
nor U9484 (N_9484,N_6384,N_6783);
nand U9485 (N_9485,N_7276,N_7361);
or U9486 (N_9486,N_6039,N_6988);
or U9487 (N_9487,N_6479,N_7768);
nand U9488 (N_9488,N_7517,N_7909);
or U9489 (N_9489,N_7549,N_6839);
nor U9490 (N_9490,N_7542,N_7877);
or U9491 (N_9491,N_6253,N_6809);
nand U9492 (N_9492,N_6730,N_7125);
nor U9493 (N_9493,N_7812,N_7344);
and U9494 (N_9494,N_7373,N_6936);
nand U9495 (N_9495,N_7556,N_6163);
or U9496 (N_9496,N_7903,N_7675);
and U9497 (N_9497,N_6829,N_6496);
or U9498 (N_9498,N_7218,N_6964);
nor U9499 (N_9499,N_6246,N_6047);
and U9500 (N_9500,N_7567,N_6680);
nand U9501 (N_9501,N_6384,N_6546);
nor U9502 (N_9502,N_6913,N_6245);
and U9503 (N_9503,N_7996,N_7884);
nand U9504 (N_9504,N_6338,N_6669);
nor U9505 (N_9505,N_6222,N_6157);
nor U9506 (N_9506,N_7798,N_6316);
and U9507 (N_9507,N_7141,N_7709);
or U9508 (N_9508,N_6248,N_6688);
and U9509 (N_9509,N_7610,N_6692);
nand U9510 (N_9510,N_6268,N_6317);
and U9511 (N_9511,N_7815,N_7847);
nand U9512 (N_9512,N_6889,N_7881);
or U9513 (N_9513,N_6908,N_7680);
and U9514 (N_9514,N_6182,N_6856);
nor U9515 (N_9515,N_6977,N_6347);
and U9516 (N_9516,N_6987,N_6906);
or U9517 (N_9517,N_7079,N_7094);
nand U9518 (N_9518,N_6492,N_7339);
or U9519 (N_9519,N_7285,N_7331);
and U9520 (N_9520,N_6119,N_7020);
nand U9521 (N_9521,N_6059,N_7470);
and U9522 (N_9522,N_6135,N_7417);
nand U9523 (N_9523,N_7469,N_7674);
nand U9524 (N_9524,N_7626,N_6537);
and U9525 (N_9525,N_7094,N_7674);
and U9526 (N_9526,N_7724,N_6263);
nor U9527 (N_9527,N_7805,N_7885);
nor U9528 (N_9528,N_7985,N_7879);
xor U9529 (N_9529,N_7991,N_7222);
nor U9530 (N_9530,N_6970,N_7016);
xnor U9531 (N_9531,N_7626,N_6207);
nor U9532 (N_9532,N_7819,N_6273);
nor U9533 (N_9533,N_7703,N_7224);
nor U9534 (N_9534,N_7845,N_6198);
nand U9535 (N_9535,N_6580,N_7614);
nand U9536 (N_9536,N_7651,N_7963);
and U9537 (N_9537,N_6285,N_7543);
or U9538 (N_9538,N_6976,N_7070);
or U9539 (N_9539,N_6341,N_7286);
and U9540 (N_9540,N_6558,N_7671);
or U9541 (N_9541,N_7013,N_7919);
xnor U9542 (N_9542,N_7983,N_7057);
and U9543 (N_9543,N_7620,N_6594);
nand U9544 (N_9544,N_6006,N_7422);
and U9545 (N_9545,N_6426,N_7343);
nor U9546 (N_9546,N_7266,N_7269);
nor U9547 (N_9547,N_7511,N_6886);
and U9548 (N_9548,N_7685,N_7190);
and U9549 (N_9549,N_6234,N_7348);
or U9550 (N_9550,N_7269,N_6631);
nor U9551 (N_9551,N_6142,N_7209);
and U9552 (N_9552,N_7561,N_7424);
or U9553 (N_9553,N_6559,N_7406);
or U9554 (N_9554,N_6897,N_7290);
nand U9555 (N_9555,N_7177,N_6667);
nor U9556 (N_9556,N_6238,N_6855);
xor U9557 (N_9557,N_6487,N_6287);
or U9558 (N_9558,N_7697,N_6098);
and U9559 (N_9559,N_6758,N_6519);
nor U9560 (N_9560,N_6321,N_7521);
nand U9561 (N_9561,N_7556,N_6564);
xnor U9562 (N_9562,N_7790,N_7050);
or U9563 (N_9563,N_7989,N_7752);
nand U9564 (N_9564,N_7686,N_6267);
or U9565 (N_9565,N_7843,N_6267);
nand U9566 (N_9566,N_6017,N_6678);
or U9567 (N_9567,N_6053,N_7368);
nand U9568 (N_9568,N_7122,N_6939);
and U9569 (N_9569,N_6163,N_7278);
and U9570 (N_9570,N_7525,N_7385);
nor U9571 (N_9571,N_6733,N_6343);
nor U9572 (N_9572,N_6809,N_7529);
nor U9573 (N_9573,N_6987,N_7859);
nand U9574 (N_9574,N_6776,N_6205);
nand U9575 (N_9575,N_7058,N_6867);
nand U9576 (N_9576,N_6129,N_6602);
nand U9577 (N_9577,N_6684,N_7064);
nor U9578 (N_9578,N_7910,N_7991);
nand U9579 (N_9579,N_7131,N_6529);
nor U9580 (N_9580,N_6413,N_7276);
nand U9581 (N_9581,N_7292,N_7347);
nand U9582 (N_9582,N_7972,N_6072);
and U9583 (N_9583,N_7488,N_6517);
nor U9584 (N_9584,N_7582,N_6728);
nand U9585 (N_9585,N_6820,N_6150);
nor U9586 (N_9586,N_7412,N_6070);
and U9587 (N_9587,N_6169,N_7777);
nand U9588 (N_9588,N_6554,N_7234);
or U9589 (N_9589,N_6248,N_6526);
nand U9590 (N_9590,N_7870,N_6232);
nor U9591 (N_9591,N_6950,N_6786);
nor U9592 (N_9592,N_7314,N_6280);
and U9593 (N_9593,N_6696,N_7518);
nor U9594 (N_9594,N_7312,N_6555);
nor U9595 (N_9595,N_6135,N_6188);
xor U9596 (N_9596,N_7928,N_6353);
and U9597 (N_9597,N_7005,N_7448);
or U9598 (N_9598,N_6182,N_6537);
nand U9599 (N_9599,N_6346,N_7930);
xor U9600 (N_9600,N_7211,N_7131);
and U9601 (N_9601,N_7026,N_7856);
nor U9602 (N_9602,N_6197,N_6184);
nor U9603 (N_9603,N_7362,N_7769);
nor U9604 (N_9604,N_7152,N_7833);
nand U9605 (N_9605,N_7855,N_6185);
or U9606 (N_9606,N_6965,N_6371);
nor U9607 (N_9607,N_7174,N_6981);
nor U9608 (N_9608,N_7084,N_7907);
or U9609 (N_9609,N_7072,N_7486);
nand U9610 (N_9610,N_6427,N_6111);
or U9611 (N_9611,N_7473,N_6197);
nor U9612 (N_9612,N_6145,N_7851);
and U9613 (N_9613,N_7247,N_6172);
or U9614 (N_9614,N_6276,N_6257);
nor U9615 (N_9615,N_7776,N_6960);
xnor U9616 (N_9616,N_7599,N_7353);
nor U9617 (N_9617,N_6701,N_7328);
nand U9618 (N_9618,N_6517,N_7901);
nand U9619 (N_9619,N_6223,N_7320);
nor U9620 (N_9620,N_7175,N_7258);
and U9621 (N_9621,N_6226,N_6642);
nand U9622 (N_9622,N_6570,N_6406);
nand U9623 (N_9623,N_7777,N_7854);
and U9624 (N_9624,N_7880,N_6002);
or U9625 (N_9625,N_7325,N_6113);
or U9626 (N_9626,N_6406,N_6478);
and U9627 (N_9627,N_6248,N_6340);
nand U9628 (N_9628,N_6074,N_6648);
and U9629 (N_9629,N_6451,N_6208);
xnor U9630 (N_9630,N_7122,N_6203);
nor U9631 (N_9631,N_7084,N_7522);
and U9632 (N_9632,N_6070,N_6302);
nand U9633 (N_9633,N_7378,N_7939);
nor U9634 (N_9634,N_6276,N_6987);
or U9635 (N_9635,N_6105,N_6587);
and U9636 (N_9636,N_6612,N_7185);
nand U9637 (N_9637,N_7557,N_7769);
or U9638 (N_9638,N_7418,N_6357);
nor U9639 (N_9639,N_7950,N_7669);
or U9640 (N_9640,N_7293,N_6123);
and U9641 (N_9641,N_6396,N_6269);
nand U9642 (N_9642,N_7852,N_7189);
nand U9643 (N_9643,N_6688,N_6588);
nor U9644 (N_9644,N_6842,N_6671);
and U9645 (N_9645,N_7721,N_6848);
and U9646 (N_9646,N_7448,N_6924);
or U9647 (N_9647,N_7206,N_7910);
and U9648 (N_9648,N_7241,N_6190);
or U9649 (N_9649,N_6432,N_7991);
or U9650 (N_9650,N_6095,N_6476);
xor U9651 (N_9651,N_7342,N_7062);
and U9652 (N_9652,N_6660,N_7509);
nor U9653 (N_9653,N_6422,N_6618);
or U9654 (N_9654,N_6889,N_6461);
and U9655 (N_9655,N_6664,N_7957);
nand U9656 (N_9656,N_7689,N_6078);
or U9657 (N_9657,N_7380,N_6755);
nor U9658 (N_9658,N_6135,N_6832);
or U9659 (N_9659,N_7431,N_7883);
or U9660 (N_9660,N_7002,N_7303);
nor U9661 (N_9661,N_6522,N_6177);
and U9662 (N_9662,N_6548,N_7743);
or U9663 (N_9663,N_7144,N_6497);
or U9664 (N_9664,N_6781,N_6739);
or U9665 (N_9665,N_6428,N_7344);
or U9666 (N_9666,N_7189,N_7566);
and U9667 (N_9667,N_6707,N_7679);
or U9668 (N_9668,N_6083,N_6586);
or U9669 (N_9669,N_7786,N_7021);
or U9670 (N_9670,N_6625,N_6851);
nand U9671 (N_9671,N_6414,N_6671);
xor U9672 (N_9672,N_6738,N_7366);
and U9673 (N_9673,N_6339,N_6613);
and U9674 (N_9674,N_7380,N_6896);
and U9675 (N_9675,N_6613,N_7831);
nand U9676 (N_9676,N_6914,N_6700);
nor U9677 (N_9677,N_6783,N_7830);
or U9678 (N_9678,N_7790,N_6965);
nor U9679 (N_9679,N_6270,N_6978);
and U9680 (N_9680,N_7060,N_7445);
nor U9681 (N_9681,N_6448,N_6427);
nand U9682 (N_9682,N_7943,N_6140);
or U9683 (N_9683,N_6069,N_6792);
nand U9684 (N_9684,N_7503,N_6204);
and U9685 (N_9685,N_6155,N_6995);
nor U9686 (N_9686,N_7667,N_7159);
nand U9687 (N_9687,N_7803,N_6121);
nor U9688 (N_9688,N_7858,N_7869);
nor U9689 (N_9689,N_7162,N_6258);
nand U9690 (N_9690,N_6242,N_6985);
or U9691 (N_9691,N_7608,N_7167);
and U9692 (N_9692,N_6067,N_6347);
xor U9693 (N_9693,N_7496,N_6836);
and U9694 (N_9694,N_6075,N_7866);
nor U9695 (N_9695,N_7764,N_7630);
nand U9696 (N_9696,N_6605,N_7953);
nor U9697 (N_9697,N_6316,N_6297);
and U9698 (N_9698,N_7427,N_7901);
nand U9699 (N_9699,N_7247,N_7793);
nand U9700 (N_9700,N_6644,N_7808);
and U9701 (N_9701,N_6361,N_7849);
or U9702 (N_9702,N_7331,N_7376);
or U9703 (N_9703,N_6916,N_7369);
nor U9704 (N_9704,N_6785,N_7857);
nor U9705 (N_9705,N_6088,N_6708);
and U9706 (N_9706,N_6006,N_6715);
or U9707 (N_9707,N_7805,N_7329);
nor U9708 (N_9708,N_7897,N_6769);
and U9709 (N_9709,N_6021,N_6074);
and U9710 (N_9710,N_6704,N_7285);
and U9711 (N_9711,N_6219,N_6916);
nand U9712 (N_9712,N_6400,N_6933);
or U9713 (N_9713,N_6299,N_7365);
and U9714 (N_9714,N_6829,N_7255);
nor U9715 (N_9715,N_6461,N_7528);
and U9716 (N_9716,N_6302,N_6145);
nor U9717 (N_9717,N_7149,N_7441);
or U9718 (N_9718,N_7181,N_6024);
nor U9719 (N_9719,N_6688,N_7014);
nor U9720 (N_9720,N_7944,N_7770);
xor U9721 (N_9721,N_6202,N_7469);
or U9722 (N_9722,N_7109,N_6654);
nand U9723 (N_9723,N_6763,N_7619);
or U9724 (N_9724,N_6131,N_7763);
nand U9725 (N_9725,N_6220,N_7135);
nand U9726 (N_9726,N_7599,N_6898);
or U9727 (N_9727,N_7179,N_7365);
and U9728 (N_9728,N_6518,N_6849);
and U9729 (N_9729,N_6581,N_7742);
nand U9730 (N_9730,N_7733,N_6572);
xor U9731 (N_9731,N_7138,N_6497);
or U9732 (N_9732,N_7934,N_6870);
and U9733 (N_9733,N_6530,N_6988);
nand U9734 (N_9734,N_6757,N_7288);
nor U9735 (N_9735,N_7386,N_7318);
or U9736 (N_9736,N_7618,N_7195);
nand U9737 (N_9737,N_6109,N_7833);
and U9738 (N_9738,N_6228,N_7095);
nor U9739 (N_9739,N_6928,N_7980);
nor U9740 (N_9740,N_6298,N_7524);
nor U9741 (N_9741,N_7373,N_7454);
nor U9742 (N_9742,N_7066,N_7841);
or U9743 (N_9743,N_7076,N_6595);
or U9744 (N_9744,N_7804,N_6897);
and U9745 (N_9745,N_6856,N_7199);
nor U9746 (N_9746,N_6303,N_6960);
or U9747 (N_9747,N_7595,N_7551);
nand U9748 (N_9748,N_7824,N_6918);
nand U9749 (N_9749,N_6676,N_6347);
or U9750 (N_9750,N_7954,N_6113);
and U9751 (N_9751,N_6120,N_6546);
nor U9752 (N_9752,N_7715,N_6491);
nor U9753 (N_9753,N_7853,N_6789);
and U9754 (N_9754,N_7305,N_7999);
nand U9755 (N_9755,N_7630,N_7809);
nor U9756 (N_9756,N_6924,N_6851);
or U9757 (N_9757,N_6366,N_7466);
nand U9758 (N_9758,N_7549,N_6665);
and U9759 (N_9759,N_6814,N_6431);
or U9760 (N_9760,N_6554,N_6184);
nor U9761 (N_9761,N_7781,N_6197);
or U9762 (N_9762,N_7503,N_7831);
or U9763 (N_9763,N_6938,N_7886);
and U9764 (N_9764,N_7567,N_6993);
or U9765 (N_9765,N_7008,N_6597);
nand U9766 (N_9766,N_7635,N_7273);
xor U9767 (N_9767,N_7575,N_6571);
nor U9768 (N_9768,N_7022,N_6915);
nor U9769 (N_9769,N_7614,N_6890);
and U9770 (N_9770,N_7433,N_6476);
nand U9771 (N_9771,N_6761,N_7482);
nor U9772 (N_9772,N_6235,N_6038);
nor U9773 (N_9773,N_7454,N_6127);
nand U9774 (N_9774,N_6646,N_7362);
nand U9775 (N_9775,N_6940,N_6716);
nand U9776 (N_9776,N_7475,N_6865);
and U9777 (N_9777,N_6117,N_6628);
or U9778 (N_9778,N_7237,N_6303);
or U9779 (N_9779,N_6050,N_7853);
nand U9780 (N_9780,N_7652,N_6987);
or U9781 (N_9781,N_6801,N_6892);
and U9782 (N_9782,N_7801,N_6213);
nor U9783 (N_9783,N_6188,N_7840);
nor U9784 (N_9784,N_6342,N_6260);
and U9785 (N_9785,N_7940,N_6636);
nand U9786 (N_9786,N_7246,N_7060);
nand U9787 (N_9787,N_6159,N_6802);
nor U9788 (N_9788,N_7766,N_6406);
or U9789 (N_9789,N_7956,N_7331);
and U9790 (N_9790,N_7592,N_7654);
nand U9791 (N_9791,N_6472,N_7760);
nand U9792 (N_9792,N_6681,N_6162);
nand U9793 (N_9793,N_6188,N_6979);
nand U9794 (N_9794,N_6063,N_6120);
nand U9795 (N_9795,N_7616,N_6764);
nand U9796 (N_9796,N_6261,N_6212);
nor U9797 (N_9797,N_6403,N_7525);
nor U9798 (N_9798,N_7985,N_6828);
nor U9799 (N_9799,N_6562,N_7894);
xnor U9800 (N_9800,N_6684,N_7653);
and U9801 (N_9801,N_7777,N_7132);
or U9802 (N_9802,N_7378,N_6072);
or U9803 (N_9803,N_6426,N_6657);
and U9804 (N_9804,N_6510,N_7929);
and U9805 (N_9805,N_6353,N_6786);
xor U9806 (N_9806,N_7341,N_6265);
nor U9807 (N_9807,N_7981,N_7361);
nor U9808 (N_9808,N_6672,N_6907);
and U9809 (N_9809,N_6588,N_6855);
and U9810 (N_9810,N_7674,N_6345);
or U9811 (N_9811,N_6960,N_6085);
or U9812 (N_9812,N_6018,N_6758);
nor U9813 (N_9813,N_7206,N_7923);
nand U9814 (N_9814,N_7396,N_7706);
and U9815 (N_9815,N_7665,N_6778);
and U9816 (N_9816,N_7674,N_7464);
and U9817 (N_9817,N_6758,N_6608);
or U9818 (N_9818,N_6429,N_6094);
or U9819 (N_9819,N_7621,N_7706);
and U9820 (N_9820,N_7793,N_7105);
and U9821 (N_9821,N_7411,N_6588);
or U9822 (N_9822,N_7389,N_7682);
or U9823 (N_9823,N_7705,N_6427);
nor U9824 (N_9824,N_7154,N_7400);
or U9825 (N_9825,N_6903,N_6428);
nand U9826 (N_9826,N_7939,N_7209);
nand U9827 (N_9827,N_6235,N_6924);
and U9828 (N_9828,N_7812,N_6393);
or U9829 (N_9829,N_7345,N_6174);
or U9830 (N_9830,N_6449,N_7710);
nor U9831 (N_9831,N_7152,N_6010);
or U9832 (N_9832,N_7891,N_6399);
or U9833 (N_9833,N_7291,N_7616);
or U9834 (N_9834,N_7793,N_6639);
or U9835 (N_9835,N_6212,N_6195);
and U9836 (N_9836,N_6658,N_7666);
or U9837 (N_9837,N_6796,N_6716);
nor U9838 (N_9838,N_7943,N_6793);
or U9839 (N_9839,N_7497,N_7118);
and U9840 (N_9840,N_7475,N_6574);
or U9841 (N_9841,N_7990,N_7876);
nand U9842 (N_9842,N_7557,N_7932);
nor U9843 (N_9843,N_7217,N_6121);
nor U9844 (N_9844,N_6602,N_6725);
or U9845 (N_9845,N_7760,N_7510);
and U9846 (N_9846,N_7364,N_7717);
and U9847 (N_9847,N_6328,N_6678);
nand U9848 (N_9848,N_7145,N_7357);
nand U9849 (N_9849,N_6303,N_7072);
or U9850 (N_9850,N_6256,N_6697);
nand U9851 (N_9851,N_7346,N_7135);
nor U9852 (N_9852,N_7348,N_7990);
nor U9853 (N_9853,N_6138,N_6264);
nand U9854 (N_9854,N_6177,N_6360);
nand U9855 (N_9855,N_6347,N_6053);
or U9856 (N_9856,N_7315,N_6307);
nor U9857 (N_9857,N_6411,N_7933);
nor U9858 (N_9858,N_6839,N_7405);
nor U9859 (N_9859,N_7487,N_6671);
and U9860 (N_9860,N_7924,N_7642);
or U9861 (N_9861,N_6390,N_6412);
nor U9862 (N_9862,N_7341,N_7332);
and U9863 (N_9863,N_6666,N_6972);
nor U9864 (N_9864,N_6269,N_7693);
nor U9865 (N_9865,N_7063,N_6993);
nor U9866 (N_9866,N_7162,N_7094);
and U9867 (N_9867,N_6451,N_7676);
and U9868 (N_9868,N_6764,N_6869);
and U9869 (N_9869,N_7178,N_6881);
nand U9870 (N_9870,N_7464,N_6123);
nand U9871 (N_9871,N_7203,N_7543);
nand U9872 (N_9872,N_6827,N_6951);
and U9873 (N_9873,N_6389,N_6437);
or U9874 (N_9874,N_7985,N_6227);
or U9875 (N_9875,N_6656,N_6717);
or U9876 (N_9876,N_6241,N_7139);
nor U9877 (N_9877,N_7584,N_7005);
and U9878 (N_9878,N_7066,N_7527);
or U9879 (N_9879,N_6763,N_6006);
and U9880 (N_9880,N_7783,N_6236);
nand U9881 (N_9881,N_6743,N_6285);
and U9882 (N_9882,N_7674,N_6851);
and U9883 (N_9883,N_6978,N_7546);
nand U9884 (N_9884,N_6289,N_7711);
nand U9885 (N_9885,N_6124,N_6395);
or U9886 (N_9886,N_6491,N_6823);
and U9887 (N_9887,N_6630,N_7391);
nor U9888 (N_9888,N_6001,N_6516);
xnor U9889 (N_9889,N_7337,N_7865);
nor U9890 (N_9890,N_7290,N_7185);
nand U9891 (N_9891,N_6067,N_7972);
nor U9892 (N_9892,N_7034,N_6977);
and U9893 (N_9893,N_6925,N_6534);
and U9894 (N_9894,N_6724,N_6931);
nand U9895 (N_9895,N_7909,N_7014);
or U9896 (N_9896,N_6497,N_7584);
nand U9897 (N_9897,N_7318,N_6417);
nand U9898 (N_9898,N_7174,N_6386);
or U9899 (N_9899,N_6997,N_7166);
or U9900 (N_9900,N_6655,N_6145);
or U9901 (N_9901,N_6502,N_7999);
or U9902 (N_9902,N_6267,N_6930);
and U9903 (N_9903,N_6790,N_7727);
and U9904 (N_9904,N_7985,N_7666);
nor U9905 (N_9905,N_7145,N_6914);
or U9906 (N_9906,N_6943,N_6359);
or U9907 (N_9907,N_7879,N_7402);
nor U9908 (N_9908,N_7171,N_7033);
and U9909 (N_9909,N_7904,N_6601);
or U9910 (N_9910,N_6089,N_6042);
nor U9911 (N_9911,N_7962,N_7100);
nand U9912 (N_9912,N_6606,N_6982);
or U9913 (N_9913,N_7874,N_6995);
and U9914 (N_9914,N_7531,N_7392);
nand U9915 (N_9915,N_7200,N_7396);
nor U9916 (N_9916,N_6636,N_7948);
nand U9917 (N_9917,N_7658,N_7223);
and U9918 (N_9918,N_6325,N_6518);
and U9919 (N_9919,N_7347,N_7057);
or U9920 (N_9920,N_6295,N_7144);
or U9921 (N_9921,N_7300,N_6695);
nand U9922 (N_9922,N_6625,N_7221);
and U9923 (N_9923,N_6221,N_6844);
nand U9924 (N_9924,N_7570,N_7591);
nor U9925 (N_9925,N_6303,N_6763);
nor U9926 (N_9926,N_7365,N_7808);
and U9927 (N_9927,N_6706,N_6788);
nand U9928 (N_9928,N_6812,N_7717);
nor U9929 (N_9929,N_7597,N_7070);
or U9930 (N_9930,N_6560,N_7710);
nand U9931 (N_9931,N_7135,N_6100);
or U9932 (N_9932,N_7099,N_7551);
or U9933 (N_9933,N_7821,N_6355);
nand U9934 (N_9934,N_6970,N_7660);
or U9935 (N_9935,N_6885,N_6562);
and U9936 (N_9936,N_7282,N_6593);
nand U9937 (N_9937,N_6150,N_6609);
and U9938 (N_9938,N_6470,N_7730);
and U9939 (N_9939,N_6422,N_6803);
and U9940 (N_9940,N_6879,N_6116);
nand U9941 (N_9941,N_7752,N_7633);
nor U9942 (N_9942,N_7319,N_7342);
or U9943 (N_9943,N_7927,N_7379);
and U9944 (N_9944,N_6104,N_6517);
nand U9945 (N_9945,N_7339,N_7157);
nand U9946 (N_9946,N_6612,N_7298);
and U9947 (N_9947,N_7139,N_6156);
xor U9948 (N_9948,N_6374,N_7231);
nor U9949 (N_9949,N_7031,N_6523);
or U9950 (N_9950,N_6624,N_7961);
nor U9951 (N_9951,N_6308,N_7404);
nor U9952 (N_9952,N_6865,N_7257);
and U9953 (N_9953,N_7288,N_6492);
and U9954 (N_9954,N_7399,N_6021);
and U9955 (N_9955,N_6119,N_6693);
and U9956 (N_9956,N_6488,N_6636);
nor U9957 (N_9957,N_6984,N_7978);
xor U9958 (N_9958,N_6040,N_7861);
nand U9959 (N_9959,N_7982,N_7104);
nand U9960 (N_9960,N_6322,N_6767);
and U9961 (N_9961,N_6401,N_6784);
and U9962 (N_9962,N_6904,N_6145);
nor U9963 (N_9963,N_7369,N_6152);
nor U9964 (N_9964,N_7197,N_7223);
or U9965 (N_9965,N_6795,N_7229);
nor U9966 (N_9966,N_7444,N_7409);
or U9967 (N_9967,N_6367,N_6940);
nand U9968 (N_9968,N_6708,N_6213);
or U9969 (N_9969,N_6236,N_7461);
or U9970 (N_9970,N_7599,N_6104);
nor U9971 (N_9971,N_6315,N_6620);
xor U9972 (N_9972,N_6029,N_6551);
nor U9973 (N_9973,N_6188,N_6500);
nor U9974 (N_9974,N_7138,N_6415);
and U9975 (N_9975,N_6613,N_7921);
xor U9976 (N_9976,N_7641,N_7710);
and U9977 (N_9977,N_6006,N_7087);
nand U9978 (N_9978,N_6990,N_7654);
nand U9979 (N_9979,N_7399,N_6089);
and U9980 (N_9980,N_6875,N_7398);
nor U9981 (N_9981,N_6154,N_6666);
nor U9982 (N_9982,N_7785,N_7363);
nor U9983 (N_9983,N_7452,N_6951);
or U9984 (N_9984,N_6352,N_6225);
nor U9985 (N_9985,N_7783,N_7108);
or U9986 (N_9986,N_7889,N_7854);
and U9987 (N_9987,N_6514,N_6156);
and U9988 (N_9988,N_6795,N_7203);
or U9989 (N_9989,N_6881,N_6249);
nand U9990 (N_9990,N_7887,N_7496);
and U9991 (N_9991,N_6116,N_7657);
or U9992 (N_9992,N_6783,N_6346);
nor U9993 (N_9993,N_7899,N_7692);
xnor U9994 (N_9994,N_7034,N_7402);
or U9995 (N_9995,N_7372,N_7057);
or U9996 (N_9996,N_7239,N_6073);
nor U9997 (N_9997,N_7571,N_7244);
and U9998 (N_9998,N_6111,N_7781);
nand U9999 (N_9999,N_7468,N_6300);
nand UO_0 (O_0,N_8818,N_9160);
or UO_1 (O_1,N_8346,N_9705);
and UO_2 (O_2,N_8082,N_9475);
nand UO_3 (O_3,N_8380,N_9277);
and UO_4 (O_4,N_8345,N_9389);
xor UO_5 (O_5,N_8111,N_8465);
xor UO_6 (O_6,N_8398,N_9483);
nor UO_7 (O_7,N_9465,N_9262);
nor UO_8 (O_8,N_9456,N_9020);
or UO_9 (O_9,N_8130,N_8533);
nor UO_10 (O_10,N_9949,N_8745);
or UO_11 (O_11,N_9355,N_8020);
nor UO_12 (O_12,N_9528,N_9142);
or UO_13 (O_13,N_8768,N_9971);
nor UO_14 (O_14,N_9058,N_9400);
nand UO_15 (O_15,N_9302,N_8249);
or UO_16 (O_16,N_8305,N_9496);
xor UO_17 (O_17,N_9487,N_9586);
or UO_18 (O_18,N_8207,N_8522);
nand UO_19 (O_19,N_8877,N_9289);
nand UO_20 (O_20,N_9579,N_8413);
nor UO_21 (O_21,N_9741,N_8660);
nor UO_22 (O_22,N_9181,N_8667);
nor UO_23 (O_23,N_8945,N_8620);
nor UO_24 (O_24,N_9447,N_9328);
or UO_25 (O_25,N_9081,N_9342);
nor UO_26 (O_26,N_9788,N_9866);
or UO_27 (O_27,N_8725,N_8496);
nor UO_28 (O_28,N_9336,N_8903);
nand UO_29 (O_29,N_8592,N_9923);
or UO_30 (O_30,N_8555,N_8062);
nor UO_31 (O_31,N_8315,N_9958);
and UO_32 (O_32,N_8896,N_8577);
nor UO_33 (O_33,N_9761,N_8681);
nand UO_34 (O_34,N_8705,N_8858);
or UO_35 (O_35,N_8589,N_8963);
nand UO_36 (O_36,N_8976,N_8230);
nor UO_37 (O_37,N_8418,N_8754);
nand UO_38 (O_38,N_8337,N_8756);
and UO_39 (O_39,N_9733,N_9530);
nor UO_40 (O_40,N_9652,N_9934);
nand UO_41 (O_41,N_9694,N_9632);
nand UO_42 (O_42,N_8158,N_9750);
nand UO_43 (O_43,N_8536,N_8883);
nor UO_44 (O_44,N_8802,N_8987);
or UO_45 (O_45,N_9911,N_9808);
or UO_46 (O_46,N_8609,N_9050);
and UO_47 (O_47,N_8479,N_9504);
or UO_48 (O_48,N_8326,N_8659);
or UO_49 (O_49,N_8443,N_9769);
nor UO_50 (O_50,N_9674,N_8910);
and UO_51 (O_51,N_8543,N_9038);
or UO_52 (O_52,N_8211,N_8750);
or UO_53 (O_53,N_9387,N_8982);
nand UO_54 (O_54,N_9864,N_8591);
nor UO_55 (O_55,N_9977,N_9470);
nand UO_56 (O_56,N_9782,N_8539);
and UO_57 (O_57,N_8478,N_8245);
nand UO_58 (O_58,N_9485,N_9906);
or UO_59 (O_59,N_8823,N_9379);
nand UO_60 (O_60,N_8679,N_9192);
and UO_61 (O_61,N_9905,N_8734);
nor UO_62 (O_62,N_9973,N_9039);
or UO_63 (O_63,N_8237,N_8921);
nand UO_64 (O_64,N_9689,N_8269);
or UO_65 (O_65,N_8138,N_8927);
xor UO_66 (O_66,N_8957,N_9194);
nor UO_67 (O_67,N_9036,N_9871);
and UO_68 (O_68,N_8846,N_9820);
and UO_69 (O_69,N_9435,N_8144);
xnor UO_70 (O_70,N_9129,N_9372);
or UO_71 (O_71,N_9888,N_8018);
or UO_72 (O_72,N_9843,N_9857);
and UO_73 (O_73,N_8170,N_9658);
and UO_74 (O_74,N_8696,N_9356);
nand UO_75 (O_75,N_8387,N_8766);
nor UO_76 (O_76,N_8753,N_9890);
nor UO_77 (O_77,N_9933,N_9224);
and UO_78 (O_78,N_9210,N_9813);
or UO_79 (O_79,N_9320,N_9052);
nand UO_80 (O_80,N_9827,N_9089);
nand UO_81 (O_81,N_9369,N_9719);
nand UO_82 (O_82,N_9563,N_9351);
and UO_83 (O_83,N_8608,N_8419);
nand UO_84 (O_84,N_9133,N_9756);
nand UO_85 (O_85,N_9371,N_8039);
or UO_86 (O_86,N_8073,N_8509);
and UO_87 (O_87,N_8489,N_8476);
nand UO_88 (O_88,N_8325,N_9564);
or UO_89 (O_89,N_9805,N_8310);
and UO_90 (O_90,N_9197,N_9161);
and UO_91 (O_91,N_9230,N_9595);
or UO_92 (O_92,N_8410,N_8395);
nand UO_93 (O_93,N_8266,N_9625);
or UO_94 (O_94,N_8748,N_9540);
or UO_95 (O_95,N_8821,N_8164);
nand UO_96 (O_96,N_8668,N_8236);
nand UO_97 (O_97,N_9109,N_8832);
and UO_98 (O_98,N_8174,N_9294);
nor UO_99 (O_99,N_9554,N_8558);
nand UO_100 (O_100,N_9965,N_9330);
or UO_101 (O_101,N_9641,N_9265);
and UO_102 (O_102,N_9441,N_9019);
nand UO_103 (O_103,N_9031,N_8542);
xnor UO_104 (O_104,N_8778,N_9506);
and UO_105 (O_105,N_8160,N_8633);
nand UO_106 (O_106,N_9755,N_9753);
nor UO_107 (O_107,N_8001,N_8333);
and UO_108 (O_108,N_8240,N_9128);
and UO_109 (O_109,N_9253,N_9437);
nor UO_110 (O_110,N_8518,N_8669);
nand UO_111 (O_111,N_9122,N_9882);
or UO_112 (O_112,N_9489,N_9124);
or UO_113 (O_113,N_9983,N_8698);
or UO_114 (O_114,N_9850,N_8940);
and UO_115 (O_115,N_8666,N_9102);
or UO_116 (O_116,N_8391,N_8183);
and UO_117 (O_117,N_9108,N_8942);
xnor UO_118 (O_118,N_9112,N_8621);
or UO_119 (O_119,N_8168,N_8513);
and UO_120 (O_120,N_9110,N_8864);
and UO_121 (O_121,N_9413,N_8363);
or UO_122 (O_122,N_8360,N_9059);
and UO_123 (O_123,N_9130,N_9821);
and UO_124 (O_124,N_9361,N_9943);
xor UO_125 (O_125,N_8726,N_9633);
nand UO_126 (O_126,N_9023,N_8448);
nor UO_127 (O_127,N_8105,N_9026);
and UO_128 (O_128,N_8457,N_8036);
or UO_129 (O_129,N_9991,N_9681);
nor UO_130 (O_130,N_9243,N_8131);
and UO_131 (O_131,N_9469,N_9683);
or UO_132 (O_132,N_8202,N_9439);
or UO_133 (O_133,N_8133,N_9453);
nor UO_134 (O_134,N_8568,N_8220);
nor UO_135 (O_135,N_8837,N_8193);
nor UO_136 (O_136,N_8757,N_9642);
nor UO_137 (O_137,N_8838,N_8495);
nor UO_138 (O_138,N_9785,N_8070);
xnor UO_139 (O_139,N_8897,N_9378);
nor UO_140 (O_140,N_9323,N_9555);
or UO_141 (O_141,N_8525,N_8546);
nor UO_142 (O_142,N_8534,N_8190);
xor UO_143 (O_143,N_9582,N_8990);
nand UO_144 (O_144,N_8309,N_9069);
nor UO_145 (O_145,N_9819,N_9335);
nand UO_146 (O_146,N_8961,N_8150);
or UO_147 (O_147,N_9987,N_8559);
and UO_148 (O_148,N_8425,N_9478);
or UO_149 (O_149,N_8600,N_8435);
nand UO_150 (O_150,N_8129,N_9845);
and UO_151 (O_151,N_8261,N_8051);
and UO_152 (O_152,N_9182,N_8390);
or UO_153 (O_153,N_9803,N_9634);
or UO_154 (O_154,N_9666,N_9926);
or UO_155 (O_155,N_9889,N_8464);
and UO_156 (O_156,N_8694,N_8707);
nor UO_157 (O_157,N_8894,N_8421);
nor UO_158 (O_158,N_8178,N_9875);
xor UO_159 (O_159,N_8017,N_8729);
or UO_160 (O_160,N_9234,N_8724);
and UO_161 (O_161,N_8132,N_9724);
nor UO_162 (O_162,N_9045,N_8602);
nand UO_163 (O_163,N_9383,N_9732);
or UO_164 (O_164,N_9216,N_8852);
nand UO_165 (O_165,N_8644,N_9776);
nand UO_166 (O_166,N_8804,N_8598);
and UO_167 (O_167,N_9333,N_8710);
and UO_168 (O_168,N_8923,N_9362);
nand UO_169 (O_169,N_9961,N_9405);
nor UO_170 (O_170,N_9282,N_9629);
nand UO_171 (O_171,N_9848,N_9913);
nand UO_172 (O_172,N_8799,N_8011);
nor UO_173 (O_173,N_9638,N_8434);
nor UO_174 (O_174,N_8650,N_9492);
xnor UO_175 (O_175,N_8311,N_9525);
nor UO_176 (O_176,N_8503,N_9448);
or UO_177 (O_177,N_8046,N_8654);
nand UO_178 (O_178,N_8670,N_9749);
and UO_179 (O_179,N_9028,N_9591);
and UO_180 (O_180,N_8831,N_9541);
nand UO_181 (O_181,N_8480,N_9452);
nand UO_182 (O_182,N_8557,N_9752);
nor UO_183 (O_183,N_9644,N_9589);
nand UO_184 (O_184,N_8741,N_8731);
nor UO_185 (O_185,N_8102,N_9440);
nor UO_186 (O_186,N_8252,N_8426);
and UO_187 (O_187,N_8226,N_9273);
nand UO_188 (O_188,N_8357,N_9202);
nand UO_189 (O_189,N_9360,N_9715);
nor UO_190 (O_190,N_8538,N_9975);
nor UO_191 (O_191,N_9556,N_9546);
nor UO_192 (O_192,N_8115,N_9115);
or UO_193 (O_193,N_9252,N_8647);
nor UO_194 (O_194,N_9079,N_9974);
nor UO_195 (O_195,N_8449,N_9096);
or UO_196 (O_196,N_9609,N_8227);
xor UO_197 (O_197,N_8863,N_9712);
nor UO_198 (O_198,N_8442,N_8966);
or UO_199 (O_199,N_9211,N_8549);
or UO_200 (O_200,N_9946,N_9298);
nand UO_201 (O_201,N_8512,N_9764);
nand UO_202 (O_202,N_8468,N_8431);
and UO_203 (O_203,N_8689,N_8121);
or UO_204 (O_204,N_8739,N_8793);
or UO_205 (O_205,N_9463,N_8842);
nand UO_206 (O_206,N_9924,N_9256);
and UO_207 (O_207,N_9099,N_9103);
or UO_208 (O_208,N_8540,N_8165);
nand UO_209 (O_209,N_8658,N_9545);
nor UO_210 (O_210,N_8221,N_8762);
nor UO_211 (O_211,N_8347,N_8569);
or UO_212 (O_212,N_9598,N_8862);
nand UO_213 (O_213,N_9231,N_8428);
or UO_214 (O_214,N_8076,N_9114);
or UO_215 (O_215,N_9444,N_8026);
and UO_216 (O_216,N_9308,N_8447);
nor UO_217 (O_217,N_9090,N_9064);
or UO_218 (O_218,N_9482,N_9012);
nand UO_219 (O_219,N_9673,N_9338);
nor UO_220 (O_220,N_9880,N_8191);
xor UO_221 (O_221,N_9768,N_9140);
nand UO_222 (O_222,N_8673,N_9056);
or UO_223 (O_223,N_8025,N_8408);
nor UO_224 (O_224,N_8566,N_9948);
or UO_225 (O_225,N_8071,N_9604);
nor UO_226 (O_226,N_9316,N_8330);
or UO_227 (O_227,N_8157,N_8021);
nand UO_228 (O_228,N_9071,N_8350);
and UO_229 (O_229,N_8939,N_9490);
or UO_230 (O_230,N_9380,N_8833);
nand UO_231 (O_231,N_8572,N_8937);
nand UO_232 (O_232,N_9818,N_8893);
nor UO_233 (O_233,N_9570,N_9222);
nand UO_234 (O_234,N_8752,N_8914);
nor UO_235 (O_235,N_9789,N_8152);
or UO_236 (O_236,N_8275,N_9030);
or UO_237 (O_237,N_8242,N_9852);
and UO_238 (O_238,N_8367,N_8335);
nand UO_239 (O_239,N_9837,N_8235);
or UO_240 (O_240,N_9590,N_8231);
and UO_241 (O_241,N_8873,N_9895);
nor UO_242 (O_242,N_9804,N_8091);
nor UO_243 (O_243,N_9003,N_8143);
or UO_244 (O_244,N_8219,N_9557);
or UO_245 (O_245,N_8359,N_8550);
nand UO_246 (O_246,N_8086,N_9690);
and UO_247 (O_247,N_9344,N_9876);
nor UO_248 (O_248,N_8742,N_8114);
nand UO_249 (O_249,N_8388,N_8640);
nand UO_250 (O_250,N_9816,N_9858);
and UO_251 (O_251,N_8779,N_9872);
nor UO_252 (O_252,N_9739,N_9601);
or UO_253 (O_253,N_9146,N_8224);
and UO_254 (O_254,N_8173,N_9418);
nand UO_255 (O_255,N_8494,N_9951);
or UO_256 (O_256,N_9425,N_9723);
nor UO_257 (O_257,N_9502,N_8262);
nor UO_258 (O_258,N_9022,N_8188);
and UO_259 (O_259,N_9095,N_8989);
nor UO_260 (O_260,N_8321,N_8653);
or UO_261 (O_261,N_9430,N_8389);
nor UO_262 (O_262,N_9917,N_9364);
nor UO_263 (O_263,N_9429,N_9669);
nor UO_264 (O_264,N_8339,N_9029);
nand UO_265 (O_265,N_9760,N_8198);
and UO_266 (O_266,N_9794,N_9806);
or UO_267 (O_267,N_9565,N_8520);
nand UO_268 (O_268,N_8088,N_8280);
nand UO_269 (O_269,N_8394,N_9147);
nor UO_270 (O_270,N_8067,N_9834);
or UO_271 (O_271,N_8294,N_9537);
and UO_272 (O_272,N_9709,N_8850);
nor UO_273 (O_273,N_9722,N_9959);
nand UO_274 (O_274,N_9054,N_8652);
nor UO_275 (O_275,N_9840,N_8047);
or UO_276 (O_276,N_8445,N_8348);
nor UO_277 (O_277,N_8905,N_8083);
and UO_278 (O_278,N_8195,N_9393);
and UO_279 (O_279,N_8081,N_9600);
or UO_280 (O_280,N_8255,N_8740);
and UO_281 (O_281,N_9618,N_9575);
and UO_282 (O_282,N_8316,N_8570);
nor UO_283 (O_283,N_8161,N_9293);
nor UO_284 (O_284,N_8747,N_9016);
or UO_285 (O_285,N_9771,N_9377);
nor UO_286 (O_286,N_9067,N_9212);
and UO_287 (O_287,N_9568,N_8706);
nor UO_288 (O_288,N_8034,N_8743);
or UO_289 (O_289,N_8580,N_8848);
nor UO_290 (O_290,N_8898,N_9763);
and UO_291 (O_291,N_8415,N_9986);
nor UO_292 (O_292,N_8634,N_9665);
nor UO_293 (O_293,N_9126,N_9375);
and UO_294 (O_294,N_9966,N_9744);
and UO_295 (O_295,N_9676,N_9063);
nor UO_296 (O_296,N_8213,N_8909);
and UO_297 (O_297,N_9479,N_8225);
nor UO_298 (O_298,N_9711,N_8642);
or UO_299 (O_299,N_8092,N_9094);
nand UO_300 (O_300,N_9141,N_8618);
or UO_301 (O_301,N_8931,N_8474);
and UO_302 (O_302,N_9286,N_8407);
or UO_303 (O_303,N_9612,N_8506);
nor UO_304 (O_304,N_8376,N_8057);
and UO_305 (O_305,N_9886,N_8303);
nand UO_306 (O_306,N_8267,N_8635);
nor UO_307 (O_307,N_9969,N_9627);
nor UO_308 (O_308,N_9571,N_8798);
nor UO_309 (O_309,N_9457,N_8947);
nand UO_310 (O_310,N_8044,N_9793);
or UO_311 (O_311,N_9428,N_9299);
and UO_312 (O_312,N_9896,N_9326);
or UO_313 (O_313,N_9386,N_8383);
and UO_314 (O_314,N_8941,N_8682);
and UO_315 (O_315,N_9855,N_8099);
xor UO_316 (O_316,N_9092,N_8451);
nor UO_317 (O_317,N_9559,N_8994);
nor UO_318 (O_318,N_9004,N_9390);
nor UO_319 (O_319,N_8167,N_9508);
nand UO_320 (O_320,N_8192,N_8875);
nand UO_321 (O_321,N_9593,N_8194);
nor UO_322 (O_322,N_9100,N_9839);
and UO_323 (O_323,N_9828,N_8087);
nor UO_324 (O_324,N_9825,N_8065);
xor UO_325 (O_325,N_8432,N_9849);
or UO_326 (O_326,N_8764,N_9713);
nand UO_327 (O_327,N_9513,N_8678);
or UO_328 (O_328,N_9640,N_9920);
or UO_329 (O_329,N_8692,N_8677);
or UO_330 (O_330,N_8003,N_8933);
or UO_331 (O_331,N_8406,N_9259);
and UO_332 (O_332,N_8027,N_8477);
and UO_333 (O_333,N_8127,N_8908);
or UO_334 (O_334,N_8217,N_8876);
nand UO_335 (O_335,N_8530,N_9399);
nor UO_336 (O_336,N_8604,N_9416);
xor UO_337 (O_337,N_8212,N_8153);
and UO_338 (O_338,N_9310,N_9121);
nand UO_339 (O_339,N_9186,N_9879);
nor UO_340 (O_340,N_9795,N_8645);
and UO_341 (O_341,N_9280,N_8996);
nor UO_342 (O_342,N_8384,N_9410);
nand UO_343 (O_343,N_8343,N_9534);
and UO_344 (O_344,N_8505,N_8308);
or UO_345 (O_345,N_8601,N_9939);
and UO_346 (O_346,N_8603,N_9932);
or UO_347 (O_347,N_9955,N_8334);
nor UO_348 (O_348,N_9519,N_8354);
or UO_349 (O_349,N_8735,N_9321);
and UO_350 (O_350,N_8291,N_9835);
or UO_351 (O_351,N_9844,N_8560);
nor UO_352 (O_352,N_8110,N_8323);
or UO_353 (O_353,N_9236,N_8285);
or UO_354 (O_354,N_8488,N_8134);
nor UO_355 (O_355,N_8777,N_9358);
xnor UO_356 (O_356,N_9248,N_9315);
nand UO_357 (O_357,N_8769,N_9171);
and UO_358 (O_358,N_9660,N_9251);
or UO_359 (O_359,N_8938,N_8655);
nor UO_360 (O_360,N_9445,N_8935);
nor UO_361 (O_361,N_8736,N_9717);
nand UO_362 (O_362,N_8300,N_8272);
and UO_363 (O_363,N_9748,N_9376);
nor UO_364 (O_364,N_8920,N_8934);
and UO_365 (O_365,N_8946,N_8282);
or UO_366 (O_366,N_9979,N_8885);
nor UO_367 (O_367,N_9195,N_9495);
or UO_368 (O_368,N_8578,N_8830);
and UO_369 (O_369,N_9581,N_8627);
xnor UO_370 (O_370,N_9451,N_8952);
nor UO_371 (O_371,N_8562,N_8414);
or UO_372 (O_372,N_9152,N_8109);
or UO_373 (O_373,N_8890,N_9972);
or UO_374 (O_374,N_8919,N_8292);
nand UO_375 (O_375,N_9264,N_8907);
or UO_376 (O_376,N_9798,N_8761);
or UO_377 (O_377,N_8843,N_8738);
nand UO_378 (O_378,N_8624,N_9883);
nor UO_379 (O_379,N_8785,N_9068);
xor UO_380 (O_380,N_9529,N_9158);
and UO_381 (O_381,N_8077,N_9918);
nand UO_382 (O_382,N_9784,N_8712);
and UO_383 (O_383,N_8959,N_8547);
nor UO_384 (O_384,N_8500,N_8041);
and UO_385 (O_385,N_8780,N_8732);
nand UO_386 (O_386,N_8386,N_9859);
nor UO_387 (O_387,N_8416,N_9421);
nand UO_388 (O_388,N_8402,N_8064);
nor UO_389 (O_389,N_9851,N_8686);
nor UO_390 (O_390,N_9411,N_9436);
nand UO_391 (O_391,N_8140,N_9057);
and UO_392 (O_392,N_8048,N_8470);
or UO_393 (O_393,N_8800,N_9459);
or UO_394 (O_394,N_9745,N_9619);
nor UO_395 (O_395,N_9536,N_8450);
nor UO_396 (O_396,N_8597,N_9964);
nor UO_397 (O_397,N_8038,N_8299);
nand UO_398 (O_398,N_8979,N_9414);
nand UO_399 (O_399,N_8617,N_9157);
nand UO_400 (O_400,N_9381,N_8648);
or UO_401 (O_401,N_9686,N_8709);
nand UO_402 (O_402,N_9091,N_8853);
or UO_403 (O_403,N_8599,N_9936);
nand UO_404 (O_404,N_9088,N_8312);
nand UO_405 (O_405,N_8684,N_8180);
and UO_406 (O_406,N_8789,N_8290);
and UO_407 (O_407,N_9515,N_8595);
or UO_408 (O_408,N_9558,N_9624);
nor UO_409 (O_409,N_8163,N_9704);
nor UO_410 (O_410,N_8819,N_9037);
and UO_411 (O_411,N_8962,N_8454);
nand UO_412 (O_412,N_9655,N_8607);
nand UO_413 (O_413,N_9462,N_9678);
or UO_414 (O_414,N_8467,N_8004);
and UO_415 (O_415,N_9433,N_8007);
and UO_416 (O_416,N_9007,N_8593);
and UO_417 (O_417,N_9066,N_8590);
nor UO_418 (O_418,N_9040,N_8548);
nand UO_419 (O_419,N_9533,N_9909);
or UO_420 (O_420,N_9842,N_9992);
or UO_421 (O_421,N_8200,N_9269);
nand UO_422 (O_422,N_9201,N_8805);
nand UO_423 (O_423,N_8370,N_9567);
nor UO_424 (O_424,N_9867,N_8459);
nor UO_425 (O_425,N_9209,N_9925);
xor UO_426 (O_426,N_9395,N_9947);
xnor UO_427 (O_427,N_8055,N_9566);
nor UO_428 (O_428,N_8544,N_8301);
nor UO_429 (O_429,N_9297,N_9341);
nor UO_430 (O_430,N_8708,N_9935);
or UO_431 (O_431,N_9576,N_8626);
nand UO_432 (O_432,N_8377,N_9423);
or UO_433 (O_433,N_8135,N_9300);
or UO_434 (O_434,N_8998,N_8169);
and UO_435 (O_435,N_9093,N_8810);
and UO_436 (O_436,N_8795,N_8032);
nand UO_437 (O_437,N_9311,N_8835);
or UO_438 (O_438,N_8462,N_9814);
or UO_439 (O_439,N_8529,N_8953);
and UO_440 (O_440,N_8553,N_8949);
nor UO_441 (O_441,N_9370,N_8880);
nor UO_442 (O_442,N_8146,N_8671);
or UO_443 (O_443,N_8098,N_9759);
nand UO_444 (O_444,N_9501,N_9334);
or UO_445 (O_445,N_9175,N_9863);
or UO_446 (O_446,N_8571,N_8579);
and UO_447 (O_447,N_9797,N_8822);
xnor UO_448 (O_448,N_8074,N_9065);
and UO_449 (O_449,N_8867,N_9027);
and UO_450 (O_450,N_9073,N_9783);
nand UO_451 (O_451,N_8713,N_8286);
nor UO_452 (O_452,N_9017,N_9762);
nand UO_453 (O_453,N_9561,N_8006);
xnor UO_454 (O_454,N_9854,N_9348);
nand UO_455 (O_455,N_9167,N_9084);
nor UO_456 (O_456,N_8205,N_9226);
nand UO_457 (O_457,N_8924,N_8078);
and UO_458 (O_458,N_9144,N_8373);
nand UO_459 (O_459,N_9894,N_8482);
xnor UO_460 (O_460,N_9322,N_8068);
or UO_461 (O_461,N_9295,N_8155);
or UO_462 (O_462,N_8737,N_9291);
xor UO_463 (O_463,N_8702,N_9464);
nor UO_464 (O_464,N_8765,N_8711);
nor UO_465 (O_465,N_8986,N_9846);
nor UO_466 (O_466,N_9930,N_8181);
and UO_467 (O_467,N_8199,N_9373);
or UO_468 (O_468,N_9608,N_8094);
nand UO_469 (O_469,N_9931,N_9915);
nand UO_470 (O_470,N_8786,N_8050);
nor UO_471 (O_471,N_9870,N_9468);
and UO_472 (O_472,N_9869,N_8166);
nor UO_473 (O_473,N_9626,N_9309);
nand UO_474 (O_474,N_9679,N_8186);
nor UO_475 (O_475,N_9174,N_9118);
xnor UO_476 (O_476,N_8759,N_8781);
nor UO_477 (O_477,N_9580,N_8069);
nor UO_478 (O_478,N_8177,N_8632);
and UO_479 (O_479,N_8646,N_9006);
and UO_480 (O_480,N_9013,N_8535);
nor UO_481 (O_481,N_9646,N_9662);
or UO_482 (O_482,N_8507,N_8287);
and UO_483 (O_483,N_9402,N_8049);
nand UO_484 (O_484,N_9136,N_8719);
or UO_485 (O_485,N_9266,N_8714);
nor UO_486 (O_486,N_9401,N_9535);
nor UO_487 (O_487,N_8095,N_8906);
and UO_488 (O_488,N_8901,N_8733);
or UO_489 (O_489,N_8234,N_9471);
and UO_490 (O_490,N_8374,N_9737);
or UO_491 (O_491,N_8452,N_8817);
and UO_492 (O_492,N_9774,N_9912);
and UO_493 (O_493,N_9659,N_9521);
and UO_494 (O_494,N_9817,N_9275);
nor UO_495 (O_495,N_9018,N_9420);
nor UO_496 (O_496,N_8685,N_8120);
nand UO_497 (O_497,N_9283,N_9611);
nor UO_498 (O_498,N_9780,N_8970);
nor UO_499 (O_499,N_9021,N_8293);
and UO_500 (O_500,N_8090,N_8208);
nand UO_501 (O_501,N_9367,N_9494);
or UO_502 (O_502,N_9176,N_8501);
and UO_503 (O_503,N_9204,N_9578);
or UO_504 (O_504,N_8239,N_8879);
or UO_505 (O_505,N_9696,N_9384);
nor UO_506 (O_506,N_8277,N_8318);
or UO_507 (O_507,N_8241,N_8375);
nand UO_508 (O_508,N_8322,N_9688);
nor UO_509 (O_509,N_9922,N_9740);
or UO_510 (O_510,N_9183,N_9168);
nand UO_511 (O_511,N_8888,N_8815);
and UO_512 (O_512,N_9885,N_8441);
or UO_513 (O_513,N_8185,N_8420);
xor UO_514 (O_514,N_9901,N_9417);
nor UO_515 (O_515,N_9319,N_9198);
or UO_516 (O_516,N_9055,N_8466);
nand UO_517 (O_517,N_8461,N_9648);
nor UO_518 (O_518,N_9412,N_8932);
and UO_519 (O_519,N_9105,N_9488);
nand UO_520 (O_520,N_8586,N_9670);
nand UO_521 (O_521,N_9682,N_8106);
xor UO_522 (O_522,N_9592,N_9047);
and UO_523 (O_523,N_9207,N_8128);
or UO_524 (O_524,N_8997,N_8774);
and UO_525 (O_525,N_9191,N_9661);
nor UO_526 (O_526,N_8913,N_9352);
and UO_527 (O_527,N_9729,N_8954);
or UO_528 (O_528,N_9596,N_9874);
and UO_529 (O_529,N_8834,N_9200);
nand UO_530 (O_530,N_9597,N_9177);
nand UO_531 (O_531,N_9639,N_9442);
and UO_532 (O_532,N_9993,N_8688);
or UO_533 (O_533,N_8508,N_8216);
nand UO_534 (O_534,N_9426,N_8403);
or UO_535 (O_535,N_9725,N_9937);
or UO_536 (O_536,N_9053,N_8251);
nand UO_537 (O_537,N_8061,N_8612);
or UO_538 (O_538,N_9622,N_9786);
nand UO_539 (O_539,N_8904,N_8126);
nand UO_540 (O_540,N_8002,N_9125);
and UO_541 (O_541,N_8749,N_9304);
nand UO_542 (O_542,N_8382,N_8223);
nor UO_543 (O_543,N_9553,N_8453);
nor UO_544 (O_544,N_8537,N_8141);
xor UO_545 (O_545,N_8854,N_8840);
and UO_546 (O_546,N_9654,N_9233);
and UO_547 (O_547,N_9138,N_8751);
and UO_548 (O_548,N_9276,N_9657);
xor UO_549 (O_549,N_9061,N_8891);
or UO_550 (O_550,N_8259,N_9347);
and UO_551 (O_551,N_9139,N_9610);
nand UO_552 (O_552,N_8616,N_8978);
or UO_553 (O_553,N_8511,N_9847);
and UO_554 (O_554,N_8154,N_9498);
nor UO_555 (O_555,N_8699,N_8024);
nand UO_556 (O_556,N_8409,N_9223);
and UO_557 (O_557,N_9279,N_8871);
nor UO_558 (O_558,N_9271,N_9602);
and UO_559 (O_559,N_8317,N_9268);
nor UO_560 (O_560,N_8722,N_8575);
nand UO_561 (O_561,N_8967,N_9623);
nor UO_562 (O_562,N_9518,N_8147);
and UO_563 (O_563,N_8490,N_9143);
nor UO_564 (O_564,N_8826,N_8258);
nor UO_565 (O_565,N_9241,N_8148);
nand UO_566 (O_566,N_9727,N_9077);
nor UO_567 (O_567,N_9317,N_9217);
or UO_568 (O_568,N_9551,N_8964);
nand UO_569 (O_569,N_9583,N_9403);
or UO_570 (O_570,N_8497,N_8755);
nor UO_571 (O_571,N_9716,N_9116);
nand UO_572 (O_572,N_8304,N_8320);
and UO_573 (O_573,N_8005,N_9225);
nand UO_574 (O_574,N_8984,N_8878);
nor UO_575 (O_575,N_9836,N_9916);
and UO_576 (O_576,N_9550,N_9187);
nor UO_577 (O_577,N_9111,N_8456);
nand UO_578 (O_578,N_9954,N_8332);
and UO_579 (O_579,N_8839,N_8502);
nand UO_580 (O_580,N_9284,N_9621);
nor UO_581 (O_581,N_9516,N_8329);
nand UO_582 (O_582,N_9929,N_8771);
nand UO_583 (O_583,N_9824,N_9278);
or UO_584 (O_584,N_9573,N_9190);
and UO_585 (O_585,N_8022,N_9305);
nand UO_586 (O_586,N_8246,N_9878);
nand UO_587 (O_587,N_9726,N_8159);
or UO_588 (O_588,N_8981,N_9945);
nand UO_589 (O_589,N_9742,N_9684);
or UO_590 (O_590,N_8510,N_8444);
or UO_591 (O_591,N_8423,N_9856);
or UO_592 (O_592,N_8053,N_9512);
nor UO_593 (O_593,N_8123,N_8072);
and UO_594 (O_594,N_8031,N_9497);
and UO_595 (O_595,N_9014,N_8565);
and UO_596 (O_596,N_9941,N_9349);
nor UO_597 (O_597,N_8524,N_9398);
nor UO_598 (O_598,N_8895,N_8149);
nand UO_599 (O_599,N_9617,N_8767);
or UO_600 (O_600,N_8983,N_9692);
or UO_601 (O_601,N_9461,N_9354);
nand UO_602 (O_602,N_9270,N_8233);
xor UO_603 (O_603,N_8899,N_8142);
nand UO_604 (O_604,N_9049,N_9766);
nor UO_605 (O_605,N_9353,N_9877);
and UO_606 (O_606,N_9424,N_8016);
nand UO_607 (O_607,N_9048,N_9543);
or UO_608 (O_608,N_8691,N_8772);
or UO_609 (O_609,N_8232,N_9238);
nor UO_610 (O_610,N_8056,N_8860);
nand UO_611 (O_611,N_8728,N_8980);
nand UO_612 (O_612,N_8112,N_8253);
or UO_613 (O_613,N_9833,N_9113);
or UO_614 (O_614,N_8531,N_8656);
or UO_615 (O_615,N_8486,N_9892);
and UO_616 (O_616,N_9454,N_9968);
nand UO_617 (O_617,N_8201,N_9123);
nor UO_618 (O_618,N_9656,N_8008);
or UO_619 (O_619,N_8836,N_8175);
nor UO_620 (O_620,N_8930,N_9770);
nor UO_621 (O_621,N_8430,N_9032);
nor UO_622 (O_622,N_9903,N_9887);
and UO_623 (O_623,N_8107,N_9514);
nor UO_624 (O_624,N_8613,N_9976);
nor UO_625 (O_625,N_8331,N_9346);
nand UO_626 (O_626,N_8912,N_8328);
or UO_627 (O_627,N_9407,N_9097);
and UO_628 (O_628,N_8274,N_9313);
nor UO_629 (O_629,N_9082,N_8587);
nand UO_630 (O_630,N_8381,N_8424);
nand UO_631 (O_631,N_8366,N_8855);
and UO_632 (O_632,N_9891,N_9431);
nor UO_633 (O_633,N_9357,N_8715);
nand UO_634 (O_634,N_9672,N_8701);
and UO_635 (O_635,N_8922,N_8137);
nand UO_636 (O_636,N_9005,N_8372);
and UO_637 (O_637,N_8639,N_9163);
nor UO_638 (O_638,N_8972,N_9898);
nand UO_639 (O_639,N_8554,N_8187);
nor UO_640 (O_640,N_8630,N_9509);
and UO_641 (O_641,N_9967,N_9206);
xnor UO_642 (O_642,N_9606,N_8911);
and UO_643 (O_643,N_8475,N_8349);
nand UO_644 (O_644,N_9254,N_9910);
and UO_645 (O_645,N_9826,N_8787);
or UO_646 (O_646,N_9107,N_8458);
nor UO_647 (O_647,N_8481,N_9329);
nand UO_648 (O_648,N_9180,N_8276);
nand UO_649 (O_649,N_8956,N_8327);
nand UO_650 (O_650,N_8614,N_8256);
and UO_651 (O_651,N_9997,N_9466);
nand UO_652 (O_652,N_8023,N_9153);
xor UO_653 (O_653,N_9427,N_8929);
and UO_654 (O_654,N_9812,N_9246);
nand UO_655 (O_655,N_9643,N_8218);
and UO_656 (O_656,N_9574,N_8806);
nor UO_657 (O_657,N_9708,N_8857);
nor UO_658 (O_658,N_8623,N_9701);
and UO_659 (O_659,N_8561,N_9149);
nor UO_660 (O_660,N_8556,N_9337);
or UO_661 (O_661,N_9605,N_9340);
or UO_662 (O_662,N_9218,N_8564);
or UO_663 (O_663,N_8532,N_9213);
and UO_664 (O_664,N_9823,N_9060);
or UO_665 (O_665,N_8052,N_9758);
or UO_666 (O_666,N_9893,N_9781);
and UO_667 (O_667,N_8491,N_9815);
and UO_668 (O_668,N_9510,N_9307);
nor UO_669 (O_669,N_9865,N_8013);
nor UO_670 (O_670,N_9170,N_9476);
nor UO_671 (O_671,N_8030,N_8975);
and UO_672 (O_672,N_9594,N_9331);
and UO_673 (O_673,N_8324,N_8108);
nand UO_674 (O_674,N_8399,N_8369);
and UO_675 (O_675,N_8605,N_9517);
nand UO_676 (O_676,N_8664,N_8296);
nand UO_677 (O_677,N_8125,N_9085);
nor UO_678 (O_678,N_8816,N_8847);
nand UO_679 (O_679,N_9693,N_8584);
nand UO_680 (O_680,N_8117,N_8746);
nor UO_681 (O_681,N_8361,N_9985);
nand UO_682 (O_682,N_9809,N_9743);
nand UO_683 (O_683,N_8116,N_8718);
or UO_684 (O_684,N_9062,N_8631);
or UO_685 (O_685,N_9647,N_8210);
nand UO_686 (O_686,N_8948,N_8716);
and UO_687 (O_687,N_8872,N_9086);
nand UO_688 (O_688,N_8063,N_8951);
nand UO_689 (O_689,N_8636,N_9636);
and UO_690 (O_690,N_8827,N_9185);
nand UO_691 (O_691,N_8401,N_9382);
and UO_692 (O_692,N_8196,N_9703);
nor UO_693 (O_693,N_8790,N_8662);
and UO_694 (O_694,N_9950,N_8281);
nand UO_695 (O_695,N_9388,N_8574);
nand UO_696 (O_696,N_9188,N_9051);
xor UO_697 (O_697,N_8596,N_8965);
or UO_698 (O_698,N_8969,N_8791);
nand UO_699 (O_699,N_8824,N_9009);
xor UO_700 (O_700,N_9631,N_9714);
and UO_701 (O_701,N_9015,N_9687);
nand UO_702 (O_702,N_9523,N_9205);
nand UO_703 (O_703,N_8519,N_8615);
nor UO_704 (O_704,N_8045,N_8663);
and UO_705 (O_705,N_8336,N_9500);
or UO_706 (O_706,N_8368,N_9404);
and UO_707 (O_707,N_8995,N_9730);
and UO_708 (O_708,N_9982,N_9547);
nor UO_709 (O_709,N_9560,N_8378);
nand UO_710 (O_710,N_8955,N_8118);
or UO_711 (O_711,N_8573,N_8881);
and UO_712 (O_712,N_8870,N_9884);
nand UO_713 (O_713,N_8674,N_9860);
nor UO_714 (O_714,N_9902,N_9080);
nand UO_715 (O_715,N_9978,N_8676);
or UO_716 (O_716,N_9778,N_8439);
and UO_717 (O_717,N_9532,N_8567);
nor UO_718 (O_718,N_9312,N_8625);
nand UO_719 (O_719,N_9645,N_9990);
nand UO_720 (O_720,N_8926,N_9024);
or UO_721 (O_721,N_8637,N_9368);
nor UO_722 (O_722,N_9184,N_9196);
and UO_723 (O_723,N_8991,N_8340);
or UO_724 (O_724,N_9728,N_8364);
nor UO_725 (O_725,N_8882,N_8176);
nor UO_726 (O_726,N_9862,N_8298);
nand UO_727 (O_727,N_9635,N_9075);
nand UO_728 (O_728,N_9419,N_9735);
nor UO_729 (O_729,N_9791,N_8429);
or UO_730 (O_730,N_9810,N_9984);
nor UO_731 (O_731,N_9172,N_8865);
nand UO_732 (O_732,N_8284,N_8427);
and UO_733 (O_733,N_9258,N_9989);
nor UO_734 (O_734,N_9438,N_9134);
nor UO_735 (O_735,N_9106,N_9861);
nor UO_736 (O_736,N_9098,N_9000);
and UO_737 (O_737,N_8440,N_9630);
and UO_738 (O_738,N_8472,N_8244);
or UO_739 (O_739,N_8104,N_9165);
nor UO_740 (O_740,N_8629,N_8365);
xnor UO_741 (O_741,N_9043,N_9232);
nand UO_742 (O_742,N_9359,N_9928);
or UO_743 (O_743,N_8889,N_9394);
nand UO_744 (O_744,N_9117,N_9306);
nor UO_745 (O_745,N_9332,N_9408);
and UO_746 (O_746,N_9562,N_9460);
or UO_747 (O_747,N_8974,N_8887);
nand UO_748 (O_748,N_9288,N_8861);
nor UO_749 (O_749,N_9166,N_9841);
xor UO_750 (O_750,N_8059,N_9548);
nor UO_751 (O_751,N_8992,N_8319);
nand UO_752 (O_752,N_8066,N_8783);
xnor UO_753 (O_753,N_8973,N_8845);
or UO_754 (O_754,N_8516,N_8782);
xnor UO_755 (O_755,N_8156,N_9374);
nor UO_756 (O_756,N_8675,N_9220);
or UO_757 (O_757,N_9314,N_8396);
and UO_758 (O_758,N_8700,N_8796);
nand UO_759 (O_759,N_9025,N_8139);
or UO_760 (O_760,N_9801,N_9422);
and UO_761 (O_761,N_9988,N_9397);
or UO_762 (O_762,N_8900,N_9396);
nor UO_763 (O_763,N_9777,N_8079);
or UO_764 (O_764,N_8145,N_9343);
and UO_765 (O_765,N_9614,N_9503);
and UO_766 (O_766,N_8471,N_8371);
nand UO_767 (O_767,N_9587,N_9083);
nor UO_768 (O_768,N_8527,N_8763);
or UO_769 (O_769,N_8643,N_9480);
nand UO_770 (O_770,N_8197,N_8928);
or UO_771 (O_771,N_9938,N_8215);
or UO_772 (O_772,N_8801,N_9281);
or UO_773 (O_773,N_9520,N_8042);
nand UO_774 (O_774,N_8985,N_9486);
nand UO_775 (O_775,N_9907,N_9588);
nand UO_776 (O_776,N_9391,N_9119);
or UO_777 (O_777,N_9491,N_9035);
or UO_778 (O_778,N_9544,N_9292);
or UO_779 (O_779,N_9507,N_9900);
and UO_780 (O_780,N_8943,N_9267);
or UO_781 (O_781,N_8925,N_9980);
xnor UO_782 (O_782,N_9542,N_8775);
or UO_783 (O_783,N_9620,N_8999);
nand UO_784 (O_784,N_9104,N_9325);
or UO_785 (O_785,N_8264,N_9285);
and UO_786 (O_786,N_8084,N_8776);
or UO_787 (O_787,N_8868,N_9159);
nand UO_788 (O_788,N_8085,N_9237);
or UO_789 (O_789,N_9940,N_9274);
and UO_790 (O_790,N_8551,N_8270);
and UO_791 (O_791,N_8803,N_8342);
and UO_792 (O_792,N_8588,N_9150);
nand UO_793 (O_793,N_8352,N_9953);
nand UO_794 (O_794,N_8526,N_9677);
or UO_795 (O_795,N_8455,N_9339);
nand UO_796 (O_796,N_9219,N_8971);
nand UO_797 (O_797,N_9493,N_8545);
or UO_798 (O_798,N_8214,N_8385);
nand UO_799 (O_799,N_8690,N_8060);
nor UO_800 (O_800,N_9511,N_9087);
nand UO_801 (O_801,N_8841,N_8638);
nand UO_802 (O_802,N_8271,N_9245);
nand UO_803 (O_803,N_8436,N_9944);
nand UO_804 (O_804,N_9260,N_9552);
nor UO_805 (O_805,N_9822,N_9538);
nand UO_806 (O_806,N_8353,N_9415);
nor UO_807 (O_807,N_9526,N_9765);
nor UO_808 (O_808,N_9956,N_8268);
or UO_809 (O_809,N_8859,N_9718);
xor UO_810 (O_810,N_8019,N_9699);
or UO_811 (O_811,N_8243,N_8437);
and UO_812 (O_812,N_9577,N_9615);
nand UO_813 (O_813,N_8314,N_9076);
or UO_814 (O_814,N_8723,N_9042);
nand UO_815 (O_815,N_8828,N_8619);
nand UO_816 (O_816,N_8122,N_9010);
or UO_817 (O_817,N_9914,N_9838);
and UO_818 (O_818,N_9613,N_8438);
or UO_819 (O_819,N_8493,N_9754);
nand UO_820 (O_820,N_8103,N_9214);
xor UO_821 (O_821,N_8392,N_9473);
or UO_822 (O_822,N_8809,N_9215);
or UO_823 (O_823,N_9261,N_9199);
and UO_824 (O_824,N_8514,N_8043);
xor UO_825 (O_825,N_9458,N_9668);
or UO_826 (O_826,N_9481,N_9156);
and UO_827 (O_827,N_9173,N_8037);
and UO_828 (O_828,N_9522,N_9899);
or UO_829 (O_829,N_9779,N_9881);
nand UO_830 (O_830,N_8936,N_8651);
or UO_831 (O_831,N_9365,N_9235);
nor UO_832 (O_832,N_8379,N_9350);
or UO_833 (O_833,N_9527,N_9832);
and UO_834 (O_834,N_9539,N_8917);
and UO_835 (O_835,N_9145,N_8582);
nand UO_836 (O_836,N_9996,N_9710);
or UO_837 (O_837,N_9449,N_9963);
and UO_838 (O_838,N_8968,N_9101);
nor UO_839 (O_839,N_8892,N_8351);
nand UO_840 (O_840,N_8162,N_8015);
and UO_841 (O_841,N_8794,N_8697);
nand UO_842 (O_842,N_8417,N_8228);
or UO_843 (O_843,N_9164,N_9443);
or UO_844 (O_844,N_8844,N_8628);
or UO_845 (O_845,N_9607,N_8096);
nand UO_846 (O_846,N_9041,N_8788);
nand UO_847 (O_847,N_9366,N_8029);
and UO_848 (O_848,N_9650,N_8874);
and UO_849 (O_849,N_9155,N_8950);
and UO_850 (O_850,N_9675,N_9720);
nand UO_851 (O_851,N_9628,N_9734);
nor UO_852 (O_852,N_9995,N_8279);
or UO_853 (O_853,N_8209,N_8773);
and UO_854 (O_854,N_8356,N_8054);
or UO_855 (O_855,N_8720,N_8622);
and UO_856 (O_856,N_9074,N_8829);
or UO_857 (O_857,N_8641,N_8182);
or UO_858 (O_858,N_9203,N_9301);
or UO_859 (O_859,N_8229,N_8820);
and UO_860 (O_860,N_8814,N_9455);
nand UO_861 (O_861,N_9775,N_8918);
or UO_862 (O_862,N_8058,N_9653);
nand UO_863 (O_863,N_9078,N_9178);
and UO_864 (O_864,N_9998,N_9505);
or UO_865 (O_865,N_8254,N_8649);
nor UO_866 (O_866,N_9731,N_8035);
and UO_867 (O_867,N_8792,N_8869);
nand UO_868 (O_868,N_9477,N_9363);
nor UO_869 (O_869,N_9667,N_9952);
or UO_870 (O_870,N_9773,N_8247);
or UO_871 (O_871,N_9873,N_9685);
or UO_872 (O_872,N_8594,N_9290);
nand UO_873 (O_873,N_8851,N_8813);
or UO_874 (O_874,N_9970,N_9303);
or UO_875 (O_875,N_8610,N_9957);
or UO_876 (O_876,N_9651,N_9649);
nor UO_877 (O_877,N_9240,N_8528);
and UO_878 (O_878,N_9796,N_8101);
and UO_879 (O_879,N_8521,N_8797);
and UO_880 (O_880,N_9962,N_9746);
and UO_881 (O_881,N_8278,N_9008);
and UO_882 (O_882,N_8289,N_8344);
nand UO_883 (O_883,N_8412,N_9868);
nor UO_884 (O_884,N_9691,N_8886);
or UO_885 (O_885,N_9327,N_8206);
or UO_886 (O_886,N_9603,N_8393);
nand UO_887 (O_887,N_8238,N_8184);
or UO_888 (O_888,N_9738,N_8358);
and UO_889 (O_889,N_8487,N_8288);
and UO_890 (O_890,N_9385,N_8687);
nor UO_891 (O_891,N_8263,N_8657);
or UO_892 (O_892,N_8080,N_9227);
or UO_893 (O_893,N_9193,N_8257);
nor UO_894 (O_894,N_9757,N_8703);
xnor UO_895 (O_895,N_8404,N_8313);
and UO_896 (O_896,N_9830,N_8469);
or UO_897 (O_897,N_8446,N_9070);
nand UO_898 (O_898,N_8405,N_9239);
nor UO_899 (O_899,N_8136,N_9772);
or UO_900 (O_900,N_9671,N_9921);
nor UO_901 (O_901,N_9698,N_9702);
or UO_902 (O_902,N_8811,N_9033);
or UO_903 (O_903,N_9853,N_9697);
nand UO_904 (O_904,N_8204,N_9569);
nand UO_905 (O_905,N_8012,N_9706);
and UO_906 (O_906,N_9229,N_9831);
nand UO_907 (O_907,N_9120,N_8849);
nand UO_908 (O_908,N_9484,N_9467);
nand UO_909 (O_909,N_9999,N_8172);
and UO_910 (O_910,N_8902,N_8856);
and UO_911 (O_911,N_9919,N_8760);
and UO_912 (O_912,N_8014,N_9531);
or UO_913 (O_913,N_9044,N_8283);
or UO_914 (O_914,N_9751,N_9392);
or UO_915 (O_915,N_9432,N_9811);
nor UO_916 (O_916,N_8484,N_9942);
and UO_917 (O_917,N_9695,N_9799);
nor UO_918 (O_918,N_9127,N_8541);
or UO_919 (O_919,N_8680,N_9549);
nor UO_920 (O_920,N_8113,N_8362);
nand UO_921 (O_921,N_9829,N_9994);
nand UO_922 (O_922,N_8093,N_8988);
nor UO_923 (O_923,N_8784,N_9499);
or UO_924 (O_924,N_9221,N_9927);
nor UO_925 (O_925,N_9800,N_8203);
nand UO_926 (O_926,N_9707,N_9787);
and UO_927 (O_927,N_8581,N_8583);
or UO_928 (O_928,N_8222,N_9981);
xnor UO_929 (O_929,N_9616,N_8661);
or UO_930 (O_930,N_9584,N_8273);
and UO_931 (O_931,N_9446,N_8151);
nor UO_932 (O_932,N_9721,N_9897);
or UO_933 (O_933,N_8397,N_9137);
and UO_934 (O_934,N_8179,N_8515);
or UO_935 (O_935,N_9700,N_9034);
nor UO_936 (O_936,N_8189,N_8265);
nor UO_937 (O_937,N_8463,N_8807);
nor UO_938 (O_938,N_9002,N_8916);
and UO_939 (O_939,N_8606,N_9472);
and UO_940 (O_940,N_9572,N_9450);
and UO_941 (O_941,N_8552,N_8944);
or UO_942 (O_942,N_8758,N_8585);
nand UO_943 (O_943,N_8433,N_9148);
and UO_944 (O_944,N_9747,N_9263);
or UO_945 (O_945,N_8422,N_8411);
or UO_946 (O_946,N_9585,N_8884);
or UO_947 (O_947,N_8295,N_8563);
nand UO_948 (O_948,N_8040,N_9680);
or UO_949 (O_949,N_9228,N_9736);
or UO_950 (O_950,N_8730,N_8693);
nor UO_951 (O_951,N_8000,N_9663);
and UO_952 (O_952,N_8473,N_8075);
nor UO_953 (O_953,N_8958,N_8993);
and UO_954 (O_954,N_9179,N_9247);
nor UO_955 (O_955,N_8825,N_9296);
xnor UO_956 (O_956,N_9072,N_9904);
nand UO_957 (O_957,N_9908,N_8499);
nor UO_958 (O_958,N_8866,N_8808);
nand UO_959 (O_959,N_8704,N_8483);
and UO_960 (O_960,N_9250,N_8770);
and UO_961 (O_961,N_8683,N_9189);
and UO_962 (O_962,N_9287,N_8302);
and UO_963 (O_963,N_8744,N_8977);
nand UO_964 (O_964,N_9162,N_9242);
and UO_965 (O_965,N_8400,N_9208);
and UO_966 (O_966,N_9154,N_8338);
or UO_967 (O_967,N_9767,N_8960);
nand UO_968 (O_968,N_8727,N_8665);
nand UO_969 (O_969,N_8033,N_9409);
nand UO_970 (O_970,N_8717,N_8248);
nor UO_971 (O_971,N_9318,N_8672);
or UO_972 (O_972,N_9792,N_8119);
nand UO_973 (O_973,N_8721,N_8171);
nor UO_974 (O_974,N_8097,N_8307);
nor UO_975 (O_975,N_8250,N_8460);
and UO_976 (O_976,N_9406,N_8355);
and UO_977 (O_977,N_8260,N_9249);
nor UO_978 (O_978,N_8297,N_8498);
or UO_979 (O_979,N_8010,N_8504);
and UO_980 (O_980,N_9011,N_8485);
or UO_981 (O_981,N_9257,N_9960);
and UO_982 (O_982,N_8089,N_8523);
and UO_983 (O_983,N_9807,N_8100);
or UO_984 (O_984,N_9046,N_9169);
nor UO_985 (O_985,N_9131,N_8124);
nand UO_986 (O_986,N_9001,N_9244);
or UO_987 (O_987,N_8576,N_8009);
and UO_988 (O_988,N_9664,N_9132);
or UO_989 (O_989,N_9255,N_9434);
nor UO_990 (O_990,N_9599,N_8695);
and UO_991 (O_991,N_8915,N_9474);
nand UO_992 (O_992,N_8812,N_8306);
xnor UO_993 (O_993,N_9524,N_9272);
nor UO_994 (O_994,N_9135,N_8492);
nand UO_995 (O_995,N_9637,N_9802);
or UO_996 (O_996,N_9151,N_8341);
nor UO_997 (O_997,N_9790,N_8517);
or UO_998 (O_998,N_9324,N_8611);
nand UO_999 (O_999,N_9345,N_8028);
or UO_1000 (O_1000,N_8572,N_9335);
and UO_1001 (O_1001,N_8907,N_8364);
or UO_1002 (O_1002,N_8169,N_8020);
nor UO_1003 (O_1003,N_9516,N_8539);
nand UO_1004 (O_1004,N_8816,N_9532);
and UO_1005 (O_1005,N_8826,N_8479);
nor UO_1006 (O_1006,N_8786,N_9346);
or UO_1007 (O_1007,N_9182,N_9427);
xnor UO_1008 (O_1008,N_9515,N_9531);
nand UO_1009 (O_1009,N_8878,N_9788);
or UO_1010 (O_1010,N_9698,N_8428);
nand UO_1011 (O_1011,N_9615,N_9673);
nand UO_1012 (O_1012,N_8501,N_8086);
nor UO_1013 (O_1013,N_9583,N_9675);
nand UO_1014 (O_1014,N_8472,N_9549);
and UO_1015 (O_1015,N_8459,N_9292);
nor UO_1016 (O_1016,N_8876,N_9799);
nand UO_1017 (O_1017,N_9112,N_9401);
and UO_1018 (O_1018,N_9034,N_8799);
and UO_1019 (O_1019,N_9779,N_9410);
nand UO_1020 (O_1020,N_9629,N_8040);
nand UO_1021 (O_1021,N_9817,N_8912);
or UO_1022 (O_1022,N_8165,N_9859);
and UO_1023 (O_1023,N_8723,N_8705);
nor UO_1024 (O_1024,N_9706,N_9635);
nor UO_1025 (O_1025,N_8167,N_9348);
or UO_1026 (O_1026,N_9373,N_8097);
and UO_1027 (O_1027,N_8411,N_9391);
nor UO_1028 (O_1028,N_8300,N_9029);
nand UO_1029 (O_1029,N_9822,N_9743);
nand UO_1030 (O_1030,N_9957,N_8121);
nor UO_1031 (O_1031,N_8708,N_8187);
xnor UO_1032 (O_1032,N_9335,N_8729);
nand UO_1033 (O_1033,N_8971,N_8382);
and UO_1034 (O_1034,N_8857,N_8221);
or UO_1035 (O_1035,N_9432,N_8072);
and UO_1036 (O_1036,N_9001,N_8155);
nand UO_1037 (O_1037,N_9519,N_8611);
xor UO_1038 (O_1038,N_9459,N_9849);
nor UO_1039 (O_1039,N_8401,N_8941);
and UO_1040 (O_1040,N_9039,N_8663);
and UO_1041 (O_1041,N_9433,N_9974);
nand UO_1042 (O_1042,N_9332,N_8958);
or UO_1043 (O_1043,N_8640,N_8863);
nor UO_1044 (O_1044,N_8688,N_9454);
or UO_1045 (O_1045,N_9868,N_9054);
nor UO_1046 (O_1046,N_8058,N_9246);
and UO_1047 (O_1047,N_9056,N_8800);
nand UO_1048 (O_1048,N_9676,N_8236);
and UO_1049 (O_1049,N_8724,N_8856);
nor UO_1050 (O_1050,N_9615,N_8353);
or UO_1051 (O_1051,N_8446,N_9652);
nor UO_1052 (O_1052,N_9971,N_8812);
nand UO_1053 (O_1053,N_9204,N_9902);
nand UO_1054 (O_1054,N_9278,N_9933);
or UO_1055 (O_1055,N_8285,N_9647);
nand UO_1056 (O_1056,N_9922,N_9115);
or UO_1057 (O_1057,N_9505,N_8885);
nand UO_1058 (O_1058,N_8212,N_8465);
nor UO_1059 (O_1059,N_9613,N_9190);
and UO_1060 (O_1060,N_9867,N_8296);
or UO_1061 (O_1061,N_9998,N_8602);
or UO_1062 (O_1062,N_9051,N_8704);
nor UO_1063 (O_1063,N_9072,N_8254);
and UO_1064 (O_1064,N_9031,N_8617);
nand UO_1065 (O_1065,N_8574,N_8399);
nor UO_1066 (O_1066,N_8794,N_8566);
nand UO_1067 (O_1067,N_9758,N_8215);
or UO_1068 (O_1068,N_9704,N_9714);
or UO_1069 (O_1069,N_9266,N_8493);
and UO_1070 (O_1070,N_9333,N_9147);
or UO_1071 (O_1071,N_8125,N_9963);
and UO_1072 (O_1072,N_9717,N_8057);
nand UO_1073 (O_1073,N_9110,N_9822);
and UO_1074 (O_1074,N_8730,N_9488);
or UO_1075 (O_1075,N_8360,N_9865);
and UO_1076 (O_1076,N_9872,N_8230);
nand UO_1077 (O_1077,N_9923,N_9939);
and UO_1078 (O_1078,N_9410,N_9862);
or UO_1079 (O_1079,N_9366,N_9744);
or UO_1080 (O_1080,N_8219,N_8186);
nor UO_1081 (O_1081,N_9368,N_9521);
or UO_1082 (O_1082,N_8373,N_9777);
and UO_1083 (O_1083,N_9019,N_8400);
nand UO_1084 (O_1084,N_9101,N_8259);
and UO_1085 (O_1085,N_9737,N_9466);
nor UO_1086 (O_1086,N_8095,N_9105);
or UO_1087 (O_1087,N_9663,N_8774);
nand UO_1088 (O_1088,N_9938,N_9200);
or UO_1089 (O_1089,N_9366,N_8821);
or UO_1090 (O_1090,N_8857,N_8763);
xor UO_1091 (O_1091,N_9759,N_8424);
nor UO_1092 (O_1092,N_8777,N_9108);
nor UO_1093 (O_1093,N_8047,N_9396);
nor UO_1094 (O_1094,N_8642,N_8345);
xor UO_1095 (O_1095,N_9985,N_9960);
nand UO_1096 (O_1096,N_9788,N_8649);
nor UO_1097 (O_1097,N_8558,N_8348);
nor UO_1098 (O_1098,N_9107,N_9794);
nor UO_1099 (O_1099,N_9556,N_9903);
or UO_1100 (O_1100,N_9991,N_8440);
or UO_1101 (O_1101,N_8282,N_9247);
and UO_1102 (O_1102,N_9722,N_9121);
nor UO_1103 (O_1103,N_8601,N_8560);
nor UO_1104 (O_1104,N_8116,N_8300);
nand UO_1105 (O_1105,N_9359,N_9800);
or UO_1106 (O_1106,N_9490,N_8925);
nor UO_1107 (O_1107,N_9093,N_9424);
nand UO_1108 (O_1108,N_9361,N_8757);
nor UO_1109 (O_1109,N_9324,N_9746);
nor UO_1110 (O_1110,N_8126,N_9251);
nand UO_1111 (O_1111,N_9468,N_8852);
and UO_1112 (O_1112,N_9007,N_8947);
or UO_1113 (O_1113,N_9103,N_9421);
nor UO_1114 (O_1114,N_8173,N_9496);
and UO_1115 (O_1115,N_9953,N_9647);
nand UO_1116 (O_1116,N_9496,N_8733);
and UO_1117 (O_1117,N_8740,N_8378);
and UO_1118 (O_1118,N_9220,N_8277);
nand UO_1119 (O_1119,N_8608,N_8860);
or UO_1120 (O_1120,N_9477,N_8404);
or UO_1121 (O_1121,N_9375,N_9361);
nor UO_1122 (O_1122,N_8023,N_9466);
and UO_1123 (O_1123,N_9713,N_9754);
xnor UO_1124 (O_1124,N_9741,N_9651);
nand UO_1125 (O_1125,N_9564,N_9234);
nand UO_1126 (O_1126,N_8771,N_8809);
nand UO_1127 (O_1127,N_8778,N_8025);
nor UO_1128 (O_1128,N_8256,N_9125);
and UO_1129 (O_1129,N_8414,N_9936);
nor UO_1130 (O_1130,N_9674,N_8752);
and UO_1131 (O_1131,N_9658,N_9108);
or UO_1132 (O_1132,N_8559,N_8084);
or UO_1133 (O_1133,N_9829,N_9035);
or UO_1134 (O_1134,N_8470,N_8801);
or UO_1135 (O_1135,N_8180,N_8230);
xor UO_1136 (O_1136,N_8954,N_9690);
nor UO_1137 (O_1137,N_9390,N_9526);
nand UO_1138 (O_1138,N_8015,N_9444);
nor UO_1139 (O_1139,N_8316,N_8449);
or UO_1140 (O_1140,N_8357,N_8367);
or UO_1141 (O_1141,N_8489,N_9610);
or UO_1142 (O_1142,N_8377,N_8870);
or UO_1143 (O_1143,N_8575,N_8598);
nor UO_1144 (O_1144,N_9776,N_8109);
nand UO_1145 (O_1145,N_9828,N_9180);
xnor UO_1146 (O_1146,N_9365,N_8146);
xor UO_1147 (O_1147,N_9514,N_8954);
nor UO_1148 (O_1148,N_8577,N_9452);
nand UO_1149 (O_1149,N_9053,N_8068);
and UO_1150 (O_1150,N_9203,N_9938);
and UO_1151 (O_1151,N_9080,N_8687);
or UO_1152 (O_1152,N_9267,N_9385);
and UO_1153 (O_1153,N_8427,N_9763);
or UO_1154 (O_1154,N_9901,N_9701);
and UO_1155 (O_1155,N_9824,N_9439);
nor UO_1156 (O_1156,N_9236,N_9081);
nor UO_1157 (O_1157,N_9385,N_9963);
or UO_1158 (O_1158,N_9699,N_8431);
nand UO_1159 (O_1159,N_9942,N_8750);
or UO_1160 (O_1160,N_8577,N_9703);
nand UO_1161 (O_1161,N_9528,N_8941);
and UO_1162 (O_1162,N_8732,N_9280);
xnor UO_1163 (O_1163,N_8013,N_8622);
nor UO_1164 (O_1164,N_9094,N_8202);
nand UO_1165 (O_1165,N_9531,N_9975);
and UO_1166 (O_1166,N_9346,N_8713);
nand UO_1167 (O_1167,N_8354,N_8630);
and UO_1168 (O_1168,N_9331,N_8704);
or UO_1169 (O_1169,N_8730,N_9375);
and UO_1170 (O_1170,N_9598,N_8633);
or UO_1171 (O_1171,N_9534,N_8166);
nand UO_1172 (O_1172,N_9352,N_8967);
or UO_1173 (O_1173,N_8342,N_9510);
nand UO_1174 (O_1174,N_9996,N_9778);
nor UO_1175 (O_1175,N_8815,N_8316);
or UO_1176 (O_1176,N_9351,N_9245);
nand UO_1177 (O_1177,N_9837,N_8491);
nor UO_1178 (O_1178,N_8367,N_8959);
or UO_1179 (O_1179,N_8296,N_9869);
or UO_1180 (O_1180,N_9911,N_8681);
nand UO_1181 (O_1181,N_8655,N_8654);
nor UO_1182 (O_1182,N_9777,N_9472);
nand UO_1183 (O_1183,N_8545,N_9988);
nor UO_1184 (O_1184,N_8432,N_9156);
and UO_1185 (O_1185,N_8090,N_9291);
nand UO_1186 (O_1186,N_8347,N_9896);
or UO_1187 (O_1187,N_8601,N_8628);
nand UO_1188 (O_1188,N_9170,N_8334);
or UO_1189 (O_1189,N_9636,N_8019);
nand UO_1190 (O_1190,N_9939,N_9602);
and UO_1191 (O_1191,N_8160,N_9624);
nand UO_1192 (O_1192,N_9654,N_9412);
nand UO_1193 (O_1193,N_9591,N_8509);
nand UO_1194 (O_1194,N_9820,N_9130);
and UO_1195 (O_1195,N_8272,N_8454);
nor UO_1196 (O_1196,N_8521,N_8146);
nand UO_1197 (O_1197,N_9476,N_8398);
nand UO_1198 (O_1198,N_8979,N_9705);
or UO_1199 (O_1199,N_8432,N_8089);
nand UO_1200 (O_1200,N_8514,N_8438);
nor UO_1201 (O_1201,N_8465,N_8291);
nand UO_1202 (O_1202,N_9302,N_8703);
and UO_1203 (O_1203,N_9638,N_8662);
nor UO_1204 (O_1204,N_8636,N_9854);
nor UO_1205 (O_1205,N_8456,N_9995);
or UO_1206 (O_1206,N_8025,N_9634);
nand UO_1207 (O_1207,N_8215,N_9017);
nand UO_1208 (O_1208,N_8044,N_9475);
and UO_1209 (O_1209,N_8308,N_9184);
and UO_1210 (O_1210,N_9179,N_9100);
nor UO_1211 (O_1211,N_9161,N_9929);
and UO_1212 (O_1212,N_9154,N_8752);
or UO_1213 (O_1213,N_8757,N_8622);
nor UO_1214 (O_1214,N_9269,N_9758);
or UO_1215 (O_1215,N_8589,N_8468);
nand UO_1216 (O_1216,N_9063,N_9037);
and UO_1217 (O_1217,N_9961,N_8338);
xor UO_1218 (O_1218,N_8092,N_9034);
or UO_1219 (O_1219,N_9148,N_8534);
and UO_1220 (O_1220,N_8608,N_9654);
nand UO_1221 (O_1221,N_9030,N_9701);
nand UO_1222 (O_1222,N_8761,N_8518);
or UO_1223 (O_1223,N_8281,N_8782);
nor UO_1224 (O_1224,N_9622,N_9248);
or UO_1225 (O_1225,N_9198,N_9065);
and UO_1226 (O_1226,N_9878,N_8439);
or UO_1227 (O_1227,N_8276,N_9674);
nand UO_1228 (O_1228,N_8470,N_8089);
nand UO_1229 (O_1229,N_9226,N_8480);
and UO_1230 (O_1230,N_9203,N_9899);
and UO_1231 (O_1231,N_9892,N_8834);
nand UO_1232 (O_1232,N_9281,N_8456);
and UO_1233 (O_1233,N_9232,N_8662);
or UO_1234 (O_1234,N_8447,N_8934);
or UO_1235 (O_1235,N_8189,N_9035);
nor UO_1236 (O_1236,N_8841,N_9397);
nor UO_1237 (O_1237,N_9277,N_9038);
nand UO_1238 (O_1238,N_8686,N_9982);
nand UO_1239 (O_1239,N_9099,N_8585);
nand UO_1240 (O_1240,N_8104,N_8669);
and UO_1241 (O_1241,N_8356,N_8651);
and UO_1242 (O_1242,N_9607,N_9742);
and UO_1243 (O_1243,N_8591,N_8394);
and UO_1244 (O_1244,N_8867,N_9568);
or UO_1245 (O_1245,N_8207,N_8099);
and UO_1246 (O_1246,N_9432,N_9516);
or UO_1247 (O_1247,N_8450,N_8903);
xor UO_1248 (O_1248,N_9577,N_9402);
nor UO_1249 (O_1249,N_8496,N_9979);
nand UO_1250 (O_1250,N_9558,N_9245);
nor UO_1251 (O_1251,N_8960,N_9880);
nor UO_1252 (O_1252,N_8187,N_8189);
nor UO_1253 (O_1253,N_9895,N_8380);
nand UO_1254 (O_1254,N_9710,N_9569);
and UO_1255 (O_1255,N_8643,N_9171);
and UO_1256 (O_1256,N_8682,N_8201);
and UO_1257 (O_1257,N_8621,N_8804);
or UO_1258 (O_1258,N_8139,N_9343);
nor UO_1259 (O_1259,N_8006,N_8517);
nor UO_1260 (O_1260,N_8148,N_8356);
nand UO_1261 (O_1261,N_8675,N_8323);
and UO_1262 (O_1262,N_9577,N_8460);
nor UO_1263 (O_1263,N_8789,N_9964);
nor UO_1264 (O_1264,N_9635,N_8619);
and UO_1265 (O_1265,N_8228,N_8203);
nor UO_1266 (O_1266,N_9941,N_8165);
and UO_1267 (O_1267,N_8947,N_9232);
nor UO_1268 (O_1268,N_9039,N_8602);
and UO_1269 (O_1269,N_9886,N_8123);
and UO_1270 (O_1270,N_9849,N_9632);
and UO_1271 (O_1271,N_8260,N_8571);
or UO_1272 (O_1272,N_9683,N_8121);
or UO_1273 (O_1273,N_9469,N_8530);
nand UO_1274 (O_1274,N_8380,N_9142);
and UO_1275 (O_1275,N_8738,N_8017);
and UO_1276 (O_1276,N_9567,N_9985);
or UO_1277 (O_1277,N_9443,N_9125);
nand UO_1278 (O_1278,N_8177,N_9499);
and UO_1279 (O_1279,N_8468,N_8987);
and UO_1280 (O_1280,N_8813,N_9543);
or UO_1281 (O_1281,N_8410,N_8924);
nand UO_1282 (O_1282,N_9011,N_8403);
or UO_1283 (O_1283,N_8444,N_9822);
or UO_1284 (O_1284,N_9647,N_9883);
nor UO_1285 (O_1285,N_9983,N_8083);
xnor UO_1286 (O_1286,N_8849,N_8949);
and UO_1287 (O_1287,N_8586,N_8122);
nand UO_1288 (O_1288,N_8355,N_9066);
nand UO_1289 (O_1289,N_8619,N_9146);
or UO_1290 (O_1290,N_9775,N_8532);
or UO_1291 (O_1291,N_9669,N_8420);
nor UO_1292 (O_1292,N_9720,N_8762);
nand UO_1293 (O_1293,N_9872,N_8572);
nor UO_1294 (O_1294,N_8114,N_9354);
nor UO_1295 (O_1295,N_8528,N_8444);
nand UO_1296 (O_1296,N_9533,N_9745);
or UO_1297 (O_1297,N_8296,N_9532);
or UO_1298 (O_1298,N_9362,N_9178);
nor UO_1299 (O_1299,N_9209,N_8629);
and UO_1300 (O_1300,N_9495,N_9728);
nand UO_1301 (O_1301,N_8232,N_8376);
nor UO_1302 (O_1302,N_8811,N_8948);
and UO_1303 (O_1303,N_9432,N_8883);
or UO_1304 (O_1304,N_8518,N_8474);
and UO_1305 (O_1305,N_9521,N_9059);
or UO_1306 (O_1306,N_8419,N_8369);
nor UO_1307 (O_1307,N_9495,N_8294);
nor UO_1308 (O_1308,N_9911,N_8179);
and UO_1309 (O_1309,N_9955,N_9867);
or UO_1310 (O_1310,N_8892,N_8416);
nor UO_1311 (O_1311,N_8034,N_8144);
or UO_1312 (O_1312,N_8780,N_8989);
and UO_1313 (O_1313,N_8898,N_9659);
or UO_1314 (O_1314,N_8746,N_9432);
and UO_1315 (O_1315,N_8873,N_8680);
nor UO_1316 (O_1316,N_8108,N_9725);
nor UO_1317 (O_1317,N_9230,N_8527);
or UO_1318 (O_1318,N_9405,N_8315);
nor UO_1319 (O_1319,N_9302,N_8954);
or UO_1320 (O_1320,N_9844,N_9444);
nand UO_1321 (O_1321,N_8769,N_9440);
and UO_1322 (O_1322,N_9233,N_8597);
or UO_1323 (O_1323,N_8601,N_9636);
or UO_1324 (O_1324,N_8536,N_8442);
and UO_1325 (O_1325,N_8589,N_9483);
nor UO_1326 (O_1326,N_8138,N_8513);
xnor UO_1327 (O_1327,N_8089,N_9227);
nor UO_1328 (O_1328,N_8594,N_9429);
or UO_1329 (O_1329,N_9160,N_8521);
or UO_1330 (O_1330,N_9226,N_9142);
and UO_1331 (O_1331,N_8272,N_8589);
nor UO_1332 (O_1332,N_9129,N_8263);
nor UO_1333 (O_1333,N_8766,N_8648);
and UO_1334 (O_1334,N_9798,N_9207);
nor UO_1335 (O_1335,N_8090,N_8910);
nand UO_1336 (O_1336,N_9542,N_8644);
nand UO_1337 (O_1337,N_9031,N_9848);
nor UO_1338 (O_1338,N_9333,N_9279);
nor UO_1339 (O_1339,N_8693,N_9446);
xor UO_1340 (O_1340,N_8815,N_9868);
and UO_1341 (O_1341,N_9895,N_9032);
nand UO_1342 (O_1342,N_8939,N_9369);
or UO_1343 (O_1343,N_9659,N_9635);
and UO_1344 (O_1344,N_9596,N_8808);
or UO_1345 (O_1345,N_9832,N_8025);
or UO_1346 (O_1346,N_9809,N_9988);
nand UO_1347 (O_1347,N_8495,N_9181);
nand UO_1348 (O_1348,N_8477,N_8110);
nand UO_1349 (O_1349,N_9407,N_8418);
nand UO_1350 (O_1350,N_8029,N_8456);
xor UO_1351 (O_1351,N_9928,N_9730);
nor UO_1352 (O_1352,N_9569,N_9507);
nor UO_1353 (O_1353,N_9214,N_8076);
or UO_1354 (O_1354,N_9956,N_9753);
nor UO_1355 (O_1355,N_8987,N_8496);
nand UO_1356 (O_1356,N_8112,N_9008);
or UO_1357 (O_1357,N_9172,N_8807);
nor UO_1358 (O_1358,N_8612,N_8701);
and UO_1359 (O_1359,N_8448,N_9045);
and UO_1360 (O_1360,N_9185,N_9162);
and UO_1361 (O_1361,N_8345,N_9319);
nand UO_1362 (O_1362,N_9639,N_8428);
nand UO_1363 (O_1363,N_8239,N_8515);
nor UO_1364 (O_1364,N_9246,N_9218);
nand UO_1365 (O_1365,N_8875,N_9825);
and UO_1366 (O_1366,N_9213,N_9130);
nand UO_1367 (O_1367,N_8674,N_8139);
nand UO_1368 (O_1368,N_9287,N_9555);
nor UO_1369 (O_1369,N_9572,N_8739);
and UO_1370 (O_1370,N_8281,N_9261);
nand UO_1371 (O_1371,N_9542,N_9533);
and UO_1372 (O_1372,N_8953,N_8249);
nand UO_1373 (O_1373,N_9951,N_9947);
or UO_1374 (O_1374,N_8138,N_8652);
and UO_1375 (O_1375,N_9876,N_8268);
or UO_1376 (O_1376,N_8805,N_9596);
nor UO_1377 (O_1377,N_9836,N_9823);
nand UO_1378 (O_1378,N_8911,N_9213);
nor UO_1379 (O_1379,N_9577,N_9926);
and UO_1380 (O_1380,N_8595,N_9623);
nor UO_1381 (O_1381,N_8657,N_8108);
nor UO_1382 (O_1382,N_9934,N_9292);
nor UO_1383 (O_1383,N_9678,N_8495);
or UO_1384 (O_1384,N_9195,N_9202);
or UO_1385 (O_1385,N_8933,N_8214);
nand UO_1386 (O_1386,N_8834,N_8068);
xor UO_1387 (O_1387,N_9483,N_9445);
or UO_1388 (O_1388,N_9309,N_8691);
and UO_1389 (O_1389,N_8574,N_9968);
nand UO_1390 (O_1390,N_9884,N_8807);
or UO_1391 (O_1391,N_9109,N_8427);
and UO_1392 (O_1392,N_9295,N_8654);
and UO_1393 (O_1393,N_8611,N_8706);
xor UO_1394 (O_1394,N_9594,N_8906);
nor UO_1395 (O_1395,N_9944,N_8285);
or UO_1396 (O_1396,N_8656,N_8459);
nand UO_1397 (O_1397,N_9218,N_9939);
and UO_1398 (O_1398,N_9281,N_8448);
and UO_1399 (O_1399,N_9664,N_8841);
or UO_1400 (O_1400,N_8953,N_8891);
nor UO_1401 (O_1401,N_9971,N_9110);
or UO_1402 (O_1402,N_9075,N_9418);
and UO_1403 (O_1403,N_8740,N_9466);
nand UO_1404 (O_1404,N_8726,N_8472);
or UO_1405 (O_1405,N_9252,N_8745);
and UO_1406 (O_1406,N_8349,N_8479);
nor UO_1407 (O_1407,N_9935,N_9120);
nor UO_1408 (O_1408,N_8641,N_9149);
or UO_1409 (O_1409,N_9998,N_8370);
and UO_1410 (O_1410,N_8649,N_8632);
or UO_1411 (O_1411,N_8121,N_8438);
nor UO_1412 (O_1412,N_9708,N_9518);
nor UO_1413 (O_1413,N_9490,N_9566);
nor UO_1414 (O_1414,N_9112,N_9389);
nor UO_1415 (O_1415,N_8203,N_9525);
or UO_1416 (O_1416,N_8504,N_8013);
and UO_1417 (O_1417,N_9355,N_9576);
nor UO_1418 (O_1418,N_9928,N_8975);
and UO_1419 (O_1419,N_8829,N_8367);
or UO_1420 (O_1420,N_9195,N_8854);
and UO_1421 (O_1421,N_9860,N_8467);
and UO_1422 (O_1422,N_8126,N_8794);
nand UO_1423 (O_1423,N_9240,N_8096);
or UO_1424 (O_1424,N_9404,N_9377);
or UO_1425 (O_1425,N_9246,N_9684);
or UO_1426 (O_1426,N_9816,N_9885);
nand UO_1427 (O_1427,N_9176,N_8826);
or UO_1428 (O_1428,N_8645,N_8982);
nand UO_1429 (O_1429,N_9430,N_8448);
nand UO_1430 (O_1430,N_8096,N_8441);
and UO_1431 (O_1431,N_8243,N_9003);
nor UO_1432 (O_1432,N_8807,N_9732);
nor UO_1433 (O_1433,N_9429,N_9582);
nor UO_1434 (O_1434,N_8749,N_8810);
nand UO_1435 (O_1435,N_9295,N_8614);
nand UO_1436 (O_1436,N_9797,N_8128);
or UO_1437 (O_1437,N_8430,N_9812);
nor UO_1438 (O_1438,N_8207,N_9542);
or UO_1439 (O_1439,N_9487,N_9420);
nor UO_1440 (O_1440,N_8811,N_9618);
nand UO_1441 (O_1441,N_8416,N_8321);
and UO_1442 (O_1442,N_9376,N_9545);
or UO_1443 (O_1443,N_8852,N_8882);
or UO_1444 (O_1444,N_8708,N_8595);
nand UO_1445 (O_1445,N_9927,N_8406);
nand UO_1446 (O_1446,N_8898,N_9756);
and UO_1447 (O_1447,N_8786,N_8416);
and UO_1448 (O_1448,N_8119,N_9203);
and UO_1449 (O_1449,N_8027,N_8128);
nand UO_1450 (O_1450,N_9600,N_8850);
nor UO_1451 (O_1451,N_9966,N_8762);
nor UO_1452 (O_1452,N_8206,N_8055);
xor UO_1453 (O_1453,N_8173,N_9779);
nand UO_1454 (O_1454,N_8876,N_9578);
or UO_1455 (O_1455,N_8942,N_8966);
and UO_1456 (O_1456,N_9720,N_9230);
and UO_1457 (O_1457,N_8255,N_9934);
and UO_1458 (O_1458,N_9653,N_8577);
nand UO_1459 (O_1459,N_9773,N_8668);
nand UO_1460 (O_1460,N_9632,N_9616);
nand UO_1461 (O_1461,N_9202,N_8419);
and UO_1462 (O_1462,N_9670,N_8916);
nand UO_1463 (O_1463,N_9320,N_8769);
and UO_1464 (O_1464,N_8513,N_8780);
or UO_1465 (O_1465,N_8053,N_8416);
nand UO_1466 (O_1466,N_9734,N_9008);
and UO_1467 (O_1467,N_9149,N_8361);
or UO_1468 (O_1468,N_9566,N_8191);
and UO_1469 (O_1469,N_9652,N_9516);
and UO_1470 (O_1470,N_9839,N_8598);
and UO_1471 (O_1471,N_8202,N_9773);
nor UO_1472 (O_1472,N_8260,N_9979);
or UO_1473 (O_1473,N_8550,N_9058);
nand UO_1474 (O_1474,N_8978,N_8737);
and UO_1475 (O_1475,N_9079,N_8967);
or UO_1476 (O_1476,N_8756,N_9884);
nor UO_1477 (O_1477,N_9353,N_9082);
nand UO_1478 (O_1478,N_8165,N_9297);
and UO_1479 (O_1479,N_9538,N_8502);
and UO_1480 (O_1480,N_9627,N_9863);
nand UO_1481 (O_1481,N_9049,N_9324);
nor UO_1482 (O_1482,N_8906,N_9105);
or UO_1483 (O_1483,N_9111,N_9420);
or UO_1484 (O_1484,N_8519,N_9938);
nor UO_1485 (O_1485,N_9035,N_9259);
or UO_1486 (O_1486,N_9674,N_8698);
or UO_1487 (O_1487,N_9670,N_8748);
nor UO_1488 (O_1488,N_9272,N_9301);
nand UO_1489 (O_1489,N_9930,N_9213);
and UO_1490 (O_1490,N_8655,N_8062);
nor UO_1491 (O_1491,N_9114,N_8095);
or UO_1492 (O_1492,N_9128,N_9258);
nor UO_1493 (O_1493,N_9939,N_8492);
nand UO_1494 (O_1494,N_8935,N_9245);
nand UO_1495 (O_1495,N_8954,N_8348);
and UO_1496 (O_1496,N_9136,N_8199);
nor UO_1497 (O_1497,N_9308,N_8830);
nand UO_1498 (O_1498,N_9974,N_9216);
nor UO_1499 (O_1499,N_9956,N_8995);
endmodule