module basic_3000_30000_3500_30_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_794,In_638);
or U1 (N_1,In_1640,In_1290);
nor U2 (N_2,In_975,In_2404);
or U3 (N_3,In_1865,In_579);
or U4 (N_4,In_1429,In_2470);
nand U5 (N_5,In_2097,In_2661);
nor U6 (N_6,In_2045,In_2444);
or U7 (N_7,In_1957,In_1079);
xor U8 (N_8,In_1104,In_611);
or U9 (N_9,In_362,In_1676);
nor U10 (N_10,In_1075,In_1762);
nand U11 (N_11,In_880,In_1219);
xor U12 (N_12,In_2071,In_542);
nand U13 (N_13,In_2802,In_1503);
nand U14 (N_14,In_1664,In_5);
and U15 (N_15,In_1673,In_2084);
nand U16 (N_16,In_2903,In_2359);
and U17 (N_17,In_81,In_262);
or U18 (N_18,In_712,In_2032);
and U19 (N_19,In_2707,In_2273);
xor U20 (N_20,In_1462,In_408);
nand U21 (N_21,In_657,In_1354);
or U22 (N_22,In_1502,In_2892);
xor U23 (N_23,In_2431,In_1214);
and U24 (N_24,In_2539,In_387);
or U25 (N_25,In_1090,In_833);
or U26 (N_26,In_2252,In_1115);
nand U27 (N_27,In_1006,In_233);
nor U28 (N_28,In_1187,In_2468);
xor U29 (N_29,In_799,In_1776);
and U30 (N_30,In_2569,In_1301);
nand U31 (N_31,In_2805,In_516);
xnor U32 (N_32,In_868,In_2472);
or U33 (N_33,In_2495,In_163);
nand U34 (N_34,In_140,In_1695);
and U35 (N_35,In_1207,In_1518);
nor U36 (N_36,In_1517,In_1400);
nor U37 (N_37,In_1575,In_2837);
xor U38 (N_38,In_2755,In_1094);
nor U39 (N_39,In_416,In_2374);
nand U40 (N_40,In_876,In_1661);
nand U41 (N_41,In_1372,In_1936);
and U42 (N_42,In_1925,In_505);
xnor U43 (N_43,In_1060,In_40);
or U44 (N_44,In_1362,In_2192);
xnor U45 (N_45,In_2363,In_1922);
nand U46 (N_46,In_2435,In_1168);
xnor U47 (N_47,In_2749,In_1701);
xnor U48 (N_48,In_1789,In_2390);
or U49 (N_49,In_2686,In_1844);
or U50 (N_50,In_513,In_2684);
and U51 (N_51,In_575,In_822);
nand U52 (N_52,In_2937,In_1063);
xor U53 (N_53,In_2635,In_2051);
nand U54 (N_54,In_1396,In_2382);
nor U55 (N_55,In_2112,In_1847);
nor U56 (N_56,In_1178,In_2486);
xnor U57 (N_57,In_115,In_1623);
xor U58 (N_58,In_308,In_874);
or U59 (N_59,In_1221,In_1620);
xnor U60 (N_60,In_2588,In_652);
nand U61 (N_61,In_1458,In_1333);
or U62 (N_62,In_1113,In_1938);
or U63 (N_63,In_2777,In_1583);
xor U64 (N_64,In_2441,In_2584);
and U65 (N_65,In_2070,In_73);
and U66 (N_66,In_1249,In_654);
xnor U67 (N_67,In_2741,In_711);
or U68 (N_68,In_690,In_2080);
nand U69 (N_69,In_390,In_1770);
nor U70 (N_70,In_2909,In_2411);
or U71 (N_71,In_31,In_1618);
xor U72 (N_72,In_1379,In_627);
xor U73 (N_73,In_924,In_576);
nand U74 (N_74,In_2625,In_174);
nor U75 (N_75,In_2939,In_2908);
nand U76 (N_76,In_77,In_2832);
nor U77 (N_77,In_97,In_2973);
and U78 (N_78,In_46,In_2406);
nand U79 (N_79,In_2245,In_148);
nand U80 (N_80,In_2813,In_34);
and U81 (N_81,In_1752,In_866);
and U82 (N_82,In_374,In_15);
or U83 (N_83,In_20,In_852);
xor U84 (N_84,In_2963,In_38);
nand U85 (N_85,In_412,In_2602);
xor U86 (N_86,In_2727,In_1794);
or U87 (N_87,In_2942,In_2887);
xor U88 (N_88,In_1526,In_1826);
nor U89 (N_89,In_62,In_592);
nand U90 (N_90,In_443,In_996);
xnor U91 (N_91,In_2189,In_1255);
and U92 (N_92,In_1270,In_2241);
nor U93 (N_93,In_1982,In_184);
nor U94 (N_94,In_1602,In_2293);
nand U95 (N_95,In_1629,In_2559);
xor U96 (N_96,In_2193,In_561);
or U97 (N_97,In_2361,In_171);
and U98 (N_98,In_29,In_1325);
nor U99 (N_99,In_104,In_2166);
xor U100 (N_100,In_94,In_2428);
and U101 (N_101,In_206,In_748);
or U102 (N_102,In_2692,In_353);
and U103 (N_103,In_1148,In_1487);
xor U104 (N_104,In_2422,In_51);
and U105 (N_105,In_2175,In_1814);
xor U106 (N_106,In_2966,In_2483);
or U107 (N_107,In_1857,In_2348);
nor U108 (N_108,In_284,In_970);
or U109 (N_109,In_2880,In_753);
xnor U110 (N_110,In_187,In_277);
or U111 (N_111,In_615,In_2249);
nand U112 (N_112,In_2121,In_767);
or U113 (N_113,In_2247,In_2573);
nor U114 (N_114,In_2415,In_2377);
and U115 (N_115,In_1264,In_1283);
nor U116 (N_116,In_774,In_2122);
xor U117 (N_117,In_1638,In_333);
or U118 (N_118,In_2144,In_1659);
xor U119 (N_119,In_380,In_2794);
xor U120 (N_120,In_1973,In_2442);
nor U121 (N_121,In_1646,In_203);
nor U122 (N_122,In_1692,In_1342);
xnor U123 (N_123,In_1564,In_2772);
or U124 (N_124,In_1535,In_901);
or U125 (N_125,In_2980,In_85);
xnor U126 (N_126,In_817,In_1945);
and U127 (N_127,In_1078,In_2745);
or U128 (N_128,In_1439,In_2268);
nand U129 (N_129,In_1477,In_398);
xnor U130 (N_130,In_2465,In_1765);
and U131 (N_131,In_2593,In_1709);
nor U132 (N_132,In_2231,In_2388);
or U133 (N_133,In_2952,In_1771);
xor U134 (N_134,In_1978,In_1025);
and U135 (N_135,In_677,In_662);
nor U136 (N_136,In_1469,In_628);
nor U137 (N_137,In_1190,In_323);
xor U138 (N_138,In_1642,In_481);
and U139 (N_139,In_1251,In_1086);
nor U140 (N_140,In_2039,In_2488);
or U141 (N_141,In_776,In_1277);
or U142 (N_142,In_2111,In_2067);
nor U143 (N_143,In_1314,In_125);
xor U144 (N_144,In_182,In_1530);
nand U145 (N_145,In_824,In_2726);
and U146 (N_146,In_2683,In_2585);
xor U147 (N_147,In_1010,In_1934);
nor U148 (N_148,In_1316,In_2910);
xor U149 (N_149,In_2804,In_2793);
nor U150 (N_150,In_80,In_137);
nor U151 (N_151,In_1622,In_2645);
or U152 (N_152,In_2133,In_2524);
nor U153 (N_153,In_1533,In_446);
nor U154 (N_154,In_2792,In_1445);
and U155 (N_155,In_2314,In_605);
and U156 (N_156,In_1838,In_2556);
and U157 (N_157,In_1900,In_1624);
or U158 (N_158,In_631,In_340);
or U159 (N_159,In_888,In_2616);
or U160 (N_160,In_704,In_2222);
and U161 (N_161,In_733,In_2362);
nand U162 (N_162,In_166,In_1778);
xnor U163 (N_163,In_514,In_781);
or U164 (N_164,In_1785,In_1202);
nand U165 (N_165,In_2353,In_2852);
nand U166 (N_166,In_702,In_836);
or U167 (N_167,In_2103,In_2279);
or U168 (N_168,In_2370,In_1805);
nor U169 (N_169,In_70,In_1364);
nand U170 (N_170,In_264,In_1741);
xor U171 (N_171,In_1143,In_1757);
and U172 (N_172,In_986,In_1134);
and U173 (N_173,In_1605,In_2970);
nor U174 (N_174,In_2449,In_1706);
xnor U175 (N_175,In_293,In_2494);
and U176 (N_176,In_1554,In_509);
or U177 (N_177,In_1157,In_2376);
or U178 (N_178,In_2038,In_512);
xnor U179 (N_179,In_687,In_21);
nand U180 (N_180,In_1939,In_1877);
xor U181 (N_181,In_1881,In_665);
xor U182 (N_182,In_908,In_1022);
and U183 (N_183,In_604,In_895);
or U184 (N_184,In_987,In_1894);
and U185 (N_185,In_943,In_2708);
or U186 (N_186,In_2839,In_1068);
nor U187 (N_187,In_1118,In_2479);
or U188 (N_188,In_1643,In_810);
and U189 (N_189,In_1798,In_1296);
xor U190 (N_190,In_188,In_950);
or U191 (N_191,In_2060,In_982);
and U192 (N_192,In_1841,In_263);
or U193 (N_193,In_260,In_164);
or U194 (N_194,In_1192,In_301);
xor U195 (N_195,In_2326,In_138);
or U196 (N_196,In_1371,In_1558);
nor U197 (N_197,In_332,In_739);
nor U198 (N_198,In_230,In_1424);
xnor U199 (N_199,In_2047,In_2607);
nor U200 (N_200,In_2198,In_2007);
nand U201 (N_201,In_152,In_113);
nand U202 (N_202,In_2110,In_771);
nand U203 (N_203,In_1217,In_355);
or U204 (N_204,In_2427,In_2578);
and U205 (N_205,In_2102,In_2250);
and U206 (N_206,In_1723,In_1966);
nor U207 (N_207,In_238,In_1200);
nor U208 (N_208,In_1402,In_1779);
xnor U209 (N_209,In_843,In_201);
xnor U210 (N_210,In_2203,In_2010);
or U211 (N_211,In_597,In_1811);
nand U212 (N_212,In_458,In_122);
and U213 (N_213,In_2054,In_2294);
or U214 (N_214,In_2734,In_2959);
nor U215 (N_215,In_2156,In_2905);
and U216 (N_216,In_2629,In_2787);
xor U217 (N_217,In_251,In_966);
nor U218 (N_218,In_258,In_224);
xor U219 (N_219,In_1413,In_837);
xnor U220 (N_220,In_2810,In_1786);
and U221 (N_221,In_1896,In_1230);
nor U222 (N_222,In_879,In_1756);
nor U223 (N_223,In_2209,In_777);
and U224 (N_224,In_1790,In_2606);
or U225 (N_225,In_1084,In_1349);
nor U226 (N_226,In_2098,In_2710);
nand U227 (N_227,In_732,In_2534);
xor U228 (N_228,In_1274,In_211);
nand U229 (N_229,In_2763,In_270);
and U230 (N_230,In_2740,In_1758);
nor U231 (N_231,In_779,In_1476);
or U232 (N_232,In_1842,In_2036);
xnor U233 (N_233,In_2058,In_2276);
xnor U234 (N_234,In_2628,In_2788);
nand U235 (N_235,In_2219,In_830);
xnor U236 (N_236,In_2315,In_2519);
xnor U237 (N_237,In_865,In_2379);
and U238 (N_238,In_176,In_1797);
nand U239 (N_239,In_2693,In_2828);
nand U240 (N_240,In_2420,In_2263);
nand U241 (N_241,In_1281,In_1014);
and U242 (N_242,In_2134,In_1815);
xor U243 (N_243,In_1699,In_205);
nand U244 (N_244,In_992,In_1679);
nand U245 (N_245,In_643,In_891);
or U246 (N_246,In_1598,In_1403);
nand U247 (N_247,In_2639,In_582);
or U248 (N_248,In_750,In_2471);
and U249 (N_249,In_1715,In_647);
nand U250 (N_250,In_1943,In_1233);
nor U251 (N_251,In_2844,In_1980);
xnor U252 (N_252,In_745,In_477);
or U253 (N_253,In_2696,In_2083);
or U254 (N_254,In_1466,In_802);
and U255 (N_255,In_2667,In_35);
or U256 (N_256,In_2354,In_821);
nor U257 (N_257,In_2278,In_839);
nor U258 (N_258,In_25,In_524);
nor U259 (N_259,In_1066,In_2824);
xnor U260 (N_260,In_305,In_2413);
nor U261 (N_261,In_1431,In_2316);
xnor U262 (N_262,In_328,In_705);
xnor U263 (N_263,In_1338,In_1917);
xor U264 (N_264,In_1220,In_816);
nand U265 (N_265,In_571,In_2408);
and U266 (N_266,In_186,In_159);
and U267 (N_267,In_1250,In_50);
and U268 (N_268,In_1451,In_2831);
and U269 (N_269,In_1702,In_1289);
xor U270 (N_270,In_939,In_1500);
xor U271 (N_271,In_2691,In_2850);
and U272 (N_272,In_404,In_1528);
or U273 (N_273,In_2758,In_2474);
and U274 (N_274,In_1018,In_1240);
nand U275 (N_275,In_2637,In_2120);
and U276 (N_276,In_2630,In_2168);
nand U277 (N_277,In_1392,In_553);
xnor U278 (N_278,In_1522,In_9);
and U279 (N_279,In_2600,In_2995);
nor U280 (N_280,In_533,In_283);
nor U281 (N_281,In_1262,In_1100);
nand U282 (N_282,In_2176,In_324);
or U283 (N_283,In_1196,In_1426);
xor U284 (N_284,In_2753,In_1843);
or U285 (N_285,In_2105,In_902);
or U286 (N_286,In_2025,In_2738);
and U287 (N_287,In_2631,In_850);
xnor U288 (N_288,In_1700,In_2685);
nor U289 (N_289,In_1043,In_1156);
nand U290 (N_290,In_1026,In_1136);
nor U291 (N_291,In_194,In_2565);
and U292 (N_292,In_851,In_1739);
or U293 (N_293,In_912,In_1944);
nor U294 (N_294,In_1208,In_2152);
xor U295 (N_295,In_56,In_2711);
nand U296 (N_296,In_2267,In_1658);
nand U297 (N_297,In_800,In_783);
nand U298 (N_298,In_2881,In_536);
nand U299 (N_299,In_146,In_1218);
xnor U300 (N_300,In_1963,In_2902);
nand U301 (N_301,In_75,In_884);
nor U302 (N_302,In_1335,In_727);
or U303 (N_303,In_956,In_2643);
or U304 (N_304,In_2649,In_8);
xnor U305 (N_305,In_2022,In_2681);
xnor U306 (N_306,In_1641,In_473);
xor U307 (N_307,In_1886,In_2337);
and U308 (N_308,In_466,In_1572);
or U309 (N_309,In_2533,In_2938);
or U310 (N_310,In_18,In_2956);
nand U311 (N_311,In_2634,In_285);
nand U312 (N_312,In_1997,In_341);
xor U313 (N_313,In_756,In_2392);
xor U314 (N_314,In_204,In_2733);
and U315 (N_315,In_2971,In_2418);
or U316 (N_316,In_2598,In_2170);
or U317 (N_317,In_2447,In_1935);
xnor U318 (N_318,In_2975,In_2679);
and U319 (N_319,In_242,In_2188);
nor U320 (N_320,In_927,In_2013);
and U321 (N_321,In_580,In_2827);
or U322 (N_322,In_1989,In_2243);
nor U323 (N_323,In_2695,In_1749);
or U324 (N_324,In_1671,In_424);
nor U325 (N_325,In_2087,In_1009);
nor U326 (N_326,In_2046,In_620);
and U327 (N_327,In_2384,In_805);
nor U328 (N_328,In_1269,In_1428);
or U329 (N_329,In_2065,In_2211);
nor U330 (N_330,In_1260,In_1390);
and U331 (N_331,In_502,In_141);
nand U332 (N_332,In_1649,In_814);
and U333 (N_333,In_2445,In_1236);
and U334 (N_334,In_602,In_2836);
nand U335 (N_335,In_2311,In_2508);
and U336 (N_336,In_2342,In_467);
xnor U337 (N_337,In_2339,In_2993);
or U338 (N_338,In_1962,In_2303);
xnor U339 (N_339,In_1635,In_557);
nand U340 (N_340,In_2964,In_735);
nand U341 (N_341,In_958,In_474);
and U342 (N_342,In_2870,In_2988);
or U343 (N_343,In_618,In_63);
nor U344 (N_344,In_128,In_2147);
and U345 (N_345,In_860,In_2597);
nor U346 (N_346,In_2857,In_1703);
xnor U347 (N_347,In_1806,In_483);
nand U348 (N_348,In_1918,In_650);
xnor U349 (N_349,In_1680,In_731);
xor U350 (N_350,In_2346,In_1222);
and U351 (N_351,In_679,In_798);
nor U352 (N_352,In_292,In_1122);
xnor U353 (N_353,In_2797,In_1440);
or U354 (N_354,In_2401,In_1740);
and U355 (N_355,In_708,In_1373);
or U356 (N_356,In_476,In_624);
and U357 (N_357,In_1135,In_736);
or U358 (N_358,In_1870,In_295);
nand U359 (N_359,In_2658,In_887);
or U360 (N_360,In_1824,In_1527);
and U361 (N_361,In_1686,In_243);
xnor U362 (N_362,In_1430,In_232);
nor U363 (N_363,In_2555,In_2089);
and U364 (N_364,In_1246,In_2666);
nand U365 (N_365,In_933,In_2771);
or U366 (N_366,In_2095,In_1461);
nand U367 (N_367,In_1543,In_910);
nand U368 (N_368,In_1017,In_1952);
xnor U369 (N_369,In_478,In_1307);
xor U370 (N_370,In_2414,In_2889);
or U371 (N_371,In_856,In_2702);
nor U372 (N_372,In_2609,In_2397);
nand U373 (N_373,In_655,In_2101);
or U374 (N_374,In_1186,In_758);
or U375 (N_375,In_683,In_1975);
and U376 (N_376,In_2642,In_1394);
and U377 (N_377,In_1556,In_1463);
or U378 (N_378,In_425,In_2715);
and U379 (N_379,In_1615,In_1887);
nor U380 (N_380,In_1099,In_161);
nor U381 (N_381,In_1675,In_1407);
xnor U382 (N_382,In_2227,In_511);
or U383 (N_383,In_1873,In_707);
nor U384 (N_384,In_1631,In_2405);
and U385 (N_385,In_281,In_2736);
or U386 (N_386,In_119,In_2823);
nand U387 (N_387,In_1545,In_1532);
and U388 (N_388,In_364,In_931);
and U389 (N_389,In_2754,In_178);
xor U390 (N_390,In_768,In_1879);
nand U391 (N_391,In_578,In_1915);
xnor U392 (N_392,In_92,In_2553);
or U393 (N_393,In_1601,In_1357);
nand U394 (N_394,In_1866,In_2714);
xnor U395 (N_395,In_2750,In_1415);
and U396 (N_396,In_436,In_330);
and U397 (N_397,In_1884,In_619);
nand U398 (N_398,In_1688,In_2400);
or U399 (N_399,In_2603,In_2983);
or U400 (N_400,In_1140,In_1667);
nand U401 (N_401,In_2871,In_2561);
or U402 (N_402,In_2946,In_2931);
xnor U403 (N_403,In_1232,In_318);
or U404 (N_404,In_319,In_1689);
nand U405 (N_405,In_2622,In_2847);
or U406 (N_406,In_2184,In_2527);
or U407 (N_407,In_2493,In_1107);
nand U408 (N_408,In_863,In_2873);
or U409 (N_409,In_722,In_1607);
or U410 (N_410,In_2459,In_2672);
nor U411 (N_411,In_279,In_1245);
nand U412 (N_412,In_367,In_1990);
nor U413 (N_413,In_1549,In_1044);
nand U414 (N_414,In_1998,In_2506);
and U415 (N_415,In_124,In_72);
and U416 (N_416,In_2320,In_660);
and U417 (N_417,In_378,In_1254);
and U418 (N_418,In_2497,In_598);
xor U419 (N_419,In_7,In_445);
nor U420 (N_420,In_1423,In_623);
xor U421 (N_421,In_28,In_60);
and U422 (N_422,In_2854,In_2976);
xnor U423 (N_423,In_2996,In_475);
xor U424 (N_424,In_2372,In_1344);
nand U425 (N_425,In_532,In_2720);
nor U426 (N_426,In_1243,In_2572);
nor U427 (N_427,In_2632,In_1442);
xnor U428 (N_428,In_947,In_1382);
or U429 (N_429,In_2288,In_2920);
and U430 (N_430,In_273,In_2577);
nor U431 (N_431,In_1361,In_1621);
nand U432 (N_432,In_2846,In_1585);
xnor U433 (N_433,In_1694,In_1375);
xor U434 (N_434,In_1080,In_1803);
nor U435 (N_435,In_2653,In_2657);
xor U436 (N_436,In_1946,In_401);
or U437 (N_437,In_131,In_1011);
nor U438 (N_438,In_1923,In_2344);
xnor U439 (N_439,In_200,In_221);
xor U440 (N_440,In_156,In_1057);
xnor U441 (N_441,In_2402,In_529);
nor U442 (N_442,In_1184,In_773);
nand U443 (N_443,In_1225,In_2762);
nand U444 (N_444,In_1512,In_608);
and U445 (N_445,In_459,In_796);
and U446 (N_446,In_759,In_1332);
and U447 (N_447,In_1566,In_2820);
nand U448 (N_448,In_645,In_2214);
nand U449 (N_449,In_1496,In_2778);
xor U450 (N_450,In_2950,In_2324);
nand U451 (N_451,In_954,In_434);
xor U452 (N_452,In_897,In_2333);
and U453 (N_453,In_1224,In_78);
nand U454 (N_454,In_1813,In_1846);
or U455 (N_455,In_701,In_2535);
and U456 (N_456,In_2335,In_2285);
and U457 (N_457,In_2255,In_1855);
and U458 (N_458,In_2869,In_1048);
nand U459 (N_459,In_1279,In_1452);
and U460 (N_460,In_2389,In_1397);
xor U461 (N_461,In_2257,In_621);
or U462 (N_462,In_1529,In_2298);
and U463 (N_463,In_1016,In_1328);
nand U464 (N_464,In_1125,In_1172);
or U465 (N_465,In_2197,In_634);
and U466 (N_466,In_872,In_272);
and U467 (N_467,In_246,In_422);
nor U468 (N_468,In_1213,In_937);
or U469 (N_469,In_1718,In_244);
or U470 (N_470,In_180,In_261);
xor U471 (N_471,In_2489,In_2246);
nor U472 (N_472,In_1376,In_1151);
or U473 (N_473,In_2928,In_1031);
nor U474 (N_474,In_2064,In_1345);
and U475 (N_475,In_222,In_2932);
and U476 (N_476,In_2941,In_312);
or U477 (N_477,In_407,In_554);
and U478 (N_478,In_2367,In_2399);
or U479 (N_479,In_2023,In_1298);
nor U480 (N_480,In_1895,In_157);
xor U481 (N_481,In_2703,In_2688);
xor U482 (N_482,In_2248,In_1901);
or U483 (N_483,In_878,In_2934);
and U484 (N_484,In_1059,In_1809);
nor U485 (N_485,In_453,In_955);
nand U486 (N_486,In_1636,In_2562);
xnor U487 (N_487,In_2586,In_1924);
nand U488 (N_488,In_2242,In_1652);
nand U489 (N_489,In_1907,In_26);
nand U490 (N_490,In_1105,In_1697);
xnor U491 (N_491,In_565,In_550);
and U492 (N_492,In_2664,In_253);
nand U493 (N_493,In_1331,In_2464);
nor U494 (N_494,In_2003,In_1453);
nor U495 (N_495,In_1698,In_2500);
nor U496 (N_496,In_1893,In_573);
nand U497 (N_497,In_2393,In_1589);
nor U498 (N_498,In_2879,In_2386);
nand U499 (N_499,In_1177,In_684);
or U500 (N_500,In_544,In_754);
or U501 (N_501,In_537,In_946);
or U502 (N_502,In_350,In_2712);
nor U503 (N_503,In_1696,In_593);
nand U504 (N_504,In_2138,In_462);
xor U505 (N_505,In_1787,In_1121);
and U506 (N_506,In_2648,In_1253);
xor U507 (N_507,In_1903,In_339);
xor U508 (N_508,In_1103,In_479);
or U509 (N_509,In_2041,In_2108);
nand U510 (N_510,In_1102,In_760);
xnor U511 (N_511,In_455,In_1318);
xor U512 (N_512,In_334,In_36);
and U513 (N_513,In_2014,In_2544);
xor U514 (N_514,In_1420,In_236);
and U515 (N_515,In_1353,In_2528);
nor U516 (N_516,In_1406,In_2765);
nand U517 (N_517,In_807,In_1761);
or U518 (N_518,In_2646,In_1651);
and U519 (N_519,In_1821,In_452);
or U520 (N_520,In_1954,In_749);
and U521 (N_521,In_2300,In_2016);
or U522 (N_522,In_2725,In_197);
xnor U523 (N_523,In_248,In_2998);
nand U524 (N_524,In_496,In_2476);
and U525 (N_525,In_2615,In_315);
nand U526 (N_526,In_642,In_686);
xor U527 (N_527,In_1619,In_415);
nand U528 (N_528,In_158,In_1021);
and U529 (N_529,In_2742,In_361);
nand U530 (N_530,In_1486,In_2469);
or U531 (N_531,In_109,In_2546);
and U532 (N_532,In_2453,In_2129);
nor U533 (N_533,In_173,In_1065);
nand U534 (N_534,In_465,In_1860);
or U535 (N_535,In_357,In_151);
nand U536 (N_536,In_820,In_2721);
xor U537 (N_537,In_162,In_1764);
and U538 (N_538,In_929,In_1111);
or U539 (N_539,In_2764,In_1091);
and U540 (N_540,In_86,In_2150);
or U541 (N_541,In_2332,In_2724);
nor U542 (N_542,In_170,In_1053);
nand U543 (N_543,In_1662,In_1263);
or U544 (N_544,In_1323,In_2874);
nor U545 (N_545,In_2309,In_1563);
or U546 (N_546,In_2394,In_2204);
or U547 (N_547,In_1835,In_2660);
and U548 (N_548,In_2699,In_2548);
or U549 (N_549,In_789,In_603);
xnor U550 (N_550,In_1479,In_2958);
nand U551 (N_551,In_2334,In_82);
nor U552 (N_552,In_2957,In_2760);
and U553 (N_553,In_1355,In_1432);
nand U554 (N_554,In_2000,In_111);
and U555 (N_555,In_2074,In_241);
nor U556 (N_556,In_2767,In_2997);
nand U557 (N_557,In_1546,In_2811);
or U558 (N_558,In_1816,In_1443);
or U559 (N_559,In_2930,In_1005);
xnor U560 (N_560,In_198,In_1913);
or U561 (N_561,In_1366,In_1215);
or U562 (N_562,In_2929,In_2365);
or U563 (N_563,In_1271,In_1926);
xor U564 (N_564,In_1802,In_1120);
and U565 (N_565,In_595,In_1465);
and U566 (N_566,In_2321,In_2872);
nor U567 (N_567,In_1704,In_14);
nor U568 (N_568,In_527,In_44);
or U569 (N_569,In_1773,In_2913);
nor U570 (N_570,In_2062,In_793);
nand U571 (N_571,In_922,In_2944);
and U572 (N_572,In_234,In_217);
or U573 (N_573,In_486,In_226);
xnor U574 (N_574,In_349,In_1650);
or U575 (N_575,In_1677,In_1197);
or U576 (N_576,In_1109,In_1174);
nor U577 (N_577,In_2601,In_2160);
nor U578 (N_578,In_2803,In_2918);
xor U579 (N_579,In_1448,In_2893);
xor U580 (N_580,In_1726,In_2713);
nand U581 (N_581,In_1474,In_2654);
and U582 (N_582,In_165,In_1470);
nor U583 (N_583,In_2269,In_1534);
or U584 (N_584,In_406,In_437);
and U585 (N_585,In_1827,In_2571);
nor U586 (N_586,In_2056,In_1788);
or U587 (N_587,In_1804,In_2868);
and U588 (N_588,In_1507,In_2436);
nor U589 (N_589,In_1123,In_2167);
nand U590 (N_590,In_2270,In_1904);
and U591 (N_591,In_99,In_2936);
xor U592 (N_592,In_1385,In_2723);
and U593 (N_593,In_2730,In_2251);
nor U594 (N_594,In_2757,In_175);
and U595 (N_595,In_2927,In_2935);
or U596 (N_596,In_39,In_57);
or U597 (N_597,In_267,In_2130);
xnor U598 (N_598,In_2682,In_2888);
and U599 (N_599,In_47,In_150);
nor U600 (N_600,In_1672,In_930);
or U601 (N_601,In_1129,In_1164);
nor U602 (N_602,In_321,In_360);
nand U603 (N_603,In_2650,In_555);
or U604 (N_604,In_1288,In_1515);
xor U605 (N_605,In_915,In_2829);
or U606 (N_606,In_1456,In_2747);
nand U607 (N_607,In_52,In_1818);
nor U608 (N_608,In_2208,In_1096);
nor U609 (N_609,In_117,In_2878);
nand U610 (N_610,In_2545,In_2283);
xor U611 (N_611,In_490,In_549);
nor U612 (N_612,In_2200,In_2542);
or U613 (N_613,In_1750,In_289);
xnor U614 (N_614,In_1062,In_659);
nand U615 (N_615,In_1961,In_2086);
or U616 (N_616,In_1040,In_2035);
nor U617 (N_617,In_1892,In_2511);
xor U618 (N_618,In_2391,In_400);
and U619 (N_619,In_144,In_2912);
and U620 (N_620,In_1359,In_1013);
or U621 (N_621,In_1074,In_2502);
or U622 (N_622,In_646,In_2592);
or U623 (N_623,In_885,In_358);
or U624 (N_624,In_488,In_2510);
xnor U625 (N_625,In_801,In_2233);
nor U626 (N_626,In_2705,In_2700);
and U627 (N_627,In_935,In_1731);
nand U628 (N_628,In_2604,In_1126);
nand U629 (N_629,In_2323,In_2865);
and U630 (N_630,In_2969,In_869);
nand U631 (N_631,In_1684,In_2948);
xnor U632 (N_632,In_1446,In_2785);
nor U633 (N_633,In_2991,In_2890);
and U634 (N_634,In_1971,In_1226);
nor U635 (N_635,In_1380,In_1348);
and U636 (N_636,In_2475,In_2729);
and U637 (N_637,In_2017,In_316);
and U638 (N_638,In_2328,In_697);
and U639 (N_639,In_1334,In_2148);
or U640 (N_640,In_2662,In_2774);
nor U641 (N_641,In_567,In_706);
nand U642 (N_642,In_531,In_983);
xor U643 (N_643,In_1438,In_351);
and U644 (N_644,In_974,In_1329);
nand U645 (N_645,In_240,In_2419);
nor U646 (N_646,In_1436,In_1574);
nor U647 (N_647,In_1682,In_76);
nor U648 (N_648,In_829,In_2589);
nor U649 (N_649,In_2478,In_2355);
nand U650 (N_650,In_469,In_1656);
nand U651 (N_651,In_2302,In_700);
xnor U652 (N_652,In_1852,In_1520);
and U653 (N_653,In_120,In_786);
and U654 (N_654,In_959,In_584);
nand U655 (N_655,In_2430,In_32);
nand U656 (N_656,In_1193,In_2432);
xnor U657 (N_657,In_1007,In_1488);
or U658 (N_658,In_636,In_395);
xnor U659 (N_659,In_2306,In_430);
nand U660 (N_660,In_1210,In_309);
nand U661 (N_661,In_2732,In_381);
nor U662 (N_662,In_2443,In_649);
and U663 (N_663,In_772,In_494);
nor U664 (N_664,In_84,In_1189);
or U665 (N_665,In_581,In_1861);
xor U666 (N_666,In_2537,In_278);
nand U667 (N_667,In_656,In_2775);
or U668 (N_668,In_218,In_726);
nor U669 (N_669,In_2153,In_2911);
or U670 (N_670,In_1464,In_1198);
nor U671 (N_671,In_24,In_2951);
and U672 (N_672,In_1599,In_2610);
nand U673 (N_673,In_681,In_859);
or U674 (N_674,In_2137,In_2675);
or U675 (N_675,In_1015,In_460);
or U676 (N_676,In_641,In_1906);
or U677 (N_677,In_1045,In_1781);
xnor U678 (N_678,In_1911,In_1559);
xor U679 (N_679,In_670,In_426);
xnor U680 (N_680,In_121,In_1191);
xor U681 (N_681,In_2079,In_609);
or U682 (N_682,In_944,In_300);
xor U683 (N_683,In_2919,In_1336);
or U684 (N_684,In_2531,In_1685);
and U685 (N_685,In_1085,In_761);
nand U686 (N_686,In_2694,In_2456);
or U687 (N_687,In_385,In_2641);
and U688 (N_688,In_2451,In_738);
or U689 (N_689,In_1547,In_2238);
and U690 (N_690,In_55,In_1733);
xor U691 (N_691,In_1795,In_988);
xnor U692 (N_692,In_2006,In_1964);
xor U693 (N_693,In_181,In_905);
or U694 (N_694,In_397,In_600);
nand U695 (N_695,In_396,In_2135);
and U696 (N_696,In_1889,In_1665);
xor U697 (N_697,In_457,In_552);
xnor U698 (N_698,In_714,In_2141);
nand U699 (N_699,In_1227,In_136);
xnor U700 (N_700,In_2244,In_2987);
nand U701 (N_701,In_965,In_721);
nor U702 (N_702,In_518,In_41);
nor U703 (N_703,In_2599,In_2549);
nand U704 (N_704,In_1064,In_2515);
xnor U705 (N_705,In_2295,In_2517);
nor U706 (N_706,In_1727,In_2968);
or U707 (N_707,In_1095,In_1774);
or U708 (N_708,In_168,In_2292);
nand U709 (N_709,In_1050,In_2024);
and U710 (N_710,In_1993,In_538);
xnor U711 (N_711,In_1669,In_1106);
and U712 (N_712,In_1169,In_2652);
nand U713 (N_713,In_413,In_971);
and U714 (N_714,In_1616,In_147);
and U715 (N_715,In_1083,In_2450);
or U716 (N_716,In_2026,In_717);
xor U717 (N_717,In_33,In_2199);
or U718 (N_718,In_1504,In_2155);
and U719 (N_719,In_2448,In_1159);
and U720 (N_720,In_352,In_782);
xor U721 (N_721,In_421,In_666);
or U722 (N_722,In_2043,In_853);
or U723 (N_723,In_2050,In_2186);
or U724 (N_724,In_214,In_2136);
xnor U725 (N_725,In_2,In_2072);
or U726 (N_726,In_1327,In_1216);
xnor U727 (N_727,In_689,In_337);
nor U728 (N_728,In_2808,In_2818);
nand U729 (N_729,In_2627,In_149);
xor U730 (N_730,In_228,In_1768);
xor U731 (N_731,In_2687,In_1967);
nand U732 (N_732,In_2063,In_989);
nor U733 (N_733,In_2690,In_2636);
nor U734 (N_734,In_491,In_2570);
xor U735 (N_735,In_2618,In_1141);
and U736 (N_736,In_508,In_811);
nor U737 (N_737,In_2566,In_110);
or U738 (N_738,In_1712,In_2191);
xnor U739 (N_739,In_6,In_2433);
nor U740 (N_740,In_813,In_2115);
xnor U741 (N_741,In_1383,In_2773);
nor U742 (N_742,In_1237,In_1940);
and U743 (N_743,In_2274,In_2287);
and U744 (N_744,In_2018,In_1139);
nand U745 (N_745,In_815,In_2206);
or U746 (N_746,In_2260,In_133);
or U747 (N_747,In_42,In_2312);
nor U748 (N_748,In_1239,In_1020);
and U749 (N_749,In_1265,In_1751);
or U750 (N_750,In_828,In_1165);
nand U751 (N_751,In_2259,In_2842);
and U752 (N_752,In_2825,In_2329);
and U753 (N_753,In_784,In_2856);
nor U754 (N_754,In_210,In_1707);
nand U755 (N_755,In_972,In_685);
nand U756 (N_756,In_495,In_2579);
and U757 (N_757,In_1377,In_728);
nand U758 (N_758,In_569,In_88);
xnor U759 (N_759,In_37,In_1584);
or U760 (N_760,In_108,In_1155);
nand U761 (N_761,In_1769,In_64);
and U762 (N_762,In_209,In_2516);
xnor U763 (N_763,In_1266,In_2743);
nand U764 (N_764,In_545,In_410);
nor U765 (N_765,In_461,In_93);
and U766 (N_766,In_202,In_572);
nor U767 (N_767,In_1295,In_1509);
nor U768 (N_768,In_368,In_2965);
and U769 (N_769,In_441,In_2947);
nand U770 (N_770,In_227,In_612);
or U771 (N_771,In_2776,In_299);
and U772 (N_772,In_2077,In_2822);
nand U773 (N_773,In_53,In_2179);
nor U774 (N_774,In_1663,In_1082);
nand U775 (N_775,In_2340,In_719);
and U776 (N_776,In_2132,In_2819);
nand U777 (N_777,In_2375,In_2106);
or U778 (N_778,In_1745,In_1600);
and U779 (N_779,In_806,In_2633);
nand U780 (N_780,In_1833,In_456);
and U781 (N_781,In_635,In_2815);
xor U782 (N_782,In_2945,In_1931);
xnor U783 (N_783,In_1203,In_448);
xnor U784 (N_784,In_2482,In_1738);
and U785 (N_785,In_566,In_1389);
and U786 (N_786,In_2124,In_1365);
or U787 (N_787,In_129,In_1648);
and U788 (N_788,In_2884,In_320);
and U789 (N_789,In_2900,In_586);
and U790 (N_790,In_2547,In_2368);
nand U791 (N_791,In_2795,In_2605);
xnor U792 (N_792,In_59,In_43);
or U793 (N_793,In_2378,In_2620);
xor U794 (N_794,In_919,In_123);
nand U795 (N_795,In_118,In_2655);
xnor U796 (N_796,In_2205,In_2434);
and U797 (N_797,In_855,In_2756);
or U798 (N_798,In_2149,In_1987);
or U799 (N_799,In_2439,In_716);
or U800 (N_800,In_2505,In_858);
nor U801 (N_801,In_2100,In_2780);
nand U802 (N_802,In_329,In_2037);
nor U803 (N_803,In_1983,In_629);
or U804 (N_804,In_1792,In_1897);
and U805 (N_805,In_747,In_2480);
nor U806 (N_806,In_2728,In_2689);
and U807 (N_807,In_2853,In_2182);
xnor U808 (N_808,In_492,In_673);
nor U809 (N_809,In_237,In_640);
nand U810 (N_810,In_1358,In_2560);
nand U811 (N_811,In_1539,In_2943);
xnor U812 (N_812,In_1668,In_1984);
or U813 (N_813,In_1916,In_1248);
and U814 (N_814,In_1885,In_1201);
xor U815 (N_815,In_1181,In_484);
nor U816 (N_816,In_2789,In_1419);
or U817 (N_817,In_2452,In_1932);
or U818 (N_818,In_2090,In_2118);
nand U819 (N_819,In_2088,In_2875);
and U820 (N_820,In_1951,In_2313);
or U821 (N_821,In_2580,In_2256);
or U822 (N_822,In_1627,In_2145);
and U823 (N_823,In_142,In_1163);
xnor U824 (N_824,In_1324,In_219);
nor U825 (N_825,In_1483,In_345);
and U826 (N_826,In_2009,In_464);
nand U827 (N_827,In_577,In_2224);
xor U828 (N_828,In_519,In_2647);
xor U829 (N_829,In_1754,In_1137);
or U830 (N_830,In_1175,In_1497);
or U831 (N_831,In_1597,In_1511);
nand U832 (N_832,In_1368,In_1965);
or U833 (N_833,In_2640,In_2099);
xnor U834 (N_834,In_613,In_962);
nand U835 (N_835,In_599,In_130);
nor U836 (N_836,In_2463,In_419);
xnor U837 (N_837,In_112,In_2005);
nor U838 (N_838,In_1859,In_1853);
xor U839 (N_839,In_2752,In_1880);
xnor U840 (N_840,In_1729,In_1205);
nand U841 (N_841,In_1772,In_2240);
xnor U842 (N_842,In_2261,In_2665);
xor U843 (N_843,In_1055,In_191);
xor U844 (N_844,In_501,In_1591);
or U845 (N_845,In_849,In_2053);
nand U846 (N_846,In_723,In_105);
nor U847 (N_847,In_1576,In_2915);
nand U848 (N_848,In_1493,In_625);
or U849 (N_849,In_1150,In_1273);
nand U850 (N_850,In_766,In_1211);
or U851 (N_851,In_757,In_1114);
and U852 (N_852,In_1153,In_985);
or U853 (N_853,In_563,In_369);
nand U854 (N_854,In_953,In_1812);
and U855 (N_855,In_2237,In_936);
or U856 (N_856,In_275,In_1959);
and U857 (N_857,In_322,In_1450);
nor U858 (N_858,In_2187,In_420);
xnor U859 (N_859,In_1728,In_16);
nand U860 (N_860,In_622,In_2859);
or U861 (N_861,In_1721,In_2425);
or U862 (N_862,In_2751,In_2520);
and U863 (N_863,In_1297,In_2759);
xor U864 (N_864,In_1851,In_1544);
nand U865 (N_865,In_1542,In_2458);
nor U866 (N_866,In_1612,In_1073);
and U867 (N_867,In_1995,In_1747);
xor U868 (N_868,In_2461,In_2611);
and U869 (N_869,In_1401,In_500);
nor U870 (N_870,In_1410,In_791);
or U871 (N_871,In_383,In_135);
and U872 (N_872,In_993,In_154);
xor U873 (N_873,In_2624,In_957);
and U874 (N_874,In_1161,In_2575);
or U875 (N_875,In_564,In_2181);
and U876 (N_876,In_83,In_1969);
nor U877 (N_877,In_2669,In_695);
or U878 (N_878,In_2216,In_2011);
and U879 (N_879,In_2862,In_2989);
and U880 (N_880,In_2194,In_1902);
nand U881 (N_881,In_2894,In_2381);
xor U882 (N_882,In_1832,In_1282);
and U883 (N_883,In_1571,In_2671);
xnor U884 (N_884,In_1199,In_12);
and U885 (N_885,In_2901,In_179);
and U886 (N_886,In_831,In_216);
nor U887 (N_887,In_2612,In_1570);
and U888 (N_888,In_1760,In_1108);
xor U889 (N_889,In_1145,In_11);
nor U890 (N_890,In_1505,In_2863);
nand U891 (N_891,In_2748,In_2092);
nor U892 (N_892,In_2040,In_239);
and U893 (N_893,In_2659,In_1834);
nand U894 (N_894,In_2477,In_298);
or U895 (N_895,In_730,In_797);
and U896 (N_896,In_2437,In_409);
xor U897 (N_897,In_1124,In_2582);
xor U898 (N_898,In_1647,In_2698);
or U899 (N_899,In_2504,In_1819);
and U900 (N_900,In_1351,In_1553);
xnor U901 (N_901,In_1304,In_2351);
xor U902 (N_902,In_1491,In_1996);
nand U903 (N_903,In_468,In_2999);
and U904 (N_904,In_1093,In_1725);
xor U905 (N_905,In_1801,In_2885);
and U906 (N_906,In_720,In_1370);
nand U907 (N_907,In_2008,In_2159);
and U908 (N_908,In_432,In_1793);
nor U909 (N_909,In_941,In_2417);
nand U910 (N_910,In_507,In_2343);
xor U911 (N_911,In_2981,In_1791);
xor U912 (N_912,In_2151,In_746);
nand U913 (N_913,In_2262,In_1632);
nand U914 (N_914,In_1625,In_675);
nor U915 (N_915,In_2498,In_1555);
nor U916 (N_916,In_389,In_2921);
xnor U917 (N_917,In_1350,In_393);
xnor U918 (N_918,In_2232,In_2522);
nand U919 (N_919,In_914,In_1711);
nand U920 (N_920,In_1732,In_1352);
xnor U921 (N_921,In_1910,In_2078);
xnor U922 (N_922,In_1929,In_1565);
nand U923 (N_923,In_403,In_1092);
nand U924 (N_924,In_1742,In_1828);
xor U925 (N_925,In_1927,In_790);
and U926 (N_926,In_900,In_963);
nor U927 (N_927,In_269,In_778);
nand U928 (N_928,In_2277,In_427);
or U929 (N_929,In_2673,In_1330);
nor U930 (N_930,In_848,In_1994);
or U931 (N_931,In_1501,In_984);
nor U932 (N_932,In_1414,In_1367);
xnor U933 (N_933,In_414,In_1593);
or U934 (N_934,In_1343,In_1259);
xnor U935 (N_935,In_2737,In_2395);
or U936 (N_936,In_1590,In_819);
nand U937 (N_937,In_2532,In_1595);
nand U938 (N_938,In_2552,In_1149);
and U939 (N_939,In_973,In_1069);
nand U940 (N_940,In_980,In_2977);
and U941 (N_941,In_2557,In_864);
nor U942 (N_942,In_296,In_1468);
nor U943 (N_943,In_692,In_2923);
and U944 (N_944,In_1473,In_1034);
and U945 (N_945,In_2530,In_2855);
xor U946 (N_946,In_1098,In_160);
or U947 (N_947,In_291,In_1404);
nand U948 (N_948,In_540,In_2183);
nor U949 (N_949,In_2066,In_1611);
nand U950 (N_950,In_663,In_1128);
and U951 (N_951,In_1999,In_235);
xnor U952 (N_952,In_2140,In_2234);
or U953 (N_953,In_1862,In_548);
or U954 (N_954,In_1538,In_177);
xor U955 (N_955,In_648,In_1876);
xor U956 (N_956,In_2364,In_1630);
xnor U957 (N_957,In_522,In_268);
xor U958 (N_958,In_1374,In_2860);
or U959 (N_959,In_1484,In_431);
and U960 (N_960,In_840,In_225);
nand U961 (N_961,In_2499,In_762);
or U962 (N_962,In_1868,In_703);
xnor U963 (N_963,In_857,In_1028);
nor U964 (N_964,In_1449,In_1056);
and U965 (N_965,In_392,In_1550);
nor U966 (N_966,In_2409,In_1);
and U967 (N_967,In_423,In_2492);
nand U968 (N_968,In_2651,In_2897);
xnor U969 (N_969,In_2851,In_2157);
and U970 (N_970,In_2407,In_2307);
nor U971 (N_971,In_470,In_388);
xor U972 (N_972,In_2718,In_2460);
xnor U973 (N_973,In_2143,In_1582);
nand U974 (N_974,In_2380,In_809);
or U975 (N_975,In_2591,In_1687);
and U976 (N_976,In_1489,In_2094);
xnor U977 (N_977,In_698,In_1810);
and U978 (N_978,In_1052,In_812);
nand U979 (N_979,In_568,In_1280);
or U980 (N_980,In_1974,In_2796);
nor U981 (N_981,In_2812,In_132);
xor U982 (N_982,In_2028,In_1460);
nor U983 (N_983,In_1660,In_639);
xor U984 (N_984,In_886,In_116);
xor U985 (N_985,In_1767,In_651);
and U986 (N_986,In_2325,In_882);
nand U987 (N_987,In_2523,In_2906);
nor U988 (N_988,In_2848,In_384);
or U989 (N_989,In_2596,In_2926);
xor U990 (N_990,In_2426,In_1617);
nand U991 (N_991,In_1278,In_2518);
and U992 (N_992,In_2761,In_2896);
xor U993 (N_993,In_1387,In_49);
nor U994 (N_994,In_1386,In_2223);
or U995 (N_995,In_2264,In_1131);
xor U996 (N_996,In_755,In_2429);
nor U997 (N_997,In_967,In_2960);
nand U998 (N_998,In_861,In_2412);
nand U999 (N_999,In_923,In_1655);
nand U1000 (N_1000,N_650,N_356);
or U1001 (N_1001,N_418,In_1427);
nand U1002 (N_1002,N_141,In_213);
and U1003 (N_1003,In_1033,N_182);
nor U1004 (N_1004,N_961,In_1132);
and U1005 (N_1005,In_288,In_2961);
or U1006 (N_1006,N_572,In_2073);
xor U1007 (N_1007,In_1146,In_1633);
nor U1008 (N_1008,In_832,N_382);
xnor U1009 (N_1009,N_478,In_303);
nor U1010 (N_1010,N_488,N_213);
xnor U1011 (N_1011,N_968,N_530);
or U1012 (N_1012,N_482,N_712);
xor U1013 (N_1013,N_468,N_722);
nand U1014 (N_1014,N_810,N_53);
and U1015 (N_1015,In_1054,In_2174);
nor U1016 (N_1016,N_593,N_937);
nand U1017 (N_1017,In_489,In_1956);
nand U1018 (N_1018,N_951,In_1981);
xor U1019 (N_1019,In_1716,N_533);
nor U1020 (N_1020,N_241,In_2543);
nor U1021 (N_1021,In_1369,N_280);
nand U1022 (N_1022,In_22,In_79);
nor U1023 (N_1023,In_402,In_2403);
nand U1024 (N_1024,N_105,In_2834);
nand U1025 (N_1025,In_189,In_2784);
and U1026 (N_1026,N_667,In_979);
xnor U1027 (N_1027,In_2907,In_1454);
nand U1028 (N_1028,In_114,N_313);
nand U1029 (N_1029,In_2424,N_691);
nand U1030 (N_1030,N_491,In_1719);
nand U1031 (N_1031,In_190,In_911);
nor U1032 (N_1032,N_877,N_658);
nand U1033 (N_1033,N_481,In_19);
nand U1034 (N_1034,In_1637,N_946);
nor U1035 (N_1035,In_2817,N_957);
xnor U1036 (N_1036,N_557,In_287);
nand U1037 (N_1037,N_293,In_1234);
xnor U1038 (N_1038,In_2195,In_2158);
xnor U1039 (N_1039,N_311,N_870);
nor U1040 (N_1040,In_2816,N_58);
or U1041 (N_1041,N_731,In_2680);
and U1042 (N_1042,In_2704,N_355);
nor U1043 (N_1043,N_871,In_1953);
nand U1044 (N_1044,In_1840,In_2861);
and U1045 (N_1045,N_333,In_1730);
nor U1046 (N_1046,In_282,In_1171);
or U1047 (N_1047,N_25,In_667);
nand U1048 (N_1048,In_1097,N_436);
or U1049 (N_1049,N_329,N_913);
xnor U1050 (N_1050,N_749,In_1303);
xor U1051 (N_1051,In_1471,N_684);
and U1052 (N_1052,In_2798,In_2165);
xor U1053 (N_1053,In_2169,In_2623);
and U1054 (N_1054,In_952,In_2801);
or U1055 (N_1055,In_1596,N_37);
or U1056 (N_1056,In_1003,In_780);
nor U1057 (N_1057,N_338,N_264);
or U1058 (N_1058,In_2877,In_1848);
or U1059 (N_1059,In_229,N_575);
nor U1060 (N_1060,N_671,In_925);
nor U1061 (N_1061,In_336,N_55);
xnor U1062 (N_1062,N_72,N_199);
nand U1063 (N_1063,In_2826,N_99);
and U1064 (N_1064,N_291,In_1548);
nand U1065 (N_1065,In_1268,In_1825);
and U1066 (N_1066,In_854,In_668);
xor U1067 (N_1067,In_674,In_881);
nor U1068 (N_1068,In_399,N_860);
or U1069 (N_1069,N_143,In_1780);
or U1070 (N_1070,In_976,In_2104);
nand U1071 (N_1071,N_197,N_777);
and U1072 (N_1072,In_1144,In_1569);
xor U1073 (N_1073,N_726,In_867);
nor U1074 (N_1074,In_153,In_338);
nand U1075 (N_1075,In_493,In_271);
and U1076 (N_1076,In_317,N_997);
nor U1077 (N_1077,N_505,In_2608);
nand U1078 (N_1078,N_545,In_61);
and U1079 (N_1079,In_66,In_2766);
xnor U1080 (N_1080,In_1152,N_631);
nand U1081 (N_1081,N_346,N_496);
or U1082 (N_1082,N_406,In_1039);
and U1083 (N_1083,In_2142,In_1775);
and U1084 (N_1084,In_2914,N_112);
nor U1085 (N_1085,In_877,N_295);
or U1086 (N_1086,N_179,N_170);
or U1087 (N_1087,In_827,In_354);
or U1088 (N_1088,N_286,N_399);
nor U1089 (N_1089,In_450,N_230);
nor U1090 (N_1090,N_655,N_892);
xor U1091 (N_1091,N_857,N_816);
and U1092 (N_1092,In_626,N_362);
and U1093 (N_1093,N_50,N_300);
and U1094 (N_1094,N_190,N_967);
nand U1095 (N_1095,In_2678,In_741);
nand U1096 (N_1096,In_2536,N_643);
xnor U1097 (N_1097,In_1519,N_63);
xnor U1098 (N_1098,N_890,N_259);
or U1099 (N_1099,N_164,In_257);
and U1100 (N_1100,N_128,In_556);
nor U1101 (N_1101,In_1580,In_617);
and U1102 (N_1102,N_352,In_2421);
or U1103 (N_1103,In_1294,N_886);
or U1104 (N_1104,In_1717,N_983);
nand U1105 (N_1105,In_1499,N_483);
nand U1106 (N_1106,In_1820,In_1856);
nand U1107 (N_1107,In_688,In_2438);
nand U1108 (N_1108,N_249,In_1890);
and U1109 (N_1109,N_203,In_883);
nand U1110 (N_1110,N_470,N_462);
nand U1111 (N_1111,N_990,In_525);
nand U1112 (N_1112,In_1101,N_986);
or U1113 (N_1113,N_570,In_2201);
or U1114 (N_1114,In_1162,In_1284);
nor U1115 (N_1115,In_744,N_15);
nand U1116 (N_1116,In_934,N_153);
or U1117 (N_1117,In_2282,N_282);
and U1118 (N_1118,In_2782,In_1817);
or U1119 (N_1119,In_1170,N_206);
and U1120 (N_1120,In_1223,In_2266);
nand U1121 (N_1121,N_212,N_517);
nor U1122 (N_1122,In_2296,In_2746);
xnor U1123 (N_1123,N_148,In_1919);
xor U1124 (N_1124,N_652,In_17);
xor U1125 (N_1125,In_2614,N_633);
nand U1126 (N_1126,N_863,In_499);
or U1127 (N_1127,In_331,In_1312);
or U1128 (N_1128,N_439,In_1858);
nor U1129 (N_1129,In_1495,N_165);
nor U1130 (N_1130,In_1299,N_403);
xnor U1131 (N_1131,In_671,N_82);
nor U1132 (N_1132,N_534,In_2202);
nand U1133 (N_1133,In_1276,N_867);
or U1134 (N_1134,In_589,In_1356);
or U1135 (N_1135,In_1185,N_939);
and U1136 (N_1136,In_0,N_642);
and U1137 (N_1137,N_612,In_1783);
and U1138 (N_1138,In_134,N_261);
xnor U1139 (N_1139,In_607,In_918);
or U1140 (N_1140,N_198,In_2481);
xor U1141 (N_1141,N_582,N_86);
or U1142 (N_1142,In_1531,In_348);
nand U1143 (N_1143,N_68,In_1614);
xor U1144 (N_1144,In_826,In_1206);
xor U1145 (N_1145,In_1455,N_525);
nor U1146 (N_1146,In_2117,In_1076);
nor U1147 (N_1147,N_150,In_1763);
xnor U1148 (N_1148,N_678,In_2514);
or U1149 (N_1149,In_2484,N_52);
or U1150 (N_1150,In_969,N_620);
nor U1151 (N_1151,N_617,N_467);
nand U1152 (N_1152,In_2904,N_409);
and U1153 (N_1153,In_596,N_110);
or U1154 (N_1154,In_2239,N_976);
nor U1155 (N_1155,N_878,In_48);
and U1156 (N_1156,N_495,N_696);
xor U1157 (N_1157,N_922,N_542);
xnor U1158 (N_1158,In_346,N_127);
nor U1159 (N_1159,In_2131,In_1933);
nor U1160 (N_1160,In_1204,In_2347);
nand U1161 (N_1161,N_24,In_680);
and U1162 (N_1162,In_2076,In_307);
or U1163 (N_1163,In_2213,N_125);
and U1164 (N_1164,N_370,In_102);
nor U1165 (N_1165,In_2509,N_502);
nor U1166 (N_1166,N_429,In_2161);
and U1167 (N_1167,N_35,N_423);
or U1168 (N_1168,N_891,N_885);
nor U1169 (N_1169,N_758,N_227);
xor U1170 (N_1170,In_1072,In_2085);
or U1171 (N_1171,In_1231,N_447);
and U1172 (N_1172,In_2416,N_177);
nand U1173 (N_1173,N_514,N_69);
nor U1174 (N_1174,In_2621,N_753);
or U1175 (N_1175,N_699,N_999);
and U1176 (N_1176,In_2581,In_1425);
xnor U1177 (N_1177,N_724,N_969);
xor U1178 (N_1178,In_2226,In_2109);
nor U1179 (N_1179,In_1908,In_1722);
nor U1180 (N_1180,In_1408,In_1928);
nor U1181 (N_1181,In_610,N_623);
or U1182 (N_1182,In_825,N_377);
nand U1183 (N_1183,In_765,N_791);
and U1184 (N_1184,N_680,N_441);
nor U1185 (N_1185,In_664,N_469);
or U1186 (N_1186,N_613,In_2677);
or U1187 (N_1187,N_344,In_1592);
nor U1188 (N_1188,In_842,N_659);
nand U1189 (N_1189,N_269,N_693);
nor U1190 (N_1190,In_570,N_500);
or U1191 (N_1191,N_455,N_140);
nor U1192 (N_1192,N_532,In_920);
xnor U1193 (N_1193,In_435,In_1242);
and U1194 (N_1194,N_40,In_1322);
or U1195 (N_1195,In_1070,N_319);
nand U1196 (N_1196,N_543,N_540);
or U1197 (N_1197,N_389,N_639);
xor U1198 (N_1198,N_769,In_65);
nand U1199 (N_1199,In_2551,In_551);
nor U1200 (N_1200,N_2,N_45);
and U1201 (N_1201,N_689,In_325);
xor U1202 (N_1202,N_762,In_382);
and U1203 (N_1203,N_49,N_460);
nor U1204 (N_1204,In_2059,In_2770);
or U1205 (N_1205,In_2030,In_310);
and U1206 (N_1206,N_438,N_87);
xnor U1207 (N_1207,In_2272,N_579);
nor U1208 (N_1208,N_827,In_1326);
nand U1209 (N_1209,N_20,N_85);
or U1210 (N_1210,In_1705,N_137);
nand U1211 (N_1211,N_771,In_921);
and U1212 (N_1212,In_245,N_869);
or U1213 (N_1213,In_1127,In_637);
xor U1214 (N_1214,In_2410,N_337);
and U1215 (N_1215,In_1004,N_432);
nor U1216 (N_1216,N_942,In_803);
nand U1217 (N_1217,In_2992,N_255);
and U1218 (N_1218,In_1209,In_2457);
nor U1219 (N_1219,N_826,N_126);
xor U1220 (N_1220,N_121,N_604);
nor U1221 (N_1221,N_861,N_859);
or U1222 (N_1222,N_433,N_506);
and U1223 (N_1223,In_1800,In_904);
xor U1224 (N_1224,In_1160,In_2744);
xnor U1225 (N_1225,N_768,In_1409);
and U1226 (N_1226,In_907,N_359);
or U1227 (N_1227,N_167,In_1513);
xnor U1228 (N_1228,N_131,In_2564);
and U1229 (N_1229,In_1467,N_522);
nor U1230 (N_1230,N_960,N_666);
xor U1231 (N_1231,In_1293,In_1681);
xnor U1232 (N_1232,In_526,N_600);
nand U1233 (N_1233,N_598,In_787);
xor U1234 (N_1234,In_1182,N_340);
and U1235 (N_1235,N_60,In_559);
nor U1236 (N_1236,N_833,N_318);
nor U1237 (N_1237,In_2783,In_503);
and U1238 (N_1238,N_670,In_2924);
and U1239 (N_1239,In_2349,In_896);
nor U1240 (N_1240,N_966,In_1937);
xor U1241 (N_1241,In_440,In_2982);
nor U1242 (N_1242,N_511,N_220);
and U1243 (N_1243,In_1829,N_654);
xnor U1244 (N_1244,N_825,In_280);
nor U1245 (N_1245,In_1228,In_1972);
and U1246 (N_1246,N_166,N_673);
and U1247 (N_1247,In_909,In_2841);
or U1248 (N_1248,N_915,In_2933);
or U1249 (N_1249,In_515,N_453);
nor U1250 (N_1250,In_2215,In_2674);
and U1251 (N_1251,In_2833,N_668);
or U1252 (N_1252,N_706,N_805);
or U1253 (N_1253,In_143,N_710);
or U1254 (N_1254,In_223,In_2503);
and U1255 (N_1255,N_408,N_773);
xor U1256 (N_1256,N_809,In_2978);
or U1257 (N_1257,N_501,N_836);
nor U1258 (N_1258,In_1645,N_747);
nand U1259 (N_1259,N_569,N_265);
nand U1260 (N_1260,N_837,In_1305);
and U1261 (N_1261,N_750,N_430);
nand U1262 (N_1262,In_2383,N_367);
nor U1263 (N_1263,N_729,In_2538);
or U1264 (N_1264,In_2164,N_289);
xnor U1265 (N_1265,In_977,In_1176);
and U1266 (N_1266,In_1674,In_2305);
nor U1267 (N_1267,N_178,N_743);
nor U1268 (N_1268,In_1766,In_1378);
and U1269 (N_1269,In_107,In_614);
nand U1270 (N_1270,N_214,In_2883);
or U1271 (N_1271,N_740,In_785);
nand U1272 (N_1272,In_968,In_1654);
and U1273 (N_1273,In_2235,In_1837);
nor U1274 (N_1274,N_473,N_70);
or U1275 (N_1275,N_134,In_926);
or U1276 (N_1276,In_1110,N_897);
and U1277 (N_1277,In_1759,N_927);
and U1278 (N_1278,N_701,In_1823);
xor U1279 (N_1279,In_1272,N_681);
or U1280 (N_1280,In_903,In_1058);
xnor U1281 (N_1281,In_302,In_1942);
nand U1282 (N_1282,In_1950,In_2318);
or U1283 (N_1283,N_84,N_518);
nor U1284 (N_1284,In_2554,N_814);
xnor U1285 (N_1285,N_285,In_1836);
and U1286 (N_1286,N_815,N_649);
or U1287 (N_1287,In_2027,In_1909);
nand U1288 (N_1288,N_57,N_147);
xor U1289 (N_1289,N_764,N_237);
nand U1290 (N_1290,In_429,In_2986);
nor U1291 (N_1291,N_417,In_1256);
nor U1292 (N_1292,In_1560,N_508);
or U1293 (N_1293,N_267,In_2521);
and U1294 (N_1294,N_779,N_477);
nand U1295 (N_1295,N_383,In_1077);
and U1296 (N_1296,N_537,In_2864);
or U1297 (N_1297,In_2455,N_395);
nand U1298 (N_1298,N_761,N_988);
or U1299 (N_1299,In_764,In_1678);
and U1300 (N_1300,In_710,In_2922);
and U1301 (N_1301,N_314,In_2626);
nor U1302 (N_1302,In_1808,N_923);
xnor U1303 (N_1303,In_2594,In_1395);
or U1304 (N_1304,N_309,In_949);
or U1305 (N_1305,In_742,N_95);
xor U1306 (N_1306,N_963,N_81);
nand U1307 (N_1307,In_2352,In_999);
nand U1308 (N_1308,In_1905,In_405);
or U1309 (N_1309,N_235,N_982);
nand U1310 (N_1310,N_958,N_19);
xor U1311 (N_1311,N_822,In_1541);
and U1312 (N_1312,In_601,N_407);
and U1313 (N_1313,In_990,N_748);
nor U1314 (N_1314,In_1291,N_933);
and U1315 (N_1315,N_26,In_546);
nand U1316 (N_1316,N_79,In_2886);
nor U1317 (N_1317,In_2146,N_201);
and U1318 (N_1318,N_145,In_2955);
xnor U1319 (N_1319,N_3,N_411);
nand U1320 (N_1320,N_956,In_196);
or U1321 (N_1321,In_737,N_798);
nand U1322 (N_1322,In_1708,N_901);
nor U1323 (N_1323,N_828,N_276);
or U1324 (N_1324,N_363,N_328);
xor U1325 (N_1325,N_16,N_852);
nor U1326 (N_1326,N_422,N_219);
nand U1327 (N_1327,N_938,In_375);
nor U1328 (N_1328,N_766,In_734);
and U1329 (N_1329,In_2075,N_419);
and U1330 (N_1330,N_862,N_312);
nor U1331 (N_1331,N_576,N_161);
and U1332 (N_1332,N_676,N_256);
and U1333 (N_1333,In_2526,N_76);
xnor U1334 (N_1334,In_1315,In_1417);
and U1335 (N_1335,N_531,In_1914);
nand U1336 (N_1336,N_848,N_817);
nor U1337 (N_1337,In_2485,In_709);
nand U1338 (N_1338,In_1606,N_799);
and U1339 (N_1339,In_1029,N_10);
and U1340 (N_1340,In_1023,N_794);
nand U1341 (N_1341,In_2331,N_847);
and U1342 (N_1342,In_1744,N_741);
or U1343 (N_1343,In_2979,In_2466);
nand U1344 (N_1344,N_465,N_171);
or U1345 (N_1345,N_484,N_638);
nor U1346 (N_1346,N_583,N_959);
and U1347 (N_1347,In_1799,N_947);
or U1348 (N_1348,In_1958,N_451);
or U1349 (N_1349,In_69,In_1433);
xnor U1350 (N_1350,N_776,In_1036);
or U1351 (N_1351,N_672,In_2507);
nor U1352 (N_1352,In_359,N_30);
xnor U1353 (N_1353,N_251,In_2180);
and U1354 (N_1354,N_571,In_2275);
and U1355 (N_1355,N_122,In_2253);
xor U1356 (N_1356,In_998,In_2467);
nand U1357 (N_1357,In_2280,N_751);
nand U1358 (N_1358,N_562,In_2048);
and U1359 (N_1359,In_480,In_729);
or U1360 (N_1360,In_1609,N_77);
xnor U1361 (N_1361,In_1536,N_846);
and U1362 (N_1362,N_12,N_866);
xor U1363 (N_1363,N_519,In_68);
nor U1364 (N_1364,In_1713,In_981);
and U1365 (N_1365,In_2029,In_1753);
and U1366 (N_1366,In_1653,N_239);
nand U1367 (N_1367,In_1610,In_1089);
xnor U1368 (N_1368,In_2396,In_1051);
or U1369 (N_1369,N_431,In_2002);
xor U1370 (N_1370,In_304,N_152);
nor U1371 (N_1371,In_2617,N_43);
or U1372 (N_1372,In_2849,N_281);
nor U1373 (N_1373,N_962,N_559);
and U1374 (N_1374,In_1046,N_173);
nor U1375 (N_1375,N_108,N_415);
and U1376 (N_1376,In_2356,N_479);
or U1377 (N_1377,In_335,N_648);
nand U1378 (N_1378,N_725,N_926);
nor U1379 (N_1379,N_989,N_868);
nand U1380 (N_1380,N_558,N_709);
or U1381 (N_1381,N_42,N_443);
nor U1382 (N_1382,In_220,In_694);
nand U1383 (N_1383,N_552,In_1421);
xnor U1384 (N_1384,In_2781,In_2015);
and U1385 (N_1385,In_2128,N_420);
or U1386 (N_1386,In_2722,In_472);
xnor U1387 (N_1387,N_629,In_1521);
or U1388 (N_1388,N_183,N_807);
nor U1389 (N_1389,N_644,N_772);
nand U1390 (N_1390,N_107,In_978);
nor U1391 (N_1391,In_2291,N_635);
xnor U1392 (N_1392,In_2440,In_1830);
or U1393 (N_1393,In_249,In_1435);
nand U1394 (N_1394,N_687,N_471);
nand U1395 (N_1395,In_2327,N_169);
xnor U1396 (N_1396,In_344,N_384);
or U1397 (N_1397,In_192,In_938);
xnor U1398 (N_1398,N_556,N_573);
xnor U1399 (N_1399,In_2563,In_889);
nand U1400 (N_1400,In_1238,In_2297);
and U1401 (N_1401,In_482,In_1166);
nand U1402 (N_1402,N_247,In_2491);
or U1403 (N_1403,N_299,In_2972);
nor U1404 (N_1404,N_755,N_48);
nand U1405 (N_1405,N_945,N_955);
or U1406 (N_1406,N_831,N_760);
xor U1407 (N_1407,In_2385,In_1088);
xnor U1408 (N_1408,In_510,In_951);
and U1409 (N_1409,N_541,N_647);
nor U1410 (N_1410,N_711,In_2177);
and U1411 (N_1411,In_2171,In_497);
nand U1412 (N_1412,In_1977,N_935);
xnor U1413 (N_1413,N_361,In_1292);
or U1414 (N_1414,In_945,N_921);
or U1415 (N_1415,In_2212,In_838);
or U1416 (N_1416,In_1000,In_574);
nand U1417 (N_1417,In_845,N_733);
or U1418 (N_1418,N_290,N_527);
nand U1419 (N_1419,N_321,N_824);
and U1420 (N_1420,N_719,In_1478);
and U1421 (N_1421,N_450,N_250);
and U1422 (N_1422,N_795,N_896);
or U1423 (N_1423,In_1724,In_1970);
xnor U1424 (N_1424,In_417,In_539);
or U1425 (N_1425,N_426,In_1796);
or U1426 (N_1426,In_2207,N_626);
nor U1427 (N_1427,In_487,In_2322);
nor U1428 (N_1428,In_2360,N_208);
and U1429 (N_1429,N_334,In_2876);
nor U1430 (N_1430,N_609,N_325);
or U1431 (N_1431,In_2487,In_606);
xor U1432 (N_1432,In_266,N_596);
or U1433 (N_1433,In_2925,In_1321);
xor U1434 (N_1434,In_2838,In_2990);
xnor U1435 (N_1435,N_396,N_224);
or U1436 (N_1436,In_1743,In_1398);
nor U1437 (N_1437,N_932,In_2595);
and U1438 (N_1438,In_294,In_1822);
nor U1439 (N_1439,In_1457,In_1346);
or U1440 (N_1440,In_1494,N_243);
or U1441 (N_1441,N_965,N_305);
nand U1442 (N_1442,In_376,N_713);
and U1443 (N_1443,In_371,N_223);
and U1444 (N_1444,In_2304,In_808);
xor U1445 (N_1445,N_914,N_645);
or U1446 (N_1446,In_2091,N_222);
and U1447 (N_1447,N_630,N_390);
or U1448 (N_1448,N_97,In_835);
nand U1449 (N_1449,In_255,N_565);
nor U1450 (N_1450,N_138,N_353);
and U1451 (N_1451,N_184,In_195);
or U1452 (N_1452,N_607,In_2114);
and U1453 (N_1453,In_2716,In_691);
nor U1454 (N_1454,N_61,In_2550);
and U1455 (N_1455,N_440,N_936);
xor U1456 (N_1456,In_1247,N_374);
nand U1457 (N_1457,In_1537,N_308);
nand U1458 (N_1458,In_1588,In_894);
and U1459 (N_1459,In_2123,N_841);
nor U1460 (N_1460,N_516,N_278);
nand U1461 (N_1461,In_672,N_675);
nand U1462 (N_1462,In_2049,N_258);
nor U1463 (N_1463,In_433,N_563);
xnor U1464 (N_1464,In_795,In_1666);
or U1465 (N_1465,In_2154,In_1634);
or U1466 (N_1466,N_372,In_2172);
nand U1467 (N_1467,In_2791,In_2800);
nor U1468 (N_1468,N_187,In_1850);
nand U1469 (N_1469,N_387,In_1363);
xnor U1470 (N_1470,N_929,In_718);
and U1471 (N_1471,N_102,In_1948);
xnor U1472 (N_1472,N_819,In_1188);
or U1473 (N_1473,N_876,N_685);
xor U1474 (N_1474,In_1310,N_434);
nand U1475 (N_1475,In_183,In_517);
and U1476 (N_1476,In_1081,In_2119);
or U1477 (N_1477,In_169,N_641);
and U1478 (N_1478,N_476,In_1872);
xor U1479 (N_1479,N_975,N_274);
xnor U1480 (N_1480,In_2096,In_792);
xnor U1481 (N_1481,In_871,In_2229);
or U1482 (N_1482,In_1302,N_784);
nand U1483 (N_1483,N_549,In_616);
xor U1484 (N_1484,N_326,N_188);
or U1485 (N_1485,N_715,N_744);
and U1486 (N_1486,N_221,In_1737);
and U1487 (N_1487,N_262,N_931);
nor U1488 (N_1488,N_304,N_474);
or U1489 (N_1489,N_628,N_83);
and U1490 (N_1490,In_669,N_632);
or U1491 (N_1491,In_1071,N_925);
or U1492 (N_1492,In_1482,In_13);
nor U1493 (N_1493,In_2357,In_2717);
or U1494 (N_1494,In_1613,In_530);
xnor U1495 (N_1495,In_155,In_2012);
and U1496 (N_1496,N_978,In_2567);
or U1497 (N_1497,In_1490,N_918);
xnor U1498 (N_1498,In_2345,In_1603);
nor U1499 (N_1499,In_2082,N_44);
xor U1500 (N_1500,N_765,In_1112);
and U1501 (N_1501,N_820,In_1891);
nand U1502 (N_1502,N_435,N_920);
nor U1503 (N_1503,In_2949,N_21);
and U1504 (N_1504,N_194,In_2525);
xor U1505 (N_1505,N_332,N_720);
xnor U1506 (N_1506,N_492,N_4);
and U1507 (N_1507,In_256,N_580);
or U1508 (N_1508,In_2217,N_564);
or U1509 (N_1509,In_2809,In_1195);
nand U1510 (N_1510,In_1388,N_899);
and U1511 (N_1511,In_1030,In_1579);
nor U1512 (N_1512,In_442,N_456);
nor U1513 (N_1513,N_268,N_123);
nor U1514 (N_1514,In_870,N_839);
and U1515 (N_1515,In_847,In_1180);
and U1516 (N_1516,N_158,N_661);
nor U1517 (N_1517,N_378,N_211);
nand U1518 (N_1518,N_887,N_879);
nand U1519 (N_1519,In_696,N_924);
nand U1520 (N_1520,N_590,In_2116);
nand U1521 (N_1521,N_62,In_1736);
nor U1522 (N_1522,N_908,In_2731);
xnor U1523 (N_1523,In_326,In_377);
or U1524 (N_1524,N_485,In_1047);
xnor U1525 (N_1525,In_311,N_428);
nand U1526 (N_1526,In_818,In_1179);
xor U1527 (N_1527,In_942,N_977);
and U1528 (N_1528,In_2286,In_2541);
nand U1529 (N_1529,In_463,N_51);
and U1530 (N_1530,In_2768,In_2835);
or U1531 (N_1531,N_283,In_447);
xor U1532 (N_1532,In_1807,N_195);
or U1533 (N_1533,In_740,In_875);
and U1534 (N_1534,In_1042,N_210);
nand U1535 (N_1535,N_875,In_1087);
nand U1536 (N_1536,In_2656,In_2513);
xor U1537 (N_1537,N_103,In_2590);
xor U1538 (N_1538,In_2290,N_246);
and U1539 (N_1539,N_8,N_578);
or U1540 (N_1540,In_1320,N_277);
xor U1541 (N_1541,N_59,In_991);
nand U1542 (N_1542,In_2271,N_746);
or U1543 (N_1543,N_987,N_331);
xnor U1544 (N_1544,N_364,N_911);
xor U1545 (N_1545,In_893,N_515);
nor U1546 (N_1546,N_756,In_2501);
nor U1547 (N_1547,In_1061,In_1992);
nand U1548 (N_1548,In_2081,In_391);
xor U1549 (N_1549,In_1562,In_994);
nor U1550 (N_1550,In_208,In_1117);
nor U1551 (N_1551,In_1921,N_216);
xnor U1552 (N_1552,N_544,In_1525);
xor U1553 (N_1553,In_2387,N_585);
or U1554 (N_1554,N_493,N_736);
or U1555 (N_1555,N_392,N_104);
nand U1556 (N_1556,N_682,N_65);
and U1557 (N_1557,In_1154,In_1391);
and U1558 (N_1558,N_149,In_862);
or U1559 (N_1559,In_1252,In_90);
xnor U1560 (N_1560,N_714,N_553);
nand U1561 (N_1561,N_480,N_366);
nand U1562 (N_1562,In_653,N_560);
or U1563 (N_1563,In_1573,N_253);
xor U1564 (N_1564,In_960,In_10);
and U1565 (N_1565,N_909,In_2840);
xor U1566 (N_1566,N_32,N_853);
or U1567 (N_1567,In_1746,N_738);
xor U1568 (N_1568,N_622,In_1244);
or U1569 (N_1569,In_591,In_543);
xnor U1570 (N_1570,N_793,N_373);
nor U1571 (N_1571,N_574,N_546);
nor U1572 (N_1572,N_347,N_884);
and U1573 (N_1573,N_88,In_1049);
nor U1574 (N_1574,N_448,In_365);
nand U1575 (N_1575,N_466,N_917);
or U1576 (N_1576,N_883,In_106);
and U1577 (N_1577,In_1229,In_1755);
nand U1578 (N_1578,N_310,N_36);
or U1579 (N_1579,In_1258,N_705);
and U1580 (N_1580,N_446,N_494);
or U1581 (N_1581,In_1735,N_664);
and U1582 (N_1582,In_1340,In_770);
or U1583 (N_1583,N_207,N_529);
nor U1584 (N_1584,N_774,N_513);
xor U1585 (N_1585,N_444,In_997);
and U1586 (N_1586,N_114,N_818);
or U1587 (N_1587,In_2638,N_78);
nand U1588 (N_1588,N_790,In_2954);
nor U1589 (N_1589,N_974,N_934);
xor U1590 (N_1590,In_290,In_1317);
nor U1591 (N_1591,N_349,In_2373);
nor U1592 (N_1592,N_606,N_452);
or U1593 (N_1593,N_627,In_2568);
nand U1594 (N_1594,In_379,N_634);
and U1595 (N_1595,N_536,In_2953);
nand U1596 (N_1596,In_366,N_586);
xor U1597 (N_1597,N_812,In_1657);
nor U1598 (N_1598,N_555,N_136);
nor U1599 (N_1599,N_916,N_71);
or U1600 (N_1600,In_1119,N_385);
nand U1601 (N_1601,N_144,In_95);
xor U1602 (N_1602,N_163,N_350);
nor U1603 (N_1603,In_2917,In_2891);
xnor U1604 (N_1604,N_636,N_806);
and U1605 (N_1605,N_716,In_1644);
nand U1606 (N_1606,N_284,In_1871);
and U1607 (N_1607,N_880,In_2210);
or U1608 (N_1608,In_2676,In_1441);
nor U1609 (N_1609,N_757,In_167);
or U1610 (N_1610,N_581,N_154);
nor U1611 (N_1611,N_92,N_489);
and U1612 (N_1612,N_910,N_17);
xor U1613 (N_1613,In_1422,In_678);
nand U1614 (N_1614,In_2967,In_1399);
xnor U1615 (N_1615,N_379,In_2185);
nand U1616 (N_1616,N_252,N_610);
nor U1617 (N_1617,In_411,N_708);
or U1618 (N_1618,In_1241,In_1524);
nand U1619 (N_1619,In_2221,In_2052);
or U1620 (N_1620,N_694,In_2821);
xnor U1621 (N_1621,N_602,N_297);
nand U1622 (N_1622,In_2697,In_2330);
xor U1623 (N_1623,In_1472,In_2031);
xnor U1624 (N_1624,N_994,N_952);
xor U1625 (N_1625,In_1514,In_1949);
nand U1626 (N_1626,In_535,N_591);
nand U1627 (N_1627,In_906,N_509);
nand U1628 (N_1628,N_840,In_313);
xor U1629 (N_1629,N_619,In_276);
or U1630 (N_1630,In_2127,N_118);
nand U1631 (N_1631,In_373,N_339);
nor U1632 (N_1632,N_375,N_679);
nand U1633 (N_1633,N_90,In_2985);
and U1634 (N_1634,N_662,N_674);
nand U1635 (N_1635,N_614,N_745);
nor U1636 (N_1636,In_1437,N_204);
nand U1637 (N_1637,In_247,N_162);
xnor U1638 (N_1638,N_767,In_1986);
nor U1639 (N_1639,N_189,In_1481);
nand U1640 (N_1640,N_376,N_73);
xnor U1641 (N_1641,N_646,N_215);
nor U1642 (N_1642,In_2126,In_1710);
nand U1643 (N_1643,In_1459,N_225);
or U1644 (N_1644,N_306,N_245);
nand U1645 (N_1645,N_587,N_980);
nand U1646 (N_1646,N_651,N_844);
and U1647 (N_1647,N_226,N_1);
xor U1648 (N_1648,In_1869,In_1540);
xnor U1649 (N_1649,In_1968,N_547);
xor U1650 (N_1650,In_1777,In_682);
xor U1651 (N_1651,In_2769,In_658);
xnor U1652 (N_1652,N_728,N_159);
or U1653 (N_1653,In_87,N_991);
xor U1654 (N_1654,In_2706,N_804);
nor U1655 (N_1655,In_899,In_1412);
nor U1656 (N_1656,N_98,In_71);
or U1657 (N_1657,In_1628,In_1067);
and U1658 (N_1658,N_393,N_130);
xnor U1659 (N_1659,In_1882,N_803);
and U1660 (N_1660,N_146,N_96);
nand U1661 (N_1661,N_566,In_286);
xnor U1662 (N_1662,In_1261,In_306);
xor U1663 (N_1663,N_902,N_524);
nor U1664 (N_1664,In_1167,In_418);
nor U1665 (N_1665,N_832,In_100);
or U1666 (N_1666,In_917,In_2619);
nor U1667 (N_1667,N_704,In_2061);
xnor U1668 (N_1668,N_739,N_919);
nor U1669 (N_1669,N_688,N_907);
and U1670 (N_1670,In_2299,N_13);
nor U1671 (N_1671,N_100,In_74);
xor U1672 (N_1672,N_272,In_2668);
or U1673 (N_1673,In_103,N_787);
or U1674 (N_1674,In_1286,In_1480);
or U1675 (N_1675,In_1888,N_343);
nand U1676 (N_1676,In_1510,N_229);
nor U1677 (N_1677,N_603,In_250);
nand U1678 (N_1678,N_66,In_67);
nand U1679 (N_1679,In_743,N_781);
and U1680 (N_1680,N_873,In_2055);
nand U1681 (N_1681,In_2162,In_1138);
and U1682 (N_1682,In_2786,N_775);
or U1683 (N_1683,N_139,N_717);
and U1684 (N_1684,N_595,In_4);
nor U1685 (N_1685,In_372,In_1720);
and U1686 (N_1686,N_157,N_416);
xnor U1687 (N_1687,In_54,N_464);
xnor U1688 (N_1688,N_335,N_47);
nand U1689 (N_1689,In_2125,N_46);
and U1690 (N_1690,In_1867,In_2371);
or U1691 (N_1691,N_882,In_2962);
xor U1692 (N_1692,In_2576,N_979);
xnor U1693 (N_1693,In_2512,N_414);
nand U1694 (N_1694,N_234,N_507);
and U1695 (N_1695,In_1863,In_199);
and U1696 (N_1696,In_1183,N_971);
or U1697 (N_1697,N_906,N_271);
nor U1698 (N_1698,N_270,In_2107);
nand U1699 (N_1699,N_369,In_127);
or U1700 (N_1700,N_984,N_486);
xor U1701 (N_1701,In_2163,N_109);
nor U1702 (N_1702,In_2984,N_718);
xor U1703 (N_1703,In_1411,N_193);
xor U1704 (N_1704,N_117,N_248);
and U1705 (N_1705,N_218,In_1784);
and U1706 (N_1706,N_964,N_330);
and U1707 (N_1707,In_995,In_1492);
nand U1708 (N_1708,N_653,In_1976);
xnor U1709 (N_1709,N_551,In_449);
xor U1710 (N_1710,N_616,In_1985);
nand U1711 (N_1711,N_855,In_2019);
nand U1712 (N_1712,In_2663,In_2044);
xor U1713 (N_1713,N_18,N_835);
and U1714 (N_1714,N_770,N_348);
xor U1715 (N_1715,In_2196,N_763);
nor U1716 (N_1716,In_1194,In_1032);
nand U1717 (N_1717,N_307,N_124);
nand U1718 (N_1718,In_715,In_1552);
nor U1719 (N_1719,N_412,In_1988);
xnor U1720 (N_1720,In_1748,N_973);
nand U1721 (N_1721,In_769,N_33);
and U1722 (N_1722,N_29,N_302);
nand U1723 (N_1723,In_185,In_1920);
xor U1724 (N_1724,In_948,N_260);
or U1725 (N_1725,N_327,N_802);
or U1726 (N_1726,N_782,N_677);
nor U1727 (N_1727,N_151,In_1594);
and U1728 (N_1728,In_2220,N_279);
nand U1729 (N_1729,In_2583,In_2301);
or U1730 (N_1730,In_1498,In_1849);
xor U1731 (N_1731,In_2916,N_663);
nor U1732 (N_1732,In_342,N_941);
xor U1733 (N_1733,N_797,N_594);
or U1734 (N_1734,In_2558,N_637);
nor U1735 (N_1735,In_1347,In_91);
nand U1736 (N_1736,N_116,In_1319);
nand U1737 (N_1737,N_669,N_940);
nor U1738 (N_1738,N_864,N_993);
nand U1739 (N_1739,N_567,N_953);
and U1740 (N_1740,In_1360,N_238);
and U1741 (N_1741,N_930,N_954);
nand U1742 (N_1742,In_2974,N_357);
and U1743 (N_1743,N_449,N_475);
and U1744 (N_1744,N_912,N_22);
nand U1745 (N_1745,In_2807,N_577);
or U1746 (N_1746,In_583,N_657);
and U1747 (N_1747,N_801,N_296);
or U1748 (N_1748,N_698,N_548);
nor U1749 (N_1749,N_721,In_2587);
and U1750 (N_1750,In_1991,N_174);
xor U1751 (N_1751,In_823,N_618);
xor U1752 (N_1752,N_135,N_115);
nor U1753 (N_1753,In_172,In_2895);
or U1754 (N_1754,N_23,N_294);
nand U1755 (N_1755,N_874,N_800);
or U1756 (N_1756,N_181,N_792);
nand U1757 (N_1757,N_523,N_742);
nor U1758 (N_1758,In_1670,In_126);
or U1759 (N_1759,N_754,In_1561);
xnor U1760 (N_1760,N_28,N_113);
or U1761 (N_1761,N_683,In_1604);
xor U1762 (N_1762,N_202,N_410);
or U1763 (N_1763,N_849,In_1158);
nor U1764 (N_1764,In_841,In_2473);
and U1765 (N_1765,N_457,In_1475);
and U1766 (N_1766,In_752,N_838);
xor U1767 (N_1767,In_1955,In_2236);
nor U1768 (N_1768,In_693,In_1142);
and U1769 (N_1769,In_2454,In_587);
nor U1770 (N_1770,N_74,N_345);
nand U1771 (N_1771,N_700,In_1300);
and U1772 (N_1772,In_1516,N_752);
or U1773 (N_1773,N_402,N_240);
nor U1774 (N_1774,N_39,In_193);
nand U1775 (N_1775,In_1027,In_534);
or U1776 (N_1776,N_950,N_316);
nand U1777 (N_1777,In_964,N_200);
nor U1778 (N_1778,N_881,N_111);
xor U1779 (N_1779,In_428,N_292);
nor U1780 (N_1780,In_713,In_844);
nand U1781 (N_1781,N_487,In_2613);
nand U1782 (N_1782,N_723,N_900);
nand U1783 (N_1783,N_472,In_438);
or U1784 (N_1784,In_231,N_425);
xnor U1785 (N_1785,N_554,N_903);
or U1786 (N_1786,N_811,N_156);
nor U1787 (N_1787,In_1405,In_212);
nor U1788 (N_1788,N_231,In_892);
xnor U1789 (N_1789,In_1690,N_759);
nor U1790 (N_1790,N_499,In_775);
and U1791 (N_1791,N_142,N_324);
xor U1792 (N_1792,N_888,In_1912);
and U1793 (N_1793,In_356,N_7);
and U1794 (N_1794,In_2806,In_1567);
nand U1795 (N_1795,N_597,N_894);
or U1796 (N_1796,In_2940,N_512);
and U1797 (N_1797,N_244,In_630);
nor U1798 (N_1798,In_1235,In_2021);
nand U1799 (N_1799,N_611,In_1782);
nand U1800 (N_1800,N_398,In_2423);
and U1801 (N_1801,In_2093,N_301);
nand U1802 (N_1802,N_236,In_2034);
nand U1803 (N_1803,In_2994,In_504);
and U1804 (N_1804,In_588,N_34);
xor U1805 (N_1805,N_365,In_1012);
xor U1806 (N_1806,N_780,In_1626);
xnor U1807 (N_1807,In_2284,N_67);
nand U1808 (N_1808,N_320,N_160);
nand U1809 (N_1809,N_834,In_485);
nor U1810 (N_1810,In_2779,In_1285);
and U1811 (N_1811,In_1037,In_751);
xor U1812 (N_1812,In_2004,In_1691);
xnor U1813 (N_1813,In_2033,In_528);
nand U1814 (N_1814,N_788,N_191);
xor U1815 (N_1815,In_98,In_2898);
or U1816 (N_1816,In_1384,N_404);
nor U1817 (N_1817,In_1212,In_632);
nor U1818 (N_1818,N_14,N_850);
nor U1819 (N_1819,N_133,In_763);
or U1820 (N_1820,In_928,In_2490);
or U1821 (N_1821,In_2369,In_1133);
xor U1822 (N_1822,In_2178,In_2719);
nand U1823 (N_1823,N_829,In_699);
and U1824 (N_1824,In_498,In_1308);
nand U1825 (N_1825,In_1930,N_454);
and U1826 (N_1826,In_2845,In_932);
xor U1827 (N_1827,In_2899,N_27);
and U1828 (N_1828,N_397,N_129);
xor U1829 (N_1829,N_526,In_1506);
nand U1830 (N_1830,In_506,In_2496);
nand U1831 (N_1831,N_490,N_342);
or U1832 (N_1832,In_1508,N_605);
and U1833 (N_1833,In_1341,N_360);
nor U1834 (N_1834,In_2830,In_252);
nor U1835 (N_1835,N_119,In_2843);
nor U1836 (N_1836,N_371,In_2228);
or U1837 (N_1837,N_703,N_427);
and U1838 (N_1838,In_451,In_96);
nor U1839 (N_1839,N_601,In_1683);
or U1840 (N_1840,N_778,N_80);
nand U1841 (N_1841,N_172,N_168);
nor U1842 (N_1842,N_889,N_180);
and U1843 (N_1843,In_2866,In_2644);
xnor U1844 (N_1844,N_695,In_1551);
or U1845 (N_1845,In_265,N_400);
xor U1846 (N_1846,N_120,In_2358);
and U1847 (N_1847,In_644,N_970);
nor U1848 (N_1848,N_789,In_1041);
nor U1849 (N_1849,In_2858,N_588);
or U1850 (N_1850,N_998,N_783);
or U1851 (N_1851,N_656,In_2350);
and U1852 (N_1852,N_535,In_2289);
nand U1853 (N_1853,N_75,N_101);
nand U1854 (N_1854,N_707,In_1339);
nor U1855 (N_1855,In_1878,N_727);
nand U1856 (N_1856,In_1883,N_735);
or U1857 (N_1857,N_205,N_336);
or U1858 (N_1858,In_1313,In_834);
or U1859 (N_1859,N_56,N_459);
nand U1860 (N_1860,In_1639,N_275);
xor U1861 (N_1861,N_510,N_538);
xor U1862 (N_1862,N_528,In_1875);
nor U1863 (N_1863,N_89,N_854);
xor U1864 (N_1864,In_1693,In_145);
nand U1865 (N_1865,In_444,N_185);
xor U1866 (N_1866,In_1024,In_725);
xor U1867 (N_1867,In_1845,In_2462);
and U1868 (N_1868,In_585,N_391);
and U1869 (N_1869,In_1586,In_1434);
and U1870 (N_1870,In_1275,In_471);
and U1871 (N_1871,In_2139,In_2069);
and U1872 (N_1872,In_2338,N_584);
xnor U1873 (N_1873,N_697,In_1831);
nand U1874 (N_1874,In_1578,N_93);
or U1875 (N_1875,In_547,N_266);
or U1876 (N_1876,N_257,In_1418);
xor U1877 (N_1877,N_94,In_560);
nand U1878 (N_1878,N_830,N_341);
xor U1879 (N_1879,N_730,N_0);
or U1880 (N_1880,In_2529,N_405);
and U1881 (N_1881,N_31,In_1979);
xor U1882 (N_1882,N_845,N_992);
and U1883 (N_1883,In_520,N_599);
or U1884 (N_1884,In_1287,In_521);
nand U1885 (N_1885,In_2254,In_1557);
xnor U1886 (N_1886,N_6,In_2540);
or U1887 (N_1887,N_11,In_940);
and U1888 (N_1888,N_521,In_523);
nand U1889 (N_1889,In_913,In_2310);
or U1890 (N_1890,In_2739,In_2701);
nand U1891 (N_1891,In_1267,N_858);
and U1892 (N_1892,N_944,In_594);
or U1893 (N_1893,N_539,N_228);
and U1894 (N_1894,In_386,In_259);
and U1895 (N_1895,In_1173,In_724);
nand U1896 (N_1896,N_315,In_1899);
nor U1897 (N_1897,N_665,N_298);
nor U1898 (N_1898,N_38,In_1306);
xor U1899 (N_1899,N_904,N_808);
xnor U1900 (N_1900,N_380,In_1839);
nand U1901 (N_1901,In_2057,N_893);
nand U1902 (N_1902,N_734,In_27);
and U1903 (N_1903,In_676,In_439);
nand U1904 (N_1904,N_786,In_2218);
xor U1905 (N_1905,N_785,In_661);
or U1906 (N_1906,In_890,In_2336);
or U1907 (N_1907,N_351,N_981);
xnor U1908 (N_1908,In_343,In_1444);
and U1909 (N_1909,N_624,In_1381);
xor U1910 (N_1910,In_2867,N_354);
or U1911 (N_1911,N_254,N_702);
or U1912 (N_1912,In_873,N_176);
nand U1913 (N_1913,N_842,In_2020);
and U1914 (N_1914,N_155,In_254);
xor U1915 (N_1915,N_192,In_347);
and U1916 (N_1916,In_1941,N_851);
xor U1917 (N_1917,N_856,N_520);
nor U1918 (N_1918,In_1581,N_209);
or U1919 (N_1919,In_2814,N_401);
or U1920 (N_1920,In_1568,In_23);
or U1921 (N_1921,N_568,N_461);
or U1922 (N_1922,N_358,In_633);
xor U1923 (N_1923,N_233,In_1393);
xnor U1924 (N_1924,In_2265,In_1008);
nor U1925 (N_1925,In_314,N_217);
or U1926 (N_1926,In_961,N_732);
or U1927 (N_1927,N_317,In_1035);
xnor U1928 (N_1928,In_2790,In_2001);
and U1929 (N_1929,N_381,N_287);
nand U1930 (N_1930,N_497,In_2068);
or U1931 (N_1931,N_394,N_843);
nand U1932 (N_1932,In_1874,In_370);
and U1933 (N_1933,N_323,In_3);
and U1934 (N_1934,N_692,N_640);
and U1935 (N_1935,N_503,N_865);
nor U1936 (N_1936,In_207,N_621);
nand U1937 (N_1937,N_615,N_561);
nor U1938 (N_1938,In_1960,N_368);
nand U1939 (N_1939,In_1608,N_196);
or U1940 (N_1940,N_424,N_550);
nand U1941 (N_1941,In_1416,N_943);
nor U1942 (N_1942,N_625,In_1002);
nor U1943 (N_1943,In_45,In_1485);
nand U1944 (N_1944,In_1447,In_2735);
and U1945 (N_1945,In_1864,In_2341);
xor U1946 (N_1946,In_2799,In_30);
xor U1947 (N_1947,In_2366,In_1019);
nor U1948 (N_1948,In_2230,N_949);
or U1949 (N_1949,N_996,N_995);
or U1950 (N_1950,In_1947,In_1337);
and U1951 (N_1951,In_788,N_737);
xor U1952 (N_1952,N_928,N_388);
xor U1953 (N_1953,In_2281,In_916);
xor U1954 (N_1954,In_558,In_297);
or U1955 (N_1955,In_2225,N_823);
nand U1956 (N_1956,In_2574,N_463);
nand U1957 (N_1957,In_2113,N_288);
and U1958 (N_1958,In_2398,N_660);
and U1959 (N_1959,N_686,N_175);
nor U1960 (N_1960,N_106,N_273);
nor U1961 (N_1961,N_898,N_421);
nand U1962 (N_1962,N_608,N_796);
nor U1963 (N_1963,N_895,In_2319);
xor U1964 (N_1964,N_498,In_1257);
and U1965 (N_1965,In_1577,N_413);
nand U1966 (N_1966,N_9,N_504);
xor U1967 (N_1967,N_589,In_1734);
or U1968 (N_1968,In_2882,In_274);
or U1969 (N_1969,N_872,N_41);
xnor U1970 (N_1970,In_2709,In_454);
and U1971 (N_1971,In_1587,In_101);
or U1972 (N_1972,In_2446,N_132);
xor U1973 (N_1973,In_1311,In_2190);
xnor U1974 (N_1974,N_985,N_5);
nand U1975 (N_1975,N_821,In_89);
nor U1976 (N_1976,N_54,In_804);
xor U1977 (N_1977,In_327,N_813);
and U1978 (N_1978,In_1116,In_2317);
nor U1979 (N_1979,In_1714,N_322);
and U1980 (N_1980,In_363,In_394);
nor U1981 (N_1981,N_458,N_303);
xnor U1982 (N_1982,In_590,N_64);
or U1983 (N_1983,In_1898,In_898);
xor U1984 (N_1984,In_2308,N_592);
or U1985 (N_1985,In_1523,N_948);
or U1986 (N_1986,In_541,In_2258);
nor U1987 (N_1987,In_215,In_2670);
nor U1988 (N_1988,In_2042,In_58);
or U1989 (N_1989,N_386,In_1130);
nand U1990 (N_1990,N_263,N_437);
nor U1991 (N_1991,In_562,In_1309);
nand U1992 (N_1992,N_905,N_445);
and U1993 (N_1993,In_1854,N_232);
nor U1994 (N_1994,N_242,N_186);
xor U1995 (N_1995,N_972,In_846);
and U1996 (N_1996,In_139,In_1001);
or U1997 (N_1997,In_2173,In_1038);
nor U1998 (N_1998,N_91,N_442);
nand U1999 (N_1999,N_690,In_1147);
nor U2000 (N_2000,N_1647,N_1104);
or U2001 (N_2001,N_1106,N_1037);
or U2002 (N_2002,N_1930,N_1812);
xor U2003 (N_2003,N_1762,N_1826);
nand U2004 (N_2004,N_1565,N_1452);
xor U2005 (N_2005,N_1983,N_1063);
or U2006 (N_2006,N_1966,N_1373);
nor U2007 (N_2007,N_1878,N_1094);
and U2008 (N_2008,N_1308,N_1659);
and U2009 (N_2009,N_1204,N_1665);
nor U2010 (N_2010,N_1376,N_1239);
or U2011 (N_2011,N_1331,N_1099);
or U2012 (N_2012,N_1107,N_1971);
xor U2013 (N_2013,N_1705,N_1864);
nor U2014 (N_2014,N_1747,N_1183);
or U2015 (N_2015,N_1334,N_1506);
and U2016 (N_2016,N_1509,N_1141);
xnor U2017 (N_2017,N_1843,N_1207);
xnor U2018 (N_2018,N_1296,N_1065);
nand U2019 (N_2019,N_1952,N_1816);
and U2020 (N_2020,N_1160,N_1608);
xor U2021 (N_2021,N_1850,N_1682);
nor U2022 (N_2022,N_1643,N_1466);
or U2023 (N_2023,N_1152,N_1679);
and U2024 (N_2024,N_1410,N_1751);
and U2025 (N_2025,N_1711,N_1748);
nor U2026 (N_2026,N_1162,N_1198);
xor U2027 (N_2027,N_1592,N_1793);
nor U2028 (N_2028,N_1265,N_1990);
or U2029 (N_2029,N_1332,N_1633);
xor U2030 (N_2030,N_1859,N_1758);
xnor U2031 (N_2031,N_1272,N_1144);
nor U2032 (N_2032,N_1507,N_1440);
nor U2033 (N_2033,N_1785,N_1362);
or U2034 (N_2034,N_1087,N_1210);
nand U2035 (N_2035,N_1354,N_1525);
nor U2036 (N_2036,N_1310,N_1380);
or U2037 (N_2037,N_1432,N_1753);
or U2038 (N_2038,N_1025,N_1865);
or U2039 (N_2039,N_1283,N_1177);
nor U2040 (N_2040,N_1417,N_1825);
nand U2041 (N_2041,N_1042,N_1407);
and U2042 (N_2042,N_1480,N_1512);
or U2043 (N_2043,N_1021,N_1866);
and U2044 (N_2044,N_1384,N_1600);
or U2045 (N_2045,N_1858,N_1796);
xor U2046 (N_2046,N_1357,N_1847);
nand U2047 (N_2047,N_1472,N_1009);
nor U2048 (N_2048,N_1536,N_1423);
nor U2049 (N_2049,N_1015,N_1074);
nor U2050 (N_2050,N_1415,N_1095);
and U2051 (N_2051,N_1911,N_1539);
nor U2052 (N_2052,N_1285,N_1403);
xnor U2053 (N_2053,N_1834,N_1400);
nand U2054 (N_2054,N_1733,N_1564);
nand U2055 (N_2055,N_1427,N_1098);
xor U2056 (N_2056,N_1398,N_1041);
and U2057 (N_2057,N_1253,N_1542);
nor U2058 (N_2058,N_1430,N_1982);
or U2059 (N_2059,N_1991,N_1620);
nand U2060 (N_2060,N_1302,N_1093);
or U2061 (N_2061,N_1245,N_1563);
or U2062 (N_2062,N_1612,N_1721);
or U2063 (N_2063,N_1264,N_1585);
nor U2064 (N_2064,N_1809,N_1129);
and U2065 (N_2065,N_1562,N_1914);
or U2066 (N_2066,N_1717,N_1341);
or U2067 (N_2067,N_1737,N_1677);
nand U2068 (N_2068,N_1327,N_1981);
and U2069 (N_2069,N_1589,N_1352);
or U2070 (N_2070,N_1372,N_1220);
nor U2071 (N_2071,N_1580,N_1568);
or U2072 (N_2072,N_1856,N_1353);
or U2073 (N_2073,N_1078,N_1441);
nor U2074 (N_2074,N_1374,N_1576);
nand U2075 (N_2075,N_1479,N_1201);
nor U2076 (N_2076,N_1181,N_1393);
nor U2077 (N_2077,N_1953,N_1544);
and U2078 (N_2078,N_1840,N_1686);
nand U2079 (N_2079,N_1942,N_1891);
xnor U2080 (N_2080,N_1744,N_1892);
nor U2081 (N_2081,N_1028,N_1454);
nand U2082 (N_2082,N_1014,N_1829);
and U2083 (N_2083,N_1926,N_1326);
or U2084 (N_2084,N_1121,N_1456);
xnor U2085 (N_2085,N_1727,N_1408);
nor U2086 (N_2086,N_1993,N_1382);
nor U2087 (N_2087,N_1111,N_1738);
nor U2088 (N_2088,N_1746,N_1928);
xnor U2089 (N_2089,N_1668,N_1969);
and U2090 (N_2090,N_1084,N_1126);
nor U2091 (N_2091,N_1795,N_1309);
or U2092 (N_2092,N_1208,N_1103);
nor U2093 (N_2093,N_1279,N_1157);
nor U2094 (N_2094,N_1205,N_1061);
or U2095 (N_2095,N_1258,N_1560);
nand U2096 (N_2096,N_1096,N_1236);
or U2097 (N_2097,N_1473,N_1321);
and U2098 (N_2098,N_1378,N_1765);
nand U2099 (N_2099,N_1277,N_1559);
nor U2100 (N_2100,N_1940,N_1798);
nand U2101 (N_2101,N_1588,N_1889);
nor U2102 (N_2102,N_1617,N_1616);
nand U2103 (N_2103,N_1995,N_1792);
and U2104 (N_2104,N_1537,N_1081);
xnor U2105 (N_2105,N_1155,N_1964);
nor U2106 (N_2106,N_1805,N_1092);
and U2107 (N_2107,N_1857,N_1573);
nand U2108 (N_2108,N_1045,N_1819);
and U2109 (N_2109,N_1048,N_1924);
nor U2110 (N_2110,N_1178,N_1505);
nand U2111 (N_2111,N_1956,N_1476);
or U2112 (N_2112,N_1718,N_1218);
or U2113 (N_2113,N_1271,N_1574);
or U2114 (N_2114,N_1289,N_1607);
xor U2115 (N_2115,N_1534,N_1246);
and U2116 (N_2116,N_1681,N_1128);
or U2117 (N_2117,N_1312,N_1197);
xor U2118 (N_2118,N_1471,N_1123);
xor U2119 (N_2119,N_1292,N_1330);
nand U2120 (N_2120,N_1324,N_1269);
nand U2121 (N_2121,N_1381,N_1527);
nor U2122 (N_2122,N_1058,N_1595);
nor U2123 (N_2123,N_1869,N_1791);
or U2124 (N_2124,N_1596,N_1338);
nor U2125 (N_2125,N_1550,N_1010);
xor U2126 (N_2126,N_1775,N_1194);
and U2127 (N_2127,N_1119,N_1115);
nand U2128 (N_2128,N_1019,N_1364);
nand U2129 (N_2129,N_1555,N_1346);
or U2130 (N_2130,N_1614,N_1667);
or U2131 (N_2131,N_1174,N_1363);
xnor U2132 (N_2132,N_1091,N_1619);
nand U2133 (N_2133,N_1200,N_1979);
and U2134 (N_2134,N_1250,N_1469);
or U2135 (N_2135,N_1672,N_1919);
xor U2136 (N_2136,N_1811,N_1033);
nand U2137 (N_2137,N_1286,N_1556);
and U2138 (N_2138,N_1514,N_1824);
nand U2139 (N_2139,N_1779,N_1149);
or U2140 (N_2140,N_1913,N_1146);
or U2141 (N_2141,N_1377,N_1077);
xnor U2142 (N_2142,N_1387,N_1728);
xnor U2143 (N_2143,N_1951,N_1941);
nand U2144 (N_2144,N_1526,N_1613);
nor U2145 (N_2145,N_1599,N_1117);
or U2146 (N_2146,N_1970,N_1611);
and U2147 (N_2147,N_1029,N_1267);
and U2148 (N_2148,N_1213,N_1138);
xor U2149 (N_2149,N_1158,N_1333);
nor U2150 (N_2150,N_1597,N_1909);
nor U2151 (N_2151,N_1217,N_1317);
nand U2152 (N_2152,N_1495,N_1233);
xor U2153 (N_2153,N_1939,N_1402);
nand U2154 (N_2154,N_1242,N_1523);
nand U2155 (N_2155,N_1630,N_1713);
nor U2156 (N_2156,N_1463,N_1957);
xnor U2157 (N_2157,N_1692,N_1335);
nor U2158 (N_2158,N_1262,N_1827);
nor U2159 (N_2159,N_1499,N_1591);
nand U2160 (N_2160,N_1813,N_1579);
and U2161 (N_2161,N_1229,N_1276);
nand U2162 (N_2162,N_1492,N_1488);
xor U2163 (N_2163,N_1192,N_1846);
or U2164 (N_2164,N_1967,N_1422);
or U2165 (N_2165,N_1431,N_1936);
and U2166 (N_2166,N_1294,N_1777);
xnor U2167 (N_2167,N_1419,N_1797);
nand U2168 (N_2168,N_1132,N_1114);
or U2169 (N_2169,N_1026,N_1343);
nor U2170 (N_2170,N_1671,N_1424);
nor U2171 (N_2171,N_1848,N_1604);
and U2172 (N_2172,N_1949,N_1266);
nand U2173 (N_2173,N_1501,N_1112);
nand U2174 (N_2174,N_1133,N_1071);
or U2175 (N_2175,N_1822,N_1036);
or U2176 (N_2176,N_1828,N_1224);
xor U2177 (N_2177,N_1358,N_1912);
and U2178 (N_2178,N_1085,N_1195);
xnor U2179 (N_2179,N_1586,N_1366);
nor U2180 (N_2180,N_1237,N_1690);
nor U2181 (N_2181,N_1487,N_1925);
nor U2182 (N_2182,N_1089,N_1004);
or U2183 (N_2183,N_1278,N_1223);
nand U2184 (N_2184,N_1803,N_1216);
and U2185 (N_2185,N_1170,N_1470);
nor U2186 (N_2186,N_1039,N_1626);
nor U2187 (N_2187,N_1287,N_1761);
nor U2188 (N_2188,N_1247,N_1165);
nand U2189 (N_2189,N_1528,N_1888);
nand U2190 (N_2190,N_1994,N_1388);
nand U2191 (N_2191,N_1898,N_1068);
and U2192 (N_2192,N_1518,N_1072);
nand U2193 (N_2193,N_1464,N_1038);
xnor U2194 (N_2194,N_1052,N_1179);
or U2195 (N_2195,N_1437,N_1306);
nor U2196 (N_2196,N_1290,N_1548);
or U2197 (N_2197,N_1734,N_1116);
nor U2198 (N_2198,N_1769,N_1807);
xor U2199 (N_2199,N_1188,N_1663);
or U2200 (N_2200,N_1154,N_1273);
nand U2201 (N_2201,N_1571,N_1902);
nand U2202 (N_2202,N_1557,N_1947);
nor U2203 (N_2203,N_1907,N_1999);
nand U2204 (N_2204,N_1203,N_1259);
and U2205 (N_2205,N_1148,N_1315);
nand U2206 (N_2206,N_1897,N_1496);
xor U2207 (N_2207,N_1301,N_1590);
or U2208 (N_2208,N_1593,N_1745);
or U2209 (N_2209,N_1685,N_1102);
or U2210 (N_2210,N_1067,N_1356);
nand U2211 (N_2211,N_1521,N_1135);
xnor U2212 (N_2212,N_1655,N_1875);
and U2213 (N_2213,N_1639,N_1678);
nand U2214 (N_2214,N_1455,N_1405);
xnor U2215 (N_2215,N_1768,N_1411);
xnor U2216 (N_2216,N_1531,N_1238);
xnor U2217 (N_2217,N_1989,N_1386);
and U2218 (N_2218,N_1013,N_1212);
and U2219 (N_2219,N_1069,N_1905);
xor U2220 (N_2220,N_1664,N_1908);
nor U2221 (N_2221,N_1697,N_1871);
and U2222 (N_2222,N_1752,N_1529);
nor U2223 (N_2223,N_1687,N_1484);
nor U2224 (N_2224,N_1513,N_1642);
nand U2225 (N_2225,N_1541,N_1756);
nand U2226 (N_2226,N_1142,N_1426);
nor U2227 (N_2227,N_1156,N_1644);
or U2228 (N_2228,N_1396,N_1901);
nor U2229 (N_2229,N_1347,N_1182);
or U2230 (N_2230,N_1307,N_1749);
and U2231 (N_2231,N_1771,N_1360);
nand U2232 (N_2232,N_1992,N_1836);
and U2233 (N_2233,N_1050,N_1683);
or U2234 (N_2234,N_1319,N_1927);
or U2235 (N_2235,N_1741,N_1448);
nand U2236 (N_2236,N_1553,N_1399);
or U2237 (N_2237,N_1566,N_1732);
or U2238 (N_2238,N_1802,N_1654);
nand U2239 (N_2239,N_1657,N_1652);
and U2240 (N_2240,N_1660,N_1249);
nand U2241 (N_2241,N_1783,N_1497);
or U2242 (N_2242,N_1511,N_1710);
nand U2243 (N_2243,N_1046,N_1412);
nor U2244 (N_2244,N_1638,N_1552);
xnor U2245 (N_2245,N_1228,N_1578);
or U2246 (N_2246,N_1298,N_1351);
or U2247 (N_2247,N_1180,N_1975);
or U2248 (N_2248,N_1674,N_1478);
nand U2249 (N_2249,N_1945,N_1770);
xor U2250 (N_2250,N_1572,N_1445);
xor U2251 (N_2251,N_1887,N_1450);
xnor U2252 (N_2252,N_1823,N_1120);
nor U2253 (N_2253,N_1972,N_1057);
nand U2254 (N_2254,N_1766,N_1680);
nor U2255 (N_2255,N_1708,N_1371);
and U2256 (N_2256,N_1461,N_1449);
nand U2257 (N_2257,N_1299,N_1845);
nand U2258 (N_2258,N_1903,N_1706);
and U2259 (N_2259,N_1375,N_1997);
or U2260 (N_2260,N_1695,N_1561);
and U2261 (N_2261,N_1577,N_1842);
xor U2262 (N_2262,N_1881,N_1263);
nand U2263 (N_2263,N_1524,N_1109);
nor U2264 (N_2264,N_1694,N_1754);
nand U2265 (N_2265,N_1244,N_1870);
and U2266 (N_2266,N_1090,N_1428);
xnor U2267 (N_2267,N_1776,N_1284);
or U2268 (N_2268,N_1429,N_1457);
nand U2269 (N_2269,N_1214,N_1206);
and U2270 (N_2270,N_1367,N_1520);
nand U2271 (N_2271,N_1621,N_1786);
xor U2272 (N_2272,N_1545,N_1606);
or U2273 (N_2273,N_1814,N_1305);
xor U2274 (N_2274,N_1917,N_1641);
xor U2275 (N_2275,N_1465,N_1804);
or U2276 (N_2276,N_1627,N_1973);
nor U2277 (N_2277,N_1635,N_1549);
xor U2278 (N_2278,N_1603,N_1027);
xor U2279 (N_2279,N_1689,N_1159);
nor U2280 (N_2280,N_1369,N_1199);
xor U2281 (N_2281,N_1086,N_1533);
or U2282 (N_2282,N_1515,N_1872);
nand U2283 (N_2283,N_1699,N_1838);
and U2284 (N_2284,N_1631,N_1637);
nor U2285 (N_2285,N_1740,N_1118);
and U2286 (N_2286,N_1110,N_1349);
nand U2287 (N_2287,N_1304,N_1161);
nand U2288 (N_2288,N_1772,N_1462);
or U2289 (N_2289,N_1730,N_1782);
or U2290 (N_2290,N_1731,N_1551);
nand U2291 (N_2291,N_1137,N_1409);
and U2292 (N_2292,N_1918,N_1879);
xor U2293 (N_2293,N_1017,N_1934);
nand U2294 (N_2294,N_1849,N_1168);
or U2295 (N_2295,N_1368,N_1629);
and U2296 (N_2296,N_1893,N_1007);
nand U2297 (N_2297,N_1517,N_1191);
and U2298 (N_2298,N_1764,N_1535);
or U2299 (N_2299,N_1379,N_1288);
or U2300 (N_2300,N_1890,N_1609);
nor U2301 (N_2301,N_1024,N_1774);
nand U2302 (N_2302,N_1260,N_1211);
or U2303 (N_2303,N_1724,N_1504);
and U2304 (N_2304,N_1185,N_1988);
nand U2305 (N_2305,N_1035,N_1002);
xnor U2306 (N_2306,N_1006,N_1906);
nand U2307 (N_2307,N_1575,N_1459);
nand U2308 (N_2308,N_1817,N_1538);
xor U2309 (N_2309,N_1040,N_1801);
and U2310 (N_2310,N_1325,N_1636);
xnor U2311 (N_2311,N_1662,N_1789);
nor U2312 (N_2312,N_1446,N_1406);
or U2313 (N_2313,N_1581,N_1831);
or U2314 (N_2314,N_1060,N_1145);
xnor U2315 (N_2315,N_1532,N_1187);
nand U2316 (N_2316,N_1498,N_1799);
nand U2317 (N_2317,N_1383,N_1190);
xnor U2318 (N_2318,N_1780,N_1340);
nand U2319 (N_2319,N_1656,N_1915);
xor U2320 (N_2320,N_1500,N_1011);
or U2321 (N_2321,N_1618,N_1108);
nor U2322 (N_2322,N_1083,N_1790);
xor U2323 (N_2323,N_1297,N_1202);
xnor U2324 (N_2324,N_1980,N_1894);
nor U2325 (N_2325,N_1696,N_1337);
nand U2326 (N_2326,N_1863,N_1163);
or U2327 (N_2327,N_1714,N_1583);
xor U2328 (N_2328,N_1698,N_1008);
nand U2329 (N_2329,N_1522,N_1645);
nor U2330 (N_2330,N_1853,N_1916);
nand U2331 (N_2331,N_1056,N_1003);
or U2332 (N_2332,N_1291,N_1510);
xor U2333 (N_2333,N_1231,N_1131);
xnor U2334 (N_2334,N_1508,N_1054);
xor U2335 (N_2335,N_1490,N_1808);
xnor U2336 (N_2336,N_1059,N_1391);
nand U2337 (N_2337,N_1725,N_1830);
nand U2338 (N_2338,N_1723,N_1987);
or U2339 (N_2339,N_1164,N_1860);
nand U2340 (N_2340,N_1361,N_1359);
nor U2341 (N_2341,N_1821,N_1895);
nand U2342 (N_2342,N_1904,N_1719);
nand U2343 (N_2343,N_1787,N_1222);
and U2344 (N_2344,N_1547,N_1018);
xor U2345 (N_2345,N_1255,N_1675);
and U2346 (N_2346,N_1064,N_1955);
nor U2347 (N_2347,N_1855,N_1920);
and U2348 (N_2348,N_1034,N_1491);
nor U2349 (N_2349,N_1311,N_1420);
and U2350 (N_2350,N_1839,N_1666);
xor U2351 (N_2351,N_1241,N_1702);
nor U2352 (N_2352,N_1570,N_1569);
or U2353 (N_2353,N_1234,N_1493);
xnor U2354 (N_2354,N_1720,N_1582);
nand U2355 (N_2355,N_1257,N_1806);
xor U2356 (N_2356,N_1862,N_1055);
or U2357 (N_2357,N_1075,N_1240);
nor U2358 (N_2358,N_1605,N_1700);
xor U2359 (N_2359,N_1944,N_1482);
nor U2360 (N_2360,N_1062,N_1225);
nor U2361 (N_2361,N_1467,N_1530);
nor U2362 (N_2362,N_1594,N_1800);
nand U2363 (N_2363,N_1416,N_1778);
nand U2364 (N_2364,N_1043,N_1100);
and U2365 (N_2365,N_1113,N_1709);
and U2366 (N_2366,N_1598,N_1935);
nand U2367 (N_2367,N_1243,N_1844);
nor U2368 (N_2368,N_1625,N_1961);
nand U2369 (N_2369,N_1610,N_1623);
and U2370 (N_2370,N_1884,N_1820);
or U2371 (N_2371,N_1044,N_1477);
nor U2372 (N_2372,N_1397,N_1189);
and U2373 (N_2373,N_1166,N_1837);
and U2374 (N_2374,N_1923,N_1485);
or U2375 (N_2375,N_1968,N_1143);
xnor U2376 (N_2376,N_1221,N_1948);
or U2377 (N_2377,N_1784,N_1707);
xnor U2378 (N_2378,N_1339,N_1835);
or U2379 (N_2379,N_1877,N_1962);
and U2380 (N_2380,N_1395,N_1996);
or U2381 (N_2381,N_1688,N_1632);
or U2382 (N_2382,N_1474,N_1701);
or U2383 (N_2383,N_1703,N_1984);
xor U2384 (N_2384,N_1601,N_1818);
and U2385 (N_2385,N_1886,N_1757);
or U2386 (N_2386,N_1932,N_1281);
or U2387 (N_2387,N_1175,N_1938);
and U2388 (N_2388,N_1634,N_1053);
and U2389 (N_2389,N_1885,N_1444);
or U2390 (N_2390,N_1503,N_1676);
and U2391 (N_2391,N_1615,N_1350);
nand U2392 (N_2392,N_1646,N_1540);
nand U2393 (N_2393,N_1439,N_1254);
xnor U2394 (N_2394,N_1303,N_1554);
xnor U2395 (N_2395,N_1451,N_1767);
xor U2396 (N_2396,N_1959,N_1314);
nand U2397 (N_2397,N_1841,N_1481);
nor U2398 (N_2398,N_1355,N_1453);
xnor U2399 (N_2399,N_1082,N_1810);
nand U2400 (N_2400,N_1150,N_1963);
or U2401 (N_2401,N_1097,N_1759);
nand U2402 (N_2402,N_1125,N_1729);
nand U2403 (N_2403,N_1370,N_1316);
xnor U2404 (N_2404,N_1670,N_1122);
and U2405 (N_2405,N_1425,N_1684);
xor U2406 (N_2406,N_1587,N_1788);
xnor U2407 (N_2407,N_1256,N_1105);
nor U2408 (N_2408,N_1421,N_1235);
nand U2409 (N_2409,N_1280,N_1519);
xor U2410 (N_2410,N_1943,N_1976);
nand U2411 (N_2411,N_1910,N_1602);
or U2412 (N_2412,N_1502,N_1342);
nor U2413 (N_2413,N_1950,N_1344);
or U2414 (N_2414,N_1650,N_1124);
nor U2415 (N_2415,N_1404,N_1193);
xnor U2416 (N_2416,N_1322,N_1365);
nand U2417 (N_2417,N_1268,N_1139);
nand U2418 (N_2418,N_1815,N_1032);
and U2419 (N_2419,N_1049,N_1385);
xor U2420 (N_2420,N_1153,N_1318);
xor U2421 (N_2421,N_1394,N_1167);
or U2422 (N_2422,N_1232,N_1435);
nor U2423 (N_2423,N_1329,N_1931);
and U2424 (N_2424,N_1735,N_1833);
xor U2425 (N_2425,N_1442,N_1691);
nor U2426 (N_2426,N_1274,N_1030);
or U2427 (N_2427,N_1209,N_1750);
xor U2428 (N_2428,N_1022,N_1543);
nand U2429 (N_2429,N_1640,N_1899);
nand U2430 (N_2430,N_1494,N_1704);
or U2431 (N_2431,N_1261,N_1101);
or U2432 (N_2432,N_1624,N_1715);
xor U2433 (N_2433,N_1726,N_1127);
nand U2434 (N_2434,N_1293,N_1475);
nor U2435 (N_2435,N_1076,N_1755);
nor U2436 (N_2436,N_1693,N_1389);
nor U2437 (N_2437,N_1900,N_1743);
nand U2438 (N_2438,N_1300,N_1653);
nor U2439 (N_2439,N_1978,N_1584);
or U2440 (N_2440,N_1066,N_1854);
and U2441 (N_2441,N_1434,N_1418);
xor U2442 (N_2442,N_1960,N_1649);
nand U2443 (N_2443,N_1020,N_1661);
or U2444 (N_2444,N_1781,N_1328);
and U2445 (N_2445,N_1001,N_1673);
and U2446 (N_2446,N_1937,N_1794);
xor U2447 (N_2447,N_1929,N_1736);
nand U2448 (N_2448,N_1998,N_1985);
or U2449 (N_2449,N_1414,N_1739);
nand U2450 (N_2450,N_1176,N_1186);
xor U2451 (N_2451,N_1447,N_1742);
nor U2452 (N_2452,N_1251,N_1669);
and U2453 (N_2453,N_1443,N_1882);
nand U2454 (N_2454,N_1868,N_1047);
xor U2455 (N_2455,N_1468,N_1005);
or U2456 (N_2456,N_1016,N_1436);
nand U2457 (N_2457,N_1295,N_1883);
nand U2458 (N_2458,N_1977,N_1546);
xnor U2459 (N_2459,N_1896,N_1248);
nor U2460 (N_2460,N_1712,N_1348);
nor U2461 (N_2461,N_1852,N_1215);
xor U2462 (N_2462,N_1147,N_1974);
and U2463 (N_2463,N_1320,N_1282);
or U2464 (N_2464,N_1012,N_1861);
xnor U2465 (N_2465,N_1965,N_1169);
xnor U2466 (N_2466,N_1413,N_1716);
and U2467 (N_2467,N_1933,N_1134);
and U2468 (N_2468,N_1252,N_1313);
or U2469 (N_2469,N_1323,N_1227);
xnor U2470 (N_2470,N_1986,N_1458);
xor U2471 (N_2471,N_1401,N_1184);
or U2472 (N_2472,N_1088,N_1275);
nand U2473 (N_2473,N_1651,N_1130);
nand U2474 (N_2474,N_1873,N_1219);
or U2475 (N_2475,N_1151,N_1345);
nand U2476 (N_2476,N_1628,N_1070);
and U2477 (N_2477,N_1230,N_1390);
or U2478 (N_2478,N_1773,N_1079);
and U2479 (N_2479,N_1874,N_1648);
nor U2480 (N_2480,N_1483,N_1946);
nand U2481 (N_2481,N_1876,N_1392);
nor U2482 (N_2482,N_1460,N_1954);
nand U2483 (N_2483,N_1880,N_1173);
nor U2484 (N_2484,N_1763,N_1226);
nand U2485 (N_2485,N_1558,N_1336);
xor U2486 (N_2486,N_1438,N_1080);
xnor U2487 (N_2487,N_1722,N_1867);
xnor U2488 (N_2488,N_1622,N_1433);
nor U2489 (N_2489,N_1136,N_1270);
nand U2490 (N_2490,N_1172,N_1760);
xor U2491 (N_2491,N_1486,N_1171);
xor U2492 (N_2492,N_1958,N_1921);
nor U2493 (N_2493,N_1073,N_1023);
nor U2494 (N_2494,N_1851,N_1140);
nand U2495 (N_2495,N_1516,N_1196);
and U2496 (N_2496,N_1567,N_1658);
xnor U2497 (N_2497,N_1051,N_1489);
or U2498 (N_2498,N_1000,N_1922);
and U2499 (N_2499,N_1031,N_1832);
and U2500 (N_2500,N_1677,N_1990);
nor U2501 (N_2501,N_1475,N_1832);
xor U2502 (N_2502,N_1615,N_1510);
xor U2503 (N_2503,N_1113,N_1662);
and U2504 (N_2504,N_1734,N_1474);
or U2505 (N_2505,N_1676,N_1609);
xor U2506 (N_2506,N_1445,N_1484);
xor U2507 (N_2507,N_1349,N_1522);
or U2508 (N_2508,N_1490,N_1322);
nand U2509 (N_2509,N_1284,N_1381);
xnor U2510 (N_2510,N_1758,N_1383);
nor U2511 (N_2511,N_1775,N_1695);
xnor U2512 (N_2512,N_1396,N_1490);
and U2513 (N_2513,N_1003,N_1742);
or U2514 (N_2514,N_1192,N_1888);
nand U2515 (N_2515,N_1941,N_1535);
xnor U2516 (N_2516,N_1390,N_1247);
nand U2517 (N_2517,N_1591,N_1934);
or U2518 (N_2518,N_1421,N_1946);
nand U2519 (N_2519,N_1642,N_1424);
nor U2520 (N_2520,N_1205,N_1534);
nand U2521 (N_2521,N_1727,N_1180);
nand U2522 (N_2522,N_1159,N_1084);
nand U2523 (N_2523,N_1069,N_1634);
nor U2524 (N_2524,N_1041,N_1167);
or U2525 (N_2525,N_1192,N_1702);
and U2526 (N_2526,N_1956,N_1727);
xor U2527 (N_2527,N_1121,N_1612);
and U2528 (N_2528,N_1659,N_1052);
or U2529 (N_2529,N_1876,N_1305);
or U2530 (N_2530,N_1977,N_1648);
nand U2531 (N_2531,N_1622,N_1068);
or U2532 (N_2532,N_1282,N_1180);
nor U2533 (N_2533,N_1508,N_1645);
xor U2534 (N_2534,N_1607,N_1026);
or U2535 (N_2535,N_1157,N_1915);
and U2536 (N_2536,N_1503,N_1006);
or U2537 (N_2537,N_1826,N_1141);
nand U2538 (N_2538,N_1567,N_1117);
and U2539 (N_2539,N_1674,N_1788);
nand U2540 (N_2540,N_1235,N_1894);
and U2541 (N_2541,N_1482,N_1519);
and U2542 (N_2542,N_1621,N_1717);
xnor U2543 (N_2543,N_1717,N_1122);
xor U2544 (N_2544,N_1761,N_1870);
or U2545 (N_2545,N_1080,N_1532);
or U2546 (N_2546,N_1138,N_1096);
nand U2547 (N_2547,N_1070,N_1439);
and U2548 (N_2548,N_1536,N_1040);
and U2549 (N_2549,N_1054,N_1483);
xnor U2550 (N_2550,N_1452,N_1826);
or U2551 (N_2551,N_1190,N_1339);
nand U2552 (N_2552,N_1841,N_1247);
or U2553 (N_2553,N_1540,N_1340);
xor U2554 (N_2554,N_1821,N_1963);
xnor U2555 (N_2555,N_1902,N_1117);
xor U2556 (N_2556,N_1055,N_1845);
or U2557 (N_2557,N_1194,N_1899);
xor U2558 (N_2558,N_1936,N_1332);
or U2559 (N_2559,N_1359,N_1496);
nand U2560 (N_2560,N_1098,N_1299);
and U2561 (N_2561,N_1314,N_1780);
xnor U2562 (N_2562,N_1084,N_1468);
and U2563 (N_2563,N_1041,N_1859);
nand U2564 (N_2564,N_1265,N_1795);
nor U2565 (N_2565,N_1934,N_1663);
xnor U2566 (N_2566,N_1214,N_1529);
nor U2567 (N_2567,N_1271,N_1120);
nand U2568 (N_2568,N_1199,N_1209);
or U2569 (N_2569,N_1348,N_1097);
or U2570 (N_2570,N_1756,N_1810);
nand U2571 (N_2571,N_1230,N_1081);
or U2572 (N_2572,N_1953,N_1897);
xor U2573 (N_2573,N_1000,N_1611);
xor U2574 (N_2574,N_1915,N_1024);
or U2575 (N_2575,N_1902,N_1164);
and U2576 (N_2576,N_1336,N_1467);
and U2577 (N_2577,N_1601,N_1724);
xnor U2578 (N_2578,N_1095,N_1029);
nand U2579 (N_2579,N_1659,N_1314);
and U2580 (N_2580,N_1185,N_1647);
nor U2581 (N_2581,N_1623,N_1065);
or U2582 (N_2582,N_1744,N_1019);
xor U2583 (N_2583,N_1690,N_1867);
nor U2584 (N_2584,N_1071,N_1017);
or U2585 (N_2585,N_1318,N_1872);
xnor U2586 (N_2586,N_1695,N_1353);
or U2587 (N_2587,N_1071,N_1918);
xor U2588 (N_2588,N_1740,N_1959);
and U2589 (N_2589,N_1493,N_1118);
nand U2590 (N_2590,N_1264,N_1966);
or U2591 (N_2591,N_1438,N_1613);
and U2592 (N_2592,N_1530,N_1472);
xor U2593 (N_2593,N_1592,N_1647);
nand U2594 (N_2594,N_1198,N_1343);
nor U2595 (N_2595,N_1942,N_1531);
nand U2596 (N_2596,N_1739,N_1631);
or U2597 (N_2597,N_1728,N_1312);
and U2598 (N_2598,N_1844,N_1163);
and U2599 (N_2599,N_1111,N_1283);
nor U2600 (N_2600,N_1348,N_1869);
nor U2601 (N_2601,N_1313,N_1483);
xnor U2602 (N_2602,N_1832,N_1406);
or U2603 (N_2603,N_1211,N_1225);
nor U2604 (N_2604,N_1999,N_1438);
nand U2605 (N_2605,N_1627,N_1436);
or U2606 (N_2606,N_1040,N_1254);
or U2607 (N_2607,N_1750,N_1239);
and U2608 (N_2608,N_1968,N_1528);
and U2609 (N_2609,N_1110,N_1224);
and U2610 (N_2610,N_1631,N_1885);
and U2611 (N_2611,N_1824,N_1699);
xnor U2612 (N_2612,N_1838,N_1041);
nand U2613 (N_2613,N_1235,N_1123);
or U2614 (N_2614,N_1678,N_1827);
nand U2615 (N_2615,N_1332,N_1135);
nand U2616 (N_2616,N_1092,N_1713);
xor U2617 (N_2617,N_1731,N_1100);
nor U2618 (N_2618,N_1641,N_1632);
nor U2619 (N_2619,N_1959,N_1673);
or U2620 (N_2620,N_1219,N_1035);
nor U2621 (N_2621,N_1947,N_1262);
xor U2622 (N_2622,N_1416,N_1326);
and U2623 (N_2623,N_1943,N_1893);
nand U2624 (N_2624,N_1093,N_1208);
and U2625 (N_2625,N_1228,N_1672);
nor U2626 (N_2626,N_1504,N_1147);
nand U2627 (N_2627,N_1205,N_1903);
xor U2628 (N_2628,N_1842,N_1346);
xor U2629 (N_2629,N_1645,N_1662);
nor U2630 (N_2630,N_1612,N_1855);
or U2631 (N_2631,N_1182,N_1934);
nand U2632 (N_2632,N_1106,N_1641);
and U2633 (N_2633,N_1814,N_1246);
nor U2634 (N_2634,N_1972,N_1107);
nor U2635 (N_2635,N_1166,N_1065);
or U2636 (N_2636,N_1882,N_1478);
nand U2637 (N_2637,N_1738,N_1928);
nand U2638 (N_2638,N_1398,N_1300);
or U2639 (N_2639,N_1004,N_1110);
or U2640 (N_2640,N_1742,N_1907);
or U2641 (N_2641,N_1074,N_1364);
and U2642 (N_2642,N_1382,N_1665);
nand U2643 (N_2643,N_1076,N_1645);
nor U2644 (N_2644,N_1623,N_1287);
or U2645 (N_2645,N_1284,N_1966);
nor U2646 (N_2646,N_1442,N_1278);
and U2647 (N_2647,N_1137,N_1008);
nor U2648 (N_2648,N_1035,N_1608);
or U2649 (N_2649,N_1483,N_1752);
xnor U2650 (N_2650,N_1013,N_1361);
nand U2651 (N_2651,N_1113,N_1931);
or U2652 (N_2652,N_1093,N_1107);
xnor U2653 (N_2653,N_1711,N_1717);
nor U2654 (N_2654,N_1139,N_1507);
or U2655 (N_2655,N_1688,N_1488);
or U2656 (N_2656,N_1111,N_1035);
nor U2657 (N_2657,N_1339,N_1149);
nor U2658 (N_2658,N_1323,N_1869);
or U2659 (N_2659,N_1977,N_1068);
or U2660 (N_2660,N_1982,N_1758);
nand U2661 (N_2661,N_1022,N_1128);
xor U2662 (N_2662,N_1652,N_1490);
and U2663 (N_2663,N_1324,N_1774);
xnor U2664 (N_2664,N_1091,N_1956);
nand U2665 (N_2665,N_1256,N_1882);
nor U2666 (N_2666,N_1165,N_1133);
nor U2667 (N_2667,N_1634,N_1012);
and U2668 (N_2668,N_1202,N_1642);
xor U2669 (N_2669,N_1101,N_1005);
nor U2670 (N_2670,N_1334,N_1057);
or U2671 (N_2671,N_1518,N_1066);
nor U2672 (N_2672,N_1851,N_1936);
nand U2673 (N_2673,N_1300,N_1657);
or U2674 (N_2674,N_1184,N_1690);
nor U2675 (N_2675,N_1886,N_1846);
or U2676 (N_2676,N_1847,N_1480);
or U2677 (N_2677,N_1771,N_1288);
and U2678 (N_2678,N_1842,N_1859);
xnor U2679 (N_2679,N_1349,N_1253);
nor U2680 (N_2680,N_1964,N_1853);
nor U2681 (N_2681,N_1457,N_1785);
nand U2682 (N_2682,N_1653,N_1800);
nor U2683 (N_2683,N_1381,N_1032);
and U2684 (N_2684,N_1597,N_1893);
and U2685 (N_2685,N_1126,N_1272);
and U2686 (N_2686,N_1221,N_1457);
or U2687 (N_2687,N_1373,N_1119);
nand U2688 (N_2688,N_1276,N_1857);
xor U2689 (N_2689,N_1084,N_1606);
or U2690 (N_2690,N_1747,N_1979);
or U2691 (N_2691,N_1938,N_1365);
xnor U2692 (N_2692,N_1493,N_1669);
and U2693 (N_2693,N_1377,N_1621);
xnor U2694 (N_2694,N_1833,N_1893);
xnor U2695 (N_2695,N_1266,N_1388);
xor U2696 (N_2696,N_1608,N_1206);
nor U2697 (N_2697,N_1982,N_1485);
or U2698 (N_2698,N_1556,N_1115);
xnor U2699 (N_2699,N_1276,N_1380);
and U2700 (N_2700,N_1501,N_1786);
nor U2701 (N_2701,N_1927,N_1027);
and U2702 (N_2702,N_1103,N_1240);
or U2703 (N_2703,N_1977,N_1167);
and U2704 (N_2704,N_1421,N_1556);
and U2705 (N_2705,N_1519,N_1693);
and U2706 (N_2706,N_1343,N_1460);
nand U2707 (N_2707,N_1754,N_1208);
or U2708 (N_2708,N_1780,N_1332);
nand U2709 (N_2709,N_1950,N_1015);
nand U2710 (N_2710,N_1526,N_1869);
nand U2711 (N_2711,N_1778,N_1043);
xnor U2712 (N_2712,N_1527,N_1728);
nand U2713 (N_2713,N_1389,N_1841);
nand U2714 (N_2714,N_1423,N_1215);
and U2715 (N_2715,N_1860,N_1382);
nor U2716 (N_2716,N_1926,N_1039);
or U2717 (N_2717,N_1475,N_1869);
nor U2718 (N_2718,N_1859,N_1629);
xor U2719 (N_2719,N_1537,N_1740);
nor U2720 (N_2720,N_1215,N_1925);
or U2721 (N_2721,N_1958,N_1076);
and U2722 (N_2722,N_1438,N_1516);
nor U2723 (N_2723,N_1303,N_1498);
xnor U2724 (N_2724,N_1054,N_1201);
nor U2725 (N_2725,N_1328,N_1471);
nand U2726 (N_2726,N_1195,N_1050);
nand U2727 (N_2727,N_1403,N_1602);
and U2728 (N_2728,N_1827,N_1117);
or U2729 (N_2729,N_1936,N_1075);
or U2730 (N_2730,N_1073,N_1425);
and U2731 (N_2731,N_1120,N_1570);
xnor U2732 (N_2732,N_1613,N_1140);
nor U2733 (N_2733,N_1960,N_1973);
nand U2734 (N_2734,N_1463,N_1695);
xor U2735 (N_2735,N_1766,N_1188);
or U2736 (N_2736,N_1096,N_1205);
xor U2737 (N_2737,N_1902,N_1904);
xor U2738 (N_2738,N_1126,N_1182);
nor U2739 (N_2739,N_1268,N_1252);
nand U2740 (N_2740,N_1196,N_1904);
or U2741 (N_2741,N_1915,N_1331);
nor U2742 (N_2742,N_1867,N_1897);
or U2743 (N_2743,N_1199,N_1509);
xnor U2744 (N_2744,N_1994,N_1548);
or U2745 (N_2745,N_1582,N_1256);
and U2746 (N_2746,N_1678,N_1999);
or U2747 (N_2747,N_1221,N_1323);
and U2748 (N_2748,N_1467,N_1604);
nand U2749 (N_2749,N_1057,N_1419);
or U2750 (N_2750,N_1833,N_1216);
xor U2751 (N_2751,N_1876,N_1427);
nand U2752 (N_2752,N_1877,N_1191);
or U2753 (N_2753,N_1002,N_1569);
xor U2754 (N_2754,N_1354,N_1487);
or U2755 (N_2755,N_1059,N_1707);
nand U2756 (N_2756,N_1241,N_1726);
nor U2757 (N_2757,N_1243,N_1101);
or U2758 (N_2758,N_1597,N_1814);
nor U2759 (N_2759,N_1079,N_1997);
nand U2760 (N_2760,N_1248,N_1716);
xor U2761 (N_2761,N_1037,N_1036);
and U2762 (N_2762,N_1281,N_1342);
or U2763 (N_2763,N_1026,N_1218);
and U2764 (N_2764,N_1826,N_1937);
xnor U2765 (N_2765,N_1838,N_1621);
nand U2766 (N_2766,N_1890,N_1316);
and U2767 (N_2767,N_1819,N_1118);
xnor U2768 (N_2768,N_1476,N_1801);
xnor U2769 (N_2769,N_1888,N_1325);
nor U2770 (N_2770,N_1362,N_1838);
nor U2771 (N_2771,N_1928,N_1608);
and U2772 (N_2772,N_1305,N_1233);
or U2773 (N_2773,N_1641,N_1517);
or U2774 (N_2774,N_1961,N_1798);
or U2775 (N_2775,N_1785,N_1672);
nand U2776 (N_2776,N_1616,N_1935);
nor U2777 (N_2777,N_1992,N_1534);
nor U2778 (N_2778,N_1441,N_1889);
xor U2779 (N_2779,N_1080,N_1629);
and U2780 (N_2780,N_1062,N_1643);
xor U2781 (N_2781,N_1040,N_1682);
or U2782 (N_2782,N_1574,N_1960);
nand U2783 (N_2783,N_1331,N_1761);
nand U2784 (N_2784,N_1325,N_1693);
or U2785 (N_2785,N_1267,N_1591);
nor U2786 (N_2786,N_1826,N_1329);
nand U2787 (N_2787,N_1499,N_1717);
xor U2788 (N_2788,N_1547,N_1106);
xor U2789 (N_2789,N_1854,N_1572);
nand U2790 (N_2790,N_1852,N_1973);
xnor U2791 (N_2791,N_1886,N_1856);
or U2792 (N_2792,N_1800,N_1343);
xnor U2793 (N_2793,N_1154,N_1183);
nor U2794 (N_2794,N_1445,N_1630);
or U2795 (N_2795,N_1261,N_1928);
and U2796 (N_2796,N_1592,N_1439);
and U2797 (N_2797,N_1110,N_1121);
or U2798 (N_2798,N_1052,N_1515);
and U2799 (N_2799,N_1441,N_1052);
or U2800 (N_2800,N_1607,N_1918);
nand U2801 (N_2801,N_1718,N_1196);
or U2802 (N_2802,N_1518,N_1824);
and U2803 (N_2803,N_1279,N_1524);
nand U2804 (N_2804,N_1338,N_1409);
nand U2805 (N_2805,N_1269,N_1094);
nor U2806 (N_2806,N_1239,N_1546);
nand U2807 (N_2807,N_1402,N_1673);
nand U2808 (N_2808,N_1113,N_1412);
xor U2809 (N_2809,N_1948,N_1456);
and U2810 (N_2810,N_1368,N_1753);
nor U2811 (N_2811,N_1549,N_1569);
nand U2812 (N_2812,N_1949,N_1603);
nand U2813 (N_2813,N_1750,N_1119);
nor U2814 (N_2814,N_1253,N_1067);
and U2815 (N_2815,N_1758,N_1954);
nor U2816 (N_2816,N_1954,N_1449);
nor U2817 (N_2817,N_1050,N_1361);
nand U2818 (N_2818,N_1918,N_1147);
nor U2819 (N_2819,N_1156,N_1247);
xnor U2820 (N_2820,N_1805,N_1317);
or U2821 (N_2821,N_1699,N_1320);
nor U2822 (N_2822,N_1963,N_1773);
nor U2823 (N_2823,N_1265,N_1449);
nor U2824 (N_2824,N_1613,N_1059);
xor U2825 (N_2825,N_1128,N_1135);
and U2826 (N_2826,N_1113,N_1009);
and U2827 (N_2827,N_1105,N_1341);
or U2828 (N_2828,N_1068,N_1930);
nor U2829 (N_2829,N_1240,N_1269);
or U2830 (N_2830,N_1427,N_1073);
or U2831 (N_2831,N_1811,N_1853);
nand U2832 (N_2832,N_1836,N_1060);
nand U2833 (N_2833,N_1712,N_1743);
xnor U2834 (N_2834,N_1573,N_1504);
nor U2835 (N_2835,N_1624,N_1350);
xnor U2836 (N_2836,N_1889,N_1140);
nand U2837 (N_2837,N_1511,N_1130);
nand U2838 (N_2838,N_1781,N_1736);
or U2839 (N_2839,N_1618,N_1664);
nor U2840 (N_2840,N_1787,N_1617);
xor U2841 (N_2841,N_1650,N_1010);
and U2842 (N_2842,N_1792,N_1813);
nor U2843 (N_2843,N_1654,N_1723);
nand U2844 (N_2844,N_1848,N_1189);
or U2845 (N_2845,N_1573,N_1937);
or U2846 (N_2846,N_1390,N_1232);
or U2847 (N_2847,N_1409,N_1135);
nor U2848 (N_2848,N_1595,N_1933);
and U2849 (N_2849,N_1162,N_1438);
nor U2850 (N_2850,N_1047,N_1912);
or U2851 (N_2851,N_1544,N_1429);
and U2852 (N_2852,N_1343,N_1455);
nor U2853 (N_2853,N_1209,N_1292);
or U2854 (N_2854,N_1239,N_1917);
and U2855 (N_2855,N_1197,N_1971);
and U2856 (N_2856,N_1473,N_1135);
xor U2857 (N_2857,N_1939,N_1771);
xnor U2858 (N_2858,N_1057,N_1533);
and U2859 (N_2859,N_1048,N_1469);
xnor U2860 (N_2860,N_1620,N_1689);
nand U2861 (N_2861,N_1003,N_1894);
nand U2862 (N_2862,N_1538,N_1745);
nor U2863 (N_2863,N_1158,N_1641);
or U2864 (N_2864,N_1390,N_1079);
xor U2865 (N_2865,N_1584,N_1398);
xor U2866 (N_2866,N_1895,N_1921);
xor U2867 (N_2867,N_1379,N_1088);
xor U2868 (N_2868,N_1512,N_1638);
xnor U2869 (N_2869,N_1941,N_1175);
and U2870 (N_2870,N_1260,N_1730);
or U2871 (N_2871,N_1408,N_1970);
and U2872 (N_2872,N_1690,N_1296);
nor U2873 (N_2873,N_1311,N_1209);
and U2874 (N_2874,N_1166,N_1600);
nand U2875 (N_2875,N_1204,N_1407);
or U2876 (N_2876,N_1181,N_1283);
xor U2877 (N_2877,N_1002,N_1453);
nor U2878 (N_2878,N_1472,N_1511);
nor U2879 (N_2879,N_1426,N_1266);
xor U2880 (N_2880,N_1397,N_1191);
or U2881 (N_2881,N_1350,N_1874);
nand U2882 (N_2882,N_1188,N_1978);
nor U2883 (N_2883,N_1307,N_1058);
and U2884 (N_2884,N_1299,N_1499);
or U2885 (N_2885,N_1034,N_1773);
nor U2886 (N_2886,N_1017,N_1552);
and U2887 (N_2887,N_1495,N_1825);
and U2888 (N_2888,N_1013,N_1932);
nand U2889 (N_2889,N_1963,N_1003);
or U2890 (N_2890,N_1392,N_1140);
nand U2891 (N_2891,N_1236,N_1467);
and U2892 (N_2892,N_1000,N_1703);
and U2893 (N_2893,N_1780,N_1330);
or U2894 (N_2894,N_1210,N_1864);
nand U2895 (N_2895,N_1618,N_1977);
nor U2896 (N_2896,N_1556,N_1273);
nor U2897 (N_2897,N_1812,N_1609);
or U2898 (N_2898,N_1887,N_1520);
and U2899 (N_2899,N_1266,N_1716);
or U2900 (N_2900,N_1262,N_1370);
nor U2901 (N_2901,N_1682,N_1772);
xnor U2902 (N_2902,N_1345,N_1020);
nor U2903 (N_2903,N_1173,N_1850);
nor U2904 (N_2904,N_1066,N_1341);
or U2905 (N_2905,N_1169,N_1438);
nor U2906 (N_2906,N_1056,N_1300);
nor U2907 (N_2907,N_1876,N_1057);
xor U2908 (N_2908,N_1563,N_1178);
xor U2909 (N_2909,N_1659,N_1471);
nand U2910 (N_2910,N_1371,N_1256);
nor U2911 (N_2911,N_1151,N_1154);
or U2912 (N_2912,N_1477,N_1808);
and U2913 (N_2913,N_1825,N_1947);
nor U2914 (N_2914,N_1176,N_1771);
nor U2915 (N_2915,N_1086,N_1929);
xnor U2916 (N_2916,N_1540,N_1293);
and U2917 (N_2917,N_1251,N_1323);
or U2918 (N_2918,N_1779,N_1026);
and U2919 (N_2919,N_1061,N_1252);
nand U2920 (N_2920,N_1706,N_1788);
nor U2921 (N_2921,N_1701,N_1755);
xor U2922 (N_2922,N_1878,N_1038);
xor U2923 (N_2923,N_1221,N_1446);
or U2924 (N_2924,N_1623,N_1988);
nor U2925 (N_2925,N_1105,N_1832);
xor U2926 (N_2926,N_1199,N_1262);
nand U2927 (N_2927,N_1260,N_1406);
and U2928 (N_2928,N_1695,N_1364);
nand U2929 (N_2929,N_1946,N_1923);
nand U2930 (N_2930,N_1815,N_1607);
or U2931 (N_2931,N_1751,N_1464);
nand U2932 (N_2932,N_1178,N_1676);
nor U2933 (N_2933,N_1934,N_1337);
and U2934 (N_2934,N_1097,N_1715);
nand U2935 (N_2935,N_1824,N_1952);
or U2936 (N_2936,N_1984,N_1411);
or U2937 (N_2937,N_1877,N_1216);
xor U2938 (N_2938,N_1454,N_1560);
nand U2939 (N_2939,N_1391,N_1513);
and U2940 (N_2940,N_1991,N_1862);
nand U2941 (N_2941,N_1992,N_1382);
and U2942 (N_2942,N_1199,N_1653);
nand U2943 (N_2943,N_1702,N_1366);
nor U2944 (N_2944,N_1485,N_1096);
xnor U2945 (N_2945,N_1719,N_1349);
nor U2946 (N_2946,N_1724,N_1221);
or U2947 (N_2947,N_1424,N_1589);
or U2948 (N_2948,N_1084,N_1986);
or U2949 (N_2949,N_1924,N_1505);
and U2950 (N_2950,N_1068,N_1069);
xnor U2951 (N_2951,N_1464,N_1298);
or U2952 (N_2952,N_1152,N_1294);
and U2953 (N_2953,N_1649,N_1444);
and U2954 (N_2954,N_1611,N_1682);
nor U2955 (N_2955,N_1020,N_1089);
nor U2956 (N_2956,N_1492,N_1242);
xor U2957 (N_2957,N_1494,N_1445);
xor U2958 (N_2958,N_1424,N_1681);
xor U2959 (N_2959,N_1084,N_1509);
nor U2960 (N_2960,N_1635,N_1041);
or U2961 (N_2961,N_1042,N_1923);
nor U2962 (N_2962,N_1261,N_1672);
xor U2963 (N_2963,N_1077,N_1857);
and U2964 (N_2964,N_1705,N_1327);
or U2965 (N_2965,N_1446,N_1671);
xnor U2966 (N_2966,N_1180,N_1602);
nand U2967 (N_2967,N_1242,N_1598);
nand U2968 (N_2968,N_1005,N_1835);
or U2969 (N_2969,N_1934,N_1598);
or U2970 (N_2970,N_1487,N_1462);
xor U2971 (N_2971,N_1925,N_1705);
and U2972 (N_2972,N_1869,N_1403);
nor U2973 (N_2973,N_1995,N_1597);
xnor U2974 (N_2974,N_1113,N_1035);
nand U2975 (N_2975,N_1835,N_1819);
xnor U2976 (N_2976,N_1784,N_1010);
nand U2977 (N_2977,N_1582,N_1882);
and U2978 (N_2978,N_1904,N_1776);
xor U2979 (N_2979,N_1324,N_1299);
or U2980 (N_2980,N_1610,N_1660);
nor U2981 (N_2981,N_1078,N_1199);
and U2982 (N_2982,N_1669,N_1195);
nand U2983 (N_2983,N_1346,N_1144);
nor U2984 (N_2984,N_1650,N_1602);
nand U2985 (N_2985,N_1000,N_1295);
nor U2986 (N_2986,N_1376,N_1392);
or U2987 (N_2987,N_1667,N_1124);
nand U2988 (N_2988,N_1428,N_1078);
or U2989 (N_2989,N_1555,N_1917);
nor U2990 (N_2990,N_1570,N_1965);
nand U2991 (N_2991,N_1436,N_1609);
xor U2992 (N_2992,N_1716,N_1040);
nand U2993 (N_2993,N_1302,N_1249);
nor U2994 (N_2994,N_1828,N_1979);
nand U2995 (N_2995,N_1268,N_1059);
and U2996 (N_2996,N_1302,N_1253);
and U2997 (N_2997,N_1462,N_1193);
nor U2998 (N_2998,N_1543,N_1807);
nor U2999 (N_2999,N_1995,N_1929);
nor U3000 (N_3000,N_2638,N_2179);
nor U3001 (N_3001,N_2618,N_2234);
nand U3002 (N_3002,N_2743,N_2015);
nor U3003 (N_3003,N_2485,N_2938);
and U3004 (N_3004,N_2439,N_2251);
xor U3005 (N_3005,N_2785,N_2929);
xnor U3006 (N_3006,N_2865,N_2242);
nor U3007 (N_3007,N_2308,N_2620);
xnor U3008 (N_3008,N_2721,N_2367);
and U3009 (N_3009,N_2222,N_2874);
and U3010 (N_3010,N_2417,N_2004);
nor U3011 (N_3011,N_2952,N_2023);
nor U3012 (N_3012,N_2059,N_2118);
or U3013 (N_3013,N_2724,N_2800);
or U3014 (N_3014,N_2748,N_2052);
xnor U3015 (N_3015,N_2986,N_2840);
and U3016 (N_3016,N_2925,N_2658);
and U3017 (N_3017,N_2038,N_2003);
xor U3018 (N_3018,N_2745,N_2751);
and U3019 (N_3019,N_2292,N_2821);
nand U3020 (N_3020,N_2582,N_2138);
or U3021 (N_3021,N_2271,N_2685);
nor U3022 (N_3022,N_2306,N_2054);
or U3023 (N_3023,N_2686,N_2568);
or U3024 (N_3024,N_2274,N_2924);
or U3025 (N_3025,N_2894,N_2550);
or U3026 (N_3026,N_2132,N_2285);
nand U3027 (N_3027,N_2590,N_2882);
and U3028 (N_3028,N_2357,N_2825);
and U3029 (N_3029,N_2915,N_2127);
or U3030 (N_3030,N_2290,N_2967);
xnor U3031 (N_3031,N_2476,N_2622);
or U3032 (N_3032,N_2948,N_2223);
or U3033 (N_3033,N_2573,N_2598);
nand U3034 (N_3034,N_2906,N_2364);
or U3035 (N_3035,N_2529,N_2885);
and U3036 (N_3036,N_2642,N_2451);
and U3037 (N_3037,N_2407,N_2495);
or U3038 (N_3038,N_2551,N_2481);
xor U3039 (N_3039,N_2231,N_2062);
nor U3040 (N_3040,N_2478,N_2207);
and U3041 (N_3041,N_2419,N_2266);
and U3042 (N_3042,N_2583,N_2810);
xor U3043 (N_3043,N_2695,N_2258);
nand U3044 (N_3044,N_2414,N_2307);
nor U3045 (N_3045,N_2471,N_2098);
nor U3046 (N_3046,N_2103,N_2682);
nand U3047 (N_3047,N_2169,N_2978);
nand U3048 (N_3048,N_2775,N_2280);
or U3049 (N_3049,N_2377,N_2097);
and U3050 (N_3050,N_2965,N_2617);
and U3051 (N_3051,N_2596,N_2764);
or U3052 (N_3052,N_2216,N_2613);
nand U3053 (N_3053,N_2463,N_2755);
or U3054 (N_3054,N_2096,N_2650);
and U3055 (N_3055,N_2700,N_2786);
or U3056 (N_3056,N_2574,N_2387);
and U3057 (N_3057,N_2698,N_2637);
xnor U3058 (N_3058,N_2202,N_2589);
nand U3059 (N_3059,N_2022,N_2697);
nor U3060 (N_3060,N_2465,N_2099);
nor U3061 (N_3061,N_2656,N_2475);
nor U3062 (N_3062,N_2887,N_2790);
nor U3063 (N_3063,N_2851,N_2980);
or U3064 (N_3064,N_2789,N_2516);
or U3065 (N_3065,N_2181,N_2832);
and U3066 (N_3066,N_2296,N_2368);
or U3067 (N_3067,N_2560,N_2146);
and U3068 (N_3068,N_2005,N_2160);
and U3069 (N_3069,N_2892,N_2229);
and U3070 (N_3070,N_2442,N_2415);
nand U3071 (N_3071,N_2241,N_2677);
nor U3072 (N_3072,N_2195,N_2544);
xnor U3073 (N_3073,N_2384,N_2155);
nor U3074 (N_3074,N_2166,N_2014);
nor U3075 (N_3075,N_2016,N_2288);
and U3076 (N_3076,N_2131,N_2346);
and U3077 (N_3077,N_2089,N_2467);
nor U3078 (N_3078,N_2802,N_2689);
nand U3079 (N_3079,N_2171,N_2740);
nor U3080 (N_3080,N_2612,N_2850);
xnor U3081 (N_3081,N_2629,N_2591);
xor U3082 (N_3082,N_2873,N_2900);
nand U3083 (N_3083,N_2153,N_2259);
and U3084 (N_3084,N_2219,N_2683);
nand U3085 (N_3085,N_2774,N_2738);
xnor U3086 (N_3086,N_2453,N_2142);
or U3087 (N_3087,N_2607,N_2049);
and U3088 (N_3088,N_2730,N_2958);
xor U3089 (N_3089,N_2326,N_2483);
nand U3090 (N_3090,N_2860,N_2902);
or U3091 (N_3091,N_2907,N_2389);
xnor U3092 (N_3092,N_2606,N_2563);
xor U3093 (N_3093,N_2211,N_2408);
or U3094 (N_3094,N_2325,N_2149);
and U3095 (N_3095,N_2917,N_2007);
xnor U3096 (N_3096,N_2982,N_2659);
and U3097 (N_3097,N_2263,N_2634);
nor U3098 (N_3098,N_2916,N_2898);
or U3099 (N_3099,N_2939,N_2203);
nand U3100 (N_3100,N_2192,N_2517);
and U3101 (N_3101,N_2176,N_2469);
xor U3102 (N_3102,N_2552,N_2283);
nor U3103 (N_3103,N_2889,N_2114);
or U3104 (N_3104,N_2556,N_2024);
nand U3105 (N_3105,N_2742,N_2672);
and U3106 (N_3106,N_2433,N_2117);
xnor U3107 (N_3107,N_2933,N_2331);
nor U3108 (N_3108,N_2947,N_2190);
xor U3109 (N_3109,N_2776,N_2757);
or U3110 (N_3110,N_2173,N_2457);
and U3111 (N_3111,N_2979,N_2651);
or U3112 (N_3112,N_2150,N_2163);
xnor U3113 (N_3113,N_2093,N_2466);
xnor U3114 (N_3114,N_2393,N_2489);
or U3115 (N_3115,N_2675,N_2124);
nor U3116 (N_3116,N_2781,N_2328);
and U3117 (N_3117,N_2901,N_2218);
or U3118 (N_3118,N_2392,N_2069);
nand U3119 (N_3119,N_2831,N_2666);
nand U3120 (N_3120,N_2960,N_2238);
or U3121 (N_3121,N_2449,N_2320);
xnor U3122 (N_3122,N_2426,N_2652);
nand U3123 (N_3123,N_2968,N_2654);
xor U3124 (N_3124,N_2406,N_2541);
or U3125 (N_3125,N_2336,N_2795);
or U3126 (N_3126,N_2269,N_2196);
nor U3127 (N_3127,N_2010,N_2587);
xnor U3128 (N_3128,N_2987,N_2239);
nand U3129 (N_3129,N_2520,N_2311);
nor U3130 (N_3130,N_2429,N_2701);
and U3131 (N_3131,N_2177,N_2482);
xor U3132 (N_3132,N_2116,N_2107);
and U3133 (N_3133,N_2291,N_2298);
and U3134 (N_3134,N_2558,N_2995);
or U3135 (N_3135,N_2398,N_2616);
or U3136 (N_3136,N_2812,N_2625);
xnor U3137 (N_3137,N_2732,N_2914);
and U3138 (N_3138,N_2268,N_2610);
or U3139 (N_3139,N_2067,N_2145);
and U3140 (N_3140,N_2048,N_2773);
xnor U3141 (N_3141,N_2385,N_2567);
xnor U3142 (N_3142,N_2343,N_2856);
nand U3143 (N_3143,N_2646,N_2849);
or U3144 (N_3144,N_2147,N_2335);
nand U3145 (N_3145,N_2524,N_2603);
xor U3146 (N_3146,N_2782,N_2744);
and U3147 (N_3147,N_2382,N_2221);
nor U3148 (N_3148,N_2302,N_2655);
nor U3149 (N_3149,N_2844,N_2588);
nand U3150 (N_3150,N_2704,N_2746);
nand U3151 (N_3151,N_2926,N_2383);
nand U3152 (N_3152,N_2991,N_2714);
or U3153 (N_3153,N_2080,N_2792);
nor U3154 (N_3154,N_2324,N_2121);
and U3155 (N_3155,N_2394,N_2920);
nor U3156 (N_3156,N_2428,N_2454);
nor U3157 (N_3157,N_2162,N_2747);
nor U3158 (N_3158,N_2318,N_2521);
and U3159 (N_3159,N_2240,N_2799);
nor U3160 (N_3160,N_2531,N_2972);
nand U3161 (N_3161,N_2867,N_2621);
xnor U3162 (N_3162,N_2911,N_2858);
nand U3163 (N_3163,N_2963,N_2805);
or U3164 (N_3164,N_2673,N_2233);
nand U3165 (N_3165,N_2707,N_2758);
nand U3166 (N_3166,N_2660,N_2633);
xor U3167 (N_3167,N_2154,N_2962);
nand U3168 (N_3168,N_2055,N_2494);
and U3169 (N_3169,N_2643,N_2913);
and U3170 (N_3170,N_2694,N_2100);
and U3171 (N_3171,N_2768,N_2230);
nor U3172 (N_3172,N_2870,N_2314);
and U3173 (N_3173,N_2703,N_2039);
nor U3174 (N_3174,N_2820,N_2572);
or U3175 (N_3175,N_2455,N_2827);
or U3176 (N_3176,N_2985,N_2631);
or U3177 (N_3177,N_2272,N_2585);
and U3178 (N_3178,N_2853,N_2395);
xnor U3179 (N_3179,N_2593,N_2226);
and U3180 (N_3180,N_2510,N_2749);
nand U3181 (N_3181,N_2586,N_2765);
xor U3182 (N_3182,N_2305,N_2649);
and U3183 (N_3183,N_2896,N_2157);
and U3184 (N_3184,N_2555,N_2828);
or U3185 (N_3185,N_2668,N_2794);
and U3186 (N_3186,N_2605,N_2891);
and U3187 (N_3187,N_2813,N_2082);
and U3188 (N_3188,N_2806,N_2189);
nor U3189 (N_3189,N_2739,N_2206);
nand U3190 (N_3190,N_2514,N_2225);
nand U3191 (N_3191,N_2158,N_2340);
nor U3192 (N_3192,N_2111,N_2954);
or U3193 (N_3193,N_2198,N_2736);
nand U3194 (N_3194,N_2168,N_2330);
nand U3195 (N_3195,N_2945,N_2502);
xor U3196 (N_3196,N_2294,N_2281);
and U3197 (N_3197,N_2019,N_2456);
xor U3198 (N_3198,N_2361,N_2161);
xnor U3199 (N_3199,N_2632,N_2935);
nand U3200 (N_3200,N_2425,N_2974);
and U3201 (N_3201,N_2159,N_2505);
and U3202 (N_3202,N_2396,N_2791);
or U3203 (N_3203,N_2209,N_2122);
nand U3204 (N_3204,N_2872,N_2078);
or U3205 (N_3205,N_2577,N_2369);
nand U3206 (N_3206,N_2602,N_2033);
nand U3207 (N_3207,N_2303,N_2513);
or U3208 (N_3208,N_2255,N_2106);
xor U3209 (N_3209,N_2955,N_2564);
or U3210 (N_3210,N_2815,N_2741);
or U3211 (N_3211,N_2354,N_2769);
xnor U3212 (N_3212,N_2895,N_2623);
nand U3213 (N_3213,N_2446,N_2880);
nor U3214 (N_3214,N_2187,N_2058);
nand U3215 (N_3215,N_2112,N_2247);
xor U3216 (N_3216,N_2737,N_2923);
nand U3217 (N_3217,N_2075,N_2674);
and U3218 (N_3218,N_2254,N_2930);
xnor U3219 (N_3219,N_2983,N_2542);
or U3220 (N_3220,N_2752,N_2543);
nor U3221 (N_3221,N_2709,N_2105);
xnor U3222 (N_3222,N_2829,N_2879);
xor U3223 (N_3223,N_2708,N_2260);
or U3224 (N_3224,N_2057,N_2072);
xor U3225 (N_3225,N_2412,N_2964);
xnor U3226 (N_3226,N_2423,N_2779);
and U3227 (N_3227,N_2180,N_2569);
or U3228 (N_3228,N_2017,N_2140);
nor U3229 (N_3229,N_2644,N_2584);
and U3230 (N_3230,N_2422,N_2323);
nand U3231 (N_3231,N_2418,N_2990);
nand U3232 (N_3232,N_2546,N_2338);
xor U3233 (N_3233,N_2282,N_2904);
nor U3234 (N_3234,N_2090,N_2201);
or U3235 (N_3235,N_2042,N_2188);
or U3236 (N_3236,N_2277,N_2778);
and U3237 (N_3237,N_2988,N_2215);
xor U3238 (N_3238,N_2110,N_2854);
or U3239 (N_3239,N_2946,N_2380);
and U3240 (N_3240,N_2224,N_2375);
nor U3241 (N_3241,N_2819,N_2735);
nand U3242 (N_3242,N_2753,N_2044);
nand U3243 (N_3243,N_2886,N_2594);
nor U3244 (N_3244,N_2909,N_2399);
nand U3245 (N_3245,N_2578,N_2706);
or U3246 (N_3246,N_2458,N_2762);
xor U3247 (N_3247,N_2557,N_2506);
or U3248 (N_3248,N_2186,N_2763);
xnor U3249 (N_3249,N_2109,N_2966);
xor U3250 (N_3250,N_2645,N_2043);
nor U3251 (N_3251,N_2339,N_2691);
and U3252 (N_3252,N_2358,N_2403);
nand U3253 (N_3253,N_2562,N_2237);
or U3254 (N_3254,N_2136,N_2348);
and U3255 (N_3255,N_2848,N_2092);
nor U3256 (N_3256,N_2194,N_2671);
or U3257 (N_3257,N_2869,N_2611);
and U3258 (N_3258,N_2852,N_2085);
or U3259 (N_3259,N_2474,N_2797);
nand U3260 (N_3260,N_2178,N_2592);
and U3261 (N_3261,N_2728,N_2046);
nor U3262 (N_3262,N_2137,N_2530);
nor U3263 (N_3263,N_2711,N_2826);
and U3264 (N_3264,N_2910,N_2329);
nor U3265 (N_3265,N_2624,N_2445);
nor U3266 (N_3266,N_2197,N_2688);
nand U3267 (N_3267,N_2793,N_2528);
and U3268 (N_3268,N_2293,N_2888);
and U3269 (N_3269,N_2859,N_2717);
nand U3270 (N_3270,N_2006,N_2317);
or U3271 (N_3271,N_2561,N_2868);
and U3272 (N_3272,N_2811,N_2319);
or U3273 (N_3273,N_2554,N_2413);
nor U3274 (N_3274,N_2051,N_2205);
xor U3275 (N_3275,N_2961,N_2356);
and U3276 (N_3276,N_2518,N_2432);
xor U3277 (N_3277,N_2897,N_2835);
or U3278 (N_3278,N_2345,N_2472);
or U3279 (N_3279,N_2648,N_2934);
and U3280 (N_3280,N_2265,N_2928);
nor U3281 (N_3281,N_2441,N_2352);
and U3282 (N_3282,N_2210,N_2595);
nor U3283 (N_3283,N_2580,N_2628);
nor U3284 (N_3284,N_2719,N_2289);
and U3285 (N_3285,N_2350,N_2376);
xnor U3286 (N_3286,N_2499,N_2064);
and U3287 (N_3287,N_2599,N_2532);
and U3288 (N_3288,N_2712,N_2501);
or U3289 (N_3289,N_2937,N_2152);
nand U3290 (N_3290,N_2065,N_2264);
xnor U3291 (N_3291,N_2436,N_2809);
nor U3292 (N_3292,N_2362,N_2244);
and U3293 (N_3293,N_2492,N_2372);
nand U3294 (N_3294,N_2309,N_2861);
nor U3295 (N_3295,N_2081,N_2504);
nor U3296 (N_3296,N_2262,N_2784);
or U3297 (N_3297,N_2316,N_2705);
nor U3298 (N_3298,N_2940,N_2034);
nor U3299 (N_3299,N_2438,N_2866);
xnor U3300 (N_3300,N_2679,N_2273);
nand U3301 (N_3301,N_2883,N_2333);
nor U3302 (N_3302,N_2975,N_2678);
nor U3303 (N_3303,N_2559,N_2626);
and U3304 (N_3304,N_2077,N_2535);
nor U3305 (N_3305,N_2257,N_2723);
or U3306 (N_3306,N_2733,N_2400);
xnor U3307 (N_3307,N_2846,N_2956);
or U3308 (N_3308,N_2808,N_2295);
nand U3309 (N_3309,N_2663,N_2130);
nor U3310 (N_3310,N_2253,N_2175);
and U3311 (N_3311,N_2404,N_2847);
or U3312 (N_3312,N_2102,N_2839);
nor U3313 (N_3313,N_2227,N_2248);
xnor U3314 (N_3314,N_2969,N_2000);
and U3315 (N_3315,N_2619,N_2547);
and U3316 (N_3316,N_2029,N_2243);
or U3317 (N_3317,N_2087,N_2165);
nor U3318 (N_3318,N_2434,N_2878);
and U3319 (N_3319,N_2718,N_2405);
and U3320 (N_3320,N_2115,N_2018);
and U3321 (N_3321,N_2681,N_2026);
and U3322 (N_3322,N_2957,N_2025);
or U3323 (N_3323,N_2997,N_2921);
or U3324 (N_3324,N_2391,N_2579);
nand U3325 (N_3325,N_2630,N_2807);
nand U3326 (N_3326,N_2079,N_2374);
nand U3327 (N_3327,N_2250,N_2002);
nor U3328 (N_3328,N_2437,N_2056);
nor U3329 (N_3329,N_2031,N_2101);
xnor U3330 (N_3330,N_2713,N_2074);
xnor U3331 (N_3331,N_2804,N_2470);
nor U3332 (N_3332,N_2443,N_2040);
and U3333 (N_3333,N_2687,N_2095);
xor U3334 (N_3334,N_2801,N_2798);
xor U3335 (N_3335,N_2070,N_2959);
or U3336 (N_3336,N_2484,N_2788);
nor U3337 (N_3337,N_2028,N_2304);
nand U3338 (N_3338,N_2609,N_2460);
nand U3339 (N_3339,N_2770,N_2526);
or U3340 (N_3340,N_2351,N_2702);
xnor U3341 (N_3341,N_2855,N_2533);
or U3342 (N_3342,N_2690,N_2999);
nand U3343 (N_3343,N_2669,N_2783);
nand U3344 (N_3344,N_2134,N_2148);
or U3345 (N_3345,N_2608,N_2508);
nor U3346 (N_3346,N_2063,N_2943);
nand U3347 (N_3347,N_2989,N_2692);
and U3348 (N_3348,N_2837,N_2893);
nand U3349 (N_3349,N_2754,N_2780);
nor U3350 (N_3350,N_2060,N_2875);
and U3351 (N_3351,N_2498,N_2971);
nand U3352 (N_3352,N_2313,N_2994);
nand U3353 (N_3353,N_2139,N_2734);
nand U3354 (N_3354,N_2341,N_2667);
and U3355 (N_3355,N_2512,N_2693);
nor U3356 (N_3356,N_2636,N_2008);
and U3357 (N_3357,N_2486,N_2640);
and U3358 (N_3358,N_2843,N_2310);
or U3359 (N_3359,N_2193,N_2722);
xnor U3360 (N_3360,N_2565,N_2036);
nand U3361 (N_3361,N_2899,N_2604);
nand U3362 (N_3362,N_2750,N_2315);
and U3363 (N_3363,N_2684,N_2927);
and U3364 (N_3364,N_2427,N_2390);
nor U3365 (N_3365,N_2830,N_2842);
and U3366 (N_3366,N_2661,N_2477);
nand U3367 (N_3367,N_2386,N_2918);
nor U3368 (N_3368,N_2818,N_2353);
and U3369 (N_3369,N_2912,N_2037);
nor U3370 (N_3370,N_2450,N_2321);
nor U3371 (N_3371,N_2877,N_2084);
xnor U3372 (N_3372,N_2094,N_2941);
or U3373 (N_3373,N_2803,N_2297);
or U3374 (N_3374,N_2027,N_2720);
nand U3375 (N_3375,N_2614,N_2267);
or U3376 (N_3376,N_2515,N_2462);
xnor U3377 (N_3377,N_2824,N_2410);
and U3378 (N_3378,N_2371,N_2355);
nor U3379 (N_3379,N_2639,N_2030);
or U3380 (N_3380,N_2772,N_2756);
and U3381 (N_3381,N_2548,N_2647);
and U3382 (N_3382,N_2020,N_2487);
nor U3383 (N_3383,N_2841,N_2170);
xnor U3384 (N_3384,N_2236,N_2256);
xnor U3385 (N_3385,N_2976,N_2232);
nor U3386 (N_3386,N_2699,N_2120);
or U3387 (N_3387,N_2409,N_2401);
nand U3388 (N_3388,N_2480,N_2836);
nor U3389 (N_3389,N_2083,N_2597);
nand U3390 (N_3390,N_2665,N_2823);
nor U3391 (N_3391,N_2086,N_2050);
nand U3392 (N_3392,N_2276,N_2342);
xor U3393 (N_3393,N_2519,N_2381);
nor U3394 (N_3394,N_2715,N_2123);
nand U3395 (N_3395,N_2523,N_2726);
xnor U3396 (N_3396,N_2220,N_2838);
and U3397 (N_3397,N_2863,N_2128);
xor U3398 (N_3398,N_2834,N_2950);
nor U3399 (N_3399,N_2235,N_2500);
xnor U3400 (N_3400,N_2932,N_2104);
nand U3401 (N_3401,N_2534,N_2164);
nor U3402 (N_3402,N_2490,N_2435);
or U3403 (N_3403,N_2379,N_2664);
nor U3404 (N_3404,N_2088,N_2261);
and U3405 (N_3405,N_2729,N_2581);
and U3406 (N_3406,N_2013,N_2766);
nand U3407 (N_3407,N_2141,N_2670);
nand U3408 (N_3408,N_2497,N_2571);
and U3409 (N_3409,N_2953,N_2144);
nand U3410 (N_3410,N_2973,N_2076);
or U3411 (N_3411,N_2172,N_2459);
nand U3412 (N_3412,N_2071,N_2047);
and U3413 (N_3413,N_2252,N_2759);
xor U3414 (N_3414,N_2213,N_2566);
or U3415 (N_3415,N_2993,N_2822);
or U3416 (N_3416,N_2249,N_2817);
and U3417 (N_3417,N_2491,N_2627);
xor U3418 (N_3418,N_2760,N_2922);
nand U3419 (N_3419,N_2214,N_2167);
and U3420 (N_3420,N_2464,N_2021);
or U3421 (N_3421,N_2833,N_2496);
xor U3422 (N_3422,N_2507,N_2287);
and U3423 (N_3423,N_2903,N_2332);
nor U3424 (N_3424,N_2536,N_2996);
nor U3425 (N_3425,N_2777,N_2951);
nand U3426 (N_3426,N_2091,N_2440);
xor U3427 (N_3427,N_2284,N_2397);
and U3428 (N_3428,N_2761,N_2725);
nor U3429 (N_3429,N_2312,N_2217);
nor U3430 (N_3430,N_2347,N_2931);
or U3431 (N_3431,N_2864,N_2402);
or U3432 (N_3432,N_2977,N_2191);
and U3433 (N_3433,N_2113,N_2431);
and U3434 (N_3434,N_2862,N_2151);
nand U3435 (N_3435,N_2411,N_2421);
nor U3436 (N_3436,N_2905,N_2108);
nor U3437 (N_3437,N_2981,N_2270);
nor U3438 (N_3438,N_2185,N_2334);
nor U3439 (N_3439,N_2388,N_2696);
or U3440 (N_3440,N_2119,N_2493);
and U3441 (N_3441,N_2444,N_2045);
nor U3442 (N_3442,N_2657,N_2327);
xnor U3443 (N_3443,N_2448,N_2365);
nand U3444 (N_3444,N_2452,N_2992);
or U3445 (N_3445,N_2299,N_2884);
nand U3446 (N_3446,N_2488,N_2416);
xnor U3447 (N_3447,N_2970,N_2944);
nor U3448 (N_3448,N_2787,N_2600);
and U3449 (N_3449,N_2461,N_2182);
and U3450 (N_3450,N_2143,N_2125);
xor U3451 (N_3451,N_2322,N_2731);
nand U3452 (N_3452,N_2522,N_2919);
xor U3453 (N_3453,N_2908,N_2936);
nand U3454 (N_3454,N_2009,N_2503);
and U3455 (N_3455,N_2540,N_2012);
xnor U3456 (N_3456,N_2337,N_2871);
or U3457 (N_3457,N_2635,N_2300);
or U3458 (N_3458,N_2156,N_2881);
nand U3459 (N_3459,N_2473,N_2615);
and U3460 (N_3460,N_2570,N_2001);
xor U3461 (N_3461,N_2998,N_2727);
nand U3462 (N_3462,N_2245,N_2525);
nor U3463 (N_3463,N_2890,N_2349);
nand U3464 (N_3464,N_2378,N_2068);
nor U3465 (N_3465,N_2553,N_2796);
and U3466 (N_3466,N_2228,N_2066);
xnor U3467 (N_3467,N_2479,N_2549);
and U3468 (N_3468,N_2041,N_2246);
nor U3469 (N_3469,N_2199,N_2344);
nor U3470 (N_3470,N_2816,N_2279);
and U3471 (N_3471,N_2876,N_2575);
nand U3472 (N_3472,N_2537,N_2576);
and U3473 (N_3473,N_2011,N_2183);
nand U3474 (N_3474,N_2468,N_2509);
nor U3475 (N_3475,N_2942,N_2949);
xor U3476 (N_3476,N_2301,N_2716);
and U3477 (N_3477,N_2545,N_2133);
or U3478 (N_3478,N_2073,N_2129);
nor U3479 (N_3479,N_2035,N_2135);
xnor U3480 (N_3480,N_2126,N_2538);
xor U3481 (N_3481,N_2366,N_2208);
nand U3482 (N_3482,N_2527,N_2373);
and U3483 (N_3483,N_2275,N_2680);
and U3484 (N_3484,N_2204,N_2662);
and U3485 (N_3485,N_2424,N_2710);
xnor U3486 (N_3486,N_2601,N_2061);
or U3487 (N_3487,N_2767,N_2200);
and U3488 (N_3488,N_2771,N_2984);
xnor U3489 (N_3489,N_2359,N_2641);
xor U3490 (N_3490,N_2370,N_2286);
or U3491 (N_3491,N_2184,N_2420);
nor U3492 (N_3492,N_2857,N_2278);
xor U3493 (N_3493,N_2653,N_2430);
and U3494 (N_3494,N_2676,N_2212);
nand U3495 (N_3495,N_2814,N_2845);
nor U3496 (N_3496,N_2360,N_2447);
and U3497 (N_3497,N_2363,N_2539);
nand U3498 (N_3498,N_2174,N_2511);
nand U3499 (N_3499,N_2032,N_2053);
or U3500 (N_3500,N_2293,N_2309);
nand U3501 (N_3501,N_2274,N_2353);
xnor U3502 (N_3502,N_2967,N_2024);
xnor U3503 (N_3503,N_2573,N_2936);
xnor U3504 (N_3504,N_2017,N_2477);
and U3505 (N_3505,N_2588,N_2605);
and U3506 (N_3506,N_2517,N_2827);
and U3507 (N_3507,N_2939,N_2091);
xnor U3508 (N_3508,N_2842,N_2677);
nand U3509 (N_3509,N_2771,N_2621);
or U3510 (N_3510,N_2298,N_2672);
and U3511 (N_3511,N_2988,N_2385);
nand U3512 (N_3512,N_2176,N_2734);
nand U3513 (N_3513,N_2132,N_2053);
nand U3514 (N_3514,N_2714,N_2064);
nand U3515 (N_3515,N_2732,N_2064);
or U3516 (N_3516,N_2769,N_2301);
nand U3517 (N_3517,N_2378,N_2025);
xnor U3518 (N_3518,N_2390,N_2041);
and U3519 (N_3519,N_2738,N_2987);
and U3520 (N_3520,N_2157,N_2646);
nand U3521 (N_3521,N_2479,N_2147);
or U3522 (N_3522,N_2704,N_2101);
or U3523 (N_3523,N_2635,N_2813);
or U3524 (N_3524,N_2359,N_2031);
nand U3525 (N_3525,N_2291,N_2717);
nand U3526 (N_3526,N_2146,N_2187);
nor U3527 (N_3527,N_2723,N_2851);
xnor U3528 (N_3528,N_2863,N_2557);
or U3529 (N_3529,N_2510,N_2514);
nand U3530 (N_3530,N_2337,N_2016);
or U3531 (N_3531,N_2366,N_2825);
or U3532 (N_3532,N_2291,N_2067);
or U3533 (N_3533,N_2569,N_2918);
or U3534 (N_3534,N_2648,N_2921);
nor U3535 (N_3535,N_2108,N_2045);
xnor U3536 (N_3536,N_2658,N_2390);
xor U3537 (N_3537,N_2250,N_2942);
or U3538 (N_3538,N_2852,N_2003);
and U3539 (N_3539,N_2095,N_2412);
nand U3540 (N_3540,N_2998,N_2808);
and U3541 (N_3541,N_2677,N_2065);
and U3542 (N_3542,N_2152,N_2650);
nand U3543 (N_3543,N_2207,N_2536);
nand U3544 (N_3544,N_2632,N_2220);
xnor U3545 (N_3545,N_2633,N_2618);
xnor U3546 (N_3546,N_2155,N_2064);
nand U3547 (N_3547,N_2893,N_2189);
xor U3548 (N_3548,N_2771,N_2160);
xor U3549 (N_3549,N_2871,N_2780);
and U3550 (N_3550,N_2907,N_2915);
and U3551 (N_3551,N_2673,N_2452);
nor U3552 (N_3552,N_2231,N_2084);
nor U3553 (N_3553,N_2094,N_2945);
xor U3554 (N_3554,N_2540,N_2737);
xor U3555 (N_3555,N_2563,N_2771);
nor U3556 (N_3556,N_2001,N_2410);
nand U3557 (N_3557,N_2306,N_2599);
xor U3558 (N_3558,N_2274,N_2778);
nor U3559 (N_3559,N_2424,N_2196);
nor U3560 (N_3560,N_2175,N_2542);
nor U3561 (N_3561,N_2375,N_2343);
and U3562 (N_3562,N_2526,N_2772);
xor U3563 (N_3563,N_2965,N_2804);
nand U3564 (N_3564,N_2571,N_2514);
and U3565 (N_3565,N_2322,N_2937);
or U3566 (N_3566,N_2089,N_2712);
nor U3567 (N_3567,N_2217,N_2714);
and U3568 (N_3568,N_2803,N_2656);
and U3569 (N_3569,N_2614,N_2208);
xnor U3570 (N_3570,N_2904,N_2284);
nand U3571 (N_3571,N_2111,N_2504);
xnor U3572 (N_3572,N_2526,N_2769);
nor U3573 (N_3573,N_2582,N_2796);
xor U3574 (N_3574,N_2378,N_2562);
and U3575 (N_3575,N_2692,N_2797);
or U3576 (N_3576,N_2824,N_2244);
and U3577 (N_3577,N_2956,N_2977);
nand U3578 (N_3578,N_2450,N_2114);
or U3579 (N_3579,N_2776,N_2223);
nor U3580 (N_3580,N_2566,N_2541);
and U3581 (N_3581,N_2768,N_2886);
nand U3582 (N_3582,N_2794,N_2670);
or U3583 (N_3583,N_2666,N_2987);
nor U3584 (N_3584,N_2428,N_2043);
nand U3585 (N_3585,N_2883,N_2084);
or U3586 (N_3586,N_2149,N_2822);
and U3587 (N_3587,N_2088,N_2428);
xor U3588 (N_3588,N_2111,N_2011);
or U3589 (N_3589,N_2767,N_2280);
and U3590 (N_3590,N_2280,N_2190);
nor U3591 (N_3591,N_2982,N_2266);
or U3592 (N_3592,N_2486,N_2279);
or U3593 (N_3593,N_2810,N_2775);
and U3594 (N_3594,N_2644,N_2520);
nor U3595 (N_3595,N_2393,N_2029);
nand U3596 (N_3596,N_2506,N_2976);
xor U3597 (N_3597,N_2660,N_2945);
xnor U3598 (N_3598,N_2113,N_2905);
and U3599 (N_3599,N_2132,N_2407);
xor U3600 (N_3600,N_2951,N_2470);
or U3601 (N_3601,N_2827,N_2602);
nand U3602 (N_3602,N_2530,N_2823);
nand U3603 (N_3603,N_2125,N_2298);
or U3604 (N_3604,N_2631,N_2420);
xnor U3605 (N_3605,N_2138,N_2878);
or U3606 (N_3606,N_2630,N_2223);
nor U3607 (N_3607,N_2329,N_2741);
or U3608 (N_3608,N_2207,N_2584);
or U3609 (N_3609,N_2116,N_2201);
xnor U3610 (N_3610,N_2915,N_2701);
and U3611 (N_3611,N_2507,N_2774);
or U3612 (N_3612,N_2054,N_2311);
nand U3613 (N_3613,N_2966,N_2961);
nor U3614 (N_3614,N_2727,N_2571);
xor U3615 (N_3615,N_2715,N_2142);
or U3616 (N_3616,N_2470,N_2011);
and U3617 (N_3617,N_2787,N_2882);
nor U3618 (N_3618,N_2517,N_2592);
and U3619 (N_3619,N_2704,N_2142);
nor U3620 (N_3620,N_2268,N_2042);
nand U3621 (N_3621,N_2506,N_2459);
nor U3622 (N_3622,N_2167,N_2679);
nor U3623 (N_3623,N_2805,N_2544);
xnor U3624 (N_3624,N_2141,N_2677);
nor U3625 (N_3625,N_2094,N_2595);
or U3626 (N_3626,N_2880,N_2098);
nand U3627 (N_3627,N_2238,N_2613);
xor U3628 (N_3628,N_2113,N_2859);
and U3629 (N_3629,N_2712,N_2122);
or U3630 (N_3630,N_2136,N_2402);
nor U3631 (N_3631,N_2078,N_2245);
nor U3632 (N_3632,N_2411,N_2423);
or U3633 (N_3633,N_2747,N_2222);
nand U3634 (N_3634,N_2346,N_2380);
xor U3635 (N_3635,N_2763,N_2849);
nor U3636 (N_3636,N_2035,N_2159);
xnor U3637 (N_3637,N_2618,N_2482);
xnor U3638 (N_3638,N_2361,N_2957);
or U3639 (N_3639,N_2579,N_2838);
nand U3640 (N_3640,N_2274,N_2055);
nor U3641 (N_3641,N_2745,N_2121);
or U3642 (N_3642,N_2729,N_2580);
and U3643 (N_3643,N_2476,N_2109);
nand U3644 (N_3644,N_2594,N_2531);
and U3645 (N_3645,N_2657,N_2237);
xor U3646 (N_3646,N_2022,N_2794);
or U3647 (N_3647,N_2415,N_2703);
or U3648 (N_3648,N_2590,N_2182);
nor U3649 (N_3649,N_2059,N_2686);
nand U3650 (N_3650,N_2085,N_2771);
xor U3651 (N_3651,N_2283,N_2874);
xnor U3652 (N_3652,N_2315,N_2900);
nand U3653 (N_3653,N_2453,N_2801);
or U3654 (N_3654,N_2761,N_2964);
nor U3655 (N_3655,N_2644,N_2289);
nor U3656 (N_3656,N_2491,N_2192);
nand U3657 (N_3657,N_2935,N_2930);
nor U3658 (N_3658,N_2132,N_2139);
and U3659 (N_3659,N_2252,N_2268);
and U3660 (N_3660,N_2568,N_2507);
nand U3661 (N_3661,N_2676,N_2369);
or U3662 (N_3662,N_2127,N_2300);
or U3663 (N_3663,N_2761,N_2013);
and U3664 (N_3664,N_2650,N_2506);
xor U3665 (N_3665,N_2511,N_2918);
nor U3666 (N_3666,N_2910,N_2720);
xnor U3667 (N_3667,N_2837,N_2043);
and U3668 (N_3668,N_2553,N_2033);
xnor U3669 (N_3669,N_2489,N_2116);
and U3670 (N_3670,N_2066,N_2328);
or U3671 (N_3671,N_2057,N_2376);
xor U3672 (N_3672,N_2538,N_2961);
nand U3673 (N_3673,N_2133,N_2526);
and U3674 (N_3674,N_2971,N_2993);
xnor U3675 (N_3675,N_2431,N_2412);
xnor U3676 (N_3676,N_2486,N_2416);
nand U3677 (N_3677,N_2427,N_2029);
and U3678 (N_3678,N_2815,N_2166);
nand U3679 (N_3679,N_2261,N_2958);
xor U3680 (N_3680,N_2625,N_2637);
nor U3681 (N_3681,N_2946,N_2148);
nor U3682 (N_3682,N_2338,N_2940);
and U3683 (N_3683,N_2148,N_2350);
or U3684 (N_3684,N_2403,N_2143);
nand U3685 (N_3685,N_2611,N_2797);
nor U3686 (N_3686,N_2840,N_2967);
nor U3687 (N_3687,N_2286,N_2907);
and U3688 (N_3688,N_2250,N_2487);
xor U3689 (N_3689,N_2259,N_2034);
and U3690 (N_3690,N_2277,N_2791);
nand U3691 (N_3691,N_2384,N_2443);
or U3692 (N_3692,N_2297,N_2458);
xnor U3693 (N_3693,N_2938,N_2441);
xor U3694 (N_3694,N_2961,N_2337);
or U3695 (N_3695,N_2036,N_2360);
xor U3696 (N_3696,N_2290,N_2308);
xnor U3697 (N_3697,N_2079,N_2486);
nand U3698 (N_3698,N_2353,N_2325);
xnor U3699 (N_3699,N_2713,N_2337);
xnor U3700 (N_3700,N_2633,N_2307);
or U3701 (N_3701,N_2196,N_2011);
nor U3702 (N_3702,N_2255,N_2797);
xor U3703 (N_3703,N_2069,N_2244);
or U3704 (N_3704,N_2750,N_2580);
nand U3705 (N_3705,N_2921,N_2890);
or U3706 (N_3706,N_2144,N_2358);
xnor U3707 (N_3707,N_2137,N_2561);
and U3708 (N_3708,N_2935,N_2188);
and U3709 (N_3709,N_2808,N_2674);
xnor U3710 (N_3710,N_2354,N_2897);
xnor U3711 (N_3711,N_2412,N_2486);
nand U3712 (N_3712,N_2171,N_2855);
nand U3713 (N_3713,N_2795,N_2494);
or U3714 (N_3714,N_2447,N_2568);
or U3715 (N_3715,N_2699,N_2790);
nor U3716 (N_3716,N_2536,N_2085);
nor U3717 (N_3717,N_2167,N_2432);
and U3718 (N_3718,N_2592,N_2974);
or U3719 (N_3719,N_2409,N_2317);
xnor U3720 (N_3720,N_2622,N_2749);
nor U3721 (N_3721,N_2250,N_2235);
nor U3722 (N_3722,N_2595,N_2543);
or U3723 (N_3723,N_2758,N_2345);
or U3724 (N_3724,N_2870,N_2203);
xor U3725 (N_3725,N_2302,N_2700);
xor U3726 (N_3726,N_2157,N_2774);
nor U3727 (N_3727,N_2032,N_2831);
and U3728 (N_3728,N_2939,N_2844);
nand U3729 (N_3729,N_2480,N_2131);
xor U3730 (N_3730,N_2629,N_2944);
nand U3731 (N_3731,N_2659,N_2559);
or U3732 (N_3732,N_2460,N_2748);
and U3733 (N_3733,N_2446,N_2801);
and U3734 (N_3734,N_2013,N_2783);
xnor U3735 (N_3735,N_2378,N_2377);
nor U3736 (N_3736,N_2963,N_2482);
xor U3737 (N_3737,N_2887,N_2220);
nand U3738 (N_3738,N_2591,N_2544);
nand U3739 (N_3739,N_2584,N_2152);
nor U3740 (N_3740,N_2543,N_2658);
or U3741 (N_3741,N_2748,N_2589);
nor U3742 (N_3742,N_2471,N_2127);
nand U3743 (N_3743,N_2882,N_2085);
xor U3744 (N_3744,N_2051,N_2397);
and U3745 (N_3745,N_2178,N_2388);
nand U3746 (N_3746,N_2222,N_2724);
and U3747 (N_3747,N_2107,N_2279);
and U3748 (N_3748,N_2740,N_2721);
and U3749 (N_3749,N_2777,N_2514);
nor U3750 (N_3750,N_2667,N_2157);
nor U3751 (N_3751,N_2606,N_2981);
nor U3752 (N_3752,N_2875,N_2779);
nor U3753 (N_3753,N_2407,N_2720);
or U3754 (N_3754,N_2764,N_2663);
nor U3755 (N_3755,N_2137,N_2882);
nand U3756 (N_3756,N_2111,N_2331);
nand U3757 (N_3757,N_2323,N_2514);
or U3758 (N_3758,N_2073,N_2734);
or U3759 (N_3759,N_2800,N_2581);
nand U3760 (N_3760,N_2009,N_2895);
or U3761 (N_3761,N_2009,N_2491);
xnor U3762 (N_3762,N_2023,N_2586);
nand U3763 (N_3763,N_2234,N_2777);
nand U3764 (N_3764,N_2051,N_2019);
or U3765 (N_3765,N_2317,N_2430);
nand U3766 (N_3766,N_2451,N_2486);
and U3767 (N_3767,N_2948,N_2851);
xnor U3768 (N_3768,N_2180,N_2337);
nand U3769 (N_3769,N_2069,N_2631);
and U3770 (N_3770,N_2708,N_2083);
or U3771 (N_3771,N_2432,N_2065);
nor U3772 (N_3772,N_2680,N_2300);
or U3773 (N_3773,N_2195,N_2299);
nand U3774 (N_3774,N_2084,N_2403);
nor U3775 (N_3775,N_2406,N_2034);
nand U3776 (N_3776,N_2320,N_2730);
and U3777 (N_3777,N_2217,N_2735);
nor U3778 (N_3778,N_2819,N_2367);
xnor U3779 (N_3779,N_2937,N_2713);
and U3780 (N_3780,N_2379,N_2729);
xnor U3781 (N_3781,N_2578,N_2699);
and U3782 (N_3782,N_2201,N_2703);
nand U3783 (N_3783,N_2924,N_2160);
or U3784 (N_3784,N_2283,N_2350);
xor U3785 (N_3785,N_2824,N_2760);
or U3786 (N_3786,N_2611,N_2214);
nor U3787 (N_3787,N_2460,N_2286);
and U3788 (N_3788,N_2276,N_2460);
xor U3789 (N_3789,N_2424,N_2571);
xnor U3790 (N_3790,N_2241,N_2142);
and U3791 (N_3791,N_2744,N_2528);
nor U3792 (N_3792,N_2165,N_2011);
or U3793 (N_3793,N_2634,N_2380);
or U3794 (N_3794,N_2093,N_2939);
or U3795 (N_3795,N_2287,N_2518);
xor U3796 (N_3796,N_2772,N_2056);
and U3797 (N_3797,N_2825,N_2336);
nand U3798 (N_3798,N_2002,N_2502);
nand U3799 (N_3799,N_2430,N_2539);
and U3800 (N_3800,N_2253,N_2070);
and U3801 (N_3801,N_2996,N_2883);
and U3802 (N_3802,N_2908,N_2632);
and U3803 (N_3803,N_2405,N_2666);
nor U3804 (N_3804,N_2786,N_2075);
or U3805 (N_3805,N_2071,N_2462);
and U3806 (N_3806,N_2424,N_2499);
and U3807 (N_3807,N_2263,N_2257);
or U3808 (N_3808,N_2694,N_2674);
or U3809 (N_3809,N_2486,N_2995);
xnor U3810 (N_3810,N_2217,N_2812);
and U3811 (N_3811,N_2711,N_2796);
or U3812 (N_3812,N_2505,N_2109);
xor U3813 (N_3813,N_2108,N_2333);
xnor U3814 (N_3814,N_2107,N_2227);
nand U3815 (N_3815,N_2984,N_2369);
or U3816 (N_3816,N_2532,N_2682);
or U3817 (N_3817,N_2681,N_2705);
nand U3818 (N_3818,N_2789,N_2386);
or U3819 (N_3819,N_2299,N_2559);
or U3820 (N_3820,N_2545,N_2661);
nand U3821 (N_3821,N_2260,N_2499);
xor U3822 (N_3822,N_2264,N_2974);
nor U3823 (N_3823,N_2359,N_2006);
and U3824 (N_3824,N_2165,N_2817);
nand U3825 (N_3825,N_2580,N_2537);
xnor U3826 (N_3826,N_2178,N_2998);
nand U3827 (N_3827,N_2518,N_2895);
and U3828 (N_3828,N_2647,N_2504);
or U3829 (N_3829,N_2566,N_2496);
or U3830 (N_3830,N_2892,N_2160);
nor U3831 (N_3831,N_2450,N_2043);
and U3832 (N_3832,N_2783,N_2758);
and U3833 (N_3833,N_2520,N_2484);
xor U3834 (N_3834,N_2831,N_2859);
xnor U3835 (N_3835,N_2077,N_2277);
nor U3836 (N_3836,N_2893,N_2635);
nand U3837 (N_3837,N_2494,N_2655);
xor U3838 (N_3838,N_2994,N_2065);
nand U3839 (N_3839,N_2958,N_2280);
xnor U3840 (N_3840,N_2522,N_2966);
nand U3841 (N_3841,N_2865,N_2278);
nand U3842 (N_3842,N_2534,N_2513);
xor U3843 (N_3843,N_2569,N_2017);
and U3844 (N_3844,N_2411,N_2970);
or U3845 (N_3845,N_2781,N_2334);
nor U3846 (N_3846,N_2163,N_2702);
and U3847 (N_3847,N_2406,N_2771);
nand U3848 (N_3848,N_2247,N_2398);
nor U3849 (N_3849,N_2317,N_2931);
and U3850 (N_3850,N_2137,N_2206);
nor U3851 (N_3851,N_2310,N_2134);
nor U3852 (N_3852,N_2630,N_2804);
nand U3853 (N_3853,N_2660,N_2520);
nand U3854 (N_3854,N_2914,N_2615);
nand U3855 (N_3855,N_2111,N_2949);
nor U3856 (N_3856,N_2804,N_2638);
nor U3857 (N_3857,N_2842,N_2144);
nor U3858 (N_3858,N_2986,N_2749);
and U3859 (N_3859,N_2066,N_2651);
nand U3860 (N_3860,N_2372,N_2466);
nor U3861 (N_3861,N_2976,N_2310);
and U3862 (N_3862,N_2903,N_2924);
xnor U3863 (N_3863,N_2304,N_2327);
or U3864 (N_3864,N_2430,N_2884);
nor U3865 (N_3865,N_2890,N_2624);
nand U3866 (N_3866,N_2498,N_2098);
nor U3867 (N_3867,N_2417,N_2888);
and U3868 (N_3868,N_2159,N_2122);
xnor U3869 (N_3869,N_2287,N_2442);
nand U3870 (N_3870,N_2285,N_2844);
nand U3871 (N_3871,N_2707,N_2575);
and U3872 (N_3872,N_2481,N_2797);
or U3873 (N_3873,N_2045,N_2104);
nand U3874 (N_3874,N_2467,N_2095);
xnor U3875 (N_3875,N_2609,N_2254);
xnor U3876 (N_3876,N_2893,N_2871);
or U3877 (N_3877,N_2655,N_2698);
nand U3878 (N_3878,N_2974,N_2230);
nor U3879 (N_3879,N_2320,N_2169);
nand U3880 (N_3880,N_2233,N_2848);
nor U3881 (N_3881,N_2859,N_2038);
xnor U3882 (N_3882,N_2341,N_2494);
nor U3883 (N_3883,N_2912,N_2334);
nand U3884 (N_3884,N_2379,N_2061);
or U3885 (N_3885,N_2043,N_2545);
or U3886 (N_3886,N_2362,N_2956);
nor U3887 (N_3887,N_2122,N_2205);
and U3888 (N_3888,N_2383,N_2794);
nand U3889 (N_3889,N_2671,N_2621);
or U3890 (N_3890,N_2685,N_2351);
nor U3891 (N_3891,N_2609,N_2927);
nand U3892 (N_3892,N_2941,N_2360);
nor U3893 (N_3893,N_2017,N_2914);
or U3894 (N_3894,N_2984,N_2918);
and U3895 (N_3895,N_2604,N_2885);
or U3896 (N_3896,N_2373,N_2544);
or U3897 (N_3897,N_2603,N_2914);
or U3898 (N_3898,N_2696,N_2950);
nand U3899 (N_3899,N_2794,N_2172);
or U3900 (N_3900,N_2626,N_2740);
or U3901 (N_3901,N_2601,N_2387);
or U3902 (N_3902,N_2823,N_2662);
nor U3903 (N_3903,N_2000,N_2001);
nand U3904 (N_3904,N_2753,N_2149);
nand U3905 (N_3905,N_2342,N_2302);
nor U3906 (N_3906,N_2276,N_2103);
nand U3907 (N_3907,N_2984,N_2777);
or U3908 (N_3908,N_2960,N_2388);
nand U3909 (N_3909,N_2479,N_2624);
or U3910 (N_3910,N_2579,N_2661);
and U3911 (N_3911,N_2236,N_2890);
or U3912 (N_3912,N_2228,N_2790);
xor U3913 (N_3913,N_2483,N_2303);
nor U3914 (N_3914,N_2513,N_2520);
xor U3915 (N_3915,N_2244,N_2874);
and U3916 (N_3916,N_2427,N_2740);
xnor U3917 (N_3917,N_2704,N_2053);
nor U3918 (N_3918,N_2966,N_2319);
nand U3919 (N_3919,N_2836,N_2966);
and U3920 (N_3920,N_2867,N_2389);
and U3921 (N_3921,N_2085,N_2401);
and U3922 (N_3922,N_2434,N_2324);
and U3923 (N_3923,N_2828,N_2940);
or U3924 (N_3924,N_2830,N_2368);
and U3925 (N_3925,N_2307,N_2773);
or U3926 (N_3926,N_2178,N_2980);
and U3927 (N_3927,N_2499,N_2452);
nand U3928 (N_3928,N_2450,N_2276);
xor U3929 (N_3929,N_2588,N_2317);
nor U3930 (N_3930,N_2732,N_2275);
and U3931 (N_3931,N_2900,N_2971);
nand U3932 (N_3932,N_2872,N_2136);
xor U3933 (N_3933,N_2824,N_2937);
or U3934 (N_3934,N_2721,N_2689);
nor U3935 (N_3935,N_2218,N_2326);
nand U3936 (N_3936,N_2297,N_2165);
xor U3937 (N_3937,N_2023,N_2452);
nor U3938 (N_3938,N_2096,N_2235);
xnor U3939 (N_3939,N_2921,N_2195);
nand U3940 (N_3940,N_2231,N_2425);
nand U3941 (N_3941,N_2231,N_2141);
xor U3942 (N_3942,N_2126,N_2897);
nor U3943 (N_3943,N_2144,N_2412);
xor U3944 (N_3944,N_2067,N_2795);
nand U3945 (N_3945,N_2655,N_2540);
or U3946 (N_3946,N_2568,N_2254);
or U3947 (N_3947,N_2521,N_2349);
and U3948 (N_3948,N_2078,N_2876);
nand U3949 (N_3949,N_2111,N_2805);
nor U3950 (N_3950,N_2215,N_2024);
and U3951 (N_3951,N_2325,N_2760);
or U3952 (N_3952,N_2257,N_2105);
nand U3953 (N_3953,N_2943,N_2725);
and U3954 (N_3954,N_2294,N_2058);
or U3955 (N_3955,N_2978,N_2738);
nor U3956 (N_3956,N_2018,N_2430);
and U3957 (N_3957,N_2064,N_2834);
xnor U3958 (N_3958,N_2865,N_2731);
xor U3959 (N_3959,N_2391,N_2121);
nor U3960 (N_3960,N_2216,N_2968);
and U3961 (N_3961,N_2670,N_2776);
xor U3962 (N_3962,N_2885,N_2810);
or U3963 (N_3963,N_2328,N_2060);
nor U3964 (N_3964,N_2251,N_2772);
and U3965 (N_3965,N_2579,N_2516);
or U3966 (N_3966,N_2221,N_2095);
nand U3967 (N_3967,N_2098,N_2067);
nor U3968 (N_3968,N_2899,N_2096);
nor U3969 (N_3969,N_2896,N_2201);
nor U3970 (N_3970,N_2649,N_2977);
xor U3971 (N_3971,N_2986,N_2245);
and U3972 (N_3972,N_2705,N_2582);
or U3973 (N_3973,N_2080,N_2527);
nand U3974 (N_3974,N_2177,N_2257);
and U3975 (N_3975,N_2480,N_2443);
or U3976 (N_3976,N_2793,N_2500);
and U3977 (N_3977,N_2497,N_2549);
and U3978 (N_3978,N_2730,N_2312);
nor U3979 (N_3979,N_2598,N_2253);
and U3980 (N_3980,N_2879,N_2032);
or U3981 (N_3981,N_2404,N_2257);
nand U3982 (N_3982,N_2457,N_2692);
nor U3983 (N_3983,N_2567,N_2609);
xnor U3984 (N_3984,N_2424,N_2811);
nor U3985 (N_3985,N_2690,N_2282);
or U3986 (N_3986,N_2112,N_2610);
or U3987 (N_3987,N_2094,N_2830);
and U3988 (N_3988,N_2074,N_2732);
nor U3989 (N_3989,N_2328,N_2431);
nor U3990 (N_3990,N_2889,N_2628);
xor U3991 (N_3991,N_2232,N_2156);
nor U3992 (N_3992,N_2316,N_2466);
nand U3993 (N_3993,N_2382,N_2328);
nand U3994 (N_3994,N_2866,N_2794);
nor U3995 (N_3995,N_2622,N_2500);
nand U3996 (N_3996,N_2230,N_2902);
or U3997 (N_3997,N_2852,N_2792);
nand U3998 (N_3998,N_2177,N_2434);
and U3999 (N_3999,N_2070,N_2082);
nor U4000 (N_4000,N_3332,N_3954);
or U4001 (N_4001,N_3425,N_3681);
or U4002 (N_4002,N_3684,N_3898);
or U4003 (N_4003,N_3367,N_3643);
nor U4004 (N_4004,N_3473,N_3544);
and U4005 (N_4005,N_3509,N_3378);
nor U4006 (N_4006,N_3598,N_3104);
xnor U4007 (N_4007,N_3629,N_3686);
or U4008 (N_4008,N_3034,N_3190);
nand U4009 (N_4009,N_3679,N_3476);
or U4010 (N_4010,N_3398,N_3581);
xnor U4011 (N_4011,N_3966,N_3567);
nand U4012 (N_4012,N_3053,N_3251);
and U4013 (N_4013,N_3268,N_3244);
or U4014 (N_4014,N_3957,N_3566);
nor U4015 (N_4015,N_3380,N_3064);
nand U4016 (N_4016,N_3394,N_3140);
or U4017 (N_4017,N_3208,N_3722);
or U4018 (N_4018,N_3627,N_3225);
xnor U4019 (N_4019,N_3763,N_3186);
nor U4020 (N_4020,N_3114,N_3014);
xnor U4021 (N_4021,N_3285,N_3257);
and U4022 (N_4022,N_3060,N_3365);
or U4023 (N_4023,N_3249,N_3075);
and U4024 (N_4024,N_3716,N_3795);
or U4025 (N_4025,N_3650,N_3265);
or U4026 (N_4026,N_3870,N_3562);
xor U4027 (N_4027,N_3555,N_3608);
and U4028 (N_4028,N_3443,N_3305);
or U4029 (N_4029,N_3464,N_3557);
and U4030 (N_4030,N_3044,N_3669);
and U4031 (N_4031,N_3338,N_3712);
and U4032 (N_4032,N_3886,N_3009);
nor U4033 (N_4033,N_3573,N_3214);
nor U4034 (N_4034,N_3328,N_3692);
xnor U4035 (N_4035,N_3011,N_3304);
and U4036 (N_4036,N_3325,N_3177);
nand U4037 (N_4037,N_3522,N_3196);
or U4038 (N_4038,N_3657,N_3537);
and U4039 (N_4039,N_3729,N_3262);
or U4040 (N_4040,N_3178,N_3027);
xor U4041 (N_4041,N_3919,N_3368);
nand U4042 (N_4042,N_3575,N_3090);
nand U4043 (N_4043,N_3652,N_3023);
and U4044 (N_4044,N_3559,N_3069);
xor U4045 (N_4045,N_3970,N_3730);
and U4046 (N_4046,N_3182,N_3642);
and U4047 (N_4047,N_3995,N_3930);
and U4048 (N_4048,N_3732,N_3098);
nor U4049 (N_4049,N_3632,N_3582);
and U4050 (N_4050,N_3113,N_3740);
xnor U4051 (N_4051,N_3517,N_3736);
xnor U4052 (N_4052,N_3000,N_3396);
nor U4053 (N_4053,N_3314,N_3370);
nor U4054 (N_4054,N_3625,N_3383);
nor U4055 (N_4055,N_3040,N_3645);
and U4056 (N_4056,N_3032,N_3424);
or U4057 (N_4057,N_3761,N_3153);
or U4058 (N_4058,N_3269,N_3174);
nand U4059 (N_4059,N_3228,N_3707);
and U4060 (N_4060,N_3809,N_3323);
nor U4061 (N_4061,N_3083,N_3039);
xor U4062 (N_4062,N_3960,N_3796);
nor U4063 (N_4063,N_3733,N_3918);
and U4064 (N_4064,N_3911,N_3086);
nand U4065 (N_4065,N_3916,N_3454);
or U4066 (N_4066,N_3980,N_3242);
nand U4067 (N_4067,N_3051,N_3926);
nand U4068 (N_4068,N_3913,N_3955);
nor U4069 (N_4069,N_3709,N_3194);
or U4070 (N_4070,N_3179,N_3158);
or U4071 (N_4071,N_3151,N_3865);
nand U4072 (N_4072,N_3883,N_3601);
xor U4073 (N_4073,N_3308,N_3626);
and U4074 (N_4074,N_3620,N_3395);
xor U4075 (N_4075,N_3165,N_3436);
and U4076 (N_4076,N_3691,N_3584);
xnor U4077 (N_4077,N_3910,N_3070);
nand U4078 (N_4078,N_3611,N_3986);
nor U4079 (N_4079,N_3570,N_3175);
or U4080 (N_4080,N_3506,N_3696);
nand U4081 (N_4081,N_3357,N_3654);
nor U4082 (N_4082,N_3977,N_3416);
and U4083 (N_4083,N_3503,N_3329);
or U4084 (N_4084,N_3100,N_3591);
nor U4085 (N_4085,N_3124,N_3350);
and U4086 (N_4086,N_3539,N_3271);
or U4087 (N_4087,N_3298,N_3132);
and U4088 (N_4088,N_3699,N_3273);
nor U4089 (N_4089,N_3291,N_3264);
and U4090 (N_4090,N_3518,N_3402);
nor U4091 (N_4091,N_3355,N_3448);
nand U4092 (N_4092,N_3888,N_3203);
nand U4093 (N_4093,N_3906,N_3167);
nand U4094 (N_4094,N_3658,N_3183);
or U4095 (N_4095,N_3289,N_3659);
or U4096 (N_4096,N_3205,N_3471);
nor U4097 (N_4097,N_3318,N_3845);
nand U4098 (N_4098,N_3768,N_3337);
and U4099 (N_4099,N_3045,N_3817);
nand U4100 (N_4100,N_3411,N_3832);
xor U4101 (N_4101,N_3912,N_3997);
or U4102 (N_4102,N_3780,N_3811);
nand U4103 (N_4103,N_3420,N_3248);
and U4104 (N_4104,N_3621,N_3920);
nor U4105 (N_4105,N_3301,N_3585);
nor U4106 (N_4106,N_3335,N_3223);
or U4107 (N_4107,N_3360,N_3147);
nand U4108 (N_4108,N_3802,N_3532);
xnor U4109 (N_4109,N_3117,N_3494);
or U4110 (N_4110,N_3161,N_3874);
nand U4111 (N_4111,N_3837,N_3836);
and U4112 (N_4112,N_3879,N_3450);
xor U4113 (N_4113,N_3859,N_3036);
xnor U4114 (N_4114,N_3094,N_3030);
xnor U4115 (N_4115,N_3597,N_3530);
xor U4116 (N_4116,N_3340,N_3102);
and U4117 (N_4117,N_3202,N_3979);
xnor U4118 (N_4118,N_3789,N_3422);
or U4119 (N_4119,N_3284,N_3862);
and U4120 (N_4120,N_3680,N_3108);
and U4121 (N_4121,N_3613,N_3583);
nand U4122 (N_4122,N_3245,N_3770);
or U4123 (N_4123,N_3541,N_3666);
or U4124 (N_4124,N_3618,N_3595);
or U4125 (N_4125,N_3373,N_3737);
xor U4126 (N_4126,N_3491,N_3451);
nand U4127 (N_4127,N_3376,N_3351);
nor U4128 (N_4128,N_3118,N_3093);
xnor U4129 (N_4129,N_3745,N_3538);
and U4130 (N_4130,N_3099,N_3974);
and U4131 (N_4131,N_3333,N_3061);
nand U4132 (N_4132,N_3002,N_3753);
and U4133 (N_4133,N_3885,N_3881);
and U4134 (N_4134,N_3379,N_3587);
nand U4135 (N_4135,N_3812,N_3341);
or U4136 (N_4136,N_3472,N_3143);
and U4137 (N_4137,N_3689,N_3079);
nand U4138 (N_4138,N_3950,N_3195);
xor U4139 (N_4139,N_3279,N_3602);
and U4140 (N_4140,N_3739,N_3087);
or U4141 (N_4141,N_3460,N_3667);
or U4142 (N_4142,N_3746,N_3880);
nor U4143 (N_4143,N_3687,N_3144);
nor U4144 (N_4144,N_3330,N_3052);
nand U4145 (N_4145,N_3496,N_3864);
xnor U4146 (N_4146,N_3320,N_3369);
or U4147 (N_4147,N_3821,N_3578);
and U4148 (N_4148,N_3005,N_3944);
xnor U4149 (N_4149,N_3572,N_3071);
nand U4150 (N_4150,N_3311,N_3742);
and U4151 (N_4151,N_3478,N_3965);
or U4152 (N_4152,N_3492,N_3232);
and U4153 (N_4153,N_3825,N_3220);
or U4154 (N_4154,N_3366,N_3788);
xor U4155 (N_4155,N_3767,N_3515);
nand U4156 (N_4156,N_3731,N_3154);
nor U4157 (N_4157,N_3527,N_3142);
and U4158 (N_4158,N_3949,N_3828);
and U4159 (N_4159,N_3294,N_3551);
nor U4160 (N_4160,N_3038,N_3619);
or U4161 (N_4161,N_3839,N_3672);
nand U4162 (N_4162,N_3028,N_3967);
or U4163 (N_4163,N_3213,N_3212);
xor U4164 (N_4164,N_3306,N_3004);
and U4165 (N_4165,N_3259,N_3031);
nand U4166 (N_4166,N_3197,N_3651);
nor U4167 (N_4167,N_3495,N_3917);
nor U4168 (N_4168,N_3807,N_3711);
xnor U4169 (N_4169,N_3336,N_3590);
and U4170 (N_4170,N_3525,N_3890);
nor U4171 (N_4171,N_3393,N_3531);
nor U4172 (N_4172,N_3207,N_3412);
nor U4173 (N_4173,N_3488,N_3349);
nor U4174 (N_4174,N_3941,N_3634);
nor U4175 (N_4175,N_3637,N_3067);
or U4176 (N_4176,N_3932,N_3863);
nor U4177 (N_4177,N_3256,N_3748);
nor U4178 (N_4178,N_3106,N_3655);
xnor U4179 (N_4179,N_3033,N_3516);
and U4180 (N_4180,N_3157,N_3682);
or U4181 (N_4181,N_3484,N_3947);
and U4182 (N_4182,N_3550,N_3247);
xnor U4183 (N_4183,N_3857,N_3107);
nand U4184 (N_4184,N_3713,N_3180);
and U4185 (N_4185,N_3007,N_3814);
nor U4186 (N_4186,N_3677,N_3364);
xnor U4187 (N_4187,N_3407,N_3794);
and U4188 (N_4188,N_3047,N_3674);
xnor U4189 (N_4189,N_3465,N_3191);
or U4190 (N_4190,N_3813,N_3347);
and U4191 (N_4191,N_3635,N_3700);
nor U4192 (N_4192,N_3482,N_3925);
nand U4193 (N_4193,N_3199,N_3169);
nand U4194 (N_4194,N_3483,N_3066);
or U4195 (N_4195,N_3641,N_3111);
nor U4196 (N_4196,N_3705,N_3803);
and U4197 (N_4197,N_3101,N_3639);
and U4198 (N_4198,N_3082,N_3133);
or U4199 (N_4199,N_3410,N_3307);
nand U4200 (N_4200,N_3904,N_3384);
nor U4201 (N_4201,N_3580,N_3356);
nor U4202 (N_4202,N_3283,N_3440);
or U4203 (N_4203,N_3016,N_3694);
nand U4204 (N_4204,N_3791,N_3239);
and U4205 (N_4205,N_3022,N_3848);
or U4206 (N_4206,N_3734,N_3078);
and U4207 (N_4207,N_3948,N_3850);
xor U4208 (N_4208,N_3348,N_3263);
and U4209 (N_4209,N_3468,N_3596);
and U4210 (N_4210,N_3479,N_3240);
or U4211 (N_4211,N_3735,N_3775);
and U4212 (N_4212,N_3185,N_3827);
nand U4213 (N_4213,N_3852,N_3217);
or U4214 (N_4214,N_3467,N_3280);
xnor U4215 (N_4215,N_3564,N_3971);
or U4216 (N_4216,N_3988,N_3103);
or U4217 (N_4217,N_3149,N_3112);
nor U4218 (N_4218,N_3976,N_3310);
and U4219 (N_4219,N_3676,N_3871);
or U4220 (N_4220,N_3673,N_3431);
xnor U4221 (N_4221,N_3594,N_3293);
nor U4222 (N_4222,N_3609,N_3046);
xor U4223 (N_4223,N_3710,N_3875);
nand U4224 (N_4224,N_3838,N_3400);
nor U4225 (N_4225,N_3084,N_3276);
nor U4226 (N_4226,N_3095,N_3610);
and U4227 (N_4227,N_3354,N_3432);
nor U4228 (N_4228,N_3678,N_3893);
or U4229 (N_4229,N_3818,N_3923);
xor U4230 (N_4230,N_3612,N_3915);
and U4231 (N_4231,N_3160,N_3470);
xor U4232 (N_4232,N_3778,N_3312);
nand U4233 (N_4233,N_3670,N_3987);
xor U4234 (N_4234,N_3958,N_3545);
xor U4235 (N_4235,N_3173,N_3937);
nor U4236 (N_4236,N_3128,N_3286);
and U4237 (N_4237,N_3781,N_3092);
or U4238 (N_4238,N_3415,N_3116);
or U4239 (N_4239,N_3258,N_3556);
xor U4240 (N_4240,N_3091,N_3317);
xnor U4241 (N_4241,N_3403,N_3938);
xor U4242 (N_4242,N_3622,N_3469);
or U4243 (N_4243,N_3576,N_3757);
nand U4244 (N_4244,N_3894,N_3466);
xnor U4245 (N_4245,N_3222,N_3404);
or U4246 (N_4246,N_3392,N_3631);
and U4247 (N_4247,N_3952,N_3773);
nor U4248 (N_4248,N_3607,N_3024);
nor U4249 (N_4249,N_3990,N_3656);
nor U4250 (N_4250,N_3418,N_3524);
xnor U4251 (N_4251,N_3801,N_3513);
xnor U4252 (N_4252,N_3302,N_3640);
nor U4253 (N_4253,N_3299,N_3772);
nand U4254 (N_4254,N_3127,N_3824);
or U4255 (N_4255,N_3449,N_3633);
nand U4256 (N_4256,N_3428,N_3565);
nor U4257 (N_4257,N_3810,N_3981);
or U4258 (N_4258,N_3750,N_3339);
nor U4259 (N_4259,N_3994,N_3907);
or U4260 (N_4260,N_3292,N_3444);
xor U4261 (N_4261,N_3387,N_3546);
and U4262 (N_4262,N_3624,N_3287);
or U4263 (N_4263,N_3343,N_3401);
or U4264 (N_4264,N_3714,N_3385);
nand U4265 (N_4265,N_3800,N_3390);
xnor U4266 (N_4266,N_3296,N_3507);
and U4267 (N_4267,N_3822,N_3744);
and U4268 (N_4268,N_3535,N_3371);
or U4269 (N_4269,N_3897,N_3446);
nor U4270 (N_4270,N_3936,N_3989);
nand U4271 (N_4271,N_3074,N_3521);
and U4272 (N_4272,N_3876,N_3475);
or U4273 (N_4273,N_3511,N_3255);
and U4274 (N_4274,N_3520,N_3297);
nand U4275 (N_4275,N_3927,N_3783);
xor U4276 (N_4276,N_3833,N_3145);
or U4277 (N_4277,N_3758,N_3695);
nor U4278 (N_4278,N_3685,N_3499);
xor U4279 (N_4279,N_3972,N_3353);
nand U4280 (N_4280,N_3771,N_3130);
xor U4281 (N_4281,N_3463,N_3561);
nor U4282 (N_4282,N_3899,N_3569);
xnor U4283 (N_4283,N_3221,N_3549);
xnor U4284 (N_4284,N_3326,N_3526);
xnor U4285 (N_4285,N_3480,N_3945);
or U4286 (N_4286,N_3999,N_3261);
xnor U4287 (N_4287,N_3181,N_3344);
and U4288 (N_4288,N_3072,N_3246);
xnor U4289 (N_4289,N_3018,N_3148);
xor U4290 (N_4290,N_3188,N_3458);
nor U4291 (N_4291,N_3152,N_3715);
nor U4292 (N_4292,N_3278,N_3909);
nand U4293 (N_4293,N_3804,N_3738);
or U4294 (N_4294,N_3843,N_3363);
nor U4295 (N_4295,N_3547,N_3946);
nand U4296 (N_4296,N_3589,N_3834);
or U4297 (N_4297,N_3868,N_3056);
nand U4298 (N_4298,N_3536,N_3029);
and U4299 (N_4299,N_3374,N_3514);
and U4300 (N_4300,N_3943,N_3840);
and U4301 (N_4301,N_3275,N_3021);
nand U4302 (N_4302,N_3043,N_3501);
xor U4303 (N_4303,N_3122,N_3236);
and U4304 (N_4304,N_3540,N_3996);
nor U4305 (N_4305,N_3049,N_3984);
and U4306 (N_4306,N_3372,N_3935);
xnor U4307 (N_4307,N_3717,N_3964);
xor U4308 (N_4308,N_3166,N_3688);
and U4309 (N_4309,N_3200,N_3505);
or U4310 (N_4310,N_3361,N_3426);
xnor U4311 (N_4311,N_3962,N_3327);
and U4312 (N_4312,N_3777,N_3170);
xnor U4313 (N_4313,N_3577,N_3787);
or U4314 (N_4314,N_3959,N_3054);
nor U4315 (N_4315,N_3728,N_3846);
or U4316 (N_4316,N_3755,N_3358);
or U4317 (N_4317,N_3055,N_3088);
xor U4318 (N_4318,N_3017,N_3851);
xor U4319 (N_4319,N_3797,N_3421);
or U4320 (N_4320,N_3588,N_3866);
nand U4321 (N_4321,N_3929,N_3542);
and U4322 (N_4322,N_3939,N_3847);
xor U4323 (N_4323,N_3529,N_3209);
nor U4324 (N_4324,N_3453,N_3616);
nor U4325 (N_4325,N_3841,N_3720);
nor U4326 (N_4326,N_3835,N_3992);
nor U4327 (N_4327,N_3235,N_3139);
or U4328 (N_4328,N_3172,N_3940);
nand U4329 (N_4329,N_3487,N_3983);
nor U4330 (N_4330,N_3563,N_3623);
nand U4331 (N_4331,N_3784,N_3806);
nor U4332 (N_4332,N_3605,N_3900);
nand U4333 (N_4333,N_3126,N_3131);
or U4334 (N_4334,N_3969,N_3718);
nor U4335 (N_4335,N_3123,N_3164);
nand U4336 (N_4336,N_3891,N_3331);
nand U4337 (N_4337,N_3553,N_3884);
nor U4338 (N_4338,N_3644,N_3638);
or U4339 (N_4339,N_3922,N_3193);
nor U4340 (N_4340,N_3747,N_3115);
nor U4341 (N_4341,N_3050,N_3942);
and U4342 (N_4342,N_3887,N_3241);
or U4343 (N_4343,N_3903,N_3933);
and U4344 (N_4344,N_3408,N_3552);
nand U4345 (N_4345,N_3189,N_3346);
xnor U4346 (N_4346,N_3238,N_3041);
xnor U4347 (N_4347,N_3816,N_3211);
xnor U4348 (N_4348,N_3704,N_3413);
nor U4349 (N_4349,N_3362,N_3156);
and U4350 (N_4350,N_3764,N_3250);
nor U4351 (N_4351,N_3010,N_3274);
xnor U4352 (N_4352,N_3855,N_3759);
xnor U4353 (N_4353,N_3437,N_3405);
or U4354 (N_4354,N_3754,N_3697);
nand U4355 (N_4355,N_3219,N_3726);
and U4356 (N_4356,N_3381,N_3786);
nor U4357 (N_4357,N_3889,N_3234);
nor U4358 (N_4358,N_3216,N_3604);
or U4359 (N_4359,N_3617,N_3653);
or U4360 (N_4360,N_3081,N_3504);
nand U4361 (N_4361,N_3253,N_3908);
or U4362 (N_4362,N_3430,N_3928);
nor U4363 (N_4363,N_3110,N_3433);
and U4364 (N_4364,N_3741,N_3769);
nor U4365 (N_4365,N_3215,N_3951);
xor U4366 (N_4366,N_3441,N_3877);
nand U4367 (N_4367,N_3058,N_3872);
or U4368 (N_4368,N_3978,N_3490);
and U4369 (N_4369,N_3309,N_3452);
nor U4370 (N_4370,N_3956,N_3701);
nand U4371 (N_4371,N_3042,N_3120);
nand U4372 (N_4372,N_3792,N_3417);
nand U4373 (N_4373,N_3793,N_3141);
and U4374 (N_4374,N_3603,N_3661);
nor U4375 (N_4375,N_3727,N_3853);
xor U4376 (N_4376,N_3226,N_3150);
xor U4377 (N_4377,N_3295,N_3319);
nand U4378 (N_4378,N_3324,N_3752);
and U4379 (N_4379,N_3204,N_3805);
nand U4380 (N_4380,N_3077,N_3762);
nand U4381 (N_4381,N_3035,N_3934);
and U4382 (N_4382,N_3649,N_3477);
or U4383 (N_4383,N_3210,N_3630);
nor U4384 (N_4384,N_3008,N_3121);
nor U4385 (N_4385,N_3869,N_3931);
nand U4386 (N_4386,N_3636,N_3963);
or U4387 (N_4387,N_3288,N_3137);
nand U4388 (N_4388,N_3006,N_3830);
and U4389 (N_4389,N_3628,N_3533);
xor U4390 (N_4390,N_3386,N_3878);
nand U4391 (N_4391,N_3399,N_3724);
or U4392 (N_4392,N_3968,N_3861);
or U4393 (N_4393,N_3719,N_3012);
xor U4394 (N_4394,N_3798,N_3860);
or U4395 (N_4395,N_3671,N_3282);
nand U4396 (N_4396,N_3260,N_3749);
xor U4397 (N_4397,N_3001,N_3665);
nand U4398 (N_4398,N_3062,N_3435);
nand U4399 (N_4399,N_3799,N_3647);
and U4400 (N_4400,N_3723,N_3873);
nand U4401 (N_4401,N_3442,N_3277);
nand U4402 (N_4402,N_3543,N_3760);
nor U4403 (N_4403,N_3406,N_3765);
xnor U4404 (N_4404,N_3815,N_3162);
and U4405 (N_4405,N_3683,N_3119);
or U4406 (N_4406,N_3447,N_3831);
and U4407 (N_4407,N_3300,N_3842);
nand U4408 (N_4408,N_3315,N_3895);
nand U4409 (N_4409,N_3455,N_3706);
nor U4410 (N_4410,N_3474,N_3489);
xor U4411 (N_4411,N_3334,N_3389);
xnor U4412 (N_4412,N_3303,N_3037);
or U4413 (N_4413,N_3057,N_3003);
and U4414 (N_4414,N_3013,N_3743);
nand U4415 (N_4415,N_3243,N_3290);
nand U4416 (N_4416,N_3456,N_3660);
nand U4417 (N_4417,N_3159,N_3019);
nor U4418 (N_4418,N_3388,N_3663);
nor U4419 (N_4419,N_3391,N_3858);
nand U4420 (N_4420,N_3892,N_3134);
or U4421 (N_4421,N_3322,N_3272);
nor U4422 (N_4422,N_3342,N_3206);
nor U4423 (N_4423,N_3097,N_3497);
nand U4424 (N_4424,N_3461,N_3703);
nor U4425 (N_4425,N_3698,N_3606);
or U4426 (N_4426,N_3592,N_3423);
xor U4427 (N_4427,N_3096,N_3026);
and U4428 (N_4428,N_3721,N_3924);
nand U4429 (N_4429,N_3856,N_3534);
or U4430 (N_4430,N_3345,N_3176);
or U4431 (N_4431,N_3690,N_3218);
nor U4432 (N_4432,N_3693,N_3059);
and U4433 (N_4433,N_3599,N_3998);
nand U4434 (N_4434,N_3579,N_3819);
nor U4435 (N_4435,N_3560,N_3020);
and U4436 (N_4436,N_3015,N_3528);
nand U4437 (N_4437,N_3414,N_3993);
nor U4438 (N_4438,N_3462,N_3025);
xnor U4439 (N_4439,N_3574,N_3267);
nor U4440 (N_4440,N_3820,N_3313);
nor U4441 (N_4441,N_3921,N_3063);
nor U4442 (N_4442,N_3048,N_3481);
and U4443 (N_4443,N_3136,N_3359);
xor U4444 (N_4444,N_3548,N_3080);
xnor U4445 (N_4445,N_3187,N_3668);
nand U4446 (N_4446,N_3896,N_3615);
xor U4447 (N_4447,N_3829,N_3854);
or U4448 (N_4448,N_3961,N_3849);
nand U4449 (N_4449,N_3500,N_3163);
xor U4450 (N_4450,N_3675,N_3725);
and U4451 (N_4451,N_3146,N_3397);
xnor U4452 (N_4452,N_3593,N_3168);
nand U4453 (N_4453,N_3138,N_3201);
xor U4454 (N_4454,N_3085,N_3985);
nor U4455 (N_4455,N_3129,N_3905);
nand U4456 (N_4456,N_3646,N_3519);
nand U4457 (N_4457,N_3568,N_3254);
xnor U4458 (N_4458,N_3224,N_3068);
or U4459 (N_4459,N_3523,N_3776);
and U4460 (N_4460,N_3252,N_3266);
nand U4461 (N_4461,N_3486,N_3382);
nand U4462 (N_4462,N_3766,N_3171);
and U4463 (N_4463,N_3192,N_3459);
or U4464 (N_4464,N_3230,N_3227);
and U4465 (N_4465,N_3375,N_3233);
xor U4466 (N_4466,N_3105,N_3902);
nand U4467 (N_4467,N_3427,N_3409);
nor U4468 (N_4468,N_3377,N_3554);
nand U4469 (N_4469,N_3558,N_3751);
nor U4470 (N_4470,N_3439,N_3512);
nor U4471 (N_4471,N_3502,N_3457);
or U4472 (N_4472,N_3914,N_3434);
nor U4473 (N_4473,N_3493,N_3508);
or U4474 (N_4474,N_3571,N_3429);
and U4475 (N_4475,N_3586,N_3109);
xor U4476 (N_4476,N_3316,N_3756);
xnor U4477 (N_4477,N_3844,N_3982);
nand U4478 (N_4478,N_3198,N_3882);
nor U4479 (N_4479,N_3774,N_3237);
nand U4480 (N_4480,N_3073,N_3953);
and U4481 (N_4481,N_3785,N_3867);
or U4482 (N_4482,N_3662,N_3510);
or U4483 (N_4483,N_3135,N_3498);
nand U4484 (N_4484,N_3184,N_3790);
and U4485 (N_4485,N_3782,N_3352);
nor U4486 (N_4486,N_3419,N_3485);
xor U4487 (N_4487,N_3708,N_3648);
nor U4488 (N_4488,N_3089,N_3702);
and U4489 (N_4489,N_3901,N_3445);
xor U4490 (N_4490,N_3779,N_3229);
nand U4491 (N_4491,N_3614,N_3808);
nor U4492 (N_4492,N_3975,N_3321);
xnor U4493 (N_4493,N_3973,N_3823);
nor U4494 (N_4494,N_3231,N_3155);
or U4495 (N_4495,N_3991,N_3065);
nand U4496 (N_4496,N_3438,N_3664);
nor U4497 (N_4497,N_3076,N_3281);
and U4498 (N_4498,N_3600,N_3270);
and U4499 (N_4499,N_3826,N_3125);
and U4500 (N_4500,N_3358,N_3454);
and U4501 (N_4501,N_3044,N_3731);
and U4502 (N_4502,N_3908,N_3224);
or U4503 (N_4503,N_3651,N_3787);
and U4504 (N_4504,N_3413,N_3316);
xnor U4505 (N_4505,N_3525,N_3433);
or U4506 (N_4506,N_3032,N_3493);
nand U4507 (N_4507,N_3954,N_3353);
nor U4508 (N_4508,N_3713,N_3465);
or U4509 (N_4509,N_3857,N_3126);
and U4510 (N_4510,N_3827,N_3839);
xor U4511 (N_4511,N_3265,N_3524);
and U4512 (N_4512,N_3802,N_3321);
xnor U4513 (N_4513,N_3645,N_3473);
nor U4514 (N_4514,N_3174,N_3013);
nor U4515 (N_4515,N_3545,N_3832);
or U4516 (N_4516,N_3443,N_3876);
or U4517 (N_4517,N_3507,N_3676);
nor U4518 (N_4518,N_3436,N_3272);
or U4519 (N_4519,N_3012,N_3374);
or U4520 (N_4520,N_3211,N_3501);
nor U4521 (N_4521,N_3276,N_3481);
nand U4522 (N_4522,N_3336,N_3386);
xnor U4523 (N_4523,N_3900,N_3648);
or U4524 (N_4524,N_3232,N_3171);
or U4525 (N_4525,N_3018,N_3851);
nor U4526 (N_4526,N_3176,N_3108);
nor U4527 (N_4527,N_3316,N_3652);
or U4528 (N_4528,N_3260,N_3204);
xor U4529 (N_4529,N_3230,N_3200);
nor U4530 (N_4530,N_3636,N_3578);
nor U4531 (N_4531,N_3203,N_3651);
nand U4532 (N_4532,N_3467,N_3000);
xor U4533 (N_4533,N_3290,N_3827);
or U4534 (N_4534,N_3075,N_3968);
xnor U4535 (N_4535,N_3151,N_3221);
nor U4536 (N_4536,N_3849,N_3110);
or U4537 (N_4537,N_3200,N_3779);
xor U4538 (N_4538,N_3776,N_3238);
and U4539 (N_4539,N_3467,N_3697);
nand U4540 (N_4540,N_3179,N_3801);
nor U4541 (N_4541,N_3928,N_3086);
or U4542 (N_4542,N_3399,N_3422);
xnor U4543 (N_4543,N_3423,N_3827);
nand U4544 (N_4544,N_3421,N_3101);
or U4545 (N_4545,N_3181,N_3816);
nor U4546 (N_4546,N_3711,N_3477);
or U4547 (N_4547,N_3746,N_3870);
and U4548 (N_4548,N_3918,N_3974);
nor U4549 (N_4549,N_3171,N_3724);
nor U4550 (N_4550,N_3890,N_3719);
xnor U4551 (N_4551,N_3157,N_3863);
nand U4552 (N_4552,N_3660,N_3587);
nand U4553 (N_4553,N_3315,N_3387);
xor U4554 (N_4554,N_3680,N_3703);
and U4555 (N_4555,N_3075,N_3103);
and U4556 (N_4556,N_3699,N_3346);
nand U4557 (N_4557,N_3023,N_3150);
nand U4558 (N_4558,N_3235,N_3938);
or U4559 (N_4559,N_3657,N_3854);
nor U4560 (N_4560,N_3381,N_3537);
nor U4561 (N_4561,N_3416,N_3507);
nor U4562 (N_4562,N_3271,N_3366);
xnor U4563 (N_4563,N_3725,N_3041);
and U4564 (N_4564,N_3513,N_3537);
xnor U4565 (N_4565,N_3029,N_3635);
and U4566 (N_4566,N_3392,N_3316);
nand U4567 (N_4567,N_3128,N_3768);
and U4568 (N_4568,N_3057,N_3790);
nor U4569 (N_4569,N_3172,N_3870);
and U4570 (N_4570,N_3533,N_3442);
xor U4571 (N_4571,N_3096,N_3191);
nor U4572 (N_4572,N_3201,N_3891);
or U4573 (N_4573,N_3348,N_3681);
or U4574 (N_4574,N_3735,N_3537);
nor U4575 (N_4575,N_3937,N_3474);
nand U4576 (N_4576,N_3892,N_3962);
nor U4577 (N_4577,N_3080,N_3845);
and U4578 (N_4578,N_3676,N_3411);
and U4579 (N_4579,N_3846,N_3370);
or U4580 (N_4580,N_3220,N_3040);
and U4581 (N_4581,N_3573,N_3607);
or U4582 (N_4582,N_3215,N_3156);
xor U4583 (N_4583,N_3798,N_3839);
or U4584 (N_4584,N_3463,N_3994);
nor U4585 (N_4585,N_3986,N_3348);
or U4586 (N_4586,N_3904,N_3024);
xnor U4587 (N_4587,N_3901,N_3354);
xnor U4588 (N_4588,N_3844,N_3572);
and U4589 (N_4589,N_3030,N_3119);
xnor U4590 (N_4590,N_3821,N_3035);
xor U4591 (N_4591,N_3986,N_3804);
nor U4592 (N_4592,N_3097,N_3684);
or U4593 (N_4593,N_3974,N_3045);
nand U4594 (N_4594,N_3332,N_3449);
nand U4595 (N_4595,N_3692,N_3119);
or U4596 (N_4596,N_3600,N_3526);
xnor U4597 (N_4597,N_3471,N_3570);
nor U4598 (N_4598,N_3869,N_3057);
nand U4599 (N_4599,N_3987,N_3909);
xnor U4600 (N_4600,N_3742,N_3450);
xnor U4601 (N_4601,N_3152,N_3178);
and U4602 (N_4602,N_3612,N_3480);
nor U4603 (N_4603,N_3833,N_3252);
xnor U4604 (N_4604,N_3562,N_3698);
nor U4605 (N_4605,N_3571,N_3895);
or U4606 (N_4606,N_3151,N_3528);
xor U4607 (N_4607,N_3576,N_3214);
nor U4608 (N_4608,N_3977,N_3351);
and U4609 (N_4609,N_3336,N_3310);
or U4610 (N_4610,N_3627,N_3356);
or U4611 (N_4611,N_3888,N_3379);
nand U4612 (N_4612,N_3960,N_3443);
nand U4613 (N_4613,N_3266,N_3168);
nand U4614 (N_4614,N_3830,N_3808);
and U4615 (N_4615,N_3294,N_3218);
and U4616 (N_4616,N_3948,N_3328);
nand U4617 (N_4617,N_3216,N_3330);
or U4618 (N_4618,N_3653,N_3544);
or U4619 (N_4619,N_3063,N_3829);
xnor U4620 (N_4620,N_3307,N_3818);
or U4621 (N_4621,N_3322,N_3666);
and U4622 (N_4622,N_3579,N_3432);
and U4623 (N_4623,N_3990,N_3137);
nor U4624 (N_4624,N_3148,N_3356);
nand U4625 (N_4625,N_3753,N_3544);
or U4626 (N_4626,N_3786,N_3005);
xor U4627 (N_4627,N_3910,N_3794);
xnor U4628 (N_4628,N_3178,N_3851);
nand U4629 (N_4629,N_3197,N_3400);
nand U4630 (N_4630,N_3387,N_3620);
and U4631 (N_4631,N_3048,N_3378);
xnor U4632 (N_4632,N_3832,N_3679);
nor U4633 (N_4633,N_3978,N_3095);
or U4634 (N_4634,N_3637,N_3087);
and U4635 (N_4635,N_3249,N_3740);
xor U4636 (N_4636,N_3949,N_3255);
and U4637 (N_4637,N_3692,N_3444);
and U4638 (N_4638,N_3188,N_3577);
and U4639 (N_4639,N_3628,N_3084);
and U4640 (N_4640,N_3561,N_3817);
or U4641 (N_4641,N_3379,N_3261);
nand U4642 (N_4642,N_3171,N_3013);
nand U4643 (N_4643,N_3980,N_3191);
and U4644 (N_4644,N_3047,N_3847);
nand U4645 (N_4645,N_3655,N_3584);
nor U4646 (N_4646,N_3600,N_3631);
xor U4647 (N_4647,N_3449,N_3679);
nand U4648 (N_4648,N_3460,N_3683);
nor U4649 (N_4649,N_3663,N_3351);
nand U4650 (N_4650,N_3235,N_3730);
or U4651 (N_4651,N_3067,N_3296);
nor U4652 (N_4652,N_3260,N_3273);
nor U4653 (N_4653,N_3936,N_3981);
and U4654 (N_4654,N_3770,N_3431);
nand U4655 (N_4655,N_3136,N_3612);
and U4656 (N_4656,N_3483,N_3453);
nor U4657 (N_4657,N_3151,N_3845);
nor U4658 (N_4658,N_3870,N_3086);
xnor U4659 (N_4659,N_3898,N_3795);
and U4660 (N_4660,N_3105,N_3318);
nand U4661 (N_4661,N_3111,N_3733);
xor U4662 (N_4662,N_3345,N_3435);
xnor U4663 (N_4663,N_3926,N_3038);
xnor U4664 (N_4664,N_3557,N_3334);
or U4665 (N_4665,N_3639,N_3370);
nor U4666 (N_4666,N_3115,N_3988);
nand U4667 (N_4667,N_3646,N_3431);
or U4668 (N_4668,N_3368,N_3921);
nand U4669 (N_4669,N_3178,N_3731);
nor U4670 (N_4670,N_3126,N_3928);
or U4671 (N_4671,N_3981,N_3260);
xnor U4672 (N_4672,N_3110,N_3132);
and U4673 (N_4673,N_3546,N_3275);
or U4674 (N_4674,N_3165,N_3396);
and U4675 (N_4675,N_3389,N_3328);
xnor U4676 (N_4676,N_3551,N_3068);
or U4677 (N_4677,N_3382,N_3734);
nor U4678 (N_4678,N_3092,N_3064);
or U4679 (N_4679,N_3583,N_3916);
nand U4680 (N_4680,N_3117,N_3880);
nand U4681 (N_4681,N_3705,N_3598);
and U4682 (N_4682,N_3069,N_3987);
and U4683 (N_4683,N_3829,N_3465);
nor U4684 (N_4684,N_3941,N_3398);
or U4685 (N_4685,N_3200,N_3480);
or U4686 (N_4686,N_3856,N_3748);
nor U4687 (N_4687,N_3947,N_3577);
xnor U4688 (N_4688,N_3611,N_3420);
nor U4689 (N_4689,N_3853,N_3645);
or U4690 (N_4690,N_3801,N_3593);
nor U4691 (N_4691,N_3729,N_3679);
nor U4692 (N_4692,N_3234,N_3496);
nor U4693 (N_4693,N_3493,N_3849);
or U4694 (N_4694,N_3309,N_3290);
or U4695 (N_4695,N_3164,N_3471);
nand U4696 (N_4696,N_3234,N_3269);
or U4697 (N_4697,N_3963,N_3755);
xor U4698 (N_4698,N_3782,N_3902);
nor U4699 (N_4699,N_3199,N_3950);
or U4700 (N_4700,N_3995,N_3054);
and U4701 (N_4701,N_3285,N_3077);
or U4702 (N_4702,N_3770,N_3300);
nor U4703 (N_4703,N_3266,N_3154);
nor U4704 (N_4704,N_3890,N_3562);
nand U4705 (N_4705,N_3814,N_3752);
nand U4706 (N_4706,N_3200,N_3774);
nor U4707 (N_4707,N_3174,N_3666);
nor U4708 (N_4708,N_3872,N_3082);
or U4709 (N_4709,N_3308,N_3299);
nand U4710 (N_4710,N_3171,N_3706);
or U4711 (N_4711,N_3354,N_3156);
or U4712 (N_4712,N_3522,N_3649);
nor U4713 (N_4713,N_3093,N_3328);
or U4714 (N_4714,N_3970,N_3097);
nand U4715 (N_4715,N_3963,N_3067);
xor U4716 (N_4716,N_3008,N_3075);
nand U4717 (N_4717,N_3964,N_3296);
or U4718 (N_4718,N_3749,N_3366);
and U4719 (N_4719,N_3327,N_3589);
xnor U4720 (N_4720,N_3835,N_3193);
nand U4721 (N_4721,N_3137,N_3517);
nand U4722 (N_4722,N_3174,N_3358);
nor U4723 (N_4723,N_3514,N_3315);
nor U4724 (N_4724,N_3378,N_3651);
or U4725 (N_4725,N_3047,N_3414);
nor U4726 (N_4726,N_3992,N_3798);
xor U4727 (N_4727,N_3777,N_3873);
nor U4728 (N_4728,N_3566,N_3685);
nor U4729 (N_4729,N_3821,N_3499);
or U4730 (N_4730,N_3283,N_3864);
nor U4731 (N_4731,N_3155,N_3881);
and U4732 (N_4732,N_3392,N_3116);
and U4733 (N_4733,N_3290,N_3662);
or U4734 (N_4734,N_3569,N_3818);
xor U4735 (N_4735,N_3192,N_3446);
nor U4736 (N_4736,N_3486,N_3399);
nor U4737 (N_4737,N_3224,N_3230);
or U4738 (N_4738,N_3675,N_3201);
nand U4739 (N_4739,N_3747,N_3015);
nand U4740 (N_4740,N_3874,N_3577);
nand U4741 (N_4741,N_3405,N_3580);
and U4742 (N_4742,N_3991,N_3256);
and U4743 (N_4743,N_3817,N_3324);
or U4744 (N_4744,N_3266,N_3039);
or U4745 (N_4745,N_3576,N_3516);
xnor U4746 (N_4746,N_3182,N_3262);
nand U4747 (N_4747,N_3501,N_3870);
nand U4748 (N_4748,N_3752,N_3200);
nand U4749 (N_4749,N_3924,N_3604);
nand U4750 (N_4750,N_3763,N_3428);
nand U4751 (N_4751,N_3022,N_3335);
xnor U4752 (N_4752,N_3146,N_3084);
nand U4753 (N_4753,N_3774,N_3300);
or U4754 (N_4754,N_3571,N_3064);
nand U4755 (N_4755,N_3721,N_3991);
xor U4756 (N_4756,N_3107,N_3015);
xnor U4757 (N_4757,N_3626,N_3189);
xor U4758 (N_4758,N_3004,N_3192);
nand U4759 (N_4759,N_3944,N_3335);
xnor U4760 (N_4760,N_3980,N_3566);
nor U4761 (N_4761,N_3758,N_3965);
nor U4762 (N_4762,N_3699,N_3456);
or U4763 (N_4763,N_3434,N_3060);
nand U4764 (N_4764,N_3164,N_3350);
nand U4765 (N_4765,N_3643,N_3596);
and U4766 (N_4766,N_3254,N_3438);
xnor U4767 (N_4767,N_3325,N_3014);
nor U4768 (N_4768,N_3193,N_3844);
xnor U4769 (N_4769,N_3310,N_3699);
xnor U4770 (N_4770,N_3339,N_3182);
or U4771 (N_4771,N_3482,N_3878);
xor U4772 (N_4772,N_3492,N_3243);
xor U4773 (N_4773,N_3054,N_3281);
xor U4774 (N_4774,N_3540,N_3056);
or U4775 (N_4775,N_3392,N_3344);
nor U4776 (N_4776,N_3924,N_3224);
or U4777 (N_4777,N_3604,N_3764);
xor U4778 (N_4778,N_3287,N_3325);
xor U4779 (N_4779,N_3372,N_3527);
or U4780 (N_4780,N_3981,N_3773);
and U4781 (N_4781,N_3347,N_3645);
xnor U4782 (N_4782,N_3714,N_3483);
or U4783 (N_4783,N_3628,N_3113);
and U4784 (N_4784,N_3373,N_3953);
nor U4785 (N_4785,N_3383,N_3533);
or U4786 (N_4786,N_3480,N_3494);
nor U4787 (N_4787,N_3109,N_3416);
nand U4788 (N_4788,N_3585,N_3745);
nand U4789 (N_4789,N_3098,N_3224);
nand U4790 (N_4790,N_3127,N_3566);
xnor U4791 (N_4791,N_3332,N_3593);
and U4792 (N_4792,N_3162,N_3317);
and U4793 (N_4793,N_3376,N_3374);
xnor U4794 (N_4794,N_3197,N_3584);
and U4795 (N_4795,N_3723,N_3180);
nor U4796 (N_4796,N_3591,N_3414);
and U4797 (N_4797,N_3237,N_3442);
and U4798 (N_4798,N_3998,N_3285);
or U4799 (N_4799,N_3417,N_3330);
nor U4800 (N_4800,N_3643,N_3268);
xor U4801 (N_4801,N_3854,N_3727);
or U4802 (N_4802,N_3561,N_3928);
or U4803 (N_4803,N_3180,N_3853);
and U4804 (N_4804,N_3203,N_3701);
and U4805 (N_4805,N_3397,N_3305);
nand U4806 (N_4806,N_3909,N_3398);
or U4807 (N_4807,N_3719,N_3886);
and U4808 (N_4808,N_3374,N_3819);
and U4809 (N_4809,N_3404,N_3007);
nor U4810 (N_4810,N_3270,N_3645);
and U4811 (N_4811,N_3485,N_3424);
nand U4812 (N_4812,N_3402,N_3829);
xnor U4813 (N_4813,N_3977,N_3209);
nand U4814 (N_4814,N_3811,N_3557);
or U4815 (N_4815,N_3905,N_3509);
and U4816 (N_4816,N_3884,N_3377);
xnor U4817 (N_4817,N_3195,N_3209);
nand U4818 (N_4818,N_3815,N_3261);
nor U4819 (N_4819,N_3274,N_3717);
nor U4820 (N_4820,N_3626,N_3515);
and U4821 (N_4821,N_3513,N_3172);
or U4822 (N_4822,N_3916,N_3745);
xor U4823 (N_4823,N_3748,N_3827);
and U4824 (N_4824,N_3518,N_3678);
nand U4825 (N_4825,N_3950,N_3974);
nor U4826 (N_4826,N_3345,N_3313);
or U4827 (N_4827,N_3270,N_3079);
or U4828 (N_4828,N_3426,N_3776);
nor U4829 (N_4829,N_3291,N_3593);
nand U4830 (N_4830,N_3888,N_3643);
and U4831 (N_4831,N_3777,N_3320);
or U4832 (N_4832,N_3907,N_3949);
or U4833 (N_4833,N_3907,N_3685);
or U4834 (N_4834,N_3408,N_3290);
nor U4835 (N_4835,N_3556,N_3521);
and U4836 (N_4836,N_3239,N_3531);
xor U4837 (N_4837,N_3290,N_3089);
nor U4838 (N_4838,N_3162,N_3484);
and U4839 (N_4839,N_3681,N_3299);
xor U4840 (N_4840,N_3257,N_3855);
or U4841 (N_4841,N_3903,N_3180);
and U4842 (N_4842,N_3866,N_3272);
or U4843 (N_4843,N_3631,N_3592);
or U4844 (N_4844,N_3753,N_3831);
nor U4845 (N_4845,N_3188,N_3718);
or U4846 (N_4846,N_3559,N_3404);
nor U4847 (N_4847,N_3841,N_3592);
nand U4848 (N_4848,N_3555,N_3407);
or U4849 (N_4849,N_3879,N_3781);
nor U4850 (N_4850,N_3030,N_3172);
and U4851 (N_4851,N_3937,N_3065);
nor U4852 (N_4852,N_3354,N_3416);
nand U4853 (N_4853,N_3805,N_3617);
nand U4854 (N_4854,N_3993,N_3253);
nand U4855 (N_4855,N_3557,N_3473);
or U4856 (N_4856,N_3054,N_3876);
nand U4857 (N_4857,N_3179,N_3660);
or U4858 (N_4858,N_3076,N_3720);
xor U4859 (N_4859,N_3551,N_3224);
nor U4860 (N_4860,N_3854,N_3745);
nor U4861 (N_4861,N_3119,N_3838);
and U4862 (N_4862,N_3272,N_3445);
nor U4863 (N_4863,N_3899,N_3660);
and U4864 (N_4864,N_3922,N_3006);
xnor U4865 (N_4865,N_3739,N_3111);
or U4866 (N_4866,N_3984,N_3973);
or U4867 (N_4867,N_3314,N_3320);
and U4868 (N_4868,N_3743,N_3074);
xnor U4869 (N_4869,N_3900,N_3700);
or U4870 (N_4870,N_3471,N_3493);
nor U4871 (N_4871,N_3927,N_3454);
xor U4872 (N_4872,N_3676,N_3851);
or U4873 (N_4873,N_3766,N_3824);
xor U4874 (N_4874,N_3052,N_3049);
nand U4875 (N_4875,N_3802,N_3398);
nand U4876 (N_4876,N_3763,N_3741);
nand U4877 (N_4877,N_3414,N_3659);
and U4878 (N_4878,N_3746,N_3026);
xnor U4879 (N_4879,N_3475,N_3493);
xnor U4880 (N_4880,N_3519,N_3585);
nand U4881 (N_4881,N_3565,N_3766);
xor U4882 (N_4882,N_3866,N_3895);
xor U4883 (N_4883,N_3695,N_3773);
xor U4884 (N_4884,N_3659,N_3425);
or U4885 (N_4885,N_3031,N_3777);
nor U4886 (N_4886,N_3792,N_3846);
nand U4887 (N_4887,N_3116,N_3781);
nand U4888 (N_4888,N_3057,N_3954);
and U4889 (N_4889,N_3566,N_3665);
and U4890 (N_4890,N_3381,N_3593);
or U4891 (N_4891,N_3607,N_3892);
and U4892 (N_4892,N_3587,N_3053);
and U4893 (N_4893,N_3944,N_3129);
or U4894 (N_4894,N_3946,N_3802);
nor U4895 (N_4895,N_3184,N_3705);
nand U4896 (N_4896,N_3473,N_3872);
and U4897 (N_4897,N_3002,N_3626);
or U4898 (N_4898,N_3762,N_3074);
or U4899 (N_4899,N_3892,N_3037);
and U4900 (N_4900,N_3021,N_3377);
xor U4901 (N_4901,N_3132,N_3307);
nand U4902 (N_4902,N_3000,N_3293);
nor U4903 (N_4903,N_3128,N_3025);
and U4904 (N_4904,N_3474,N_3686);
and U4905 (N_4905,N_3047,N_3271);
or U4906 (N_4906,N_3057,N_3257);
and U4907 (N_4907,N_3141,N_3381);
nor U4908 (N_4908,N_3196,N_3769);
or U4909 (N_4909,N_3699,N_3759);
nand U4910 (N_4910,N_3475,N_3796);
nor U4911 (N_4911,N_3431,N_3025);
nand U4912 (N_4912,N_3178,N_3989);
or U4913 (N_4913,N_3557,N_3006);
nand U4914 (N_4914,N_3908,N_3789);
or U4915 (N_4915,N_3742,N_3928);
and U4916 (N_4916,N_3028,N_3091);
and U4917 (N_4917,N_3923,N_3091);
xor U4918 (N_4918,N_3916,N_3680);
xor U4919 (N_4919,N_3209,N_3851);
nand U4920 (N_4920,N_3209,N_3534);
and U4921 (N_4921,N_3528,N_3037);
nor U4922 (N_4922,N_3009,N_3609);
nor U4923 (N_4923,N_3654,N_3436);
xnor U4924 (N_4924,N_3863,N_3742);
nand U4925 (N_4925,N_3611,N_3482);
nand U4926 (N_4926,N_3157,N_3635);
or U4927 (N_4927,N_3732,N_3581);
nor U4928 (N_4928,N_3453,N_3773);
and U4929 (N_4929,N_3770,N_3230);
nand U4930 (N_4930,N_3111,N_3609);
xnor U4931 (N_4931,N_3105,N_3802);
xor U4932 (N_4932,N_3204,N_3136);
xnor U4933 (N_4933,N_3244,N_3015);
xnor U4934 (N_4934,N_3954,N_3389);
and U4935 (N_4935,N_3398,N_3035);
or U4936 (N_4936,N_3593,N_3745);
or U4937 (N_4937,N_3989,N_3084);
or U4938 (N_4938,N_3026,N_3158);
and U4939 (N_4939,N_3964,N_3672);
nor U4940 (N_4940,N_3882,N_3184);
xor U4941 (N_4941,N_3708,N_3623);
and U4942 (N_4942,N_3985,N_3371);
xnor U4943 (N_4943,N_3533,N_3207);
nand U4944 (N_4944,N_3568,N_3271);
xor U4945 (N_4945,N_3913,N_3702);
and U4946 (N_4946,N_3659,N_3266);
and U4947 (N_4947,N_3834,N_3880);
nand U4948 (N_4948,N_3203,N_3970);
nor U4949 (N_4949,N_3131,N_3928);
and U4950 (N_4950,N_3565,N_3811);
nand U4951 (N_4951,N_3628,N_3797);
or U4952 (N_4952,N_3163,N_3161);
xnor U4953 (N_4953,N_3149,N_3936);
nand U4954 (N_4954,N_3728,N_3125);
and U4955 (N_4955,N_3849,N_3306);
and U4956 (N_4956,N_3858,N_3738);
nand U4957 (N_4957,N_3188,N_3602);
and U4958 (N_4958,N_3755,N_3689);
nand U4959 (N_4959,N_3952,N_3116);
nand U4960 (N_4960,N_3136,N_3077);
nand U4961 (N_4961,N_3810,N_3145);
or U4962 (N_4962,N_3673,N_3105);
or U4963 (N_4963,N_3618,N_3141);
nor U4964 (N_4964,N_3639,N_3276);
and U4965 (N_4965,N_3245,N_3799);
nand U4966 (N_4966,N_3137,N_3621);
or U4967 (N_4967,N_3829,N_3542);
or U4968 (N_4968,N_3070,N_3591);
nand U4969 (N_4969,N_3583,N_3371);
nor U4970 (N_4970,N_3665,N_3614);
and U4971 (N_4971,N_3134,N_3957);
or U4972 (N_4972,N_3633,N_3366);
nor U4973 (N_4973,N_3125,N_3571);
nand U4974 (N_4974,N_3803,N_3112);
nor U4975 (N_4975,N_3248,N_3259);
nand U4976 (N_4976,N_3812,N_3406);
or U4977 (N_4977,N_3240,N_3728);
xnor U4978 (N_4978,N_3173,N_3614);
xor U4979 (N_4979,N_3923,N_3646);
xor U4980 (N_4980,N_3688,N_3810);
or U4981 (N_4981,N_3376,N_3086);
nor U4982 (N_4982,N_3543,N_3174);
nand U4983 (N_4983,N_3371,N_3643);
nand U4984 (N_4984,N_3649,N_3811);
xnor U4985 (N_4985,N_3573,N_3869);
or U4986 (N_4986,N_3382,N_3946);
and U4987 (N_4987,N_3637,N_3927);
nor U4988 (N_4988,N_3110,N_3673);
nand U4989 (N_4989,N_3038,N_3726);
and U4990 (N_4990,N_3046,N_3767);
and U4991 (N_4991,N_3922,N_3126);
and U4992 (N_4992,N_3315,N_3695);
and U4993 (N_4993,N_3096,N_3424);
or U4994 (N_4994,N_3462,N_3040);
xnor U4995 (N_4995,N_3172,N_3962);
or U4996 (N_4996,N_3346,N_3818);
and U4997 (N_4997,N_3164,N_3149);
and U4998 (N_4998,N_3491,N_3965);
and U4999 (N_4999,N_3253,N_3668);
nor U5000 (N_5000,N_4968,N_4399);
or U5001 (N_5001,N_4070,N_4899);
and U5002 (N_5002,N_4699,N_4118);
xor U5003 (N_5003,N_4570,N_4471);
or U5004 (N_5004,N_4370,N_4334);
xor U5005 (N_5005,N_4257,N_4622);
or U5006 (N_5006,N_4931,N_4454);
and U5007 (N_5007,N_4295,N_4706);
or U5008 (N_5008,N_4646,N_4615);
nand U5009 (N_5009,N_4209,N_4550);
and U5010 (N_5010,N_4269,N_4344);
xor U5011 (N_5011,N_4720,N_4562);
xnor U5012 (N_5012,N_4945,N_4494);
nor U5013 (N_5013,N_4530,N_4178);
xnor U5014 (N_5014,N_4115,N_4382);
nand U5015 (N_5015,N_4329,N_4145);
and U5016 (N_5016,N_4221,N_4608);
nor U5017 (N_5017,N_4187,N_4419);
and U5018 (N_5018,N_4875,N_4110);
nand U5019 (N_5019,N_4514,N_4149);
or U5020 (N_5020,N_4620,N_4338);
nor U5021 (N_5021,N_4279,N_4464);
xnor U5022 (N_5022,N_4981,N_4618);
and U5023 (N_5023,N_4708,N_4166);
nand U5024 (N_5024,N_4631,N_4974);
or U5025 (N_5025,N_4098,N_4971);
nor U5026 (N_5026,N_4687,N_4616);
nand U5027 (N_5027,N_4964,N_4565);
and U5028 (N_5028,N_4319,N_4633);
and U5029 (N_5029,N_4259,N_4006);
nand U5030 (N_5030,N_4685,N_4223);
nand U5031 (N_5031,N_4249,N_4365);
and U5032 (N_5032,N_4676,N_4171);
and U5033 (N_5033,N_4340,N_4424);
nand U5034 (N_5034,N_4917,N_4815);
and U5035 (N_5035,N_4861,N_4750);
nand U5036 (N_5036,N_4043,N_4129);
xor U5037 (N_5037,N_4577,N_4053);
and U5038 (N_5038,N_4734,N_4077);
nor U5039 (N_5039,N_4341,N_4665);
nand U5040 (N_5040,N_4793,N_4818);
or U5041 (N_5041,N_4575,N_4356);
and U5042 (N_5042,N_4366,N_4813);
xnor U5043 (N_5043,N_4262,N_4359);
and U5044 (N_5044,N_4052,N_4589);
nand U5045 (N_5045,N_4939,N_4950);
xnor U5046 (N_5046,N_4501,N_4039);
xnor U5047 (N_5047,N_4659,N_4679);
xor U5048 (N_5048,N_4474,N_4605);
nand U5049 (N_5049,N_4585,N_4300);
nand U5050 (N_5050,N_4814,N_4060);
xnor U5051 (N_5051,N_4122,N_4536);
nand U5052 (N_5052,N_4477,N_4282);
and U5053 (N_5053,N_4229,N_4730);
nand U5054 (N_5054,N_4508,N_4606);
xnor U5055 (N_5055,N_4363,N_4292);
or U5056 (N_5056,N_4690,N_4709);
nand U5057 (N_5057,N_4417,N_4998);
xnor U5058 (N_5058,N_4179,N_4151);
or U5059 (N_5059,N_4503,N_4152);
xnor U5060 (N_5060,N_4147,N_4901);
and U5061 (N_5061,N_4448,N_4877);
or U5062 (N_5062,N_4138,N_4624);
or U5063 (N_5063,N_4369,N_4302);
nor U5064 (N_5064,N_4032,N_4410);
nand U5065 (N_5065,N_4397,N_4509);
xor U5066 (N_5066,N_4444,N_4207);
or U5067 (N_5067,N_4788,N_4046);
nand U5068 (N_5068,N_4809,N_4507);
xnor U5069 (N_5069,N_4858,N_4271);
nand U5070 (N_5070,N_4041,N_4342);
or U5071 (N_5071,N_4924,N_4090);
nor U5072 (N_5072,N_4218,N_4353);
xnor U5073 (N_5073,N_4026,N_4495);
or U5074 (N_5074,N_4653,N_4119);
nor U5075 (N_5075,N_4607,N_4848);
xnor U5076 (N_5076,N_4718,N_4893);
and U5077 (N_5077,N_4673,N_4777);
and U5078 (N_5078,N_4787,N_4439);
or U5079 (N_5079,N_4648,N_4322);
nand U5080 (N_5080,N_4016,N_4386);
and U5081 (N_5081,N_4120,N_4521);
xor U5082 (N_5082,N_4746,N_4908);
nand U5083 (N_5083,N_4754,N_4104);
and U5084 (N_5084,N_4933,N_4668);
nor U5085 (N_5085,N_4472,N_4484);
xor U5086 (N_5086,N_4458,N_4447);
or U5087 (N_5087,N_4594,N_4581);
and U5088 (N_5088,N_4107,N_4599);
nand U5089 (N_5089,N_4505,N_4498);
nand U5090 (N_5090,N_4543,N_4211);
or U5091 (N_5091,N_4527,N_4891);
or U5092 (N_5092,N_4412,N_4136);
nor U5093 (N_5093,N_4422,N_4853);
nand U5094 (N_5094,N_4388,N_4973);
nor U5095 (N_5095,N_4379,N_4184);
xor U5096 (N_5096,N_4666,N_4975);
and U5097 (N_5097,N_4267,N_4871);
nor U5098 (N_5098,N_4384,N_4354);
and U5099 (N_5099,N_4450,N_4492);
and U5100 (N_5100,N_4092,N_4644);
xor U5101 (N_5101,N_4522,N_4431);
and U5102 (N_5102,N_4663,N_4314);
nand U5103 (N_5103,N_4545,N_4897);
xor U5104 (N_5104,N_4266,N_4284);
or U5105 (N_5105,N_4827,N_4778);
or U5106 (N_5106,N_4892,N_4160);
nand U5107 (N_5107,N_4159,N_4729);
nand U5108 (N_5108,N_4671,N_4153);
nand U5109 (N_5109,N_4781,N_4792);
nand U5110 (N_5110,N_4086,N_4749);
or U5111 (N_5111,N_4985,N_4047);
or U5112 (N_5112,N_4073,N_4829);
xor U5113 (N_5113,N_4807,N_4889);
nor U5114 (N_5114,N_4611,N_4768);
and U5115 (N_5115,N_4662,N_4614);
nor U5116 (N_5116,N_4632,N_4854);
or U5117 (N_5117,N_4506,N_4958);
and U5118 (N_5118,N_4802,N_4499);
or U5119 (N_5119,N_4025,N_4113);
nand U5120 (N_5120,N_4967,N_4842);
and U5121 (N_5121,N_4918,N_4031);
and U5122 (N_5122,N_4825,N_4940);
nand U5123 (N_5123,N_4771,N_4821);
or U5124 (N_5124,N_4833,N_4131);
or U5125 (N_5125,N_4672,N_4411);
and U5126 (N_5126,N_4641,N_4057);
nor U5127 (N_5127,N_4828,N_4701);
nor U5128 (N_5128,N_4488,N_4146);
or U5129 (N_5129,N_4045,N_4216);
or U5130 (N_5130,N_4097,N_4868);
xor U5131 (N_5131,N_4072,N_4879);
nand U5132 (N_5132,N_4112,N_4761);
and U5133 (N_5133,N_4519,N_4517);
nor U5134 (N_5134,N_4582,N_4831);
and U5135 (N_5135,N_4638,N_4075);
nor U5136 (N_5136,N_4540,N_4288);
xor U5137 (N_5137,N_4834,N_4215);
nand U5138 (N_5138,N_4776,N_4172);
nand U5139 (N_5139,N_4553,N_4297);
or U5140 (N_5140,N_4111,N_4142);
or U5141 (N_5141,N_4051,N_4261);
nor U5142 (N_5142,N_4883,N_4602);
xnor U5143 (N_5143,N_4976,N_4376);
xnor U5144 (N_5144,N_4515,N_4301);
and U5145 (N_5145,N_4253,N_4005);
or U5146 (N_5146,N_4936,N_4489);
and U5147 (N_5147,N_4626,N_4712);
xnor U5148 (N_5148,N_4955,N_4516);
nand U5149 (N_5149,N_4476,N_4555);
and U5150 (N_5150,N_4841,N_4832);
and U5151 (N_5151,N_4204,N_4198);
or U5152 (N_5152,N_4925,N_4798);
nor U5153 (N_5153,N_4093,N_4739);
nor U5154 (N_5154,N_4935,N_4972);
xor U5155 (N_5155,N_4715,N_4742);
and U5156 (N_5156,N_4135,N_4629);
or U5157 (N_5157,N_4281,N_4864);
nand U5158 (N_5158,N_4014,N_4174);
or U5159 (N_5159,N_4381,N_4083);
or U5160 (N_5160,N_4374,N_4460);
nand U5161 (N_5161,N_4330,N_4843);
xor U5162 (N_5162,N_4256,N_4878);
and U5163 (N_5163,N_4466,N_4678);
nand U5164 (N_5164,N_4909,N_4817);
nand U5165 (N_5165,N_4361,N_4535);
xnor U5166 (N_5166,N_4423,N_4429);
nand U5167 (N_5167,N_4716,N_4590);
xnor U5168 (N_5168,N_4378,N_4385);
nand U5169 (N_5169,N_4510,N_4013);
and U5170 (N_5170,N_4857,N_4299);
or U5171 (N_5171,N_4231,N_4636);
or U5172 (N_5172,N_4681,N_4686);
nand U5173 (N_5173,N_4811,N_4040);
or U5174 (N_5174,N_4309,N_4785);
or U5175 (N_5175,N_4542,N_4453);
nor U5176 (N_5176,N_4434,N_4698);
or U5177 (N_5177,N_4760,N_4664);
xnor U5178 (N_5178,N_4283,N_4426);
or U5179 (N_5179,N_4779,N_4557);
nand U5180 (N_5180,N_4921,N_4068);
or U5181 (N_5181,N_4108,N_4258);
or U5182 (N_5182,N_4658,N_4015);
xor U5183 (N_5183,N_4081,N_4490);
xor U5184 (N_5184,N_4969,N_4089);
nor U5185 (N_5185,N_4774,N_4316);
or U5186 (N_5186,N_4121,N_4881);
nor U5187 (N_5187,N_4613,N_4306);
nand U5188 (N_5188,N_4865,N_4475);
nor U5189 (N_5189,N_4473,N_4004);
xnor U5190 (N_5190,N_4034,N_4688);
nand U5191 (N_5191,N_4723,N_4794);
and U5192 (N_5192,N_4806,N_4949);
nand U5193 (N_5193,N_4704,N_4165);
nand U5194 (N_5194,N_4263,N_4226);
or U5195 (N_5195,N_4091,N_4591);
and U5196 (N_5196,N_4801,N_4994);
nand U5197 (N_5197,N_4937,N_4371);
nand U5198 (N_5198,N_4018,N_4445);
or U5199 (N_5199,N_4406,N_4189);
xnor U5200 (N_5200,N_4639,N_4546);
xnor U5201 (N_5201,N_4775,N_4846);
xnor U5202 (N_5202,N_4059,N_4244);
nand U5203 (N_5203,N_4427,N_4769);
nand U5204 (N_5204,N_4696,N_4432);
nor U5205 (N_5205,N_4640,N_4048);
nor U5206 (N_5206,N_4368,N_4758);
or U5207 (N_5207,N_4010,N_4180);
nand U5208 (N_5208,N_4078,N_4027);
xnor U5209 (N_5209,N_4951,N_4736);
xnor U5210 (N_5210,N_4114,N_4310);
xor U5211 (N_5211,N_4126,N_4812);
and U5212 (N_5212,N_4906,N_4117);
and U5213 (N_5213,N_4203,N_4210);
nand U5214 (N_5214,N_4408,N_4182);
nand U5215 (N_5215,N_4481,N_4360);
xor U5216 (N_5216,N_4199,N_4772);
nor U5217 (N_5217,N_4325,N_4420);
nand U5218 (N_5218,N_4103,N_4230);
and U5219 (N_5219,N_4645,N_4929);
nor U5220 (N_5220,N_4217,N_4449);
nor U5221 (N_5221,N_4849,N_4732);
or U5222 (N_5222,N_4988,N_4030);
nor U5223 (N_5223,N_4038,N_4235);
nand U5224 (N_5224,N_4795,N_4441);
or U5225 (N_5225,N_4593,N_4710);
nand U5226 (N_5226,N_4377,N_4500);
or U5227 (N_5227,N_4446,N_4493);
nor U5228 (N_5228,N_4695,N_4328);
and U5229 (N_5229,N_4173,N_4661);
or U5230 (N_5230,N_4744,N_4437);
or U5231 (N_5231,N_4511,N_4124);
or U5232 (N_5232,N_4600,N_4127);
nand U5233 (N_5233,N_4332,N_4394);
xnor U5234 (N_5234,N_4947,N_4693);
or U5235 (N_5235,N_4396,N_4919);
nor U5236 (N_5236,N_4874,N_4689);
nand U5237 (N_5237,N_4331,N_4095);
xnor U5238 (N_5238,N_4029,N_4375);
or U5239 (N_5239,N_4414,N_4277);
nor U5240 (N_5240,N_4860,N_4986);
xor U5241 (N_5241,N_4738,N_4085);
xor U5242 (N_5242,N_4764,N_4824);
or U5243 (N_5243,N_4934,N_4028);
xor U5244 (N_5244,N_4212,N_4803);
xor U5245 (N_5245,N_4531,N_4911);
nand U5246 (N_5246,N_4463,N_4670);
or U5247 (N_5247,N_4999,N_4957);
and U5248 (N_5248,N_4836,N_4402);
and U5249 (N_5249,N_4168,N_4479);
nand U5250 (N_5250,N_4887,N_4024);
and U5251 (N_5251,N_4483,N_4697);
nor U5252 (N_5252,N_4966,N_4992);
nand U5253 (N_5253,N_4962,N_4808);
xor U5254 (N_5254,N_4596,N_4260);
and U5255 (N_5255,N_4035,N_4003);
nor U5256 (N_5256,N_4274,N_4862);
or U5257 (N_5257,N_4819,N_4926);
and U5258 (N_5258,N_4601,N_4286);
nor U5259 (N_5259,N_4873,N_4755);
nand U5260 (N_5260,N_4389,N_4222);
xor U5261 (N_5261,N_4433,N_4461);
nand U5262 (N_5262,N_4592,N_4337);
nand U5263 (N_5263,N_4496,N_4728);
nor U5264 (N_5264,N_4948,N_4418);
xnor U5265 (N_5265,N_4191,N_4684);
and U5266 (N_5266,N_4336,N_4882);
nor U5267 (N_5267,N_4206,N_4416);
nor U5268 (N_5268,N_4692,N_4225);
nand U5269 (N_5269,N_4847,N_4304);
or U5270 (N_5270,N_4019,N_4886);
and U5271 (N_5271,N_4036,N_4838);
nor U5272 (N_5272,N_4980,N_4573);
or U5273 (N_5273,N_4691,N_4387);
nand U5274 (N_5274,N_4339,N_4109);
xor U5275 (N_5275,N_4317,N_4063);
and U5276 (N_5276,N_4910,N_4140);
and U5277 (N_5277,N_4480,N_4486);
or U5278 (N_5278,N_4265,N_4845);
and U5279 (N_5279,N_4752,N_4558);
nand U5280 (N_5280,N_4170,N_4804);
and U5281 (N_5281,N_4438,N_4922);
and U5282 (N_5282,N_4128,N_4588);
nor U5283 (N_5283,N_4916,N_4737);
xor U5284 (N_5284,N_4786,N_4780);
and U5285 (N_5285,N_4912,N_4246);
xor U5286 (N_5286,N_4428,N_4435);
xnor U5287 (N_5287,N_4401,N_4395);
and U5288 (N_5288,N_4991,N_4625);
and U5289 (N_5289,N_4082,N_4997);
and U5290 (N_5290,N_4323,N_4350);
nor U5291 (N_5291,N_4042,N_4959);
nor U5292 (N_5292,N_4799,N_4660);
nand U5293 (N_5293,N_4062,N_4826);
or U5294 (N_5294,N_4245,N_4456);
and U5295 (N_5295,N_4134,N_4789);
nor U5296 (N_5296,N_4133,N_4551);
xor U5297 (N_5297,N_4055,N_4890);
or U5298 (N_5298,N_4465,N_4528);
xnor U5299 (N_5299,N_4087,N_4296);
nand U5300 (N_5300,N_4023,N_4213);
and U5301 (N_5301,N_4067,N_4782);
nand U5302 (N_5302,N_4642,N_4044);
and U5303 (N_5303,N_4102,N_4054);
or U5304 (N_5304,N_4280,N_4584);
nor U5305 (N_5305,N_4995,N_4870);
or U5306 (N_5306,N_4930,N_4987);
nand U5307 (N_5307,N_4759,N_4587);
and U5308 (N_5308,N_4567,N_4711);
nand U5309 (N_5309,N_4240,N_4571);
and U5310 (N_5310,N_4020,N_4193);
or U5311 (N_5311,N_4079,N_4726);
nor U5312 (N_5312,N_4655,N_4150);
nor U5313 (N_5313,N_4520,N_4201);
nor U5314 (N_5314,N_4970,N_4275);
nand U5315 (N_5315,N_4667,N_4993);
nor U5316 (N_5316,N_4462,N_4220);
nor U5317 (N_5317,N_4276,N_4148);
or U5318 (N_5318,N_4255,N_4233);
or U5319 (N_5319,N_4219,N_4548);
nor U5320 (N_5320,N_4169,N_4457);
nor U5321 (N_5321,N_4717,N_4863);
xnor U5322 (N_5322,N_4907,N_4816);
nand U5323 (N_5323,N_4652,N_4132);
nor U5324 (N_5324,N_4268,N_4425);
xnor U5325 (N_5325,N_4982,N_4311);
xor U5326 (N_5326,N_4157,N_4796);
nand U5327 (N_5327,N_4544,N_4525);
xnor U5328 (N_5328,N_4161,N_4894);
and U5329 (N_5329,N_4287,N_4290);
nand U5330 (N_5330,N_4383,N_4139);
xor U5331 (N_5331,N_4351,N_4609);
nor U5332 (N_5332,N_4700,N_4162);
nand U5333 (N_5333,N_4393,N_4637);
nand U5334 (N_5334,N_4564,N_4867);
and U5335 (N_5335,N_4000,N_4852);
and U5336 (N_5336,N_4011,N_4630);
and U5337 (N_5337,N_4523,N_4569);
xor U5338 (N_5338,N_4578,N_4927);
nor U5339 (N_5339,N_4651,N_4756);
and U5340 (N_5340,N_4953,N_4214);
or U5341 (N_5341,N_4731,N_4634);
nor U5342 (N_5342,N_4294,N_4099);
nor U5343 (N_5343,N_4568,N_4763);
and U5344 (N_5344,N_4176,N_4197);
nor U5345 (N_5345,N_4324,N_4713);
or U5346 (N_5346,N_4724,N_4491);
and U5347 (N_5347,N_4076,N_4977);
or U5348 (N_5348,N_4898,N_4748);
or U5349 (N_5349,N_4621,N_4289);
xor U5350 (N_5350,N_4529,N_4022);
nand U5351 (N_5351,N_4757,N_4745);
nor U5352 (N_5352,N_4009,N_4954);
and U5353 (N_5353,N_4270,N_4037);
or U5354 (N_5354,N_4733,N_4141);
or U5355 (N_5355,N_4367,N_4404);
or U5356 (N_5356,N_4236,N_4595);
nand U5357 (N_5357,N_4888,N_4163);
nor U5358 (N_5358,N_4380,N_4627);
nand U5359 (N_5359,N_4762,N_4468);
nand U5360 (N_5360,N_4313,N_4061);
nor U5361 (N_5361,N_4398,N_4784);
and U5362 (N_5362,N_4071,N_4561);
nor U5363 (N_5363,N_4979,N_4840);
nor U5364 (N_5364,N_4537,N_4707);
nor U5365 (N_5365,N_4583,N_4566);
nand U5366 (N_5366,N_4407,N_4196);
or U5367 (N_5367,N_4409,N_4272);
or U5368 (N_5368,N_4326,N_4872);
xnor U5369 (N_5369,N_4923,N_4783);
nor U5370 (N_5370,N_4164,N_4250);
nand U5371 (N_5371,N_4443,N_4241);
xnor U5372 (N_5372,N_4088,N_4526);
and U5373 (N_5373,N_4065,N_4597);
xor U5374 (N_5374,N_4403,N_4539);
xnor U5375 (N_5375,N_4790,N_4205);
xor U5376 (N_5376,N_4952,N_4239);
nor U5377 (N_5377,N_4001,N_4946);
or U5378 (N_5378,N_4895,N_4248);
nand U5379 (N_5379,N_4185,N_4303);
nand U5380 (N_5380,N_4069,N_4188);
nor U5381 (N_5381,N_4617,N_4649);
and U5382 (N_5382,N_4643,N_4703);
or U5383 (N_5383,N_4033,N_4612);
nor U5384 (N_5384,N_4459,N_4603);
xnor U5385 (N_5385,N_4116,N_4358);
or U5386 (N_5386,N_4859,N_4130);
and U5387 (N_5387,N_4904,N_4232);
nor U5388 (N_5388,N_4186,N_4208);
or U5389 (N_5389,N_4346,N_4680);
and U5390 (N_5390,N_4961,N_4635);
nor U5391 (N_5391,N_4751,N_4293);
and U5392 (N_5392,N_4347,N_4470);
and U5393 (N_5393,N_4579,N_4357);
xnor U5394 (N_5394,N_4559,N_4856);
or U5395 (N_5395,N_4512,N_4155);
or U5396 (N_5396,N_4064,N_4234);
and U5397 (N_5397,N_4254,N_4541);
xnor U5398 (N_5398,N_4298,N_4056);
nand U5399 (N_5399,N_4123,N_4880);
nand U5400 (N_5400,N_4321,N_4805);
and U5401 (N_5401,N_4143,N_4308);
nand U5402 (N_5402,N_4532,N_4960);
and U5403 (N_5403,N_4440,N_4725);
and U5404 (N_5404,N_4080,N_4905);
xor U5405 (N_5405,N_4200,N_4556);
xnor U5406 (N_5406,N_4333,N_4741);
xnor U5407 (N_5407,N_4482,N_4167);
xor U5408 (N_5408,N_4549,N_4442);
xnor U5409 (N_5409,N_4942,N_4177);
or U5410 (N_5410,N_4066,N_4851);
nor U5411 (N_5411,N_4604,N_4944);
or U5412 (N_5412,N_4903,N_4106);
nand U5413 (N_5413,N_4291,N_4273);
nor U5414 (N_5414,N_4855,N_4158);
nor U5415 (N_5415,N_4547,N_4913);
xnor U5416 (N_5416,N_4021,N_4978);
xnor U5417 (N_5417,N_4839,N_4343);
nor U5418 (N_5418,N_4914,N_4983);
or U5419 (N_5419,N_4413,N_4320);
or U5420 (N_5420,N_4312,N_4674);
xnor U5421 (N_5421,N_4996,N_4721);
nor U5422 (N_5422,N_4694,N_4610);
nand U5423 (N_5423,N_4770,N_4896);
and U5424 (N_5424,N_4227,N_4392);
and U5425 (N_5425,N_4372,N_4183);
or U5426 (N_5426,N_4049,N_4647);
xnor U5427 (N_5427,N_4956,N_4574);
and U5428 (N_5428,N_4554,N_4364);
nand U5429 (N_5429,N_4192,N_4727);
nand U5430 (N_5430,N_4181,N_4485);
or U5431 (N_5431,N_4823,N_4251);
nand U5432 (N_5432,N_4105,N_4753);
nand U5433 (N_5433,N_4791,N_4683);
or U5434 (N_5434,N_4100,N_4619);
nor U5435 (N_5435,N_4675,N_4315);
and U5436 (N_5436,N_4349,N_4224);
and U5437 (N_5437,N_4096,N_4285);
xor U5438 (N_5438,N_4144,N_4190);
nand U5439 (N_5439,N_4747,N_4467);
nand U5440 (N_5440,N_4497,N_4405);
nand U5441 (N_5441,N_4345,N_4628);
xnor U5442 (N_5442,N_4534,N_4352);
nand U5443 (N_5443,N_4943,N_4125);
or U5444 (N_5444,N_4538,N_4002);
and U5445 (N_5445,N_4650,N_4237);
xnor U5446 (N_5446,N_4576,N_4810);
or U5447 (N_5447,N_4572,N_4264);
nand U5448 (N_5448,N_4885,N_4735);
xnor U5449 (N_5449,N_4902,N_4705);
and U5450 (N_5450,N_4436,N_4252);
nand U5451 (N_5451,N_4932,N_4502);
nor U5452 (N_5452,N_4469,N_4421);
or U5453 (N_5453,N_4563,N_4714);
and U5454 (N_5454,N_4362,N_4580);
or U5455 (N_5455,N_4175,N_4307);
or U5456 (N_5456,N_4765,N_4669);
nand U5457 (N_5457,N_4154,N_4722);
xnor U5458 (N_5458,N_4202,N_4656);
nor U5459 (N_5459,N_4318,N_4900);
and U5460 (N_5460,N_4355,N_4920);
or U5461 (N_5461,N_4194,N_4156);
nor U5462 (N_5462,N_4820,N_4844);
xnor U5463 (N_5463,N_4050,N_4984);
nor U5464 (N_5464,N_4335,N_4007);
nor U5465 (N_5465,N_4012,N_4586);
nand U5466 (N_5466,N_4504,N_4195);
nand U5467 (N_5467,N_4869,N_4084);
nor U5468 (N_5468,N_4518,N_4876);
nand U5469 (N_5469,N_4822,N_4835);
and U5470 (N_5470,N_4390,N_4800);
nand U5471 (N_5471,N_4963,N_4391);
xnor U5472 (N_5472,N_4915,N_4008);
nand U5473 (N_5473,N_4415,N_4400);
or U5474 (N_5474,N_4941,N_4552);
nand U5475 (N_5475,N_4094,N_4623);
xor U5476 (N_5476,N_4017,N_4451);
nor U5477 (N_5477,N_4058,N_4767);
and U5478 (N_5478,N_4990,N_4487);
and U5479 (N_5479,N_4965,N_4137);
or U5480 (N_5480,N_4478,N_4850);
or U5481 (N_5481,N_4702,N_4657);
and U5482 (N_5482,N_4513,N_4560);
or U5483 (N_5483,N_4305,N_4884);
and U5484 (N_5484,N_4989,N_4773);
or U5485 (N_5485,N_4719,N_4278);
nand U5486 (N_5486,N_4654,N_4430);
xor U5487 (N_5487,N_4074,N_4452);
and U5488 (N_5488,N_4242,N_4327);
nor U5489 (N_5489,N_4837,N_4797);
xnor U5490 (N_5490,N_4677,N_4938);
xor U5491 (N_5491,N_4866,N_4247);
and U5492 (N_5492,N_4348,N_4524);
and U5493 (N_5493,N_4533,N_4682);
nand U5494 (N_5494,N_4243,N_4766);
nor U5495 (N_5495,N_4455,N_4373);
xnor U5496 (N_5496,N_4228,N_4101);
or U5497 (N_5497,N_4598,N_4830);
and U5498 (N_5498,N_4740,N_4928);
nand U5499 (N_5499,N_4238,N_4743);
or U5500 (N_5500,N_4463,N_4712);
or U5501 (N_5501,N_4513,N_4614);
or U5502 (N_5502,N_4271,N_4155);
or U5503 (N_5503,N_4316,N_4910);
or U5504 (N_5504,N_4256,N_4789);
nand U5505 (N_5505,N_4838,N_4852);
nor U5506 (N_5506,N_4525,N_4005);
nand U5507 (N_5507,N_4035,N_4297);
nor U5508 (N_5508,N_4173,N_4910);
xnor U5509 (N_5509,N_4929,N_4637);
xor U5510 (N_5510,N_4497,N_4702);
or U5511 (N_5511,N_4123,N_4158);
and U5512 (N_5512,N_4364,N_4136);
xnor U5513 (N_5513,N_4649,N_4476);
xor U5514 (N_5514,N_4585,N_4965);
nand U5515 (N_5515,N_4375,N_4197);
xor U5516 (N_5516,N_4722,N_4993);
xnor U5517 (N_5517,N_4696,N_4929);
nand U5518 (N_5518,N_4766,N_4257);
nor U5519 (N_5519,N_4543,N_4126);
xnor U5520 (N_5520,N_4284,N_4547);
or U5521 (N_5521,N_4627,N_4224);
xor U5522 (N_5522,N_4582,N_4808);
and U5523 (N_5523,N_4137,N_4638);
nor U5524 (N_5524,N_4542,N_4042);
or U5525 (N_5525,N_4958,N_4999);
or U5526 (N_5526,N_4606,N_4749);
and U5527 (N_5527,N_4216,N_4553);
or U5528 (N_5528,N_4274,N_4391);
and U5529 (N_5529,N_4959,N_4691);
nor U5530 (N_5530,N_4940,N_4460);
and U5531 (N_5531,N_4185,N_4422);
or U5532 (N_5532,N_4830,N_4784);
nor U5533 (N_5533,N_4742,N_4421);
xor U5534 (N_5534,N_4073,N_4876);
or U5535 (N_5535,N_4259,N_4760);
nand U5536 (N_5536,N_4038,N_4923);
xnor U5537 (N_5537,N_4150,N_4279);
and U5538 (N_5538,N_4227,N_4366);
or U5539 (N_5539,N_4137,N_4087);
or U5540 (N_5540,N_4516,N_4632);
nand U5541 (N_5541,N_4464,N_4889);
nand U5542 (N_5542,N_4615,N_4345);
or U5543 (N_5543,N_4600,N_4847);
and U5544 (N_5544,N_4919,N_4499);
and U5545 (N_5545,N_4658,N_4945);
xor U5546 (N_5546,N_4007,N_4597);
nor U5547 (N_5547,N_4214,N_4375);
nor U5548 (N_5548,N_4318,N_4130);
or U5549 (N_5549,N_4782,N_4197);
xnor U5550 (N_5550,N_4167,N_4453);
nand U5551 (N_5551,N_4925,N_4381);
and U5552 (N_5552,N_4725,N_4972);
nand U5553 (N_5553,N_4057,N_4649);
nor U5554 (N_5554,N_4548,N_4687);
and U5555 (N_5555,N_4505,N_4343);
xnor U5556 (N_5556,N_4378,N_4821);
and U5557 (N_5557,N_4207,N_4130);
nor U5558 (N_5558,N_4386,N_4653);
nor U5559 (N_5559,N_4414,N_4973);
or U5560 (N_5560,N_4400,N_4797);
nand U5561 (N_5561,N_4510,N_4249);
xor U5562 (N_5562,N_4916,N_4609);
and U5563 (N_5563,N_4711,N_4267);
nor U5564 (N_5564,N_4981,N_4876);
xnor U5565 (N_5565,N_4803,N_4642);
and U5566 (N_5566,N_4958,N_4844);
or U5567 (N_5567,N_4892,N_4324);
nor U5568 (N_5568,N_4849,N_4167);
and U5569 (N_5569,N_4663,N_4036);
xnor U5570 (N_5570,N_4510,N_4204);
xnor U5571 (N_5571,N_4137,N_4356);
and U5572 (N_5572,N_4291,N_4896);
nand U5573 (N_5573,N_4210,N_4080);
xnor U5574 (N_5574,N_4186,N_4171);
xnor U5575 (N_5575,N_4286,N_4464);
nand U5576 (N_5576,N_4795,N_4520);
xnor U5577 (N_5577,N_4071,N_4773);
or U5578 (N_5578,N_4247,N_4577);
or U5579 (N_5579,N_4868,N_4331);
and U5580 (N_5580,N_4961,N_4107);
nor U5581 (N_5581,N_4907,N_4719);
and U5582 (N_5582,N_4339,N_4411);
xor U5583 (N_5583,N_4955,N_4787);
xnor U5584 (N_5584,N_4361,N_4836);
nand U5585 (N_5585,N_4985,N_4450);
nor U5586 (N_5586,N_4587,N_4574);
nor U5587 (N_5587,N_4158,N_4307);
xor U5588 (N_5588,N_4396,N_4326);
nand U5589 (N_5589,N_4756,N_4455);
nand U5590 (N_5590,N_4335,N_4853);
and U5591 (N_5591,N_4662,N_4526);
or U5592 (N_5592,N_4147,N_4308);
or U5593 (N_5593,N_4366,N_4961);
nor U5594 (N_5594,N_4050,N_4063);
xnor U5595 (N_5595,N_4860,N_4018);
xor U5596 (N_5596,N_4402,N_4157);
nand U5597 (N_5597,N_4619,N_4889);
nor U5598 (N_5598,N_4845,N_4843);
nand U5599 (N_5599,N_4172,N_4391);
or U5600 (N_5600,N_4894,N_4041);
nand U5601 (N_5601,N_4245,N_4151);
nand U5602 (N_5602,N_4003,N_4946);
or U5603 (N_5603,N_4211,N_4334);
or U5604 (N_5604,N_4510,N_4456);
and U5605 (N_5605,N_4929,N_4239);
and U5606 (N_5606,N_4008,N_4180);
or U5607 (N_5607,N_4753,N_4320);
and U5608 (N_5608,N_4692,N_4752);
or U5609 (N_5609,N_4371,N_4225);
xnor U5610 (N_5610,N_4367,N_4183);
nor U5611 (N_5611,N_4790,N_4965);
xnor U5612 (N_5612,N_4042,N_4043);
and U5613 (N_5613,N_4538,N_4625);
xnor U5614 (N_5614,N_4875,N_4125);
nor U5615 (N_5615,N_4383,N_4336);
or U5616 (N_5616,N_4134,N_4731);
and U5617 (N_5617,N_4396,N_4425);
and U5618 (N_5618,N_4273,N_4332);
and U5619 (N_5619,N_4524,N_4929);
and U5620 (N_5620,N_4397,N_4064);
or U5621 (N_5621,N_4227,N_4554);
or U5622 (N_5622,N_4955,N_4965);
nor U5623 (N_5623,N_4089,N_4973);
nand U5624 (N_5624,N_4727,N_4415);
and U5625 (N_5625,N_4739,N_4844);
xor U5626 (N_5626,N_4269,N_4867);
and U5627 (N_5627,N_4438,N_4533);
nor U5628 (N_5628,N_4323,N_4769);
or U5629 (N_5629,N_4850,N_4504);
xnor U5630 (N_5630,N_4767,N_4370);
nor U5631 (N_5631,N_4351,N_4489);
xnor U5632 (N_5632,N_4311,N_4737);
or U5633 (N_5633,N_4716,N_4361);
and U5634 (N_5634,N_4982,N_4261);
xnor U5635 (N_5635,N_4240,N_4263);
nand U5636 (N_5636,N_4935,N_4355);
nand U5637 (N_5637,N_4159,N_4268);
nand U5638 (N_5638,N_4422,N_4170);
xnor U5639 (N_5639,N_4050,N_4205);
nor U5640 (N_5640,N_4511,N_4220);
or U5641 (N_5641,N_4230,N_4049);
xor U5642 (N_5642,N_4824,N_4170);
or U5643 (N_5643,N_4340,N_4410);
or U5644 (N_5644,N_4889,N_4120);
nor U5645 (N_5645,N_4640,N_4672);
or U5646 (N_5646,N_4621,N_4555);
and U5647 (N_5647,N_4864,N_4938);
nand U5648 (N_5648,N_4085,N_4293);
nand U5649 (N_5649,N_4247,N_4287);
nor U5650 (N_5650,N_4179,N_4642);
and U5651 (N_5651,N_4737,N_4156);
and U5652 (N_5652,N_4758,N_4605);
xor U5653 (N_5653,N_4118,N_4673);
nor U5654 (N_5654,N_4253,N_4394);
nor U5655 (N_5655,N_4661,N_4632);
and U5656 (N_5656,N_4459,N_4149);
or U5657 (N_5657,N_4903,N_4328);
and U5658 (N_5658,N_4002,N_4368);
or U5659 (N_5659,N_4924,N_4240);
or U5660 (N_5660,N_4029,N_4755);
and U5661 (N_5661,N_4674,N_4990);
xor U5662 (N_5662,N_4079,N_4978);
or U5663 (N_5663,N_4802,N_4212);
and U5664 (N_5664,N_4067,N_4049);
nor U5665 (N_5665,N_4281,N_4138);
nor U5666 (N_5666,N_4352,N_4300);
or U5667 (N_5667,N_4357,N_4832);
and U5668 (N_5668,N_4090,N_4164);
and U5669 (N_5669,N_4171,N_4978);
and U5670 (N_5670,N_4911,N_4860);
nand U5671 (N_5671,N_4972,N_4728);
nor U5672 (N_5672,N_4104,N_4202);
nand U5673 (N_5673,N_4572,N_4893);
nand U5674 (N_5674,N_4759,N_4082);
nor U5675 (N_5675,N_4288,N_4546);
xor U5676 (N_5676,N_4173,N_4105);
and U5677 (N_5677,N_4530,N_4561);
xor U5678 (N_5678,N_4351,N_4682);
xnor U5679 (N_5679,N_4107,N_4276);
nor U5680 (N_5680,N_4694,N_4361);
and U5681 (N_5681,N_4964,N_4423);
and U5682 (N_5682,N_4505,N_4356);
or U5683 (N_5683,N_4540,N_4718);
nor U5684 (N_5684,N_4387,N_4175);
nor U5685 (N_5685,N_4648,N_4441);
nor U5686 (N_5686,N_4891,N_4622);
xnor U5687 (N_5687,N_4077,N_4545);
nand U5688 (N_5688,N_4876,N_4688);
nand U5689 (N_5689,N_4488,N_4042);
nor U5690 (N_5690,N_4836,N_4662);
xnor U5691 (N_5691,N_4472,N_4841);
or U5692 (N_5692,N_4944,N_4654);
xnor U5693 (N_5693,N_4101,N_4100);
and U5694 (N_5694,N_4802,N_4466);
and U5695 (N_5695,N_4995,N_4177);
or U5696 (N_5696,N_4803,N_4196);
or U5697 (N_5697,N_4175,N_4932);
xor U5698 (N_5698,N_4444,N_4220);
nor U5699 (N_5699,N_4812,N_4865);
and U5700 (N_5700,N_4816,N_4163);
nor U5701 (N_5701,N_4029,N_4593);
and U5702 (N_5702,N_4349,N_4918);
or U5703 (N_5703,N_4142,N_4029);
or U5704 (N_5704,N_4477,N_4116);
xnor U5705 (N_5705,N_4298,N_4019);
and U5706 (N_5706,N_4647,N_4803);
nand U5707 (N_5707,N_4841,N_4354);
or U5708 (N_5708,N_4905,N_4893);
xor U5709 (N_5709,N_4465,N_4288);
nor U5710 (N_5710,N_4431,N_4493);
and U5711 (N_5711,N_4375,N_4866);
or U5712 (N_5712,N_4335,N_4487);
xor U5713 (N_5713,N_4735,N_4757);
and U5714 (N_5714,N_4647,N_4318);
xnor U5715 (N_5715,N_4183,N_4055);
nand U5716 (N_5716,N_4088,N_4197);
nand U5717 (N_5717,N_4670,N_4019);
or U5718 (N_5718,N_4031,N_4758);
nor U5719 (N_5719,N_4532,N_4941);
xor U5720 (N_5720,N_4409,N_4022);
xnor U5721 (N_5721,N_4332,N_4846);
nor U5722 (N_5722,N_4471,N_4637);
and U5723 (N_5723,N_4959,N_4069);
and U5724 (N_5724,N_4943,N_4401);
or U5725 (N_5725,N_4501,N_4247);
xor U5726 (N_5726,N_4808,N_4568);
xnor U5727 (N_5727,N_4886,N_4662);
or U5728 (N_5728,N_4146,N_4313);
or U5729 (N_5729,N_4543,N_4071);
nor U5730 (N_5730,N_4306,N_4123);
or U5731 (N_5731,N_4051,N_4210);
xnor U5732 (N_5732,N_4704,N_4439);
and U5733 (N_5733,N_4287,N_4099);
or U5734 (N_5734,N_4820,N_4483);
nor U5735 (N_5735,N_4210,N_4776);
xor U5736 (N_5736,N_4045,N_4700);
or U5737 (N_5737,N_4907,N_4002);
xnor U5738 (N_5738,N_4149,N_4030);
xor U5739 (N_5739,N_4489,N_4736);
and U5740 (N_5740,N_4353,N_4596);
or U5741 (N_5741,N_4386,N_4122);
xor U5742 (N_5742,N_4658,N_4938);
or U5743 (N_5743,N_4585,N_4785);
xor U5744 (N_5744,N_4957,N_4237);
xor U5745 (N_5745,N_4203,N_4581);
or U5746 (N_5746,N_4780,N_4468);
xnor U5747 (N_5747,N_4008,N_4510);
or U5748 (N_5748,N_4151,N_4993);
and U5749 (N_5749,N_4706,N_4722);
nor U5750 (N_5750,N_4553,N_4071);
and U5751 (N_5751,N_4603,N_4567);
or U5752 (N_5752,N_4274,N_4460);
nor U5753 (N_5753,N_4542,N_4868);
xor U5754 (N_5754,N_4923,N_4645);
or U5755 (N_5755,N_4490,N_4559);
xor U5756 (N_5756,N_4663,N_4735);
and U5757 (N_5757,N_4294,N_4394);
nor U5758 (N_5758,N_4292,N_4516);
nor U5759 (N_5759,N_4791,N_4180);
and U5760 (N_5760,N_4918,N_4729);
nor U5761 (N_5761,N_4336,N_4897);
xnor U5762 (N_5762,N_4721,N_4890);
and U5763 (N_5763,N_4767,N_4904);
and U5764 (N_5764,N_4465,N_4998);
xor U5765 (N_5765,N_4006,N_4125);
nand U5766 (N_5766,N_4867,N_4790);
nor U5767 (N_5767,N_4739,N_4165);
nand U5768 (N_5768,N_4917,N_4911);
or U5769 (N_5769,N_4724,N_4599);
or U5770 (N_5770,N_4626,N_4304);
and U5771 (N_5771,N_4650,N_4895);
and U5772 (N_5772,N_4320,N_4670);
nor U5773 (N_5773,N_4361,N_4610);
or U5774 (N_5774,N_4322,N_4086);
nand U5775 (N_5775,N_4319,N_4349);
nor U5776 (N_5776,N_4880,N_4514);
nor U5777 (N_5777,N_4370,N_4371);
or U5778 (N_5778,N_4878,N_4377);
and U5779 (N_5779,N_4049,N_4254);
nor U5780 (N_5780,N_4650,N_4911);
nor U5781 (N_5781,N_4046,N_4795);
nor U5782 (N_5782,N_4408,N_4346);
or U5783 (N_5783,N_4153,N_4323);
xnor U5784 (N_5784,N_4789,N_4552);
xnor U5785 (N_5785,N_4793,N_4254);
xnor U5786 (N_5786,N_4497,N_4083);
and U5787 (N_5787,N_4653,N_4203);
xnor U5788 (N_5788,N_4338,N_4914);
nand U5789 (N_5789,N_4335,N_4684);
nor U5790 (N_5790,N_4487,N_4896);
nor U5791 (N_5791,N_4774,N_4132);
xor U5792 (N_5792,N_4090,N_4820);
nor U5793 (N_5793,N_4547,N_4575);
xor U5794 (N_5794,N_4103,N_4216);
nand U5795 (N_5795,N_4078,N_4915);
or U5796 (N_5796,N_4424,N_4910);
nand U5797 (N_5797,N_4158,N_4441);
nand U5798 (N_5798,N_4086,N_4227);
or U5799 (N_5799,N_4868,N_4696);
nor U5800 (N_5800,N_4308,N_4036);
nand U5801 (N_5801,N_4316,N_4124);
nor U5802 (N_5802,N_4118,N_4068);
nor U5803 (N_5803,N_4641,N_4211);
and U5804 (N_5804,N_4904,N_4839);
or U5805 (N_5805,N_4129,N_4757);
or U5806 (N_5806,N_4123,N_4339);
nand U5807 (N_5807,N_4956,N_4373);
or U5808 (N_5808,N_4284,N_4781);
xor U5809 (N_5809,N_4662,N_4923);
or U5810 (N_5810,N_4748,N_4993);
xnor U5811 (N_5811,N_4378,N_4256);
nand U5812 (N_5812,N_4016,N_4068);
or U5813 (N_5813,N_4071,N_4221);
or U5814 (N_5814,N_4505,N_4322);
and U5815 (N_5815,N_4727,N_4990);
nand U5816 (N_5816,N_4609,N_4983);
and U5817 (N_5817,N_4791,N_4042);
nor U5818 (N_5818,N_4757,N_4783);
nor U5819 (N_5819,N_4105,N_4548);
nand U5820 (N_5820,N_4399,N_4778);
nand U5821 (N_5821,N_4959,N_4338);
nor U5822 (N_5822,N_4305,N_4714);
nand U5823 (N_5823,N_4665,N_4269);
nor U5824 (N_5824,N_4588,N_4229);
and U5825 (N_5825,N_4070,N_4361);
xnor U5826 (N_5826,N_4966,N_4186);
xor U5827 (N_5827,N_4552,N_4710);
nand U5828 (N_5828,N_4658,N_4139);
nand U5829 (N_5829,N_4167,N_4360);
xnor U5830 (N_5830,N_4861,N_4757);
or U5831 (N_5831,N_4871,N_4045);
and U5832 (N_5832,N_4913,N_4077);
and U5833 (N_5833,N_4726,N_4514);
nand U5834 (N_5834,N_4360,N_4345);
and U5835 (N_5835,N_4217,N_4195);
xor U5836 (N_5836,N_4289,N_4247);
xnor U5837 (N_5837,N_4827,N_4834);
and U5838 (N_5838,N_4650,N_4280);
xor U5839 (N_5839,N_4393,N_4381);
and U5840 (N_5840,N_4352,N_4740);
and U5841 (N_5841,N_4976,N_4231);
xnor U5842 (N_5842,N_4564,N_4323);
and U5843 (N_5843,N_4560,N_4282);
xnor U5844 (N_5844,N_4779,N_4840);
nor U5845 (N_5845,N_4943,N_4452);
and U5846 (N_5846,N_4801,N_4965);
or U5847 (N_5847,N_4113,N_4613);
nand U5848 (N_5848,N_4068,N_4555);
nor U5849 (N_5849,N_4464,N_4332);
or U5850 (N_5850,N_4693,N_4819);
and U5851 (N_5851,N_4440,N_4803);
or U5852 (N_5852,N_4042,N_4684);
nor U5853 (N_5853,N_4708,N_4707);
or U5854 (N_5854,N_4509,N_4193);
or U5855 (N_5855,N_4590,N_4696);
nand U5856 (N_5856,N_4302,N_4459);
xor U5857 (N_5857,N_4539,N_4713);
xor U5858 (N_5858,N_4405,N_4502);
nor U5859 (N_5859,N_4354,N_4082);
and U5860 (N_5860,N_4515,N_4941);
xnor U5861 (N_5861,N_4765,N_4285);
xor U5862 (N_5862,N_4875,N_4873);
and U5863 (N_5863,N_4117,N_4779);
and U5864 (N_5864,N_4764,N_4170);
and U5865 (N_5865,N_4814,N_4666);
and U5866 (N_5866,N_4300,N_4531);
xor U5867 (N_5867,N_4546,N_4315);
nor U5868 (N_5868,N_4791,N_4704);
nor U5869 (N_5869,N_4748,N_4740);
xor U5870 (N_5870,N_4173,N_4439);
and U5871 (N_5871,N_4548,N_4959);
xnor U5872 (N_5872,N_4851,N_4210);
nor U5873 (N_5873,N_4088,N_4816);
nor U5874 (N_5874,N_4910,N_4990);
and U5875 (N_5875,N_4136,N_4240);
nand U5876 (N_5876,N_4965,N_4185);
nand U5877 (N_5877,N_4640,N_4741);
xnor U5878 (N_5878,N_4267,N_4748);
and U5879 (N_5879,N_4570,N_4561);
xor U5880 (N_5880,N_4114,N_4654);
and U5881 (N_5881,N_4269,N_4427);
and U5882 (N_5882,N_4468,N_4305);
xnor U5883 (N_5883,N_4682,N_4110);
xor U5884 (N_5884,N_4097,N_4492);
nor U5885 (N_5885,N_4129,N_4178);
and U5886 (N_5886,N_4828,N_4780);
xor U5887 (N_5887,N_4664,N_4120);
or U5888 (N_5888,N_4010,N_4424);
nor U5889 (N_5889,N_4679,N_4399);
nand U5890 (N_5890,N_4894,N_4824);
nor U5891 (N_5891,N_4056,N_4970);
nand U5892 (N_5892,N_4012,N_4378);
nand U5893 (N_5893,N_4707,N_4038);
nand U5894 (N_5894,N_4398,N_4495);
or U5895 (N_5895,N_4309,N_4557);
or U5896 (N_5896,N_4464,N_4424);
nor U5897 (N_5897,N_4436,N_4565);
and U5898 (N_5898,N_4048,N_4140);
nand U5899 (N_5899,N_4516,N_4237);
nand U5900 (N_5900,N_4821,N_4854);
nor U5901 (N_5901,N_4773,N_4586);
and U5902 (N_5902,N_4753,N_4856);
nand U5903 (N_5903,N_4009,N_4761);
nand U5904 (N_5904,N_4685,N_4768);
nand U5905 (N_5905,N_4338,N_4664);
nand U5906 (N_5906,N_4739,N_4113);
nand U5907 (N_5907,N_4048,N_4388);
xnor U5908 (N_5908,N_4909,N_4033);
nand U5909 (N_5909,N_4181,N_4944);
nor U5910 (N_5910,N_4938,N_4720);
xor U5911 (N_5911,N_4180,N_4016);
xor U5912 (N_5912,N_4966,N_4830);
nor U5913 (N_5913,N_4840,N_4781);
nor U5914 (N_5914,N_4062,N_4718);
xnor U5915 (N_5915,N_4305,N_4115);
nand U5916 (N_5916,N_4552,N_4413);
nand U5917 (N_5917,N_4889,N_4772);
and U5918 (N_5918,N_4414,N_4912);
nor U5919 (N_5919,N_4224,N_4375);
nand U5920 (N_5920,N_4012,N_4762);
nor U5921 (N_5921,N_4003,N_4602);
nand U5922 (N_5922,N_4426,N_4608);
and U5923 (N_5923,N_4909,N_4641);
or U5924 (N_5924,N_4481,N_4355);
or U5925 (N_5925,N_4777,N_4122);
nor U5926 (N_5926,N_4076,N_4345);
and U5927 (N_5927,N_4811,N_4903);
and U5928 (N_5928,N_4709,N_4343);
or U5929 (N_5929,N_4372,N_4276);
xor U5930 (N_5930,N_4235,N_4979);
or U5931 (N_5931,N_4907,N_4495);
nand U5932 (N_5932,N_4915,N_4464);
or U5933 (N_5933,N_4603,N_4082);
and U5934 (N_5934,N_4633,N_4675);
nor U5935 (N_5935,N_4769,N_4060);
or U5936 (N_5936,N_4514,N_4600);
nand U5937 (N_5937,N_4216,N_4210);
and U5938 (N_5938,N_4061,N_4947);
xor U5939 (N_5939,N_4379,N_4739);
and U5940 (N_5940,N_4633,N_4463);
xor U5941 (N_5941,N_4816,N_4599);
nor U5942 (N_5942,N_4592,N_4410);
and U5943 (N_5943,N_4915,N_4848);
nor U5944 (N_5944,N_4818,N_4095);
xnor U5945 (N_5945,N_4463,N_4977);
and U5946 (N_5946,N_4425,N_4286);
nand U5947 (N_5947,N_4777,N_4319);
nor U5948 (N_5948,N_4668,N_4681);
nor U5949 (N_5949,N_4529,N_4203);
xor U5950 (N_5950,N_4856,N_4068);
and U5951 (N_5951,N_4474,N_4152);
or U5952 (N_5952,N_4303,N_4903);
nand U5953 (N_5953,N_4827,N_4107);
nor U5954 (N_5954,N_4727,N_4480);
or U5955 (N_5955,N_4387,N_4564);
xnor U5956 (N_5956,N_4959,N_4169);
nand U5957 (N_5957,N_4457,N_4070);
xnor U5958 (N_5958,N_4639,N_4326);
nor U5959 (N_5959,N_4306,N_4662);
nor U5960 (N_5960,N_4540,N_4873);
nor U5961 (N_5961,N_4744,N_4742);
xor U5962 (N_5962,N_4664,N_4226);
or U5963 (N_5963,N_4833,N_4491);
and U5964 (N_5964,N_4662,N_4204);
xor U5965 (N_5965,N_4939,N_4618);
and U5966 (N_5966,N_4005,N_4739);
xnor U5967 (N_5967,N_4380,N_4083);
and U5968 (N_5968,N_4629,N_4727);
or U5969 (N_5969,N_4721,N_4153);
and U5970 (N_5970,N_4305,N_4230);
nand U5971 (N_5971,N_4115,N_4297);
nand U5972 (N_5972,N_4619,N_4245);
nor U5973 (N_5973,N_4981,N_4821);
or U5974 (N_5974,N_4905,N_4977);
or U5975 (N_5975,N_4576,N_4138);
nand U5976 (N_5976,N_4500,N_4227);
or U5977 (N_5977,N_4330,N_4114);
xnor U5978 (N_5978,N_4653,N_4421);
nand U5979 (N_5979,N_4068,N_4735);
nor U5980 (N_5980,N_4692,N_4186);
xnor U5981 (N_5981,N_4885,N_4383);
nor U5982 (N_5982,N_4183,N_4245);
or U5983 (N_5983,N_4672,N_4015);
nand U5984 (N_5984,N_4669,N_4956);
xnor U5985 (N_5985,N_4060,N_4965);
nor U5986 (N_5986,N_4527,N_4946);
xor U5987 (N_5987,N_4655,N_4129);
or U5988 (N_5988,N_4025,N_4585);
nor U5989 (N_5989,N_4995,N_4496);
or U5990 (N_5990,N_4973,N_4208);
nand U5991 (N_5991,N_4728,N_4430);
nand U5992 (N_5992,N_4470,N_4273);
nand U5993 (N_5993,N_4353,N_4192);
xnor U5994 (N_5994,N_4904,N_4854);
nor U5995 (N_5995,N_4669,N_4110);
or U5996 (N_5996,N_4531,N_4839);
xor U5997 (N_5997,N_4266,N_4894);
nor U5998 (N_5998,N_4413,N_4004);
xnor U5999 (N_5999,N_4466,N_4765);
nand U6000 (N_6000,N_5869,N_5034);
or U6001 (N_6001,N_5752,N_5690);
nor U6002 (N_6002,N_5632,N_5358);
nand U6003 (N_6003,N_5853,N_5812);
xnor U6004 (N_6004,N_5930,N_5422);
xor U6005 (N_6005,N_5190,N_5597);
nor U6006 (N_6006,N_5113,N_5759);
and U6007 (N_6007,N_5010,N_5799);
nor U6008 (N_6008,N_5165,N_5865);
nand U6009 (N_6009,N_5757,N_5886);
xor U6010 (N_6010,N_5257,N_5827);
and U6011 (N_6011,N_5933,N_5687);
nand U6012 (N_6012,N_5565,N_5848);
or U6013 (N_6013,N_5161,N_5000);
xnor U6014 (N_6014,N_5919,N_5052);
xnor U6015 (N_6015,N_5800,N_5427);
nand U6016 (N_6016,N_5828,N_5809);
and U6017 (N_6017,N_5775,N_5735);
xor U6018 (N_6018,N_5247,N_5670);
nor U6019 (N_6019,N_5469,N_5328);
nor U6020 (N_6020,N_5350,N_5103);
nor U6021 (N_6021,N_5156,N_5850);
xnor U6022 (N_6022,N_5254,N_5645);
xnor U6023 (N_6023,N_5666,N_5399);
xor U6024 (N_6024,N_5763,N_5626);
and U6025 (N_6025,N_5734,N_5088);
and U6026 (N_6026,N_5346,N_5871);
xnor U6027 (N_6027,N_5798,N_5824);
nor U6028 (N_6028,N_5196,N_5563);
nand U6029 (N_6029,N_5635,N_5630);
or U6030 (N_6030,N_5599,N_5602);
nand U6031 (N_6031,N_5108,N_5045);
xor U6032 (N_6032,N_5104,N_5948);
and U6033 (N_6033,N_5888,N_5494);
or U6034 (N_6034,N_5406,N_5720);
nand U6035 (N_6035,N_5061,N_5875);
xor U6036 (N_6036,N_5892,N_5905);
and U6037 (N_6037,N_5958,N_5496);
nand U6038 (N_6038,N_5683,N_5056);
or U6039 (N_6039,N_5242,N_5130);
or U6040 (N_6040,N_5843,N_5992);
nor U6041 (N_6041,N_5898,N_5493);
and U6042 (N_6042,N_5213,N_5331);
nor U6043 (N_6043,N_5567,N_5319);
or U6044 (N_6044,N_5721,N_5530);
nor U6045 (N_6045,N_5259,N_5680);
nor U6046 (N_6046,N_5516,N_5437);
or U6047 (N_6047,N_5556,N_5162);
xor U6048 (N_6048,N_5481,N_5004);
or U6049 (N_6049,N_5068,N_5013);
xor U6050 (N_6050,N_5248,N_5194);
and U6051 (N_6051,N_5105,N_5694);
nor U6052 (N_6052,N_5455,N_5138);
nor U6053 (N_6053,N_5994,N_5750);
nand U6054 (N_6054,N_5911,N_5198);
nand U6055 (N_6055,N_5753,N_5758);
xor U6056 (N_6056,N_5250,N_5405);
xnor U6057 (N_6057,N_5560,N_5989);
nand U6058 (N_6058,N_5665,N_5701);
xor U6059 (N_6059,N_5795,N_5012);
nor U6060 (N_6060,N_5741,N_5927);
nor U6061 (N_6061,N_5803,N_5225);
xor U6062 (N_6062,N_5649,N_5745);
and U6063 (N_6063,N_5480,N_5212);
and U6064 (N_6064,N_5233,N_5878);
or U6065 (N_6065,N_5561,N_5302);
and U6066 (N_6066,N_5421,N_5710);
nand U6067 (N_6067,N_5120,N_5778);
or U6068 (N_6068,N_5479,N_5523);
or U6069 (N_6069,N_5021,N_5788);
xnor U6070 (N_6070,N_5901,N_5849);
nor U6071 (N_6071,N_5434,N_5880);
nand U6072 (N_6072,N_5551,N_5451);
nor U6073 (N_6073,N_5844,N_5145);
nand U6074 (N_6074,N_5614,N_5224);
nor U6075 (N_6075,N_5566,N_5595);
and U6076 (N_6076,N_5305,N_5049);
and U6077 (N_6077,N_5274,N_5218);
or U6078 (N_6078,N_5385,N_5386);
xor U6079 (N_6079,N_5847,N_5430);
nor U6080 (N_6080,N_5015,N_5404);
nand U6081 (N_6081,N_5728,N_5545);
nand U6082 (N_6082,N_5137,N_5431);
or U6083 (N_6083,N_5851,N_5375);
nor U6084 (N_6084,N_5292,N_5967);
and U6085 (N_6085,N_5365,N_5963);
xnor U6086 (N_6086,N_5519,N_5277);
or U6087 (N_6087,N_5280,N_5588);
nor U6088 (N_6088,N_5085,N_5529);
or U6089 (N_6089,N_5636,N_5581);
or U6090 (N_6090,N_5546,N_5727);
or U6091 (N_6091,N_5158,N_5644);
xor U6092 (N_6092,N_5604,N_5355);
xor U6093 (N_6093,N_5662,N_5990);
nand U6094 (N_6094,N_5019,N_5063);
and U6095 (N_6095,N_5732,N_5999);
or U6096 (N_6096,N_5100,N_5939);
or U6097 (N_6097,N_5463,N_5641);
nor U6098 (N_6098,N_5653,N_5656);
nor U6099 (N_6099,N_5368,N_5957);
nor U6100 (N_6100,N_5440,N_5243);
xor U6101 (N_6101,N_5907,N_5226);
xnor U6102 (N_6102,N_5598,N_5407);
nand U6103 (N_6103,N_5920,N_5262);
nor U6104 (N_6104,N_5023,N_5220);
xnor U6105 (N_6105,N_5180,N_5383);
nand U6106 (N_6106,N_5971,N_5184);
or U6107 (N_6107,N_5922,N_5209);
or U6108 (N_6108,N_5719,N_5181);
nand U6109 (N_6109,N_5472,N_5522);
xor U6110 (N_6110,N_5286,N_5584);
and U6111 (N_6111,N_5390,N_5748);
or U6112 (N_6112,N_5637,N_5805);
or U6113 (N_6113,N_5294,N_5378);
and U6114 (N_6114,N_5039,N_5981);
nor U6115 (N_6115,N_5362,N_5816);
xor U6116 (N_6116,N_5715,N_5084);
and U6117 (N_6117,N_5921,N_5620);
or U6118 (N_6118,N_5706,N_5051);
xor U6119 (N_6119,N_5944,N_5035);
or U6120 (N_6120,N_5001,N_5514);
or U6121 (N_6121,N_5608,N_5578);
nand U6122 (N_6122,N_5449,N_5348);
nand U6123 (N_6123,N_5606,N_5552);
xor U6124 (N_6124,N_5325,N_5961);
nand U6125 (N_6125,N_5539,N_5767);
nor U6126 (N_6126,N_5965,N_5738);
nor U6127 (N_6127,N_5582,N_5908);
or U6128 (N_6128,N_5167,N_5903);
nor U6129 (N_6129,N_5548,N_5031);
nand U6130 (N_6130,N_5490,N_5647);
and U6131 (N_6131,N_5609,N_5760);
or U6132 (N_6132,N_5183,N_5866);
or U6133 (N_6133,N_5766,N_5192);
nand U6134 (N_6134,N_5893,N_5322);
nand U6135 (N_6135,N_5364,N_5263);
xnor U6136 (N_6136,N_5371,N_5401);
or U6137 (N_6137,N_5697,N_5462);
or U6138 (N_6138,N_5897,N_5366);
xnor U6139 (N_6139,N_5078,N_5555);
and U6140 (N_6140,N_5557,N_5815);
and U6141 (N_6141,N_5011,N_5150);
or U6142 (N_6142,N_5834,N_5478);
xor U6143 (N_6143,N_5515,N_5311);
or U6144 (N_6144,N_5792,N_5255);
nand U6145 (N_6145,N_5381,N_5685);
and U6146 (N_6146,N_5070,N_5205);
xor U6147 (N_6147,N_5742,N_5396);
xor U6148 (N_6148,N_5206,N_5842);
and U6149 (N_6149,N_5442,N_5112);
or U6150 (N_6150,N_5170,N_5510);
nand U6151 (N_6151,N_5855,N_5146);
nor U6152 (N_6152,N_5682,N_5291);
nand U6153 (N_6153,N_5982,N_5193);
and U6154 (N_6154,N_5997,N_5195);
or U6155 (N_6155,N_5352,N_5029);
and U6156 (N_6156,N_5335,N_5411);
xnor U6157 (N_6157,N_5786,N_5391);
and U6158 (N_6158,N_5504,N_5435);
nor U6159 (N_6159,N_5819,N_5336);
nand U6160 (N_6160,N_5367,N_5153);
xnor U6161 (N_6161,N_5749,N_5283);
nor U6162 (N_6162,N_5909,N_5361);
or U6163 (N_6163,N_5596,N_5338);
and U6164 (N_6164,N_5591,N_5902);
and U6165 (N_6165,N_5400,N_5703);
or U6166 (N_6166,N_5033,N_5507);
nand U6167 (N_6167,N_5345,N_5432);
nand U6168 (N_6168,N_5973,N_5906);
and U6169 (N_6169,N_5932,N_5107);
nor U6170 (N_6170,N_5429,N_5762);
xnor U6171 (N_6171,N_5144,N_5221);
or U6172 (N_6172,N_5298,N_5201);
or U6173 (N_6173,N_5873,N_5458);
xnor U6174 (N_6174,N_5398,N_5534);
or U6175 (N_6175,N_5952,N_5688);
xor U6176 (N_6176,N_5453,N_5299);
xor U6177 (N_6177,N_5076,N_5590);
xnor U6178 (N_6178,N_5896,N_5468);
nor U6179 (N_6179,N_5172,N_5258);
nand U6180 (N_6180,N_5704,N_5950);
nand U6181 (N_6181,N_5253,N_5940);
xnor U6182 (N_6182,N_5773,N_5115);
and U6183 (N_6183,N_5633,N_5038);
and U6184 (N_6184,N_5502,N_5718);
xnor U6185 (N_6185,N_5946,N_5082);
xnor U6186 (N_6186,N_5511,N_5282);
xor U6187 (N_6187,N_5452,N_5969);
xnor U6188 (N_6188,N_5776,N_5730);
or U6189 (N_6189,N_5392,N_5116);
or U6190 (N_6190,N_5910,N_5796);
nor U6191 (N_6191,N_5712,N_5295);
nand U6192 (N_6192,N_5945,N_5168);
and U6193 (N_6193,N_5729,N_5240);
xor U6194 (N_6194,N_5060,N_5974);
nor U6195 (N_6195,N_5954,N_5203);
and U6196 (N_6196,N_5527,N_5814);
nand U6197 (N_6197,N_5985,N_5147);
xnor U6198 (N_6198,N_5267,N_5313);
and U6199 (N_6199,N_5794,N_5420);
and U6200 (N_6200,N_5071,N_5132);
or U6201 (N_6201,N_5895,N_5042);
and U6202 (N_6202,N_5333,N_5369);
nor U6203 (N_6203,N_5210,N_5624);
and U6204 (N_6204,N_5312,N_5017);
nand U6205 (N_6205,N_5572,N_5676);
nand U6206 (N_6206,N_5217,N_5883);
xor U6207 (N_6207,N_5326,N_5416);
and U6208 (N_6208,N_5651,N_5913);
or U6209 (N_6209,N_5664,N_5062);
xnor U6210 (N_6210,N_5733,N_5185);
nor U6211 (N_6211,N_5395,N_5306);
nor U6212 (N_6212,N_5860,N_5900);
xor U6213 (N_6213,N_5993,N_5852);
and U6214 (N_6214,N_5186,N_5592);
nor U6215 (N_6215,N_5722,N_5931);
or U6216 (N_6216,N_5117,N_5204);
xor U6217 (N_6217,N_5571,N_5002);
and U6218 (N_6218,N_5495,N_5155);
xor U6219 (N_6219,N_5074,N_5488);
nand U6220 (N_6220,N_5857,N_5465);
nor U6221 (N_6221,N_5711,N_5093);
or U6222 (N_6222,N_5443,N_5297);
or U6223 (N_6223,N_5811,N_5657);
xnor U6224 (N_6224,N_5915,N_5055);
or U6225 (N_6225,N_5744,N_5215);
and U6226 (N_6226,N_5419,N_5768);
or U6227 (N_6227,N_5309,N_5314);
and U6228 (N_6228,N_5081,N_5164);
and U6229 (N_6229,N_5177,N_5838);
xor U6230 (N_6230,N_5133,N_5569);
nor U6231 (N_6231,N_5926,N_5445);
and U6232 (N_6232,N_5822,N_5271);
or U6233 (N_6233,N_5652,N_5618);
or U6234 (N_6234,N_5040,N_5579);
nor U6235 (N_6235,N_5166,N_5157);
xnor U6236 (N_6236,N_5027,N_5791);
or U6237 (N_6237,N_5470,N_5245);
xnor U6238 (N_6238,N_5885,N_5043);
nand U6239 (N_6239,N_5717,N_5764);
nor U6240 (N_6240,N_5576,N_5675);
xnor U6241 (N_6241,N_5438,N_5547);
or U6242 (N_6242,N_5272,N_5223);
or U6243 (N_6243,N_5409,N_5134);
or U6244 (N_6244,N_5308,N_5935);
nor U6245 (N_6245,N_5631,N_5667);
xnor U6246 (N_6246,N_5949,N_5376);
xnor U6247 (N_6247,N_5817,N_5991);
nand U6248 (N_6248,N_5526,N_5136);
nor U6249 (N_6249,N_5238,N_5197);
nor U6250 (N_6250,N_5268,N_5171);
nor U6251 (N_6251,N_5394,N_5508);
nor U6252 (N_6252,N_5387,N_5782);
nand U6253 (N_6253,N_5877,N_5363);
xor U6254 (N_6254,N_5293,N_5629);
and U6255 (N_6255,N_5050,N_5191);
or U6256 (N_6256,N_5784,N_5347);
and U6257 (N_6257,N_5269,N_5106);
nand U6258 (N_6258,N_5700,N_5779);
and U6259 (N_6259,N_5261,N_5536);
nand U6260 (N_6260,N_5899,N_5343);
nand U6261 (N_6261,N_5216,N_5611);
xnor U6262 (N_6262,N_5114,N_5473);
nand U6263 (N_6263,N_5554,N_5639);
nor U6264 (N_6264,N_5677,N_5109);
nand U6265 (N_6265,N_5660,N_5845);
and U6266 (N_6266,N_5131,N_5393);
or U6267 (N_6267,N_5389,N_5270);
nand U6268 (N_6268,N_5320,N_5005);
or U6269 (N_6269,N_5339,N_5781);
nand U6270 (N_6270,N_5861,N_5266);
and U6271 (N_6271,N_5679,N_5457);
xor U6272 (N_6272,N_5708,N_5160);
and U6273 (N_6273,N_5709,N_5083);
xnor U6274 (N_6274,N_5057,N_5780);
xor U6275 (N_6275,N_5998,N_5564);
nor U6276 (N_6276,N_5489,N_5149);
or U6277 (N_6277,N_5518,N_5524);
nand U6278 (N_6278,N_5917,N_5332);
xnor U6279 (N_6279,N_5324,N_5765);
or U6280 (N_6280,N_5249,N_5265);
and U6281 (N_6281,N_5317,N_5832);
or U6282 (N_6282,N_5342,N_5787);
and U6283 (N_6283,N_5691,N_5408);
or U6284 (N_6284,N_5976,N_5761);
nand U6285 (N_6285,N_5925,N_5737);
or U6286 (N_6286,N_5918,N_5370);
or U6287 (N_6287,N_5531,N_5276);
or U6288 (N_6288,N_5505,N_5092);
xnor U6289 (N_6289,N_5777,N_5436);
or U6290 (N_6290,N_5121,N_5640);
and U6291 (N_6291,N_5517,N_5125);
nor U6292 (N_6292,N_5123,N_5256);
nor U6293 (N_6293,N_5549,N_5696);
xor U6294 (N_6294,N_5059,N_5846);
or U6295 (N_6295,N_5028,N_5329);
or U6296 (N_6296,N_5065,N_5219);
xnor U6297 (N_6297,N_5410,N_5154);
and U6298 (N_6298,N_5327,N_5627);
nand U6299 (N_6299,N_5942,N_5980);
or U6300 (N_6300,N_5542,N_5067);
nand U6301 (N_6301,N_5541,N_5099);
nand U6302 (N_6302,N_5377,N_5884);
nand U6303 (N_6303,N_5953,N_5222);
nor U6304 (N_6304,N_5736,N_5924);
nor U6305 (N_6305,N_5111,N_5743);
nor U6306 (N_6306,N_5208,N_5009);
xor U6307 (N_6307,N_5829,N_5941);
nand U6308 (N_6308,N_5474,N_5615);
nand U6309 (N_6309,N_5574,N_5937);
xnor U6310 (N_6310,N_5354,N_5890);
nand U6311 (N_6311,N_5623,N_5374);
xor U6312 (N_6312,N_5705,N_5402);
and U6313 (N_6313,N_5178,N_5127);
and U6314 (N_6314,N_5372,N_5673);
and U6315 (N_6315,N_5251,N_5616);
and U6316 (N_6316,N_5678,N_5353);
nor U6317 (N_6317,N_5968,N_5373);
xnor U6318 (N_6318,N_5577,N_5466);
nand U6319 (N_6319,N_5807,N_5642);
nor U6320 (N_6320,N_5983,N_5868);
and U6321 (N_6321,N_5064,N_5097);
or U6322 (N_6322,N_5862,N_5036);
or U6323 (N_6323,N_5840,N_5612);
nor U6324 (N_6324,N_5101,N_5936);
and U6325 (N_6325,N_5234,N_5498);
and U6326 (N_6326,N_5129,N_5972);
xnor U6327 (N_6327,N_5955,N_5521);
nor U6328 (N_6328,N_5499,N_5228);
and U6329 (N_6329,N_5625,N_5301);
nand U6330 (N_6330,N_5412,N_5058);
nand U6331 (N_6331,N_5140,N_5079);
and U6332 (N_6332,N_5091,N_5724);
nand U6333 (N_6333,N_5315,N_5638);
or U6334 (N_6334,N_5648,N_5200);
and U6335 (N_6335,N_5772,N_5573);
nand U6336 (N_6336,N_5321,N_5006);
and U6337 (N_6337,N_5996,N_5535);
and U6338 (N_6338,N_5956,N_5199);
and U6339 (N_6339,N_5622,N_5513);
or U6340 (N_6340,N_5553,N_5471);
nand U6341 (N_6341,N_5538,N_5882);
or U6342 (N_6342,N_5500,N_5041);
or U6343 (N_6343,N_5634,N_5966);
and U6344 (N_6344,N_5929,N_5303);
xor U6345 (N_6345,N_5163,N_5951);
or U6346 (N_6346,N_5413,N_5273);
xnor U6347 (N_6347,N_5987,N_5143);
or U6348 (N_6348,N_5230,N_5239);
nor U6349 (N_6349,N_5241,N_5693);
nand U6350 (N_6350,N_5859,N_5820);
or U6351 (N_6351,N_5689,N_5018);
xnor U6352 (N_6352,N_5543,N_5054);
or U6353 (N_6353,N_5349,N_5872);
nand U6354 (N_6354,N_5189,N_5148);
or U6355 (N_6355,N_5380,N_5278);
nor U6356 (N_6356,N_5528,N_5580);
xnor U6357 (N_6357,N_5447,N_5714);
or U6358 (N_6358,N_5341,N_5894);
xnor U6359 (N_6359,N_5053,N_5986);
nor U6360 (N_6360,N_5975,N_5232);
and U6361 (N_6361,N_5141,N_5889);
and U6362 (N_6362,N_5159,N_5310);
and U6363 (N_6363,N_5594,N_5044);
nor U6364 (N_6364,N_5831,N_5483);
and U6365 (N_6365,N_5094,N_5628);
or U6366 (N_6366,N_5537,N_5207);
nor U6367 (N_6367,N_5175,N_5231);
or U6368 (N_6368,N_5544,N_5279);
or U6369 (N_6369,N_5876,N_5450);
nand U6370 (N_6370,N_5692,N_5605);
and U6371 (N_6371,N_5142,N_5236);
nor U6372 (N_6372,N_5964,N_5771);
or U6373 (N_6373,N_5864,N_5979);
or U6374 (N_6374,N_5448,N_5713);
or U6375 (N_6375,N_5669,N_5977);
xor U6376 (N_6376,N_5340,N_5804);
nor U6377 (N_6377,N_5655,N_5891);
and U6378 (N_6378,N_5562,N_5533);
or U6379 (N_6379,N_5790,N_5188);
xor U6380 (N_6380,N_5532,N_5858);
and U6381 (N_6381,N_5075,N_5459);
nand U6382 (N_6382,N_5095,N_5839);
nand U6383 (N_6383,N_5439,N_5444);
and U6384 (N_6384,N_5619,N_5912);
xor U6385 (N_6385,N_5492,N_5202);
xnor U6386 (N_6386,N_5661,N_5032);
and U6387 (N_6387,N_5995,N_5770);
xor U6388 (N_6388,N_5607,N_5414);
nor U6389 (N_6389,N_5096,N_5621);
nor U6390 (N_6390,N_5069,N_5454);
or U6391 (N_6391,N_5403,N_5586);
or U6392 (N_6392,N_5318,N_5938);
nor U6393 (N_6393,N_5600,N_5214);
nand U6394 (N_6394,N_5003,N_5384);
and U6395 (N_6395,N_5122,N_5360);
or U6396 (N_6396,N_5643,N_5476);
xnor U6397 (N_6397,N_5260,N_5356);
nor U6398 (N_6398,N_5988,N_5187);
or U6399 (N_6399,N_5151,N_5836);
nor U6400 (N_6400,N_5016,N_5307);
nor U6401 (N_6401,N_5030,N_5086);
xor U6402 (N_6402,N_5482,N_5570);
or U6403 (N_6403,N_5126,N_5962);
nor U6404 (N_6404,N_5789,N_5854);
or U6405 (N_6405,N_5072,N_5022);
or U6406 (N_6406,N_5731,N_5477);
nand U6407 (N_6407,N_5382,N_5802);
nand U6408 (N_6408,N_5984,N_5684);
xnor U6409 (N_6409,N_5135,N_5726);
nand U6410 (N_6410,N_5934,N_5746);
xor U6411 (N_6411,N_5585,N_5020);
nand U6412 (N_6412,N_5415,N_5014);
xnor U6413 (N_6413,N_5601,N_5501);
nor U6414 (N_6414,N_5264,N_5589);
or U6415 (N_6415,N_5874,N_5698);
nand U6416 (N_6416,N_5281,N_5304);
nand U6417 (N_6417,N_5785,N_5793);
nor U6418 (N_6418,N_5833,N_5102);
or U6419 (N_6419,N_5124,N_5491);
nand U6420 (N_6420,N_5837,N_5550);
and U6421 (N_6421,N_5176,N_5007);
nand U6422 (N_6422,N_5856,N_5716);
xor U6423 (N_6423,N_5486,N_5699);
nor U6424 (N_6424,N_5351,N_5046);
and U6425 (N_6425,N_5928,N_5073);
nor U6426 (N_6426,N_5610,N_5467);
nor U6427 (N_6427,N_5593,N_5870);
or U6428 (N_6428,N_5098,N_5497);
xnor U6429 (N_6429,N_5821,N_5300);
nand U6430 (N_6430,N_5288,N_5090);
nand U6431 (N_6431,N_5025,N_5674);
xor U6432 (N_6432,N_5914,N_5671);
nand U6433 (N_6433,N_5460,N_5139);
nand U6434 (N_6434,N_5128,N_5428);
nor U6435 (N_6435,N_5418,N_5048);
and U6436 (N_6436,N_5960,N_5603);
and U6437 (N_6437,N_5484,N_5289);
nand U6438 (N_6438,N_5344,N_5379);
nor U6439 (N_6439,N_5179,N_5559);
xor U6440 (N_6440,N_5417,N_5723);
nand U6441 (N_6441,N_5774,N_5330);
nand U6442 (N_6442,N_5801,N_5182);
and U6443 (N_6443,N_5237,N_5863);
nand U6444 (N_6444,N_5923,N_5316);
nor U6445 (N_6445,N_5754,N_5066);
and U6446 (N_6446,N_5797,N_5087);
and U6447 (N_6447,N_5227,N_5174);
xor U6448 (N_6448,N_5568,N_5235);
nand U6449 (N_6449,N_5725,N_5575);
nor U6450 (N_6450,N_5806,N_5613);
nor U6451 (N_6451,N_5818,N_5978);
and U6452 (N_6452,N_5485,N_5841);
nand U6453 (N_6453,N_5441,N_5287);
and U6454 (N_6454,N_5808,N_5357);
nand U6455 (N_6455,N_5702,N_5707);
xnor U6456 (N_6456,N_5118,N_5830);
and U6457 (N_6457,N_5668,N_5756);
or U6458 (N_6458,N_5211,N_5681);
and U6459 (N_6459,N_5089,N_5037);
nand U6460 (N_6460,N_5397,N_5540);
nor U6461 (N_6461,N_5077,N_5024);
nor U6462 (N_6462,N_5252,N_5509);
xor U6463 (N_6463,N_5654,N_5887);
nor U6464 (N_6464,N_5740,N_5823);
xor U6465 (N_6465,N_5290,N_5296);
and U6466 (N_6466,N_5388,N_5423);
nand U6467 (N_6467,N_5867,N_5080);
nor U6468 (N_6468,N_5658,N_5672);
or U6469 (N_6469,N_5152,N_5244);
xor U6470 (N_6470,N_5904,N_5959);
nand U6471 (N_6471,N_5026,N_5229);
xnor U6472 (N_6472,N_5587,N_5047);
nor U6473 (N_6473,N_5464,N_5881);
xnor U6474 (N_6474,N_5947,N_5739);
or U6475 (N_6475,N_5323,N_5119);
or U6476 (N_6476,N_5813,N_5512);
and U6477 (N_6477,N_5558,N_5173);
xnor U6478 (N_6478,N_5783,N_5835);
nand U6479 (N_6479,N_5246,N_5284);
nand U6480 (N_6480,N_5169,N_5769);
and U6481 (N_6481,N_5008,N_5424);
nand U6482 (N_6482,N_5686,N_5487);
nand U6483 (N_6483,N_5426,N_5285);
and U6484 (N_6484,N_5826,N_5583);
and U6485 (N_6485,N_5110,N_5970);
xnor U6486 (N_6486,N_5751,N_5663);
nand U6487 (N_6487,N_5695,N_5617);
or U6488 (N_6488,N_5879,N_5825);
xor U6489 (N_6489,N_5943,N_5461);
nor U6490 (N_6490,N_5506,N_5503);
nand U6491 (N_6491,N_5520,N_5650);
xnor U6492 (N_6492,N_5359,N_5337);
xor U6493 (N_6493,N_5334,N_5433);
and U6494 (N_6494,N_5446,N_5755);
nand U6495 (N_6495,N_5425,N_5475);
and U6496 (N_6496,N_5916,N_5659);
nand U6497 (N_6497,N_5810,N_5275);
or U6498 (N_6498,N_5747,N_5456);
nor U6499 (N_6499,N_5646,N_5525);
xor U6500 (N_6500,N_5579,N_5614);
or U6501 (N_6501,N_5177,N_5713);
nor U6502 (N_6502,N_5053,N_5788);
or U6503 (N_6503,N_5864,N_5762);
or U6504 (N_6504,N_5613,N_5970);
xor U6505 (N_6505,N_5787,N_5784);
xor U6506 (N_6506,N_5644,N_5832);
and U6507 (N_6507,N_5413,N_5525);
xnor U6508 (N_6508,N_5864,N_5552);
or U6509 (N_6509,N_5227,N_5676);
nor U6510 (N_6510,N_5314,N_5210);
and U6511 (N_6511,N_5176,N_5759);
nor U6512 (N_6512,N_5918,N_5906);
or U6513 (N_6513,N_5013,N_5819);
nand U6514 (N_6514,N_5681,N_5989);
and U6515 (N_6515,N_5540,N_5314);
nand U6516 (N_6516,N_5864,N_5983);
and U6517 (N_6517,N_5343,N_5691);
xnor U6518 (N_6518,N_5815,N_5532);
or U6519 (N_6519,N_5131,N_5315);
nor U6520 (N_6520,N_5428,N_5895);
and U6521 (N_6521,N_5046,N_5051);
nor U6522 (N_6522,N_5083,N_5572);
nand U6523 (N_6523,N_5424,N_5373);
nor U6524 (N_6524,N_5254,N_5672);
xor U6525 (N_6525,N_5407,N_5912);
and U6526 (N_6526,N_5770,N_5017);
nand U6527 (N_6527,N_5783,N_5446);
nor U6528 (N_6528,N_5454,N_5824);
and U6529 (N_6529,N_5425,N_5800);
xor U6530 (N_6530,N_5215,N_5053);
or U6531 (N_6531,N_5227,N_5777);
and U6532 (N_6532,N_5404,N_5684);
nor U6533 (N_6533,N_5941,N_5913);
xor U6534 (N_6534,N_5854,N_5265);
xnor U6535 (N_6535,N_5036,N_5321);
or U6536 (N_6536,N_5424,N_5681);
nor U6537 (N_6537,N_5049,N_5927);
xnor U6538 (N_6538,N_5880,N_5426);
nor U6539 (N_6539,N_5936,N_5319);
xnor U6540 (N_6540,N_5919,N_5463);
nand U6541 (N_6541,N_5856,N_5616);
and U6542 (N_6542,N_5436,N_5278);
xor U6543 (N_6543,N_5679,N_5815);
xnor U6544 (N_6544,N_5866,N_5619);
nand U6545 (N_6545,N_5993,N_5262);
xor U6546 (N_6546,N_5580,N_5400);
or U6547 (N_6547,N_5287,N_5561);
nand U6548 (N_6548,N_5380,N_5816);
nand U6549 (N_6549,N_5834,N_5549);
xor U6550 (N_6550,N_5188,N_5173);
nor U6551 (N_6551,N_5826,N_5942);
or U6552 (N_6552,N_5684,N_5927);
or U6553 (N_6553,N_5279,N_5497);
or U6554 (N_6554,N_5380,N_5226);
xnor U6555 (N_6555,N_5525,N_5216);
and U6556 (N_6556,N_5746,N_5853);
or U6557 (N_6557,N_5390,N_5244);
or U6558 (N_6558,N_5978,N_5143);
xnor U6559 (N_6559,N_5341,N_5807);
or U6560 (N_6560,N_5355,N_5108);
xor U6561 (N_6561,N_5521,N_5490);
xor U6562 (N_6562,N_5300,N_5301);
nor U6563 (N_6563,N_5327,N_5828);
or U6564 (N_6564,N_5570,N_5940);
nor U6565 (N_6565,N_5456,N_5359);
nand U6566 (N_6566,N_5548,N_5995);
or U6567 (N_6567,N_5213,N_5023);
nand U6568 (N_6568,N_5863,N_5334);
nand U6569 (N_6569,N_5703,N_5198);
and U6570 (N_6570,N_5138,N_5340);
nand U6571 (N_6571,N_5867,N_5147);
nand U6572 (N_6572,N_5264,N_5218);
or U6573 (N_6573,N_5265,N_5828);
nand U6574 (N_6574,N_5361,N_5884);
xnor U6575 (N_6575,N_5240,N_5260);
xor U6576 (N_6576,N_5570,N_5034);
and U6577 (N_6577,N_5093,N_5500);
nand U6578 (N_6578,N_5155,N_5152);
nand U6579 (N_6579,N_5620,N_5723);
nor U6580 (N_6580,N_5932,N_5594);
nand U6581 (N_6581,N_5994,N_5560);
and U6582 (N_6582,N_5650,N_5980);
nand U6583 (N_6583,N_5160,N_5287);
nand U6584 (N_6584,N_5626,N_5408);
nand U6585 (N_6585,N_5907,N_5430);
nor U6586 (N_6586,N_5475,N_5915);
nor U6587 (N_6587,N_5124,N_5925);
or U6588 (N_6588,N_5093,N_5805);
nor U6589 (N_6589,N_5950,N_5923);
nor U6590 (N_6590,N_5739,N_5664);
xor U6591 (N_6591,N_5154,N_5833);
xor U6592 (N_6592,N_5764,N_5699);
or U6593 (N_6593,N_5907,N_5574);
xor U6594 (N_6594,N_5818,N_5471);
nor U6595 (N_6595,N_5385,N_5482);
xnor U6596 (N_6596,N_5134,N_5732);
and U6597 (N_6597,N_5034,N_5335);
or U6598 (N_6598,N_5293,N_5482);
or U6599 (N_6599,N_5197,N_5970);
or U6600 (N_6600,N_5508,N_5595);
and U6601 (N_6601,N_5411,N_5906);
nor U6602 (N_6602,N_5928,N_5814);
or U6603 (N_6603,N_5949,N_5636);
or U6604 (N_6604,N_5132,N_5415);
or U6605 (N_6605,N_5467,N_5447);
nor U6606 (N_6606,N_5326,N_5322);
or U6607 (N_6607,N_5048,N_5470);
and U6608 (N_6608,N_5834,N_5953);
or U6609 (N_6609,N_5873,N_5172);
nor U6610 (N_6610,N_5523,N_5387);
and U6611 (N_6611,N_5664,N_5283);
xnor U6612 (N_6612,N_5443,N_5365);
or U6613 (N_6613,N_5621,N_5748);
and U6614 (N_6614,N_5352,N_5743);
xnor U6615 (N_6615,N_5891,N_5448);
and U6616 (N_6616,N_5678,N_5361);
or U6617 (N_6617,N_5906,N_5279);
and U6618 (N_6618,N_5007,N_5996);
nor U6619 (N_6619,N_5499,N_5478);
or U6620 (N_6620,N_5817,N_5986);
xor U6621 (N_6621,N_5838,N_5870);
xnor U6622 (N_6622,N_5810,N_5623);
or U6623 (N_6623,N_5931,N_5685);
and U6624 (N_6624,N_5838,N_5207);
xnor U6625 (N_6625,N_5954,N_5415);
and U6626 (N_6626,N_5353,N_5962);
nor U6627 (N_6627,N_5498,N_5813);
and U6628 (N_6628,N_5991,N_5005);
xor U6629 (N_6629,N_5818,N_5251);
nand U6630 (N_6630,N_5715,N_5100);
xor U6631 (N_6631,N_5073,N_5137);
nand U6632 (N_6632,N_5063,N_5615);
or U6633 (N_6633,N_5852,N_5350);
xor U6634 (N_6634,N_5256,N_5501);
nor U6635 (N_6635,N_5303,N_5484);
nor U6636 (N_6636,N_5576,N_5252);
or U6637 (N_6637,N_5906,N_5761);
xnor U6638 (N_6638,N_5063,N_5530);
xnor U6639 (N_6639,N_5572,N_5386);
and U6640 (N_6640,N_5286,N_5825);
xor U6641 (N_6641,N_5427,N_5494);
and U6642 (N_6642,N_5708,N_5448);
nor U6643 (N_6643,N_5162,N_5778);
and U6644 (N_6644,N_5836,N_5118);
and U6645 (N_6645,N_5425,N_5804);
xor U6646 (N_6646,N_5332,N_5851);
and U6647 (N_6647,N_5402,N_5079);
nor U6648 (N_6648,N_5262,N_5558);
nand U6649 (N_6649,N_5393,N_5473);
nand U6650 (N_6650,N_5384,N_5733);
nand U6651 (N_6651,N_5300,N_5934);
xor U6652 (N_6652,N_5143,N_5465);
or U6653 (N_6653,N_5690,N_5788);
and U6654 (N_6654,N_5553,N_5391);
xor U6655 (N_6655,N_5443,N_5849);
nand U6656 (N_6656,N_5738,N_5983);
xor U6657 (N_6657,N_5122,N_5870);
nand U6658 (N_6658,N_5833,N_5151);
nand U6659 (N_6659,N_5746,N_5369);
or U6660 (N_6660,N_5992,N_5723);
or U6661 (N_6661,N_5427,N_5919);
or U6662 (N_6662,N_5712,N_5358);
nand U6663 (N_6663,N_5568,N_5698);
nand U6664 (N_6664,N_5837,N_5548);
or U6665 (N_6665,N_5115,N_5667);
or U6666 (N_6666,N_5833,N_5426);
nor U6667 (N_6667,N_5092,N_5617);
and U6668 (N_6668,N_5827,N_5491);
and U6669 (N_6669,N_5275,N_5477);
nand U6670 (N_6670,N_5439,N_5960);
nor U6671 (N_6671,N_5054,N_5725);
xnor U6672 (N_6672,N_5704,N_5859);
nor U6673 (N_6673,N_5019,N_5582);
nand U6674 (N_6674,N_5121,N_5112);
xor U6675 (N_6675,N_5418,N_5262);
xnor U6676 (N_6676,N_5385,N_5928);
and U6677 (N_6677,N_5039,N_5182);
xor U6678 (N_6678,N_5180,N_5503);
and U6679 (N_6679,N_5003,N_5529);
nor U6680 (N_6680,N_5852,N_5425);
nor U6681 (N_6681,N_5068,N_5142);
nand U6682 (N_6682,N_5039,N_5142);
nand U6683 (N_6683,N_5739,N_5991);
nand U6684 (N_6684,N_5395,N_5969);
xnor U6685 (N_6685,N_5244,N_5588);
xnor U6686 (N_6686,N_5187,N_5851);
or U6687 (N_6687,N_5402,N_5401);
xnor U6688 (N_6688,N_5133,N_5298);
nor U6689 (N_6689,N_5702,N_5146);
nand U6690 (N_6690,N_5141,N_5706);
and U6691 (N_6691,N_5201,N_5490);
and U6692 (N_6692,N_5371,N_5058);
nor U6693 (N_6693,N_5776,N_5417);
nor U6694 (N_6694,N_5330,N_5520);
and U6695 (N_6695,N_5230,N_5584);
nor U6696 (N_6696,N_5766,N_5792);
nand U6697 (N_6697,N_5108,N_5594);
and U6698 (N_6698,N_5112,N_5988);
nand U6699 (N_6699,N_5649,N_5931);
or U6700 (N_6700,N_5925,N_5745);
nor U6701 (N_6701,N_5546,N_5908);
or U6702 (N_6702,N_5991,N_5408);
nor U6703 (N_6703,N_5542,N_5142);
and U6704 (N_6704,N_5845,N_5521);
nor U6705 (N_6705,N_5444,N_5991);
xnor U6706 (N_6706,N_5773,N_5841);
and U6707 (N_6707,N_5582,N_5808);
nor U6708 (N_6708,N_5215,N_5029);
and U6709 (N_6709,N_5803,N_5202);
or U6710 (N_6710,N_5442,N_5361);
or U6711 (N_6711,N_5384,N_5184);
or U6712 (N_6712,N_5643,N_5310);
nand U6713 (N_6713,N_5851,N_5492);
or U6714 (N_6714,N_5002,N_5526);
nor U6715 (N_6715,N_5305,N_5677);
xnor U6716 (N_6716,N_5957,N_5149);
or U6717 (N_6717,N_5211,N_5725);
nand U6718 (N_6718,N_5011,N_5156);
nand U6719 (N_6719,N_5241,N_5031);
and U6720 (N_6720,N_5961,N_5629);
and U6721 (N_6721,N_5631,N_5033);
xnor U6722 (N_6722,N_5835,N_5349);
xor U6723 (N_6723,N_5623,N_5005);
and U6724 (N_6724,N_5610,N_5640);
nor U6725 (N_6725,N_5981,N_5288);
xor U6726 (N_6726,N_5619,N_5281);
nor U6727 (N_6727,N_5005,N_5581);
or U6728 (N_6728,N_5339,N_5017);
xnor U6729 (N_6729,N_5903,N_5611);
xnor U6730 (N_6730,N_5783,N_5116);
nor U6731 (N_6731,N_5737,N_5405);
or U6732 (N_6732,N_5104,N_5906);
xor U6733 (N_6733,N_5624,N_5443);
and U6734 (N_6734,N_5760,N_5116);
or U6735 (N_6735,N_5334,N_5012);
xnor U6736 (N_6736,N_5363,N_5316);
nor U6737 (N_6737,N_5117,N_5314);
and U6738 (N_6738,N_5436,N_5438);
nor U6739 (N_6739,N_5189,N_5779);
and U6740 (N_6740,N_5479,N_5354);
or U6741 (N_6741,N_5329,N_5376);
nand U6742 (N_6742,N_5682,N_5659);
nor U6743 (N_6743,N_5679,N_5887);
nand U6744 (N_6744,N_5774,N_5278);
or U6745 (N_6745,N_5872,N_5903);
nor U6746 (N_6746,N_5453,N_5069);
or U6747 (N_6747,N_5364,N_5499);
xor U6748 (N_6748,N_5510,N_5687);
nand U6749 (N_6749,N_5632,N_5171);
nor U6750 (N_6750,N_5067,N_5395);
nor U6751 (N_6751,N_5337,N_5907);
xnor U6752 (N_6752,N_5934,N_5588);
or U6753 (N_6753,N_5737,N_5335);
nor U6754 (N_6754,N_5796,N_5899);
nand U6755 (N_6755,N_5439,N_5064);
and U6756 (N_6756,N_5347,N_5296);
or U6757 (N_6757,N_5991,N_5538);
nand U6758 (N_6758,N_5724,N_5294);
xnor U6759 (N_6759,N_5172,N_5972);
xor U6760 (N_6760,N_5836,N_5541);
xor U6761 (N_6761,N_5181,N_5977);
nor U6762 (N_6762,N_5929,N_5830);
xor U6763 (N_6763,N_5105,N_5719);
xnor U6764 (N_6764,N_5052,N_5889);
nand U6765 (N_6765,N_5554,N_5370);
nor U6766 (N_6766,N_5942,N_5339);
and U6767 (N_6767,N_5548,N_5619);
and U6768 (N_6768,N_5929,N_5869);
nand U6769 (N_6769,N_5663,N_5639);
and U6770 (N_6770,N_5220,N_5824);
nand U6771 (N_6771,N_5216,N_5933);
xor U6772 (N_6772,N_5347,N_5362);
and U6773 (N_6773,N_5196,N_5221);
or U6774 (N_6774,N_5729,N_5096);
nand U6775 (N_6775,N_5377,N_5129);
xor U6776 (N_6776,N_5716,N_5931);
nor U6777 (N_6777,N_5621,N_5887);
nor U6778 (N_6778,N_5134,N_5388);
nand U6779 (N_6779,N_5824,N_5055);
nand U6780 (N_6780,N_5267,N_5254);
and U6781 (N_6781,N_5963,N_5878);
and U6782 (N_6782,N_5116,N_5986);
xor U6783 (N_6783,N_5930,N_5007);
nand U6784 (N_6784,N_5230,N_5282);
xor U6785 (N_6785,N_5708,N_5319);
nand U6786 (N_6786,N_5379,N_5538);
or U6787 (N_6787,N_5653,N_5476);
nand U6788 (N_6788,N_5842,N_5950);
nand U6789 (N_6789,N_5062,N_5895);
or U6790 (N_6790,N_5616,N_5003);
nor U6791 (N_6791,N_5432,N_5192);
nand U6792 (N_6792,N_5584,N_5635);
or U6793 (N_6793,N_5902,N_5866);
nor U6794 (N_6794,N_5560,N_5397);
nand U6795 (N_6795,N_5772,N_5490);
nand U6796 (N_6796,N_5839,N_5628);
xor U6797 (N_6797,N_5694,N_5815);
nand U6798 (N_6798,N_5204,N_5486);
and U6799 (N_6799,N_5116,N_5972);
and U6800 (N_6800,N_5199,N_5393);
nand U6801 (N_6801,N_5636,N_5059);
and U6802 (N_6802,N_5398,N_5938);
nor U6803 (N_6803,N_5748,N_5753);
xor U6804 (N_6804,N_5099,N_5895);
or U6805 (N_6805,N_5062,N_5686);
xor U6806 (N_6806,N_5820,N_5787);
or U6807 (N_6807,N_5540,N_5672);
nand U6808 (N_6808,N_5542,N_5135);
nand U6809 (N_6809,N_5675,N_5061);
xnor U6810 (N_6810,N_5452,N_5588);
nor U6811 (N_6811,N_5094,N_5411);
or U6812 (N_6812,N_5944,N_5453);
or U6813 (N_6813,N_5864,N_5660);
nand U6814 (N_6814,N_5189,N_5737);
and U6815 (N_6815,N_5908,N_5288);
and U6816 (N_6816,N_5975,N_5516);
nor U6817 (N_6817,N_5616,N_5454);
xor U6818 (N_6818,N_5743,N_5313);
and U6819 (N_6819,N_5511,N_5603);
and U6820 (N_6820,N_5751,N_5306);
or U6821 (N_6821,N_5752,N_5854);
nor U6822 (N_6822,N_5110,N_5266);
nor U6823 (N_6823,N_5033,N_5168);
xor U6824 (N_6824,N_5713,N_5123);
and U6825 (N_6825,N_5098,N_5942);
nor U6826 (N_6826,N_5139,N_5103);
nand U6827 (N_6827,N_5352,N_5603);
xnor U6828 (N_6828,N_5766,N_5235);
nor U6829 (N_6829,N_5647,N_5428);
nor U6830 (N_6830,N_5920,N_5165);
xor U6831 (N_6831,N_5612,N_5153);
or U6832 (N_6832,N_5682,N_5579);
nand U6833 (N_6833,N_5442,N_5487);
nor U6834 (N_6834,N_5178,N_5828);
nand U6835 (N_6835,N_5245,N_5591);
and U6836 (N_6836,N_5761,N_5668);
or U6837 (N_6837,N_5260,N_5898);
nor U6838 (N_6838,N_5770,N_5719);
or U6839 (N_6839,N_5627,N_5663);
nand U6840 (N_6840,N_5602,N_5323);
or U6841 (N_6841,N_5063,N_5669);
and U6842 (N_6842,N_5237,N_5412);
nand U6843 (N_6843,N_5341,N_5808);
or U6844 (N_6844,N_5451,N_5970);
nand U6845 (N_6845,N_5440,N_5431);
nor U6846 (N_6846,N_5984,N_5183);
or U6847 (N_6847,N_5594,N_5869);
nand U6848 (N_6848,N_5084,N_5585);
xor U6849 (N_6849,N_5493,N_5977);
nor U6850 (N_6850,N_5236,N_5534);
nor U6851 (N_6851,N_5027,N_5409);
nand U6852 (N_6852,N_5949,N_5293);
or U6853 (N_6853,N_5954,N_5116);
or U6854 (N_6854,N_5604,N_5709);
or U6855 (N_6855,N_5943,N_5287);
and U6856 (N_6856,N_5455,N_5731);
and U6857 (N_6857,N_5032,N_5414);
nor U6858 (N_6858,N_5587,N_5430);
or U6859 (N_6859,N_5872,N_5266);
nand U6860 (N_6860,N_5134,N_5286);
or U6861 (N_6861,N_5098,N_5422);
xnor U6862 (N_6862,N_5851,N_5432);
or U6863 (N_6863,N_5309,N_5329);
nand U6864 (N_6864,N_5363,N_5624);
or U6865 (N_6865,N_5710,N_5822);
and U6866 (N_6866,N_5836,N_5339);
and U6867 (N_6867,N_5838,N_5070);
nand U6868 (N_6868,N_5322,N_5320);
and U6869 (N_6869,N_5830,N_5379);
nand U6870 (N_6870,N_5084,N_5338);
nand U6871 (N_6871,N_5547,N_5105);
xnor U6872 (N_6872,N_5324,N_5064);
nor U6873 (N_6873,N_5009,N_5924);
nand U6874 (N_6874,N_5605,N_5606);
xor U6875 (N_6875,N_5912,N_5365);
and U6876 (N_6876,N_5936,N_5471);
nor U6877 (N_6877,N_5820,N_5487);
nand U6878 (N_6878,N_5888,N_5236);
or U6879 (N_6879,N_5643,N_5580);
nand U6880 (N_6880,N_5888,N_5437);
nand U6881 (N_6881,N_5667,N_5164);
nand U6882 (N_6882,N_5670,N_5249);
nand U6883 (N_6883,N_5774,N_5828);
nor U6884 (N_6884,N_5082,N_5370);
nor U6885 (N_6885,N_5194,N_5813);
nor U6886 (N_6886,N_5469,N_5423);
nand U6887 (N_6887,N_5084,N_5371);
and U6888 (N_6888,N_5456,N_5539);
xor U6889 (N_6889,N_5950,N_5733);
or U6890 (N_6890,N_5600,N_5735);
or U6891 (N_6891,N_5824,N_5699);
nor U6892 (N_6892,N_5660,N_5807);
and U6893 (N_6893,N_5923,N_5560);
or U6894 (N_6894,N_5580,N_5890);
nor U6895 (N_6895,N_5755,N_5638);
nor U6896 (N_6896,N_5262,N_5966);
nand U6897 (N_6897,N_5731,N_5584);
nand U6898 (N_6898,N_5608,N_5070);
and U6899 (N_6899,N_5447,N_5726);
nand U6900 (N_6900,N_5874,N_5516);
xnor U6901 (N_6901,N_5362,N_5014);
or U6902 (N_6902,N_5598,N_5784);
nand U6903 (N_6903,N_5678,N_5990);
nor U6904 (N_6904,N_5201,N_5339);
xnor U6905 (N_6905,N_5107,N_5544);
xnor U6906 (N_6906,N_5087,N_5381);
or U6907 (N_6907,N_5622,N_5558);
nand U6908 (N_6908,N_5433,N_5203);
or U6909 (N_6909,N_5051,N_5052);
xor U6910 (N_6910,N_5903,N_5411);
or U6911 (N_6911,N_5274,N_5164);
and U6912 (N_6912,N_5477,N_5249);
xor U6913 (N_6913,N_5929,N_5874);
nor U6914 (N_6914,N_5971,N_5741);
or U6915 (N_6915,N_5319,N_5689);
xor U6916 (N_6916,N_5180,N_5855);
nor U6917 (N_6917,N_5528,N_5390);
and U6918 (N_6918,N_5320,N_5153);
xor U6919 (N_6919,N_5043,N_5247);
nand U6920 (N_6920,N_5720,N_5150);
xor U6921 (N_6921,N_5489,N_5116);
and U6922 (N_6922,N_5438,N_5034);
or U6923 (N_6923,N_5215,N_5884);
or U6924 (N_6924,N_5995,N_5670);
or U6925 (N_6925,N_5684,N_5300);
nand U6926 (N_6926,N_5028,N_5411);
or U6927 (N_6927,N_5564,N_5774);
or U6928 (N_6928,N_5567,N_5201);
nor U6929 (N_6929,N_5909,N_5359);
nor U6930 (N_6930,N_5559,N_5153);
xor U6931 (N_6931,N_5970,N_5554);
nor U6932 (N_6932,N_5823,N_5892);
xor U6933 (N_6933,N_5428,N_5485);
nand U6934 (N_6934,N_5682,N_5007);
xnor U6935 (N_6935,N_5378,N_5638);
or U6936 (N_6936,N_5631,N_5930);
nor U6937 (N_6937,N_5920,N_5249);
xnor U6938 (N_6938,N_5812,N_5655);
nor U6939 (N_6939,N_5460,N_5095);
nor U6940 (N_6940,N_5987,N_5635);
and U6941 (N_6941,N_5562,N_5030);
xor U6942 (N_6942,N_5726,N_5245);
nand U6943 (N_6943,N_5658,N_5278);
or U6944 (N_6944,N_5136,N_5840);
and U6945 (N_6945,N_5144,N_5813);
or U6946 (N_6946,N_5544,N_5141);
nor U6947 (N_6947,N_5894,N_5353);
nand U6948 (N_6948,N_5519,N_5937);
nor U6949 (N_6949,N_5363,N_5990);
xnor U6950 (N_6950,N_5084,N_5915);
xnor U6951 (N_6951,N_5450,N_5464);
nor U6952 (N_6952,N_5206,N_5800);
nor U6953 (N_6953,N_5455,N_5100);
nand U6954 (N_6954,N_5951,N_5333);
xnor U6955 (N_6955,N_5139,N_5637);
or U6956 (N_6956,N_5360,N_5085);
nor U6957 (N_6957,N_5316,N_5019);
xnor U6958 (N_6958,N_5662,N_5230);
or U6959 (N_6959,N_5997,N_5232);
nand U6960 (N_6960,N_5288,N_5029);
and U6961 (N_6961,N_5947,N_5926);
and U6962 (N_6962,N_5767,N_5881);
xnor U6963 (N_6963,N_5901,N_5752);
and U6964 (N_6964,N_5210,N_5588);
and U6965 (N_6965,N_5954,N_5615);
nor U6966 (N_6966,N_5720,N_5665);
xnor U6967 (N_6967,N_5840,N_5213);
and U6968 (N_6968,N_5174,N_5173);
xor U6969 (N_6969,N_5119,N_5240);
or U6970 (N_6970,N_5997,N_5763);
or U6971 (N_6971,N_5911,N_5692);
nand U6972 (N_6972,N_5431,N_5562);
or U6973 (N_6973,N_5716,N_5768);
and U6974 (N_6974,N_5865,N_5125);
or U6975 (N_6975,N_5198,N_5995);
nor U6976 (N_6976,N_5994,N_5990);
nor U6977 (N_6977,N_5013,N_5063);
and U6978 (N_6978,N_5239,N_5969);
nand U6979 (N_6979,N_5231,N_5575);
xor U6980 (N_6980,N_5576,N_5958);
and U6981 (N_6981,N_5290,N_5363);
or U6982 (N_6982,N_5190,N_5869);
or U6983 (N_6983,N_5726,N_5561);
xnor U6984 (N_6984,N_5901,N_5333);
nand U6985 (N_6985,N_5226,N_5323);
nor U6986 (N_6986,N_5591,N_5497);
xor U6987 (N_6987,N_5561,N_5842);
xor U6988 (N_6988,N_5738,N_5815);
nand U6989 (N_6989,N_5743,N_5243);
xor U6990 (N_6990,N_5024,N_5453);
or U6991 (N_6991,N_5483,N_5944);
and U6992 (N_6992,N_5034,N_5386);
xnor U6993 (N_6993,N_5437,N_5719);
nor U6994 (N_6994,N_5536,N_5712);
and U6995 (N_6995,N_5100,N_5816);
and U6996 (N_6996,N_5662,N_5776);
or U6997 (N_6997,N_5517,N_5605);
or U6998 (N_6998,N_5335,N_5104);
nand U6999 (N_6999,N_5908,N_5906);
nor U7000 (N_7000,N_6296,N_6693);
and U7001 (N_7001,N_6670,N_6940);
or U7002 (N_7002,N_6671,N_6688);
or U7003 (N_7003,N_6981,N_6139);
xnor U7004 (N_7004,N_6014,N_6637);
nand U7005 (N_7005,N_6140,N_6512);
nand U7006 (N_7006,N_6681,N_6542);
nand U7007 (N_7007,N_6739,N_6357);
xnor U7008 (N_7008,N_6582,N_6327);
and U7009 (N_7009,N_6137,N_6768);
or U7010 (N_7010,N_6146,N_6600);
and U7011 (N_7011,N_6998,N_6079);
nor U7012 (N_7012,N_6969,N_6439);
xor U7013 (N_7013,N_6385,N_6813);
nand U7014 (N_7014,N_6366,N_6571);
nor U7015 (N_7015,N_6594,N_6817);
and U7016 (N_7016,N_6651,N_6982);
nor U7017 (N_7017,N_6658,N_6728);
or U7018 (N_7018,N_6446,N_6313);
and U7019 (N_7019,N_6212,N_6973);
and U7020 (N_7020,N_6548,N_6599);
nor U7021 (N_7021,N_6369,N_6622);
or U7022 (N_7022,N_6669,N_6545);
or U7023 (N_7023,N_6523,N_6463);
xor U7024 (N_7024,N_6855,N_6227);
or U7025 (N_7025,N_6776,N_6844);
and U7026 (N_7026,N_6726,N_6390);
or U7027 (N_7027,N_6355,N_6980);
nor U7028 (N_7028,N_6265,N_6574);
or U7029 (N_7029,N_6051,N_6967);
nor U7030 (N_7030,N_6904,N_6462);
or U7031 (N_7031,N_6121,N_6602);
or U7032 (N_7032,N_6011,N_6849);
nand U7033 (N_7033,N_6577,N_6065);
and U7034 (N_7034,N_6499,N_6229);
nor U7035 (N_7035,N_6340,N_6775);
nor U7036 (N_7036,N_6573,N_6682);
nand U7037 (N_7037,N_6906,N_6226);
or U7038 (N_7038,N_6230,N_6092);
xor U7039 (N_7039,N_6762,N_6984);
nand U7040 (N_7040,N_6037,N_6897);
nand U7041 (N_7041,N_6114,N_6828);
nor U7042 (N_7042,N_6736,N_6552);
and U7043 (N_7043,N_6514,N_6405);
nand U7044 (N_7044,N_6960,N_6052);
and U7045 (N_7045,N_6246,N_6947);
and U7046 (N_7046,N_6862,N_6206);
xor U7047 (N_7047,N_6713,N_6101);
nor U7048 (N_7048,N_6287,N_6363);
and U7049 (N_7049,N_6319,N_6174);
nor U7050 (N_7050,N_6742,N_6565);
nor U7051 (N_7051,N_6173,N_6288);
and U7052 (N_7052,N_6664,N_6223);
or U7053 (N_7053,N_6667,N_6692);
nand U7054 (N_7054,N_6239,N_6961);
or U7055 (N_7055,N_6335,N_6394);
xnor U7056 (N_7056,N_6191,N_6730);
and U7057 (N_7057,N_6911,N_6816);
nand U7058 (N_7058,N_6080,N_6978);
nor U7059 (N_7059,N_6497,N_6533);
and U7060 (N_7060,N_6604,N_6541);
nor U7061 (N_7061,N_6386,N_6245);
nor U7062 (N_7062,N_6469,N_6814);
xnor U7063 (N_7063,N_6216,N_6401);
or U7064 (N_7064,N_6777,N_6719);
nor U7065 (N_7065,N_6506,N_6889);
or U7066 (N_7066,N_6979,N_6425);
xor U7067 (N_7067,N_6735,N_6916);
or U7068 (N_7068,N_6704,N_6259);
xor U7069 (N_7069,N_6192,N_6220);
nand U7070 (N_7070,N_6486,N_6913);
or U7071 (N_7071,N_6010,N_6822);
nand U7072 (N_7072,N_6878,N_6528);
and U7073 (N_7073,N_6891,N_6679);
nand U7074 (N_7074,N_6718,N_6027);
nand U7075 (N_7075,N_6881,N_6242);
nor U7076 (N_7076,N_6299,N_6927);
xnor U7077 (N_7077,N_6605,N_6185);
or U7078 (N_7078,N_6617,N_6663);
xnor U7079 (N_7079,N_6968,N_6078);
nor U7080 (N_7080,N_6427,N_6801);
or U7081 (N_7081,N_6122,N_6187);
xor U7082 (N_7082,N_6473,N_6767);
nand U7083 (N_7083,N_6616,N_6323);
nor U7084 (N_7084,N_6962,N_6503);
or U7085 (N_7085,N_6148,N_6654);
and U7086 (N_7086,N_6361,N_6731);
xor U7087 (N_7087,N_6983,N_6966);
and U7088 (N_7088,N_6064,N_6636);
and U7089 (N_7089,N_6102,N_6289);
xor U7090 (N_7090,N_6831,N_6930);
nor U7091 (N_7091,N_6184,N_6786);
and U7092 (N_7092,N_6826,N_6224);
or U7093 (N_7093,N_6527,N_6235);
nor U7094 (N_7094,N_6537,N_6627);
and U7095 (N_7095,N_6346,N_6359);
nand U7096 (N_7096,N_6181,N_6870);
nand U7097 (N_7097,N_6766,N_6480);
nand U7098 (N_7098,N_6465,N_6393);
or U7099 (N_7099,N_6408,N_6155);
xnor U7100 (N_7100,N_6632,N_6494);
nand U7101 (N_7101,N_6807,N_6917);
and U7102 (N_7102,N_6186,N_6270);
nand U7103 (N_7103,N_6492,N_6772);
or U7104 (N_7104,N_6232,N_6406);
xnor U7105 (N_7105,N_6213,N_6596);
nor U7106 (N_7106,N_6205,N_6662);
xor U7107 (N_7107,N_6708,N_6721);
xor U7108 (N_7108,N_6672,N_6055);
and U7109 (N_7109,N_6188,N_6524);
xor U7110 (N_7110,N_6628,N_6788);
nor U7111 (N_7111,N_6928,N_6309);
nand U7112 (N_7112,N_6081,N_6536);
and U7113 (N_7113,N_6857,N_6034);
nand U7114 (N_7114,N_6303,N_6901);
nand U7115 (N_7115,N_6260,N_6661);
nand U7116 (N_7116,N_6564,N_6640);
nand U7117 (N_7117,N_6091,N_6566);
and U7118 (N_7118,N_6532,N_6020);
and U7119 (N_7119,N_6105,N_6488);
or U7120 (N_7120,N_6630,N_6858);
nand U7121 (N_7121,N_6032,N_6097);
xnor U7122 (N_7122,N_6515,N_6885);
and U7123 (N_7123,N_6058,N_6539);
xnor U7124 (N_7124,N_6448,N_6107);
nor U7125 (N_7125,N_6601,N_6478);
xor U7126 (N_7126,N_6316,N_6135);
nor U7127 (N_7127,N_6644,N_6291);
or U7128 (N_7128,N_6421,N_6936);
or U7129 (N_7129,N_6625,N_6496);
nor U7130 (N_7130,N_6687,N_6209);
and U7131 (N_7131,N_6322,N_6996);
nand U7132 (N_7132,N_6540,N_6021);
xnor U7133 (N_7133,N_6873,N_6908);
nor U7134 (N_7134,N_6030,N_6505);
nor U7135 (N_7135,N_6903,N_6576);
and U7136 (N_7136,N_6202,N_6723);
nor U7137 (N_7137,N_6290,N_6389);
nand U7138 (N_7138,N_6061,N_6685);
and U7139 (N_7139,N_6986,N_6578);
nand U7140 (N_7140,N_6441,N_6697);
and U7141 (N_7141,N_6128,N_6038);
xnor U7142 (N_7142,N_6162,N_6821);
xor U7143 (N_7143,N_6145,N_6074);
or U7144 (N_7144,N_6431,N_6626);
nor U7145 (N_7145,N_6902,N_6294);
xnor U7146 (N_7146,N_6161,N_6467);
or U7147 (N_7147,N_6362,N_6694);
xnor U7148 (N_7148,N_6069,N_6219);
nand U7149 (N_7149,N_6832,N_6396);
nand U7150 (N_7150,N_6470,N_6588);
nor U7151 (N_7151,N_6563,N_6138);
or U7152 (N_7152,N_6603,N_6942);
and U7153 (N_7153,N_6867,N_6975);
and U7154 (N_7154,N_6676,N_6567);
xor U7155 (N_7155,N_6634,N_6825);
or U7156 (N_7156,N_6189,N_6113);
xor U7157 (N_7157,N_6999,N_6424);
and U7158 (N_7158,N_6190,N_6195);
and U7159 (N_7159,N_6006,N_6874);
or U7160 (N_7160,N_6060,N_6400);
nor U7161 (N_7161,N_6391,N_6823);
xnor U7162 (N_7162,N_6647,N_6877);
xnor U7163 (N_7163,N_6865,N_6453);
and U7164 (N_7164,N_6244,N_6798);
or U7165 (N_7165,N_6144,N_6194);
nor U7166 (N_7166,N_6554,N_6824);
nand U7167 (N_7167,N_6325,N_6447);
and U7168 (N_7168,N_6853,N_6268);
xnor U7169 (N_7169,N_6458,N_6845);
nand U7170 (N_7170,N_6311,N_6909);
xor U7171 (N_7171,N_6922,N_6300);
nor U7172 (N_7172,N_6710,N_6784);
nor U7173 (N_7173,N_6292,N_6587);
xnor U7174 (N_7174,N_6175,N_6379);
nor U7175 (N_7175,N_6275,N_6864);
or U7176 (N_7176,N_6987,N_6787);
and U7177 (N_7177,N_6521,N_6802);
nand U7178 (N_7178,N_6062,N_6182);
nor U7179 (N_7179,N_6507,N_6934);
nor U7180 (N_7180,N_6314,N_6561);
nor U7181 (N_7181,N_6785,N_6403);
nor U7182 (N_7182,N_6696,N_6875);
nor U7183 (N_7183,N_6352,N_6752);
nor U7184 (N_7184,N_6493,N_6104);
and U7185 (N_7185,N_6840,N_6477);
xnor U7186 (N_7186,N_6757,N_6770);
or U7187 (N_7187,N_6007,N_6673);
or U7188 (N_7188,N_6129,N_6738);
or U7189 (N_7189,N_6252,N_6336);
nor U7190 (N_7190,N_6758,N_6029);
nand U7191 (N_7191,N_6337,N_6141);
xnor U7192 (N_7192,N_6277,N_6177);
nand U7193 (N_7193,N_6332,N_6256);
or U7194 (N_7194,N_6549,N_6273);
or U7195 (N_7195,N_6261,N_6197);
xor U7196 (N_7196,N_6172,N_6407);
or U7197 (N_7197,N_6955,N_6033);
nand U7198 (N_7198,N_6056,N_6364);
xor U7199 (N_7199,N_6354,N_6608);
and U7200 (N_7200,N_6452,N_6003);
xor U7201 (N_7201,N_6759,N_6618);
xor U7202 (N_7202,N_6717,N_6779);
xor U7203 (N_7203,N_6057,N_6409);
xnor U7204 (N_7204,N_6009,N_6484);
or U7205 (N_7205,N_6151,N_6147);
nor U7206 (N_7206,N_6333,N_6529);
or U7207 (N_7207,N_6843,N_6882);
nor U7208 (N_7208,N_6025,N_6035);
xnor U7209 (N_7209,N_6948,N_6015);
nor U7210 (N_7210,N_6995,N_6675);
and U7211 (N_7211,N_6378,N_6559);
nor U7212 (N_7212,N_6491,N_6411);
nor U7213 (N_7213,N_6839,N_6570);
nor U7214 (N_7214,N_6076,N_6709);
nand U7215 (N_7215,N_6422,N_6159);
nor U7216 (N_7216,N_6350,N_6872);
or U7217 (N_7217,N_6520,N_6650);
xor U7218 (N_7218,N_6956,N_6516);
nor U7219 (N_7219,N_6106,N_6339);
nand U7220 (N_7220,N_6879,N_6169);
or U7221 (N_7221,N_6417,N_6412);
nor U7222 (N_7222,N_6535,N_6615);
nor U7223 (N_7223,N_6763,N_6351);
nor U7224 (N_7224,N_6939,N_6464);
nor U7225 (N_7225,N_6899,N_6435);
or U7226 (N_7226,N_6328,N_6755);
nor U7227 (N_7227,N_6374,N_6795);
nand U7228 (N_7228,N_6444,N_6683);
nor U7229 (N_7229,N_6321,N_6228);
nand U7230 (N_7230,N_6584,N_6164);
nor U7231 (N_7231,N_6049,N_6012);
nor U7232 (N_7232,N_6171,N_6812);
nor U7233 (N_7233,N_6093,N_6249);
or U7234 (N_7234,N_6343,N_6384);
nand U7235 (N_7235,N_6474,N_6263);
and U7236 (N_7236,N_6883,N_6088);
nand U7237 (N_7237,N_6149,N_6099);
nand U7238 (N_7238,N_6744,N_6952);
xor U7239 (N_7239,N_6715,N_6748);
xor U7240 (N_7240,N_6741,N_6375);
nor U7241 (N_7241,N_6954,N_6648);
xor U7242 (N_7242,N_6156,N_6481);
or U7243 (N_7243,N_6876,N_6214);
or U7244 (N_7244,N_6130,N_6415);
nor U7245 (N_7245,N_6179,N_6946);
nand U7246 (N_7246,N_6923,N_6666);
xor U7247 (N_7247,N_6943,N_6756);
nand U7248 (N_7248,N_6132,N_6706);
and U7249 (N_7249,N_6863,N_6438);
and U7250 (N_7250,N_6067,N_6614);
nor U7251 (N_7251,N_6087,N_6115);
and U7252 (N_7252,N_6783,N_6789);
nor U7253 (N_7253,N_6991,N_6167);
xor U7254 (N_7254,N_6944,N_6200);
xnor U7255 (N_7255,N_6160,N_6041);
nand U7256 (N_7256,N_6722,N_6456);
or U7257 (N_7257,N_6047,N_6429);
xor U7258 (N_7258,N_6774,N_6659);
or U7259 (N_7259,N_6691,N_6714);
xnor U7260 (N_7260,N_6811,N_6898);
xnor U7261 (N_7261,N_6780,N_6804);
xor U7262 (N_7262,N_6368,N_6546);
or U7263 (N_7263,N_6264,N_6075);
or U7264 (N_7264,N_6108,N_6869);
and U7265 (N_7265,N_6024,N_6941);
or U7266 (N_7266,N_6937,N_6633);
and U7267 (N_7267,N_6284,N_6312);
nand U7268 (N_7268,N_6805,N_6639);
nor U7269 (N_7269,N_6851,N_6656);
and U7270 (N_7270,N_6377,N_6315);
xor U7271 (N_7271,N_6689,N_6419);
and U7272 (N_7272,N_6436,N_6086);
nor U7273 (N_7273,N_6836,N_6490);
or U7274 (N_7274,N_6157,N_6797);
nand U7275 (N_7275,N_6178,N_6233);
and U7276 (N_7276,N_6476,N_6008);
and U7277 (N_7277,N_6992,N_6070);
and U7278 (N_7278,N_6660,N_6761);
xor U7279 (N_7279,N_6001,N_6818);
nand U7280 (N_7280,N_6042,N_6276);
xor U7281 (N_7281,N_6402,N_6084);
or U7282 (N_7282,N_6282,N_6207);
nand U7283 (N_7283,N_6382,N_6153);
or U7284 (N_7284,N_6243,N_6211);
and U7285 (N_7285,N_6489,N_6248);
nand U7286 (N_7286,N_6513,N_6353);
or U7287 (N_7287,N_6950,N_6054);
and U7288 (N_7288,N_6238,N_6504);
xnor U7289 (N_7289,N_6281,N_6861);
or U7290 (N_7290,N_6305,N_6236);
nand U7291 (N_7291,N_6482,N_6330);
nor U7292 (N_7292,N_6932,N_6050);
and U7293 (N_7293,N_6707,N_6732);
nand U7294 (N_7294,N_6990,N_6307);
or U7295 (N_7295,N_6974,N_6695);
xnor U7296 (N_7296,N_6652,N_6460);
or U7297 (N_7297,N_6395,N_6338);
nand U7298 (N_7298,N_6257,N_6686);
xor U7299 (N_7299,N_6077,N_6136);
xor U7300 (N_7300,N_6066,N_6479);
and U7301 (N_7301,N_6829,N_6308);
xor U7302 (N_7302,N_6631,N_6269);
and U7303 (N_7303,N_6331,N_6320);
and U7304 (N_7304,N_6053,N_6705);
and U7305 (N_7305,N_6028,N_6373);
xor U7306 (N_7306,N_6886,N_6684);
or U7307 (N_7307,N_6971,N_6933);
xor U7308 (N_7308,N_6534,N_6773);
nor U7309 (N_7309,N_6716,N_6519);
or U7310 (N_7310,N_6502,N_6550);
nor U7311 (N_7311,N_6977,N_6002);
nand U7312 (N_7312,N_6963,N_6013);
nor U7313 (N_7313,N_6094,N_6753);
nand U7314 (N_7314,N_6517,N_6884);
xor U7315 (N_7315,N_6531,N_6000);
xor U7316 (N_7316,N_6349,N_6597);
and U7317 (N_7317,N_6645,N_6820);
or U7318 (N_7318,N_6310,N_6880);
and U7319 (N_7319,N_6388,N_6063);
and U7320 (N_7320,N_6860,N_6116);
nor U7321 (N_7321,N_6183,N_6085);
or U7322 (N_7322,N_6555,N_6449);
xnor U7323 (N_7323,N_6737,N_6914);
nand U7324 (N_7324,N_6170,N_6833);
and U7325 (N_7325,N_6293,N_6225);
xnor U7326 (N_7326,N_6609,N_6043);
nand U7327 (N_7327,N_6237,N_6165);
and U7328 (N_7328,N_6953,N_6272);
and U7329 (N_7329,N_6642,N_6110);
or U7330 (N_7330,N_6838,N_6126);
nor U7331 (N_7331,N_6124,N_6750);
or U7332 (N_7332,N_6036,N_6118);
nand U7333 (N_7333,N_6111,N_6796);
nor U7334 (N_7334,N_6887,N_6964);
nor U7335 (N_7335,N_6910,N_6215);
nor U7336 (N_7336,N_6103,N_6204);
or U7337 (N_7337,N_6278,N_6892);
nand U7338 (N_7338,N_6180,N_6583);
xor U7339 (N_7339,N_6468,N_6455);
nand U7340 (N_7340,N_6176,N_6734);
nor U7341 (N_7341,N_6747,N_6510);
and U7342 (N_7342,N_6380,N_6120);
or U7343 (N_7343,N_6302,N_6585);
nand U7344 (N_7344,N_6595,N_6044);
nor U7345 (N_7345,N_6568,N_6341);
nand U7346 (N_7346,N_6262,N_6589);
xnor U7347 (N_7347,N_6433,N_6201);
xor U7348 (N_7348,N_6629,N_6856);
nor U7349 (N_7349,N_6295,N_6808);
xor U7350 (N_7350,N_6100,N_6921);
nand U7351 (N_7351,N_6965,N_6834);
nor U7352 (N_7352,N_6434,N_6500);
or U7353 (N_7353,N_6022,N_6749);
or U7354 (N_7354,N_6657,N_6929);
xnor U7355 (N_7355,N_6071,N_6778);
or U7356 (N_7356,N_6347,N_6286);
nand U7357 (N_7357,N_6945,N_6859);
and U7358 (N_7358,N_6591,N_6871);
xor U7359 (N_7359,N_6210,N_6699);
nor U7360 (N_7360,N_6285,N_6931);
or U7361 (N_7361,N_6509,N_6745);
and U7362 (N_7362,N_6746,N_6810);
nand U7363 (N_7363,N_6994,N_6250);
nor U7364 (N_7364,N_6538,N_6727);
or U7365 (N_7365,N_6612,N_6231);
nand U7366 (N_7366,N_6815,N_6381);
or U7367 (N_7367,N_6485,N_6607);
or U7368 (N_7368,N_6472,N_6866);
and U7369 (N_7369,N_6251,N_6487);
and U7370 (N_7370,N_6483,N_6610);
xnor U7371 (N_7371,N_6641,N_6729);
nand U7372 (N_7372,N_6023,N_6765);
or U7373 (N_7373,N_6039,N_6740);
or U7374 (N_7374,N_6653,N_6544);
nor U7375 (N_7375,N_6743,N_6298);
xor U7376 (N_7376,N_6301,N_6279);
nor U7377 (N_7377,N_6495,N_6970);
or U7378 (N_7378,N_6416,N_6125);
and U7379 (N_7379,N_6306,N_6621);
or U7380 (N_7380,N_6575,N_6720);
or U7381 (N_7381,N_6397,N_6827);
and U7382 (N_7382,N_6551,N_6809);
nor U7383 (N_7383,N_6420,N_6724);
xnor U7384 (N_7384,N_6649,N_6674);
xnor U7385 (N_7385,N_6957,N_6131);
or U7386 (N_7386,N_6370,N_6016);
or U7387 (N_7387,N_6846,N_6329);
xor U7388 (N_7388,N_6234,N_6418);
nor U7389 (N_7389,N_6525,N_6972);
nand U7390 (N_7390,N_6127,N_6793);
nand U7391 (N_7391,N_6893,N_6771);
nand U7392 (N_7392,N_6912,N_6345);
and U7393 (N_7393,N_6764,N_6799);
and U7394 (N_7394,N_6915,N_6083);
and U7395 (N_7395,N_6547,N_6119);
or U7396 (N_7396,N_6526,N_6508);
nand U7397 (N_7397,N_6073,N_6404);
xnor U7398 (N_7398,N_6989,N_6133);
nand U7399 (N_7399,N_6045,N_6518);
nor U7400 (N_7400,N_6976,N_6890);
nand U7401 (N_7401,N_6095,N_6348);
and U7402 (N_7402,N_6665,N_6459);
xnor U7403 (N_7403,N_6475,N_6018);
or U7404 (N_7404,N_6635,N_6530);
or U7405 (N_7405,N_6040,N_6701);
and U7406 (N_7406,N_6847,N_6437);
nor U7407 (N_7407,N_6163,N_6297);
nand U7408 (N_7408,N_6203,N_6598);
xor U7409 (N_7409,N_6754,N_6951);
xor U7410 (N_7410,N_6152,N_6304);
nor U7411 (N_7411,N_6623,N_6274);
nand U7412 (N_7412,N_6558,N_6668);
or U7413 (N_7413,N_6918,N_6949);
nor U7414 (N_7414,N_6240,N_6854);
xnor U7415 (N_7415,N_6935,N_6562);
or U7416 (N_7416,N_6218,N_6794);
or U7417 (N_7417,N_6895,N_6166);
xor U7418 (N_7418,N_6254,N_6572);
and U7419 (N_7419,N_6253,N_6619);
or U7420 (N_7420,N_6371,N_6586);
nand U7421 (N_7421,N_6900,N_6241);
and U7422 (N_7422,N_6781,N_6466);
nor U7423 (N_7423,N_6581,N_6090);
nor U7424 (N_7424,N_6142,N_6046);
or U7425 (N_7425,N_6606,N_6208);
and U7426 (N_7426,N_6806,N_6432);
nand U7427 (N_7427,N_6702,N_6392);
and U7428 (N_7428,N_6959,N_6848);
and U7429 (N_7429,N_6198,N_6026);
nand U7430 (N_7430,N_6579,N_6267);
and U7431 (N_7431,N_6926,N_6993);
and U7432 (N_7432,N_6005,N_6017);
nor U7433 (N_7433,N_6888,N_6399);
nor U7434 (N_7434,N_6703,N_6850);
or U7435 (N_7435,N_6553,N_6678);
xor U7436 (N_7436,N_6620,N_6098);
nand U7437 (N_7437,N_6830,N_6398);
nand U7438 (N_7438,N_6638,N_6072);
nor U7439 (N_7439,N_6255,N_6199);
or U7440 (N_7440,N_6988,N_6360);
and U7441 (N_7441,N_6443,N_6450);
nor U7442 (N_7442,N_6791,N_6868);
nand U7443 (N_7443,N_6342,N_6894);
nor U7444 (N_7444,N_6283,N_6089);
and U7445 (N_7445,N_6247,N_6593);
or U7446 (N_7446,N_6383,N_6150);
nor U7447 (N_7447,N_6690,N_6997);
xor U7448 (N_7448,N_6358,N_6985);
nand U7449 (N_7449,N_6019,N_6511);
and U7450 (N_7450,N_6258,N_6498);
nand U7451 (N_7451,N_6501,N_6317);
and U7452 (N_7452,N_6733,N_6117);
and U7453 (N_7453,N_6096,N_6445);
nor U7454 (N_7454,N_6410,N_6698);
nor U7455 (N_7455,N_6896,N_6451);
or U7456 (N_7456,N_6471,N_6677);
xnor U7457 (N_7457,N_6280,N_6082);
nor U7458 (N_7458,N_6454,N_6143);
nand U7459 (N_7459,N_6580,N_6196);
and U7460 (N_7460,N_6837,N_6592);
xnor U7461 (N_7461,N_6938,N_6543);
and U7462 (N_7462,N_6819,N_6711);
nor U7463 (N_7463,N_6413,N_6751);
and U7464 (N_7464,N_6123,N_6387);
nor U7465 (N_7465,N_6442,N_6222);
and U7466 (N_7466,N_6643,N_6134);
xnor U7467 (N_7467,N_6318,N_6430);
or U7468 (N_7468,N_6655,N_6919);
nand U7469 (N_7469,N_6367,N_6792);
xnor U7470 (N_7470,N_6556,N_6423);
and U7471 (N_7471,N_6769,N_6376);
and U7472 (N_7472,N_6154,N_6068);
nand U7473 (N_7473,N_6031,N_6557);
xnor U7474 (N_7474,N_6461,N_6109);
and U7475 (N_7475,N_6905,N_6712);
or U7476 (N_7476,N_6790,N_6356);
nor U7477 (N_7477,N_6217,N_6457);
nand U7478 (N_7478,N_6613,N_6924);
nor U7479 (N_7479,N_6611,N_6271);
nand U7480 (N_7480,N_6344,N_6590);
nand U7481 (N_7481,N_6725,N_6193);
xor U7482 (N_7482,N_6059,N_6920);
nor U7483 (N_7483,N_6842,N_6522);
nor U7484 (N_7484,N_6560,N_6841);
nor U7485 (N_7485,N_6112,N_6048);
xor U7486 (N_7486,N_6852,N_6334);
nand U7487 (N_7487,N_6624,N_6428);
xor U7488 (N_7488,N_6158,N_6221);
xnor U7489 (N_7489,N_6569,N_6266);
and U7490 (N_7490,N_6326,N_6440);
xnor U7491 (N_7491,N_6680,N_6365);
nor U7492 (N_7492,N_6835,N_6324);
or U7493 (N_7493,N_6372,N_6760);
nor U7494 (N_7494,N_6782,N_6646);
xor U7495 (N_7495,N_6168,N_6426);
or U7496 (N_7496,N_6800,N_6004);
and U7497 (N_7497,N_6907,N_6414);
or U7498 (N_7498,N_6700,N_6958);
and U7499 (N_7499,N_6925,N_6803);
nor U7500 (N_7500,N_6167,N_6985);
or U7501 (N_7501,N_6403,N_6356);
nor U7502 (N_7502,N_6353,N_6051);
or U7503 (N_7503,N_6829,N_6703);
nand U7504 (N_7504,N_6116,N_6091);
and U7505 (N_7505,N_6383,N_6956);
or U7506 (N_7506,N_6615,N_6020);
and U7507 (N_7507,N_6812,N_6498);
or U7508 (N_7508,N_6391,N_6205);
or U7509 (N_7509,N_6371,N_6866);
and U7510 (N_7510,N_6777,N_6918);
or U7511 (N_7511,N_6695,N_6259);
nand U7512 (N_7512,N_6823,N_6838);
or U7513 (N_7513,N_6788,N_6954);
nand U7514 (N_7514,N_6932,N_6856);
xor U7515 (N_7515,N_6725,N_6353);
or U7516 (N_7516,N_6982,N_6852);
xor U7517 (N_7517,N_6332,N_6603);
and U7518 (N_7518,N_6522,N_6676);
and U7519 (N_7519,N_6381,N_6233);
nand U7520 (N_7520,N_6646,N_6522);
and U7521 (N_7521,N_6174,N_6134);
nor U7522 (N_7522,N_6067,N_6733);
xor U7523 (N_7523,N_6393,N_6851);
nand U7524 (N_7524,N_6375,N_6747);
nor U7525 (N_7525,N_6966,N_6102);
and U7526 (N_7526,N_6522,N_6563);
and U7527 (N_7527,N_6647,N_6381);
and U7528 (N_7528,N_6282,N_6883);
and U7529 (N_7529,N_6835,N_6032);
or U7530 (N_7530,N_6325,N_6973);
nor U7531 (N_7531,N_6316,N_6665);
or U7532 (N_7532,N_6283,N_6806);
nand U7533 (N_7533,N_6643,N_6934);
or U7534 (N_7534,N_6693,N_6034);
or U7535 (N_7535,N_6967,N_6764);
nor U7536 (N_7536,N_6418,N_6465);
or U7537 (N_7537,N_6465,N_6390);
or U7538 (N_7538,N_6779,N_6791);
nor U7539 (N_7539,N_6515,N_6447);
or U7540 (N_7540,N_6990,N_6871);
nor U7541 (N_7541,N_6815,N_6058);
nor U7542 (N_7542,N_6976,N_6684);
nand U7543 (N_7543,N_6344,N_6866);
and U7544 (N_7544,N_6964,N_6205);
xor U7545 (N_7545,N_6327,N_6753);
nand U7546 (N_7546,N_6954,N_6385);
nand U7547 (N_7547,N_6766,N_6897);
xor U7548 (N_7548,N_6391,N_6629);
and U7549 (N_7549,N_6057,N_6347);
or U7550 (N_7550,N_6772,N_6730);
or U7551 (N_7551,N_6030,N_6777);
xor U7552 (N_7552,N_6956,N_6047);
xor U7553 (N_7553,N_6558,N_6127);
xnor U7554 (N_7554,N_6934,N_6191);
or U7555 (N_7555,N_6075,N_6699);
and U7556 (N_7556,N_6582,N_6409);
or U7557 (N_7557,N_6160,N_6272);
or U7558 (N_7558,N_6423,N_6802);
nor U7559 (N_7559,N_6306,N_6311);
or U7560 (N_7560,N_6995,N_6433);
or U7561 (N_7561,N_6167,N_6846);
nand U7562 (N_7562,N_6809,N_6649);
nor U7563 (N_7563,N_6984,N_6286);
nor U7564 (N_7564,N_6778,N_6990);
nand U7565 (N_7565,N_6119,N_6579);
and U7566 (N_7566,N_6412,N_6141);
or U7567 (N_7567,N_6219,N_6343);
or U7568 (N_7568,N_6490,N_6594);
and U7569 (N_7569,N_6536,N_6305);
or U7570 (N_7570,N_6943,N_6561);
or U7571 (N_7571,N_6419,N_6618);
nand U7572 (N_7572,N_6078,N_6618);
or U7573 (N_7573,N_6075,N_6798);
and U7574 (N_7574,N_6745,N_6044);
nand U7575 (N_7575,N_6997,N_6000);
nand U7576 (N_7576,N_6793,N_6074);
and U7577 (N_7577,N_6466,N_6192);
nand U7578 (N_7578,N_6089,N_6229);
and U7579 (N_7579,N_6499,N_6150);
or U7580 (N_7580,N_6851,N_6748);
xnor U7581 (N_7581,N_6841,N_6147);
nand U7582 (N_7582,N_6842,N_6388);
and U7583 (N_7583,N_6269,N_6193);
or U7584 (N_7584,N_6296,N_6910);
xnor U7585 (N_7585,N_6732,N_6272);
and U7586 (N_7586,N_6877,N_6870);
nand U7587 (N_7587,N_6007,N_6418);
nor U7588 (N_7588,N_6755,N_6442);
nand U7589 (N_7589,N_6308,N_6157);
or U7590 (N_7590,N_6173,N_6492);
or U7591 (N_7591,N_6700,N_6367);
and U7592 (N_7592,N_6142,N_6927);
nand U7593 (N_7593,N_6824,N_6279);
nand U7594 (N_7594,N_6713,N_6091);
nand U7595 (N_7595,N_6600,N_6241);
and U7596 (N_7596,N_6767,N_6107);
or U7597 (N_7597,N_6343,N_6266);
nand U7598 (N_7598,N_6419,N_6925);
and U7599 (N_7599,N_6267,N_6435);
nand U7600 (N_7600,N_6151,N_6370);
nor U7601 (N_7601,N_6919,N_6806);
xor U7602 (N_7602,N_6026,N_6024);
nor U7603 (N_7603,N_6444,N_6633);
or U7604 (N_7604,N_6433,N_6200);
and U7605 (N_7605,N_6160,N_6583);
and U7606 (N_7606,N_6740,N_6097);
xnor U7607 (N_7607,N_6258,N_6455);
nand U7608 (N_7608,N_6451,N_6166);
and U7609 (N_7609,N_6438,N_6490);
nor U7610 (N_7610,N_6032,N_6344);
or U7611 (N_7611,N_6196,N_6334);
or U7612 (N_7612,N_6016,N_6699);
nand U7613 (N_7613,N_6185,N_6453);
xnor U7614 (N_7614,N_6050,N_6327);
and U7615 (N_7615,N_6981,N_6006);
nor U7616 (N_7616,N_6383,N_6208);
and U7617 (N_7617,N_6398,N_6567);
and U7618 (N_7618,N_6902,N_6516);
xor U7619 (N_7619,N_6132,N_6099);
nand U7620 (N_7620,N_6900,N_6650);
or U7621 (N_7621,N_6609,N_6683);
nor U7622 (N_7622,N_6621,N_6758);
or U7623 (N_7623,N_6299,N_6745);
nor U7624 (N_7624,N_6912,N_6355);
nor U7625 (N_7625,N_6579,N_6598);
xnor U7626 (N_7626,N_6750,N_6386);
or U7627 (N_7627,N_6693,N_6328);
and U7628 (N_7628,N_6219,N_6526);
nor U7629 (N_7629,N_6954,N_6742);
nor U7630 (N_7630,N_6721,N_6338);
nor U7631 (N_7631,N_6974,N_6275);
xnor U7632 (N_7632,N_6168,N_6450);
xnor U7633 (N_7633,N_6833,N_6343);
nor U7634 (N_7634,N_6470,N_6749);
nand U7635 (N_7635,N_6267,N_6117);
nor U7636 (N_7636,N_6905,N_6316);
or U7637 (N_7637,N_6766,N_6922);
and U7638 (N_7638,N_6270,N_6380);
xor U7639 (N_7639,N_6584,N_6831);
nand U7640 (N_7640,N_6116,N_6581);
nor U7641 (N_7641,N_6576,N_6532);
nand U7642 (N_7642,N_6186,N_6552);
or U7643 (N_7643,N_6462,N_6848);
xnor U7644 (N_7644,N_6775,N_6227);
nand U7645 (N_7645,N_6368,N_6198);
xnor U7646 (N_7646,N_6859,N_6185);
nand U7647 (N_7647,N_6422,N_6482);
nand U7648 (N_7648,N_6988,N_6639);
or U7649 (N_7649,N_6857,N_6257);
and U7650 (N_7650,N_6277,N_6007);
nor U7651 (N_7651,N_6730,N_6793);
and U7652 (N_7652,N_6925,N_6825);
nor U7653 (N_7653,N_6712,N_6430);
and U7654 (N_7654,N_6807,N_6599);
or U7655 (N_7655,N_6587,N_6934);
and U7656 (N_7656,N_6708,N_6981);
and U7657 (N_7657,N_6396,N_6657);
xor U7658 (N_7658,N_6689,N_6722);
or U7659 (N_7659,N_6379,N_6604);
nor U7660 (N_7660,N_6783,N_6753);
xnor U7661 (N_7661,N_6668,N_6580);
nor U7662 (N_7662,N_6076,N_6961);
and U7663 (N_7663,N_6764,N_6224);
xor U7664 (N_7664,N_6272,N_6595);
and U7665 (N_7665,N_6276,N_6289);
nand U7666 (N_7666,N_6827,N_6880);
nor U7667 (N_7667,N_6862,N_6353);
nand U7668 (N_7668,N_6528,N_6219);
or U7669 (N_7669,N_6705,N_6374);
xnor U7670 (N_7670,N_6330,N_6149);
nand U7671 (N_7671,N_6680,N_6383);
xnor U7672 (N_7672,N_6458,N_6974);
and U7673 (N_7673,N_6252,N_6040);
xnor U7674 (N_7674,N_6078,N_6282);
nand U7675 (N_7675,N_6960,N_6188);
or U7676 (N_7676,N_6454,N_6152);
xnor U7677 (N_7677,N_6382,N_6307);
or U7678 (N_7678,N_6119,N_6570);
and U7679 (N_7679,N_6692,N_6277);
or U7680 (N_7680,N_6155,N_6132);
xnor U7681 (N_7681,N_6322,N_6999);
or U7682 (N_7682,N_6078,N_6847);
xnor U7683 (N_7683,N_6601,N_6429);
nor U7684 (N_7684,N_6969,N_6772);
xor U7685 (N_7685,N_6920,N_6946);
nor U7686 (N_7686,N_6298,N_6231);
or U7687 (N_7687,N_6951,N_6116);
xor U7688 (N_7688,N_6688,N_6488);
or U7689 (N_7689,N_6636,N_6518);
or U7690 (N_7690,N_6299,N_6837);
and U7691 (N_7691,N_6718,N_6280);
nand U7692 (N_7692,N_6240,N_6440);
and U7693 (N_7693,N_6136,N_6790);
nor U7694 (N_7694,N_6051,N_6810);
xnor U7695 (N_7695,N_6987,N_6960);
nor U7696 (N_7696,N_6836,N_6166);
xor U7697 (N_7697,N_6698,N_6186);
nor U7698 (N_7698,N_6916,N_6478);
nor U7699 (N_7699,N_6853,N_6520);
nor U7700 (N_7700,N_6358,N_6602);
and U7701 (N_7701,N_6558,N_6555);
xor U7702 (N_7702,N_6856,N_6926);
or U7703 (N_7703,N_6466,N_6213);
nor U7704 (N_7704,N_6231,N_6441);
nand U7705 (N_7705,N_6715,N_6368);
or U7706 (N_7706,N_6977,N_6309);
and U7707 (N_7707,N_6439,N_6400);
and U7708 (N_7708,N_6885,N_6768);
and U7709 (N_7709,N_6179,N_6804);
nand U7710 (N_7710,N_6925,N_6863);
nand U7711 (N_7711,N_6399,N_6367);
nor U7712 (N_7712,N_6253,N_6441);
or U7713 (N_7713,N_6562,N_6400);
and U7714 (N_7714,N_6499,N_6767);
and U7715 (N_7715,N_6667,N_6723);
and U7716 (N_7716,N_6180,N_6430);
xor U7717 (N_7717,N_6900,N_6518);
or U7718 (N_7718,N_6305,N_6917);
nand U7719 (N_7719,N_6280,N_6744);
nor U7720 (N_7720,N_6098,N_6357);
nand U7721 (N_7721,N_6996,N_6543);
nor U7722 (N_7722,N_6098,N_6984);
and U7723 (N_7723,N_6986,N_6577);
xor U7724 (N_7724,N_6725,N_6175);
xor U7725 (N_7725,N_6536,N_6945);
or U7726 (N_7726,N_6444,N_6766);
or U7727 (N_7727,N_6980,N_6163);
nor U7728 (N_7728,N_6382,N_6425);
nand U7729 (N_7729,N_6063,N_6317);
and U7730 (N_7730,N_6127,N_6332);
or U7731 (N_7731,N_6927,N_6822);
and U7732 (N_7732,N_6111,N_6719);
nor U7733 (N_7733,N_6207,N_6932);
nor U7734 (N_7734,N_6373,N_6300);
or U7735 (N_7735,N_6740,N_6464);
and U7736 (N_7736,N_6346,N_6883);
and U7737 (N_7737,N_6420,N_6761);
xor U7738 (N_7738,N_6250,N_6889);
and U7739 (N_7739,N_6652,N_6432);
nand U7740 (N_7740,N_6063,N_6657);
nor U7741 (N_7741,N_6838,N_6578);
or U7742 (N_7742,N_6694,N_6947);
xnor U7743 (N_7743,N_6303,N_6523);
or U7744 (N_7744,N_6114,N_6862);
nand U7745 (N_7745,N_6434,N_6274);
nand U7746 (N_7746,N_6729,N_6867);
or U7747 (N_7747,N_6463,N_6705);
or U7748 (N_7748,N_6368,N_6772);
xor U7749 (N_7749,N_6488,N_6709);
nor U7750 (N_7750,N_6079,N_6636);
nand U7751 (N_7751,N_6730,N_6650);
nand U7752 (N_7752,N_6086,N_6793);
xnor U7753 (N_7753,N_6424,N_6676);
or U7754 (N_7754,N_6682,N_6514);
or U7755 (N_7755,N_6273,N_6664);
nand U7756 (N_7756,N_6654,N_6384);
or U7757 (N_7757,N_6349,N_6619);
nor U7758 (N_7758,N_6212,N_6746);
and U7759 (N_7759,N_6548,N_6021);
nand U7760 (N_7760,N_6168,N_6858);
or U7761 (N_7761,N_6708,N_6310);
xor U7762 (N_7762,N_6850,N_6476);
nand U7763 (N_7763,N_6946,N_6408);
nor U7764 (N_7764,N_6344,N_6453);
xnor U7765 (N_7765,N_6460,N_6845);
and U7766 (N_7766,N_6179,N_6108);
or U7767 (N_7767,N_6620,N_6190);
and U7768 (N_7768,N_6564,N_6790);
and U7769 (N_7769,N_6164,N_6753);
nor U7770 (N_7770,N_6295,N_6353);
nor U7771 (N_7771,N_6752,N_6866);
and U7772 (N_7772,N_6983,N_6846);
nand U7773 (N_7773,N_6200,N_6898);
and U7774 (N_7774,N_6704,N_6172);
nand U7775 (N_7775,N_6881,N_6817);
xor U7776 (N_7776,N_6199,N_6078);
and U7777 (N_7777,N_6405,N_6421);
nand U7778 (N_7778,N_6655,N_6621);
and U7779 (N_7779,N_6301,N_6715);
xor U7780 (N_7780,N_6589,N_6930);
or U7781 (N_7781,N_6939,N_6123);
nand U7782 (N_7782,N_6161,N_6075);
or U7783 (N_7783,N_6646,N_6924);
nor U7784 (N_7784,N_6083,N_6332);
and U7785 (N_7785,N_6386,N_6526);
or U7786 (N_7786,N_6042,N_6086);
and U7787 (N_7787,N_6474,N_6448);
nand U7788 (N_7788,N_6257,N_6151);
nand U7789 (N_7789,N_6325,N_6031);
nand U7790 (N_7790,N_6597,N_6123);
nand U7791 (N_7791,N_6518,N_6207);
nand U7792 (N_7792,N_6430,N_6230);
xor U7793 (N_7793,N_6383,N_6388);
or U7794 (N_7794,N_6639,N_6656);
nor U7795 (N_7795,N_6572,N_6500);
xor U7796 (N_7796,N_6360,N_6943);
xnor U7797 (N_7797,N_6175,N_6766);
and U7798 (N_7798,N_6825,N_6420);
nand U7799 (N_7799,N_6005,N_6445);
xor U7800 (N_7800,N_6542,N_6688);
and U7801 (N_7801,N_6226,N_6181);
xnor U7802 (N_7802,N_6294,N_6037);
nor U7803 (N_7803,N_6328,N_6625);
and U7804 (N_7804,N_6828,N_6466);
nor U7805 (N_7805,N_6888,N_6254);
and U7806 (N_7806,N_6698,N_6136);
nand U7807 (N_7807,N_6696,N_6233);
nor U7808 (N_7808,N_6294,N_6140);
nor U7809 (N_7809,N_6411,N_6401);
and U7810 (N_7810,N_6640,N_6626);
and U7811 (N_7811,N_6832,N_6189);
nor U7812 (N_7812,N_6118,N_6856);
and U7813 (N_7813,N_6065,N_6205);
or U7814 (N_7814,N_6352,N_6944);
nand U7815 (N_7815,N_6337,N_6217);
xor U7816 (N_7816,N_6338,N_6377);
and U7817 (N_7817,N_6027,N_6147);
nand U7818 (N_7818,N_6251,N_6792);
and U7819 (N_7819,N_6680,N_6851);
nor U7820 (N_7820,N_6125,N_6027);
and U7821 (N_7821,N_6538,N_6298);
and U7822 (N_7822,N_6825,N_6976);
xnor U7823 (N_7823,N_6253,N_6462);
xnor U7824 (N_7824,N_6180,N_6382);
nand U7825 (N_7825,N_6755,N_6421);
nor U7826 (N_7826,N_6110,N_6407);
or U7827 (N_7827,N_6094,N_6858);
nor U7828 (N_7828,N_6909,N_6943);
and U7829 (N_7829,N_6570,N_6565);
nor U7830 (N_7830,N_6176,N_6781);
xor U7831 (N_7831,N_6177,N_6818);
and U7832 (N_7832,N_6775,N_6042);
nand U7833 (N_7833,N_6034,N_6690);
nand U7834 (N_7834,N_6539,N_6070);
xor U7835 (N_7835,N_6692,N_6354);
and U7836 (N_7836,N_6223,N_6188);
nand U7837 (N_7837,N_6224,N_6087);
xnor U7838 (N_7838,N_6708,N_6274);
or U7839 (N_7839,N_6390,N_6878);
nor U7840 (N_7840,N_6886,N_6519);
nand U7841 (N_7841,N_6539,N_6455);
or U7842 (N_7842,N_6865,N_6473);
or U7843 (N_7843,N_6282,N_6114);
and U7844 (N_7844,N_6687,N_6115);
xor U7845 (N_7845,N_6294,N_6086);
xnor U7846 (N_7846,N_6990,N_6552);
xor U7847 (N_7847,N_6342,N_6322);
and U7848 (N_7848,N_6656,N_6829);
nand U7849 (N_7849,N_6402,N_6539);
xnor U7850 (N_7850,N_6049,N_6204);
nor U7851 (N_7851,N_6474,N_6769);
and U7852 (N_7852,N_6399,N_6785);
xnor U7853 (N_7853,N_6543,N_6986);
xor U7854 (N_7854,N_6232,N_6699);
nor U7855 (N_7855,N_6606,N_6366);
xnor U7856 (N_7856,N_6759,N_6813);
nor U7857 (N_7857,N_6955,N_6880);
and U7858 (N_7858,N_6795,N_6476);
xor U7859 (N_7859,N_6171,N_6612);
or U7860 (N_7860,N_6096,N_6816);
xor U7861 (N_7861,N_6341,N_6265);
xnor U7862 (N_7862,N_6131,N_6467);
nor U7863 (N_7863,N_6833,N_6865);
nor U7864 (N_7864,N_6577,N_6193);
xor U7865 (N_7865,N_6405,N_6196);
nand U7866 (N_7866,N_6148,N_6635);
nand U7867 (N_7867,N_6619,N_6492);
or U7868 (N_7868,N_6675,N_6971);
and U7869 (N_7869,N_6688,N_6537);
or U7870 (N_7870,N_6282,N_6712);
nor U7871 (N_7871,N_6912,N_6236);
nor U7872 (N_7872,N_6544,N_6320);
nor U7873 (N_7873,N_6017,N_6141);
and U7874 (N_7874,N_6428,N_6590);
or U7875 (N_7875,N_6843,N_6860);
xor U7876 (N_7876,N_6021,N_6608);
or U7877 (N_7877,N_6537,N_6841);
nor U7878 (N_7878,N_6346,N_6464);
or U7879 (N_7879,N_6427,N_6312);
xor U7880 (N_7880,N_6819,N_6619);
or U7881 (N_7881,N_6676,N_6034);
or U7882 (N_7882,N_6125,N_6128);
xnor U7883 (N_7883,N_6331,N_6998);
or U7884 (N_7884,N_6231,N_6794);
nor U7885 (N_7885,N_6849,N_6943);
nand U7886 (N_7886,N_6889,N_6816);
nand U7887 (N_7887,N_6740,N_6126);
nor U7888 (N_7888,N_6210,N_6033);
nor U7889 (N_7889,N_6963,N_6918);
nor U7890 (N_7890,N_6141,N_6547);
xnor U7891 (N_7891,N_6218,N_6223);
xor U7892 (N_7892,N_6243,N_6466);
and U7893 (N_7893,N_6678,N_6425);
xnor U7894 (N_7894,N_6607,N_6660);
nor U7895 (N_7895,N_6314,N_6318);
and U7896 (N_7896,N_6685,N_6349);
and U7897 (N_7897,N_6552,N_6946);
xnor U7898 (N_7898,N_6071,N_6050);
and U7899 (N_7899,N_6944,N_6772);
and U7900 (N_7900,N_6829,N_6171);
xor U7901 (N_7901,N_6725,N_6517);
and U7902 (N_7902,N_6336,N_6836);
nor U7903 (N_7903,N_6886,N_6731);
nand U7904 (N_7904,N_6728,N_6363);
nor U7905 (N_7905,N_6326,N_6571);
nand U7906 (N_7906,N_6938,N_6961);
nand U7907 (N_7907,N_6886,N_6195);
or U7908 (N_7908,N_6387,N_6667);
and U7909 (N_7909,N_6528,N_6692);
nor U7910 (N_7910,N_6222,N_6792);
nand U7911 (N_7911,N_6539,N_6515);
nor U7912 (N_7912,N_6424,N_6357);
or U7913 (N_7913,N_6808,N_6310);
and U7914 (N_7914,N_6005,N_6586);
nor U7915 (N_7915,N_6170,N_6183);
nor U7916 (N_7916,N_6238,N_6172);
xor U7917 (N_7917,N_6524,N_6375);
and U7918 (N_7918,N_6054,N_6899);
nor U7919 (N_7919,N_6478,N_6127);
nand U7920 (N_7920,N_6528,N_6982);
and U7921 (N_7921,N_6992,N_6306);
xor U7922 (N_7922,N_6942,N_6473);
nand U7923 (N_7923,N_6950,N_6242);
nor U7924 (N_7924,N_6273,N_6268);
nand U7925 (N_7925,N_6785,N_6569);
and U7926 (N_7926,N_6277,N_6160);
nor U7927 (N_7927,N_6909,N_6356);
nand U7928 (N_7928,N_6438,N_6245);
xor U7929 (N_7929,N_6777,N_6937);
or U7930 (N_7930,N_6780,N_6365);
xor U7931 (N_7931,N_6426,N_6121);
and U7932 (N_7932,N_6949,N_6590);
and U7933 (N_7933,N_6305,N_6130);
nor U7934 (N_7934,N_6417,N_6823);
and U7935 (N_7935,N_6920,N_6807);
nor U7936 (N_7936,N_6447,N_6631);
nor U7937 (N_7937,N_6284,N_6135);
xor U7938 (N_7938,N_6247,N_6459);
xnor U7939 (N_7939,N_6906,N_6649);
nor U7940 (N_7940,N_6608,N_6173);
nor U7941 (N_7941,N_6929,N_6143);
nand U7942 (N_7942,N_6221,N_6714);
xnor U7943 (N_7943,N_6957,N_6521);
or U7944 (N_7944,N_6929,N_6271);
nor U7945 (N_7945,N_6592,N_6603);
nand U7946 (N_7946,N_6488,N_6287);
or U7947 (N_7947,N_6620,N_6825);
and U7948 (N_7948,N_6371,N_6438);
nand U7949 (N_7949,N_6826,N_6735);
xnor U7950 (N_7950,N_6070,N_6317);
and U7951 (N_7951,N_6608,N_6899);
and U7952 (N_7952,N_6520,N_6132);
nor U7953 (N_7953,N_6094,N_6207);
nor U7954 (N_7954,N_6821,N_6887);
xor U7955 (N_7955,N_6242,N_6727);
and U7956 (N_7956,N_6680,N_6195);
or U7957 (N_7957,N_6667,N_6441);
nor U7958 (N_7958,N_6804,N_6066);
and U7959 (N_7959,N_6143,N_6887);
or U7960 (N_7960,N_6814,N_6745);
and U7961 (N_7961,N_6913,N_6934);
nor U7962 (N_7962,N_6029,N_6992);
xor U7963 (N_7963,N_6415,N_6933);
nor U7964 (N_7964,N_6857,N_6085);
xnor U7965 (N_7965,N_6079,N_6188);
or U7966 (N_7966,N_6326,N_6123);
nor U7967 (N_7967,N_6149,N_6209);
and U7968 (N_7968,N_6413,N_6726);
nor U7969 (N_7969,N_6689,N_6681);
nand U7970 (N_7970,N_6158,N_6389);
or U7971 (N_7971,N_6260,N_6852);
and U7972 (N_7972,N_6939,N_6482);
and U7973 (N_7973,N_6625,N_6282);
or U7974 (N_7974,N_6499,N_6936);
or U7975 (N_7975,N_6605,N_6430);
nand U7976 (N_7976,N_6931,N_6761);
or U7977 (N_7977,N_6967,N_6195);
nor U7978 (N_7978,N_6865,N_6536);
nand U7979 (N_7979,N_6871,N_6835);
and U7980 (N_7980,N_6355,N_6621);
nand U7981 (N_7981,N_6447,N_6858);
xnor U7982 (N_7982,N_6654,N_6247);
or U7983 (N_7983,N_6348,N_6667);
or U7984 (N_7984,N_6717,N_6056);
xor U7985 (N_7985,N_6435,N_6724);
nor U7986 (N_7986,N_6386,N_6491);
and U7987 (N_7987,N_6643,N_6586);
xnor U7988 (N_7988,N_6293,N_6086);
and U7989 (N_7989,N_6973,N_6394);
xor U7990 (N_7990,N_6893,N_6935);
nor U7991 (N_7991,N_6799,N_6569);
xnor U7992 (N_7992,N_6386,N_6190);
xnor U7993 (N_7993,N_6296,N_6456);
xnor U7994 (N_7994,N_6276,N_6405);
nor U7995 (N_7995,N_6045,N_6552);
nand U7996 (N_7996,N_6860,N_6694);
xnor U7997 (N_7997,N_6769,N_6650);
xor U7998 (N_7998,N_6565,N_6960);
nor U7999 (N_7999,N_6698,N_6563);
nor U8000 (N_8000,N_7667,N_7002);
nand U8001 (N_8001,N_7124,N_7337);
and U8002 (N_8002,N_7536,N_7292);
and U8003 (N_8003,N_7024,N_7349);
nand U8004 (N_8004,N_7128,N_7638);
xor U8005 (N_8005,N_7906,N_7261);
nand U8006 (N_8006,N_7407,N_7262);
xnor U8007 (N_8007,N_7937,N_7230);
or U8008 (N_8008,N_7883,N_7926);
xnor U8009 (N_8009,N_7988,N_7466);
and U8010 (N_8010,N_7393,N_7049);
nor U8011 (N_8011,N_7963,N_7138);
or U8012 (N_8012,N_7485,N_7625);
xnor U8013 (N_8013,N_7998,N_7192);
xor U8014 (N_8014,N_7175,N_7953);
or U8015 (N_8015,N_7809,N_7389);
nand U8016 (N_8016,N_7641,N_7981);
nand U8017 (N_8017,N_7879,N_7609);
xor U8018 (N_8018,N_7721,N_7909);
nand U8019 (N_8019,N_7283,N_7557);
nor U8020 (N_8020,N_7312,N_7394);
nor U8021 (N_8021,N_7488,N_7975);
and U8022 (N_8022,N_7022,N_7596);
and U8023 (N_8023,N_7701,N_7733);
nor U8024 (N_8024,N_7472,N_7922);
nand U8025 (N_8025,N_7116,N_7195);
nor U8026 (N_8026,N_7282,N_7848);
nor U8027 (N_8027,N_7779,N_7388);
nand U8028 (N_8028,N_7546,N_7374);
xnor U8029 (N_8029,N_7839,N_7852);
nor U8030 (N_8030,N_7765,N_7269);
nor U8031 (N_8031,N_7057,N_7121);
nor U8032 (N_8032,N_7058,N_7265);
nand U8033 (N_8033,N_7530,N_7592);
or U8034 (N_8034,N_7547,N_7004);
nor U8035 (N_8035,N_7228,N_7371);
nor U8036 (N_8036,N_7956,N_7664);
nor U8037 (N_8037,N_7548,N_7935);
xor U8038 (N_8038,N_7226,N_7558);
and U8039 (N_8039,N_7213,N_7015);
and U8040 (N_8040,N_7660,N_7204);
xnor U8041 (N_8041,N_7986,N_7595);
or U8042 (N_8042,N_7353,N_7768);
or U8043 (N_8043,N_7869,N_7481);
and U8044 (N_8044,N_7785,N_7523);
nand U8045 (N_8045,N_7056,N_7403);
xnor U8046 (N_8046,N_7632,N_7657);
nand U8047 (N_8047,N_7377,N_7460);
nor U8048 (N_8048,N_7902,N_7987);
xor U8049 (N_8049,N_7506,N_7527);
and U8050 (N_8050,N_7362,N_7894);
nor U8051 (N_8051,N_7888,N_7997);
and U8052 (N_8052,N_7199,N_7617);
or U8053 (N_8053,N_7504,N_7147);
or U8054 (N_8054,N_7202,N_7402);
nand U8055 (N_8055,N_7691,N_7767);
nor U8056 (N_8056,N_7095,N_7300);
nand U8057 (N_8057,N_7003,N_7214);
nor U8058 (N_8058,N_7092,N_7396);
nor U8059 (N_8059,N_7811,N_7989);
xnor U8060 (N_8060,N_7410,N_7212);
xnor U8061 (N_8061,N_7191,N_7984);
and U8062 (N_8062,N_7821,N_7099);
nand U8063 (N_8063,N_7359,N_7755);
and U8064 (N_8064,N_7112,N_7052);
and U8065 (N_8065,N_7620,N_7045);
nor U8066 (N_8066,N_7316,N_7978);
or U8067 (N_8067,N_7338,N_7919);
and U8068 (N_8068,N_7610,N_7562);
nand U8069 (N_8069,N_7067,N_7738);
xnor U8070 (N_8070,N_7034,N_7794);
and U8071 (N_8071,N_7850,N_7746);
nand U8072 (N_8072,N_7231,N_7341);
xnor U8073 (N_8073,N_7583,N_7211);
nand U8074 (N_8074,N_7133,N_7429);
and U8075 (N_8075,N_7822,N_7440);
nor U8076 (N_8076,N_7135,N_7812);
xnor U8077 (N_8077,N_7859,N_7387);
xnor U8078 (N_8078,N_7705,N_7019);
and U8079 (N_8079,N_7758,N_7828);
xor U8080 (N_8080,N_7729,N_7892);
or U8081 (N_8081,N_7025,N_7790);
or U8082 (N_8082,N_7877,N_7509);
or U8083 (N_8083,N_7478,N_7216);
and U8084 (N_8084,N_7791,N_7062);
nor U8085 (N_8085,N_7853,N_7073);
nor U8086 (N_8086,N_7136,N_7115);
and U8087 (N_8087,N_7637,N_7661);
or U8088 (N_8088,N_7111,N_7678);
xnor U8089 (N_8089,N_7459,N_7898);
or U8090 (N_8090,N_7305,N_7087);
nand U8091 (N_8091,N_7273,N_7177);
and U8092 (N_8092,N_7905,N_7081);
and U8093 (N_8093,N_7965,N_7865);
xor U8094 (N_8094,N_7278,N_7958);
xor U8095 (N_8095,N_7421,N_7125);
nor U8096 (N_8096,N_7489,N_7614);
xor U8097 (N_8097,N_7172,N_7653);
or U8098 (N_8098,N_7659,N_7837);
xnor U8099 (N_8099,N_7722,N_7361);
xnor U8100 (N_8100,N_7581,N_7411);
nand U8101 (N_8101,N_7232,N_7078);
xor U8102 (N_8102,N_7076,N_7616);
and U8103 (N_8103,N_7517,N_7684);
nand U8104 (N_8104,N_7268,N_7151);
or U8105 (N_8105,N_7996,N_7071);
and U8106 (N_8106,N_7130,N_7090);
or U8107 (N_8107,N_7566,N_7166);
and U8108 (N_8108,N_7249,N_7760);
and U8109 (N_8109,N_7612,N_7658);
and U8110 (N_8110,N_7887,N_7759);
and U8111 (N_8111,N_7134,N_7082);
and U8112 (N_8112,N_7035,N_7027);
and U8113 (N_8113,N_7943,N_7161);
and U8114 (N_8114,N_7408,N_7505);
and U8115 (N_8115,N_7551,N_7868);
or U8116 (N_8116,N_7744,N_7171);
or U8117 (N_8117,N_7123,N_7590);
and U8118 (N_8118,N_7193,N_7330);
and U8119 (N_8119,N_7301,N_7126);
xnor U8120 (N_8120,N_7322,N_7069);
and U8121 (N_8121,N_7014,N_7054);
nor U8122 (N_8122,N_7732,N_7236);
nor U8123 (N_8123,N_7375,N_7923);
nor U8124 (N_8124,N_7252,N_7325);
and U8125 (N_8125,N_7257,N_7155);
nor U8126 (N_8126,N_7565,N_7425);
or U8127 (N_8127,N_7016,N_7702);
nor U8128 (N_8128,N_7063,N_7917);
nand U8129 (N_8129,N_7468,N_7441);
nand U8130 (N_8130,N_7493,N_7890);
nand U8131 (N_8131,N_7381,N_7855);
xnor U8132 (N_8132,N_7949,N_7320);
or U8133 (N_8133,N_7552,N_7836);
and U8134 (N_8134,N_7588,N_7689);
nand U8135 (N_8135,N_7480,N_7223);
and U8136 (N_8136,N_7060,N_7818);
or U8137 (N_8137,N_7178,N_7766);
or U8138 (N_8138,N_7247,N_7823);
nor U8139 (N_8139,N_7699,N_7947);
and U8140 (N_8140,N_7379,N_7229);
nand U8141 (N_8141,N_7927,N_7439);
xnor U8142 (N_8142,N_7961,N_7384);
or U8143 (N_8143,N_7576,N_7113);
nand U8144 (N_8144,N_7347,N_7187);
nand U8145 (N_8145,N_7146,N_7365);
or U8146 (N_8146,N_7307,N_7652);
and U8147 (N_8147,N_7860,N_7769);
or U8148 (N_8148,N_7311,N_7535);
and U8149 (N_8149,N_7011,N_7041);
and U8150 (N_8150,N_7655,N_7646);
or U8151 (N_8151,N_7777,N_7948);
and U8152 (N_8152,N_7462,N_7005);
and U8153 (N_8153,N_7143,N_7977);
nor U8154 (N_8154,N_7200,N_7197);
xor U8155 (N_8155,N_7773,N_7241);
and U8156 (N_8156,N_7453,N_7914);
and U8157 (N_8157,N_7020,N_7053);
nand U8158 (N_8158,N_7662,N_7033);
xnor U8159 (N_8159,N_7284,N_7974);
and U8160 (N_8160,N_7788,N_7635);
nand U8161 (N_8161,N_7569,N_7825);
nor U8162 (N_8162,N_7762,N_7544);
or U8163 (N_8163,N_7194,N_7712);
nor U8164 (N_8164,N_7999,N_7055);
nor U8165 (N_8165,N_7954,N_7532);
nor U8166 (N_8166,N_7931,N_7929);
nor U8167 (N_8167,N_7404,N_7382);
and U8168 (N_8168,N_7108,N_7918);
nand U8169 (N_8169,N_7477,N_7862);
nor U8170 (N_8170,N_7237,N_7405);
nand U8171 (N_8171,N_7272,N_7973);
nand U8172 (N_8172,N_7910,N_7626);
xor U8173 (N_8173,N_7484,N_7771);
xnor U8174 (N_8174,N_7531,N_7824);
or U8175 (N_8175,N_7219,N_7838);
nor U8176 (N_8176,N_7805,N_7520);
nand U8177 (N_8177,N_7577,N_7538);
xnor U8178 (N_8178,N_7797,N_7217);
xor U8179 (N_8179,N_7619,N_7242);
nor U8180 (N_8180,N_7623,N_7679);
xor U8181 (N_8181,N_7795,N_7461);
or U8182 (N_8182,N_7445,N_7735);
or U8183 (N_8183,N_7117,N_7802);
or U8184 (N_8184,N_7604,N_7843);
and U8185 (N_8185,N_7238,N_7700);
or U8186 (N_8186,N_7324,N_7438);
xor U8187 (N_8187,N_7145,N_7206);
nand U8188 (N_8188,N_7751,N_7499);
or U8189 (N_8189,N_7378,N_7329);
xor U8190 (N_8190,N_7666,N_7179);
and U8191 (N_8191,N_7141,N_7781);
or U8192 (N_8192,N_7876,N_7363);
or U8193 (N_8193,N_7064,N_7940);
or U8194 (N_8194,N_7186,N_7743);
xnor U8195 (N_8195,N_7774,N_7118);
nand U8196 (N_8196,N_7415,N_7456);
xnor U8197 (N_8197,N_7803,N_7398);
xnor U8198 (N_8198,N_7101,N_7793);
and U8199 (N_8199,N_7358,N_7075);
and U8200 (N_8200,N_7782,N_7938);
and U8201 (N_8201,N_7518,N_7649);
nor U8202 (N_8202,N_7114,N_7490);
nor U8203 (N_8203,N_7224,N_7611);
and U8204 (N_8204,N_7740,N_7454);
nor U8205 (N_8205,N_7783,N_7367);
and U8206 (N_8206,N_7512,N_7209);
or U8207 (N_8207,N_7185,N_7571);
nor U8208 (N_8208,N_7482,N_7920);
or U8209 (N_8209,N_7713,N_7264);
nand U8210 (N_8210,N_7068,N_7295);
nand U8211 (N_8211,N_7745,N_7776);
and U8212 (N_8212,N_7182,N_7763);
and U8213 (N_8213,N_7469,N_7846);
nor U8214 (N_8214,N_7475,N_7871);
and U8215 (N_8215,N_7503,N_7613);
nand U8216 (N_8216,N_7624,N_7521);
or U8217 (N_8217,N_7281,N_7435);
or U8218 (N_8218,N_7559,N_7266);
nor U8219 (N_8219,N_7110,N_7899);
or U8220 (N_8220,N_7663,N_7184);
nor U8221 (N_8221,N_7234,N_7519);
nor U8222 (N_8222,N_7640,N_7208);
nand U8223 (N_8223,N_7677,N_7934);
nor U8224 (N_8224,N_7010,N_7980);
nand U8225 (N_8225,N_7293,N_7796);
or U8226 (N_8226,N_7957,N_7951);
nand U8227 (N_8227,N_7921,N_7545);
and U8228 (N_8228,N_7176,N_7434);
xor U8229 (N_8229,N_7391,N_7636);
nand U8230 (N_8230,N_7644,N_7443);
xnor U8231 (N_8231,N_7697,N_7842);
xor U8232 (N_8232,N_7497,N_7753);
and U8233 (N_8233,N_7400,N_7979);
and U8234 (N_8234,N_7599,N_7908);
nor U8235 (N_8235,N_7085,N_7676);
nor U8236 (N_8236,N_7294,N_7152);
or U8237 (N_8237,N_7775,N_7080);
nand U8238 (N_8238,N_7856,N_7383);
xor U8239 (N_8239,N_7083,N_7798);
nor U8240 (N_8240,N_7685,N_7985);
and U8241 (N_8241,N_7983,N_7476);
or U8242 (N_8242,N_7972,N_7864);
and U8243 (N_8243,N_7031,N_7356);
and U8244 (N_8244,N_7895,N_7502);
nor U8245 (N_8245,N_7140,N_7522);
nand U8246 (N_8246,N_7752,N_7707);
xnor U8247 (N_8247,N_7982,N_7030);
nor U8248 (N_8248,N_7335,N_7444);
xor U8249 (N_8249,N_7501,N_7603);
or U8250 (N_8250,N_7556,N_7575);
xor U8251 (N_8251,N_7040,N_7343);
and U8252 (N_8252,N_7719,N_7274);
nand U8253 (N_8253,N_7107,N_7368);
or U8254 (N_8254,N_7627,N_7584);
and U8255 (N_8255,N_7065,N_7225);
nor U8256 (N_8256,N_7715,N_7933);
xor U8257 (N_8257,N_7156,N_7296);
or U8258 (N_8258,N_7749,N_7723);
nor U8259 (N_8259,N_7543,N_7392);
and U8260 (N_8260,N_7006,N_7098);
xor U8261 (N_8261,N_7017,N_7542);
nand U8262 (N_8262,N_7704,N_7994);
and U8263 (N_8263,N_7650,N_7059);
nand U8264 (N_8264,N_7180,N_7406);
xnor U8265 (N_8265,N_7734,N_7420);
nand U8266 (N_8266,N_7448,N_7739);
nand U8267 (N_8267,N_7834,N_7881);
and U8268 (N_8268,N_7670,N_7630);
nand U8269 (N_8269,N_7433,N_7345);
nand U8270 (N_8270,N_7750,N_7880);
or U8271 (N_8271,N_7409,N_7157);
nor U8272 (N_8272,N_7473,N_7800);
nand U8273 (N_8273,N_7297,N_7449);
nand U8274 (N_8274,N_7539,N_7928);
nor U8275 (N_8275,N_7939,N_7164);
and U8276 (N_8276,N_7742,N_7037);
nor U8277 (N_8277,N_7789,N_7196);
nand U8278 (N_8278,N_7276,N_7074);
nand U8279 (N_8279,N_7446,N_7875);
and U8280 (N_8280,N_7084,N_7605);
or U8281 (N_8281,N_7256,N_7622);
nor U8282 (N_8282,N_7572,N_7807);
xnor U8283 (N_8283,N_7683,N_7799);
xnor U8284 (N_8284,N_7525,N_7465);
xnor U8285 (N_8285,N_7631,N_7245);
and U8286 (N_8286,N_7203,N_7183);
xnor U8287 (N_8287,N_7866,N_7587);
and U8288 (N_8288,N_7221,N_7680);
and U8289 (N_8289,N_7317,N_7220);
or U8290 (N_8290,N_7896,N_7510);
or U8291 (N_8291,N_7645,N_7351);
nor U8292 (N_8292,N_7528,N_7873);
and U8293 (N_8293,N_7168,N_7306);
and U8294 (N_8294,N_7971,N_7309);
or U8295 (N_8295,N_7814,N_7968);
nand U8296 (N_8296,N_7629,N_7390);
nand U8297 (N_8297,N_7819,N_7500);
and U8298 (N_8298,N_7903,N_7861);
nand U8299 (N_8299,N_7808,N_7711);
xor U8300 (N_8300,N_7780,N_7131);
nand U8301 (N_8301,N_7354,N_7801);
nor U8302 (N_8302,N_7120,N_7048);
nor U8303 (N_8303,N_7360,N_7741);
nor U8304 (N_8304,N_7319,N_7654);
or U8305 (N_8305,N_7254,N_7737);
nand U8306 (N_8306,N_7827,N_7149);
nor U8307 (N_8307,N_7792,N_7553);
nand U8308 (N_8308,N_7430,N_7893);
xor U8309 (N_8309,N_7416,N_7215);
nor U8310 (N_8310,N_7298,N_7244);
or U8311 (N_8311,N_7561,N_7778);
or U8312 (N_8312,N_7915,N_7962);
xnor U8313 (N_8313,N_7452,N_7032);
or U8314 (N_8314,N_7942,N_7847);
and U8315 (N_8315,N_7537,N_7447);
and U8316 (N_8316,N_7727,N_7255);
and U8317 (N_8317,N_7376,N_7686);
or U8318 (N_8318,N_7508,N_7946);
and U8319 (N_8319,N_7450,N_7813);
nor U8320 (N_8320,N_7582,N_7573);
or U8321 (N_8321,N_7026,N_7227);
and U8322 (N_8322,N_7872,N_7162);
xnor U8323 (N_8323,N_7882,N_7633);
xor U8324 (N_8324,N_7089,N_7607);
nor U8325 (N_8325,N_7285,N_7279);
and U8326 (N_8326,N_7784,N_7886);
or U8327 (N_8327,N_7851,N_7606);
nand U8328 (N_8328,N_7050,N_7369);
and U8329 (N_8329,N_7594,N_7253);
or U8330 (N_8330,N_7129,N_7529);
nand U8331 (N_8331,N_7471,N_7457);
nand U8332 (N_8332,N_7580,N_7039);
and U8333 (N_8333,N_7695,N_7431);
xnor U8334 (N_8334,N_7170,N_7831);
nand U8335 (N_8335,N_7786,N_7419);
xnor U8336 (N_8336,N_7534,N_7109);
and U8337 (N_8337,N_7844,N_7275);
xnor U8338 (N_8338,N_7878,N_7668);
nand U8339 (N_8339,N_7731,N_7857);
nand U8340 (N_8340,N_7366,N_7397);
nor U8341 (N_8341,N_7648,N_7401);
nand U8342 (N_8342,N_7380,N_7013);
xor U8343 (N_8343,N_7900,N_7474);
nand U8344 (N_8344,N_7698,N_7845);
and U8345 (N_8345,N_7976,N_7100);
xnor U8346 (N_8346,N_7029,N_7190);
xor U8347 (N_8347,N_7944,N_7491);
or U8348 (N_8348,N_7153,N_7990);
xnor U8349 (N_8349,N_7672,N_7163);
nand U8350 (N_8350,N_7674,N_7656);
nand U8351 (N_8351,N_7086,N_7849);
xnor U8352 (N_8352,N_7270,N_7969);
xor U8353 (N_8353,N_7286,N_7097);
and U8354 (N_8354,N_7250,N_7725);
xor U8355 (N_8355,N_7486,N_7077);
xor U8356 (N_8356,N_7139,N_7515);
nand U8357 (N_8357,N_7174,N_7321);
or U8358 (N_8358,N_7967,N_7618);
or U8359 (N_8359,N_7925,N_7966);
nand U8360 (N_8360,N_7159,N_7291);
nand U8361 (N_8361,N_7315,N_7806);
or U8362 (N_8362,N_7012,N_7327);
and U8363 (N_8363,N_7889,N_7709);
and U8364 (N_8364,N_7042,N_7567);
nand U8365 (N_8365,N_7413,N_7717);
nor U8366 (N_8366,N_7198,N_7804);
and U8367 (N_8367,N_7564,N_7008);
xor U8368 (N_8368,N_7550,N_7395);
and U8369 (N_8369,N_7385,N_7260);
nand U8370 (N_8370,N_7830,N_7201);
and U8371 (N_8371,N_7991,N_7826);
or U8372 (N_8372,N_7370,N_7568);
xor U8373 (N_8373,N_7043,N_7833);
or U8374 (N_8374,N_7458,N_7549);
xnor U8375 (N_8375,N_7348,N_7835);
xor U8376 (N_8376,N_7287,N_7858);
xor U8377 (N_8377,N_7554,N_7102);
and U8378 (N_8378,N_7589,N_7621);
xor U8379 (N_8379,N_7907,N_7952);
xnor U8380 (N_8380,N_7716,N_7820);
or U8381 (N_8381,N_7601,N_7258);
or U8382 (N_8382,N_7336,N_7093);
xor U8383 (N_8383,N_7516,N_7682);
nor U8384 (N_8384,N_7579,N_7280);
or U8385 (N_8385,N_7277,N_7574);
or U8386 (N_8386,N_7945,N_7941);
nand U8387 (N_8387,N_7710,N_7148);
nor U8388 (N_8388,N_7451,N_7426);
and U8389 (N_8389,N_7960,N_7639);
nor U8390 (N_8390,N_7496,N_7593);
nand U8391 (N_8391,N_7038,N_7912);
nor U8392 (N_8392,N_7891,N_7181);
nor U8393 (N_8393,N_7119,N_7787);
xnor U8394 (N_8394,N_7165,N_7955);
and U8395 (N_8395,N_7160,N_7748);
nand U8396 (N_8396,N_7044,N_7690);
or U8397 (N_8397,N_7494,N_7096);
nand U8398 (N_8398,N_7829,N_7331);
and U8399 (N_8399,N_7205,N_7364);
nand U8400 (N_8400,N_7688,N_7671);
and U8401 (N_8401,N_7418,N_7757);
nand U8402 (N_8402,N_7313,N_7854);
nand U8403 (N_8403,N_7863,N_7665);
nand U8404 (N_8404,N_7916,N_7021);
and U8405 (N_8405,N_7009,N_7597);
and U8406 (N_8406,N_7332,N_7832);
or U8407 (N_8407,N_7483,N_7870);
or U8408 (N_8408,N_7207,N_7417);
nor U8409 (N_8409,N_7414,N_7724);
and U8410 (N_8410,N_7728,N_7467);
or U8411 (N_8411,N_7289,N_7687);
xnor U8412 (N_8412,N_7911,N_7072);
or U8413 (N_8413,N_7154,N_7372);
nor U8414 (N_8414,N_7647,N_7105);
and U8415 (N_8415,N_7188,N_7079);
and U8416 (N_8416,N_7326,N_7770);
or U8417 (N_8417,N_7602,N_7259);
xor U8418 (N_8418,N_7142,N_7328);
nor U8419 (N_8419,N_7578,N_7930);
nor U8420 (N_8420,N_7304,N_7675);
or U8421 (N_8421,N_7036,N_7708);
and U8422 (N_8422,N_7498,N_7959);
nor U8423 (N_8423,N_7964,N_7924);
nand U8424 (N_8424,N_7094,N_7233);
and U8425 (N_8425,N_7103,N_7586);
xnor U8426 (N_8426,N_7761,N_7669);
and U8427 (N_8427,N_7189,N_7560);
xnor U8428 (N_8428,N_7422,N_7437);
and U8429 (N_8429,N_7106,N_7681);
xor U8430 (N_8430,N_7692,N_7507);
xnor U8431 (N_8431,N_7218,N_7495);
or U8432 (N_8432,N_7703,N_7563);
and U8433 (N_8433,N_7432,N_7302);
and U8434 (N_8434,N_7714,N_7066);
nand U8435 (N_8435,N_7513,N_7314);
or U8436 (N_8436,N_7600,N_7841);
xnor U8437 (N_8437,N_7399,N_7696);
and U8438 (N_8438,N_7323,N_7993);
xor U8439 (N_8439,N_7334,N_7455);
xnor U8440 (N_8440,N_7167,N_7673);
nor U8441 (N_8441,N_7464,N_7246);
or U8442 (N_8442,N_7339,N_7222);
nor U8443 (N_8443,N_7061,N_7344);
or U8444 (N_8444,N_7070,N_7570);
xnor U8445 (N_8445,N_7526,N_7355);
or U8446 (N_8446,N_7436,N_7511);
nand U8447 (N_8447,N_7815,N_7651);
nand U8448 (N_8448,N_7754,N_7144);
or U8449 (N_8449,N_7897,N_7290);
nand U8450 (N_8450,N_7747,N_7137);
nor U8451 (N_8451,N_7904,N_7634);
nand U8452 (N_8452,N_7352,N_7913);
nor U8453 (N_8453,N_7463,N_7018);
and U8454 (N_8454,N_7357,N_7240);
or U8455 (N_8455,N_7540,N_7303);
and U8456 (N_8456,N_7427,N_7251);
and U8457 (N_8457,N_7487,N_7840);
and U8458 (N_8458,N_7694,N_7693);
or U8459 (N_8459,N_7541,N_7642);
nor U8460 (N_8460,N_7350,N_7127);
nand U8461 (N_8461,N_7643,N_7318);
nand U8462 (N_8462,N_7428,N_7412);
and U8463 (N_8463,N_7023,N_7342);
nand U8464 (N_8464,N_7970,N_7591);
and U8465 (N_8465,N_7000,N_7091);
or U8466 (N_8466,N_7104,N_7299);
and U8467 (N_8467,N_7001,N_7901);
and U8468 (N_8468,N_7346,N_7340);
and U8469 (N_8469,N_7243,N_7210);
xor U8470 (N_8470,N_7874,N_7817);
nand U8471 (N_8471,N_7235,N_7533);
xnor U8472 (N_8472,N_7585,N_7288);
nor U8473 (N_8473,N_7726,N_7628);
xnor U8474 (N_8474,N_7992,N_7470);
and U8475 (N_8475,N_7706,N_7936);
or U8476 (N_8476,N_7122,N_7263);
and U8477 (N_8477,N_7047,N_7730);
nand U8478 (N_8478,N_7884,N_7615);
and U8479 (N_8479,N_7028,N_7950);
nand U8480 (N_8480,N_7386,N_7173);
nor U8481 (N_8481,N_7308,N_7046);
and U8482 (N_8482,N_7885,N_7756);
nand U8483 (N_8483,N_7810,N_7555);
nand U8484 (N_8484,N_7271,N_7310);
nand U8485 (N_8485,N_7423,N_7816);
or U8486 (N_8486,N_7995,N_7492);
or U8487 (N_8487,N_7608,N_7333);
nand U8488 (N_8488,N_7267,N_7424);
or U8489 (N_8489,N_7720,N_7373);
nor U8490 (N_8490,N_7442,N_7088);
and U8491 (N_8491,N_7736,N_7867);
xor U8492 (N_8492,N_7239,N_7150);
nor U8493 (N_8493,N_7514,N_7932);
xnor U8494 (N_8494,N_7007,N_7169);
xor U8495 (N_8495,N_7764,N_7718);
xnor U8496 (N_8496,N_7598,N_7524);
xor U8497 (N_8497,N_7051,N_7248);
and U8498 (N_8498,N_7158,N_7772);
or U8499 (N_8499,N_7479,N_7132);
and U8500 (N_8500,N_7037,N_7270);
or U8501 (N_8501,N_7817,N_7735);
nand U8502 (N_8502,N_7027,N_7123);
or U8503 (N_8503,N_7369,N_7883);
nand U8504 (N_8504,N_7009,N_7722);
nand U8505 (N_8505,N_7369,N_7176);
and U8506 (N_8506,N_7038,N_7885);
nand U8507 (N_8507,N_7040,N_7151);
nor U8508 (N_8508,N_7909,N_7439);
and U8509 (N_8509,N_7844,N_7544);
nand U8510 (N_8510,N_7612,N_7569);
and U8511 (N_8511,N_7434,N_7534);
xor U8512 (N_8512,N_7552,N_7062);
xnor U8513 (N_8513,N_7139,N_7560);
or U8514 (N_8514,N_7073,N_7571);
or U8515 (N_8515,N_7940,N_7208);
and U8516 (N_8516,N_7542,N_7939);
or U8517 (N_8517,N_7388,N_7325);
nand U8518 (N_8518,N_7681,N_7945);
nor U8519 (N_8519,N_7224,N_7862);
or U8520 (N_8520,N_7971,N_7623);
nand U8521 (N_8521,N_7202,N_7631);
xnor U8522 (N_8522,N_7401,N_7755);
or U8523 (N_8523,N_7804,N_7377);
nand U8524 (N_8524,N_7970,N_7363);
nand U8525 (N_8525,N_7398,N_7922);
nor U8526 (N_8526,N_7631,N_7139);
and U8527 (N_8527,N_7708,N_7234);
nor U8528 (N_8528,N_7525,N_7841);
nor U8529 (N_8529,N_7750,N_7396);
xnor U8530 (N_8530,N_7829,N_7800);
and U8531 (N_8531,N_7022,N_7475);
and U8532 (N_8532,N_7216,N_7148);
or U8533 (N_8533,N_7609,N_7409);
xnor U8534 (N_8534,N_7337,N_7764);
xor U8535 (N_8535,N_7920,N_7969);
nor U8536 (N_8536,N_7473,N_7197);
xnor U8537 (N_8537,N_7570,N_7834);
or U8538 (N_8538,N_7120,N_7211);
or U8539 (N_8539,N_7748,N_7369);
or U8540 (N_8540,N_7065,N_7670);
xnor U8541 (N_8541,N_7038,N_7922);
nor U8542 (N_8542,N_7288,N_7418);
or U8543 (N_8543,N_7509,N_7005);
nor U8544 (N_8544,N_7147,N_7317);
xor U8545 (N_8545,N_7058,N_7116);
and U8546 (N_8546,N_7981,N_7837);
or U8547 (N_8547,N_7866,N_7493);
or U8548 (N_8548,N_7370,N_7463);
or U8549 (N_8549,N_7195,N_7723);
xnor U8550 (N_8550,N_7610,N_7725);
nor U8551 (N_8551,N_7611,N_7997);
xor U8552 (N_8552,N_7386,N_7438);
and U8553 (N_8553,N_7213,N_7059);
nand U8554 (N_8554,N_7220,N_7623);
or U8555 (N_8555,N_7657,N_7644);
or U8556 (N_8556,N_7638,N_7760);
nor U8557 (N_8557,N_7845,N_7984);
xor U8558 (N_8558,N_7855,N_7436);
or U8559 (N_8559,N_7203,N_7005);
xor U8560 (N_8560,N_7387,N_7183);
xnor U8561 (N_8561,N_7935,N_7347);
nand U8562 (N_8562,N_7326,N_7020);
or U8563 (N_8563,N_7684,N_7259);
nand U8564 (N_8564,N_7638,N_7291);
xnor U8565 (N_8565,N_7413,N_7830);
or U8566 (N_8566,N_7213,N_7014);
nor U8567 (N_8567,N_7313,N_7192);
xor U8568 (N_8568,N_7026,N_7608);
xor U8569 (N_8569,N_7438,N_7757);
and U8570 (N_8570,N_7177,N_7631);
nand U8571 (N_8571,N_7014,N_7565);
xnor U8572 (N_8572,N_7621,N_7882);
xor U8573 (N_8573,N_7771,N_7187);
nor U8574 (N_8574,N_7656,N_7526);
xor U8575 (N_8575,N_7979,N_7507);
xor U8576 (N_8576,N_7248,N_7158);
and U8577 (N_8577,N_7528,N_7583);
nand U8578 (N_8578,N_7655,N_7313);
nor U8579 (N_8579,N_7783,N_7791);
xor U8580 (N_8580,N_7040,N_7016);
or U8581 (N_8581,N_7595,N_7025);
xor U8582 (N_8582,N_7761,N_7642);
nand U8583 (N_8583,N_7348,N_7639);
or U8584 (N_8584,N_7315,N_7292);
nand U8585 (N_8585,N_7813,N_7752);
nor U8586 (N_8586,N_7151,N_7781);
xor U8587 (N_8587,N_7348,N_7957);
xor U8588 (N_8588,N_7666,N_7410);
and U8589 (N_8589,N_7128,N_7805);
and U8590 (N_8590,N_7225,N_7169);
nand U8591 (N_8591,N_7910,N_7977);
or U8592 (N_8592,N_7513,N_7761);
or U8593 (N_8593,N_7736,N_7700);
or U8594 (N_8594,N_7399,N_7096);
or U8595 (N_8595,N_7476,N_7242);
and U8596 (N_8596,N_7207,N_7078);
and U8597 (N_8597,N_7422,N_7967);
nor U8598 (N_8598,N_7307,N_7299);
nand U8599 (N_8599,N_7246,N_7620);
nand U8600 (N_8600,N_7847,N_7800);
nor U8601 (N_8601,N_7733,N_7184);
xor U8602 (N_8602,N_7697,N_7542);
or U8603 (N_8603,N_7018,N_7336);
nor U8604 (N_8604,N_7693,N_7596);
nor U8605 (N_8605,N_7249,N_7360);
nor U8606 (N_8606,N_7238,N_7086);
nand U8607 (N_8607,N_7435,N_7255);
and U8608 (N_8608,N_7796,N_7626);
nor U8609 (N_8609,N_7835,N_7813);
xnor U8610 (N_8610,N_7273,N_7609);
and U8611 (N_8611,N_7774,N_7473);
xor U8612 (N_8612,N_7840,N_7971);
nand U8613 (N_8613,N_7296,N_7165);
nand U8614 (N_8614,N_7589,N_7369);
xnor U8615 (N_8615,N_7405,N_7794);
nand U8616 (N_8616,N_7411,N_7371);
nor U8617 (N_8617,N_7992,N_7245);
xnor U8618 (N_8618,N_7671,N_7718);
nor U8619 (N_8619,N_7128,N_7550);
or U8620 (N_8620,N_7758,N_7867);
nor U8621 (N_8621,N_7386,N_7572);
xor U8622 (N_8622,N_7209,N_7780);
and U8623 (N_8623,N_7413,N_7028);
or U8624 (N_8624,N_7142,N_7593);
nor U8625 (N_8625,N_7834,N_7827);
nand U8626 (N_8626,N_7365,N_7566);
nand U8627 (N_8627,N_7928,N_7900);
nor U8628 (N_8628,N_7110,N_7526);
xor U8629 (N_8629,N_7953,N_7824);
or U8630 (N_8630,N_7532,N_7956);
and U8631 (N_8631,N_7645,N_7690);
or U8632 (N_8632,N_7718,N_7090);
and U8633 (N_8633,N_7289,N_7405);
and U8634 (N_8634,N_7201,N_7707);
nor U8635 (N_8635,N_7334,N_7742);
nand U8636 (N_8636,N_7325,N_7155);
nand U8637 (N_8637,N_7521,N_7142);
nand U8638 (N_8638,N_7189,N_7329);
nand U8639 (N_8639,N_7477,N_7041);
nand U8640 (N_8640,N_7087,N_7977);
xor U8641 (N_8641,N_7456,N_7136);
or U8642 (N_8642,N_7204,N_7929);
or U8643 (N_8643,N_7264,N_7881);
nand U8644 (N_8644,N_7190,N_7711);
and U8645 (N_8645,N_7118,N_7795);
nor U8646 (N_8646,N_7617,N_7765);
or U8647 (N_8647,N_7692,N_7537);
or U8648 (N_8648,N_7599,N_7697);
and U8649 (N_8649,N_7222,N_7697);
or U8650 (N_8650,N_7335,N_7783);
and U8651 (N_8651,N_7986,N_7427);
nor U8652 (N_8652,N_7008,N_7134);
nand U8653 (N_8653,N_7804,N_7313);
and U8654 (N_8654,N_7130,N_7901);
or U8655 (N_8655,N_7146,N_7832);
nand U8656 (N_8656,N_7609,N_7564);
and U8657 (N_8657,N_7661,N_7021);
nand U8658 (N_8658,N_7223,N_7436);
nand U8659 (N_8659,N_7609,N_7475);
and U8660 (N_8660,N_7923,N_7381);
nor U8661 (N_8661,N_7939,N_7351);
xnor U8662 (N_8662,N_7113,N_7120);
nand U8663 (N_8663,N_7268,N_7260);
xor U8664 (N_8664,N_7985,N_7687);
and U8665 (N_8665,N_7792,N_7222);
nand U8666 (N_8666,N_7324,N_7861);
nand U8667 (N_8667,N_7795,N_7191);
xor U8668 (N_8668,N_7616,N_7688);
nand U8669 (N_8669,N_7152,N_7037);
nand U8670 (N_8670,N_7666,N_7929);
nor U8671 (N_8671,N_7282,N_7131);
xnor U8672 (N_8672,N_7284,N_7511);
nor U8673 (N_8673,N_7354,N_7827);
nor U8674 (N_8674,N_7693,N_7717);
nand U8675 (N_8675,N_7777,N_7314);
xnor U8676 (N_8676,N_7489,N_7162);
and U8677 (N_8677,N_7815,N_7267);
nand U8678 (N_8678,N_7413,N_7796);
xnor U8679 (N_8679,N_7700,N_7220);
nor U8680 (N_8680,N_7380,N_7228);
and U8681 (N_8681,N_7690,N_7593);
nand U8682 (N_8682,N_7149,N_7094);
xnor U8683 (N_8683,N_7079,N_7944);
and U8684 (N_8684,N_7956,N_7540);
xnor U8685 (N_8685,N_7965,N_7580);
or U8686 (N_8686,N_7761,N_7073);
and U8687 (N_8687,N_7255,N_7750);
xnor U8688 (N_8688,N_7447,N_7523);
xnor U8689 (N_8689,N_7529,N_7814);
or U8690 (N_8690,N_7156,N_7510);
or U8691 (N_8691,N_7808,N_7854);
or U8692 (N_8692,N_7326,N_7336);
nand U8693 (N_8693,N_7657,N_7145);
nand U8694 (N_8694,N_7453,N_7696);
or U8695 (N_8695,N_7107,N_7287);
nand U8696 (N_8696,N_7943,N_7472);
xor U8697 (N_8697,N_7429,N_7857);
xor U8698 (N_8698,N_7088,N_7322);
nor U8699 (N_8699,N_7025,N_7648);
xor U8700 (N_8700,N_7502,N_7536);
and U8701 (N_8701,N_7252,N_7159);
or U8702 (N_8702,N_7717,N_7924);
or U8703 (N_8703,N_7089,N_7191);
xnor U8704 (N_8704,N_7237,N_7888);
nor U8705 (N_8705,N_7919,N_7191);
nand U8706 (N_8706,N_7836,N_7411);
nand U8707 (N_8707,N_7460,N_7269);
and U8708 (N_8708,N_7903,N_7553);
or U8709 (N_8709,N_7768,N_7506);
or U8710 (N_8710,N_7220,N_7505);
nand U8711 (N_8711,N_7056,N_7999);
and U8712 (N_8712,N_7947,N_7983);
xnor U8713 (N_8713,N_7200,N_7178);
xor U8714 (N_8714,N_7329,N_7451);
and U8715 (N_8715,N_7402,N_7239);
and U8716 (N_8716,N_7598,N_7789);
xor U8717 (N_8717,N_7510,N_7534);
nor U8718 (N_8718,N_7898,N_7732);
nand U8719 (N_8719,N_7267,N_7087);
xor U8720 (N_8720,N_7297,N_7739);
or U8721 (N_8721,N_7210,N_7781);
and U8722 (N_8722,N_7033,N_7642);
nand U8723 (N_8723,N_7581,N_7526);
and U8724 (N_8724,N_7574,N_7890);
nand U8725 (N_8725,N_7143,N_7387);
xnor U8726 (N_8726,N_7242,N_7841);
or U8727 (N_8727,N_7463,N_7540);
or U8728 (N_8728,N_7642,N_7105);
and U8729 (N_8729,N_7731,N_7359);
or U8730 (N_8730,N_7162,N_7039);
or U8731 (N_8731,N_7012,N_7692);
nand U8732 (N_8732,N_7239,N_7816);
xnor U8733 (N_8733,N_7811,N_7346);
nand U8734 (N_8734,N_7907,N_7214);
nor U8735 (N_8735,N_7159,N_7166);
xor U8736 (N_8736,N_7893,N_7524);
nor U8737 (N_8737,N_7019,N_7938);
nor U8738 (N_8738,N_7431,N_7269);
xnor U8739 (N_8739,N_7630,N_7227);
or U8740 (N_8740,N_7538,N_7961);
and U8741 (N_8741,N_7151,N_7471);
and U8742 (N_8742,N_7140,N_7643);
nand U8743 (N_8743,N_7983,N_7912);
xor U8744 (N_8744,N_7023,N_7629);
nor U8745 (N_8745,N_7803,N_7668);
and U8746 (N_8746,N_7487,N_7452);
or U8747 (N_8747,N_7275,N_7494);
or U8748 (N_8748,N_7168,N_7823);
nor U8749 (N_8749,N_7355,N_7725);
xnor U8750 (N_8750,N_7324,N_7388);
nor U8751 (N_8751,N_7018,N_7626);
and U8752 (N_8752,N_7600,N_7073);
nand U8753 (N_8753,N_7453,N_7350);
xor U8754 (N_8754,N_7091,N_7794);
or U8755 (N_8755,N_7698,N_7713);
xnor U8756 (N_8756,N_7080,N_7151);
or U8757 (N_8757,N_7447,N_7592);
xnor U8758 (N_8758,N_7932,N_7448);
nor U8759 (N_8759,N_7199,N_7870);
and U8760 (N_8760,N_7845,N_7932);
nand U8761 (N_8761,N_7873,N_7278);
or U8762 (N_8762,N_7019,N_7338);
xnor U8763 (N_8763,N_7320,N_7345);
nor U8764 (N_8764,N_7009,N_7905);
and U8765 (N_8765,N_7245,N_7879);
nand U8766 (N_8766,N_7396,N_7887);
and U8767 (N_8767,N_7088,N_7410);
and U8768 (N_8768,N_7113,N_7774);
nand U8769 (N_8769,N_7943,N_7738);
xor U8770 (N_8770,N_7041,N_7868);
xor U8771 (N_8771,N_7009,N_7222);
nor U8772 (N_8772,N_7426,N_7840);
or U8773 (N_8773,N_7899,N_7314);
nand U8774 (N_8774,N_7856,N_7127);
nor U8775 (N_8775,N_7189,N_7059);
and U8776 (N_8776,N_7274,N_7257);
or U8777 (N_8777,N_7012,N_7245);
or U8778 (N_8778,N_7254,N_7128);
xnor U8779 (N_8779,N_7536,N_7632);
xnor U8780 (N_8780,N_7004,N_7828);
or U8781 (N_8781,N_7288,N_7666);
nor U8782 (N_8782,N_7305,N_7601);
and U8783 (N_8783,N_7935,N_7940);
nand U8784 (N_8784,N_7341,N_7979);
nand U8785 (N_8785,N_7649,N_7041);
or U8786 (N_8786,N_7497,N_7819);
and U8787 (N_8787,N_7402,N_7358);
xor U8788 (N_8788,N_7900,N_7735);
nand U8789 (N_8789,N_7715,N_7559);
nand U8790 (N_8790,N_7854,N_7517);
nor U8791 (N_8791,N_7821,N_7073);
nor U8792 (N_8792,N_7148,N_7726);
nor U8793 (N_8793,N_7994,N_7566);
xor U8794 (N_8794,N_7696,N_7592);
xnor U8795 (N_8795,N_7064,N_7133);
xnor U8796 (N_8796,N_7664,N_7802);
nor U8797 (N_8797,N_7173,N_7424);
xnor U8798 (N_8798,N_7222,N_7466);
or U8799 (N_8799,N_7471,N_7955);
nor U8800 (N_8800,N_7779,N_7351);
nor U8801 (N_8801,N_7885,N_7726);
nor U8802 (N_8802,N_7394,N_7764);
nor U8803 (N_8803,N_7921,N_7468);
nor U8804 (N_8804,N_7289,N_7379);
and U8805 (N_8805,N_7319,N_7415);
or U8806 (N_8806,N_7357,N_7189);
nand U8807 (N_8807,N_7043,N_7858);
or U8808 (N_8808,N_7480,N_7891);
nor U8809 (N_8809,N_7253,N_7911);
nand U8810 (N_8810,N_7223,N_7394);
or U8811 (N_8811,N_7413,N_7112);
xnor U8812 (N_8812,N_7509,N_7487);
nand U8813 (N_8813,N_7940,N_7480);
or U8814 (N_8814,N_7554,N_7806);
or U8815 (N_8815,N_7245,N_7047);
or U8816 (N_8816,N_7403,N_7199);
or U8817 (N_8817,N_7126,N_7974);
nand U8818 (N_8818,N_7028,N_7498);
nand U8819 (N_8819,N_7007,N_7065);
nor U8820 (N_8820,N_7069,N_7221);
and U8821 (N_8821,N_7273,N_7400);
and U8822 (N_8822,N_7887,N_7330);
nor U8823 (N_8823,N_7502,N_7355);
and U8824 (N_8824,N_7474,N_7178);
and U8825 (N_8825,N_7452,N_7081);
xor U8826 (N_8826,N_7504,N_7387);
nor U8827 (N_8827,N_7740,N_7731);
or U8828 (N_8828,N_7434,N_7319);
xor U8829 (N_8829,N_7026,N_7535);
xor U8830 (N_8830,N_7019,N_7656);
nand U8831 (N_8831,N_7654,N_7253);
nand U8832 (N_8832,N_7613,N_7241);
or U8833 (N_8833,N_7928,N_7706);
nor U8834 (N_8834,N_7888,N_7803);
nor U8835 (N_8835,N_7907,N_7364);
nor U8836 (N_8836,N_7479,N_7266);
and U8837 (N_8837,N_7910,N_7922);
nor U8838 (N_8838,N_7835,N_7830);
nand U8839 (N_8839,N_7758,N_7458);
nor U8840 (N_8840,N_7122,N_7633);
or U8841 (N_8841,N_7363,N_7250);
or U8842 (N_8842,N_7781,N_7737);
xor U8843 (N_8843,N_7966,N_7315);
nand U8844 (N_8844,N_7927,N_7171);
or U8845 (N_8845,N_7767,N_7491);
xor U8846 (N_8846,N_7068,N_7512);
xor U8847 (N_8847,N_7864,N_7478);
or U8848 (N_8848,N_7328,N_7258);
xor U8849 (N_8849,N_7601,N_7443);
or U8850 (N_8850,N_7295,N_7528);
and U8851 (N_8851,N_7777,N_7507);
nor U8852 (N_8852,N_7348,N_7010);
xnor U8853 (N_8853,N_7708,N_7427);
and U8854 (N_8854,N_7889,N_7145);
and U8855 (N_8855,N_7605,N_7826);
xor U8856 (N_8856,N_7945,N_7162);
nor U8857 (N_8857,N_7178,N_7641);
nor U8858 (N_8858,N_7366,N_7513);
and U8859 (N_8859,N_7129,N_7415);
xor U8860 (N_8860,N_7892,N_7795);
nand U8861 (N_8861,N_7846,N_7603);
xor U8862 (N_8862,N_7814,N_7023);
xor U8863 (N_8863,N_7423,N_7546);
xnor U8864 (N_8864,N_7795,N_7862);
and U8865 (N_8865,N_7052,N_7823);
nand U8866 (N_8866,N_7001,N_7080);
xnor U8867 (N_8867,N_7023,N_7325);
nand U8868 (N_8868,N_7879,N_7538);
xor U8869 (N_8869,N_7058,N_7144);
and U8870 (N_8870,N_7560,N_7041);
nor U8871 (N_8871,N_7379,N_7718);
xnor U8872 (N_8872,N_7634,N_7579);
nand U8873 (N_8873,N_7859,N_7696);
nand U8874 (N_8874,N_7448,N_7557);
xor U8875 (N_8875,N_7666,N_7561);
xnor U8876 (N_8876,N_7090,N_7756);
and U8877 (N_8877,N_7722,N_7218);
nor U8878 (N_8878,N_7387,N_7501);
or U8879 (N_8879,N_7043,N_7072);
nand U8880 (N_8880,N_7166,N_7132);
and U8881 (N_8881,N_7589,N_7902);
xnor U8882 (N_8882,N_7187,N_7020);
or U8883 (N_8883,N_7283,N_7108);
or U8884 (N_8884,N_7840,N_7281);
xnor U8885 (N_8885,N_7089,N_7982);
or U8886 (N_8886,N_7010,N_7166);
nand U8887 (N_8887,N_7454,N_7603);
nor U8888 (N_8888,N_7063,N_7218);
nor U8889 (N_8889,N_7297,N_7709);
nor U8890 (N_8890,N_7563,N_7079);
nand U8891 (N_8891,N_7897,N_7050);
xnor U8892 (N_8892,N_7737,N_7120);
or U8893 (N_8893,N_7304,N_7526);
or U8894 (N_8894,N_7952,N_7841);
nand U8895 (N_8895,N_7485,N_7030);
nand U8896 (N_8896,N_7661,N_7857);
xnor U8897 (N_8897,N_7035,N_7587);
and U8898 (N_8898,N_7736,N_7144);
and U8899 (N_8899,N_7760,N_7652);
and U8900 (N_8900,N_7949,N_7939);
or U8901 (N_8901,N_7779,N_7092);
nand U8902 (N_8902,N_7839,N_7906);
nor U8903 (N_8903,N_7170,N_7112);
xor U8904 (N_8904,N_7952,N_7775);
nand U8905 (N_8905,N_7361,N_7633);
nor U8906 (N_8906,N_7980,N_7473);
or U8907 (N_8907,N_7469,N_7980);
or U8908 (N_8908,N_7053,N_7925);
nor U8909 (N_8909,N_7070,N_7265);
or U8910 (N_8910,N_7765,N_7177);
nand U8911 (N_8911,N_7107,N_7778);
nand U8912 (N_8912,N_7452,N_7928);
or U8913 (N_8913,N_7916,N_7608);
nor U8914 (N_8914,N_7262,N_7529);
nor U8915 (N_8915,N_7686,N_7156);
nor U8916 (N_8916,N_7419,N_7489);
xnor U8917 (N_8917,N_7913,N_7953);
nand U8918 (N_8918,N_7669,N_7373);
nor U8919 (N_8919,N_7055,N_7251);
and U8920 (N_8920,N_7472,N_7935);
xor U8921 (N_8921,N_7788,N_7594);
nand U8922 (N_8922,N_7456,N_7791);
and U8923 (N_8923,N_7103,N_7989);
nand U8924 (N_8924,N_7238,N_7204);
nand U8925 (N_8925,N_7130,N_7865);
or U8926 (N_8926,N_7547,N_7061);
and U8927 (N_8927,N_7324,N_7745);
nand U8928 (N_8928,N_7011,N_7929);
nand U8929 (N_8929,N_7666,N_7398);
and U8930 (N_8930,N_7112,N_7636);
and U8931 (N_8931,N_7677,N_7251);
nor U8932 (N_8932,N_7046,N_7352);
xor U8933 (N_8933,N_7802,N_7060);
or U8934 (N_8934,N_7420,N_7763);
nor U8935 (N_8935,N_7149,N_7702);
and U8936 (N_8936,N_7125,N_7730);
xor U8937 (N_8937,N_7844,N_7863);
nor U8938 (N_8938,N_7665,N_7874);
or U8939 (N_8939,N_7033,N_7396);
nand U8940 (N_8940,N_7122,N_7561);
nand U8941 (N_8941,N_7753,N_7167);
nor U8942 (N_8942,N_7178,N_7393);
or U8943 (N_8943,N_7495,N_7550);
nand U8944 (N_8944,N_7824,N_7983);
xor U8945 (N_8945,N_7852,N_7977);
or U8946 (N_8946,N_7674,N_7271);
and U8947 (N_8947,N_7564,N_7383);
nand U8948 (N_8948,N_7780,N_7614);
nand U8949 (N_8949,N_7940,N_7712);
xnor U8950 (N_8950,N_7133,N_7950);
nor U8951 (N_8951,N_7431,N_7362);
nor U8952 (N_8952,N_7879,N_7748);
and U8953 (N_8953,N_7507,N_7032);
nand U8954 (N_8954,N_7643,N_7290);
or U8955 (N_8955,N_7709,N_7695);
xnor U8956 (N_8956,N_7062,N_7563);
or U8957 (N_8957,N_7279,N_7622);
nand U8958 (N_8958,N_7434,N_7528);
xor U8959 (N_8959,N_7956,N_7048);
nor U8960 (N_8960,N_7257,N_7350);
nand U8961 (N_8961,N_7271,N_7801);
nor U8962 (N_8962,N_7491,N_7697);
nand U8963 (N_8963,N_7975,N_7818);
and U8964 (N_8964,N_7166,N_7972);
nor U8965 (N_8965,N_7566,N_7469);
or U8966 (N_8966,N_7994,N_7506);
or U8967 (N_8967,N_7607,N_7187);
or U8968 (N_8968,N_7697,N_7620);
xnor U8969 (N_8969,N_7797,N_7365);
or U8970 (N_8970,N_7246,N_7140);
xor U8971 (N_8971,N_7355,N_7541);
and U8972 (N_8972,N_7534,N_7153);
xnor U8973 (N_8973,N_7082,N_7092);
or U8974 (N_8974,N_7045,N_7228);
nand U8975 (N_8975,N_7629,N_7910);
xor U8976 (N_8976,N_7374,N_7169);
xnor U8977 (N_8977,N_7674,N_7205);
nand U8978 (N_8978,N_7097,N_7382);
nor U8979 (N_8979,N_7618,N_7483);
or U8980 (N_8980,N_7929,N_7631);
nor U8981 (N_8981,N_7138,N_7509);
nor U8982 (N_8982,N_7558,N_7330);
nor U8983 (N_8983,N_7215,N_7041);
or U8984 (N_8984,N_7025,N_7168);
or U8985 (N_8985,N_7747,N_7507);
xnor U8986 (N_8986,N_7193,N_7271);
and U8987 (N_8987,N_7277,N_7805);
or U8988 (N_8988,N_7258,N_7787);
nor U8989 (N_8989,N_7303,N_7240);
xnor U8990 (N_8990,N_7100,N_7630);
nand U8991 (N_8991,N_7878,N_7421);
and U8992 (N_8992,N_7917,N_7019);
nand U8993 (N_8993,N_7989,N_7051);
nand U8994 (N_8994,N_7160,N_7546);
xor U8995 (N_8995,N_7595,N_7392);
nor U8996 (N_8996,N_7036,N_7977);
nand U8997 (N_8997,N_7652,N_7628);
and U8998 (N_8998,N_7337,N_7366);
nand U8999 (N_8999,N_7274,N_7394);
and U9000 (N_9000,N_8947,N_8618);
nand U9001 (N_9001,N_8382,N_8563);
xnor U9002 (N_9002,N_8379,N_8906);
nand U9003 (N_9003,N_8247,N_8227);
or U9004 (N_9004,N_8104,N_8323);
and U9005 (N_9005,N_8194,N_8029);
or U9006 (N_9006,N_8035,N_8437);
xnor U9007 (N_9007,N_8388,N_8102);
xnor U9008 (N_9008,N_8123,N_8335);
nand U9009 (N_9009,N_8549,N_8474);
or U9010 (N_9010,N_8584,N_8446);
and U9011 (N_9011,N_8482,N_8377);
and U9012 (N_9012,N_8415,N_8978);
nand U9013 (N_9013,N_8321,N_8418);
and U9014 (N_9014,N_8856,N_8435);
or U9015 (N_9015,N_8938,N_8538);
nand U9016 (N_9016,N_8897,N_8334);
nor U9017 (N_9017,N_8671,N_8070);
xor U9018 (N_9018,N_8619,N_8966);
nor U9019 (N_9019,N_8801,N_8440);
xnor U9020 (N_9020,N_8279,N_8343);
xor U9021 (N_9021,N_8506,N_8078);
nor U9022 (N_9022,N_8065,N_8235);
nor U9023 (N_9023,N_8698,N_8502);
nor U9024 (N_9024,N_8775,N_8848);
xnor U9025 (N_9025,N_8133,N_8011);
or U9026 (N_9026,N_8080,N_8036);
and U9027 (N_9027,N_8816,N_8489);
and U9028 (N_9028,N_8909,N_8164);
nor U9029 (N_9029,N_8114,N_8545);
xnor U9030 (N_9030,N_8772,N_8854);
xor U9031 (N_9031,N_8749,N_8900);
or U9032 (N_9032,N_8041,N_8789);
or U9033 (N_9033,N_8186,N_8941);
nand U9034 (N_9034,N_8218,N_8771);
and U9035 (N_9035,N_8627,N_8615);
or U9036 (N_9036,N_8439,N_8295);
nor U9037 (N_9037,N_8332,N_8600);
nand U9038 (N_9038,N_8449,N_8794);
and U9039 (N_9039,N_8460,N_8139);
or U9040 (N_9040,N_8048,N_8250);
nand U9041 (N_9041,N_8324,N_8406);
xor U9042 (N_9042,N_8173,N_8575);
xnor U9043 (N_9043,N_8708,N_8758);
xor U9044 (N_9044,N_8249,N_8242);
or U9045 (N_9045,N_8361,N_8371);
and U9046 (N_9046,N_8790,N_8764);
nor U9047 (N_9047,N_8229,N_8488);
nor U9048 (N_9048,N_8896,N_8980);
or U9049 (N_9049,N_8682,N_8369);
xnor U9050 (N_9050,N_8314,N_8889);
nand U9051 (N_9051,N_8714,N_8509);
and U9052 (N_9052,N_8798,N_8689);
or U9053 (N_9053,N_8562,N_8198);
nor U9054 (N_9054,N_8762,N_8113);
nand U9055 (N_9055,N_8776,N_8414);
nand U9056 (N_9056,N_8498,N_8802);
nor U9057 (N_9057,N_8731,N_8998);
and U9058 (N_9058,N_8788,N_8974);
xor U9059 (N_9059,N_8018,N_8803);
xnor U9060 (N_9060,N_8475,N_8611);
nand U9061 (N_9061,N_8092,N_8009);
nand U9062 (N_9062,N_8432,N_8521);
nand U9063 (N_9063,N_8337,N_8320);
and U9064 (N_9064,N_8958,N_8470);
nor U9065 (N_9065,N_8156,N_8913);
xor U9066 (N_9066,N_8777,N_8466);
xnor U9067 (N_9067,N_8716,N_8318);
and U9068 (N_9068,N_8541,N_8002);
and U9069 (N_9069,N_8677,N_8734);
nor U9070 (N_9070,N_8365,N_8039);
and U9071 (N_9071,N_8944,N_8328);
xor U9072 (N_9072,N_8037,N_8251);
xor U9073 (N_9073,N_8945,N_8725);
or U9074 (N_9074,N_8915,N_8931);
nor U9075 (N_9075,N_8225,N_8632);
nor U9076 (N_9076,N_8574,N_8026);
nor U9077 (N_9077,N_8867,N_8427);
or U9078 (N_9078,N_8013,N_8601);
xnor U9079 (N_9079,N_8292,N_8840);
and U9080 (N_9080,N_8955,N_8588);
xnor U9081 (N_9081,N_8638,N_8366);
and U9082 (N_9082,N_8479,N_8294);
xnor U9083 (N_9083,N_8110,N_8951);
and U9084 (N_9084,N_8461,N_8315);
nor U9085 (N_9085,N_8701,N_8697);
nand U9086 (N_9086,N_8744,N_8643);
nor U9087 (N_9087,N_8252,N_8617);
nor U9088 (N_9088,N_8103,N_8399);
and U9089 (N_9089,N_8231,N_8878);
or U9090 (N_9090,N_8120,N_8407);
nor U9091 (N_9091,N_8880,N_8519);
xnor U9092 (N_9092,N_8357,N_8203);
nor U9093 (N_9093,N_8747,N_8968);
or U9094 (N_9094,N_8850,N_8459);
nor U9095 (N_9095,N_8016,N_8137);
xnor U9096 (N_9096,N_8637,N_8278);
nor U9097 (N_9097,N_8926,N_8171);
and U9098 (N_9098,N_8759,N_8547);
or U9099 (N_9099,N_8993,N_8580);
or U9100 (N_9100,N_8924,N_8756);
nand U9101 (N_9101,N_8720,N_8391);
nor U9102 (N_9102,N_8319,N_8515);
xor U9103 (N_9103,N_8675,N_8626);
nand U9104 (N_9104,N_8015,N_8606);
and U9105 (N_9105,N_8179,N_8864);
nor U9106 (N_9106,N_8115,N_8411);
xor U9107 (N_9107,N_8471,N_8478);
nand U9108 (N_9108,N_8034,N_8674);
and U9109 (N_9109,N_8565,N_8290);
nor U9110 (N_9110,N_8276,N_8654);
nor U9111 (N_9111,N_8151,N_8539);
and U9112 (N_9112,N_8793,N_8526);
xor U9113 (N_9113,N_8973,N_8902);
and U9114 (N_9114,N_8395,N_8901);
nor U9115 (N_9115,N_8346,N_8063);
nand U9116 (N_9116,N_8212,N_8508);
or U9117 (N_9117,N_8283,N_8281);
nor U9118 (N_9118,N_8397,N_8305);
or U9119 (N_9119,N_8594,N_8722);
nand U9120 (N_9120,N_8327,N_8806);
nand U9121 (N_9121,N_8069,N_8903);
xor U9122 (N_9122,N_8686,N_8936);
and U9123 (N_9123,N_8707,N_8717);
or U9124 (N_9124,N_8792,N_8704);
or U9125 (N_9125,N_8797,N_8359);
xnor U9126 (N_9126,N_8917,N_8303);
or U9127 (N_9127,N_8165,N_8271);
and U9128 (N_9128,N_8989,N_8001);
xor U9129 (N_9129,N_8969,N_8044);
nor U9130 (N_9130,N_8946,N_8831);
nor U9131 (N_9131,N_8464,N_8954);
or U9132 (N_9132,N_8991,N_8086);
nand U9133 (N_9133,N_8378,N_8807);
xor U9134 (N_9134,N_8025,N_8429);
nand U9135 (N_9135,N_8064,N_8384);
or U9136 (N_9136,N_8804,N_8809);
nand U9137 (N_9137,N_8649,N_8140);
xor U9138 (N_9138,N_8970,N_8887);
nor U9139 (N_9139,N_8465,N_8648);
nand U9140 (N_9140,N_8373,N_8669);
and U9141 (N_9141,N_8061,N_8285);
nand U9142 (N_9142,N_8702,N_8472);
nand U9143 (N_9143,N_8892,N_8483);
and U9144 (N_9144,N_8254,N_8665);
or U9145 (N_9145,N_8490,N_8263);
nand U9146 (N_9146,N_8260,N_8265);
nor U9147 (N_9147,N_8999,N_8268);
nor U9148 (N_9148,N_8270,N_8888);
and U9149 (N_9149,N_8839,N_8197);
and U9150 (N_9150,N_8525,N_8233);
nor U9151 (N_9151,N_8814,N_8501);
or U9152 (N_9152,N_8659,N_8841);
nor U9153 (N_9153,N_8972,N_8885);
or U9154 (N_9154,N_8925,N_8031);
nor U9155 (N_9155,N_8291,N_8004);
and U9156 (N_9156,N_8293,N_8134);
or U9157 (N_9157,N_8201,N_8129);
nor U9158 (N_9158,N_8805,N_8554);
or U9159 (N_9159,N_8929,N_8769);
or U9160 (N_9160,N_8213,N_8605);
or U9161 (N_9161,N_8612,N_8530);
and U9162 (N_9162,N_8275,N_8083);
nor U9163 (N_9163,N_8799,N_8193);
xnor U9164 (N_9164,N_8907,N_8985);
and U9165 (N_9165,N_8301,N_8053);
xnor U9166 (N_9166,N_8299,N_8891);
nand U9167 (N_9167,N_8076,N_8322);
and U9168 (N_9168,N_8564,N_8842);
nand U9169 (N_9169,N_8154,N_8094);
nor U9170 (N_9170,N_8352,N_8658);
xnor U9171 (N_9171,N_8264,N_8934);
or U9172 (N_9172,N_8633,N_8215);
and U9173 (N_9173,N_8082,N_8870);
nand U9174 (N_9174,N_8780,N_8400);
or U9175 (N_9175,N_8224,N_8810);
nand U9176 (N_9176,N_8098,N_8222);
or U9177 (N_9177,N_8928,N_8317);
nand U9178 (N_9178,N_8485,N_8454);
nand U9179 (N_9179,N_8298,N_8830);
xor U9180 (N_9180,N_8623,N_8005);
or U9181 (N_9181,N_8206,N_8784);
nand U9182 (N_9182,N_8024,N_8835);
nor U9183 (N_9183,N_8811,N_8676);
and U9184 (N_9184,N_8308,N_8650);
and U9185 (N_9185,N_8239,N_8862);
or U9186 (N_9186,N_8117,N_8656);
and U9187 (N_9187,N_8057,N_8942);
nor U9188 (N_9188,N_8097,N_8138);
nor U9189 (N_9189,N_8095,N_8107);
nand U9190 (N_9190,N_8067,N_8778);
or U9191 (N_9191,N_8188,N_8863);
nor U9192 (N_9192,N_8723,N_8681);
xor U9193 (N_9193,N_8006,N_8949);
and U9194 (N_9194,N_8458,N_8306);
or U9195 (N_9195,N_8948,N_8937);
or U9196 (N_9196,N_8499,N_8345);
or U9197 (N_9197,N_8886,N_8693);
and U9198 (N_9198,N_8423,N_8826);
nor U9199 (N_9199,N_8409,N_8073);
nand U9200 (N_9200,N_8122,N_8551);
or U9201 (N_9201,N_8195,N_8401);
xnor U9202 (N_9202,N_8592,N_8553);
or U9203 (N_9203,N_8713,N_8899);
or U9204 (N_9204,N_8130,N_8010);
and U9205 (N_9205,N_8914,N_8438);
xnor U9206 (N_9206,N_8149,N_8680);
or U9207 (N_9207,N_8843,N_8868);
nor U9208 (N_9208,N_8786,N_8480);
and U9209 (N_9209,N_8209,N_8641);
and U9210 (N_9210,N_8736,N_8576);
nor U9211 (N_9211,N_8694,N_8766);
and U9212 (N_9212,N_8000,N_8703);
nand U9213 (N_9213,N_8939,N_8277);
nor U9214 (N_9214,N_8017,N_8834);
xor U9215 (N_9215,N_8516,N_8248);
xor U9216 (N_9216,N_8963,N_8211);
nor U9217 (N_9217,N_8597,N_8524);
nor U9218 (N_9218,N_8548,N_8404);
xor U9219 (N_9219,N_8071,N_8774);
xor U9220 (N_9220,N_8598,N_8770);
and U9221 (N_9221,N_8696,N_8312);
or U9222 (N_9222,N_8257,N_8640);
xnor U9223 (N_9223,N_8241,N_8685);
nand U9224 (N_9224,N_8090,N_8416);
or U9225 (N_9225,N_8741,N_8825);
nand U9226 (N_9226,N_8559,N_8486);
nand U9227 (N_9227,N_8495,N_8746);
and U9228 (N_9228,N_8660,N_8583);
or U9229 (N_9229,N_8136,N_8145);
nor U9230 (N_9230,N_8922,N_8787);
nand U9231 (N_9231,N_8668,N_8497);
nand U9232 (N_9232,N_8040,N_8341);
nor U9233 (N_9233,N_8255,N_8779);
and U9234 (N_9234,N_8355,N_8300);
nor U9235 (N_9235,N_8818,N_8331);
xor U9236 (N_9236,N_8829,N_8628);
nor U9237 (N_9237,N_8467,N_8520);
and U9238 (N_9238,N_8441,N_8182);
or U9239 (N_9239,N_8170,N_8531);
xor U9240 (N_9240,N_8661,N_8977);
or U9241 (N_9241,N_8216,N_8108);
and U9242 (N_9242,N_8493,N_8473);
or U9243 (N_9243,N_8570,N_8023);
and U9244 (N_9244,N_8236,N_8603);
nor U9245 (N_9245,N_8128,N_8160);
nor U9246 (N_9246,N_8566,N_8838);
and U9247 (N_9247,N_8911,N_8819);
xnor U9248 (N_9248,N_8121,N_8262);
or U9249 (N_9249,N_8066,N_8940);
and U9250 (N_9250,N_8372,N_8056);
nand U9251 (N_9251,N_8782,N_8672);
or U9252 (N_9252,N_8463,N_8032);
nor U9253 (N_9253,N_8246,N_8020);
or U9254 (N_9254,N_8043,N_8979);
and U9255 (N_9255,N_8150,N_8709);
or U9256 (N_9256,N_8118,N_8853);
or U9257 (N_9257,N_8394,N_8177);
and U9258 (N_9258,N_8132,N_8943);
nand U9259 (N_9259,N_8904,N_8923);
or U9260 (N_9260,N_8217,N_8971);
and U9261 (N_9261,N_8599,N_8112);
or U9262 (N_9262,N_8296,N_8921);
or U9263 (N_9263,N_8072,N_8214);
and U9264 (N_9264,N_8815,N_8935);
and U9265 (N_9265,N_8109,N_8760);
nand U9266 (N_9266,N_8748,N_8166);
and U9267 (N_9267,N_8644,N_8191);
xor U9268 (N_9268,N_8105,N_8253);
or U9269 (N_9269,N_8402,N_8245);
or U9270 (N_9270,N_8106,N_8865);
xnor U9271 (N_9271,N_8712,N_8930);
and U9272 (N_9272,N_8392,N_8230);
nor U9273 (N_9273,N_8890,N_8845);
nand U9274 (N_9274,N_8424,N_8325);
nor U9275 (N_9275,N_8101,N_8536);
nor U9276 (N_9276,N_8386,N_8522);
nor U9277 (N_9277,N_8837,N_8153);
xnor U9278 (N_9278,N_8161,N_8577);
nor U9279 (N_9279,N_8645,N_8302);
nand U9280 (N_9280,N_8898,N_8857);
or U9281 (N_9281,N_8822,N_8695);
and U9282 (N_9282,N_8091,N_8965);
nor U9283 (N_9283,N_8368,N_8569);
or U9284 (N_9284,N_8162,N_8381);
or U9285 (N_9285,N_8148,N_8204);
xor U9286 (N_9286,N_8436,N_8316);
nor U9287 (N_9287,N_8986,N_8718);
xnor U9288 (N_9288,N_8492,N_8705);
xnor U9289 (N_9289,N_8866,N_8087);
nand U9290 (N_9290,N_8403,N_8421);
and U9291 (N_9291,N_8221,N_8052);
and U9292 (N_9292,N_8950,N_8593);
nor U9293 (N_9293,N_8196,N_8019);
or U9294 (N_9294,N_8434,N_8131);
xnor U9295 (N_9295,N_8340,N_8860);
nand U9296 (N_9296,N_8846,N_8568);
nor U9297 (N_9297,N_8651,N_8126);
nand U9298 (N_9298,N_8587,N_8510);
nand U9299 (N_9299,N_8163,N_8099);
or U9300 (N_9300,N_8243,N_8550);
and U9301 (N_9301,N_8363,N_8918);
nand U9302 (N_9302,N_8710,N_8393);
nor U9303 (N_9303,N_8096,N_8742);
and U9304 (N_9304,N_8721,N_8111);
xor U9305 (N_9305,N_8932,N_8625);
nor U9306 (N_9306,N_8679,N_8876);
xor U9307 (N_9307,N_8518,N_8062);
xnor U9308 (N_9308,N_8635,N_8431);
nor U9309 (N_9309,N_8663,N_8175);
nor U9310 (N_9310,N_8157,N_8445);
xnor U9311 (N_9311,N_8042,N_8873);
or U9312 (N_9312,N_8706,N_8205);
nand U9313 (N_9313,N_8387,N_8074);
and U9314 (N_9314,N_8630,N_8785);
nor U9315 (N_9315,N_8389,N_8184);
or U9316 (N_9316,N_8959,N_8750);
nand U9317 (N_9317,N_8738,N_8093);
or U9318 (N_9318,N_8496,N_8961);
nand U9319 (N_9319,N_8028,N_8994);
and U9320 (N_9320,N_8084,N_8505);
xnor U9321 (N_9321,N_8622,N_8143);
nor U9322 (N_9322,N_8517,N_8513);
and U9323 (N_9323,N_8060,N_8152);
xnor U9324 (N_9324,N_8982,N_8457);
nor U9325 (N_9325,N_8220,N_8158);
xor U9326 (N_9326,N_8456,N_8621);
nand U9327 (N_9327,N_8666,N_8988);
nor U9328 (N_9328,N_8752,N_8874);
xnor U9329 (N_9329,N_8282,N_8861);
and U9330 (N_9330,N_8202,N_8311);
or U9331 (N_9331,N_8307,N_8330);
xnor U9332 (N_9332,N_8552,N_8085);
and U9333 (N_9333,N_8012,N_8425);
xnor U9334 (N_9334,N_8884,N_8228);
xnor U9335 (N_9335,N_8375,N_8952);
nand U9336 (N_9336,N_8178,N_8992);
nand U9337 (N_9337,N_8767,N_8054);
nand U9338 (N_9338,N_8956,N_8269);
xnor U9339 (N_9339,N_8560,N_8356);
xnor U9340 (N_9340,N_8181,N_8444);
nand U9341 (N_9341,N_8849,N_8894);
nor U9342 (N_9342,N_8667,N_8983);
nand U9343 (N_9343,N_8507,N_8288);
or U9344 (N_9344,N_8544,N_8755);
and U9345 (N_9345,N_8610,N_8730);
xor U9346 (N_9346,N_8629,N_8116);
nor U9347 (N_9347,N_8207,N_8075);
or U9348 (N_9348,N_8670,N_8146);
xor U9349 (N_9349,N_8477,N_8620);
or U9350 (N_9350,N_8646,N_8996);
and U9351 (N_9351,N_8326,N_8180);
nand U9352 (N_9352,N_8573,N_8190);
and U9353 (N_9353,N_8699,N_8364);
xnor U9354 (N_9354,N_8280,N_8881);
xnor U9355 (N_9355,N_8155,N_8183);
nor U9356 (N_9356,N_8591,N_8127);
nand U9357 (N_9357,N_8763,N_8455);
xor U9358 (N_9358,N_8021,N_8125);
or U9359 (N_9359,N_8244,N_8273);
or U9360 (N_9360,N_8419,N_8259);
xor U9361 (N_9361,N_8827,N_8266);
xnor U9362 (N_9362,N_8187,N_8624);
and U9363 (N_9363,N_8893,N_8284);
nor U9364 (N_9364,N_8199,N_8022);
nor U9365 (N_9365,N_8543,N_8791);
nor U9366 (N_9366,N_8310,N_8313);
xnor U9367 (N_9367,N_8351,N_8353);
xor U9368 (N_9368,N_8586,N_8726);
nand U9369 (N_9369,N_8567,N_8049);
nand U9370 (N_9370,N_8875,N_8967);
or U9371 (N_9371,N_8529,N_8634);
nand U9372 (N_9372,N_8542,N_8494);
nand U9373 (N_9373,N_8727,N_8561);
and U9374 (N_9374,N_8412,N_8754);
xnor U9375 (N_9375,N_8582,N_8579);
and U9376 (N_9376,N_8813,N_8908);
nor U9377 (N_9377,N_8200,N_8339);
or U9378 (N_9378,N_8267,N_8329);
and U9379 (N_9379,N_8426,N_8050);
and U9380 (N_9380,N_8773,N_8558);
and U9381 (N_9381,N_8410,N_8442);
xnor U9382 (N_9382,N_8398,N_8528);
xnor U9383 (N_9383,N_8079,N_8927);
nand U9384 (N_9384,N_8910,N_8783);
or U9385 (N_9385,N_8383,N_8503);
or U9386 (N_9386,N_8468,N_8385);
xnor U9387 (N_9387,N_8333,N_8589);
xor U9388 (N_9388,N_8405,N_8688);
nand U9389 (N_9389,N_8167,N_8858);
xnor U9390 (N_9390,N_8417,N_8443);
nor U9391 (N_9391,N_8557,N_8657);
nand U9392 (N_9392,N_8274,N_8692);
and U9393 (N_9393,N_8662,N_8124);
and U9394 (N_9394,N_8871,N_8823);
nor U9395 (N_9395,N_8609,N_8844);
nand U9396 (N_9396,N_8367,N_8537);
nand U9397 (N_9397,N_8753,N_8350);
nand U9398 (N_9398,N_8691,N_8481);
nor U9399 (N_9399,N_8751,N_8534);
nor U9400 (N_9400,N_8261,N_8344);
and U9401 (N_9401,N_8141,N_8514);
xor U9402 (N_9402,N_8487,N_8176);
nor U9403 (N_9403,N_8990,N_8309);
and U9404 (N_9404,N_8757,N_8639);
nand U9405 (N_9405,N_8504,N_8362);
nor U9406 (N_9406,N_8882,N_8739);
nand U9407 (N_9407,N_8919,N_8135);
and U9408 (N_9408,N_8500,N_8808);
or U9409 (N_9409,N_8546,N_8354);
or U9410 (N_9410,N_8535,N_8533);
and U9411 (N_9411,N_8761,N_8572);
and U9412 (N_9412,N_8690,N_8172);
nor U9413 (N_9413,N_8003,N_8453);
xnor U9414 (N_9414,N_8046,N_8684);
nand U9415 (N_9415,N_8348,N_8824);
nand U9416 (N_9416,N_8912,N_8030);
or U9417 (N_9417,N_8119,N_8008);
nor U9418 (N_9418,N_8847,N_8523);
or U9419 (N_9419,N_8995,N_8859);
nand U9420 (N_9420,N_8740,N_8223);
and U9421 (N_9421,N_8142,N_8174);
and U9422 (N_9422,N_8879,N_8719);
or U9423 (N_9423,N_8532,N_8984);
or U9424 (N_9424,N_8877,N_8540);
and U9425 (N_9425,N_8219,N_8745);
nor U9426 (N_9426,N_8883,N_8976);
nor U9427 (N_9427,N_8484,N_8964);
or U9428 (N_9428,N_8595,N_8447);
nor U9429 (N_9429,N_8608,N_8555);
and U9430 (N_9430,N_8855,N_8578);
nor U9431 (N_9431,N_8590,N_8981);
nor U9432 (N_9432,N_8338,N_8962);
and U9433 (N_9433,N_8581,N_8408);
and U9434 (N_9434,N_8428,N_8728);
and U9435 (N_9435,N_8724,N_8729);
nand U9436 (N_9436,N_8370,N_8512);
xor U9437 (N_9437,N_8602,N_8647);
xnor U9438 (N_9438,N_8422,N_8256);
xnor U9439 (N_9439,N_8795,N_8081);
and U9440 (N_9440,N_8433,N_8452);
nand U9441 (N_9441,N_8068,N_8851);
xor U9442 (N_9442,N_8652,N_8047);
or U9443 (N_9443,N_8585,N_8869);
nand U9444 (N_9444,N_8304,N_8347);
and U9445 (N_9445,N_8413,N_8715);
and U9446 (N_9446,N_8683,N_8616);
or U9447 (N_9447,N_8975,N_8916);
and U9448 (N_9448,N_8089,N_8192);
nand U9449 (N_9449,N_8737,N_8821);
xnor U9450 (N_9450,N_8476,N_8051);
nand U9451 (N_9451,N_8933,N_8895);
nor U9452 (N_9452,N_8007,N_8655);
or U9453 (N_9453,N_8957,N_8232);
nand U9454 (N_9454,N_8058,N_8059);
nand U9455 (N_9455,N_8642,N_8358);
and U9456 (N_9456,N_8342,N_8817);
xnor U9457 (N_9457,N_8380,N_8636);
nand U9458 (N_9458,N_8297,N_8872);
and U9459 (N_9459,N_8027,N_8100);
xor U9460 (N_9460,N_8189,N_8820);
nor U9461 (N_9461,N_8376,N_8208);
and U9462 (N_9462,N_8234,N_8905);
nor U9463 (N_9463,N_8556,N_8953);
and U9464 (N_9464,N_8833,N_8613);
xnor U9465 (N_9465,N_8038,N_8077);
and U9466 (N_9466,N_8796,N_8664);
or U9467 (N_9467,N_8169,N_8604);
and U9468 (N_9468,N_8374,N_8700);
nand U9469 (N_9469,N_8287,N_8289);
or U9470 (N_9470,N_8144,N_8420);
or U9471 (N_9471,N_8055,N_8735);
or U9472 (N_9472,N_8687,N_8768);
or U9473 (N_9473,N_8360,N_8396);
and U9474 (N_9474,N_8185,N_8226);
xnor U9475 (N_9475,N_8852,N_8781);
or U9476 (N_9476,N_8448,N_8240);
or U9477 (N_9477,N_8987,N_8430);
or U9478 (N_9478,N_8765,N_8571);
nand U9479 (N_9479,N_8733,N_8653);
xor U9480 (N_9480,N_8511,N_8462);
nor U9481 (N_9481,N_8159,N_8469);
nand U9482 (N_9482,N_8147,N_8168);
nand U9483 (N_9483,N_8920,N_8491);
nor U9484 (N_9484,N_8349,N_8258);
nor U9485 (N_9485,N_8238,N_8088);
nor U9486 (N_9486,N_8596,N_8631);
or U9487 (N_9487,N_8450,N_8014);
xor U9488 (N_9488,N_8607,N_8673);
xor U9489 (N_9489,N_8960,N_8336);
nand U9490 (N_9490,N_8527,N_8237);
nand U9491 (N_9491,N_8033,N_8812);
or U9492 (N_9492,N_8800,N_8711);
nor U9493 (N_9493,N_8678,N_8210);
nand U9494 (N_9494,N_8828,N_8732);
nand U9495 (N_9495,N_8832,N_8451);
and U9496 (N_9496,N_8390,N_8743);
and U9497 (N_9497,N_8997,N_8286);
xor U9498 (N_9498,N_8614,N_8836);
nand U9499 (N_9499,N_8045,N_8272);
xor U9500 (N_9500,N_8402,N_8435);
nand U9501 (N_9501,N_8530,N_8443);
xor U9502 (N_9502,N_8157,N_8464);
and U9503 (N_9503,N_8348,N_8355);
and U9504 (N_9504,N_8364,N_8691);
xnor U9505 (N_9505,N_8919,N_8729);
xnor U9506 (N_9506,N_8206,N_8495);
xor U9507 (N_9507,N_8414,N_8105);
or U9508 (N_9508,N_8273,N_8893);
or U9509 (N_9509,N_8731,N_8780);
xor U9510 (N_9510,N_8130,N_8221);
and U9511 (N_9511,N_8152,N_8609);
and U9512 (N_9512,N_8564,N_8671);
xnor U9513 (N_9513,N_8058,N_8398);
and U9514 (N_9514,N_8848,N_8448);
xnor U9515 (N_9515,N_8816,N_8632);
nand U9516 (N_9516,N_8708,N_8956);
and U9517 (N_9517,N_8136,N_8662);
nor U9518 (N_9518,N_8465,N_8081);
or U9519 (N_9519,N_8663,N_8973);
xor U9520 (N_9520,N_8299,N_8496);
xor U9521 (N_9521,N_8217,N_8505);
and U9522 (N_9522,N_8741,N_8496);
or U9523 (N_9523,N_8667,N_8251);
nor U9524 (N_9524,N_8682,N_8886);
and U9525 (N_9525,N_8399,N_8433);
xor U9526 (N_9526,N_8952,N_8403);
or U9527 (N_9527,N_8366,N_8933);
nor U9528 (N_9528,N_8965,N_8328);
nor U9529 (N_9529,N_8265,N_8586);
nor U9530 (N_9530,N_8025,N_8897);
nand U9531 (N_9531,N_8491,N_8778);
nand U9532 (N_9532,N_8793,N_8100);
nand U9533 (N_9533,N_8906,N_8645);
or U9534 (N_9534,N_8219,N_8873);
nand U9535 (N_9535,N_8266,N_8115);
xnor U9536 (N_9536,N_8287,N_8007);
and U9537 (N_9537,N_8499,N_8481);
xnor U9538 (N_9538,N_8128,N_8215);
nand U9539 (N_9539,N_8696,N_8429);
and U9540 (N_9540,N_8134,N_8410);
or U9541 (N_9541,N_8312,N_8460);
nand U9542 (N_9542,N_8308,N_8215);
nor U9543 (N_9543,N_8454,N_8164);
xnor U9544 (N_9544,N_8844,N_8877);
and U9545 (N_9545,N_8703,N_8527);
nand U9546 (N_9546,N_8261,N_8188);
nand U9547 (N_9547,N_8764,N_8294);
xor U9548 (N_9548,N_8641,N_8005);
xnor U9549 (N_9549,N_8447,N_8765);
xnor U9550 (N_9550,N_8922,N_8460);
or U9551 (N_9551,N_8393,N_8331);
nand U9552 (N_9552,N_8685,N_8746);
nand U9553 (N_9553,N_8225,N_8979);
nor U9554 (N_9554,N_8684,N_8649);
nand U9555 (N_9555,N_8265,N_8620);
and U9556 (N_9556,N_8230,N_8662);
nand U9557 (N_9557,N_8058,N_8586);
or U9558 (N_9558,N_8620,N_8906);
or U9559 (N_9559,N_8141,N_8875);
nand U9560 (N_9560,N_8912,N_8110);
nand U9561 (N_9561,N_8232,N_8304);
nand U9562 (N_9562,N_8401,N_8104);
nand U9563 (N_9563,N_8101,N_8673);
nand U9564 (N_9564,N_8220,N_8469);
and U9565 (N_9565,N_8976,N_8280);
xor U9566 (N_9566,N_8097,N_8629);
xor U9567 (N_9567,N_8226,N_8644);
and U9568 (N_9568,N_8662,N_8691);
nand U9569 (N_9569,N_8170,N_8244);
nor U9570 (N_9570,N_8387,N_8965);
and U9571 (N_9571,N_8234,N_8422);
or U9572 (N_9572,N_8232,N_8194);
nor U9573 (N_9573,N_8094,N_8808);
nor U9574 (N_9574,N_8666,N_8068);
or U9575 (N_9575,N_8697,N_8568);
nand U9576 (N_9576,N_8144,N_8108);
or U9577 (N_9577,N_8753,N_8686);
and U9578 (N_9578,N_8106,N_8736);
nor U9579 (N_9579,N_8507,N_8109);
or U9580 (N_9580,N_8896,N_8489);
or U9581 (N_9581,N_8771,N_8968);
nand U9582 (N_9582,N_8113,N_8718);
nor U9583 (N_9583,N_8348,N_8234);
and U9584 (N_9584,N_8996,N_8099);
or U9585 (N_9585,N_8094,N_8790);
nand U9586 (N_9586,N_8526,N_8980);
nand U9587 (N_9587,N_8361,N_8054);
nand U9588 (N_9588,N_8795,N_8592);
nand U9589 (N_9589,N_8622,N_8061);
and U9590 (N_9590,N_8570,N_8958);
or U9591 (N_9591,N_8850,N_8183);
or U9592 (N_9592,N_8736,N_8586);
or U9593 (N_9593,N_8442,N_8304);
or U9594 (N_9594,N_8424,N_8500);
nor U9595 (N_9595,N_8082,N_8234);
or U9596 (N_9596,N_8865,N_8440);
nand U9597 (N_9597,N_8981,N_8226);
nor U9598 (N_9598,N_8214,N_8217);
nand U9599 (N_9599,N_8189,N_8537);
or U9600 (N_9600,N_8547,N_8837);
xor U9601 (N_9601,N_8226,N_8604);
nand U9602 (N_9602,N_8840,N_8832);
nand U9603 (N_9603,N_8738,N_8930);
and U9604 (N_9604,N_8145,N_8016);
nor U9605 (N_9605,N_8697,N_8168);
or U9606 (N_9606,N_8856,N_8739);
nor U9607 (N_9607,N_8749,N_8084);
nand U9608 (N_9608,N_8067,N_8756);
xnor U9609 (N_9609,N_8296,N_8070);
or U9610 (N_9610,N_8208,N_8463);
xor U9611 (N_9611,N_8168,N_8901);
nor U9612 (N_9612,N_8082,N_8783);
or U9613 (N_9613,N_8846,N_8680);
or U9614 (N_9614,N_8245,N_8998);
and U9615 (N_9615,N_8995,N_8797);
nand U9616 (N_9616,N_8412,N_8889);
xor U9617 (N_9617,N_8735,N_8407);
nor U9618 (N_9618,N_8473,N_8444);
nand U9619 (N_9619,N_8271,N_8849);
xnor U9620 (N_9620,N_8958,N_8006);
nand U9621 (N_9621,N_8666,N_8474);
or U9622 (N_9622,N_8299,N_8362);
nor U9623 (N_9623,N_8730,N_8864);
or U9624 (N_9624,N_8590,N_8495);
and U9625 (N_9625,N_8219,N_8306);
xnor U9626 (N_9626,N_8769,N_8826);
and U9627 (N_9627,N_8985,N_8886);
nor U9628 (N_9628,N_8332,N_8452);
xnor U9629 (N_9629,N_8982,N_8075);
nand U9630 (N_9630,N_8958,N_8416);
and U9631 (N_9631,N_8134,N_8056);
and U9632 (N_9632,N_8694,N_8742);
nand U9633 (N_9633,N_8155,N_8458);
and U9634 (N_9634,N_8982,N_8307);
nand U9635 (N_9635,N_8820,N_8379);
nand U9636 (N_9636,N_8661,N_8298);
and U9637 (N_9637,N_8668,N_8714);
nor U9638 (N_9638,N_8610,N_8366);
and U9639 (N_9639,N_8673,N_8740);
nor U9640 (N_9640,N_8399,N_8771);
or U9641 (N_9641,N_8041,N_8353);
or U9642 (N_9642,N_8147,N_8166);
nand U9643 (N_9643,N_8225,N_8103);
nand U9644 (N_9644,N_8827,N_8245);
xnor U9645 (N_9645,N_8114,N_8506);
and U9646 (N_9646,N_8404,N_8239);
xor U9647 (N_9647,N_8745,N_8135);
nand U9648 (N_9648,N_8512,N_8776);
nand U9649 (N_9649,N_8479,N_8072);
and U9650 (N_9650,N_8568,N_8820);
or U9651 (N_9651,N_8005,N_8730);
or U9652 (N_9652,N_8195,N_8917);
nor U9653 (N_9653,N_8292,N_8006);
and U9654 (N_9654,N_8851,N_8291);
xnor U9655 (N_9655,N_8895,N_8133);
and U9656 (N_9656,N_8998,N_8929);
nor U9657 (N_9657,N_8030,N_8523);
xor U9658 (N_9658,N_8346,N_8521);
nand U9659 (N_9659,N_8493,N_8484);
or U9660 (N_9660,N_8074,N_8726);
and U9661 (N_9661,N_8955,N_8238);
nor U9662 (N_9662,N_8798,N_8144);
nor U9663 (N_9663,N_8750,N_8512);
and U9664 (N_9664,N_8024,N_8415);
nand U9665 (N_9665,N_8332,N_8519);
and U9666 (N_9666,N_8760,N_8358);
xor U9667 (N_9667,N_8884,N_8414);
nor U9668 (N_9668,N_8662,N_8746);
and U9669 (N_9669,N_8603,N_8382);
xor U9670 (N_9670,N_8460,N_8808);
and U9671 (N_9671,N_8275,N_8503);
and U9672 (N_9672,N_8568,N_8292);
xnor U9673 (N_9673,N_8822,N_8517);
or U9674 (N_9674,N_8326,N_8329);
xnor U9675 (N_9675,N_8060,N_8059);
nand U9676 (N_9676,N_8263,N_8711);
xnor U9677 (N_9677,N_8642,N_8774);
nor U9678 (N_9678,N_8539,N_8528);
and U9679 (N_9679,N_8746,N_8546);
or U9680 (N_9680,N_8234,N_8854);
nand U9681 (N_9681,N_8479,N_8015);
and U9682 (N_9682,N_8641,N_8321);
or U9683 (N_9683,N_8813,N_8208);
nand U9684 (N_9684,N_8305,N_8362);
nand U9685 (N_9685,N_8351,N_8899);
and U9686 (N_9686,N_8162,N_8619);
xnor U9687 (N_9687,N_8079,N_8048);
and U9688 (N_9688,N_8864,N_8674);
and U9689 (N_9689,N_8502,N_8899);
and U9690 (N_9690,N_8838,N_8784);
nor U9691 (N_9691,N_8367,N_8847);
nand U9692 (N_9692,N_8290,N_8724);
and U9693 (N_9693,N_8949,N_8239);
or U9694 (N_9694,N_8695,N_8226);
and U9695 (N_9695,N_8323,N_8068);
nor U9696 (N_9696,N_8973,N_8361);
or U9697 (N_9697,N_8083,N_8931);
xnor U9698 (N_9698,N_8073,N_8852);
nand U9699 (N_9699,N_8598,N_8467);
nor U9700 (N_9700,N_8457,N_8243);
xnor U9701 (N_9701,N_8830,N_8984);
xor U9702 (N_9702,N_8327,N_8502);
xor U9703 (N_9703,N_8876,N_8823);
or U9704 (N_9704,N_8698,N_8936);
nor U9705 (N_9705,N_8096,N_8301);
or U9706 (N_9706,N_8032,N_8829);
xor U9707 (N_9707,N_8937,N_8880);
and U9708 (N_9708,N_8778,N_8506);
nand U9709 (N_9709,N_8833,N_8940);
nor U9710 (N_9710,N_8372,N_8533);
or U9711 (N_9711,N_8827,N_8870);
or U9712 (N_9712,N_8802,N_8806);
nor U9713 (N_9713,N_8443,N_8049);
xnor U9714 (N_9714,N_8175,N_8138);
nand U9715 (N_9715,N_8796,N_8443);
or U9716 (N_9716,N_8869,N_8380);
and U9717 (N_9717,N_8360,N_8442);
and U9718 (N_9718,N_8401,N_8421);
and U9719 (N_9719,N_8733,N_8418);
and U9720 (N_9720,N_8052,N_8365);
xnor U9721 (N_9721,N_8902,N_8008);
xnor U9722 (N_9722,N_8498,N_8257);
nor U9723 (N_9723,N_8003,N_8512);
xnor U9724 (N_9724,N_8191,N_8622);
or U9725 (N_9725,N_8226,N_8620);
nor U9726 (N_9726,N_8633,N_8905);
or U9727 (N_9727,N_8763,N_8449);
nand U9728 (N_9728,N_8137,N_8515);
or U9729 (N_9729,N_8173,N_8465);
and U9730 (N_9730,N_8111,N_8549);
nand U9731 (N_9731,N_8359,N_8563);
nor U9732 (N_9732,N_8095,N_8351);
or U9733 (N_9733,N_8602,N_8410);
nor U9734 (N_9734,N_8577,N_8826);
nor U9735 (N_9735,N_8161,N_8552);
or U9736 (N_9736,N_8996,N_8270);
nor U9737 (N_9737,N_8743,N_8420);
or U9738 (N_9738,N_8587,N_8520);
nand U9739 (N_9739,N_8644,N_8684);
nand U9740 (N_9740,N_8334,N_8618);
nor U9741 (N_9741,N_8968,N_8941);
and U9742 (N_9742,N_8018,N_8918);
or U9743 (N_9743,N_8611,N_8203);
and U9744 (N_9744,N_8548,N_8445);
or U9745 (N_9745,N_8358,N_8587);
or U9746 (N_9746,N_8138,N_8123);
or U9747 (N_9747,N_8705,N_8450);
or U9748 (N_9748,N_8108,N_8473);
nand U9749 (N_9749,N_8884,N_8400);
and U9750 (N_9750,N_8454,N_8254);
nand U9751 (N_9751,N_8657,N_8643);
nand U9752 (N_9752,N_8581,N_8497);
or U9753 (N_9753,N_8864,N_8217);
nor U9754 (N_9754,N_8986,N_8544);
or U9755 (N_9755,N_8848,N_8466);
nor U9756 (N_9756,N_8508,N_8426);
nand U9757 (N_9757,N_8927,N_8572);
and U9758 (N_9758,N_8109,N_8208);
or U9759 (N_9759,N_8255,N_8751);
xnor U9760 (N_9760,N_8522,N_8444);
xor U9761 (N_9761,N_8219,N_8906);
xor U9762 (N_9762,N_8842,N_8737);
nor U9763 (N_9763,N_8278,N_8050);
or U9764 (N_9764,N_8189,N_8366);
or U9765 (N_9765,N_8936,N_8536);
xor U9766 (N_9766,N_8495,N_8631);
and U9767 (N_9767,N_8652,N_8127);
and U9768 (N_9768,N_8647,N_8064);
nor U9769 (N_9769,N_8392,N_8220);
nand U9770 (N_9770,N_8436,N_8922);
nand U9771 (N_9771,N_8483,N_8512);
and U9772 (N_9772,N_8463,N_8101);
nor U9773 (N_9773,N_8119,N_8676);
or U9774 (N_9774,N_8142,N_8367);
xnor U9775 (N_9775,N_8076,N_8094);
and U9776 (N_9776,N_8675,N_8775);
nand U9777 (N_9777,N_8291,N_8361);
nand U9778 (N_9778,N_8982,N_8881);
nor U9779 (N_9779,N_8481,N_8190);
xor U9780 (N_9780,N_8503,N_8550);
and U9781 (N_9781,N_8458,N_8771);
xnor U9782 (N_9782,N_8195,N_8100);
nor U9783 (N_9783,N_8576,N_8906);
nand U9784 (N_9784,N_8852,N_8223);
or U9785 (N_9785,N_8774,N_8413);
and U9786 (N_9786,N_8082,N_8114);
or U9787 (N_9787,N_8049,N_8748);
or U9788 (N_9788,N_8167,N_8051);
nor U9789 (N_9789,N_8456,N_8814);
xor U9790 (N_9790,N_8923,N_8407);
nor U9791 (N_9791,N_8290,N_8505);
and U9792 (N_9792,N_8157,N_8532);
and U9793 (N_9793,N_8604,N_8241);
or U9794 (N_9794,N_8135,N_8679);
and U9795 (N_9795,N_8451,N_8176);
nor U9796 (N_9796,N_8594,N_8516);
nor U9797 (N_9797,N_8440,N_8397);
nor U9798 (N_9798,N_8013,N_8581);
and U9799 (N_9799,N_8232,N_8122);
or U9800 (N_9800,N_8475,N_8942);
or U9801 (N_9801,N_8399,N_8832);
or U9802 (N_9802,N_8148,N_8238);
xor U9803 (N_9803,N_8690,N_8131);
xor U9804 (N_9804,N_8258,N_8878);
xnor U9805 (N_9805,N_8091,N_8389);
or U9806 (N_9806,N_8259,N_8041);
nor U9807 (N_9807,N_8998,N_8420);
and U9808 (N_9808,N_8843,N_8567);
xnor U9809 (N_9809,N_8546,N_8091);
nand U9810 (N_9810,N_8695,N_8570);
and U9811 (N_9811,N_8507,N_8613);
or U9812 (N_9812,N_8017,N_8896);
or U9813 (N_9813,N_8384,N_8274);
nor U9814 (N_9814,N_8802,N_8491);
nand U9815 (N_9815,N_8814,N_8936);
nor U9816 (N_9816,N_8758,N_8016);
or U9817 (N_9817,N_8309,N_8981);
xor U9818 (N_9818,N_8472,N_8574);
nor U9819 (N_9819,N_8268,N_8541);
and U9820 (N_9820,N_8417,N_8849);
or U9821 (N_9821,N_8276,N_8227);
nand U9822 (N_9822,N_8210,N_8906);
nor U9823 (N_9823,N_8642,N_8557);
and U9824 (N_9824,N_8510,N_8319);
or U9825 (N_9825,N_8436,N_8924);
or U9826 (N_9826,N_8109,N_8037);
nand U9827 (N_9827,N_8320,N_8122);
xor U9828 (N_9828,N_8837,N_8219);
nor U9829 (N_9829,N_8137,N_8332);
or U9830 (N_9830,N_8675,N_8763);
or U9831 (N_9831,N_8229,N_8787);
xor U9832 (N_9832,N_8789,N_8388);
and U9833 (N_9833,N_8612,N_8964);
and U9834 (N_9834,N_8671,N_8287);
or U9835 (N_9835,N_8147,N_8675);
nor U9836 (N_9836,N_8963,N_8135);
xnor U9837 (N_9837,N_8739,N_8322);
or U9838 (N_9838,N_8815,N_8413);
and U9839 (N_9839,N_8096,N_8879);
xnor U9840 (N_9840,N_8255,N_8762);
or U9841 (N_9841,N_8853,N_8627);
and U9842 (N_9842,N_8545,N_8089);
and U9843 (N_9843,N_8822,N_8685);
nor U9844 (N_9844,N_8206,N_8872);
and U9845 (N_9845,N_8557,N_8804);
and U9846 (N_9846,N_8388,N_8404);
nand U9847 (N_9847,N_8714,N_8834);
and U9848 (N_9848,N_8198,N_8130);
and U9849 (N_9849,N_8361,N_8149);
nand U9850 (N_9850,N_8986,N_8423);
and U9851 (N_9851,N_8681,N_8380);
nor U9852 (N_9852,N_8233,N_8109);
nor U9853 (N_9853,N_8063,N_8252);
or U9854 (N_9854,N_8019,N_8515);
nand U9855 (N_9855,N_8879,N_8451);
and U9856 (N_9856,N_8138,N_8586);
nor U9857 (N_9857,N_8129,N_8514);
or U9858 (N_9858,N_8306,N_8350);
xor U9859 (N_9859,N_8201,N_8131);
or U9860 (N_9860,N_8398,N_8124);
nand U9861 (N_9861,N_8858,N_8067);
and U9862 (N_9862,N_8675,N_8799);
xnor U9863 (N_9863,N_8250,N_8544);
nand U9864 (N_9864,N_8942,N_8652);
and U9865 (N_9865,N_8803,N_8338);
or U9866 (N_9866,N_8269,N_8447);
and U9867 (N_9867,N_8089,N_8388);
xor U9868 (N_9868,N_8431,N_8142);
or U9869 (N_9869,N_8195,N_8825);
and U9870 (N_9870,N_8607,N_8283);
nand U9871 (N_9871,N_8981,N_8940);
or U9872 (N_9872,N_8150,N_8958);
nand U9873 (N_9873,N_8952,N_8873);
or U9874 (N_9874,N_8979,N_8190);
and U9875 (N_9875,N_8135,N_8255);
xor U9876 (N_9876,N_8939,N_8241);
and U9877 (N_9877,N_8878,N_8637);
nand U9878 (N_9878,N_8719,N_8520);
nor U9879 (N_9879,N_8966,N_8768);
and U9880 (N_9880,N_8071,N_8122);
or U9881 (N_9881,N_8719,N_8995);
and U9882 (N_9882,N_8962,N_8937);
nor U9883 (N_9883,N_8859,N_8409);
and U9884 (N_9884,N_8053,N_8251);
nor U9885 (N_9885,N_8237,N_8048);
xnor U9886 (N_9886,N_8444,N_8776);
and U9887 (N_9887,N_8940,N_8829);
or U9888 (N_9888,N_8114,N_8628);
nand U9889 (N_9889,N_8660,N_8577);
xor U9890 (N_9890,N_8078,N_8571);
nand U9891 (N_9891,N_8067,N_8328);
and U9892 (N_9892,N_8832,N_8064);
or U9893 (N_9893,N_8986,N_8459);
nor U9894 (N_9894,N_8528,N_8652);
and U9895 (N_9895,N_8390,N_8161);
nand U9896 (N_9896,N_8683,N_8575);
or U9897 (N_9897,N_8725,N_8734);
nand U9898 (N_9898,N_8802,N_8317);
xnor U9899 (N_9899,N_8954,N_8758);
nand U9900 (N_9900,N_8851,N_8387);
xnor U9901 (N_9901,N_8343,N_8113);
xnor U9902 (N_9902,N_8468,N_8182);
nand U9903 (N_9903,N_8541,N_8301);
nor U9904 (N_9904,N_8191,N_8682);
xnor U9905 (N_9905,N_8227,N_8140);
nand U9906 (N_9906,N_8718,N_8923);
nand U9907 (N_9907,N_8329,N_8434);
and U9908 (N_9908,N_8081,N_8904);
xor U9909 (N_9909,N_8083,N_8261);
and U9910 (N_9910,N_8534,N_8334);
xnor U9911 (N_9911,N_8718,N_8735);
xor U9912 (N_9912,N_8585,N_8341);
or U9913 (N_9913,N_8776,N_8318);
nand U9914 (N_9914,N_8099,N_8858);
nand U9915 (N_9915,N_8537,N_8088);
xnor U9916 (N_9916,N_8371,N_8757);
xnor U9917 (N_9917,N_8749,N_8155);
or U9918 (N_9918,N_8772,N_8280);
or U9919 (N_9919,N_8801,N_8295);
or U9920 (N_9920,N_8175,N_8418);
xor U9921 (N_9921,N_8244,N_8920);
or U9922 (N_9922,N_8956,N_8774);
and U9923 (N_9923,N_8313,N_8254);
and U9924 (N_9924,N_8416,N_8089);
nor U9925 (N_9925,N_8715,N_8984);
nor U9926 (N_9926,N_8798,N_8967);
nand U9927 (N_9927,N_8481,N_8755);
xnor U9928 (N_9928,N_8978,N_8390);
and U9929 (N_9929,N_8734,N_8803);
nor U9930 (N_9930,N_8121,N_8020);
xnor U9931 (N_9931,N_8053,N_8979);
or U9932 (N_9932,N_8307,N_8417);
and U9933 (N_9933,N_8376,N_8652);
nor U9934 (N_9934,N_8543,N_8399);
and U9935 (N_9935,N_8138,N_8612);
and U9936 (N_9936,N_8224,N_8804);
nor U9937 (N_9937,N_8704,N_8047);
and U9938 (N_9938,N_8718,N_8535);
and U9939 (N_9939,N_8330,N_8268);
nand U9940 (N_9940,N_8687,N_8031);
and U9941 (N_9941,N_8209,N_8540);
and U9942 (N_9942,N_8222,N_8746);
and U9943 (N_9943,N_8420,N_8953);
nand U9944 (N_9944,N_8621,N_8448);
nor U9945 (N_9945,N_8868,N_8503);
xor U9946 (N_9946,N_8889,N_8099);
nor U9947 (N_9947,N_8442,N_8397);
or U9948 (N_9948,N_8365,N_8798);
nor U9949 (N_9949,N_8263,N_8605);
nor U9950 (N_9950,N_8408,N_8774);
nand U9951 (N_9951,N_8331,N_8745);
xor U9952 (N_9952,N_8523,N_8876);
xor U9953 (N_9953,N_8975,N_8852);
or U9954 (N_9954,N_8099,N_8569);
xnor U9955 (N_9955,N_8582,N_8961);
nor U9956 (N_9956,N_8101,N_8121);
nor U9957 (N_9957,N_8426,N_8338);
nor U9958 (N_9958,N_8491,N_8118);
nand U9959 (N_9959,N_8859,N_8338);
nor U9960 (N_9960,N_8959,N_8227);
or U9961 (N_9961,N_8227,N_8967);
xor U9962 (N_9962,N_8998,N_8419);
nor U9963 (N_9963,N_8617,N_8758);
nor U9964 (N_9964,N_8279,N_8318);
and U9965 (N_9965,N_8500,N_8269);
nor U9966 (N_9966,N_8711,N_8447);
nand U9967 (N_9967,N_8760,N_8601);
nand U9968 (N_9968,N_8351,N_8589);
and U9969 (N_9969,N_8341,N_8223);
xor U9970 (N_9970,N_8032,N_8913);
nor U9971 (N_9971,N_8863,N_8300);
nand U9972 (N_9972,N_8140,N_8685);
and U9973 (N_9973,N_8142,N_8839);
xor U9974 (N_9974,N_8140,N_8231);
xor U9975 (N_9975,N_8248,N_8039);
and U9976 (N_9976,N_8332,N_8699);
xnor U9977 (N_9977,N_8751,N_8976);
xnor U9978 (N_9978,N_8536,N_8520);
nor U9979 (N_9979,N_8264,N_8155);
nand U9980 (N_9980,N_8212,N_8230);
nor U9981 (N_9981,N_8876,N_8451);
and U9982 (N_9982,N_8551,N_8986);
or U9983 (N_9983,N_8356,N_8663);
nand U9984 (N_9984,N_8273,N_8530);
nand U9985 (N_9985,N_8670,N_8235);
or U9986 (N_9986,N_8903,N_8709);
or U9987 (N_9987,N_8197,N_8981);
and U9988 (N_9988,N_8673,N_8392);
xnor U9989 (N_9989,N_8010,N_8262);
or U9990 (N_9990,N_8148,N_8668);
nand U9991 (N_9991,N_8809,N_8843);
xnor U9992 (N_9992,N_8673,N_8658);
or U9993 (N_9993,N_8476,N_8559);
or U9994 (N_9994,N_8280,N_8096);
xor U9995 (N_9995,N_8710,N_8022);
nor U9996 (N_9996,N_8911,N_8023);
or U9997 (N_9997,N_8288,N_8201);
nand U9998 (N_9998,N_8216,N_8692);
or U9999 (N_9999,N_8938,N_8128);
or U10000 (N_10000,N_9106,N_9221);
or U10001 (N_10001,N_9249,N_9630);
nor U10002 (N_10002,N_9827,N_9430);
nor U10003 (N_10003,N_9929,N_9072);
nor U10004 (N_10004,N_9085,N_9327);
nor U10005 (N_10005,N_9338,N_9444);
or U10006 (N_10006,N_9992,N_9349);
xnor U10007 (N_10007,N_9801,N_9450);
nor U10008 (N_10008,N_9582,N_9042);
xnor U10009 (N_10009,N_9966,N_9626);
nand U10010 (N_10010,N_9887,N_9276);
xor U10011 (N_10011,N_9086,N_9096);
xnor U10012 (N_10012,N_9885,N_9556);
nand U10013 (N_10013,N_9071,N_9238);
xnor U10014 (N_10014,N_9942,N_9167);
nand U10015 (N_10015,N_9655,N_9390);
xor U10016 (N_10016,N_9633,N_9273);
xor U10017 (N_10017,N_9542,N_9977);
or U10018 (N_10018,N_9604,N_9255);
nand U10019 (N_10019,N_9863,N_9596);
nand U10020 (N_10020,N_9839,N_9890);
xor U10021 (N_10021,N_9646,N_9415);
or U10022 (N_10022,N_9373,N_9480);
nor U10023 (N_10023,N_9826,N_9332);
xor U10024 (N_10024,N_9687,N_9728);
nor U10025 (N_10025,N_9980,N_9590);
nand U10026 (N_10026,N_9132,N_9841);
xor U10027 (N_10027,N_9207,N_9179);
nand U10028 (N_10028,N_9000,N_9139);
and U10029 (N_10029,N_9499,N_9800);
nand U10030 (N_10030,N_9472,N_9173);
nor U10031 (N_10031,N_9615,N_9700);
and U10032 (N_10032,N_9384,N_9206);
nor U10033 (N_10033,N_9934,N_9032);
or U10034 (N_10034,N_9391,N_9171);
nand U10035 (N_10035,N_9549,N_9376);
and U10036 (N_10036,N_9235,N_9906);
or U10037 (N_10037,N_9679,N_9849);
and U10038 (N_10038,N_9583,N_9240);
xnor U10039 (N_10039,N_9363,N_9857);
nand U10040 (N_10040,N_9256,N_9599);
nand U10041 (N_10041,N_9939,N_9287);
and U10042 (N_10042,N_9355,N_9014);
xor U10043 (N_10043,N_9816,N_9600);
nor U10044 (N_10044,N_9814,N_9927);
or U10045 (N_10045,N_9069,N_9214);
nand U10046 (N_10046,N_9413,N_9260);
nor U10047 (N_10047,N_9199,N_9924);
nand U10048 (N_10048,N_9794,N_9922);
nand U10049 (N_10049,N_9151,N_9428);
and U10050 (N_10050,N_9227,N_9952);
and U10051 (N_10051,N_9840,N_9452);
and U10052 (N_10052,N_9813,N_9406);
nor U10053 (N_10053,N_9719,N_9866);
or U10054 (N_10054,N_9130,N_9546);
nand U10055 (N_10055,N_9311,N_9717);
or U10056 (N_10056,N_9304,N_9682);
xnor U10057 (N_10057,N_9325,N_9523);
and U10058 (N_10058,N_9222,N_9065);
nand U10059 (N_10059,N_9121,N_9671);
or U10060 (N_10060,N_9440,N_9754);
nand U10061 (N_10061,N_9254,N_9974);
and U10062 (N_10062,N_9476,N_9050);
nand U10063 (N_10063,N_9765,N_9577);
and U10064 (N_10064,N_9458,N_9744);
nor U10065 (N_10065,N_9243,N_9821);
or U10066 (N_10066,N_9062,N_9788);
xor U10067 (N_10067,N_9503,N_9572);
or U10068 (N_10068,N_9555,N_9131);
xnor U10069 (N_10069,N_9028,N_9704);
xnor U10070 (N_10070,N_9904,N_9531);
nor U10071 (N_10071,N_9228,N_9947);
or U10072 (N_10072,N_9166,N_9519);
nand U10073 (N_10073,N_9424,N_9478);
nand U10074 (N_10074,N_9954,N_9150);
nor U10075 (N_10075,N_9508,N_9869);
xor U10076 (N_10076,N_9019,N_9799);
or U10077 (N_10077,N_9545,N_9250);
and U10078 (N_10078,N_9898,N_9477);
nor U10079 (N_10079,N_9183,N_9160);
nand U10080 (N_10080,N_9521,N_9773);
xor U10081 (N_10081,N_9181,N_9443);
nor U10082 (N_10082,N_9786,N_9012);
and U10083 (N_10083,N_9536,N_9058);
xnor U10084 (N_10084,N_9372,N_9892);
nor U10085 (N_10085,N_9627,N_9195);
nor U10086 (N_10086,N_9093,N_9446);
nor U10087 (N_10087,N_9532,N_9436);
or U10088 (N_10088,N_9259,N_9475);
xnor U10089 (N_10089,N_9855,N_9219);
nor U10090 (N_10090,N_9081,N_9798);
or U10091 (N_10091,N_9730,N_9516);
nor U10092 (N_10092,N_9133,N_9220);
and U10093 (N_10093,N_9334,N_9039);
nand U10094 (N_10094,N_9852,N_9561);
xnor U10095 (N_10095,N_9479,N_9518);
or U10096 (N_10096,N_9959,N_9422);
or U10097 (N_10097,N_9917,N_9873);
or U10098 (N_10098,N_9076,N_9336);
or U10099 (N_10099,N_9982,N_9239);
and U10100 (N_10100,N_9226,N_9994);
and U10101 (N_10101,N_9291,N_9122);
nand U10102 (N_10102,N_9416,N_9107);
nand U10103 (N_10103,N_9120,N_9374);
xor U10104 (N_10104,N_9500,N_9252);
nor U10105 (N_10105,N_9016,N_9738);
and U10106 (N_10106,N_9568,N_9379);
xnor U10107 (N_10107,N_9729,N_9027);
nand U10108 (N_10108,N_9022,N_9691);
or U10109 (N_10109,N_9741,N_9817);
or U10110 (N_10110,N_9760,N_9234);
nand U10111 (N_10111,N_9958,N_9735);
and U10112 (N_10112,N_9676,N_9914);
xor U10113 (N_10113,N_9084,N_9835);
or U10114 (N_10114,N_9736,N_9739);
or U10115 (N_10115,N_9533,N_9049);
xor U10116 (N_10116,N_9411,N_9514);
or U10117 (N_10117,N_9812,N_9956);
or U10118 (N_10118,N_9398,N_9848);
and U10119 (N_10119,N_9547,N_9108);
nand U10120 (N_10120,N_9455,N_9486);
or U10121 (N_10121,N_9811,N_9818);
and U10122 (N_10122,N_9110,N_9074);
and U10123 (N_10123,N_9351,N_9781);
or U10124 (N_10124,N_9025,N_9520);
nor U10125 (N_10125,N_9565,N_9041);
nor U10126 (N_10126,N_9292,N_9169);
nand U10127 (N_10127,N_9787,N_9511);
nor U10128 (N_10128,N_9524,N_9156);
or U10129 (N_10129,N_9347,N_9483);
or U10130 (N_10130,N_9116,N_9253);
nor U10131 (N_10131,N_9861,N_9688);
or U10132 (N_10132,N_9896,N_9441);
xnor U10133 (N_10133,N_9783,N_9002);
nor U10134 (N_10134,N_9434,N_9283);
and U10135 (N_10135,N_9468,N_9925);
or U10136 (N_10136,N_9641,N_9282);
or U10137 (N_10137,N_9916,N_9190);
and U10138 (N_10138,N_9129,N_9265);
and U10139 (N_10139,N_9609,N_9187);
nand U10140 (N_10140,N_9680,N_9601);
or U10141 (N_10141,N_9987,N_9034);
xor U10142 (N_10142,N_9011,N_9136);
nor U10143 (N_10143,N_9497,N_9236);
nor U10144 (N_10144,N_9632,N_9098);
nor U10145 (N_10145,N_9782,N_9973);
nand U10146 (N_10146,N_9057,N_9362);
and U10147 (N_10147,N_9340,N_9838);
xor U10148 (N_10148,N_9822,N_9715);
nor U10149 (N_10149,N_9141,N_9385);
or U10150 (N_10150,N_9319,N_9460);
xnor U10151 (N_10151,N_9926,N_9820);
or U10152 (N_10152,N_9261,N_9949);
nand U10153 (N_10153,N_9033,N_9749);
nand U10154 (N_10154,N_9767,N_9957);
and U10155 (N_10155,N_9123,N_9356);
xor U10156 (N_10156,N_9603,N_9854);
nand U10157 (N_10157,N_9637,N_9540);
xnor U10158 (N_10158,N_9289,N_9078);
or U10159 (N_10159,N_9874,N_9482);
nand U10160 (N_10160,N_9296,N_9274);
nand U10161 (N_10161,N_9496,N_9563);
nand U10162 (N_10162,N_9030,N_9449);
nor U10163 (N_10163,N_9277,N_9907);
xor U10164 (N_10164,N_9491,N_9879);
nand U10165 (N_10165,N_9505,N_9017);
xor U10166 (N_10166,N_9438,N_9698);
nor U10167 (N_10167,N_9001,N_9029);
or U10168 (N_10168,N_9103,N_9899);
nor U10169 (N_10169,N_9764,N_9264);
nand U10170 (N_10170,N_9803,N_9650);
and U10171 (N_10171,N_9119,N_9357);
nand U10172 (N_10172,N_9408,N_9114);
or U10173 (N_10173,N_9462,N_9795);
xor U10174 (N_10174,N_9726,N_9512);
or U10175 (N_10175,N_9614,N_9489);
nand U10176 (N_10176,N_9456,N_9653);
or U10177 (N_10177,N_9375,N_9672);
nor U10178 (N_10178,N_9968,N_9109);
nor U10179 (N_10179,N_9617,N_9059);
nand U10180 (N_10180,N_9067,N_9860);
or U10181 (N_10181,N_9297,N_9286);
xor U10182 (N_10182,N_9381,N_9364);
nand U10183 (N_10183,N_9153,N_9999);
nor U10184 (N_10184,N_9471,N_9716);
xor U10185 (N_10185,N_9570,N_9908);
nand U10186 (N_10186,N_9213,N_9905);
and U10187 (N_10187,N_9046,N_9113);
or U10188 (N_10188,N_9608,N_9643);
nor U10189 (N_10189,N_9426,N_9910);
or U10190 (N_10190,N_9223,N_9117);
nor U10191 (N_10191,N_9544,N_9099);
nor U10192 (N_10192,N_9230,N_9891);
and U10193 (N_10193,N_9248,N_9401);
or U10194 (N_10194,N_9659,N_9553);
or U10195 (N_10195,N_9089,N_9941);
xor U10196 (N_10196,N_9125,N_9163);
or U10197 (N_10197,N_9806,N_9526);
and U10198 (N_10198,N_9184,N_9453);
nand U10199 (N_10199,N_9063,N_9023);
and U10200 (N_10200,N_9083,N_9955);
nand U10201 (N_10201,N_9048,N_9769);
or U10202 (N_10202,N_9314,N_9776);
xor U10203 (N_10203,N_9707,N_9647);
xnor U10204 (N_10204,N_9872,N_9802);
xnor U10205 (N_10205,N_9578,N_9960);
xnor U10206 (N_10206,N_9146,N_9101);
or U10207 (N_10207,N_9618,N_9395);
and U10208 (N_10208,N_9901,N_9329);
nand U10209 (N_10209,N_9135,N_9881);
nand U10210 (N_10210,N_9481,N_9115);
and U10211 (N_10211,N_9305,N_9620);
nor U10212 (N_10212,N_9168,N_9851);
or U10213 (N_10213,N_9597,N_9284);
and U10214 (N_10214,N_9779,N_9231);
and U10215 (N_10215,N_9470,N_9387);
and U10216 (N_10216,N_9902,N_9918);
nand U10217 (N_10217,N_9366,N_9288);
nand U10218 (N_10218,N_9148,N_9403);
nor U10219 (N_10219,N_9341,N_9112);
nor U10220 (N_10220,N_9268,N_9429);
xnor U10221 (N_10221,N_9111,N_9492);
or U10222 (N_10222,N_9320,N_9535);
nor U10223 (N_10223,N_9409,N_9703);
xnor U10224 (N_10224,N_9212,N_9061);
and U10225 (N_10225,N_9457,N_9003);
nor U10226 (N_10226,N_9128,N_9124);
and U10227 (N_10227,N_9420,N_9105);
nand U10228 (N_10228,N_9930,N_9138);
nor U10229 (N_10229,N_9990,N_9417);
xnor U10230 (N_10230,N_9574,N_9877);
and U10231 (N_10231,N_9548,N_9629);
xor U10232 (N_10232,N_9439,N_9746);
or U10233 (N_10233,N_9689,N_9473);
nand U10234 (N_10234,N_9656,N_9678);
and U10235 (N_10235,N_9613,N_9701);
nor U10236 (N_10236,N_9290,N_9853);
and U10237 (N_10237,N_9928,N_9339);
nor U10238 (N_10238,N_9217,N_9762);
nand U10239 (N_10239,N_9090,N_9580);
or U10240 (N_10240,N_9986,N_9971);
xnor U10241 (N_10241,N_9300,N_9616);
and U10242 (N_10242,N_9984,N_9751);
or U10243 (N_10243,N_9876,N_9433);
xnor U10244 (N_10244,N_9865,N_9175);
nand U10245 (N_10245,N_9077,N_9964);
xor U10246 (N_10246,N_9976,N_9780);
xor U10247 (N_10247,N_9038,N_9224);
or U10248 (N_10248,N_9402,N_9307);
nand U10249 (N_10249,N_9504,N_9766);
and U10250 (N_10250,N_9165,N_9770);
nand U10251 (N_10251,N_9789,N_9963);
nor U10252 (N_10252,N_9658,N_9080);
nor U10253 (N_10253,N_9400,N_9317);
nor U10254 (N_10254,N_9419,N_9186);
xnor U10255 (N_10255,N_9414,N_9713);
and U10256 (N_10256,N_9652,N_9137);
and U10257 (N_10257,N_9075,N_9389);
or U10258 (N_10258,N_9588,N_9797);
nand U10259 (N_10259,N_9864,N_9975);
xor U10260 (N_10260,N_9771,N_9775);
or U10261 (N_10261,N_9528,N_9935);
nor U10262 (N_10262,N_9936,N_9353);
nor U10263 (N_10263,N_9361,N_9088);
nand U10264 (N_10264,N_9344,N_9293);
nor U10265 (N_10265,N_9551,N_9104);
xnor U10266 (N_10266,N_9829,N_9367);
nand U10267 (N_10267,N_9383,N_9335);
and U10268 (N_10268,N_9525,N_9875);
xor U10269 (N_10269,N_9645,N_9270);
or U10270 (N_10270,N_9591,N_9053);
and U10271 (N_10271,N_9534,N_9092);
or U10272 (N_10272,N_9352,N_9303);
nor U10273 (N_10273,N_9758,N_9066);
nor U10274 (N_10274,N_9218,N_9639);
xor U10275 (N_10275,N_9573,N_9785);
xnor U10276 (N_10276,N_9144,N_9040);
and U10277 (N_10277,N_9837,N_9127);
and U10278 (N_10278,N_9244,N_9602);
or U10279 (N_10279,N_9378,N_9581);
xnor U10280 (N_10280,N_9451,N_9623);
nor U10281 (N_10281,N_9233,N_9777);
nand U10282 (N_10282,N_9560,N_9878);
or U10283 (N_10283,N_9809,N_9278);
nand U10284 (N_10284,N_9683,N_9669);
xor U10285 (N_10285,N_9251,N_9463);
or U10286 (N_10286,N_9097,N_9624);
and U10287 (N_10287,N_9681,N_9094);
nand U10288 (N_10288,N_9229,N_9550);
nand U10289 (N_10289,N_9943,N_9189);
nand U10290 (N_10290,N_9972,N_9162);
and U10291 (N_10291,N_9507,N_9194);
and U10292 (N_10292,N_9043,N_9699);
xnor U10293 (N_10293,N_9421,N_9281);
and U10294 (N_10294,N_9807,N_9258);
nor U10295 (N_10295,N_9170,N_9467);
and U10296 (N_10296,N_9407,N_9537);
and U10297 (N_10297,N_9692,N_9668);
nand U10298 (N_10298,N_9981,N_9350);
and U10299 (N_10299,N_9844,N_9257);
and U10300 (N_10300,N_9161,N_9557);
and U10301 (N_10301,N_9983,N_9642);
nand U10302 (N_10302,N_9948,N_9950);
nor U10303 (N_10303,N_9628,N_9267);
or U10304 (N_10304,N_9313,N_9660);
xnor U10305 (N_10305,N_9324,N_9466);
or U10306 (N_10306,N_9510,N_9784);
nor U10307 (N_10307,N_9280,N_9894);
nor U10308 (N_10308,N_9640,N_9348);
nor U10309 (N_10309,N_9587,N_9203);
nor U10310 (N_10310,N_9010,N_9989);
nand U10311 (N_10311,N_9909,N_9454);
and U10312 (N_10312,N_9308,N_9667);
or U10313 (N_10313,N_9399,N_9006);
xor U10314 (N_10314,N_9498,N_9102);
nand U10315 (N_10315,N_9567,N_9502);
nor U10316 (N_10316,N_9586,N_9845);
nand U10317 (N_10317,N_9513,N_9595);
xor U10318 (N_10318,N_9036,N_9832);
xnor U10319 (N_10319,N_9388,N_9673);
and U10320 (N_10320,N_9299,N_9154);
nand U10321 (N_10321,N_9196,N_9805);
nor U10322 (N_10322,N_9953,N_9118);
and U10323 (N_10323,N_9810,N_9246);
xnor U10324 (N_10324,N_9843,N_9913);
and U10325 (N_10325,N_9649,N_9740);
nor U10326 (N_10326,N_9790,N_9377);
and U10327 (N_10327,N_9008,N_9490);
nand U10328 (N_10328,N_9793,N_9020);
or U10329 (N_10329,N_9263,N_9761);
or U10330 (N_10330,N_9721,N_9833);
nor U10331 (N_10331,N_9911,N_9897);
or U10332 (N_10332,N_9714,N_9745);
nand U10333 (N_10333,N_9487,N_9657);
xor U10334 (N_10334,N_9204,N_9082);
nor U10335 (N_10335,N_9285,N_9825);
and U10336 (N_10336,N_9529,N_9828);
or U10337 (N_10337,N_9705,N_9365);
and U10338 (N_10338,N_9198,N_9607);
nor U10339 (N_10339,N_9394,N_9711);
and U10340 (N_10340,N_9051,N_9946);
xor U10341 (N_10341,N_9622,N_9174);
and U10342 (N_10342,N_9882,N_9900);
or U10343 (N_10343,N_9005,N_9944);
nor U10344 (N_10344,N_9396,N_9970);
or U10345 (N_10345,N_9585,N_9675);
xor U10346 (N_10346,N_9734,N_9371);
nand U10347 (N_10347,N_9178,N_9575);
or U10348 (N_10348,N_9100,N_9185);
nand U10349 (N_10349,N_9392,N_9710);
and U10350 (N_10350,N_9893,N_9933);
nor U10351 (N_10351,N_9405,N_9743);
nor U10352 (N_10352,N_9611,N_9895);
nand U10353 (N_10353,N_9004,N_9778);
xnor U10354 (N_10354,N_9464,N_9919);
nand U10355 (N_10355,N_9862,N_9662);
xor U10356 (N_10356,N_9142,N_9880);
xor U10357 (N_10357,N_9024,N_9326);
or U10358 (N_10358,N_9241,N_9459);
nand U10359 (N_10359,N_9559,N_9988);
and U10360 (N_10360,N_9663,N_9474);
nand U10361 (N_10361,N_9359,N_9275);
nand U10362 (N_10362,N_9301,N_9808);
or U10363 (N_10363,N_9044,N_9562);
and U10364 (N_10364,N_9527,N_9007);
nor U10365 (N_10365,N_9846,N_9404);
nand U10366 (N_10366,N_9380,N_9830);
nand U10367 (N_10367,N_9593,N_9026);
or U10368 (N_10368,N_9665,N_9923);
or U10369 (N_10369,N_9576,N_9501);
nor U10370 (N_10370,N_9702,N_9644);
or U10371 (N_10371,N_9859,N_9410);
nand U10372 (N_10372,N_9469,N_9079);
nand U10373 (N_10373,N_9768,N_9262);
nand U10374 (N_10374,N_9884,N_9727);
or U10375 (N_10375,N_9427,N_9370);
nand U10376 (N_10376,N_9200,N_9965);
nand U10377 (N_10377,N_9343,N_9091);
nand U10378 (N_10378,N_9696,N_9494);
nor U10379 (N_10379,N_9791,N_9149);
and U10380 (N_10380,N_9211,N_9279);
and U10381 (N_10381,N_9152,N_9517);
and U10382 (N_10382,N_9712,N_9346);
or U10383 (N_10383,N_9932,N_9823);
nand U10384 (N_10384,N_9579,N_9636);
or U10385 (N_10385,N_9354,N_9073);
xnor U10386 (N_10386,N_9995,N_9134);
nor U10387 (N_10387,N_9232,N_9312);
nand U10388 (N_10388,N_9054,N_9316);
or U10389 (N_10389,N_9635,N_9978);
or U10390 (N_10390,N_9158,N_9328);
or U10391 (N_10391,N_9208,N_9055);
and U10392 (N_10392,N_9318,N_9831);
nand U10393 (N_10393,N_9541,N_9515);
and U10394 (N_10394,N_9940,N_9306);
nand U10395 (N_10395,N_9035,N_9192);
nand U10396 (N_10396,N_9386,N_9598);
xnor U10397 (N_10397,N_9552,N_9856);
and U10398 (N_10398,N_9045,N_9661);
xor U10399 (N_10399,N_9566,N_9432);
and U10400 (N_10400,N_9834,N_9868);
nand U10401 (N_10401,N_9605,N_9677);
nand U10402 (N_10402,N_9216,N_9755);
xnor U10403 (N_10403,N_9397,N_9493);
and U10404 (N_10404,N_9706,N_9322);
nand U10405 (N_10405,N_9920,N_9883);
nor U10406 (N_10406,N_9143,N_9488);
or U10407 (N_10407,N_9435,N_9979);
and U10408 (N_10408,N_9564,N_9245);
xnor U10409 (N_10409,N_9967,N_9210);
nor U10410 (N_10410,N_9393,N_9188);
nand U10411 (N_10411,N_9418,N_9495);
nor U10412 (N_10412,N_9589,N_9748);
or U10413 (N_10413,N_9266,N_9792);
or U10414 (N_10414,N_9962,N_9804);
xor U10415 (N_10415,N_9140,N_9724);
xnor U10416 (N_10416,N_9323,N_9201);
nand U10417 (N_10417,N_9619,N_9651);
xor U10418 (N_10418,N_9842,N_9670);
or U10419 (N_10419,N_9180,N_9506);
and U10420 (N_10420,N_9197,N_9205);
nor U10421 (N_10421,N_9737,N_9159);
and U10422 (N_10422,N_9886,N_9871);
xor U10423 (N_10423,N_9757,N_9269);
or U10424 (N_10424,N_9772,N_9068);
nor U10425 (N_10425,N_9725,N_9903);
xor U10426 (N_10426,N_9437,N_9530);
nand U10427 (N_10427,N_9177,N_9484);
xor U10428 (N_10428,N_9722,N_9945);
and U10429 (N_10429,N_9985,N_9912);
nor U10430 (N_10430,N_9708,N_9732);
and U10431 (N_10431,N_9621,N_9461);
nor U10432 (N_10432,N_9690,N_9961);
nand U10433 (N_10433,N_9191,N_9796);
and U10434 (N_10434,N_9242,N_9310);
nor U10435 (N_10435,N_9018,N_9193);
and U10436 (N_10436,N_9485,N_9571);
nand U10437 (N_10437,N_9686,N_9358);
xor U10438 (N_10438,N_9164,N_9723);
nor U10439 (N_10439,N_9951,N_9638);
nor U10440 (N_10440,N_9052,N_9237);
or U10441 (N_10441,N_9931,N_9095);
xnor U10442 (N_10442,N_9709,N_9342);
nor U10443 (N_10443,N_9448,N_9666);
xnor U10444 (N_10444,N_9697,N_9664);
nor U10445 (N_10445,N_9858,N_9147);
nor U10446 (N_10446,N_9015,N_9991);
xnor U10447 (N_10447,N_9176,N_9009);
nor U10448 (N_10448,N_9447,N_9298);
and U10449 (N_10449,N_9774,N_9921);
nor U10450 (N_10450,N_9369,N_9847);
and U10451 (N_10451,N_9215,N_9368);
nand U10452 (N_10452,N_9333,N_9694);
or U10453 (N_10453,N_9382,N_9047);
and U10454 (N_10454,N_9756,N_9888);
xnor U10455 (N_10455,N_9742,N_9315);
nand U10456 (N_10456,N_9360,N_9202);
and U10457 (N_10457,N_9425,N_9996);
and U10458 (N_10458,N_9445,N_9558);
and U10459 (N_10459,N_9674,N_9612);
xnor U10460 (N_10460,N_9272,N_9543);
and U10461 (N_10461,N_9731,N_9993);
or U10462 (N_10462,N_9969,N_9309);
and U10463 (N_10463,N_9606,N_9412);
nand U10464 (N_10464,N_9209,N_9431);
nand U10465 (N_10465,N_9836,N_9584);
and U10466 (N_10466,N_9126,N_9302);
or U10467 (N_10467,N_9155,N_9594);
and U10468 (N_10468,N_9330,N_9064);
nor U10469 (N_10469,N_9815,N_9938);
or U10470 (N_10470,N_9013,N_9648);
xor U10471 (N_10471,N_9031,N_9695);
and U10472 (N_10472,N_9592,N_9625);
xor U10473 (N_10473,N_9247,N_9539);
nor U10474 (N_10474,N_9733,N_9295);
and U10475 (N_10475,N_9634,N_9056);
or U10476 (N_10476,N_9752,N_9747);
or U10477 (N_10477,N_9509,N_9654);
nor U10478 (N_10478,N_9824,N_9750);
nand U10479 (N_10479,N_9465,N_9145);
nor U10480 (N_10480,N_9331,N_9442);
and U10481 (N_10481,N_9522,N_9819);
nor U10482 (N_10482,N_9423,N_9021);
or U10483 (N_10483,N_9569,N_9345);
xnor U10484 (N_10484,N_9867,N_9937);
xnor U10485 (N_10485,N_9610,N_9294);
xor U10486 (N_10486,N_9070,N_9182);
and U10487 (N_10487,N_9087,N_9172);
xnor U10488 (N_10488,N_9631,N_9889);
or U10489 (N_10489,N_9915,N_9720);
and U10490 (N_10490,N_9870,N_9037);
nor U10491 (N_10491,N_9753,N_9718);
and U10492 (N_10492,N_9225,N_9850);
nand U10493 (N_10493,N_9759,N_9554);
nand U10494 (N_10494,N_9271,N_9321);
or U10495 (N_10495,N_9997,N_9693);
xnor U10496 (N_10496,N_9685,N_9763);
and U10497 (N_10497,N_9337,N_9684);
nand U10498 (N_10498,N_9538,N_9998);
or U10499 (N_10499,N_9157,N_9060);
xnor U10500 (N_10500,N_9100,N_9179);
or U10501 (N_10501,N_9076,N_9577);
and U10502 (N_10502,N_9098,N_9604);
and U10503 (N_10503,N_9950,N_9063);
xnor U10504 (N_10504,N_9054,N_9272);
and U10505 (N_10505,N_9853,N_9847);
xnor U10506 (N_10506,N_9856,N_9070);
xor U10507 (N_10507,N_9298,N_9784);
nand U10508 (N_10508,N_9154,N_9530);
or U10509 (N_10509,N_9500,N_9874);
xor U10510 (N_10510,N_9083,N_9356);
and U10511 (N_10511,N_9926,N_9502);
or U10512 (N_10512,N_9728,N_9962);
and U10513 (N_10513,N_9028,N_9632);
nor U10514 (N_10514,N_9998,N_9258);
nor U10515 (N_10515,N_9528,N_9370);
nor U10516 (N_10516,N_9976,N_9982);
and U10517 (N_10517,N_9348,N_9785);
nor U10518 (N_10518,N_9129,N_9957);
nor U10519 (N_10519,N_9655,N_9187);
xnor U10520 (N_10520,N_9946,N_9198);
or U10521 (N_10521,N_9195,N_9920);
xor U10522 (N_10522,N_9773,N_9056);
and U10523 (N_10523,N_9743,N_9395);
and U10524 (N_10524,N_9224,N_9431);
nand U10525 (N_10525,N_9778,N_9157);
xor U10526 (N_10526,N_9517,N_9146);
nor U10527 (N_10527,N_9629,N_9448);
or U10528 (N_10528,N_9574,N_9044);
or U10529 (N_10529,N_9889,N_9425);
xnor U10530 (N_10530,N_9198,N_9193);
and U10531 (N_10531,N_9682,N_9578);
nor U10532 (N_10532,N_9893,N_9311);
and U10533 (N_10533,N_9947,N_9726);
nand U10534 (N_10534,N_9852,N_9331);
and U10535 (N_10535,N_9893,N_9285);
and U10536 (N_10536,N_9142,N_9561);
xnor U10537 (N_10537,N_9207,N_9216);
xor U10538 (N_10538,N_9278,N_9037);
nor U10539 (N_10539,N_9224,N_9142);
or U10540 (N_10540,N_9034,N_9493);
nor U10541 (N_10541,N_9597,N_9836);
and U10542 (N_10542,N_9060,N_9615);
xnor U10543 (N_10543,N_9256,N_9810);
xor U10544 (N_10544,N_9858,N_9055);
or U10545 (N_10545,N_9789,N_9340);
nand U10546 (N_10546,N_9480,N_9789);
xor U10547 (N_10547,N_9093,N_9533);
nand U10548 (N_10548,N_9675,N_9732);
and U10549 (N_10549,N_9831,N_9310);
xor U10550 (N_10550,N_9025,N_9146);
and U10551 (N_10551,N_9028,N_9667);
and U10552 (N_10552,N_9764,N_9219);
nand U10553 (N_10553,N_9336,N_9784);
and U10554 (N_10554,N_9275,N_9805);
nor U10555 (N_10555,N_9783,N_9882);
nor U10556 (N_10556,N_9737,N_9283);
or U10557 (N_10557,N_9042,N_9426);
nor U10558 (N_10558,N_9176,N_9143);
nand U10559 (N_10559,N_9136,N_9629);
nand U10560 (N_10560,N_9464,N_9012);
nor U10561 (N_10561,N_9984,N_9481);
and U10562 (N_10562,N_9319,N_9980);
nor U10563 (N_10563,N_9934,N_9978);
or U10564 (N_10564,N_9486,N_9974);
nand U10565 (N_10565,N_9569,N_9250);
nand U10566 (N_10566,N_9890,N_9624);
nand U10567 (N_10567,N_9100,N_9192);
or U10568 (N_10568,N_9591,N_9674);
nand U10569 (N_10569,N_9019,N_9785);
or U10570 (N_10570,N_9562,N_9371);
xnor U10571 (N_10571,N_9380,N_9483);
or U10572 (N_10572,N_9996,N_9214);
or U10573 (N_10573,N_9229,N_9978);
xor U10574 (N_10574,N_9368,N_9245);
or U10575 (N_10575,N_9853,N_9916);
nand U10576 (N_10576,N_9012,N_9103);
nand U10577 (N_10577,N_9737,N_9161);
or U10578 (N_10578,N_9961,N_9964);
or U10579 (N_10579,N_9484,N_9999);
nand U10580 (N_10580,N_9012,N_9235);
nor U10581 (N_10581,N_9870,N_9658);
nor U10582 (N_10582,N_9201,N_9026);
or U10583 (N_10583,N_9897,N_9172);
and U10584 (N_10584,N_9754,N_9240);
nor U10585 (N_10585,N_9910,N_9846);
nor U10586 (N_10586,N_9025,N_9888);
xnor U10587 (N_10587,N_9587,N_9921);
nor U10588 (N_10588,N_9126,N_9328);
nand U10589 (N_10589,N_9958,N_9585);
nor U10590 (N_10590,N_9878,N_9748);
and U10591 (N_10591,N_9246,N_9376);
and U10592 (N_10592,N_9031,N_9067);
nor U10593 (N_10593,N_9712,N_9644);
and U10594 (N_10594,N_9038,N_9192);
or U10595 (N_10595,N_9656,N_9282);
xor U10596 (N_10596,N_9122,N_9247);
nand U10597 (N_10597,N_9238,N_9652);
and U10598 (N_10598,N_9216,N_9312);
nand U10599 (N_10599,N_9289,N_9820);
nand U10600 (N_10600,N_9024,N_9034);
nor U10601 (N_10601,N_9263,N_9714);
nand U10602 (N_10602,N_9221,N_9215);
and U10603 (N_10603,N_9047,N_9731);
xnor U10604 (N_10604,N_9958,N_9906);
nand U10605 (N_10605,N_9216,N_9359);
nor U10606 (N_10606,N_9127,N_9193);
and U10607 (N_10607,N_9700,N_9663);
xnor U10608 (N_10608,N_9931,N_9752);
nor U10609 (N_10609,N_9469,N_9686);
nor U10610 (N_10610,N_9053,N_9060);
nor U10611 (N_10611,N_9245,N_9025);
or U10612 (N_10612,N_9229,N_9468);
xnor U10613 (N_10613,N_9234,N_9119);
and U10614 (N_10614,N_9314,N_9680);
or U10615 (N_10615,N_9306,N_9741);
xor U10616 (N_10616,N_9105,N_9522);
and U10617 (N_10617,N_9855,N_9381);
nor U10618 (N_10618,N_9060,N_9921);
and U10619 (N_10619,N_9743,N_9945);
and U10620 (N_10620,N_9128,N_9352);
nor U10621 (N_10621,N_9469,N_9832);
or U10622 (N_10622,N_9466,N_9725);
xnor U10623 (N_10623,N_9796,N_9824);
nand U10624 (N_10624,N_9605,N_9600);
nand U10625 (N_10625,N_9349,N_9270);
xor U10626 (N_10626,N_9176,N_9031);
xor U10627 (N_10627,N_9881,N_9553);
nand U10628 (N_10628,N_9817,N_9070);
xor U10629 (N_10629,N_9331,N_9168);
xnor U10630 (N_10630,N_9571,N_9104);
or U10631 (N_10631,N_9753,N_9527);
or U10632 (N_10632,N_9050,N_9542);
xor U10633 (N_10633,N_9698,N_9585);
xnor U10634 (N_10634,N_9458,N_9541);
nand U10635 (N_10635,N_9623,N_9791);
nand U10636 (N_10636,N_9303,N_9253);
xnor U10637 (N_10637,N_9065,N_9770);
and U10638 (N_10638,N_9876,N_9709);
nand U10639 (N_10639,N_9990,N_9652);
nand U10640 (N_10640,N_9532,N_9437);
or U10641 (N_10641,N_9615,N_9703);
and U10642 (N_10642,N_9675,N_9912);
xnor U10643 (N_10643,N_9678,N_9566);
xnor U10644 (N_10644,N_9069,N_9745);
xnor U10645 (N_10645,N_9308,N_9201);
xnor U10646 (N_10646,N_9453,N_9167);
or U10647 (N_10647,N_9003,N_9142);
nor U10648 (N_10648,N_9794,N_9242);
nand U10649 (N_10649,N_9968,N_9072);
nor U10650 (N_10650,N_9318,N_9092);
and U10651 (N_10651,N_9667,N_9097);
and U10652 (N_10652,N_9804,N_9874);
and U10653 (N_10653,N_9918,N_9787);
xnor U10654 (N_10654,N_9638,N_9821);
and U10655 (N_10655,N_9097,N_9684);
and U10656 (N_10656,N_9185,N_9919);
nor U10657 (N_10657,N_9272,N_9732);
and U10658 (N_10658,N_9288,N_9323);
or U10659 (N_10659,N_9958,N_9504);
or U10660 (N_10660,N_9590,N_9297);
nor U10661 (N_10661,N_9916,N_9646);
nand U10662 (N_10662,N_9029,N_9759);
nor U10663 (N_10663,N_9292,N_9597);
and U10664 (N_10664,N_9883,N_9304);
and U10665 (N_10665,N_9017,N_9490);
or U10666 (N_10666,N_9787,N_9380);
xnor U10667 (N_10667,N_9021,N_9851);
xor U10668 (N_10668,N_9530,N_9554);
and U10669 (N_10669,N_9677,N_9069);
nor U10670 (N_10670,N_9432,N_9141);
and U10671 (N_10671,N_9275,N_9169);
or U10672 (N_10672,N_9274,N_9523);
nand U10673 (N_10673,N_9743,N_9221);
nand U10674 (N_10674,N_9156,N_9890);
or U10675 (N_10675,N_9331,N_9552);
and U10676 (N_10676,N_9210,N_9042);
nor U10677 (N_10677,N_9233,N_9160);
nor U10678 (N_10678,N_9835,N_9868);
and U10679 (N_10679,N_9162,N_9661);
xor U10680 (N_10680,N_9446,N_9834);
and U10681 (N_10681,N_9283,N_9909);
or U10682 (N_10682,N_9668,N_9250);
nor U10683 (N_10683,N_9764,N_9268);
xnor U10684 (N_10684,N_9921,N_9976);
and U10685 (N_10685,N_9211,N_9052);
and U10686 (N_10686,N_9615,N_9937);
nor U10687 (N_10687,N_9685,N_9309);
xnor U10688 (N_10688,N_9974,N_9904);
nand U10689 (N_10689,N_9118,N_9399);
xnor U10690 (N_10690,N_9796,N_9159);
and U10691 (N_10691,N_9829,N_9520);
and U10692 (N_10692,N_9775,N_9720);
or U10693 (N_10693,N_9523,N_9576);
nor U10694 (N_10694,N_9085,N_9161);
nand U10695 (N_10695,N_9410,N_9722);
nor U10696 (N_10696,N_9479,N_9654);
xnor U10697 (N_10697,N_9891,N_9734);
and U10698 (N_10698,N_9539,N_9497);
or U10699 (N_10699,N_9776,N_9435);
or U10700 (N_10700,N_9135,N_9706);
and U10701 (N_10701,N_9072,N_9869);
and U10702 (N_10702,N_9849,N_9493);
and U10703 (N_10703,N_9901,N_9005);
and U10704 (N_10704,N_9298,N_9218);
nor U10705 (N_10705,N_9130,N_9658);
nor U10706 (N_10706,N_9437,N_9113);
and U10707 (N_10707,N_9796,N_9492);
nor U10708 (N_10708,N_9048,N_9924);
or U10709 (N_10709,N_9660,N_9829);
xnor U10710 (N_10710,N_9832,N_9646);
nor U10711 (N_10711,N_9627,N_9478);
nor U10712 (N_10712,N_9689,N_9774);
xor U10713 (N_10713,N_9285,N_9462);
or U10714 (N_10714,N_9230,N_9943);
and U10715 (N_10715,N_9571,N_9591);
and U10716 (N_10716,N_9795,N_9604);
nor U10717 (N_10717,N_9411,N_9273);
xnor U10718 (N_10718,N_9705,N_9973);
xnor U10719 (N_10719,N_9971,N_9141);
or U10720 (N_10720,N_9663,N_9560);
or U10721 (N_10721,N_9668,N_9457);
and U10722 (N_10722,N_9484,N_9965);
xor U10723 (N_10723,N_9438,N_9176);
and U10724 (N_10724,N_9310,N_9957);
nand U10725 (N_10725,N_9563,N_9772);
and U10726 (N_10726,N_9237,N_9941);
nor U10727 (N_10727,N_9935,N_9793);
and U10728 (N_10728,N_9044,N_9646);
xnor U10729 (N_10729,N_9890,N_9448);
xor U10730 (N_10730,N_9162,N_9933);
or U10731 (N_10731,N_9629,N_9815);
and U10732 (N_10732,N_9714,N_9117);
nor U10733 (N_10733,N_9553,N_9389);
and U10734 (N_10734,N_9807,N_9431);
nand U10735 (N_10735,N_9838,N_9667);
and U10736 (N_10736,N_9535,N_9824);
or U10737 (N_10737,N_9786,N_9925);
nand U10738 (N_10738,N_9490,N_9350);
xor U10739 (N_10739,N_9596,N_9571);
xnor U10740 (N_10740,N_9449,N_9389);
nor U10741 (N_10741,N_9431,N_9231);
nor U10742 (N_10742,N_9107,N_9634);
xor U10743 (N_10743,N_9854,N_9798);
nor U10744 (N_10744,N_9632,N_9326);
nand U10745 (N_10745,N_9301,N_9791);
nand U10746 (N_10746,N_9586,N_9270);
xor U10747 (N_10747,N_9145,N_9057);
nor U10748 (N_10748,N_9846,N_9984);
xnor U10749 (N_10749,N_9135,N_9580);
nor U10750 (N_10750,N_9509,N_9413);
and U10751 (N_10751,N_9898,N_9706);
nor U10752 (N_10752,N_9903,N_9931);
or U10753 (N_10753,N_9732,N_9517);
nand U10754 (N_10754,N_9012,N_9384);
nor U10755 (N_10755,N_9851,N_9148);
nor U10756 (N_10756,N_9405,N_9335);
or U10757 (N_10757,N_9048,N_9844);
nand U10758 (N_10758,N_9305,N_9381);
nand U10759 (N_10759,N_9301,N_9432);
nor U10760 (N_10760,N_9493,N_9382);
and U10761 (N_10761,N_9638,N_9492);
and U10762 (N_10762,N_9308,N_9152);
xnor U10763 (N_10763,N_9627,N_9760);
nor U10764 (N_10764,N_9142,N_9809);
nand U10765 (N_10765,N_9982,N_9439);
or U10766 (N_10766,N_9548,N_9686);
or U10767 (N_10767,N_9638,N_9029);
and U10768 (N_10768,N_9640,N_9796);
nand U10769 (N_10769,N_9653,N_9858);
or U10770 (N_10770,N_9963,N_9265);
and U10771 (N_10771,N_9313,N_9990);
nand U10772 (N_10772,N_9268,N_9640);
nand U10773 (N_10773,N_9966,N_9110);
and U10774 (N_10774,N_9065,N_9405);
or U10775 (N_10775,N_9736,N_9929);
xor U10776 (N_10776,N_9778,N_9846);
nor U10777 (N_10777,N_9190,N_9034);
nor U10778 (N_10778,N_9640,N_9093);
xnor U10779 (N_10779,N_9387,N_9636);
nor U10780 (N_10780,N_9784,N_9738);
nor U10781 (N_10781,N_9392,N_9164);
nor U10782 (N_10782,N_9181,N_9129);
and U10783 (N_10783,N_9443,N_9930);
nand U10784 (N_10784,N_9485,N_9318);
xor U10785 (N_10785,N_9218,N_9919);
and U10786 (N_10786,N_9037,N_9542);
xor U10787 (N_10787,N_9253,N_9716);
nand U10788 (N_10788,N_9071,N_9094);
xnor U10789 (N_10789,N_9911,N_9514);
nand U10790 (N_10790,N_9962,N_9916);
xor U10791 (N_10791,N_9992,N_9851);
and U10792 (N_10792,N_9174,N_9612);
nor U10793 (N_10793,N_9408,N_9644);
nor U10794 (N_10794,N_9979,N_9683);
or U10795 (N_10795,N_9127,N_9521);
nand U10796 (N_10796,N_9004,N_9317);
xor U10797 (N_10797,N_9057,N_9619);
nor U10798 (N_10798,N_9502,N_9531);
xnor U10799 (N_10799,N_9777,N_9123);
nand U10800 (N_10800,N_9843,N_9731);
and U10801 (N_10801,N_9028,N_9056);
xnor U10802 (N_10802,N_9571,N_9373);
nand U10803 (N_10803,N_9967,N_9619);
and U10804 (N_10804,N_9354,N_9589);
nor U10805 (N_10805,N_9597,N_9236);
or U10806 (N_10806,N_9031,N_9243);
or U10807 (N_10807,N_9010,N_9385);
and U10808 (N_10808,N_9816,N_9163);
xor U10809 (N_10809,N_9487,N_9666);
nor U10810 (N_10810,N_9848,N_9959);
and U10811 (N_10811,N_9560,N_9470);
xnor U10812 (N_10812,N_9417,N_9315);
or U10813 (N_10813,N_9712,N_9913);
xnor U10814 (N_10814,N_9902,N_9354);
xnor U10815 (N_10815,N_9948,N_9340);
nand U10816 (N_10816,N_9106,N_9367);
nand U10817 (N_10817,N_9740,N_9539);
xor U10818 (N_10818,N_9819,N_9431);
or U10819 (N_10819,N_9594,N_9565);
or U10820 (N_10820,N_9522,N_9344);
nand U10821 (N_10821,N_9170,N_9712);
nor U10822 (N_10822,N_9744,N_9963);
and U10823 (N_10823,N_9667,N_9076);
nand U10824 (N_10824,N_9439,N_9438);
nor U10825 (N_10825,N_9189,N_9322);
xor U10826 (N_10826,N_9444,N_9623);
nor U10827 (N_10827,N_9983,N_9837);
and U10828 (N_10828,N_9053,N_9700);
nor U10829 (N_10829,N_9900,N_9835);
xnor U10830 (N_10830,N_9407,N_9957);
xor U10831 (N_10831,N_9962,N_9068);
nand U10832 (N_10832,N_9046,N_9383);
or U10833 (N_10833,N_9545,N_9632);
nor U10834 (N_10834,N_9917,N_9967);
nand U10835 (N_10835,N_9648,N_9813);
and U10836 (N_10836,N_9511,N_9275);
nor U10837 (N_10837,N_9698,N_9242);
nor U10838 (N_10838,N_9485,N_9796);
and U10839 (N_10839,N_9631,N_9870);
nand U10840 (N_10840,N_9158,N_9209);
or U10841 (N_10841,N_9763,N_9129);
nor U10842 (N_10842,N_9053,N_9358);
nor U10843 (N_10843,N_9369,N_9216);
nor U10844 (N_10844,N_9995,N_9593);
and U10845 (N_10845,N_9861,N_9597);
xnor U10846 (N_10846,N_9807,N_9361);
nand U10847 (N_10847,N_9195,N_9815);
nand U10848 (N_10848,N_9662,N_9483);
nand U10849 (N_10849,N_9269,N_9882);
nand U10850 (N_10850,N_9781,N_9773);
and U10851 (N_10851,N_9201,N_9265);
nor U10852 (N_10852,N_9986,N_9133);
or U10853 (N_10853,N_9327,N_9850);
xor U10854 (N_10854,N_9875,N_9597);
nand U10855 (N_10855,N_9193,N_9677);
or U10856 (N_10856,N_9559,N_9235);
nor U10857 (N_10857,N_9328,N_9069);
xnor U10858 (N_10858,N_9960,N_9544);
xor U10859 (N_10859,N_9828,N_9887);
nand U10860 (N_10860,N_9502,N_9380);
nor U10861 (N_10861,N_9531,N_9837);
and U10862 (N_10862,N_9887,N_9399);
and U10863 (N_10863,N_9378,N_9274);
nor U10864 (N_10864,N_9778,N_9818);
nand U10865 (N_10865,N_9257,N_9255);
nor U10866 (N_10866,N_9989,N_9433);
and U10867 (N_10867,N_9772,N_9477);
or U10868 (N_10868,N_9174,N_9198);
nor U10869 (N_10869,N_9411,N_9496);
or U10870 (N_10870,N_9755,N_9905);
nor U10871 (N_10871,N_9551,N_9695);
or U10872 (N_10872,N_9675,N_9783);
or U10873 (N_10873,N_9233,N_9602);
nor U10874 (N_10874,N_9364,N_9399);
xor U10875 (N_10875,N_9580,N_9207);
and U10876 (N_10876,N_9010,N_9045);
or U10877 (N_10877,N_9209,N_9277);
nand U10878 (N_10878,N_9942,N_9204);
or U10879 (N_10879,N_9145,N_9542);
xnor U10880 (N_10880,N_9819,N_9451);
nand U10881 (N_10881,N_9434,N_9175);
nor U10882 (N_10882,N_9968,N_9555);
and U10883 (N_10883,N_9754,N_9566);
or U10884 (N_10884,N_9095,N_9722);
nor U10885 (N_10885,N_9567,N_9360);
or U10886 (N_10886,N_9118,N_9326);
nand U10887 (N_10887,N_9632,N_9210);
nor U10888 (N_10888,N_9425,N_9991);
and U10889 (N_10889,N_9015,N_9677);
nand U10890 (N_10890,N_9079,N_9229);
and U10891 (N_10891,N_9248,N_9211);
or U10892 (N_10892,N_9951,N_9764);
nand U10893 (N_10893,N_9509,N_9771);
xor U10894 (N_10894,N_9640,N_9673);
nand U10895 (N_10895,N_9297,N_9702);
and U10896 (N_10896,N_9344,N_9956);
nand U10897 (N_10897,N_9310,N_9811);
nand U10898 (N_10898,N_9256,N_9275);
or U10899 (N_10899,N_9829,N_9309);
or U10900 (N_10900,N_9578,N_9074);
nand U10901 (N_10901,N_9911,N_9111);
nor U10902 (N_10902,N_9054,N_9937);
nor U10903 (N_10903,N_9820,N_9131);
and U10904 (N_10904,N_9689,N_9906);
xor U10905 (N_10905,N_9140,N_9578);
nor U10906 (N_10906,N_9621,N_9478);
and U10907 (N_10907,N_9695,N_9882);
nor U10908 (N_10908,N_9912,N_9410);
and U10909 (N_10909,N_9105,N_9887);
nand U10910 (N_10910,N_9629,N_9569);
or U10911 (N_10911,N_9244,N_9252);
nand U10912 (N_10912,N_9521,N_9332);
xor U10913 (N_10913,N_9656,N_9575);
nor U10914 (N_10914,N_9355,N_9476);
or U10915 (N_10915,N_9275,N_9062);
nor U10916 (N_10916,N_9628,N_9559);
or U10917 (N_10917,N_9267,N_9541);
or U10918 (N_10918,N_9461,N_9163);
nand U10919 (N_10919,N_9897,N_9002);
and U10920 (N_10920,N_9774,N_9750);
xnor U10921 (N_10921,N_9474,N_9153);
and U10922 (N_10922,N_9702,N_9187);
or U10923 (N_10923,N_9635,N_9182);
nand U10924 (N_10924,N_9161,N_9061);
xnor U10925 (N_10925,N_9983,N_9120);
and U10926 (N_10926,N_9263,N_9015);
nand U10927 (N_10927,N_9550,N_9502);
nor U10928 (N_10928,N_9745,N_9505);
xor U10929 (N_10929,N_9910,N_9401);
nor U10930 (N_10930,N_9964,N_9115);
nor U10931 (N_10931,N_9934,N_9135);
xor U10932 (N_10932,N_9457,N_9672);
nor U10933 (N_10933,N_9867,N_9917);
xnor U10934 (N_10934,N_9011,N_9405);
or U10935 (N_10935,N_9535,N_9123);
nor U10936 (N_10936,N_9114,N_9471);
xnor U10937 (N_10937,N_9256,N_9211);
nor U10938 (N_10938,N_9924,N_9359);
and U10939 (N_10939,N_9926,N_9340);
xnor U10940 (N_10940,N_9989,N_9727);
nor U10941 (N_10941,N_9283,N_9875);
nor U10942 (N_10942,N_9947,N_9277);
nand U10943 (N_10943,N_9149,N_9015);
xnor U10944 (N_10944,N_9646,N_9685);
nand U10945 (N_10945,N_9990,N_9597);
and U10946 (N_10946,N_9722,N_9622);
nand U10947 (N_10947,N_9638,N_9587);
or U10948 (N_10948,N_9095,N_9452);
and U10949 (N_10949,N_9148,N_9887);
and U10950 (N_10950,N_9330,N_9376);
or U10951 (N_10951,N_9179,N_9519);
and U10952 (N_10952,N_9811,N_9927);
xnor U10953 (N_10953,N_9310,N_9128);
or U10954 (N_10954,N_9310,N_9991);
or U10955 (N_10955,N_9240,N_9297);
and U10956 (N_10956,N_9360,N_9459);
and U10957 (N_10957,N_9703,N_9405);
nand U10958 (N_10958,N_9240,N_9454);
nor U10959 (N_10959,N_9742,N_9737);
or U10960 (N_10960,N_9822,N_9273);
or U10961 (N_10961,N_9903,N_9193);
and U10962 (N_10962,N_9778,N_9112);
nand U10963 (N_10963,N_9246,N_9625);
and U10964 (N_10964,N_9867,N_9341);
nand U10965 (N_10965,N_9689,N_9886);
and U10966 (N_10966,N_9833,N_9216);
xor U10967 (N_10967,N_9795,N_9126);
or U10968 (N_10968,N_9181,N_9538);
xor U10969 (N_10969,N_9776,N_9100);
xnor U10970 (N_10970,N_9709,N_9575);
and U10971 (N_10971,N_9366,N_9985);
xor U10972 (N_10972,N_9649,N_9611);
nand U10973 (N_10973,N_9314,N_9538);
nor U10974 (N_10974,N_9012,N_9569);
nand U10975 (N_10975,N_9762,N_9065);
xnor U10976 (N_10976,N_9354,N_9368);
nor U10977 (N_10977,N_9103,N_9689);
and U10978 (N_10978,N_9415,N_9880);
or U10979 (N_10979,N_9027,N_9164);
or U10980 (N_10980,N_9606,N_9543);
and U10981 (N_10981,N_9850,N_9078);
or U10982 (N_10982,N_9447,N_9569);
and U10983 (N_10983,N_9630,N_9919);
nand U10984 (N_10984,N_9460,N_9693);
and U10985 (N_10985,N_9654,N_9392);
xnor U10986 (N_10986,N_9911,N_9908);
xor U10987 (N_10987,N_9028,N_9744);
or U10988 (N_10988,N_9332,N_9747);
nor U10989 (N_10989,N_9249,N_9894);
or U10990 (N_10990,N_9437,N_9501);
nor U10991 (N_10991,N_9419,N_9731);
xor U10992 (N_10992,N_9114,N_9271);
or U10993 (N_10993,N_9843,N_9016);
nor U10994 (N_10994,N_9351,N_9783);
xor U10995 (N_10995,N_9152,N_9343);
xnor U10996 (N_10996,N_9569,N_9671);
or U10997 (N_10997,N_9445,N_9513);
or U10998 (N_10998,N_9013,N_9397);
nand U10999 (N_10999,N_9936,N_9612);
and U11000 (N_11000,N_10044,N_10843);
or U11001 (N_11001,N_10102,N_10218);
and U11002 (N_11002,N_10741,N_10826);
nand U11003 (N_11003,N_10671,N_10602);
and U11004 (N_11004,N_10118,N_10417);
nor U11005 (N_11005,N_10321,N_10713);
nor U11006 (N_11006,N_10346,N_10476);
and U11007 (N_11007,N_10923,N_10556);
nand U11008 (N_11008,N_10731,N_10136);
or U11009 (N_11009,N_10469,N_10122);
or U11010 (N_11010,N_10284,N_10520);
and U11011 (N_11011,N_10060,N_10782);
nor U11012 (N_11012,N_10229,N_10088);
nor U11013 (N_11013,N_10675,N_10299);
nor U11014 (N_11014,N_10402,N_10553);
nand U11015 (N_11015,N_10623,N_10371);
xnor U11016 (N_11016,N_10811,N_10813);
and U11017 (N_11017,N_10311,N_10139);
or U11018 (N_11018,N_10726,N_10512);
or U11019 (N_11019,N_10614,N_10239);
nand U11020 (N_11020,N_10026,N_10423);
or U11021 (N_11021,N_10945,N_10651);
xor U11022 (N_11022,N_10703,N_10230);
xnor U11023 (N_11023,N_10497,N_10388);
and U11024 (N_11024,N_10027,N_10844);
and U11025 (N_11025,N_10537,N_10976);
or U11026 (N_11026,N_10415,N_10339);
nand U11027 (N_11027,N_10667,N_10117);
or U11028 (N_11028,N_10806,N_10133);
nor U11029 (N_11029,N_10361,N_10748);
xnor U11030 (N_11030,N_10808,N_10446);
xnor U11031 (N_11031,N_10149,N_10198);
and U11032 (N_11032,N_10561,N_10482);
nand U11033 (N_11033,N_10805,N_10653);
and U11034 (N_11034,N_10982,N_10751);
or U11035 (N_11035,N_10327,N_10268);
xnor U11036 (N_11036,N_10781,N_10473);
or U11037 (N_11037,N_10892,N_10453);
xnor U11038 (N_11038,N_10507,N_10522);
or U11039 (N_11039,N_10951,N_10021);
xor U11040 (N_11040,N_10169,N_10246);
and U11041 (N_11041,N_10378,N_10256);
and U11042 (N_11042,N_10664,N_10083);
xnor U11043 (N_11043,N_10160,N_10154);
or U11044 (N_11044,N_10445,N_10135);
nor U11045 (N_11045,N_10106,N_10112);
nand U11046 (N_11046,N_10514,N_10297);
or U11047 (N_11047,N_10411,N_10901);
or U11048 (N_11048,N_10931,N_10778);
nand U11049 (N_11049,N_10358,N_10184);
and U11050 (N_11050,N_10946,N_10063);
and U11051 (N_11051,N_10288,N_10221);
and U11052 (N_11052,N_10457,N_10087);
and U11053 (N_11053,N_10927,N_10168);
or U11054 (N_11054,N_10949,N_10408);
nand U11055 (N_11055,N_10206,N_10696);
xnor U11056 (N_11056,N_10144,N_10829);
or U11057 (N_11057,N_10565,N_10278);
xnor U11058 (N_11058,N_10134,N_10884);
xor U11059 (N_11059,N_10600,N_10290);
nor U11060 (N_11060,N_10503,N_10092);
nor U11061 (N_11061,N_10909,N_10627);
xnor U11062 (N_11062,N_10236,N_10666);
nand U11063 (N_11063,N_10377,N_10451);
nor U11064 (N_11064,N_10360,N_10677);
nor U11065 (N_11065,N_10131,N_10615);
and U11066 (N_11066,N_10138,N_10201);
nand U11067 (N_11067,N_10478,N_10539);
nor U11068 (N_11068,N_10430,N_10597);
and U11069 (N_11069,N_10210,N_10858);
nor U11070 (N_11070,N_10868,N_10886);
nand U11071 (N_11071,N_10672,N_10281);
nand U11072 (N_11072,N_10763,N_10213);
and U11073 (N_11073,N_10030,N_10846);
or U11074 (N_11074,N_10908,N_10783);
nand U11075 (N_11075,N_10978,N_10510);
or U11076 (N_11076,N_10744,N_10504);
xnor U11077 (N_11077,N_10424,N_10161);
xor U11078 (N_11078,N_10082,N_10799);
xnor U11079 (N_11079,N_10691,N_10412);
or U11080 (N_11080,N_10634,N_10240);
or U11081 (N_11081,N_10099,N_10014);
or U11082 (N_11082,N_10644,N_10570);
nor U11083 (N_11083,N_10456,N_10069);
and U11084 (N_11084,N_10965,N_10568);
or U11085 (N_11085,N_10295,N_10084);
nand U11086 (N_11086,N_10993,N_10436);
nor U11087 (N_11087,N_10387,N_10287);
and U11088 (N_11088,N_10598,N_10227);
or U11089 (N_11089,N_10832,N_10990);
and U11090 (N_11090,N_10324,N_10985);
or U11091 (N_11091,N_10625,N_10925);
nor U11092 (N_11092,N_10207,N_10438);
and U11093 (N_11093,N_10646,N_10753);
nor U11094 (N_11094,N_10277,N_10319);
nor U11095 (N_11095,N_10934,N_10900);
nor U11096 (N_11096,N_10015,N_10740);
nand U11097 (N_11097,N_10337,N_10831);
nor U11098 (N_11098,N_10699,N_10483);
or U11099 (N_11099,N_10242,N_10419);
and U11100 (N_11100,N_10906,N_10452);
nor U11101 (N_11101,N_10390,N_10918);
or U11102 (N_11102,N_10313,N_10120);
or U11103 (N_11103,N_10493,N_10146);
and U11104 (N_11104,N_10269,N_10340);
xnor U11105 (N_11105,N_10479,N_10992);
nor U11106 (N_11106,N_10273,N_10543);
and U11107 (N_11107,N_10717,N_10401);
nand U11108 (N_11108,N_10932,N_10279);
nand U11109 (N_11109,N_10955,N_10687);
nor U11110 (N_11110,N_10635,N_10124);
nand U11111 (N_11111,N_10797,N_10980);
and U11112 (N_11112,N_10066,N_10655);
xnor U11113 (N_11113,N_10055,N_10854);
or U11114 (N_11114,N_10305,N_10878);
and U11115 (N_11115,N_10253,N_10864);
nor U11116 (N_11116,N_10645,N_10166);
xnor U11117 (N_11117,N_10716,N_10397);
nor U11118 (N_11118,N_10839,N_10620);
nor U11119 (N_11119,N_10787,N_10053);
or U11120 (N_11120,N_10454,N_10370);
and U11121 (N_11121,N_10759,N_10243);
nor U11122 (N_11122,N_10536,N_10989);
and U11123 (N_11123,N_10865,N_10683);
nor U11124 (N_11124,N_10604,N_10622);
xor U11125 (N_11125,N_10848,N_10559);
xnor U11126 (N_11126,N_10234,N_10766);
nand U11127 (N_11127,N_10263,N_10629);
xnor U11128 (N_11128,N_10987,N_10266);
or U11129 (N_11129,N_10132,N_10040);
and U11130 (N_11130,N_10595,N_10405);
xnor U11131 (N_11131,N_10572,N_10583);
nor U11132 (N_11132,N_10289,N_10861);
xor U11133 (N_11133,N_10029,N_10914);
nor U11134 (N_11134,N_10870,N_10538);
and U11135 (N_11135,N_10472,N_10241);
nand U11136 (N_11136,N_10577,N_10286);
and U11137 (N_11137,N_10723,N_10714);
nand U11138 (N_11138,N_10163,N_10527);
or U11139 (N_11139,N_10298,N_10704);
and U11140 (N_11140,N_10558,N_10711);
xnor U11141 (N_11141,N_10755,N_10317);
xor U11142 (N_11142,N_10694,N_10150);
nor U11143 (N_11143,N_10905,N_10750);
nor U11144 (N_11144,N_10697,N_10798);
nand U11145 (N_11145,N_10056,N_10502);
xor U11146 (N_11146,N_10073,N_10208);
xnor U11147 (N_11147,N_10009,N_10462);
or U11148 (N_11148,N_10959,N_10214);
and U11149 (N_11149,N_10251,N_10676);
xor U11150 (N_11150,N_10640,N_10524);
and U11151 (N_11151,N_10369,N_10768);
or U11152 (N_11152,N_10657,N_10735);
xnor U11153 (N_11153,N_10455,N_10877);
nand U11154 (N_11154,N_10219,N_10828);
xnor U11155 (N_11155,N_10307,N_10869);
or U11156 (N_11156,N_10636,N_10506);
xnor U11157 (N_11157,N_10052,N_10283);
nand U11158 (N_11158,N_10111,N_10019);
or U11159 (N_11159,N_10167,N_10668);
nor U11160 (N_11160,N_10964,N_10833);
nor U11161 (N_11161,N_10526,N_10681);
or U11162 (N_11162,N_10101,N_10262);
nand U11163 (N_11163,N_10148,N_10164);
and U11164 (N_11164,N_10107,N_10762);
nand U11165 (N_11165,N_10173,N_10579);
nor U11166 (N_11166,N_10971,N_10116);
xnor U11167 (N_11167,N_10081,N_10587);
and U11168 (N_11168,N_10958,N_10563);
and U11169 (N_11169,N_10754,N_10724);
and U11170 (N_11170,N_10356,N_10062);
and U11171 (N_11171,N_10329,N_10090);
and U11172 (N_11172,N_10035,N_10128);
or U11173 (N_11173,N_10757,N_10810);
or U11174 (N_11174,N_10464,N_10531);
or U11175 (N_11175,N_10354,N_10274);
xnor U11176 (N_11176,N_10126,N_10873);
xnor U11177 (N_11177,N_10679,N_10431);
nand U11178 (N_11178,N_10979,N_10688);
or U11179 (N_11179,N_10143,N_10517);
nand U11180 (N_11180,N_10547,N_10937);
nor U11181 (N_11181,N_10863,N_10566);
xnor U11182 (N_11182,N_10816,N_10114);
and U11183 (N_11183,N_10626,N_10367);
nand U11184 (N_11184,N_10596,N_10859);
nor U11185 (N_11185,N_10496,N_10986);
and U11186 (N_11186,N_10049,N_10012);
xor U11187 (N_11187,N_10785,N_10141);
nand U11188 (N_11188,N_10880,N_10093);
or U11189 (N_11189,N_10187,N_10907);
or U11190 (N_11190,N_10654,N_10611);
and U11191 (N_11191,N_10048,N_10002);
nand U11192 (N_11192,N_10197,N_10612);
and U11193 (N_11193,N_10215,N_10669);
nor U11194 (N_11194,N_10818,N_10700);
xnor U11195 (N_11195,N_10020,N_10998);
nand U11196 (N_11196,N_10225,N_10732);
nand U11197 (N_11197,N_10643,N_10267);
nor U11198 (N_11198,N_10772,N_10389);
and U11199 (N_11199,N_10233,N_10638);
nand U11200 (N_11200,N_10463,N_10326);
nand U11201 (N_11201,N_10334,N_10363);
nand U11202 (N_11202,N_10328,N_10919);
or U11203 (N_11203,N_10881,N_10940);
and U11204 (N_11204,N_10871,N_10079);
xor U11205 (N_11205,N_10571,N_10933);
nor U11206 (N_11206,N_10875,N_10774);
xor U11207 (N_11207,N_10322,N_10830);
nand U11208 (N_11208,N_10071,N_10814);
and U11209 (N_11209,N_10264,N_10847);
xnor U11210 (N_11210,N_10743,N_10205);
nand U11211 (N_11211,N_10926,N_10963);
nand U11212 (N_11212,N_10862,N_10567);
nand U11213 (N_11213,N_10342,N_10249);
nor U11214 (N_11214,N_10386,N_10031);
xor U11215 (N_11215,N_10939,N_10719);
or U11216 (N_11216,N_10938,N_10656);
xnor U11217 (N_11217,N_10722,N_10248);
nor U11218 (N_11218,N_10275,N_10705);
and U11219 (N_11219,N_10038,N_10712);
xor U11220 (N_11220,N_10192,N_10997);
and U11221 (N_11221,N_10542,N_10824);
or U11222 (N_11222,N_10935,N_10776);
nor U11223 (N_11223,N_10529,N_10067);
nand U11224 (N_11224,N_10410,N_10359);
nor U11225 (N_11225,N_10085,N_10756);
or U11226 (N_11226,N_10845,N_10301);
and U11227 (N_11227,N_10994,N_10585);
or U11228 (N_11228,N_10792,N_10265);
xnor U11229 (N_11229,N_10403,N_10338);
or U11230 (N_11230,N_10609,N_10533);
or U11231 (N_11231,N_10123,N_10812);
nand U11232 (N_11232,N_10302,N_10588);
and U11233 (N_11233,N_10701,N_10057);
nand U11234 (N_11234,N_10488,N_10721);
xnor U11235 (N_11235,N_10915,N_10548);
xnor U11236 (N_11236,N_10420,N_10385);
and U11237 (N_11237,N_10380,N_10195);
and U11238 (N_11238,N_10649,N_10803);
nand U11239 (N_11239,N_10991,N_10827);
nor U11240 (N_11240,N_10639,N_10406);
or U11241 (N_11241,N_10791,N_10137);
xnor U11242 (N_11242,N_10795,N_10663);
nand U11243 (N_11243,N_10364,N_10471);
xor U11244 (N_11244,N_10530,N_10684);
nor U11245 (N_11245,N_10680,N_10760);
nor U11246 (N_11246,N_10544,N_10211);
nand U11247 (N_11247,N_10974,N_10516);
xnor U11248 (N_11248,N_10842,N_10366);
nand U11249 (N_11249,N_10292,N_10409);
or U11250 (N_11250,N_10365,N_10442);
or U11251 (N_11251,N_10037,N_10250);
or U11252 (N_11252,N_10303,N_10414);
nand U11253 (N_11253,N_10003,N_10749);
nand U11254 (N_11254,N_10383,N_10899);
and U11255 (N_11255,N_10474,N_10058);
xor U11256 (N_11256,N_10183,N_10105);
nor U11257 (N_11257,N_10500,N_10426);
or U11258 (N_11258,N_10841,N_10235);
or U11259 (N_11259,N_10551,N_10575);
or U11260 (N_11260,N_10127,N_10835);
nand U11261 (N_11261,N_10856,N_10304);
nor U11262 (N_11262,N_10059,N_10790);
nand U11263 (N_11263,N_10070,N_10441);
xnor U11264 (N_11264,N_10280,N_10220);
or U11265 (N_11265,N_10838,N_10222);
or U11266 (N_11266,N_10153,N_10590);
and U11267 (N_11267,N_10616,N_10698);
nor U11268 (N_11268,N_10204,N_10809);
or U11269 (N_11269,N_10022,N_10942);
xnor U11270 (N_11270,N_10376,N_10323);
nor U11271 (N_11271,N_10574,N_10852);
nand U11272 (N_11272,N_10891,N_10924);
or U11273 (N_11273,N_10121,N_10196);
nor U11274 (N_11274,N_10039,N_10011);
nand U11275 (N_11275,N_10580,N_10013);
or U11276 (N_11276,N_10519,N_10761);
or U11277 (N_11277,N_10586,N_10540);
or U11278 (N_11278,N_10624,N_10525);
or U11279 (N_11279,N_10076,N_10465);
and U11280 (N_11280,N_10860,N_10080);
or U11281 (N_11281,N_10557,N_10293);
xor U11282 (N_11282,N_10421,N_10996);
xor U11283 (N_11283,N_10392,N_10000);
nand U11284 (N_11284,N_10125,N_10180);
and U11285 (N_11285,N_10418,N_10975);
nand U11286 (N_11286,N_10738,N_10172);
nor U11287 (N_11287,N_10034,N_10912);
or U11288 (N_11288,N_10347,N_10470);
xnor U11289 (N_11289,N_10162,N_10458);
xor U11290 (N_11290,N_10606,N_10103);
and U11291 (N_11291,N_10486,N_10320);
and U11292 (N_11292,N_10742,N_10840);
xor U11293 (N_11293,N_10461,N_10223);
and U11294 (N_11294,N_10115,N_10023);
and U11295 (N_11295,N_10395,N_10505);
or U11296 (N_11296,N_10381,N_10678);
nor U11297 (N_11297,N_10282,N_10310);
nor U11298 (N_11298,N_10897,N_10247);
xor U11299 (N_11299,N_10564,N_10231);
xor U11300 (N_11300,N_10786,N_10895);
or U11301 (N_11301,N_10535,N_10155);
nor U11302 (N_11302,N_10447,N_10074);
nand U11303 (N_11303,N_10294,N_10186);
and U11304 (N_11304,N_10511,N_10613);
and U11305 (N_11305,N_10707,N_10552);
nand U11306 (N_11306,N_10736,N_10352);
xor U11307 (N_11307,N_10518,N_10400);
and U11308 (N_11308,N_10007,N_10882);
nor U11309 (N_11309,N_10046,N_10618);
nand U11310 (N_11310,N_10708,N_10309);
xnor U11311 (N_11311,N_10521,N_10513);
nand U11312 (N_11312,N_10212,N_10177);
and U11313 (N_11313,N_10660,N_10170);
nor U11314 (N_11314,N_10175,N_10662);
and U11315 (N_11315,N_10966,N_10728);
nand U11316 (N_11316,N_10815,N_10821);
nor U11317 (N_11317,N_10437,N_10739);
or U11318 (N_11318,N_10331,N_10043);
nand U11319 (N_11319,N_10802,N_10151);
xor U11320 (N_11320,N_10866,N_10592);
or U11321 (N_11321,N_10788,N_10481);
or U11322 (N_11322,N_10771,N_10898);
nand U11323 (N_11323,N_10355,N_10439);
and U11324 (N_11324,N_10917,N_10498);
or U11325 (N_11325,N_10382,N_10333);
nor U11326 (N_11326,N_10306,N_10147);
nor U11327 (N_11327,N_10372,N_10422);
or U11328 (N_11328,N_10335,N_10374);
nand U11329 (N_11329,N_10545,N_10819);
nand U11330 (N_11330,N_10670,N_10075);
nand U11331 (N_11331,N_10850,N_10693);
or U11332 (N_11332,N_10028,N_10836);
nand U11333 (N_11333,N_10822,N_10404);
or U11334 (N_11334,N_10984,N_10330);
and U11335 (N_11335,N_10779,N_10769);
xor U11336 (N_11336,N_10784,N_10315);
nor U11337 (N_11337,N_10129,N_10887);
and U11338 (N_11338,N_10534,N_10350);
and U11339 (N_11339,N_10199,N_10801);
nor U11340 (N_11340,N_10272,N_10006);
or U11341 (N_11341,N_10254,N_10032);
xnor U11342 (N_11342,N_10752,N_10226);
nand U11343 (N_11343,N_10632,N_10661);
nand U11344 (N_11344,N_10094,N_10921);
xor U11345 (N_11345,N_10216,N_10849);
and U11346 (N_11346,N_10176,N_10110);
nor U11347 (N_11347,N_10098,N_10398);
nand U11348 (N_11348,N_10432,N_10777);
nand U11349 (N_11349,N_10546,N_10232);
or U11350 (N_11350,N_10953,N_10560);
nor U11351 (N_11351,N_10351,N_10332);
and U11352 (N_11352,N_10394,N_10650);
nand U11353 (N_11353,N_10930,N_10158);
nor U11354 (N_11354,N_10348,N_10800);
nor U11355 (N_11355,N_10140,N_10261);
nor U11356 (N_11356,N_10448,N_10746);
or U11357 (N_11357,N_10276,N_10343);
nor U11358 (N_11358,N_10944,N_10633);
or U11359 (N_11359,N_10064,N_10922);
nor U11360 (N_11360,N_10484,N_10807);
and U11361 (N_11361,N_10692,N_10189);
nor U11362 (N_11362,N_10825,N_10314);
and U11363 (N_11363,N_10174,N_10368);
or U11364 (N_11364,N_10312,N_10036);
or U11365 (N_11365,N_10674,N_10584);
and U11366 (N_11366,N_10095,N_10960);
xnor U11367 (N_11367,N_10193,N_10157);
xor U11368 (N_11368,N_10630,N_10244);
and U11369 (N_11369,N_10467,N_10061);
or U11370 (N_11370,N_10341,N_10576);
nand U11371 (N_11371,N_10569,N_10086);
xor U11372 (N_11372,N_10523,N_10449);
and U11373 (N_11373,N_10952,N_10181);
xnor U11374 (N_11374,N_10804,N_10729);
or U11375 (N_11375,N_10549,N_10008);
and U11376 (N_11376,N_10016,N_10904);
nand U11377 (N_11377,N_10983,N_10628);
nor U11378 (N_11378,N_10109,N_10916);
or U11379 (N_11379,N_10072,N_10793);
nor U11380 (N_11380,N_10097,N_10033);
and U11381 (N_11381,N_10734,N_10658);
or U11382 (N_11382,N_10190,N_10641);
xnor U11383 (N_11383,N_10494,N_10745);
or U11384 (N_11384,N_10499,N_10685);
or U11385 (N_11385,N_10973,N_10706);
and U11386 (N_11386,N_10589,N_10608);
and U11387 (N_11387,N_10209,N_10690);
xnor U11388 (N_11388,N_10947,N_10648);
xor U11389 (N_11389,N_10045,N_10005);
xor U11390 (N_11390,N_10773,N_10902);
nor U11391 (N_11391,N_10435,N_10883);
nor U11392 (N_11392,N_10373,N_10999);
or U11393 (N_11393,N_10165,N_10637);
and U11394 (N_11394,N_10948,N_10018);
or U11395 (N_11395,N_10817,N_10528);
or U11396 (N_11396,N_10188,N_10509);
xnor U11397 (N_11397,N_10291,N_10889);
nand U11398 (N_11398,N_10078,N_10903);
nand U11399 (N_11399,N_10720,N_10349);
xor U11400 (N_11400,N_10010,N_10145);
nor U11401 (N_11401,N_10178,N_10345);
and U11402 (N_11402,N_10758,N_10182);
xor U11403 (N_11403,N_10665,N_10433);
xnor U11404 (N_11404,N_10050,N_10194);
nand U11405 (N_11405,N_10047,N_10501);
or U11406 (N_11406,N_10954,N_10968);
xor U11407 (N_11407,N_10961,N_10943);
nand U11408 (N_11408,N_10823,N_10820);
nand U11409 (N_11409,N_10936,N_10104);
nand U11410 (N_11410,N_10893,N_10967);
and U11411 (N_11411,N_10119,N_10554);
and U11412 (N_11412,N_10896,N_10775);
nand U11413 (N_11413,N_10068,N_10300);
xnor U11414 (N_11414,N_10621,N_10399);
xnor U11415 (N_11415,N_10001,N_10325);
xor U11416 (N_11416,N_10384,N_10603);
nand U11417 (N_11417,N_10054,N_10631);
xnor U11418 (N_11418,N_10673,N_10851);
nand U11419 (N_11419,N_10647,N_10591);
xnor U11420 (N_11420,N_10477,N_10780);
nand U11421 (N_11421,N_10867,N_10747);
xor U11422 (N_11422,N_10920,N_10659);
nand U11423 (N_11423,N_10890,N_10710);
nor U11424 (N_11424,N_10308,N_10489);
nor U11425 (N_11425,N_10025,N_10245);
or U11426 (N_11426,N_10407,N_10725);
or U11427 (N_11427,N_10416,N_10593);
xor U11428 (N_11428,N_10228,N_10450);
or U11429 (N_11429,N_10459,N_10879);
and U11430 (N_11430,N_10789,N_10617);
xor U11431 (N_11431,N_10834,N_10108);
and U11432 (N_11432,N_10270,N_10730);
nor U11433 (N_11433,N_10928,N_10396);
nand U11434 (N_11434,N_10362,N_10715);
nand U11435 (N_11435,N_10202,N_10764);
xor U11436 (N_11436,N_10581,N_10874);
xnor U11437 (N_11437,N_10794,N_10872);
xnor U11438 (N_11438,N_10238,N_10532);
or U11439 (N_11439,N_10042,N_10491);
and U11440 (N_11440,N_10393,N_10737);
xnor U11441 (N_11441,N_10796,N_10765);
xnor U11442 (N_11442,N_10041,N_10434);
xor U11443 (N_11443,N_10894,N_10578);
xor U11444 (N_11444,N_10237,N_10257);
and U11445 (N_11445,N_10885,N_10259);
nor U11446 (N_11446,N_10255,N_10427);
xnor U11447 (N_11447,N_10152,N_10508);
xor U11448 (N_11448,N_10857,N_10981);
and U11449 (N_11449,N_10024,N_10357);
or U11450 (N_11450,N_10130,N_10972);
or U11451 (N_11451,N_10573,N_10089);
and U11452 (N_11452,N_10492,N_10096);
nand U11453 (N_11453,N_10191,N_10142);
xnor U11454 (N_11454,N_10440,N_10495);
xnor U11455 (N_11455,N_10913,N_10619);
and U11456 (N_11456,N_10375,N_10950);
nor U11457 (N_11457,N_10336,N_10466);
and U11458 (N_11458,N_10318,N_10652);
or U11459 (N_11459,N_10601,N_10562);
nand U11460 (N_11460,N_10682,N_10468);
or U11461 (N_11461,N_10733,N_10709);
nand U11462 (N_11462,N_10702,N_10429);
nor U11463 (N_11463,N_10091,N_10258);
nor U11464 (N_11464,N_10555,N_10487);
or U11465 (N_11465,N_10217,N_10379);
xnor U11466 (N_11466,N_10910,N_10428);
nor U11467 (N_11467,N_10941,N_10017);
xnor U11468 (N_11468,N_10594,N_10969);
nor U11469 (N_11469,N_10425,N_10260);
xor U11470 (N_11470,N_10970,N_10004);
nor U11471 (N_11471,N_10444,N_10977);
nor U11472 (N_11472,N_10515,N_10460);
and U11473 (N_11473,N_10962,N_10957);
nor U11474 (N_11474,N_10718,N_10296);
nor U11475 (N_11475,N_10490,N_10686);
nor U11476 (N_11476,N_10353,N_10695);
xor U11477 (N_11477,N_10252,N_10988);
and U11478 (N_11478,N_10344,N_10605);
nor U11479 (N_11479,N_10113,N_10100);
xnor U11480 (N_11480,N_10995,N_10610);
or U11481 (N_11481,N_10727,N_10485);
xor U11482 (N_11482,N_10200,N_10285);
and U11483 (N_11483,N_10607,N_10203);
nand U11484 (N_11484,N_10642,N_10837);
or U11485 (N_11485,N_10051,N_10159);
nand U11486 (N_11486,N_10316,N_10271);
xor U11487 (N_11487,N_10956,N_10876);
xnor U11488 (N_11488,N_10185,N_10888);
xnor U11489 (N_11489,N_10853,N_10480);
nor U11490 (N_11490,N_10171,N_10065);
or U11491 (N_11491,N_10911,N_10599);
nand U11492 (N_11492,N_10541,N_10767);
nor U11493 (N_11493,N_10179,N_10929);
or U11494 (N_11494,N_10077,N_10582);
xor U11495 (N_11495,N_10855,N_10413);
or U11496 (N_11496,N_10550,N_10391);
or U11497 (N_11497,N_10689,N_10443);
nor U11498 (N_11498,N_10224,N_10770);
or U11499 (N_11499,N_10475,N_10156);
and U11500 (N_11500,N_10179,N_10661);
xnor U11501 (N_11501,N_10937,N_10814);
and U11502 (N_11502,N_10148,N_10847);
nor U11503 (N_11503,N_10103,N_10309);
xnor U11504 (N_11504,N_10997,N_10749);
nand U11505 (N_11505,N_10016,N_10087);
and U11506 (N_11506,N_10901,N_10140);
xnor U11507 (N_11507,N_10144,N_10992);
nand U11508 (N_11508,N_10959,N_10827);
and U11509 (N_11509,N_10015,N_10339);
nand U11510 (N_11510,N_10138,N_10062);
nor U11511 (N_11511,N_10480,N_10300);
nand U11512 (N_11512,N_10779,N_10849);
xnor U11513 (N_11513,N_10261,N_10928);
and U11514 (N_11514,N_10131,N_10858);
or U11515 (N_11515,N_10549,N_10084);
xor U11516 (N_11516,N_10599,N_10996);
nor U11517 (N_11517,N_10062,N_10727);
or U11518 (N_11518,N_10211,N_10984);
and U11519 (N_11519,N_10418,N_10396);
nor U11520 (N_11520,N_10356,N_10393);
and U11521 (N_11521,N_10674,N_10242);
nand U11522 (N_11522,N_10181,N_10364);
nor U11523 (N_11523,N_10274,N_10909);
nand U11524 (N_11524,N_10842,N_10593);
nor U11525 (N_11525,N_10372,N_10127);
and U11526 (N_11526,N_10938,N_10815);
nand U11527 (N_11527,N_10241,N_10797);
or U11528 (N_11528,N_10361,N_10574);
nor U11529 (N_11529,N_10559,N_10973);
nand U11530 (N_11530,N_10935,N_10985);
nor U11531 (N_11531,N_10092,N_10228);
xnor U11532 (N_11532,N_10447,N_10255);
nand U11533 (N_11533,N_10044,N_10323);
or U11534 (N_11534,N_10760,N_10934);
nor U11535 (N_11535,N_10594,N_10479);
or U11536 (N_11536,N_10506,N_10855);
xnor U11537 (N_11537,N_10651,N_10049);
or U11538 (N_11538,N_10483,N_10990);
or U11539 (N_11539,N_10835,N_10065);
xor U11540 (N_11540,N_10822,N_10684);
nand U11541 (N_11541,N_10059,N_10229);
and U11542 (N_11542,N_10005,N_10344);
xnor U11543 (N_11543,N_10027,N_10066);
and U11544 (N_11544,N_10936,N_10970);
xor U11545 (N_11545,N_10942,N_10890);
xnor U11546 (N_11546,N_10253,N_10837);
nor U11547 (N_11547,N_10521,N_10994);
nand U11548 (N_11548,N_10378,N_10076);
or U11549 (N_11549,N_10189,N_10425);
xor U11550 (N_11550,N_10574,N_10641);
or U11551 (N_11551,N_10257,N_10405);
nand U11552 (N_11552,N_10825,N_10258);
nor U11553 (N_11553,N_10324,N_10672);
xnor U11554 (N_11554,N_10672,N_10421);
nand U11555 (N_11555,N_10692,N_10945);
nand U11556 (N_11556,N_10853,N_10418);
or U11557 (N_11557,N_10846,N_10373);
or U11558 (N_11558,N_10194,N_10208);
nand U11559 (N_11559,N_10684,N_10398);
xnor U11560 (N_11560,N_10436,N_10360);
nand U11561 (N_11561,N_10680,N_10897);
xor U11562 (N_11562,N_10690,N_10312);
nor U11563 (N_11563,N_10290,N_10583);
xor U11564 (N_11564,N_10367,N_10768);
xnor U11565 (N_11565,N_10927,N_10922);
or U11566 (N_11566,N_10722,N_10163);
and U11567 (N_11567,N_10057,N_10975);
or U11568 (N_11568,N_10459,N_10521);
or U11569 (N_11569,N_10301,N_10425);
and U11570 (N_11570,N_10836,N_10498);
and U11571 (N_11571,N_10276,N_10528);
nand U11572 (N_11572,N_10878,N_10210);
or U11573 (N_11573,N_10883,N_10553);
nor U11574 (N_11574,N_10529,N_10484);
nand U11575 (N_11575,N_10702,N_10177);
and U11576 (N_11576,N_10257,N_10981);
nor U11577 (N_11577,N_10684,N_10005);
and U11578 (N_11578,N_10550,N_10069);
or U11579 (N_11579,N_10021,N_10339);
and U11580 (N_11580,N_10172,N_10043);
or U11581 (N_11581,N_10848,N_10050);
and U11582 (N_11582,N_10068,N_10323);
and U11583 (N_11583,N_10564,N_10823);
or U11584 (N_11584,N_10586,N_10396);
nand U11585 (N_11585,N_10418,N_10998);
xor U11586 (N_11586,N_10252,N_10212);
nand U11587 (N_11587,N_10744,N_10191);
nand U11588 (N_11588,N_10937,N_10302);
xor U11589 (N_11589,N_10269,N_10512);
and U11590 (N_11590,N_10089,N_10330);
nor U11591 (N_11591,N_10128,N_10656);
xor U11592 (N_11592,N_10993,N_10233);
and U11593 (N_11593,N_10635,N_10811);
nor U11594 (N_11594,N_10912,N_10015);
xnor U11595 (N_11595,N_10650,N_10084);
nor U11596 (N_11596,N_10755,N_10062);
or U11597 (N_11597,N_10815,N_10208);
xor U11598 (N_11598,N_10853,N_10223);
and U11599 (N_11599,N_10485,N_10413);
or U11600 (N_11600,N_10852,N_10289);
nand U11601 (N_11601,N_10027,N_10666);
or U11602 (N_11602,N_10920,N_10242);
or U11603 (N_11603,N_10275,N_10324);
nand U11604 (N_11604,N_10637,N_10190);
xor U11605 (N_11605,N_10433,N_10970);
nand U11606 (N_11606,N_10378,N_10383);
nand U11607 (N_11607,N_10596,N_10820);
nand U11608 (N_11608,N_10873,N_10983);
nor U11609 (N_11609,N_10149,N_10539);
nor U11610 (N_11610,N_10657,N_10898);
and U11611 (N_11611,N_10400,N_10339);
and U11612 (N_11612,N_10111,N_10945);
nor U11613 (N_11613,N_10343,N_10220);
and U11614 (N_11614,N_10067,N_10375);
nand U11615 (N_11615,N_10292,N_10285);
or U11616 (N_11616,N_10498,N_10049);
and U11617 (N_11617,N_10143,N_10865);
and U11618 (N_11618,N_10556,N_10113);
and U11619 (N_11619,N_10571,N_10910);
nor U11620 (N_11620,N_10464,N_10448);
xor U11621 (N_11621,N_10794,N_10999);
or U11622 (N_11622,N_10411,N_10971);
and U11623 (N_11623,N_10166,N_10267);
or U11624 (N_11624,N_10450,N_10459);
xnor U11625 (N_11625,N_10019,N_10068);
and U11626 (N_11626,N_10341,N_10490);
nand U11627 (N_11627,N_10961,N_10476);
nor U11628 (N_11628,N_10141,N_10192);
xnor U11629 (N_11629,N_10147,N_10542);
and U11630 (N_11630,N_10675,N_10309);
or U11631 (N_11631,N_10761,N_10128);
nor U11632 (N_11632,N_10627,N_10664);
nand U11633 (N_11633,N_10691,N_10470);
xnor U11634 (N_11634,N_10801,N_10041);
and U11635 (N_11635,N_10041,N_10098);
or U11636 (N_11636,N_10468,N_10387);
and U11637 (N_11637,N_10050,N_10525);
nand U11638 (N_11638,N_10932,N_10970);
or U11639 (N_11639,N_10053,N_10323);
or U11640 (N_11640,N_10236,N_10924);
nand U11641 (N_11641,N_10730,N_10676);
and U11642 (N_11642,N_10588,N_10863);
and U11643 (N_11643,N_10742,N_10901);
nand U11644 (N_11644,N_10873,N_10362);
xnor U11645 (N_11645,N_10619,N_10858);
xnor U11646 (N_11646,N_10650,N_10798);
nor U11647 (N_11647,N_10362,N_10756);
nand U11648 (N_11648,N_10576,N_10361);
nand U11649 (N_11649,N_10763,N_10586);
and U11650 (N_11650,N_10628,N_10574);
nor U11651 (N_11651,N_10188,N_10714);
xnor U11652 (N_11652,N_10584,N_10412);
nand U11653 (N_11653,N_10445,N_10179);
and U11654 (N_11654,N_10573,N_10565);
nand U11655 (N_11655,N_10630,N_10541);
nor U11656 (N_11656,N_10650,N_10348);
nor U11657 (N_11657,N_10802,N_10130);
nor U11658 (N_11658,N_10370,N_10319);
and U11659 (N_11659,N_10669,N_10952);
nand U11660 (N_11660,N_10617,N_10723);
xnor U11661 (N_11661,N_10585,N_10323);
and U11662 (N_11662,N_10547,N_10203);
xor U11663 (N_11663,N_10950,N_10640);
nand U11664 (N_11664,N_10261,N_10310);
xnor U11665 (N_11665,N_10079,N_10930);
nand U11666 (N_11666,N_10731,N_10896);
or U11667 (N_11667,N_10098,N_10374);
or U11668 (N_11668,N_10228,N_10618);
and U11669 (N_11669,N_10469,N_10161);
nand U11670 (N_11670,N_10285,N_10655);
and U11671 (N_11671,N_10255,N_10417);
nand U11672 (N_11672,N_10842,N_10032);
nor U11673 (N_11673,N_10070,N_10246);
nand U11674 (N_11674,N_10271,N_10701);
xnor U11675 (N_11675,N_10467,N_10185);
and U11676 (N_11676,N_10322,N_10795);
nand U11677 (N_11677,N_10429,N_10715);
xor U11678 (N_11678,N_10192,N_10664);
nand U11679 (N_11679,N_10862,N_10167);
xnor U11680 (N_11680,N_10261,N_10880);
or U11681 (N_11681,N_10998,N_10429);
nor U11682 (N_11682,N_10393,N_10361);
nor U11683 (N_11683,N_10619,N_10580);
and U11684 (N_11684,N_10464,N_10184);
nand U11685 (N_11685,N_10582,N_10269);
and U11686 (N_11686,N_10577,N_10359);
or U11687 (N_11687,N_10894,N_10003);
or U11688 (N_11688,N_10430,N_10951);
xnor U11689 (N_11689,N_10014,N_10151);
xor U11690 (N_11690,N_10925,N_10585);
and U11691 (N_11691,N_10850,N_10766);
and U11692 (N_11692,N_10221,N_10648);
xnor U11693 (N_11693,N_10898,N_10762);
or U11694 (N_11694,N_10333,N_10122);
xor U11695 (N_11695,N_10988,N_10610);
or U11696 (N_11696,N_10895,N_10061);
and U11697 (N_11697,N_10867,N_10486);
nand U11698 (N_11698,N_10044,N_10095);
nor U11699 (N_11699,N_10441,N_10877);
or U11700 (N_11700,N_10965,N_10711);
and U11701 (N_11701,N_10325,N_10478);
or U11702 (N_11702,N_10989,N_10481);
or U11703 (N_11703,N_10577,N_10054);
nor U11704 (N_11704,N_10964,N_10075);
nand U11705 (N_11705,N_10310,N_10419);
xor U11706 (N_11706,N_10258,N_10641);
xnor U11707 (N_11707,N_10774,N_10699);
and U11708 (N_11708,N_10841,N_10589);
nand U11709 (N_11709,N_10029,N_10281);
nor U11710 (N_11710,N_10909,N_10065);
and U11711 (N_11711,N_10107,N_10832);
and U11712 (N_11712,N_10033,N_10253);
xor U11713 (N_11713,N_10322,N_10839);
nor U11714 (N_11714,N_10391,N_10153);
or U11715 (N_11715,N_10596,N_10421);
xor U11716 (N_11716,N_10296,N_10996);
nor U11717 (N_11717,N_10829,N_10058);
nand U11718 (N_11718,N_10256,N_10522);
nor U11719 (N_11719,N_10337,N_10048);
or U11720 (N_11720,N_10243,N_10476);
or U11721 (N_11721,N_10615,N_10933);
nand U11722 (N_11722,N_10031,N_10059);
and U11723 (N_11723,N_10178,N_10982);
xnor U11724 (N_11724,N_10200,N_10142);
and U11725 (N_11725,N_10701,N_10651);
nand U11726 (N_11726,N_10127,N_10016);
and U11727 (N_11727,N_10932,N_10128);
xnor U11728 (N_11728,N_10552,N_10016);
or U11729 (N_11729,N_10020,N_10389);
or U11730 (N_11730,N_10965,N_10289);
nand U11731 (N_11731,N_10845,N_10895);
xnor U11732 (N_11732,N_10276,N_10301);
xor U11733 (N_11733,N_10291,N_10730);
xnor U11734 (N_11734,N_10164,N_10426);
or U11735 (N_11735,N_10366,N_10392);
nor U11736 (N_11736,N_10290,N_10921);
or U11737 (N_11737,N_10972,N_10797);
nor U11738 (N_11738,N_10661,N_10967);
nor U11739 (N_11739,N_10506,N_10905);
or U11740 (N_11740,N_10413,N_10167);
nor U11741 (N_11741,N_10612,N_10196);
or U11742 (N_11742,N_10437,N_10709);
nor U11743 (N_11743,N_10876,N_10166);
nor U11744 (N_11744,N_10351,N_10526);
and U11745 (N_11745,N_10571,N_10391);
or U11746 (N_11746,N_10362,N_10924);
and U11747 (N_11747,N_10623,N_10066);
and U11748 (N_11748,N_10934,N_10534);
nor U11749 (N_11749,N_10434,N_10063);
and U11750 (N_11750,N_10933,N_10321);
or U11751 (N_11751,N_10432,N_10744);
nand U11752 (N_11752,N_10408,N_10398);
and U11753 (N_11753,N_10576,N_10346);
xor U11754 (N_11754,N_10141,N_10190);
or U11755 (N_11755,N_10319,N_10468);
nor U11756 (N_11756,N_10937,N_10509);
and U11757 (N_11757,N_10547,N_10294);
nor U11758 (N_11758,N_10336,N_10951);
nor U11759 (N_11759,N_10675,N_10048);
nor U11760 (N_11760,N_10498,N_10854);
and U11761 (N_11761,N_10594,N_10149);
and U11762 (N_11762,N_10897,N_10444);
xnor U11763 (N_11763,N_10301,N_10008);
xor U11764 (N_11764,N_10199,N_10919);
or U11765 (N_11765,N_10099,N_10372);
nand U11766 (N_11766,N_10883,N_10002);
nor U11767 (N_11767,N_10560,N_10264);
nand U11768 (N_11768,N_10515,N_10346);
nand U11769 (N_11769,N_10471,N_10525);
or U11770 (N_11770,N_10694,N_10637);
xor U11771 (N_11771,N_10031,N_10358);
xnor U11772 (N_11772,N_10094,N_10632);
and U11773 (N_11773,N_10022,N_10436);
and U11774 (N_11774,N_10040,N_10995);
xor U11775 (N_11775,N_10900,N_10035);
or U11776 (N_11776,N_10630,N_10264);
xnor U11777 (N_11777,N_10292,N_10365);
or U11778 (N_11778,N_10235,N_10470);
nand U11779 (N_11779,N_10920,N_10572);
and U11780 (N_11780,N_10987,N_10041);
nand U11781 (N_11781,N_10779,N_10717);
and U11782 (N_11782,N_10598,N_10058);
and U11783 (N_11783,N_10148,N_10655);
or U11784 (N_11784,N_10869,N_10087);
nor U11785 (N_11785,N_10432,N_10454);
or U11786 (N_11786,N_10511,N_10059);
xnor U11787 (N_11787,N_10028,N_10193);
xor U11788 (N_11788,N_10341,N_10729);
nand U11789 (N_11789,N_10122,N_10976);
and U11790 (N_11790,N_10655,N_10886);
nand U11791 (N_11791,N_10308,N_10111);
nor U11792 (N_11792,N_10231,N_10796);
and U11793 (N_11793,N_10291,N_10354);
nor U11794 (N_11794,N_10407,N_10843);
nand U11795 (N_11795,N_10806,N_10961);
nand U11796 (N_11796,N_10346,N_10053);
nand U11797 (N_11797,N_10073,N_10553);
nor U11798 (N_11798,N_10207,N_10532);
nor U11799 (N_11799,N_10065,N_10892);
nor U11800 (N_11800,N_10525,N_10473);
or U11801 (N_11801,N_10805,N_10314);
and U11802 (N_11802,N_10748,N_10625);
nor U11803 (N_11803,N_10174,N_10765);
xnor U11804 (N_11804,N_10502,N_10581);
and U11805 (N_11805,N_10803,N_10304);
nor U11806 (N_11806,N_10288,N_10588);
nand U11807 (N_11807,N_10779,N_10104);
or U11808 (N_11808,N_10768,N_10187);
xnor U11809 (N_11809,N_10648,N_10403);
nand U11810 (N_11810,N_10532,N_10829);
and U11811 (N_11811,N_10919,N_10862);
nor U11812 (N_11812,N_10138,N_10031);
and U11813 (N_11813,N_10981,N_10909);
xor U11814 (N_11814,N_10056,N_10853);
or U11815 (N_11815,N_10637,N_10145);
nor U11816 (N_11816,N_10716,N_10166);
or U11817 (N_11817,N_10189,N_10600);
or U11818 (N_11818,N_10295,N_10579);
xnor U11819 (N_11819,N_10875,N_10751);
or U11820 (N_11820,N_10852,N_10703);
nor U11821 (N_11821,N_10256,N_10014);
xor U11822 (N_11822,N_10812,N_10639);
nor U11823 (N_11823,N_10627,N_10057);
and U11824 (N_11824,N_10599,N_10356);
nor U11825 (N_11825,N_10476,N_10591);
nor U11826 (N_11826,N_10947,N_10181);
xor U11827 (N_11827,N_10700,N_10972);
and U11828 (N_11828,N_10710,N_10974);
xnor U11829 (N_11829,N_10086,N_10472);
and U11830 (N_11830,N_10732,N_10708);
nand U11831 (N_11831,N_10204,N_10640);
or U11832 (N_11832,N_10331,N_10435);
nand U11833 (N_11833,N_10435,N_10746);
xor U11834 (N_11834,N_10656,N_10046);
xnor U11835 (N_11835,N_10625,N_10075);
and U11836 (N_11836,N_10310,N_10648);
nand U11837 (N_11837,N_10812,N_10644);
xnor U11838 (N_11838,N_10226,N_10904);
xor U11839 (N_11839,N_10227,N_10071);
nand U11840 (N_11840,N_10854,N_10948);
nor U11841 (N_11841,N_10473,N_10348);
nand U11842 (N_11842,N_10217,N_10805);
and U11843 (N_11843,N_10481,N_10112);
nand U11844 (N_11844,N_10560,N_10272);
and U11845 (N_11845,N_10483,N_10056);
or U11846 (N_11846,N_10714,N_10736);
or U11847 (N_11847,N_10651,N_10815);
or U11848 (N_11848,N_10114,N_10692);
and U11849 (N_11849,N_10903,N_10066);
nor U11850 (N_11850,N_10112,N_10663);
xnor U11851 (N_11851,N_10258,N_10098);
or U11852 (N_11852,N_10871,N_10361);
and U11853 (N_11853,N_10744,N_10879);
xnor U11854 (N_11854,N_10702,N_10838);
or U11855 (N_11855,N_10425,N_10914);
nand U11856 (N_11856,N_10111,N_10272);
nor U11857 (N_11857,N_10771,N_10732);
and U11858 (N_11858,N_10566,N_10873);
or U11859 (N_11859,N_10109,N_10204);
or U11860 (N_11860,N_10385,N_10830);
nor U11861 (N_11861,N_10066,N_10018);
or U11862 (N_11862,N_10149,N_10557);
xnor U11863 (N_11863,N_10635,N_10575);
or U11864 (N_11864,N_10587,N_10614);
xnor U11865 (N_11865,N_10661,N_10436);
xnor U11866 (N_11866,N_10040,N_10094);
or U11867 (N_11867,N_10060,N_10098);
nor U11868 (N_11868,N_10799,N_10383);
and U11869 (N_11869,N_10878,N_10769);
nand U11870 (N_11870,N_10912,N_10661);
nand U11871 (N_11871,N_10883,N_10684);
or U11872 (N_11872,N_10482,N_10955);
nor U11873 (N_11873,N_10076,N_10010);
and U11874 (N_11874,N_10708,N_10743);
and U11875 (N_11875,N_10489,N_10938);
xnor U11876 (N_11876,N_10555,N_10980);
and U11877 (N_11877,N_10669,N_10626);
nand U11878 (N_11878,N_10219,N_10817);
and U11879 (N_11879,N_10473,N_10684);
nor U11880 (N_11880,N_10841,N_10507);
nor U11881 (N_11881,N_10445,N_10743);
nand U11882 (N_11882,N_10084,N_10912);
and U11883 (N_11883,N_10131,N_10297);
or U11884 (N_11884,N_10688,N_10509);
nor U11885 (N_11885,N_10819,N_10208);
and U11886 (N_11886,N_10279,N_10614);
xor U11887 (N_11887,N_10902,N_10325);
and U11888 (N_11888,N_10391,N_10987);
nand U11889 (N_11889,N_10580,N_10154);
nand U11890 (N_11890,N_10382,N_10703);
nor U11891 (N_11891,N_10475,N_10917);
xor U11892 (N_11892,N_10692,N_10750);
nand U11893 (N_11893,N_10059,N_10479);
and U11894 (N_11894,N_10203,N_10130);
or U11895 (N_11895,N_10190,N_10663);
and U11896 (N_11896,N_10097,N_10812);
nor U11897 (N_11897,N_10076,N_10868);
nand U11898 (N_11898,N_10020,N_10486);
xnor U11899 (N_11899,N_10980,N_10316);
or U11900 (N_11900,N_10003,N_10335);
or U11901 (N_11901,N_10721,N_10821);
or U11902 (N_11902,N_10616,N_10321);
and U11903 (N_11903,N_10577,N_10152);
and U11904 (N_11904,N_10206,N_10389);
or U11905 (N_11905,N_10811,N_10206);
nand U11906 (N_11906,N_10983,N_10244);
nor U11907 (N_11907,N_10868,N_10036);
xnor U11908 (N_11908,N_10140,N_10242);
nand U11909 (N_11909,N_10044,N_10225);
nand U11910 (N_11910,N_10341,N_10023);
and U11911 (N_11911,N_10424,N_10445);
and U11912 (N_11912,N_10681,N_10236);
xnor U11913 (N_11913,N_10203,N_10059);
xnor U11914 (N_11914,N_10064,N_10180);
nand U11915 (N_11915,N_10854,N_10154);
nand U11916 (N_11916,N_10290,N_10763);
or U11917 (N_11917,N_10872,N_10560);
and U11918 (N_11918,N_10124,N_10397);
and U11919 (N_11919,N_10207,N_10648);
nand U11920 (N_11920,N_10337,N_10856);
or U11921 (N_11921,N_10196,N_10225);
or U11922 (N_11922,N_10011,N_10022);
xnor U11923 (N_11923,N_10459,N_10168);
or U11924 (N_11924,N_10536,N_10170);
nand U11925 (N_11925,N_10373,N_10901);
and U11926 (N_11926,N_10490,N_10295);
or U11927 (N_11927,N_10753,N_10116);
nand U11928 (N_11928,N_10423,N_10173);
or U11929 (N_11929,N_10127,N_10089);
or U11930 (N_11930,N_10938,N_10319);
xor U11931 (N_11931,N_10251,N_10635);
nor U11932 (N_11932,N_10130,N_10826);
xor U11933 (N_11933,N_10169,N_10887);
xnor U11934 (N_11934,N_10507,N_10457);
xnor U11935 (N_11935,N_10940,N_10177);
or U11936 (N_11936,N_10846,N_10471);
xor U11937 (N_11937,N_10354,N_10517);
xnor U11938 (N_11938,N_10520,N_10669);
or U11939 (N_11939,N_10485,N_10697);
nand U11940 (N_11940,N_10645,N_10876);
or U11941 (N_11941,N_10205,N_10260);
nor U11942 (N_11942,N_10313,N_10642);
nor U11943 (N_11943,N_10827,N_10987);
nor U11944 (N_11944,N_10686,N_10028);
or U11945 (N_11945,N_10308,N_10794);
nand U11946 (N_11946,N_10242,N_10560);
and U11947 (N_11947,N_10616,N_10344);
or U11948 (N_11948,N_10328,N_10410);
nor U11949 (N_11949,N_10621,N_10507);
or U11950 (N_11950,N_10752,N_10308);
nor U11951 (N_11951,N_10984,N_10045);
and U11952 (N_11952,N_10725,N_10113);
nor U11953 (N_11953,N_10664,N_10520);
nor U11954 (N_11954,N_10841,N_10409);
xnor U11955 (N_11955,N_10318,N_10345);
nand U11956 (N_11956,N_10434,N_10136);
and U11957 (N_11957,N_10290,N_10839);
nor U11958 (N_11958,N_10450,N_10173);
nor U11959 (N_11959,N_10688,N_10749);
xnor U11960 (N_11960,N_10478,N_10416);
xor U11961 (N_11961,N_10254,N_10409);
xnor U11962 (N_11962,N_10731,N_10319);
or U11963 (N_11963,N_10200,N_10987);
or U11964 (N_11964,N_10396,N_10294);
xor U11965 (N_11965,N_10556,N_10792);
or U11966 (N_11966,N_10472,N_10416);
nor U11967 (N_11967,N_10226,N_10182);
nand U11968 (N_11968,N_10212,N_10617);
xnor U11969 (N_11969,N_10911,N_10106);
xnor U11970 (N_11970,N_10711,N_10968);
xnor U11971 (N_11971,N_10388,N_10514);
xor U11972 (N_11972,N_10463,N_10870);
nor U11973 (N_11973,N_10084,N_10685);
or U11974 (N_11974,N_10828,N_10989);
and U11975 (N_11975,N_10420,N_10644);
nor U11976 (N_11976,N_10336,N_10684);
xnor U11977 (N_11977,N_10237,N_10059);
or U11978 (N_11978,N_10263,N_10523);
or U11979 (N_11979,N_10669,N_10653);
xor U11980 (N_11980,N_10434,N_10835);
and U11981 (N_11981,N_10587,N_10740);
and U11982 (N_11982,N_10134,N_10237);
nand U11983 (N_11983,N_10039,N_10047);
and U11984 (N_11984,N_10515,N_10958);
nand U11985 (N_11985,N_10729,N_10455);
nand U11986 (N_11986,N_10682,N_10239);
or U11987 (N_11987,N_10520,N_10752);
nand U11988 (N_11988,N_10811,N_10205);
or U11989 (N_11989,N_10083,N_10335);
nor U11990 (N_11990,N_10358,N_10961);
xor U11991 (N_11991,N_10914,N_10864);
nor U11992 (N_11992,N_10679,N_10924);
nor U11993 (N_11993,N_10116,N_10497);
nor U11994 (N_11994,N_10066,N_10173);
xnor U11995 (N_11995,N_10272,N_10441);
or U11996 (N_11996,N_10264,N_10132);
or U11997 (N_11997,N_10217,N_10100);
and U11998 (N_11998,N_10230,N_10818);
xnor U11999 (N_11999,N_10829,N_10868);
nor U12000 (N_12000,N_11174,N_11398);
or U12001 (N_12001,N_11956,N_11449);
xor U12002 (N_12002,N_11851,N_11202);
xnor U12003 (N_12003,N_11512,N_11235);
or U12004 (N_12004,N_11876,N_11704);
nor U12005 (N_12005,N_11056,N_11326);
and U12006 (N_12006,N_11253,N_11290);
and U12007 (N_12007,N_11085,N_11979);
or U12008 (N_12008,N_11213,N_11858);
nand U12009 (N_12009,N_11030,N_11259);
and U12010 (N_12010,N_11924,N_11570);
and U12011 (N_12011,N_11342,N_11165);
or U12012 (N_12012,N_11629,N_11505);
xor U12013 (N_12013,N_11172,N_11591);
and U12014 (N_12014,N_11830,N_11674);
nand U12015 (N_12015,N_11655,N_11353);
xnor U12016 (N_12016,N_11076,N_11643);
or U12017 (N_12017,N_11513,N_11891);
xor U12018 (N_12018,N_11660,N_11573);
or U12019 (N_12019,N_11256,N_11820);
and U12020 (N_12020,N_11278,N_11321);
xor U12021 (N_12021,N_11315,N_11528);
nand U12022 (N_12022,N_11988,N_11776);
nor U12023 (N_12023,N_11019,N_11833);
nor U12024 (N_12024,N_11641,N_11507);
xor U12025 (N_12025,N_11821,N_11031);
or U12026 (N_12026,N_11116,N_11407);
and U12027 (N_12027,N_11542,N_11497);
nor U12028 (N_12028,N_11831,N_11049);
or U12029 (N_12029,N_11471,N_11195);
and U12030 (N_12030,N_11399,N_11878);
or U12031 (N_12031,N_11244,N_11420);
xor U12032 (N_12032,N_11596,N_11144);
xnor U12033 (N_12033,N_11285,N_11658);
nand U12034 (N_12034,N_11852,N_11167);
xor U12035 (N_12035,N_11684,N_11675);
and U12036 (N_12036,N_11870,N_11091);
xor U12037 (N_12037,N_11063,N_11179);
or U12038 (N_12038,N_11775,N_11487);
xor U12039 (N_12039,N_11912,N_11142);
xor U12040 (N_12040,N_11316,N_11584);
nor U12041 (N_12041,N_11535,N_11360);
or U12042 (N_12042,N_11271,N_11110);
or U12043 (N_12043,N_11077,N_11927);
nand U12044 (N_12044,N_11306,N_11223);
and U12045 (N_12045,N_11765,N_11672);
nor U12046 (N_12046,N_11245,N_11190);
nor U12047 (N_12047,N_11712,N_11274);
nor U12048 (N_12048,N_11896,N_11883);
nand U12049 (N_12049,N_11414,N_11620);
nand U12050 (N_12050,N_11583,N_11832);
nand U12051 (N_12051,N_11595,N_11022);
or U12052 (N_12052,N_11818,N_11416);
or U12053 (N_12053,N_11539,N_11518);
nand U12054 (N_12054,N_11226,N_11037);
or U12055 (N_12055,N_11649,N_11705);
and U12056 (N_12056,N_11286,N_11889);
nor U12057 (N_12057,N_11425,N_11255);
nand U12058 (N_12058,N_11756,N_11141);
xnor U12059 (N_12059,N_11132,N_11622);
or U12060 (N_12060,N_11483,N_11710);
and U12061 (N_12061,N_11923,N_11362);
nand U12062 (N_12062,N_11764,N_11992);
nor U12063 (N_12063,N_11797,N_11397);
xor U12064 (N_12064,N_11948,N_11721);
xor U12065 (N_12065,N_11603,N_11667);
or U12066 (N_12066,N_11514,N_11719);
nand U12067 (N_12067,N_11477,N_11955);
or U12068 (N_12068,N_11718,N_11531);
or U12069 (N_12069,N_11947,N_11970);
nand U12070 (N_12070,N_11178,N_11388);
and U12071 (N_12071,N_11033,N_11478);
and U12072 (N_12072,N_11578,N_11925);
xor U12073 (N_12073,N_11104,N_11099);
xor U12074 (N_12074,N_11799,N_11608);
nand U12075 (N_12075,N_11424,N_11351);
or U12076 (N_12076,N_11900,N_11673);
nand U12077 (N_12077,N_11224,N_11920);
and U12078 (N_12078,N_11034,N_11100);
nand U12079 (N_12079,N_11565,N_11810);
or U12080 (N_12080,N_11071,N_11793);
and U12081 (N_12081,N_11273,N_11358);
nand U12082 (N_12082,N_11913,N_11731);
and U12083 (N_12083,N_11191,N_11472);
and U12084 (N_12084,N_11128,N_11587);
or U12085 (N_12085,N_11630,N_11111);
nand U12086 (N_12086,N_11521,N_11205);
or U12087 (N_12087,N_11064,N_11936);
or U12088 (N_12088,N_11046,N_11052);
or U12089 (N_12089,N_11967,N_11024);
nor U12090 (N_12090,N_11002,N_11401);
nand U12091 (N_12091,N_11289,N_11383);
or U12092 (N_12092,N_11059,N_11386);
or U12093 (N_12093,N_11232,N_11768);
xor U12094 (N_12094,N_11231,N_11310);
nand U12095 (N_12095,N_11998,N_11341);
nand U12096 (N_12096,N_11537,N_11060);
xor U12097 (N_12097,N_11784,N_11840);
xor U12098 (N_12098,N_11709,N_11816);
or U12099 (N_12099,N_11160,N_11857);
nand U12100 (N_12100,N_11708,N_11156);
nor U12101 (N_12101,N_11189,N_11020);
nand U12102 (N_12102,N_11890,N_11429);
nor U12103 (N_12103,N_11503,N_11538);
and U12104 (N_12104,N_11227,N_11623);
nand U12105 (N_12105,N_11819,N_11216);
nor U12106 (N_12106,N_11124,N_11467);
and U12107 (N_12107,N_11453,N_11139);
and U12108 (N_12108,N_11795,N_11934);
nor U12109 (N_12109,N_11976,N_11087);
nor U12110 (N_12110,N_11714,N_11645);
nor U12111 (N_12111,N_11119,N_11355);
and U12112 (N_12112,N_11444,N_11657);
nor U12113 (N_12113,N_11009,N_11464);
and U12114 (N_12114,N_11781,N_11592);
or U12115 (N_12115,N_11096,N_11092);
and U12116 (N_12116,N_11347,N_11440);
xor U12117 (N_12117,N_11328,N_11045);
or U12118 (N_12118,N_11579,N_11729);
and U12119 (N_12119,N_11805,N_11669);
xnor U12120 (N_12120,N_11665,N_11715);
xor U12121 (N_12121,N_11484,N_11939);
and U12122 (N_12122,N_11602,N_11391);
and U12123 (N_12123,N_11626,N_11114);
nor U12124 (N_12124,N_11375,N_11677);
and U12125 (N_12125,N_11058,N_11417);
or U12126 (N_12126,N_11777,N_11412);
or U12127 (N_12127,N_11220,N_11447);
nand U12128 (N_12128,N_11745,N_11576);
xnor U12129 (N_12129,N_11861,N_11217);
nand U12130 (N_12130,N_11164,N_11308);
nand U12131 (N_12131,N_11280,N_11561);
nor U12132 (N_12132,N_11396,N_11894);
nor U12133 (N_12133,N_11943,N_11778);
and U12134 (N_12134,N_11711,N_11498);
nand U12135 (N_12135,N_11057,N_11722);
and U12136 (N_12136,N_11515,N_11549);
nand U12137 (N_12137,N_11126,N_11061);
nand U12138 (N_12138,N_11887,N_11905);
nor U12139 (N_12139,N_11148,N_11571);
nor U12140 (N_12140,N_11109,N_11086);
or U12141 (N_12141,N_11314,N_11094);
nor U12142 (N_12142,N_11615,N_11567);
or U12143 (N_12143,N_11480,N_11185);
or U12144 (N_12144,N_11001,N_11929);
nand U12145 (N_12145,N_11661,N_11406);
or U12146 (N_12146,N_11368,N_11225);
or U12147 (N_12147,N_11517,N_11525);
nand U12148 (N_12148,N_11390,N_11151);
nor U12149 (N_12149,N_11730,N_11664);
or U12150 (N_12150,N_11311,N_11983);
and U12151 (N_12151,N_11619,N_11656);
xnor U12152 (N_12152,N_11757,N_11131);
and U12153 (N_12153,N_11874,N_11122);
nor U12154 (N_12154,N_11859,N_11736);
xor U12155 (N_12155,N_11917,N_11825);
nor U12156 (N_12156,N_11690,N_11735);
xor U12157 (N_12157,N_11125,N_11192);
nor U12158 (N_12158,N_11356,N_11526);
xor U12159 (N_12159,N_11999,N_11760);
or U12160 (N_12160,N_11828,N_11695);
nand U12161 (N_12161,N_11845,N_11968);
xnor U12162 (N_12162,N_11115,N_11215);
nand U12163 (N_12163,N_11284,N_11794);
nor U12164 (N_12164,N_11903,N_11324);
nand U12165 (N_12165,N_11588,N_11204);
xnor U12166 (N_12166,N_11636,N_11250);
nand U12167 (N_12167,N_11370,N_11670);
or U12168 (N_12168,N_11717,N_11826);
or U12169 (N_12169,N_11260,N_11303);
and U12170 (N_12170,N_11624,N_11050);
xor U12171 (N_12171,N_11837,N_11486);
or U12172 (N_12172,N_11236,N_11036);
nor U12173 (N_12173,N_11646,N_11532);
or U12174 (N_12174,N_11302,N_11989);
nand U12175 (N_12175,N_11634,N_11411);
xor U12176 (N_12176,N_11650,N_11519);
nand U12177 (N_12177,N_11864,N_11162);
nor U12178 (N_12178,N_11047,N_11027);
and U12179 (N_12179,N_11696,N_11753);
nor U12180 (N_12180,N_11644,N_11774);
nand U12181 (N_12181,N_11072,N_11582);
nand U12182 (N_12182,N_11221,N_11240);
nor U12183 (N_12183,N_11985,N_11405);
nor U12184 (N_12184,N_11557,N_11129);
nor U12185 (N_12185,N_11380,N_11566);
xnor U12186 (N_12186,N_11332,N_11612);
xor U12187 (N_12187,N_11465,N_11454);
and U12188 (N_12188,N_11491,N_11233);
nand U12189 (N_12189,N_11038,N_11367);
and U12190 (N_12190,N_11065,N_11938);
nor U12191 (N_12191,N_11522,N_11694);
xor U12192 (N_12192,N_11436,N_11434);
xnor U12193 (N_12193,N_11680,N_11427);
nor U12194 (N_12194,N_11627,N_11208);
and U12195 (N_12195,N_11536,N_11752);
and U12196 (N_12196,N_11960,N_11201);
or U12197 (N_12197,N_11652,N_11014);
xor U12198 (N_12198,N_11373,N_11010);
xnor U12199 (N_12199,N_11006,N_11868);
nor U12200 (N_12200,N_11855,N_11758);
or U12201 (N_12201,N_11210,N_11163);
and U12202 (N_12202,N_11237,N_11902);
or U12203 (N_12203,N_11681,N_11432);
nor U12204 (N_12204,N_11371,N_11150);
nand U12205 (N_12205,N_11206,N_11155);
or U12206 (N_12206,N_11666,N_11873);
nand U12207 (N_12207,N_11222,N_11331);
nor U12208 (N_12208,N_11564,N_11127);
and U12209 (N_12209,N_11972,N_11343);
or U12210 (N_12210,N_11796,N_11823);
and U12211 (N_12211,N_11435,N_11980);
xor U12212 (N_12212,N_11838,N_11700);
nand U12213 (N_12213,N_11248,N_11662);
and U12214 (N_12214,N_11850,N_11214);
and U12215 (N_12215,N_11184,N_11942);
nand U12216 (N_12216,N_11008,N_11523);
xor U12217 (N_12217,N_11910,N_11707);
xnor U12218 (N_12218,N_11875,N_11813);
nor U12219 (N_12219,N_11246,N_11978);
xnor U12220 (N_12220,N_11292,N_11767);
or U12221 (N_12221,N_11597,N_11323);
or U12222 (N_12222,N_11703,N_11806);
nor U12223 (N_12223,N_11527,N_11490);
or U12224 (N_12224,N_11384,N_11392);
nor U12225 (N_12225,N_11926,N_11935);
nor U12226 (N_12226,N_11070,N_11581);
or U12227 (N_12227,N_11689,N_11346);
nor U12228 (N_12228,N_11611,N_11473);
xor U12229 (N_12229,N_11642,N_11639);
nor U12230 (N_12230,N_11180,N_11211);
and U12231 (N_12231,N_11198,N_11575);
and U12232 (N_12232,N_11594,N_11005);
xor U12233 (N_12233,N_11339,N_11726);
nor U12234 (N_12234,N_11754,N_11789);
or U12235 (N_12235,N_11866,N_11461);
nor U12236 (N_12236,N_11511,N_11916);
or U12237 (N_12237,N_11991,N_11013);
or U12238 (N_12238,N_11157,N_11106);
nand U12239 (N_12239,N_11802,N_11145);
nand U12240 (N_12240,N_11450,N_11430);
or U12241 (N_12241,N_11170,N_11648);
or U12242 (N_12242,N_11599,N_11755);
or U12243 (N_12243,N_11904,N_11888);
nor U12244 (N_12244,N_11548,N_11906);
nand U12245 (N_12245,N_11247,N_11400);
nor U12246 (N_12246,N_11785,N_11552);
and U12247 (N_12247,N_11319,N_11137);
xnor U12248 (N_12248,N_11640,N_11897);
nand U12249 (N_12249,N_11554,N_11843);
nand U12250 (N_12250,N_11188,N_11084);
nand U12251 (N_12251,N_11974,N_11335);
and U12252 (N_12252,N_11228,N_11618);
nor U12253 (N_12253,N_11885,N_11628);
and U12254 (N_12254,N_11848,N_11817);
and U12255 (N_12255,N_11918,N_11836);
or U12256 (N_12256,N_11361,N_11293);
xnor U12257 (N_12257,N_11196,N_11422);
nor U12258 (N_12258,N_11732,N_11078);
nand U12259 (N_12259,N_11423,N_11919);
or U12260 (N_12260,N_11871,N_11746);
or U12261 (N_12261,N_11500,N_11701);
nor U12262 (N_12262,N_11359,N_11408);
nand U12263 (N_12263,N_11699,N_11495);
nand U12264 (N_12264,N_11230,N_11476);
nor U12265 (N_12265,N_11856,N_11993);
nor U12266 (N_12266,N_11772,N_11418);
or U12267 (N_12267,N_11479,N_11882);
nor U12268 (N_12268,N_11931,N_11012);
or U12269 (N_12269,N_11915,N_11908);
xor U12270 (N_12270,N_11963,N_11252);
nor U12271 (N_12271,N_11168,N_11249);
nand U12272 (N_12272,N_11763,N_11466);
nor U12273 (N_12273,N_11283,N_11445);
and U12274 (N_12274,N_11385,N_11089);
or U12275 (N_12275,N_11130,N_11040);
and U12276 (N_12276,N_11769,N_11748);
or U12277 (N_12277,N_11770,N_11562);
nor U12278 (N_12278,N_11744,N_11379);
nor U12279 (N_12279,N_11580,N_11835);
or U12280 (N_12280,N_11693,N_11724);
and U12281 (N_12281,N_11067,N_11166);
xnor U12282 (N_12282,N_11780,N_11605);
or U12283 (N_12283,N_11138,N_11725);
xnor U12284 (N_12284,N_11766,N_11510);
or U12285 (N_12285,N_11295,N_11553);
nand U12286 (N_12286,N_11529,N_11463);
and U12287 (N_12287,N_11140,N_11382);
or U12288 (N_12288,N_11403,N_11493);
or U12289 (N_12289,N_11563,N_11687);
nand U12290 (N_12290,N_11409,N_11374);
or U12291 (N_12291,N_11804,N_11921);
nor U12292 (N_12292,N_11598,N_11637);
nor U12293 (N_12293,N_11307,N_11042);
nand U12294 (N_12294,N_11426,N_11183);
nor U12295 (N_12295,N_11496,N_11073);
xnor U12296 (N_12296,N_11811,N_11325);
and U12297 (N_12297,N_11986,N_11606);
nor U12298 (N_12298,N_11800,N_11349);
nor U12299 (N_12299,N_11585,N_11499);
xor U12300 (N_12300,N_11199,N_11081);
and U12301 (N_12301,N_11683,N_11969);
or U12302 (N_12302,N_11069,N_11621);
xnor U12303 (N_12303,N_11004,N_11834);
xor U12304 (N_12304,N_11886,N_11305);
and U12305 (N_12305,N_11740,N_11193);
or U12306 (N_12306,N_11809,N_11241);
and U12307 (N_12307,N_11443,N_11485);
and U12308 (N_12308,N_11458,N_11387);
nor U12309 (N_12309,N_11299,N_11761);
or U12310 (N_12310,N_11304,N_11279);
nand U12311 (N_12311,N_11879,N_11294);
nand U12312 (N_12312,N_11750,N_11997);
xor U12313 (N_12313,N_11686,N_11971);
or U12314 (N_12314,N_11265,N_11982);
nand U12315 (N_12315,N_11317,N_11338);
nand U12316 (N_12316,N_11363,N_11134);
nor U12317 (N_12317,N_11448,N_11632);
nand U12318 (N_12318,N_11402,N_11782);
nand U12319 (N_12319,N_11635,N_11186);
or U12320 (N_12320,N_11459,N_11945);
or U12321 (N_12321,N_11203,N_11558);
nor U12322 (N_12322,N_11301,N_11079);
nor U12323 (N_12323,N_11762,N_11437);
nand U12324 (N_12324,N_11147,N_11082);
or U12325 (N_12325,N_11101,N_11136);
or U12326 (N_12326,N_11966,N_11692);
nor U12327 (N_12327,N_11815,N_11559);
nand U12328 (N_12328,N_11357,N_11604);
xnor U12329 (N_12329,N_11187,N_11759);
nor U12330 (N_12330,N_11270,N_11209);
nand U12331 (N_12331,N_11197,N_11288);
nand U12332 (N_12332,N_11007,N_11261);
xor U12333 (N_12333,N_11275,N_11039);
xor U12334 (N_12334,N_11442,N_11880);
nand U12335 (N_12335,N_11653,N_11613);
nand U12336 (N_12336,N_11572,N_11625);
and U12337 (N_12337,N_11957,N_11439);
and U12338 (N_12338,N_11313,N_11120);
nor U12339 (N_12339,N_11928,N_11600);
nor U12340 (N_12340,N_11741,N_11108);
and U12341 (N_12341,N_11702,N_11869);
and U12342 (N_12342,N_11159,N_11395);
or U12343 (N_12343,N_11451,N_11533);
or U12344 (N_12344,N_11053,N_11909);
nor U12345 (N_12345,N_11987,N_11258);
nor U12346 (N_12346,N_11846,N_11456);
nor U12347 (N_12347,N_11631,N_11952);
nor U12348 (N_12348,N_11678,N_11739);
and U12349 (N_12349,N_11685,N_11277);
and U12350 (N_12350,N_11854,N_11556);
or U12351 (N_12351,N_11751,N_11000);
or U12352 (N_12352,N_11021,N_11475);
and U12353 (N_12353,N_11062,N_11207);
and U12354 (N_12354,N_11893,N_11043);
xnor U12355 (N_12355,N_11614,N_11616);
and U12356 (N_12356,N_11494,N_11177);
nor U12357 (N_12357,N_11508,N_11105);
or U12358 (N_12358,N_11899,N_11468);
or U12359 (N_12359,N_11333,N_11814);
nor U12360 (N_12360,N_11786,N_11352);
and U12361 (N_12361,N_11822,N_11041);
or U12362 (N_12362,N_11118,N_11638);
or U12363 (N_12363,N_11066,N_11176);
nor U12364 (N_12364,N_11698,N_11433);
and U12365 (N_12365,N_11953,N_11849);
and U12366 (N_12366,N_11791,N_11334);
nand U12367 (N_12367,N_11103,N_11950);
or U12368 (N_12368,N_11607,N_11327);
and U12369 (N_12369,N_11182,N_11016);
and U12370 (N_12370,N_11080,N_11263);
and U12371 (N_12371,N_11545,N_11842);
or U12372 (N_12372,N_11941,N_11404);
nor U12373 (N_12373,N_11287,N_11577);
nand U12374 (N_12374,N_11509,N_11441);
nand U12375 (N_12375,N_11254,N_11268);
and U12376 (N_12376,N_11011,N_11589);
nor U12377 (N_12377,N_11149,N_11133);
or U12378 (N_12378,N_11200,N_11798);
and U12379 (N_12379,N_11194,N_11394);
nor U12380 (N_12380,N_11291,N_11117);
or U12381 (N_12381,N_11516,N_11651);
and U12382 (N_12382,N_11098,N_11282);
or U12383 (N_12383,N_11269,N_11853);
xor U12384 (N_12384,N_11410,N_11469);
nand U12385 (N_12385,N_11075,N_11348);
xor U12386 (N_12386,N_11029,N_11297);
and U12387 (N_12387,N_11990,N_11543);
nor U12388 (N_12388,N_11713,N_11015);
xor U12389 (N_12389,N_11337,N_11095);
xnor U12390 (N_12390,N_11551,N_11457);
nand U12391 (N_12391,N_11276,N_11884);
xor U12392 (N_12392,N_11381,N_11944);
nor U12393 (N_12393,N_11593,N_11296);
or U12394 (N_12394,N_11995,N_11688);
or U12395 (N_12395,N_11749,N_11462);
or U12396 (N_12396,N_11309,N_11173);
nor U12397 (N_12397,N_11940,N_11787);
or U12398 (N_12398,N_11738,N_11419);
xor U12399 (N_12399,N_11679,N_11068);
xor U12400 (N_12400,N_11720,N_11003);
xor U12401 (N_12401,N_11074,N_11329);
xnor U12402 (N_12402,N_11312,N_11017);
and U12403 (N_12403,N_11369,N_11376);
xor U12404 (N_12404,N_11504,N_11262);
nand U12405 (N_12405,N_11340,N_11320);
nor U12406 (N_12406,N_11937,N_11994);
nor U12407 (N_12407,N_11898,N_11169);
or U12408 (N_12408,N_11264,N_11460);
nand U12409 (N_12409,N_11336,N_11266);
nand U12410 (N_12410,N_11298,N_11737);
nor U12411 (N_12411,N_11901,N_11839);
nor U12412 (N_12412,N_11048,N_11421);
nand U12413 (N_12413,N_11365,N_11474);
xor U12414 (N_12414,N_11984,N_11668);
or U12415 (N_12415,N_11803,N_11438);
nand U12416 (N_12416,N_11452,N_11455);
and U12417 (N_12417,N_11171,N_11844);
or U12418 (N_12418,N_11257,N_11143);
nand U12419 (N_12419,N_11026,N_11601);
and U12420 (N_12420,N_11088,N_11470);
or U12421 (N_12421,N_11975,N_11541);
nand U12422 (N_12422,N_11107,N_11790);
nand U12423 (N_12423,N_11932,N_11728);
or U12424 (N_12424,N_11959,N_11716);
or U12425 (N_12425,N_11907,N_11647);
or U12426 (N_12426,N_11372,N_11102);
and U12427 (N_12427,N_11659,N_11771);
xor U12428 (N_12428,N_11862,N_11446);
nor U12429 (N_12429,N_11550,N_11218);
nand U12430 (N_12430,N_11860,N_11083);
nor U12431 (N_12431,N_11779,N_11364);
xor U12432 (N_12432,N_11530,N_11028);
or U12433 (N_12433,N_11281,N_11238);
xnor U12434 (N_12434,N_11534,N_11773);
nand U12435 (N_12435,N_11792,N_11502);
or U12436 (N_12436,N_11682,N_11824);
xor U12437 (N_12437,N_11949,N_11933);
nand U12438 (N_12438,N_11590,N_11267);
nor U12439 (N_12439,N_11243,N_11481);
nor U12440 (N_12440,N_11054,N_11234);
xnor U12441 (N_12441,N_11951,N_11569);
nand U12442 (N_12442,N_11946,N_11733);
and U12443 (N_12443,N_11175,N_11242);
xor U12444 (N_12444,N_11153,N_11930);
xnor U12445 (N_12445,N_11586,N_11025);
nand U12446 (N_12446,N_11097,N_11251);
nand U12447 (N_12447,N_11783,N_11377);
nand U12448 (N_12448,N_11892,N_11996);
nand U12449 (N_12449,N_11568,N_11807);
or U12450 (N_12450,N_11706,N_11318);
and U12451 (N_12451,N_11506,N_11389);
xor U12452 (N_12452,N_11964,N_11788);
and U12453 (N_12453,N_11547,N_11727);
nand U12454 (N_12454,N_11872,N_11428);
nor U12455 (N_12455,N_11121,N_11239);
nand U12456 (N_12456,N_11123,N_11691);
xor U12457 (N_12457,N_11090,N_11492);
or U12458 (N_12458,N_11841,N_11415);
nor U12459 (N_12459,N_11546,N_11112);
or U12460 (N_12460,N_11610,N_11847);
or U12461 (N_12461,N_11544,N_11366);
and U12462 (N_12462,N_11431,N_11023);
nor U12463 (N_12463,N_11609,N_11161);
nor U12464 (N_12464,N_11973,N_11865);
or U12465 (N_12465,N_11914,N_11158);
nor U12466 (N_12466,N_11734,N_11093);
or U12467 (N_12467,N_11676,N_11488);
nand U12468 (N_12468,N_11962,N_11867);
and U12469 (N_12469,N_11300,N_11654);
and U12470 (N_12470,N_11965,N_11354);
xor U12471 (N_12471,N_11018,N_11330);
nor U12472 (N_12472,N_11345,N_11344);
or U12473 (N_12473,N_11743,N_11981);
nand U12474 (N_12474,N_11219,N_11617);
or U12475 (N_12475,N_11958,N_11035);
xor U12476 (N_12476,N_11113,N_11742);
xnor U12477 (N_12477,N_11135,N_11413);
xor U12478 (N_12478,N_11482,N_11146);
nand U12479 (N_12479,N_11378,N_11152);
xor U12480 (N_12480,N_11633,N_11827);
nand U12481 (N_12481,N_11922,N_11489);
nand U12482 (N_12482,N_11032,N_11272);
nor U12483 (N_12483,N_11229,N_11954);
nor U12484 (N_12484,N_11829,N_11555);
and U12485 (N_12485,N_11524,N_11723);
xnor U12486 (N_12486,N_11801,N_11911);
or U12487 (N_12487,N_11560,N_11540);
and U12488 (N_12488,N_11747,N_11977);
nand U12489 (N_12489,N_11881,N_11322);
xor U12490 (N_12490,N_11154,N_11044);
nor U12491 (N_12491,N_11671,N_11350);
and U12492 (N_12492,N_11877,N_11895);
or U12493 (N_12493,N_11574,N_11212);
xnor U12494 (N_12494,N_11520,N_11051);
nand U12495 (N_12495,N_11697,N_11055);
or U12496 (N_12496,N_11812,N_11501);
xor U12497 (N_12497,N_11393,N_11863);
and U12498 (N_12498,N_11961,N_11663);
and U12499 (N_12499,N_11181,N_11808);
nor U12500 (N_12500,N_11508,N_11097);
and U12501 (N_12501,N_11187,N_11683);
nor U12502 (N_12502,N_11852,N_11845);
xor U12503 (N_12503,N_11479,N_11320);
xnor U12504 (N_12504,N_11673,N_11622);
nand U12505 (N_12505,N_11985,N_11238);
xnor U12506 (N_12506,N_11484,N_11327);
nand U12507 (N_12507,N_11971,N_11244);
nand U12508 (N_12508,N_11668,N_11301);
or U12509 (N_12509,N_11056,N_11032);
nand U12510 (N_12510,N_11396,N_11981);
xnor U12511 (N_12511,N_11744,N_11898);
xnor U12512 (N_12512,N_11024,N_11625);
nor U12513 (N_12513,N_11476,N_11871);
and U12514 (N_12514,N_11344,N_11142);
nand U12515 (N_12515,N_11276,N_11331);
and U12516 (N_12516,N_11823,N_11105);
nand U12517 (N_12517,N_11807,N_11930);
and U12518 (N_12518,N_11593,N_11904);
and U12519 (N_12519,N_11115,N_11131);
nor U12520 (N_12520,N_11120,N_11389);
or U12521 (N_12521,N_11520,N_11595);
and U12522 (N_12522,N_11807,N_11679);
nand U12523 (N_12523,N_11876,N_11477);
xnor U12524 (N_12524,N_11061,N_11431);
or U12525 (N_12525,N_11254,N_11179);
and U12526 (N_12526,N_11812,N_11621);
xnor U12527 (N_12527,N_11671,N_11704);
or U12528 (N_12528,N_11078,N_11265);
nand U12529 (N_12529,N_11975,N_11007);
or U12530 (N_12530,N_11120,N_11103);
and U12531 (N_12531,N_11516,N_11841);
or U12532 (N_12532,N_11266,N_11409);
nand U12533 (N_12533,N_11531,N_11784);
nor U12534 (N_12534,N_11064,N_11674);
nand U12535 (N_12535,N_11032,N_11165);
or U12536 (N_12536,N_11924,N_11231);
nand U12537 (N_12537,N_11214,N_11744);
and U12538 (N_12538,N_11291,N_11982);
nor U12539 (N_12539,N_11310,N_11873);
xnor U12540 (N_12540,N_11149,N_11508);
or U12541 (N_12541,N_11947,N_11816);
nand U12542 (N_12542,N_11436,N_11025);
and U12543 (N_12543,N_11366,N_11636);
or U12544 (N_12544,N_11764,N_11892);
or U12545 (N_12545,N_11001,N_11516);
or U12546 (N_12546,N_11519,N_11513);
or U12547 (N_12547,N_11550,N_11805);
nor U12548 (N_12548,N_11894,N_11255);
or U12549 (N_12549,N_11668,N_11986);
xor U12550 (N_12550,N_11199,N_11184);
and U12551 (N_12551,N_11755,N_11908);
xnor U12552 (N_12552,N_11915,N_11314);
nand U12553 (N_12553,N_11187,N_11755);
and U12554 (N_12554,N_11966,N_11224);
xor U12555 (N_12555,N_11098,N_11573);
nor U12556 (N_12556,N_11167,N_11249);
xor U12557 (N_12557,N_11253,N_11367);
nand U12558 (N_12558,N_11303,N_11637);
xnor U12559 (N_12559,N_11459,N_11468);
nor U12560 (N_12560,N_11232,N_11432);
nand U12561 (N_12561,N_11933,N_11642);
nor U12562 (N_12562,N_11513,N_11976);
nor U12563 (N_12563,N_11098,N_11222);
nor U12564 (N_12564,N_11031,N_11989);
or U12565 (N_12565,N_11840,N_11685);
nor U12566 (N_12566,N_11134,N_11515);
or U12567 (N_12567,N_11140,N_11384);
nand U12568 (N_12568,N_11228,N_11890);
nor U12569 (N_12569,N_11766,N_11194);
xor U12570 (N_12570,N_11596,N_11031);
and U12571 (N_12571,N_11011,N_11259);
nor U12572 (N_12572,N_11377,N_11223);
or U12573 (N_12573,N_11127,N_11986);
and U12574 (N_12574,N_11112,N_11864);
nor U12575 (N_12575,N_11997,N_11792);
xor U12576 (N_12576,N_11215,N_11806);
xor U12577 (N_12577,N_11589,N_11655);
nor U12578 (N_12578,N_11929,N_11245);
xnor U12579 (N_12579,N_11678,N_11086);
or U12580 (N_12580,N_11499,N_11798);
and U12581 (N_12581,N_11572,N_11252);
and U12582 (N_12582,N_11887,N_11660);
or U12583 (N_12583,N_11707,N_11690);
xnor U12584 (N_12584,N_11923,N_11828);
or U12585 (N_12585,N_11753,N_11487);
nor U12586 (N_12586,N_11583,N_11162);
xnor U12587 (N_12587,N_11696,N_11949);
nand U12588 (N_12588,N_11009,N_11237);
or U12589 (N_12589,N_11633,N_11666);
nand U12590 (N_12590,N_11888,N_11130);
and U12591 (N_12591,N_11506,N_11498);
and U12592 (N_12592,N_11519,N_11740);
xnor U12593 (N_12593,N_11968,N_11143);
or U12594 (N_12594,N_11611,N_11287);
xnor U12595 (N_12595,N_11293,N_11376);
xnor U12596 (N_12596,N_11518,N_11234);
and U12597 (N_12597,N_11537,N_11055);
and U12598 (N_12598,N_11132,N_11056);
nor U12599 (N_12599,N_11385,N_11921);
nor U12600 (N_12600,N_11477,N_11324);
xnor U12601 (N_12601,N_11406,N_11703);
nand U12602 (N_12602,N_11068,N_11219);
nor U12603 (N_12603,N_11661,N_11808);
xnor U12604 (N_12604,N_11481,N_11223);
nor U12605 (N_12605,N_11306,N_11729);
nor U12606 (N_12606,N_11747,N_11552);
xnor U12607 (N_12607,N_11528,N_11764);
xnor U12608 (N_12608,N_11687,N_11424);
xor U12609 (N_12609,N_11886,N_11360);
and U12610 (N_12610,N_11615,N_11239);
nand U12611 (N_12611,N_11755,N_11917);
or U12612 (N_12612,N_11848,N_11759);
nor U12613 (N_12613,N_11101,N_11424);
nand U12614 (N_12614,N_11504,N_11746);
and U12615 (N_12615,N_11997,N_11935);
xor U12616 (N_12616,N_11106,N_11362);
nor U12617 (N_12617,N_11159,N_11762);
or U12618 (N_12618,N_11053,N_11890);
and U12619 (N_12619,N_11541,N_11436);
nand U12620 (N_12620,N_11378,N_11547);
xnor U12621 (N_12621,N_11118,N_11405);
or U12622 (N_12622,N_11387,N_11494);
and U12623 (N_12623,N_11180,N_11004);
and U12624 (N_12624,N_11163,N_11600);
and U12625 (N_12625,N_11641,N_11302);
xnor U12626 (N_12626,N_11102,N_11458);
xor U12627 (N_12627,N_11277,N_11754);
nand U12628 (N_12628,N_11399,N_11232);
xnor U12629 (N_12629,N_11226,N_11484);
xnor U12630 (N_12630,N_11842,N_11377);
or U12631 (N_12631,N_11024,N_11265);
nor U12632 (N_12632,N_11351,N_11335);
xnor U12633 (N_12633,N_11602,N_11006);
and U12634 (N_12634,N_11250,N_11738);
or U12635 (N_12635,N_11142,N_11454);
or U12636 (N_12636,N_11364,N_11652);
nand U12637 (N_12637,N_11989,N_11803);
or U12638 (N_12638,N_11301,N_11841);
nand U12639 (N_12639,N_11107,N_11584);
xnor U12640 (N_12640,N_11137,N_11259);
and U12641 (N_12641,N_11825,N_11356);
nand U12642 (N_12642,N_11452,N_11742);
nand U12643 (N_12643,N_11010,N_11408);
and U12644 (N_12644,N_11130,N_11399);
nor U12645 (N_12645,N_11574,N_11628);
or U12646 (N_12646,N_11177,N_11534);
nor U12647 (N_12647,N_11589,N_11995);
and U12648 (N_12648,N_11965,N_11386);
or U12649 (N_12649,N_11631,N_11331);
xor U12650 (N_12650,N_11276,N_11127);
and U12651 (N_12651,N_11451,N_11832);
nor U12652 (N_12652,N_11773,N_11343);
nor U12653 (N_12653,N_11527,N_11044);
xnor U12654 (N_12654,N_11700,N_11219);
nor U12655 (N_12655,N_11081,N_11698);
nor U12656 (N_12656,N_11459,N_11967);
and U12657 (N_12657,N_11274,N_11002);
or U12658 (N_12658,N_11873,N_11511);
or U12659 (N_12659,N_11988,N_11263);
nor U12660 (N_12660,N_11579,N_11931);
and U12661 (N_12661,N_11635,N_11633);
nand U12662 (N_12662,N_11612,N_11870);
nand U12663 (N_12663,N_11163,N_11763);
or U12664 (N_12664,N_11093,N_11002);
nand U12665 (N_12665,N_11297,N_11886);
or U12666 (N_12666,N_11841,N_11766);
xor U12667 (N_12667,N_11987,N_11567);
nor U12668 (N_12668,N_11816,N_11517);
and U12669 (N_12669,N_11083,N_11174);
xnor U12670 (N_12670,N_11727,N_11709);
nand U12671 (N_12671,N_11669,N_11177);
xor U12672 (N_12672,N_11181,N_11173);
or U12673 (N_12673,N_11629,N_11981);
nor U12674 (N_12674,N_11392,N_11858);
xor U12675 (N_12675,N_11686,N_11835);
nand U12676 (N_12676,N_11420,N_11904);
nor U12677 (N_12677,N_11754,N_11191);
and U12678 (N_12678,N_11646,N_11604);
nand U12679 (N_12679,N_11285,N_11619);
and U12680 (N_12680,N_11095,N_11698);
nand U12681 (N_12681,N_11307,N_11113);
and U12682 (N_12682,N_11251,N_11386);
nand U12683 (N_12683,N_11850,N_11435);
and U12684 (N_12684,N_11525,N_11914);
nor U12685 (N_12685,N_11225,N_11743);
or U12686 (N_12686,N_11183,N_11937);
and U12687 (N_12687,N_11112,N_11105);
and U12688 (N_12688,N_11562,N_11666);
nor U12689 (N_12689,N_11509,N_11675);
and U12690 (N_12690,N_11807,N_11024);
nand U12691 (N_12691,N_11548,N_11274);
nor U12692 (N_12692,N_11508,N_11927);
and U12693 (N_12693,N_11335,N_11067);
or U12694 (N_12694,N_11404,N_11287);
xnor U12695 (N_12695,N_11990,N_11769);
nand U12696 (N_12696,N_11523,N_11044);
or U12697 (N_12697,N_11937,N_11725);
xnor U12698 (N_12698,N_11118,N_11749);
or U12699 (N_12699,N_11807,N_11663);
nand U12700 (N_12700,N_11844,N_11643);
and U12701 (N_12701,N_11164,N_11596);
xor U12702 (N_12702,N_11978,N_11574);
or U12703 (N_12703,N_11696,N_11082);
nor U12704 (N_12704,N_11333,N_11657);
nand U12705 (N_12705,N_11919,N_11283);
xnor U12706 (N_12706,N_11754,N_11384);
and U12707 (N_12707,N_11630,N_11687);
and U12708 (N_12708,N_11077,N_11596);
or U12709 (N_12709,N_11514,N_11897);
and U12710 (N_12710,N_11594,N_11375);
and U12711 (N_12711,N_11087,N_11272);
or U12712 (N_12712,N_11730,N_11843);
nor U12713 (N_12713,N_11863,N_11638);
or U12714 (N_12714,N_11463,N_11066);
or U12715 (N_12715,N_11264,N_11409);
nand U12716 (N_12716,N_11178,N_11084);
or U12717 (N_12717,N_11912,N_11213);
nor U12718 (N_12718,N_11770,N_11112);
and U12719 (N_12719,N_11375,N_11491);
nand U12720 (N_12720,N_11495,N_11230);
and U12721 (N_12721,N_11317,N_11193);
xor U12722 (N_12722,N_11632,N_11340);
and U12723 (N_12723,N_11935,N_11664);
and U12724 (N_12724,N_11472,N_11174);
and U12725 (N_12725,N_11062,N_11971);
nor U12726 (N_12726,N_11859,N_11743);
nand U12727 (N_12727,N_11985,N_11429);
and U12728 (N_12728,N_11580,N_11849);
nor U12729 (N_12729,N_11147,N_11890);
or U12730 (N_12730,N_11894,N_11301);
or U12731 (N_12731,N_11741,N_11163);
or U12732 (N_12732,N_11414,N_11854);
xnor U12733 (N_12733,N_11513,N_11138);
and U12734 (N_12734,N_11999,N_11482);
xnor U12735 (N_12735,N_11884,N_11598);
and U12736 (N_12736,N_11167,N_11110);
nand U12737 (N_12737,N_11822,N_11133);
nand U12738 (N_12738,N_11246,N_11053);
nor U12739 (N_12739,N_11894,N_11386);
nor U12740 (N_12740,N_11936,N_11542);
nor U12741 (N_12741,N_11249,N_11779);
and U12742 (N_12742,N_11218,N_11488);
and U12743 (N_12743,N_11768,N_11316);
and U12744 (N_12744,N_11243,N_11458);
nor U12745 (N_12745,N_11677,N_11206);
nor U12746 (N_12746,N_11009,N_11961);
nand U12747 (N_12747,N_11154,N_11070);
or U12748 (N_12748,N_11939,N_11788);
or U12749 (N_12749,N_11616,N_11873);
and U12750 (N_12750,N_11786,N_11812);
and U12751 (N_12751,N_11664,N_11060);
or U12752 (N_12752,N_11452,N_11515);
and U12753 (N_12753,N_11578,N_11270);
or U12754 (N_12754,N_11839,N_11129);
nor U12755 (N_12755,N_11612,N_11189);
nor U12756 (N_12756,N_11121,N_11518);
xor U12757 (N_12757,N_11148,N_11927);
nor U12758 (N_12758,N_11971,N_11148);
xor U12759 (N_12759,N_11563,N_11049);
and U12760 (N_12760,N_11263,N_11245);
or U12761 (N_12761,N_11225,N_11520);
xnor U12762 (N_12762,N_11150,N_11579);
and U12763 (N_12763,N_11693,N_11670);
or U12764 (N_12764,N_11406,N_11966);
and U12765 (N_12765,N_11894,N_11328);
xor U12766 (N_12766,N_11210,N_11284);
and U12767 (N_12767,N_11246,N_11036);
xnor U12768 (N_12768,N_11399,N_11649);
xor U12769 (N_12769,N_11814,N_11322);
or U12770 (N_12770,N_11702,N_11979);
nand U12771 (N_12771,N_11293,N_11082);
xnor U12772 (N_12772,N_11067,N_11205);
and U12773 (N_12773,N_11930,N_11437);
nor U12774 (N_12774,N_11632,N_11787);
nand U12775 (N_12775,N_11855,N_11346);
and U12776 (N_12776,N_11627,N_11796);
or U12777 (N_12777,N_11628,N_11545);
nor U12778 (N_12778,N_11757,N_11785);
nor U12779 (N_12779,N_11466,N_11928);
nor U12780 (N_12780,N_11426,N_11145);
nor U12781 (N_12781,N_11646,N_11167);
or U12782 (N_12782,N_11840,N_11036);
or U12783 (N_12783,N_11434,N_11734);
nand U12784 (N_12784,N_11760,N_11346);
nor U12785 (N_12785,N_11805,N_11287);
xor U12786 (N_12786,N_11544,N_11075);
nand U12787 (N_12787,N_11505,N_11402);
xor U12788 (N_12788,N_11045,N_11144);
and U12789 (N_12789,N_11947,N_11423);
xor U12790 (N_12790,N_11832,N_11490);
xor U12791 (N_12791,N_11607,N_11664);
or U12792 (N_12792,N_11492,N_11649);
xor U12793 (N_12793,N_11829,N_11367);
nor U12794 (N_12794,N_11158,N_11168);
xnor U12795 (N_12795,N_11068,N_11800);
and U12796 (N_12796,N_11212,N_11203);
and U12797 (N_12797,N_11082,N_11920);
or U12798 (N_12798,N_11346,N_11728);
nand U12799 (N_12799,N_11662,N_11333);
and U12800 (N_12800,N_11823,N_11362);
nand U12801 (N_12801,N_11434,N_11228);
and U12802 (N_12802,N_11640,N_11236);
and U12803 (N_12803,N_11643,N_11317);
and U12804 (N_12804,N_11387,N_11519);
and U12805 (N_12805,N_11379,N_11957);
xnor U12806 (N_12806,N_11005,N_11524);
or U12807 (N_12807,N_11231,N_11757);
and U12808 (N_12808,N_11917,N_11156);
nand U12809 (N_12809,N_11939,N_11892);
or U12810 (N_12810,N_11280,N_11741);
xnor U12811 (N_12811,N_11635,N_11582);
xnor U12812 (N_12812,N_11430,N_11211);
or U12813 (N_12813,N_11727,N_11510);
nand U12814 (N_12814,N_11781,N_11798);
or U12815 (N_12815,N_11873,N_11320);
and U12816 (N_12816,N_11643,N_11038);
nor U12817 (N_12817,N_11039,N_11613);
and U12818 (N_12818,N_11220,N_11025);
nand U12819 (N_12819,N_11658,N_11300);
nor U12820 (N_12820,N_11802,N_11958);
xnor U12821 (N_12821,N_11970,N_11335);
or U12822 (N_12822,N_11614,N_11267);
and U12823 (N_12823,N_11189,N_11804);
nor U12824 (N_12824,N_11593,N_11843);
and U12825 (N_12825,N_11271,N_11660);
xnor U12826 (N_12826,N_11996,N_11425);
or U12827 (N_12827,N_11551,N_11177);
nor U12828 (N_12828,N_11375,N_11223);
nor U12829 (N_12829,N_11902,N_11426);
nor U12830 (N_12830,N_11144,N_11022);
xnor U12831 (N_12831,N_11135,N_11412);
nand U12832 (N_12832,N_11460,N_11626);
xnor U12833 (N_12833,N_11890,N_11405);
xnor U12834 (N_12834,N_11635,N_11508);
nor U12835 (N_12835,N_11117,N_11301);
or U12836 (N_12836,N_11435,N_11012);
or U12837 (N_12837,N_11217,N_11429);
nor U12838 (N_12838,N_11389,N_11538);
or U12839 (N_12839,N_11848,N_11336);
nor U12840 (N_12840,N_11323,N_11649);
nor U12841 (N_12841,N_11403,N_11011);
and U12842 (N_12842,N_11075,N_11778);
or U12843 (N_12843,N_11192,N_11503);
nor U12844 (N_12844,N_11679,N_11868);
nor U12845 (N_12845,N_11475,N_11417);
nor U12846 (N_12846,N_11907,N_11787);
nor U12847 (N_12847,N_11091,N_11228);
xnor U12848 (N_12848,N_11943,N_11557);
xor U12849 (N_12849,N_11070,N_11208);
nor U12850 (N_12850,N_11277,N_11722);
and U12851 (N_12851,N_11224,N_11171);
nor U12852 (N_12852,N_11356,N_11155);
and U12853 (N_12853,N_11601,N_11671);
xor U12854 (N_12854,N_11629,N_11572);
and U12855 (N_12855,N_11555,N_11687);
nand U12856 (N_12856,N_11999,N_11632);
nand U12857 (N_12857,N_11593,N_11618);
or U12858 (N_12858,N_11616,N_11727);
or U12859 (N_12859,N_11241,N_11473);
or U12860 (N_12860,N_11784,N_11859);
nor U12861 (N_12861,N_11271,N_11458);
nand U12862 (N_12862,N_11271,N_11160);
xor U12863 (N_12863,N_11819,N_11837);
nand U12864 (N_12864,N_11246,N_11135);
nor U12865 (N_12865,N_11602,N_11271);
and U12866 (N_12866,N_11048,N_11208);
or U12867 (N_12867,N_11969,N_11574);
or U12868 (N_12868,N_11614,N_11589);
or U12869 (N_12869,N_11884,N_11902);
nand U12870 (N_12870,N_11483,N_11037);
xnor U12871 (N_12871,N_11243,N_11621);
and U12872 (N_12872,N_11662,N_11231);
or U12873 (N_12873,N_11469,N_11626);
and U12874 (N_12874,N_11125,N_11012);
nand U12875 (N_12875,N_11840,N_11316);
xnor U12876 (N_12876,N_11012,N_11633);
nor U12877 (N_12877,N_11580,N_11292);
xor U12878 (N_12878,N_11004,N_11088);
nor U12879 (N_12879,N_11631,N_11341);
or U12880 (N_12880,N_11527,N_11883);
nor U12881 (N_12881,N_11536,N_11259);
and U12882 (N_12882,N_11232,N_11377);
xnor U12883 (N_12883,N_11910,N_11738);
xnor U12884 (N_12884,N_11394,N_11499);
xor U12885 (N_12885,N_11414,N_11564);
or U12886 (N_12886,N_11483,N_11811);
or U12887 (N_12887,N_11823,N_11669);
and U12888 (N_12888,N_11653,N_11972);
nor U12889 (N_12889,N_11210,N_11524);
or U12890 (N_12890,N_11683,N_11769);
or U12891 (N_12891,N_11358,N_11728);
nor U12892 (N_12892,N_11352,N_11442);
nand U12893 (N_12893,N_11862,N_11468);
nand U12894 (N_12894,N_11813,N_11223);
nand U12895 (N_12895,N_11323,N_11524);
and U12896 (N_12896,N_11899,N_11557);
xor U12897 (N_12897,N_11573,N_11661);
xnor U12898 (N_12898,N_11568,N_11529);
xnor U12899 (N_12899,N_11513,N_11231);
xor U12900 (N_12900,N_11552,N_11836);
nor U12901 (N_12901,N_11023,N_11972);
and U12902 (N_12902,N_11871,N_11672);
or U12903 (N_12903,N_11901,N_11706);
or U12904 (N_12904,N_11059,N_11958);
xor U12905 (N_12905,N_11432,N_11197);
xnor U12906 (N_12906,N_11175,N_11568);
xor U12907 (N_12907,N_11203,N_11256);
or U12908 (N_12908,N_11019,N_11156);
nand U12909 (N_12909,N_11433,N_11997);
nand U12910 (N_12910,N_11502,N_11545);
nand U12911 (N_12911,N_11140,N_11086);
nor U12912 (N_12912,N_11349,N_11902);
nand U12913 (N_12913,N_11988,N_11047);
nor U12914 (N_12914,N_11724,N_11854);
and U12915 (N_12915,N_11765,N_11906);
or U12916 (N_12916,N_11933,N_11651);
and U12917 (N_12917,N_11555,N_11812);
and U12918 (N_12918,N_11564,N_11861);
xor U12919 (N_12919,N_11649,N_11089);
xnor U12920 (N_12920,N_11894,N_11176);
xnor U12921 (N_12921,N_11694,N_11902);
nand U12922 (N_12922,N_11702,N_11770);
xor U12923 (N_12923,N_11909,N_11143);
xor U12924 (N_12924,N_11321,N_11376);
nand U12925 (N_12925,N_11958,N_11191);
xnor U12926 (N_12926,N_11196,N_11485);
nor U12927 (N_12927,N_11190,N_11156);
or U12928 (N_12928,N_11021,N_11323);
nand U12929 (N_12929,N_11959,N_11079);
or U12930 (N_12930,N_11749,N_11495);
or U12931 (N_12931,N_11062,N_11599);
xor U12932 (N_12932,N_11026,N_11790);
nand U12933 (N_12933,N_11195,N_11464);
nor U12934 (N_12934,N_11319,N_11873);
and U12935 (N_12935,N_11533,N_11946);
or U12936 (N_12936,N_11608,N_11596);
nand U12937 (N_12937,N_11083,N_11206);
or U12938 (N_12938,N_11098,N_11043);
xnor U12939 (N_12939,N_11148,N_11641);
and U12940 (N_12940,N_11099,N_11628);
nor U12941 (N_12941,N_11985,N_11276);
nand U12942 (N_12942,N_11469,N_11877);
or U12943 (N_12943,N_11602,N_11694);
nor U12944 (N_12944,N_11416,N_11838);
or U12945 (N_12945,N_11232,N_11383);
xnor U12946 (N_12946,N_11311,N_11344);
nor U12947 (N_12947,N_11941,N_11178);
nand U12948 (N_12948,N_11285,N_11825);
or U12949 (N_12949,N_11593,N_11053);
or U12950 (N_12950,N_11641,N_11012);
xnor U12951 (N_12951,N_11436,N_11819);
nand U12952 (N_12952,N_11150,N_11123);
nor U12953 (N_12953,N_11827,N_11937);
nand U12954 (N_12954,N_11380,N_11855);
or U12955 (N_12955,N_11639,N_11739);
and U12956 (N_12956,N_11683,N_11267);
nand U12957 (N_12957,N_11222,N_11777);
nor U12958 (N_12958,N_11652,N_11851);
and U12959 (N_12959,N_11438,N_11347);
nand U12960 (N_12960,N_11914,N_11304);
or U12961 (N_12961,N_11987,N_11382);
xor U12962 (N_12962,N_11664,N_11232);
nand U12963 (N_12963,N_11213,N_11153);
nor U12964 (N_12964,N_11349,N_11595);
xnor U12965 (N_12965,N_11700,N_11849);
or U12966 (N_12966,N_11044,N_11601);
nor U12967 (N_12967,N_11292,N_11239);
and U12968 (N_12968,N_11345,N_11272);
or U12969 (N_12969,N_11555,N_11746);
and U12970 (N_12970,N_11471,N_11571);
or U12971 (N_12971,N_11452,N_11711);
nor U12972 (N_12972,N_11153,N_11395);
xor U12973 (N_12973,N_11718,N_11058);
nand U12974 (N_12974,N_11755,N_11999);
nand U12975 (N_12975,N_11168,N_11563);
xnor U12976 (N_12976,N_11083,N_11524);
and U12977 (N_12977,N_11190,N_11977);
nor U12978 (N_12978,N_11615,N_11854);
nand U12979 (N_12979,N_11406,N_11112);
or U12980 (N_12980,N_11192,N_11560);
nor U12981 (N_12981,N_11579,N_11950);
or U12982 (N_12982,N_11178,N_11512);
nand U12983 (N_12983,N_11745,N_11912);
and U12984 (N_12984,N_11302,N_11268);
or U12985 (N_12985,N_11110,N_11069);
nand U12986 (N_12986,N_11558,N_11623);
nand U12987 (N_12987,N_11037,N_11961);
xnor U12988 (N_12988,N_11005,N_11989);
xor U12989 (N_12989,N_11211,N_11235);
xnor U12990 (N_12990,N_11849,N_11828);
or U12991 (N_12991,N_11042,N_11879);
xor U12992 (N_12992,N_11798,N_11707);
and U12993 (N_12993,N_11853,N_11989);
or U12994 (N_12994,N_11745,N_11488);
nand U12995 (N_12995,N_11508,N_11373);
nor U12996 (N_12996,N_11210,N_11422);
nand U12997 (N_12997,N_11105,N_11945);
or U12998 (N_12998,N_11763,N_11499);
or U12999 (N_12999,N_11540,N_11481);
xor U13000 (N_13000,N_12307,N_12875);
or U13001 (N_13001,N_12415,N_12991);
xnor U13002 (N_13002,N_12715,N_12840);
and U13003 (N_13003,N_12977,N_12032);
nor U13004 (N_13004,N_12393,N_12976);
nor U13005 (N_13005,N_12544,N_12876);
and U13006 (N_13006,N_12185,N_12873);
nand U13007 (N_13007,N_12239,N_12075);
xnor U13008 (N_13008,N_12492,N_12826);
and U13009 (N_13009,N_12647,N_12731);
nand U13010 (N_13010,N_12115,N_12552);
nor U13011 (N_13011,N_12081,N_12825);
nor U13012 (N_13012,N_12313,N_12680);
nand U13013 (N_13013,N_12286,N_12665);
nor U13014 (N_13014,N_12662,N_12880);
or U13015 (N_13015,N_12163,N_12030);
nand U13016 (N_13016,N_12007,N_12975);
and U13017 (N_13017,N_12669,N_12835);
or U13018 (N_13018,N_12343,N_12518);
nand U13019 (N_13019,N_12019,N_12342);
and U13020 (N_13020,N_12214,N_12015);
nor U13021 (N_13021,N_12484,N_12747);
nand U13022 (N_13022,N_12579,N_12199);
nand U13023 (N_13023,N_12437,N_12939);
xor U13024 (N_13024,N_12570,N_12741);
xor U13025 (N_13025,N_12907,N_12009);
nand U13026 (N_13026,N_12959,N_12703);
nor U13027 (N_13027,N_12521,N_12165);
xor U13028 (N_13028,N_12141,N_12671);
nand U13029 (N_13029,N_12349,N_12330);
xor U13030 (N_13030,N_12033,N_12436);
nor U13031 (N_13031,N_12765,N_12157);
or U13032 (N_13032,N_12283,N_12445);
and U13033 (N_13033,N_12182,N_12555);
and U13034 (N_13034,N_12174,N_12225);
nand U13035 (N_13035,N_12798,N_12045);
or U13036 (N_13036,N_12859,N_12730);
and U13037 (N_13037,N_12996,N_12622);
and U13038 (N_13038,N_12125,N_12297);
or U13039 (N_13039,N_12142,N_12711);
nor U13040 (N_13040,N_12516,N_12997);
xor U13041 (N_13041,N_12598,N_12234);
nor U13042 (N_13042,N_12596,N_12001);
and U13043 (N_13043,N_12129,N_12515);
or U13044 (N_13044,N_12729,N_12233);
nor U13045 (N_13045,N_12384,N_12450);
and U13046 (N_13046,N_12970,N_12732);
and U13047 (N_13047,N_12814,N_12014);
or U13048 (N_13048,N_12633,N_12588);
or U13049 (N_13049,N_12966,N_12005);
or U13050 (N_13050,N_12774,N_12533);
nor U13051 (N_13051,N_12634,N_12938);
or U13052 (N_13052,N_12919,N_12433);
and U13053 (N_13053,N_12781,N_12797);
and U13054 (N_13054,N_12098,N_12004);
or U13055 (N_13055,N_12520,N_12368);
or U13056 (N_13056,N_12205,N_12618);
or U13057 (N_13057,N_12587,N_12183);
nand U13058 (N_13058,N_12557,N_12025);
xor U13059 (N_13059,N_12345,N_12837);
and U13060 (N_13060,N_12000,N_12497);
and U13061 (N_13061,N_12309,N_12606);
xor U13062 (N_13062,N_12910,N_12960);
nor U13063 (N_13063,N_12105,N_12325);
and U13064 (N_13064,N_12188,N_12720);
nor U13065 (N_13065,N_12827,N_12409);
and U13066 (N_13066,N_12989,N_12100);
nor U13067 (N_13067,N_12251,N_12695);
nor U13068 (N_13068,N_12628,N_12169);
or U13069 (N_13069,N_12062,N_12351);
nand U13070 (N_13070,N_12379,N_12044);
or U13071 (N_13071,N_12945,N_12698);
and U13072 (N_13072,N_12057,N_12974);
nand U13073 (N_13073,N_12672,N_12010);
and U13074 (N_13074,N_12921,N_12635);
or U13075 (N_13075,N_12365,N_12885);
and U13076 (N_13076,N_12314,N_12083);
nand U13077 (N_13077,N_12427,N_12046);
or U13078 (N_13078,N_12882,N_12853);
and U13079 (N_13079,N_12326,N_12612);
nor U13080 (N_13080,N_12712,N_12324);
nand U13081 (N_13081,N_12152,N_12318);
nor U13082 (N_13082,N_12446,N_12863);
and U13083 (N_13083,N_12375,N_12689);
nand U13084 (N_13084,N_12973,N_12095);
or U13085 (N_13085,N_12155,N_12517);
or U13086 (N_13086,N_12394,N_12551);
xor U13087 (N_13087,N_12844,N_12793);
xnor U13088 (N_13088,N_12834,N_12531);
xor U13089 (N_13089,N_12210,N_12249);
xor U13090 (N_13090,N_12762,N_12442);
and U13091 (N_13091,N_12874,N_12128);
xor U13092 (N_13092,N_12936,N_12759);
or U13093 (N_13093,N_12138,N_12684);
or U13094 (N_13094,N_12193,N_12293);
and U13095 (N_13095,N_12078,N_12702);
or U13096 (N_13096,N_12564,N_12704);
or U13097 (N_13097,N_12200,N_12982);
nor U13098 (N_13098,N_12820,N_12813);
xnor U13099 (N_13099,N_12300,N_12829);
xnor U13100 (N_13100,N_12179,N_12553);
nor U13101 (N_13101,N_12593,N_12559);
and U13102 (N_13102,N_12211,N_12920);
or U13103 (N_13103,N_12080,N_12094);
and U13104 (N_13104,N_12012,N_12257);
and U13105 (N_13105,N_12725,N_12585);
and U13106 (N_13106,N_12319,N_12385);
nand U13107 (N_13107,N_12038,N_12654);
or U13108 (N_13108,N_12726,N_12845);
xor U13109 (N_13109,N_12637,N_12605);
nor U13110 (N_13110,N_12479,N_12070);
xor U13111 (N_13111,N_12942,N_12150);
and U13112 (N_13112,N_12928,N_12487);
nor U13113 (N_13113,N_12458,N_12180);
or U13114 (N_13114,N_12438,N_12122);
or U13115 (N_13115,N_12485,N_12916);
or U13116 (N_13116,N_12740,N_12819);
nor U13117 (N_13117,N_12263,N_12491);
or U13118 (N_13118,N_12562,N_12790);
nor U13119 (N_13119,N_12443,N_12830);
and U13120 (N_13120,N_12203,N_12498);
nor U13121 (N_13121,N_12232,N_12096);
nand U13122 (N_13122,N_12746,N_12131);
nor U13123 (N_13123,N_12255,N_12031);
xor U13124 (N_13124,N_12400,N_12049);
xnor U13125 (N_13125,N_12466,N_12507);
xor U13126 (N_13126,N_12744,N_12683);
xnor U13127 (N_13127,N_12465,N_12911);
nand U13128 (N_13128,N_12550,N_12963);
or U13129 (N_13129,N_12716,N_12506);
nor U13130 (N_13130,N_12259,N_12900);
nand U13131 (N_13131,N_12463,N_12527);
nor U13132 (N_13132,N_12363,N_12888);
xnor U13133 (N_13133,N_12476,N_12164);
xnor U13134 (N_13134,N_12119,N_12364);
nand U13135 (N_13135,N_12084,N_12528);
nor U13136 (N_13136,N_12294,N_12432);
nand U13137 (N_13137,N_12993,N_12114);
nor U13138 (N_13138,N_12322,N_12962);
nand U13139 (N_13139,N_12904,N_12076);
or U13140 (N_13140,N_12664,N_12617);
or U13141 (N_13141,N_12955,N_12186);
or U13142 (N_13142,N_12435,N_12289);
nand U13143 (N_13143,N_12235,N_12786);
and U13144 (N_13144,N_12295,N_12422);
or U13145 (N_13145,N_12299,N_12511);
nand U13146 (N_13146,N_12111,N_12583);
or U13147 (N_13147,N_12120,N_12303);
xor U13148 (N_13148,N_12079,N_12493);
xnor U13149 (N_13149,N_12134,N_12275);
nand U13150 (N_13150,N_12717,N_12878);
and U13151 (N_13151,N_12469,N_12398);
or U13152 (N_13152,N_12525,N_12956);
and U13153 (N_13153,N_12983,N_12924);
xor U13154 (N_13154,N_12495,N_12316);
or U13155 (N_13155,N_12705,N_12477);
xnor U13156 (N_13156,N_12808,N_12721);
nor U13157 (N_13157,N_12344,N_12361);
xnor U13158 (N_13158,N_12104,N_12272);
nand U13159 (N_13159,N_12615,N_12737);
nand U13160 (N_13160,N_12306,N_12254);
and U13161 (N_13161,N_12906,N_12568);
or U13162 (N_13162,N_12108,N_12222);
and U13163 (N_13163,N_12018,N_12026);
and U13164 (N_13164,N_12500,N_12091);
nand U13165 (N_13165,N_12644,N_12584);
nor U13166 (N_13166,N_12686,N_12847);
or U13167 (N_13167,N_12857,N_12201);
and U13168 (N_13168,N_12632,N_12504);
nand U13169 (N_13169,N_12748,N_12688);
nor U13170 (N_13170,N_12219,N_12929);
xnor U13171 (N_13171,N_12773,N_12950);
and U13172 (N_13172,N_12374,N_12941);
and U13173 (N_13173,N_12085,N_12292);
or U13174 (N_13174,N_12238,N_12865);
nor U13175 (N_13175,N_12953,N_12943);
nand U13176 (N_13176,N_12630,N_12089);
xnor U13177 (N_13177,N_12667,N_12133);
or U13178 (N_13178,N_12170,N_12503);
nor U13179 (N_13179,N_12707,N_12571);
and U13180 (N_13180,N_12724,N_12679);
or U13181 (N_13181,N_12839,N_12020);
nor U13182 (N_13182,N_12532,N_12961);
and U13183 (N_13183,N_12397,N_12244);
xor U13184 (N_13184,N_12146,N_12126);
and U13185 (N_13185,N_12693,N_12899);
and U13186 (N_13186,N_12039,N_12358);
and U13187 (N_13187,N_12240,N_12946);
or U13188 (N_13188,N_12713,N_12988);
and U13189 (N_13189,N_12107,N_12243);
or U13190 (N_13190,N_12071,N_12855);
nand U13191 (N_13191,N_12428,N_12171);
nand U13192 (N_13192,N_12408,N_12591);
nand U13193 (N_13193,N_12843,N_12008);
or U13194 (N_13194,N_12540,N_12957);
or U13195 (N_13195,N_12246,N_12569);
nor U13196 (N_13196,N_12348,N_12984);
nand U13197 (N_13197,N_12058,N_12524);
nand U13198 (N_13198,N_12474,N_12425);
and U13199 (N_13199,N_12581,N_12601);
and U13200 (N_13200,N_12917,N_12756);
or U13201 (N_13201,N_12577,N_12710);
xnor U13202 (N_13202,N_12590,N_12831);
and U13203 (N_13203,N_12812,N_12068);
nand U13204 (N_13204,N_12992,N_12833);
and U13205 (N_13205,N_12894,N_12459);
or U13206 (N_13206,N_12224,N_12241);
and U13207 (N_13207,N_12852,N_12505);
nand U13208 (N_13208,N_12836,N_12195);
or U13209 (N_13209,N_12206,N_12770);
nor U13210 (N_13210,N_12734,N_12915);
nand U13211 (N_13211,N_12284,N_12728);
nor U13212 (N_13212,N_12228,N_12692);
or U13213 (N_13213,N_12047,N_12794);
nor U13214 (N_13214,N_12807,N_12869);
or U13215 (N_13215,N_12461,N_12420);
nand U13216 (N_13216,N_12455,N_12287);
or U13217 (N_13217,N_12952,N_12029);
nor U13218 (N_13218,N_12610,N_12714);
xnor U13219 (N_13219,N_12822,N_12566);
nand U13220 (N_13220,N_12181,N_12296);
and U13221 (N_13221,N_12271,N_12901);
and U13222 (N_13222,N_12273,N_12048);
and U13223 (N_13223,N_12609,N_12755);
xor U13224 (N_13224,N_12594,N_12607);
or U13225 (N_13225,N_12117,N_12803);
and U13226 (N_13226,N_12750,N_12061);
and U13227 (N_13227,N_12968,N_12260);
or U13228 (N_13228,N_12818,N_12456);
nand U13229 (N_13229,N_12301,N_12481);
or U13230 (N_13230,N_12460,N_12124);
nor U13231 (N_13231,N_12360,N_12371);
nor U13232 (N_13232,N_12870,N_12202);
xnor U13233 (N_13233,N_12556,N_12245);
xor U13234 (N_13234,N_12578,N_12694);
nand U13235 (N_13235,N_12060,N_12754);
or U13236 (N_13236,N_12871,N_12093);
and U13237 (N_13237,N_12337,N_12670);
or U13238 (N_13238,N_12369,N_12423);
nor U13239 (N_13239,N_12090,N_12426);
and U13240 (N_13240,N_12391,N_12884);
xor U13241 (N_13241,N_12370,N_12625);
nor U13242 (N_13242,N_12329,N_12561);
or U13243 (N_13243,N_12650,N_12646);
nor U13244 (N_13244,N_12529,N_12539);
and U13245 (N_13245,N_12783,N_12616);
xor U13246 (N_13246,N_12903,N_12810);
nand U13247 (N_13247,N_12340,N_12543);
or U13248 (N_13248,N_12066,N_12482);
nand U13249 (N_13249,N_12380,N_12655);
nand U13250 (N_13250,N_12889,N_12087);
and U13251 (N_13251,N_12995,N_12331);
nand U13252 (N_13252,N_12473,N_12334);
nor U13253 (N_13253,N_12190,N_12537);
and U13254 (N_13254,N_12549,N_12042);
nor U13255 (N_13255,N_12097,N_12651);
nand U13256 (N_13256,N_12278,N_12805);
xor U13257 (N_13257,N_12802,N_12327);
and U13258 (N_13258,N_12013,N_12502);
or U13259 (N_13259,N_12867,N_12738);
xnor U13260 (N_13260,N_12896,N_12264);
xor U13261 (N_13261,N_12512,N_12378);
nand U13262 (N_13262,N_12269,N_12868);
or U13263 (N_13263,N_12411,N_12778);
nor U13264 (N_13264,N_12769,N_12310);
xnor U13265 (N_13265,N_12513,N_12382);
or U13266 (N_13266,N_12733,N_12501);
nor U13267 (N_13267,N_12883,N_12449);
nand U13268 (N_13268,N_12902,N_12535);
nand U13269 (N_13269,N_12700,N_12653);
nor U13270 (N_13270,N_12419,N_12806);
or U13271 (N_13271,N_12627,N_12392);
and U13272 (N_13272,N_12106,N_12077);
and U13273 (N_13273,N_12898,N_12389);
xnor U13274 (N_13274,N_12777,N_12580);
and U13275 (N_13275,N_12151,N_12574);
xnor U13276 (N_13276,N_12209,N_12040);
nand U13277 (N_13277,N_12499,N_12050);
nand U13278 (N_13278,N_12242,N_12053);
xor U13279 (N_13279,N_12949,N_12230);
nor U13280 (N_13280,N_12668,N_12223);
and U13281 (N_13281,N_12288,N_12268);
and U13282 (N_13282,N_12522,N_12795);
and U13283 (N_13283,N_12123,N_12508);
xnor U13284 (N_13284,N_12624,N_12841);
nand U13285 (N_13285,N_12320,N_12130);
nand U13286 (N_13286,N_12987,N_12418);
xor U13287 (N_13287,N_12752,N_12266);
nand U13288 (N_13288,N_12173,N_12161);
and U13289 (N_13289,N_12611,N_12328);
nor U13290 (N_13290,N_12823,N_12103);
and U13291 (N_13291,N_12041,N_12879);
nor U13292 (N_13292,N_12036,N_12373);
nor U13293 (N_13293,N_12697,N_12406);
nand U13294 (N_13294,N_12069,N_12972);
nor U13295 (N_13295,N_12052,N_12118);
nor U13296 (N_13296,N_12872,N_12563);
or U13297 (N_13297,N_12399,N_12897);
nor U13298 (N_13298,N_12064,N_12467);
and U13299 (N_13299,N_12431,N_12761);
nand U13300 (N_13300,N_12191,N_12980);
and U13301 (N_13301,N_12541,N_12626);
nand U13302 (N_13302,N_12401,N_12887);
nor U13303 (N_13303,N_12699,N_12811);
nor U13304 (N_13304,N_12099,N_12035);
xor U13305 (N_13305,N_12496,N_12675);
and U13306 (N_13306,N_12908,N_12799);
nor U13307 (N_13307,N_12022,N_12247);
nand U13308 (N_13308,N_12312,N_12416);
and U13309 (N_13309,N_12560,N_12851);
or U13310 (N_13310,N_12971,N_12250);
xnor U13311 (N_13311,N_12922,N_12353);
nand U13312 (N_13312,N_12817,N_12102);
xor U13313 (N_13313,N_12367,N_12362);
nand U13314 (N_13314,N_12931,N_12457);
and U13315 (N_13315,N_12404,N_12196);
nor U13316 (N_13316,N_12753,N_12749);
nor U13317 (N_13317,N_12402,N_12153);
nor U13318 (N_13318,N_12519,N_12267);
and U13319 (N_13319,N_12780,N_12121);
or U13320 (N_13320,N_12739,N_12454);
xnor U13321 (N_13321,N_12016,N_12766);
and U13322 (N_13322,N_12494,N_12676);
or U13323 (N_13323,N_12860,N_12413);
or U13324 (N_13324,N_12387,N_12291);
nor U13325 (N_13325,N_12430,N_12735);
or U13326 (N_13326,N_12964,N_12718);
xor U13327 (N_13327,N_12421,N_12227);
nor U13328 (N_13328,N_12854,N_12926);
nor U13329 (N_13329,N_12088,N_12175);
nand U13330 (N_13330,N_12072,N_12218);
and U13331 (N_13331,N_12768,N_12376);
or U13332 (N_13332,N_12639,N_12573);
or U13333 (N_13333,N_12403,N_12471);
xnor U13334 (N_13334,N_12478,N_12663);
xnor U13335 (N_13335,N_12101,N_12192);
xor U13336 (N_13336,N_12687,N_12923);
nor U13337 (N_13337,N_12414,N_12523);
xnor U13338 (N_13338,N_12767,N_12785);
nand U13339 (N_13339,N_12816,N_12149);
nand U13340 (N_13340,N_12156,N_12339);
nor U13341 (N_13341,N_12649,N_12110);
nand U13342 (N_13342,N_12642,N_12113);
xnor U13343 (N_13343,N_12308,N_12148);
nor U13344 (N_13344,N_12440,N_12434);
or U13345 (N_13345,N_12775,N_12947);
or U13346 (N_13346,N_12074,N_12258);
or U13347 (N_13347,N_12990,N_12784);
nor U13348 (N_13348,N_12147,N_12490);
nand U13349 (N_13349,N_12510,N_12056);
or U13350 (N_13350,N_12043,N_12509);
or U13351 (N_13351,N_12444,N_12412);
xor U13352 (N_13352,N_12881,N_12981);
or U13353 (N_13353,N_12986,N_12661);
nor U13354 (N_13354,N_12178,N_12850);
nand U13355 (N_13355,N_12545,N_12127);
xor U13356 (N_13356,N_12621,N_12927);
or U13357 (N_13357,N_12930,N_12276);
and U13358 (N_13358,N_12160,N_12554);
and U13359 (N_13359,N_12613,N_12252);
xor U13360 (N_13360,N_12140,N_12690);
and U13361 (N_13361,N_12745,N_12999);
and U13362 (N_13362,N_12858,N_12547);
nand U13363 (N_13363,N_12405,N_12172);
nor U13364 (N_13364,N_12821,N_12951);
and U13365 (N_13365,N_12336,N_12281);
nand U13366 (N_13366,N_12388,N_12144);
nand U13367 (N_13367,N_12608,N_12226);
nor U13368 (N_13368,N_12448,N_12760);
nand U13369 (N_13369,N_12166,N_12204);
nand U13370 (N_13370,N_12998,N_12346);
xor U13371 (N_13371,N_12832,N_12772);
nand U13372 (N_13372,N_12789,N_12913);
or U13373 (N_13373,N_12582,N_12395);
nor U13374 (N_13374,N_12877,N_12751);
nand U13375 (N_13375,N_12441,N_12323);
and U13376 (N_13376,N_12197,N_12279);
nand U13377 (N_13377,N_12198,N_12447);
or U13378 (N_13378,N_12116,N_12154);
nand U13379 (N_13379,N_12390,N_12864);
nor U13380 (N_13380,N_12536,N_12595);
nor U13381 (N_13381,N_12534,N_12236);
or U13382 (N_13382,N_12439,N_12347);
or U13383 (N_13383,N_12640,N_12315);
xor U13384 (N_13384,N_12357,N_12727);
nor U13385 (N_13385,N_12377,N_12213);
and U13386 (N_13386,N_12429,N_12265);
and U13387 (N_13387,N_12787,N_12892);
xnor U13388 (N_13388,N_12742,N_12194);
or U13389 (N_13389,N_12037,N_12848);
nor U13390 (N_13390,N_12159,N_12514);
xnor U13391 (N_13391,N_12472,N_12335);
or U13392 (N_13392,N_12054,N_12600);
nor U13393 (N_13393,N_12862,N_12905);
xor U13394 (N_13394,N_12652,N_12464);
xnor U13395 (N_13395,N_12978,N_12912);
and U13396 (N_13396,N_12453,N_12158);
nand U13397 (N_13397,N_12207,N_12217);
xor U13398 (N_13398,N_12967,N_12352);
or U13399 (N_13399,N_12480,N_12002);
or U13400 (N_13400,N_12332,N_12708);
nand U13401 (N_13401,N_12417,N_12658);
and U13402 (N_13402,N_12576,N_12475);
xnor U13403 (N_13403,N_12709,N_12965);
or U13404 (N_13404,N_12589,N_12891);
and U13405 (N_13405,N_12462,N_12918);
nand U13406 (N_13406,N_12027,N_12304);
nor U13407 (N_13407,N_12407,N_12599);
nor U13408 (N_13408,N_12979,N_12623);
or U13409 (N_13409,N_12355,N_12909);
nand U13410 (N_13410,N_12643,N_12828);
and U13411 (N_13411,N_12678,N_12262);
or U13412 (N_13412,N_12604,N_12782);
nand U13413 (N_13413,N_12933,N_12489);
nor U13414 (N_13414,N_12452,N_12063);
and U13415 (N_13415,N_12011,N_12256);
nand U13416 (N_13416,N_12137,N_12006);
or U13417 (N_13417,N_12849,N_12285);
nand U13418 (N_13418,N_12723,N_12925);
xor U13419 (N_13419,N_12359,N_12086);
nor U13420 (N_13420,N_12856,N_12958);
xor U13421 (N_13421,N_12526,N_12162);
nor U13422 (N_13422,N_12666,N_12758);
and U13423 (N_13423,N_12937,N_12145);
and U13424 (N_13424,N_12656,N_12788);
nor U13425 (N_13425,N_12082,N_12338);
nor U13426 (N_13426,N_12602,N_12890);
nand U13427 (N_13427,N_12696,N_12270);
or U13428 (N_13428,N_12994,N_12944);
or U13429 (N_13429,N_12763,N_12935);
xor U13430 (N_13430,N_12682,N_12736);
nor U13431 (N_13431,N_12893,N_12112);
nor U13432 (N_13432,N_12815,N_12620);
nand U13433 (N_13433,N_12572,N_12645);
and U13434 (N_13434,N_12631,N_12167);
or U13435 (N_13435,N_12221,N_12567);
nor U13436 (N_13436,N_12681,N_12298);
or U13437 (N_13437,N_12317,N_12065);
xnor U13438 (N_13438,N_12757,N_12792);
or U13439 (N_13439,N_12132,N_12135);
or U13440 (N_13440,N_12673,N_12073);
and U13441 (N_13441,N_12619,N_12538);
nand U13442 (N_13442,N_12638,N_12648);
or U13443 (N_13443,N_12143,N_12597);
xnor U13444 (N_13444,N_12800,N_12470);
and U13445 (N_13445,N_12809,N_12017);
or U13446 (N_13446,N_12229,N_12176);
nor U13447 (N_13447,N_12136,N_12109);
nand U13448 (N_13448,N_12261,N_12603);
or U13449 (N_13449,N_12350,N_12764);
nor U13450 (N_13450,N_12948,N_12024);
xor U13451 (N_13451,N_12356,N_12722);
xnor U13452 (N_13452,N_12548,N_12354);
nor U13453 (N_13453,N_12023,N_12824);
nor U13454 (N_13454,N_12059,N_12629);
xor U13455 (N_13455,N_12311,N_12372);
nand U13456 (N_13456,N_12804,N_12366);
nand U13457 (N_13457,N_12614,N_12248);
nor U13458 (N_13458,N_12954,N_12895);
and U13459 (N_13459,N_12846,N_12184);
and U13460 (N_13460,N_12530,N_12341);
nand U13461 (N_13461,N_12842,N_12021);
xnor U13462 (N_13462,N_12969,N_12215);
and U13463 (N_13463,N_12657,N_12779);
xor U13464 (N_13464,N_12274,N_12383);
and U13465 (N_13465,N_12220,N_12575);
nand U13466 (N_13466,N_12838,N_12187);
nor U13467 (N_13467,N_12985,N_12189);
xnor U13468 (N_13468,N_12674,N_12028);
xnor U13469 (N_13469,N_12719,N_12791);
nor U13470 (N_13470,N_12677,N_12168);
and U13471 (N_13471,N_12691,N_12641);
or U13472 (N_13472,N_12424,N_12051);
nand U13473 (N_13473,N_12483,N_12003);
and U13474 (N_13474,N_12290,N_12801);
xnor U13475 (N_13475,N_12282,N_12636);
and U13476 (N_13476,N_12321,N_12546);
and U13477 (N_13477,N_12934,N_12706);
nand U13478 (N_13478,N_12488,N_12861);
nand U13479 (N_13479,N_12468,N_12558);
or U13480 (N_13480,N_12092,N_12659);
and U13481 (N_13481,N_12302,N_12386);
xor U13482 (N_13482,N_12743,N_12486);
nand U13483 (N_13483,N_12776,N_12586);
or U13484 (N_13484,N_12208,N_12451);
or U13485 (N_13485,N_12067,N_12231);
xor U13486 (N_13486,N_12542,N_12940);
nor U13487 (N_13487,N_12055,N_12796);
nor U13488 (N_13488,N_12914,N_12034);
or U13489 (N_13489,N_12212,N_12280);
nor U13490 (N_13490,N_12277,N_12177);
and U13491 (N_13491,N_12396,N_12701);
or U13492 (N_13492,N_12410,N_12237);
and U13493 (N_13493,N_12381,N_12660);
xor U13494 (N_13494,N_12886,N_12305);
nor U13495 (N_13495,N_12216,N_12565);
nand U13496 (N_13496,N_12685,N_12932);
and U13497 (N_13497,N_12333,N_12253);
xnor U13498 (N_13498,N_12592,N_12139);
and U13499 (N_13499,N_12866,N_12771);
xor U13500 (N_13500,N_12420,N_12986);
xor U13501 (N_13501,N_12382,N_12022);
nor U13502 (N_13502,N_12909,N_12939);
nor U13503 (N_13503,N_12333,N_12459);
nand U13504 (N_13504,N_12195,N_12617);
nor U13505 (N_13505,N_12322,N_12259);
nor U13506 (N_13506,N_12280,N_12617);
or U13507 (N_13507,N_12151,N_12381);
xnor U13508 (N_13508,N_12840,N_12763);
nand U13509 (N_13509,N_12150,N_12054);
xor U13510 (N_13510,N_12815,N_12454);
nand U13511 (N_13511,N_12689,N_12468);
xnor U13512 (N_13512,N_12759,N_12025);
and U13513 (N_13513,N_12529,N_12724);
nand U13514 (N_13514,N_12173,N_12748);
and U13515 (N_13515,N_12697,N_12567);
and U13516 (N_13516,N_12392,N_12507);
nor U13517 (N_13517,N_12931,N_12999);
nor U13518 (N_13518,N_12499,N_12219);
nand U13519 (N_13519,N_12532,N_12373);
and U13520 (N_13520,N_12602,N_12407);
and U13521 (N_13521,N_12182,N_12193);
or U13522 (N_13522,N_12791,N_12431);
xor U13523 (N_13523,N_12232,N_12968);
nor U13524 (N_13524,N_12335,N_12762);
nand U13525 (N_13525,N_12388,N_12033);
xnor U13526 (N_13526,N_12355,N_12991);
nor U13527 (N_13527,N_12785,N_12163);
and U13528 (N_13528,N_12862,N_12464);
or U13529 (N_13529,N_12327,N_12191);
xnor U13530 (N_13530,N_12494,N_12475);
nand U13531 (N_13531,N_12909,N_12739);
xor U13532 (N_13532,N_12240,N_12884);
xnor U13533 (N_13533,N_12521,N_12924);
or U13534 (N_13534,N_12893,N_12269);
xor U13535 (N_13535,N_12483,N_12499);
nor U13536 (N_13536,N_12059,N_12055);
nor U13537 (N_13537,N_12596,N_12837);
or U13538 (N_13538,N_12105,N_12122);
nor U13539 (N_13539,N_12018,N_12072);
or U13540 (N_13540,N_12657,N_12302);
xnor U13541 (N_13541,N_12749,N_12488);
and U13542 (N_13542,N_12566,N_12660);
nor U13543 (N_13543,N_12607,N_12964);
nand U13544 (N_13544,N_12148,N_12724);
xor U13545 (N_13545,N_12045,N_12561);
nor U13546 (N_13546,N_12853,N_12767);
nand U13547 (N_13547,N_12709,N_12773);
nor U13548 (N_13548,N_12341,N_12280);
nand U13549 (N_13549,N_12565,N_12760);
and U13550 (N_13550,N_12319,N_12432);
nand U13551 (N_13551,N_12542,N_12728);
nand U13552 (N_13552,N_12730,N_12491);
xnor U13553 (N_13553,N_12615,N_12123);
nand U13554 (N_13554,N_12501,N_12743);
nor U13555 (N_13555,N_12008,N_12417);
or U13556 (N_13556,N_12256,N_12849);
or U13557 (N_13557,N_12848,N_12491);
xnor U13558 (N_13558,N_12767,N_12880);
nand U13559 (N_13559,N_12051,N_12244);
or U13560 (N_13560,N_12515,N_12127);
xnor U13561 (N_13561,N_12654,N_12495);
nand U13562 (N_13562,N_12999,N_12832);
xor U13563 (N_13563,N_12374,N_12275);
nor U13564 (N_13564,N_12573,N_12464);
nor U13565 (N_13565,N_12407,N_12784);
xnor U13566 (N_13566,N_12626,N_12668);
xnor U13567 (N_13567,N_12927,N_12730);
xnor U13568 (N_13568,N_12637,N_12889);
or U13569 (N_13569,N_12140,N_12872);
or U13570 (N_13570,N_12552,N_12974);
nor U13571 (N_13571,N_12534,N_12285);
and U13572 (N_13572,N_12396,N_12851);
nor U13573 (N_13573,N_12674,N_12092);
xnor U13574 (N_13574,N_12687,N_12612);
or U13575 (N_13575,N_12720,N_12880);
nand U13576 (N_13576,N_12676,N_12952);
nor U13577 (N_13577,N_12913,N_12897);
nand U13578 (N_13578,N_12159,N_12987);
nand U13579 (N_13579,N_12172,N_12115);
or U13580 (N_13580,N_12605,N_12792);
nor U13581 (N_13581,N_12510,N_12395);
nor U13582 (N_13582,N_12427,N_12560);
nor U13583 (N_13583,N_12770,N_12480);
or U13584 (N_13584,N_12609,N_12261);
and U13585 (N_13585,N_12915,N_12645);
nand U13586 (N_13586,N_12974,N_12644);
and U13587 (N_13587,N_12473,N_12202);
nor U13588 (N_13588,N_12610,N_12460);
and U13589 (N_13589,N_12955,N_12589);
and U13590 (N_13590,N_12407,N_12862);
nand U13591 (N_13591,N_12369,N_12611);
nor U13592 (N_13592,N_12663,N_12260);
or U13593 (N_13593,N_12642,N_12832);
nor U13594 (N_13594,N_12749,N_12823);
and U13595 (N_13595,N_12324,N_12580);
or U13596 (N_13596,N_12567,N_12914);
and U13597 (N_13597,N_12372,N_12084);
or U13598 (N_13598,N_12412,N_12153);
nand U13599 (N_13599,N_12415,N_12117);
and U13600 (N_13600,N_12599,N_12796);
and U13601 (N_13601,N_12938,N_12103);
or U13602 (N_13602,N_12909,N_12902);
xnor U13603 (N_13603,N_12042,N_12809);
xor U13604 (N_13604,N_12601,N_12063);
and U13605 (N_13605,N_12632,N_12645);
nor U13606 (N_13606,N_12499,N_12317);
nand U13607 (N_13607,N_12906,N_12513);
nor U13608 (N_13608,N_12992,N_12207);
nand U13609 (N_13609,N_12864,N_12816);
xnor U13610 (N_13610,N_12446,N_12171);
nand U13611 (N_13611,N_12573,N_12069);
nand U13612 (N_13612,N_12587,N_12730);
nand U13613 (N_13613,N_12615,N_12912);
nand U13614 (N_13614,N_12966,N_12086);
and U13615 (N_13615,N_12642,N_12299);
xnor U13616 (N_13616,N_12298,N_12987);
or U13617 (N_13617,N_12319,N_12181);
xor U13618 (N_13618,N_12100,N_12577);
xor U13619 (N_13619,N_12618,N_12617);
nand U13620 (N_13620,N_12507,N_12041);
and U13621 (N_13621,N_12142,N_12559);
nand U13622 (N_13622,N_12177,N_12789);
or U13623 (N_13623,N_12757,N_12564);
or U13624 (N_13624,N_12990,N_12268);
nand U13625 (N_13625,N_12358,N_12551);
xnor U13626 (N_13626,N_12678,N_12048);
nor U13627 (N_13627,N_12003,N_12541);
and U13628 (N_13628,N_12886,N_12268);
nor U13629 (N_13629,N_12418,N_12481);
nand U13630 (N_13630,N_12512,N_12028);
or U13631 (N_13631,N_12528,N_12013);
or U13632 (N_13632,N_12188,N_12289);
nand U13633 (N_13633,N_12877,N_12658);
nor U13634 (N_13634,N_12401,N_12741);
and U13635 (N_13635,N_12015,N_12859);
or U13636 (N_13636,N_12936,N_12177);
or U13637 (N_13637,N_12261,N_12359);
and U13638 (N_13638,N_12745,N_12568);
xnor U13639 (N_13639,N_12658,N_12810);
nand U13640 (N_13640,N_12409,N_12743);
nand U13641 (N_13641,N_12105,N_12039);
nor U13642 (N_13642,N_12971,N_12625);
or U13643 (N_13643,N_12428,N_12913);
nor U13644 (N_13644,N_12975,N_12870);
xor U13645 (N_13645,N_12026,N_12234);
or U13646 (N_13646,N_12962,N_12469);
xor U13647 (N_13647,N_12826,N_12178);
xor U13648 (N_13648,N_12626,N_12760);
and U13649 (N_13649,N_12921,N_12395);
or U13650 (N_13650,N_12428,N_12053);
xnor U13651 (N_13651,N_12732,N_12875);
nand U13652 (N_13652,N_12034,N_12312);
or U13653 (N_13653,N_12059,N_12950);
xnor U13654 (N_13654,N_12133,N_12122);
or U13655 (N_13655,N_12495,N_12396);
nand U13656 (N_13656,N_12088,N_12826);
or U13657 (N_13657,N_12788,N_12650);
nor U13658 (N_13658,N_12025,N_12765);
or U13659 (N_13659,N_12945,N_12564);
nor U13660 (N_13660,N_12114,N_12132);
xnor U13661 (N_13661,N_12396,N_12957);
xor U13662 (N_13662,N_12716,N_12991);
nand U13663 (N_13663,N_12010,N_12451);
xnor U13664 (N_13664,N_12779,N_12322);
nand U13665 (N_13665,N_12823,N_12816);
nor U13666 (N_13666,N_12701,N_12402);
nor U13667 (N_13667,N_12320,N_12593);
and U13668 (N_13668,N_12660,N_12353);
nand U13669 (N_13669,N_12244,N_12678);
and U13670 (N_13670,N_12418,N_12527);
nor U13671 (N_13671,N_12285,N_12015);
nor U13672 (N_13672,N_12988,N_12361);
nor U13673 (N_13673,N_12480,N_12969);
and U13674 (N_13674,N_12935,N_12670);
nor U13675 (N_13675,N_12850,N_12137);
or U13676 (N_13676,N_12710,N_12244);
nor U13677 (N_13677,N_12471,N_12613);
xor U13678 (N_13678,N_12250,N_12560);
and U13679 (N_13679,N_12084,N_12323);
or U13680 (N_13680,N_12331,N_12083);
and U13681 (N_13681,N_12051,N_12881);
nand U13682 (N_13682,N_12701,N_12062);
xor U13683 (N_13683,N_12969,N_12899);
nor U13684 (N_13684,N_12896,N_12730);
xnor U13685 (N_13685,N_12431,N_12227);
and U13686 (N_13686,N_12753,N_12590);
or U13687 (N_13687,N_12938,N_12134);
nand U13688 (N_13688,N_12378,N_12540);
or U13689 (N_13689,N_12981,N_12475);
nand U13690 (N_13690,N_12172,N_12116);
xnor U13691 (N_13691,N_12336,N_12095);
xor U13692 (N_13692,N_12562,N_12198);
and U13693 (N_13693,N_12743,N_12840);
xnor U13694 (N_13694,N_12037,N_12038);
xnor U13695 (N_13695,N_12724,N_12916);
xnor U13696 (N_13696,N_12344,N_12889);
nand U13697 (N_13697,N_12409,N_12259);
xnor U13698 (N_13698,N_12935,N_12450);
or U13699 (N_13699,N_12326,N_12931);
and U13700 (N_13700,N_12241,N_12835);
nand U13701 (N_13701,N_12538,N_12465);
nor U13702 (N_13702,N_12798,N_12855);
or U13703 (N_13703,N_12376,N_12553);
nor U13704 (N_13704,N_12581,N_12507);
or U13705 (N_13705,N_12032,N_12948);
and U13706 (N_13706,N_12537,N_12792);
nor U13707 (N_13707,N_12386,N_12965);
and U13708 (N_13708,N_12936,N_12100);
nor U13709 (N_13709,N_12004,N_12521);
xnor U13710 (N_13710,N_12037,N_12151);
or U13711 (N_13711,N_12112,N_12650);
or U13712 (N_13712,N_12555,N_12559);
or U13713 (N_13713,N_12816,N_12087);
nand U13714 (N_13714,N_12524,N_12009);
and U13715 (N_13715,N_12464,N_12607);
or U13716 (N_13716,N_12857,N_12220);
nand U13717 (N_13717,N_12036,N_12675);
xnor U13718 (N_13718,N_12450,N_12375);
nor U13719 (N_13719,N_12944,N_12818);
xor U13720 (N_13720,N_12345,N_12733);
and U13721 (N_13721,N_12634,N_12923);
xor U13722 (N_13722,N_12063,N_12511);
and U13723 (N_13723,N_12580,N_12043);
and U13724 (N_13724,N_12437,N_12527);
or U13725 (N_13725,N_12277,N_12655);
nand U13726 (N_13726,N_12128,N_12459);
nand U13727 (N_13727,N_12746,N_12457);
xor U13728 (N_13728,N_12221,N_12594);
and U13729 (N_13729,N_12509,N_12534);
or U13730 (N_13730,N_12726,N_12715);
nor U13731 (N_13731,N_12042,N_12452);
xor U13732 (N_13732,N_12423,N_12058);
or U13733 (N_13733,N_12423,N_12690);
or U13734 (N_13734,N_12044,N_12570);
and U13735 (N_13735,N_12047,N_12950);
or U13736 (N_13736,N_12689,N_12365);
and U13737 (N_13737,N_12766,N_12984);
xor U13738 (N_13738,N_12640,N_12726);
xnor U13739 (N_13739,N_12646,N_12940);
nor U13740 (N_13740,N_12884,N_12379);
nor U13741 (N_13741,N_12865,N_12228);
nand U13742 (N_13742,N_12908,N_12225);
xor U13743 (N_13743,N_12735,N_12560);
or U13744 (N_13744,N_12374,N_12424);
and U13745 (N_13745,N_12792,N_12292);
or U13746 (N_13746,N_12939,N_12667);
xnor U13747 (N_13747,N_12498,N_12404);
nand U13748 (N_13748,N_12222,N_12788);
nand U13749 (N_13749,N_12537,N_12117);
xor U13750 (N_13750,N_12230,N_12058);
and U13751 (N_13751,N_12294,N_12935);
or U13752 (N_13752,N_12775,N_12008);
nor U13753 (N_13753,N_12311,N_12433);
nor U13754 (N_13754,N_12140,N_12981);
and U13755 (N_13755,N_12561,N_12538);
nand U13756 (N_13756,N_12302,N_12078);
xor U13757 (N_13757,N_12148,N_12101);
and U13758 (N_13758,N_12160,N_12050);
and U13759 (N_13759,N_12364,N_12187);
nor U13760 (N_13760,N_12050,N_12906);
nand U13761 (N_13761,N_12565,N_12763);
nor U13762 (N_13762,N_12690,N_12191);
and U13763 (N_13763,N_12589,N_12689);
or U13764 (N_13764,N_12998,N_12135);
and U13765 (N_13765,N_12914,N_12188);
or U13766 (N_13766,N_12930,N_12678);
nand U13767 (N_13767,N_12358,N_12547);
nand U13768 (N_13768,N_12573,N_12970);
and U13769 (N_13769,N_12240,N_12424);
nor U13770 (N_13770,N_12259,N_12575);
nand U13771 (N_13771,N_12869,N_12324);
nor U13772 (N_13772,N_12209,N_12076);
nor U13773 (N_13773,N_12754,N_12066);
nand U13774 (N_13774,N_12778,N_12044);
or U13775 (N_13775,N_12223,N_12878);
or U13776 (N_13776,N_12782,N_12785);
and U13777 (N_13777,N_12976,N_12464);
xor U13778 (N_13778,N_12822,N_12736);
nand U13779 (N_13779,N_12306,N_12792);
nor U13780 (N_13780,N_12383,N_12895);
and U13781 (N_13781,N_12934,N_12609);
and U13782 (N_13782,N_12742,N_12791);
or U13783 (N_13783,N_12881,N_12133);
or U13784 (N_13784,N_12846,N_12197);
xor U13785 (N_13785,N_12310,N_12370);
and U13786 (N_13786,N_12194,N_12630);
nor U13787 (N_13787,N_12329,N_12544);
nor U13788 (N_13788,N_12767,N_12581);
or U13789 (N_13789,N_12176,N_12025);
or U13790 (N_13790,N_12681,N_12622);
nand U13791 (N_13791,N_12687,N_12626);
nor U13792 (N_13792,N_12152,N_12253);
nand U13793 (N_13793,N_12234,N_12649);
xor U13794 (N_13794,N_12968,N_12408);
nand U13795 (N_13795,N_12305,N_12077);
or U13796 (N_13796,N_12919,N_12183);
nand U13797 (N_13797,N_12667,N_12571);
xnor U13798 (N_13798,N_12993,N_12184);
nand U13799 (N_13799,N_12132,N_12075);
xnor U13800 (N_13800,N_12054,N_12652);
nand U13801 (N_13801,N_12686,N_12019);
and U13802 (N_13802,N_12016,N_12283);
or U13803 (N_13803,N_12387,N_12687);
and U13804 (N_13804,N_12369,N_12814);
nor U13805 (N_13805,N_12436,N_12997);
or U13806 (N_13806,N_12438,N_12275);
and U13807 (N_13807,N_12071,N_12003);
and U13808 (N_13808,N_12970,N_12866);
or U13809 (N_13809,N_12318,N_12970);
and U13810 (N_13810,N_12708,N_12321);
nor U13811 (N_13811,N_12189,N_12988);
and U13812 (N_13812,N_12649,N_12153);
and U13813 (N_13813,N_12553,N_12879);
nand U13814 (N_13814,N_12775,N_12694);
or U13815 (N_13815,N_12845,N_12007);
and U13816 (N_13816,N_12685,N_12566);
xnor U13817 (N_13817,N_12912,N_12607);
xor U13818 (N_13818,N_12701,N_12609);
xnor U13819 (N_13819,N_12975,N_12240);
or U13820 (N_13820,N_12720,N_12607);
or U13821 (N_13821,N_12474,N_12872);
nand U13822 (N_13822,N_12442,N_12620);
xor U13823 (N_13823,N_12262,N_12069);
nand U13824 (N_13824,N_12295,N_12888);
and U13825 (N_13825,N_12911,N_12770);
nand U13826 (N_13826,N_12906,N_12157);
nor U13827 (N_13827,N_12228,N_12136);
nand U13828 (N_13828,N_12205,N_12908);
or U13829 (N_13829,N_12721,N_12198);
nand U13830 (N_13830,N_12124,N_12009);
and U13831 (N_13831,N_12762,N_12665);
and U13832 (N_13832,N_12624,N_12509);
or U13833 (N_13833,N_12060,N_12065);
nor U13834 (N_13834,N_12436,N_12110);
or U13835 (N_13835,N_12649,N_12431);
xor U13836 (N_13836,N_12214,N_12529);
xnor U13837 (N_13837,N_12659,N_12211);
or U13838 (N_13838,N_12038,N_12327);
and U13839 (N_13839,N_12047,N_12472);
xnor U13840 (N_13840,N_12863,N_12213);
and U13841 (N_13841,N_12158,N_12258);
xnor U13842 (N_13842,N_12409,N_12325);
and U13843 (N_13843,N_12058,N_12768);
or U13844 (N_13844,N_12483,N_12122);
and U13845 (N_13845,N_12761,N_12070);
and U13846 (N_13846,N_12994,N_12491);
or U13847 (N_13847,N_12682,N_12930);
or U13848 (N_13848,N_12471,N_12041);
xnor U13849 (N_13849,N_12389,N_12853);
nand U13850 (N_13850,N_12732,N_12773);
or U13851 (N_13851,N_12304,N_12644);
nand U13852 (N_13852,N_12571,N_12518);
xnor U13853 (N_13853,N_12814,N_12175);
and U13854 (N_13854,N_12672,N_12198);
or U13855 (N_13855,N_12372,N_12848);
or U13856 (N_13856,N_12241,N_12108);
nand U13857 (N_13857,N_12394,N_12947);
and U13858 (N_13858,N_12322,N_12741);
or U13859 (N_13859,N_12836,N_12378);
or U13860 (N_13860,N_12873,N_12807);
nand U13861 (N_13861,N_12841,N_12234);
nor U13862 (N_13862,N_12866,N_12469);
or U13863 (N_13863,N_12501,N_12663);
or U13864 (N_13864,N_12656,N_12490);
nor U13865 (N_13865,N_12944,N_12101);
and U13866 (N_13866,N_12837,N_12555);
or U13867 (N_13867,N_12759,N_12050);
or U13868 (N_13868,N_12509,N_12200);
xnor U13869 (N_13869,N_12731,N_12964);
nor U13870 (N_13870,N_12680,N_12925);
nor U13871 (N_13871,N_12290,N_12246);
nor U13872 (N_13872,N_12374,N_12171);
nand U13873 (N_13873,N_12518,N_12834);
and U13874 (N_13874,N_12497,N_12168);
or U13875 (N_13875,N_12901,N_12995);
nor U13876 (N_13876,N_12192,N_12025);
nor U13877 (N_13877,N_12289,N_12901);
xnor U13878 (N_13878,N_12482,N_12976);
or U13879 (N_13879,N_12684,N_12359);
and U13880 (N_13880,N_12869,N_12303);
nand U13881 (N_13881,N_12000,N_12173);
and U13882 (N_13882,N_12430,N_12488);
nand U13883 (N_13883,N_12197,N_12058);
xor U13884 (N_13884,N_12744,N_12607);
or U13885 (N_13885,N_12922,N_12500);
and U13886 (N_13886,N_12357,N_12327);
nor U13887 (N_13887,N_12982,N_12727);
or U13888 (N_13888,N_12260,N_12436);
nand U13889 (N_13889,N_12558,N_12360);
or U13890 (N_13890,N_12296,N_12233);
or U13891 (N_13891,N_12315,N_12962);
nor U13892 (N_13892,N_12511,N_12554);
xnor U13893 (N_13893,N_12344,N_12736);
and U13894 (N_13894,N_12288,N_12472);
nand U13895 (N_13895,N_12687,N_12240);
nor U13896 (N_13896,N_12324,N_12122);
and U13897 (N_13897,N_12686,N_12846);
nand U13898 (N_13898,N_12341,N_12771);
or U13899 (N_13899,N_12939,N_12962);
or U13900 (N_13900,N_12079,N_12205);
xor U13901 (N_13901,N_12830,N_12951);
nor U13902 (N_13902,N_12013,N_12699);
nor U13903 (N_13903,N_12773,N_12780);
xor U13904 (N_13904,N_12591,N_12910);
nand U13905 (N_13905,N_12642,N_12727);
or U13906 (N_13906,N_12004,N_12311);
nor U13907 (N_13907,N_12039,N_12578);
nor U13908 (N_13908,N_12047,N_12621);
xor U13909 (N_13909,N_12867,N_12950);
or U13910 (N_13910,N_12393,N_12630);
nor U13911 (N_13911,N_12440,N_12048);
nor U13912 (N_13912,N_12140,N_12691);
or U13913 (N_13913,N_12946,N_12978);
xnor U13914 (N_13914,N_12561,N_12808);
and U13915 (N_13915,N_12494,N_12766);
nor U13916 (N_13916,N_12512,N_12520);
nor U13917 (N_13917,N_12347,N_12328);
and U13918 (N_13918,N_12353,N_12473);
nand U13919 (N_13919,N_12860,N_12516);
nor U13920 (N_13920,N_12255,N_12551);
nor U13921 (N_13921,N_12862,N_12683);
xnor U13922 (N_13922,N_12118,N_12279);
nor U13923 (N_13923,N_12013,N_12721);
nor U13924 (N_13924,N_12761,N_12912);
nor U13925 (N_13925,N_12902,N_12438);
nor U13926 (N_13926,N_12477,N_12201);
nand U13927 (N_13927,N_12815,N_12076);
or U13928 (N_13928,N_12167,N_12906);
nand U13929 (N_13929,N_12047,N_12203);
nor U13930 (N_13930,N_12306,N_12783);
nand U13931 (N_13931,N_12676,N_12161);
nor U13932 (N_13932,N_12472,N_12705);
nor U13933 (N_13933,N_12671,N_12308);
nand U13934 (N_13934,N_12849,N_12974);
or U13935 (N_13935,N_12193,N_12045);
or U13936 (N_13936,N_12124,N_12315);
nor U13937 (N_13937,N_12919,N_12209);
xor U13938 (N_13938,N_12123,N_12008);
and U13939 (N_13939,N_12989,N_12148);
nand U13940 (N_13940,N_12076,N_12414);
nand U13941 (N_13941,N_12878,N_12408);
or U13942 (N_13942,N_12420,N_12564);
and U13943 (N_13943,N_12387,N_12164);
or U13944 (N_13944,N_12167,N_12381);
xor U13945 (N_13945,N_12311,N_12979);
nor U13946 (N_13946,N_12819,N_12636);
and U13947 (N_13947,N_12993,N_12378);
nand U13948 (N_13948,N_12980,N_12609);
or U13949 (N_13949,N_12007,N_12711);
and U13950 (N_13950,N_12652,N_12212);
xor U13951 (N_13951,N_12896,N_12771);
xnor U13952 (N_13952,N_12911,N_12492);
or U13953 (N_13953,N_12050,N_12451);
xnor U13954 (N_13954,N_12489,N_12923);
xor U13955 (N_13955,N_12316,N_12475);
or U13956 (N_13956,N_12793,N_12965);
nor U13957 (N_13957,N_12436,N_12131);
or U13958 (N_13958,N_12496,N_12369);
nor U13959 (N_13959,N_12820,N_12242);
or U13960 (N_13960,N_12389,N_12790);
or U13961 (N_13961,N_12252,N_12182);
or U13962 (N_13962,N_12503,N_12938);
or U13963 (N_13963,N_12374,N_12690);
xor U13964 (N_13964,N_12097,N_12003);
or U13965 (N_13965,N_12950,N_12019);
or U13966 (N_13966,N_12631,N_12891);
nor U13967 (N_13967,N_12747,N_12983);
and U13968 (N_13968,N_12689,N_12267);
nand U13969 (N_13969,N_12877,N_12291);
nand U13970 (N_13970,N_12684,N_12253);
nor U13971 (N_13971,N_12395,N_12217);
and U13972 (N_13972,N_12668,N_12085);
nor U13973 (N_13973,N_12409,N_12392);
or U13974 (N_13974,N_12800,N_12868);
or U13975 (N_13975,N_12170,N_12553);
and U13976 (N_13976,N_12711,N_12990);
nand U13977 (N_13977,N_12068,N_12858);
nand U13978 (N_13978,N_12257,N_12813);
nor U13979 (N_13979,N_12343,N_12775);
and U13980 (N_13980,N_12379,N_12710);
nor U13981 (N_13981,N_12222,N_12864);
xor U13982 (N_13982,N_12582,N_12396);
xor U13983 (N_13983,N_12693,N_12348);
nor U13984 (N_13984,N_12097,N_12734);
and U13985 (N_13985,N_12402,N_12424);
or U13986 (N_13986,N_12585,N_12176);
xnor U13987 (N_13987,N_12647,N_12298);
xnor U13988 (N_13988,N_12429,N_12394);
and U13989 (N_13989,N_12024,N_12548);
xor U13990 (N_13990,N_12228,N_12239);
and U13991 (N_13991,N_12901,N_12431);
xnor U13992 (N_13992,N_12540,N_12850);
xnor U13993 (N_13993,N_12870,N_12808);
and U13994 (N_13994,N_12902,N_12422);
and U13995 (N_13995,N_12130,N_12657);
nor U13996 (N_13996,N_12749,N_12992);
nand U13997 (N_13997,N_12625,N_12109);
nand U13998 (N_13998,N_12272,N_12216);
and U13999 (N_13999,N_12091,N_12063);
nor U14000 (N_14000,N_13649,N_13757);
or U14001 (N_14001,N_13527,N_13759);
or U14002 (N_14002,N_13397,N_13915);
nor U14003 (N_14003,N_13404,N_13097);
xor U14004 (N_14004,N_13356,N_13230);
or U14005 (N_14005,N_13440,N_13232);
nor U14006 (N_14006,N_13401,N_13635);
or U14007 (N_14007,N_13675,N_13383);
nor U14008 (N_14008,N_13860,N_13767);
or U14009 (N_14009,N_13198,N_13720);
xor U14010 (N_14010,N_13507,N_13896);
xor U14011 (N_14011,N_13202,N_13526);
and U14012 (N_14012,N_13529,N_13856);
nand U14013 (N_14013,N_13602,N_13519);
nand U14014 (N_14014,N_13166,N_13567);
xor U14015 (N_14015,N_13056,N_13085);
or U14016 (N_14016,N_13384,N_13872);
and U14017 (N_14017,N_13191,N_13490);
nor U14018 (N_14018,N_13006,N_13487);
nor U14019 (N_14019,N_13695,N_13964);
and U14020 (N_14020,N_13800,N_13040);
and U14021 (N_14021,N_13375,N_13335);
and U14022 (N_14022,N_13647,N_13028);
or U14023 (N_14023,N_13072,N_13779);
nand U14024 (N_14024,N_13290,N_13659);
nand U14025 (N_14025,N_13359,N_13297);
and U14026 (N_14026,N_13851,N_13233);
nand U14027 (N_14027,N_13631,N_13911);
or U14028 (N_14028,N_13338,N_13607);
xnor U14029 (N_14029,N_13476,N_13839);
and U14030 (N_14030,N_13968,N_13765);
nor U14031 (N_14031,N_13782,N_13008);
and U14032 (N_14032,N_13343,N_13702);
xor U14033 (N_14033,N_13634,N_13271);
and U14034 (N_14034,N_13745,N_13474);
nand U14035 (N_14035,N_13471,N_13433);
and U14036 (N_14036,N_13127,N_13369);
or U14037 (N_14037,N_13798,N_13252);
and U14038 (N_14038,N_13566,N_13412);
nor U14039 (N_14039,N_13350,N_13158);
or U14040 (N_14040,N_13295,N_13497);
and U14041 (N_14041,N_13123,N_13156);
nor U14042 (N_14042,N_13391,N_13447);
and U14043 (N_14043,N_13900,N_13021);
and U14044 (N_14044,N_13106,N_13682);
xor U14045 (N_14045,N_13388,N_13540);
xnor U14046 (N_14046,N_13188,N_13481);
xnor U14047 (N_14047,N_13859,N_13374);
xor U14048 (N_14048,N_13030,N_13262);
or U14049 (N_14049,N_13841,N_13928);
nor U14050 (N_14050,N_13424,N_13064);
nor U14051 (N_14051,N_13340,N_13516);
xor U14052 (N_14052,N_13070,N_13220);
or U14053 (N_14053,N_13360,N_13962);
xnor U14054 (N_14054,N_13005,N_13362);
or U14055 (N_14055,N_13414,N_13931);
nor U14056 (N_14056,N_13605,N_13842);
nor U14057 (N_14057,N_13805,N_13808);
or U14058 (N_14058,N_13865,N_13498);
and U14059 (N_14059,N_13441,N_13026);
or U14060 (N_14060,N_13282,N_13472);
nor U14061 (N_14061,N_13336,N_13439);
nand U14062 (N_14062,N_13941,N_13129);
nand U14063 (N_14063,N_13585,N_13892);
xnor U14064 (N_14064,N_13190,N_13868);
or U14065 (N_14065,N_13742,N_13069);
or U14066 (N_14066,N_13312,N_13226);
nor U14067 (N_14067,N_13053,N_13109);
and U14068 (N_14068,N_13207,N_13803);
or U14069 (N_14069,N_13161,N_13752);
or U14070 (N_14070,N_13337,N_13991);
nand U14071 (N_14071,N_13133,N_13327);
nor U14072 (N_14072,N_13572,N_13815);
xnor U14073 (N_14073,N_13619,N_13598);
nand U14074 (N_14074,N_13591,N_13366);
nor U14075 (N_14075,N_13823,N_13972);
or U14076 (N_14076,N_13817,N_13453);
nor U14077 (N_14077,N_13912,N_13797);
or U14078 (N_14078,N_13780,N_13970);
or U14079 (N_14079,N_13907,N_13843);
nand U14080 (N_14080,N_13684,N_13183);
or U14081 (N_14081,N_13247,N_13750);
or U14082 (N_14082,N_13553,N_13764);
xnor U14083 (N_14083,N_13811,N_13050);
or U14084 (N_14084,N_13969,N_13743);
or U14085 (N_14085,N_13324,N_13216);
xor U14086 (N_14086,N_13382,N_13627);
or U14087 (N_14087,N_13041,N_13011);
or U14088 (N_14088,N_13470,N_13174);
xor U14089 (N_14089,N_13826,N_13950);
or U14090 (N_14090,N_13914,N_13814);
nor U14091 (N_14091,N_13318,N_13246);
xor U14092 (N_14092,N_13584,N_13038);
and U14093 (N_14093,N_13897,N_13426);
and U14094 (N_14094,N_13092,N_13079);
nand U14095 (N_14095,N_13073,N_13119);
or U14096 (N_14096,N_13259,N_13508);
nor U14097 (N_14097,N_13319,N_13863);
and U14098 (N_14098,N_13298,N_13523);
nor U14099 (N_14099,N_13870,N_13812);
and U14100 (N_14100,N_13217,N_13266);
nor U14101 (N_14101,N_13223,N_13613);
and U14102 (N_14102,N_13427,N_13367);
xnor U14103 (N_14103,N_13451,N_13754);
xor U14104 (N_14104,N_13082,N_13245);
and U14105 (N_14105,N_13637,N_13049);
or U14106 (N_14106,N_13945,N_13729);
nand U14107 (N_14107,N_13987,N_13052);
or U14108 (N_14108,N_13836,N_13229);
xnor U14109 (N_14109,N_13032,N_13726);
xor U14110 (N_14110,N_13313,N_13775);
xnor U14111 (N_14111,N_13199,N_13840);
nor U14112 (N_14112,N_13864,N_13978);
nand U14113 (N_14113,N_13227,N_13263);
or U14114 (N_14114,N_13284,N_13601);
nand U14115 (N_14115,N_13961,N_13075);
nand U14116 (N_14116,N_13825,N_13235);
nor U14117 (N_14117,N_13953,N_13339);
xnor U14118 (N_14118,N_13048,N_13186);
nand U14119 (N_14119,N_13551,N_13499);
xnor U14120 (N_14120,N_13162,N_13163);
nor U14121 (N_14121,N_13933,N_13813);
nand U14122 (N_14122,N_13436,N_13906);
or U14123 (N_14123,N_13379,N_13091);
and U14124 (N_14124,N_13938,N_13625);
and U14125 (N_14125,N_13442,N_13107);
nand U14126 (N_14126,N_13809,N_13086);
or U14127 (N_14127,N_13460,N_13228);
and U14128 (N_14128,N_13932,N_13205);
nor U14129 (N_14129,N_13110,N_13955);
xnor U14130 (N_14130,N_13787,N_13007);
and U14131 (N_14131,N_13940,N_13939);
and U14132 (N_14132,N_13322,N_13431);
nor U14133 (N_14133,N_13889,N_13373);
and U14134 (N_14134,N_13669,N_13878);
nand U14135 (N_14135,N_13801,N_13434);
or U14136 (N_14136,N_13467,N_13323);
xor U14137 (N_14137,N_13728,N_13795);
nor U14138 (N_14138,N_13965,N_13657);
or U14139 (N_14139,N_13673,N_13828);
xnor U14140 (N_14140,N_13589,N_13884);
and U14141 (N_14141,N_13763,N_13342);
and U14142 (N_14142,N_13714,N_13586);
xnor U14143 (N_14143,N_13116,N_13139);
nor U14144 (N_14144,N_13544,N_13381);
nor U14145 (N_14145,N_13164,N_13115);
and U14146 (N_14146,N_13098,N_13036);
nor U14147 (N_14147,N_13370,N_13985);
xor U14148 (N_14148,N_13268,N_13231);
or U14149 (N_14149,N_13628,N_13665);
nand U14150 (N_14150,N_13094,N_13389);
or U14151 (N_14151,N_13909,N_13794);
nor U14152 (N_14152,N_13448,N_13495);
or U14153 (N_14153,N_13988,N_13020);
and U14154 (N_14154,N_13265,N_13352);
xnor U14155 (N_14155,N_13993,N_13305);
nand U14156 (N_14156,N_13449,N_13380);
xnor U14157 (N_14157,N_13926,N_13744);
or U14158 (N_14158,N_13640,N_13415);
or U14159 (N_14159,N_13833,N_13432);
nor U14160 (N_14160,N_13755,N_13446);
nand U14161 (N_14161,N_13942,N_13212);
nor U14162 (N_14162,N_13850,N_13936);
xnor U14163 (N_14163,N_13676,N_13986);
nand U14164 (N_14164,N_13582,N_13749);
and U14165 (N_14165,N_13893,N_13571);
nand U14166 (N_14166,N_13234,N_13479);
nor U14167 (N_14167,N_13332,N_13542);
nand U14168 (N_14168,N_13416,N_13653);
nand U14169 (N_14169,N_13705,N_13514);
nand U14170 (N_14170,N_13902,N_13810);
and U14171 (N_14171,N_13730,N_13488);
and U14172 (N_14172,N_13108,N_13089);
or U14173 (N_14173,N_13179,N_13707);
and U14174 (N_14174,N_13237,N_13771);
xnor U14175 (N_14175,N_13361,N_13600);
nand U14176 (N_14176,N_13286,N_13983);
or U14177 (N_14177,N_13022,N_13088);
nand U14178 (N_14178,N_13661,N_13610);
nand U14179 (N_14179,N_13390,N_13114);
xnor U14180 (N_14180,N_13643,N_13518);
xnor U14181 (N_14181,N_13563,N_13832);
and U14182 (N_14182,N_13505,N_13587);
or U14183 (N_14183,N_13952,N_13943);
and U14184 (N_14184,N_13078,N_13385);
nor U14185 (N_14185,N_13395,N_13666);
nor U14186 (N_14186,N_13096,N_13456);
nand U14187 (N_14187,N_13009,N_13054);
nor U14188 (N_14188,N_13792,N_13105);
nor U14189 (N_14189,N_13579,N_13748);
and U14190 (N_14190,N_13308,N_13364);
and U14191 (N_14191,N_13218,N_13534);
nor U14192 (N_14192,N_13672,N_13292);
or U14193 (N_14193,N_13269,N_13222);
or U14194 (N_14194,N_13686,N_13113);
xnor U14195 (N_14195,N_13504,N_13716);
or U14196 (N_14196,N_13291,N_13916);
xnor U14197 (N_14197,N_13816,N_13559);
and U14198 (N_14198,N_13111,N_13713);
or U14199 (N_14199,N_13777,N_13080);
nand U14200 (N_14200,N_13248,N_13894);
nor U14201 (N_14201,N_13303,N_13590);
xor U14202 (N_14202,N_13733,N_13066);
nor U14203 (N_14203,N_13844,N_13622);
nor U14204 (N_14204,N_13554,N_13651);
nand U14205 (N_14205,N_13946,N_13310);
xnor U14206 (N_14206,N_13132,N_13924);
xor U14207 (N_14207,N_13890,N_13561);
or U14208 (N_14208,N_13063,N_13219);
and U14209 (N_14209,N_13494,N_13157);
xor U14210 (N_14210,N_13029,N_13664);
and U14211 (N_14211,N_13013,N_13326);
and U14212 (N_14212,N_13573,N_13173);
nor U14213 (N_14213,N_13354,N_13934);
and U14214 (N_14214,N_13947,N_13535);
and U14215 (N_14215,N_13493,N_13891);
or U14216 (N_14216,N_13211,N_13899);
nor U14217 (N_14217,N_13037,N_13454);
or U14218 (N_14218,N_13685,N_13908);
or U14219 (N_14219,N_13429,N_13221);
xnor U14220 (N_14220,N_13057,N_13376);
and U14221 (N_14221,N_13464,N_13425);
xnor U14222 (N_14222,N_13549,N_13254);
xor U14223 (N_14223,N_13615,N_13709);
nand U14224 (N_14224,N_13790,N_13606);
xor U14225 (N_14225,N_13781,N_13570);
xor U14226 (N_14226,N_13387,N_13071);
nand U14227 (N_14227,N_13102,N_13827);
or U14228 (N_14228,N_13660,N_13363);
nand U14229 (N_14229,N_13949,N_13569);
or U14230 (N_14230,N_13294,N_13276);
nand U14231 (N_14231,N_13960,N_13999);
or U14232 (N_14232,N_13927,N_13521);
nand U14233 (N_14233,N_13545,N_13314);
nor U14234 (N_14234,N_13746,N_13239);
xor U14235 (N_14235,N_13948,N_13128);
xnor U14236 (N_14236,N_13578,N_13473);
xor U14237 (N_14237,N_13623,N_13528);
nor U14238 (N_14238,N_13648,N_13565);
and U14239 (N_14239,N_13146,N_13918);
or U14240 (N_14240,N_13512,N_13737);
xor U14241 (N_14241,N_13923,N_13193);
and U14242 (N_14242,N_13751,N_13621);
nand U14243 (N_14243,N_13277,N_13592);
xnor U14244 (N_14244,N_13365,N_13861);
nor U14245 (N_14245,N_13122,N_13419);
and U14246 (N_14246,N_13981,N_13853);
nand U14247 (N_14247,N_13806,N_13719);
xor U14248 (N_14248,N_13989,N_13616);
xnor U14249 (N_14249,N_13555,N_13099);
and U14250 (N_14250,N_13921,N_13770);
nand U14251 (N_14251,N_13074,N_13315);
and U14252 (N_14252,N_13944,N_13185);
nand U14253 (N_14253,N_13153,N_13541);
and U14254 (N_14254,N_13047,N_13533);
nand U14255 (N_14255,N_13210,N_13300);
nor U14256 (N_14256,N_13980,N_13090);
and U14257 (N_14257,N_13061,N_13140);
xnor U14258 (N_14258,N_13910,N_13402);
nand U14259 (N_14259,N_13289,N_13329);
or U14260 (N_14260,N_13929,N_13898);
or U14261 (N_14261,N_13468,N_13019);
nor U14262 (N_14262,N_13261,N_13724);
nand U14263 (N_14263,N_13564,N_13557);
nand U14264 (N_14264,N_13694,N_13148);
and U14265 (N_14265,N_13137,N_13510);
and U14266 (N_14266,N_13055,N_13633);
xor U14267 (N_14267,N_13594,N_13243);
nor U14268 (N_14268,N_13485,N_13285);
xnor U14269 (N_14269,N_13762,N_13975);
nor U14270 (N_14270,N_13309,N_13979);
and U14271 (N_14271,N_13560,N_13882);
nand U14272 (N_14272,N_13124,N_13881);
or U14273 (N_14273,N_13786,N_13636);
nand U14274 (N_14274,N_13428,N_13182);
nand U14275 (N_14275,N_13144,N_13321);
or U14276 (N_14276,N_13278,N_13283);
or U14277 (N_14277,N_13524,N_13334);
or U14278 (N_14278,N_13195,N_13435);
or U14279 (N_14279,N_13093,N_13568);
xor U14280 (N_14280,N_13793,N_13922);
and U14281 (N_14281,N_13293,N_13215);
xor U14282 (N_14282,N_13583,N_13491);
or U14283 (N_14283,N_13525,N_13152);
or U14284 (N_14284,N_13689,N_13760);
xor U14285 (N_14285,N_13679,N_13406);
nor U14286 (N_14286,N_13413,N_13735);
or U14287 (N_14287,N_13977,N_13465);
nand U14288 (N_14288,N_13353,N_13027);
xor U14289 (N_14289,N_13717,N_13176);
and U14290 (N_14290,N_13393,N_13358);
nand U14291 (N_14291,N_13046,N_13196);
nor U14292 (N_14292,N_13469,N_13788);
nor U14293 (N_14293,N_13024,N_13995);
and U14294 (N_14294,N_13203,N_13400);
or U14295 (N_14295,N_13577,N_13873);
or U14296 (N_14296,N_13200,N_13270);
nand U14297 (N_14297,N_13224,N_13194);
nor U14298 (N_14298,N_13444,N_13804);
and U14299 (N_14299,N_13260,N_13010);
nor U14300 (N_14300,N_13895,N_13250);
nand U14301 (N_14301,N_13725,N_13480);
or U14302 (N_14302,N_13104,N_13511);
xnor U14303 (N_14303,N_13160,N_13917);
xnor U14304 (N_14304,N_13189,N_13147);
nor U14305 (N_14305,N_13045,N_13708);
xor U14306 (N_14306,N_13421,N_13645);
nor U14307 (N_14307,N_13062,N_13789);
xnor U14308 (N_14308,N_13688,N_13548);
xor U14309 (N_14309,N_13409,N_13802);
xnor U14310 (N_14310,N_13067,N_13703);
and U14311 (N_14311,N_13656,N_13001);
nand U14312 (N_14312,N_13680,N_13576);
nand U14313 (N_14313,N_13149,N_13349);
nor U14314 (N_14314,N_13638,N_13483);
nand U14315 (N_14315,N_13671,N_13112);
and U14316 (N_14316,N_13697,N_13117);
nand U14317 (N_14317,N_13831,N_13463);
or U14318 (N_14318,N_13065,N_13662);
xnor U14319 (N_14319,N_13723,N_13954);
nor U14320 (N_14320,N_13502,N_13867);
nor U14321 (N_14321,N_13394,N_13888);
and U14322 (N_14322,N_13766,N_13547);
nand U14323 (N_14323,N_13768,N_13003);
or U14324 (N_14324,N_13126,N_13718);
nand U14325 (N_14325,N_13087,N_13642);
or U14326 (N_14326,N_13783,N_13994);
nor U14327 (N_14327,N_13971,N_13935);
xor U14328 (N_14328,N_13145,N_13458);
and U14329 (N_14329,N_13058,N_13438);
or U14330 (N_14330,N_13320,N_13399);
nand U14331 (N_14331,N_13866,N_13509);
and U14332 (N_14332,N_13345,N_13883);
xnor U14333 (N_14333,N_13253,N_13484);
and U14334 (N_14334,N_13609,N_13593);
nand U14335 (N_14335,N_13875,N_13251);
nand U14336 (N_14336,N_13304,N_13819);
or U14337 (N_14337,N_13151,N_13101);
nor U14338 (N_14338,N_13236,N_13175);
or U14339 (N_14339,N_13597,N_13997);
nor U14340 (N_14340,N_13588,N_13410);
nand U14341 (N_14341,N_13347,N_13240);
or U14342 (N_14342,N_13847,N_13747);
xor U14343 (N_14343,N_13919,N_13837);
nor U14344 (N_14344,N_13711,N_13558);
and U14345 (N_14345,N_13154,N_13886);
nor U14346 (N_14346,N_13887,N_13131);
nor U14347 (N_14347,N_13034,N_13552);
nor U14348 (N_14348,N_13614,N_13462);
and U14349 (N_14349,N_13655,N_13698);
xnor U14350 (N_14350,N_13807,N_13279);
nand U14351 (N_14351,N_13307,N_13341);
and U14352 (N_14352,N_13522,N_13515);
or U14353 (N_14353,N_13187,N_13876);
nand U14354 (N_14354,N_13604,N_13691);
xor U14355 (N_14355,N_13172,N_13134);
and U14356 (N_14356,N_13258,N_13141);
xnor U14357 (N_14357,N_13017,N_13517);
nor U14358 (N_14358,N_13901,N_13181);
nand U14359 (N_14359,N_13773,N_13838);
or U14360 (N_14360,N_13443,N_13328);
or U14361 (N_14361,N_13753,N_13885);
nand U14362 (N_14362,N_13903,N_13772);
xor U14363 (N_14363,N_13739,N_13854);
and U14364 (N_14364,N_13125,N_13608);
xnor U14365 (N_14365,N_13031,N_13721);
nand U14366 (N_14366,N_13958,N_13641);
nor U14367 (N_14367,N_13599,N_13184);
or U14368 (N_14368,N_13155,N_13344);
and U14369 (N_14369,N_13192,N_13492);
or U14370 (N_14370,N_13244,N_13632);
nor U14371 (N_14371,N_13877,N_13242);
nor U14372 (N_14372,N_13357,N_13241);
nor U14373 (N_14373,N_13758,N_13171);
or U14374 (N_14374,N_13818,N_13626);
nand U14375 (N_14375,N_13165,N_13209);
nor U14376 (N_14376,N_13678,N_13059);
and U14377 (N_14377,N_13422,N_13355);
xor U14378 (N_14378,N_13043,N_13450);
xnor U14379 (N_14379,N_13976,N_13734);
nor U14380 (N_14380,N_13581,N_13503);
nand U14381 (N_14381,N_13225,N_13249);
nor U14382 (N_14382,N_13774,N_13820);
nand U14383 (N_14383,N_13274,N_13084);
nor U14384 (N_14384,N_13068,N_13741);
and U14385 (N_14385,N_13317,N_13411);
nand U14386 (N_14386,N_13513,N_13998);
nor U14387 (N_14387,N_13377,N_13799);
xnor U14388 (N_14388,N_13862,N_13051);
and U14389 (N_14389,N_13667,N_13120);
or U14390 (N_14390,N_13857,N_13348);
or U14391 (N_14391,N_13296,N_13620);
nor U14392 (N_14392,N_13420,N_13858);
nor U14393 (N_14393,N_13974,N_13466);
nand U14394 (N_14394,N_13208,N_13835);
nor U14395 (N_14395,N_13596,N_13407);
and U14396 (N_14396,N_13612,N_13550);
and U14397 (N_14397,N_13452,N_13658);
and U14398 (N_14398,N_13869,N_13142);
or U14399 (N_14399,N_13712,N_13333);
or U14400 (N_14400,N_13683,N_13267);
xnor U14401 (N_14401,N_13796,N_13992);
nand U14402 (N_14402,N_13905,N_13701);
nor U14403 (N_14403,N_13670,N_13537);
and U14404 (N_14404,N_13913,N_13871);
nor U14405 (N_14405,N_13042,N_13238);
xnor U14406 (N_14406,N_13973,N_13201);
or U14407 (N_14407,N_13214,N_13081);
nor U14408 (N_14408,N_13966,N_13538);
or U14409 (N_14409,N_13178,N_13699);
nand U14410 (N_14410,N_13461,N_13874);
and U14411 (N_14411,N_13879,N_13287);
nor U14412 (N_14412,N_13710,N_13392);
or U14413 (N_14413,N_13784,N_13693);
nand U14414 (N_14414,N_13496,N_13299);
or U14415 (N_14415,N_13417,N_13846);
nand U14416 (N_14416,N_13311,N_13617);
and U14417 (N_14417,N_13372,N_13012);
xnor U14418 (N_14418,N_13834,N_13197);
and U14419 (N_14419,N_13168,N_13180);
xnor U14420 (N_14420,N_13824,N_13256);
or U14421 (N_14421,N_13982,N_13845);
xnor U14422 (N_14422,N_13506,N_13378);
or U14423 (N_14423,N_13785,N_13306);
nor U14424 (N_14424,N_13580,N_13769);
nand U14425 (N_14425,N_13677,N_13083);
nand U14426 (N_14426,N_13996,N_13130);
or U14427 (N_14427,N_13732,N_13692);
or U14428 (N_14428,N_13937,N_13967);
nand U14429 (N_14429,N_13556,N_13077);
and U14430 (N_14430,N_13629,N_13100);
nand U14431 (N_14431,N_13095,N_13076);
nor U14432 (N_14432,N_13281,N_13408);
or U14433 (N_14433,N_13302,N_13004);
nor U14434 (N_14434,N_13025,N_13275);
or U14435 (N_14435,N_13489,N_13272);
or U14436 (N_14436,N_13206,N_13630);
xnor U14437 (N_14437,N_13423,N_13700);
xnor U14438 (N_14438,N_13368,N_13830);
nor U14439 (N_14439,N_13169,N_13951);
and U14440 (N_14440,N_13213,N_13486);
and U14441 (N_14441,N_13681,N_13475);
xnor U14442 (N_14442,N_13756,N_13855);
or U14443 (N_14443,N_13445,N_13103);
nor U14444 (N_14444,N_13644,N_13500);
xnor U14445 (N_14445,N_13396,N_13990);
and U14446 (N_14446,N_13136,N_13477);
nor U14447 (N_14447,N_13204,N_13706);
nor U14448 (N_14448,N_13791,N_13135);
nor U14449 (N_14449,N_13531,N_13925);
nor U14450 (N_14450,N_13959,N_13740);
xnor U14451 (N_14451,N_13654,N_13650);
nor U14452 (N_14452,N_13646,N_13437);
nor U14453 (N_14453,N_13727,N_13738);
nand U14454 (N_14454,N_13674,N_13562);
nor U14455 (N_14455,N_13000,N_13595);
xnor U14456 (N_14456,N_13543,N_13849);
xnor U14457 (N_14457,N_13920,N_13039);
and U14458 (N_14458,N_13351,N_13418);
nand U14459 (N_14459,N_13715,N_13023);
or U14460 (N_14460,N_13829,N_13687);
nand U14461 (N_14461,N_13530,N_13690);
xor U14462 (N_14462,N_13457,N_13264);
nand U14463 (N_14463,N_13167,N_13482);
xor U14464 (N_14464,N_13611,N_13536);
or U14465 (N_14465,N_13118,N_13546);
nand U14466 (N_14466,N_13403,N_13159);
or U14467 (N_14467,N_13060,N_13273);
and U14468 (N_14468,N_13018,N_13016);
xnor U14469 (N_14469,N_13002,N_13956);
nand U14470 (N_14470,N_13736,N_13405);
nor U14471 (N_14471,N_13984,N_13822);
or U14472 (N_14472,N_13663,N_13330);
nor U14473 (N_14473,N_13668,N_13778);
nand U14474 (N_14474,N_13257,N_13624);
or U14475 (N_14475,N_13704,N_13346);
nor U14476 (N_14476,N_13574,N_13280);
nor U14477 (N_14477,N_13386,N_13014);
xnor U14478 (N_14478,N_13575,N_13138);
or U14479 (N_14479,N_13652,N_13957);
nand U14480 (N_14480,N_13618,N_13821);
nor U14481 (N_14481,N_13170,N_13015);
or U14482 (N_14482,N_13963,N_13603);
nand U14483 (N_14483,N_13880,N_13478);
nand U14484 (N_14484,N_13639,N_13430);
or U14485 (N_14485,N_13150,N_13761);
nand U14486 (N_14486,N_13044,N_13398);
xnor U14487 (N_14487,N_13776,N_13848);
nor U14488 (N_14488,N_13731,N_13904);
xor U14489 (N_14489,N_13696,N_13852);
nor U14490 (N_14490,N_13035,N_13301);
or U14491 (N_14491,N_13459,N_13520);
xor U14492 (N_14492,N_13539,N_13455);
or U14493 (N_14493,N_13501,N_13143);
nor U14494 (N_14494,N_13331,N_13532);
and U14495 (N_14495,N_13371,N_13121);
xor U14496 (N_14496,N_13930,N_13255);
nor U14497 (N_14497,N_13288,N_13722);
nand U14498 (N_14498,N_13177,N_13325);
and U14499 (N_14499,N_13316,N_13033);
or U14500 (N_14500,N_13254,N_13098);
nand U14501 (N_14501,N_13854,N_13383);
nand U14502 (N_14502,N_13449,N_13646);
nor U14503 (N_14503,N_13009,N_13179);
xnor U14504 (N_14504,N_13007,N_13415);
nor U14505 (N_14505,N_13644,N_13099);
xnor U14506 (N_14506,N_13645,N_13569);
or U14507 (N_14507,N_13455,N_13937);
and U14508 (N_14508,N_13530,N_13323);
or U14509 (N_14509,N_13835,N_13894);
nand U14510 (N_14510,N_13373,N_13289);
xor U14511 (N_14511,N_13157,N_13173);
nor U14512 (N_14512,N_13100,N_13981);
and U14513 (N_14513,N_13566,N_13802);
and U14514 (N_14514,N_13830,N_13602);
or U14515 (N_14515,N_13929,N_13539);
nor U14516 (N_14516,N_13942,N_13803);
nor U14517 (N_14517,N_13985,N_13546);
nand U14518 (N_14518,N_13895,N_13286);
nand U14519 (N_14519,N_13779,N_13862);
xor U14520 (N_14520,N_13469,N_13403);
and U14521 (N_14521,N_13597,N_13445);
nor U14522 (N_14522,N_13344,N_13090);
nand U14523 (N_14523,N_13931,N_13385);
nand U14524 (N_14524,N_13829,N_13146);
or U14525 (N_14525,N_13256,N_13318);
nand U14526 (N_14526,N_13147,N_13994);
and U14527 (N_14527,N_13092,N_13052);
and U14528 (N_14528,N_13247,N_13894);
nand U14529 (N_14529,N_13951,N_13503);
xnor U14530 (N_14530,N_13050,N_13150);
xor U14531 (N_14531,N_13726,N_13029);
and U14532 (N_14532,N_13578,N_13962);
nor U14533 (N_14533,N_13171,N_13042);
xor U14534 (N_14534,N_13329,N_13605);
and U14535 (N_14535,N_13697,N_13977);
or U14536 (N_14536,N_13370,N_13422);
and U14537 (N_14537,N_13356,N_13685);
or U14538 (N_14538,N_13433,N_13792);
or U14539 (N_14539,N_13834,N_13280);
and U14540 (N_14540,N_13461,N_13675);
or U14541 (N_14541,N_13026,N_13258);
or U14542 (N_14542,N_13299,N_13323);
xnor U14543 (N_14543,N_13642,N_13545);
and U14544 (N_14544,N_13012,N_13813);
or U14545 (N_14545,N_13422,N_13449);
or U14546 (N_14546,N_13855,N_13371);
and U14547 (N_14547,N_13620,N_13468);
nand U14548 (N_14548,N_13069,N_13659);
nand U14549 (N_14549,N_13141,N_13378);
or U14550 (N_14550,N_13299,N_13329);
and U14551 (N_14551,N_13648,N_13050);
and U14552 (N_14552,N_13811,N_13376);
or U14553 (N_14553,N_13258,N_13751);
nor U14554 (N_14554,N_13822,N_13333);
xor U14555 (N_14555,N_13999,N_13480);
nand U14556 (N_14556,N_13974,N_13887);
or U14557 (N_14557,N_13224,N_13142);
xnor U14558 (N_14558,N_13929,N_13529);
xnor U14559 (N_14559,N_13686,N_13432);
and U14560 (N_14560,N_13008,N_13416);
or U14561 (N_14561,N_13278,N_13072);
nor U14562 (N_14562,N_13462,N_13601);
nand U14563 (N_14563,N_13561,N_13752);
and U14564 (N_14564,N_13345,N_13536);
nor U14565 (N_14565,N_13364,N_13920);
or U14566 (N_14566,N_13641,N_13485);
xor U14567 (N_14567,N_13015,N_13526);
xor U14568 (N_14568,N_13631,N_13244);
xor U14569 (N_14569,N_13147,N_13363);
nor U14570 (N_14570,N_13460,N_13234);
xor U14571 (N_14571,N_13311,N_13233);
nand U14572 (N_14572,N_13336,N_13326);
and U14573 (N_14573,N_13418,N_13410);
and U14574 (N_14574,N_13378,N_13138);
xnor U14575 (N_14575,N_13895,N_13858);
and U14576 (N_14576,N_13252,N_13753);
nor U14577 (N_14577,N_13918,N_13035);
or U14578 (N_14578,N_13828,N_13797);
xor U14579 (N_14579,N_13374,N_13655);
nor U14580 (N_14580,N_13226,N_13778);
nor U14581 (N_14581,N_13602,N_13777);
nor U14582 (N_14582,N_13061,N_13284);
xor U14583 (N_14583,N_13080,N_13842);
and U14584 (N_14584,N_13090,N_13081);
or U14585 (N_14585,N_13914,N_13566);
xor U14586 (N_14586,N_13899,N_13928);
nor U14587 (N_14587,N_13212,N_13980);
nor U14588 (N_14588,N_13867,N_13574);
nor U14589 (N_14589,N_13789,N_13923);
and U14590 (N_14590,N_13484,N_13926);
or U14591 (N_14591,N_13507,N_13584);
nand U14592 (N_14592,N_13603,N_13258);
xor U14593 (N_14593,N_13659,N_13557);
nand U14594 (N_14594,N_13120,N_13104);
and U14595 (N_14595,N_13164,N_13447);
xor U14596 (N_14596,N_13180,N_13396);
xor U14597 (N_14597,N_13841,N_13981);
and U14598 (N_14598,N_13845,N_13338);
xor U14599 (N_14599,N_13754,N_13672);
and U14600 (N_14600,N_13329,N_13237);
nand U14601 (N_14601,N_13906,N_13892);
xor U14602 (N_14602,N_13732,N_13556);
xor U14603 (N_14603,N_13279,N_13381);
or U14604 (N_14604,N_13229,N_13536);
and U14605 (N_14605,N_13956,N_13489);
nand U14606 (N_14606,N_13824,N_13846);
or U14607 (N_14607,N_13367,N_13755);
and U14608 (N_14608,N_13914,N_13310);
and U14609 (N_14609,N_13565,N_13899);
nand U14610 (N_14610,N_13172,N_13617);
xnor U14611 (N_14611,N_13594,N_13330);
nor U14612 (N_14612,N_13301,N_13199);
or U14613 (N_14613,N_13438,N_13432);
nor U14614 (N_14614,N_13701,N_13776);
xnor U14615 (N_14615,N_13575,N_13950);
nand U14616 (N_14616,N_13297,N_13821);
nor U14617 (N_14617,N_13785,N_13217);
nand U14618 (N_14618,N_13974,N_13132);
nand U14619 (N_14619,N_13578,N_13636);
xor U14620 (N_14620,N_13638,N_13125);
xor U14621 (N_14621,N_13673,N_13886);
and U14622 (N_14622,N_13946,N_13779);
nand U14623 (N_14623,N_13077,N_13204);
xor U14624 (N_14624,N_13958,N_13451);
nand U14625 (N_14625,N_13462,N_13167);
nor U14626 (N_14626,N_13256,N_13314);
nor U14627 (N_14627,N_13920,N_13579);
and U14628 (N_14628,N_13034,N_13459);
nand U14629 (N_14629,N_13109,N_13383);
or U14630 (N_14630,N_13479,N_13948);
nor U14631 (N_14631,N_13246,N_13294);
and U14632 (N_14632,N_13359,N_13162);
or U14633 (N_14633,N_13395,N_13053);
or U14634 (N_14634,N_13831,N_13723);
nor U14635 (N_14635,N_13348,N_13806);
and U14636 (N_14636,N_13155,N_13474);
or U14637 (N_14637,N_13538,N_13878);
nand U14638 (N_14638,N_13884,N_13129);
xor U14639 (N_14639,N_13445,N_13532);
nand U14640 (N_14640,N_13034,N_13324);
nor U14641 (N_14641,N_13220,N_13079);
or U14642 (N_14642,N_13292,N_13746);
nand U14643 (N_14643,N_13235,N_13903);
and U14644 (N_14644,N_13051,N_13632);
or U14645 (N_14645,N_13952,N_13974);
and U14646 (N_14646,N_13418,N_13527);
nor U14647 (N_14647,N_13756,N_13474);
xor U14648 (N_14648,N_13459,N_13527);
xnor U14649 (N_14649,N_13191,N_13946);
or U14650 (N_14650,N_13663,N_13404);
nand U14651 (N_14651,N_13595,N_13775);
nand U14652 (N_14652,N_13815,N_13291);
nand U14653 (N_14653,N_13961,N_13102);
xnor U14654 (N_14654,N_13917,N_13890);
nand U14655 (N_14655,N_13798,N_13757);
nor U14656 (N_14656,N_13995,N_13441);
xor U14657 (N_14657,N_13228,N_13727);
nor U14658 (N_14658,N_13921,N_13045);
nor U14659 (N_14659,N_13530,N_13283);
nor U14660 (N_14660,N_13426,N_13056);
nand U14661 (N_14661,N_13353,N_13012);
or U14662 (N_14662,N_13073,N_13903);
and U14663 (N_14663,N_13503,N_13826);
or U14664 (N_14664,N_13685,N_13264);
and U14665 (N_14665,N_13748,N_13032);
nand U14666 (N_14666,N_13495,N_13035);
and U14667 (N_14667,N_13191,N_13412);
or U14668 (N_14668,N_13349,N_13833);
nand U14669 (N_14669,N_13491,N_13465);
nand U14670 (N_14670,N_13417,N_13165);
or U14671 (N_14671,N_13650,N_13639);
xor U14672 (N_14672,N_13586,N_13050);
nand U14673 (N_14673,N_13485,N_13574);
nand U14674 (N_14674,N_13316,N_13358);
xor U14675 (N_14675,N_13369,N_13977);
and U14676 (N_14676,N_13160,N_13508);
and U14677 (N_14677,N_13363,N_13585);
xnor U14678 (N_14678,N_13312,N_13854);
nor U14679 (N_14679,N_13500,N_13035);
xnor U14680 (N_14680,N_13747,N_13620);
or U14681 (N_14681,N_13626,N_13021);
or U14682 (N_14682,N_13194,N_13123);
nor U14683 (N_14683,N_13865,N_13511);
nor U14684 (N_14684,N_13140,N_13335);
nor U14685 (N_14685,N_13677,N_13135);
xor U14686 (N_14686,N_13091,N_13005);
xor U14687 (N_14687,N_13207,N_13127);
or U14688 (N_14688,N_13846,N_13471);
xor U14689 (N_14689,N_13589,N_13410);
or U14690 (N_14690,N_13534,N_13075);
or U14691 (N_14691,N_13369,N_13692);
nor U14692 (N_14692,N_13053,N_13088);
and U14693 (N_14693,N_13242,N_13802);
and U14694 (N_14694,N_13717,N_13771);
or U14695 (N_14695,N_13675,N_13719);
and U14696 (N_14696,N_13035,N_13853);
and U14697 (N_14697,N_13243,N_13286);
nor U14698 (N_14698,N_13432,N_13063);
nor U14699 (N_14699,N_13087,N_13699);
and U14700 (N_14700,N_13610,N_13530);
nand U14701 (N_14701,N_13079,N_13550);
xnor U14702 (N_14702,N_13636,N_13635);
or U14703 (N_14703,N_13350,N_13095);
xor U14704 (N_14704,N_13326,N_13813);
or U14705 (N_14705,N_13978,N_13894);
xnor U14706 (N_14706,N_13876,N_13777);
nand U14707 (N_14707,N_13516,N_13545);
or U14708 (N_14708,N_13826,N_13486);
nand U14709 (N_14709,N_13217,N_13724);
and U14710 (N_14710,N_13330,N_13920);
and U14711 (N_14711,N_13393,N_13444);
nor U14712 (N_14712,N_13410,N_13934);
and U14713 (N_14713,N_13055,N_13657);
xnor U14714 (N_14714,N_13629,N_13756);
nor U14715 (N_14715,N_13957,N_13509);
nor U14716 (N_14716,N_13721,N_13434);
and U14717 (N_14717,N_13328,N_13901);
nand U14718 (N_14718,N_13919,N_13299);
xor U14719 (N_14719,N_13301,N_13476);
nor U14720 (N_14720,N_13713,N_13962);
xnor U14721 (N_14721,N_13259,N_13309);
nand U14722 (N_14722,N_13735,N_13544);
or U14723 (N_14723,N_13119,N_13901);
nand U14724 (N_14724,N_13573,N_13822);
nand U14725 (N_14725,N_13171,N_13203);
or U14726 (N_14726,N_13238,N_13504);
nand U14727 (N_14727,N_13218,N_13428);
and U14728 (N_14728,N_13177,N_13033);
nand U14729 (N_14729,N_13396,N_13930);
nand U14730 (N_14730,N_13916,N_13093);
nor U14731 (N_14731,N_13322,N_13175);
and U14732 (N_14732,N_13641,N_13348);
or U14733 (N_14733,N_13336,N_13211);
nor U14734 (N_14734,N_13209,N_13806);
nor U14735 (N_14735,N_13094,N_13428);
nand U14736 (N_14736,N_13253,N_13650);
nor U14737 (N_14737,N_13575,N_13639);
nand U14738 (N_14738,N_13707,N_13966);
or U14739 (N_14739,N_13411,N_13732);
and U14740 (N_14740,N_13788,N_13911);
and U14741 (N_14741,N_13819,N_13349);
nor U14742 (N_14742,N_13366,N_13593);
and U14743 (N_14743,N_13805,N_13191);
nor U14744 (N_14744,N_13697,N_13754);
or U14745 (N_14745,N_13067,N_13158);
xnor U14746 (N_14746,N_13801,N_13908);
or U14747 (N_14747,N_13767,N_13981);
or U14748 (N_14748,N_13902,N_13384);
xnor U14749 (N_14749,N_13290,N_13588);
nor U14750 (N_14750,N_13482,N_13935);
or U14751 (N_14751,N_13148,N_13101);
nand U14752 (N_14752,N_13624,N_13844);
nand U14753 (N_14753,N_13795,N_13062);
or U14754 (N_14754,N_13767,N_13246);
nand U14755 (N_14755,N_13523,N_13434);
nor U14756 (N_14756,N_13338,N_13905);
nand U14757 (N_14757,N_13338,N_13705);
nand U14758 (N_14758,N_13737,N_13665);
or U14759 (N_14759,N_13483,N_13604);
and U14760 (N_14760,N_13228,N_13435);
nand U14761 (N_14761,N_13101,N_13338);
nor U14762 (N_14762,N_13244,N_13922);
or U14763 (N_14763,N_13714,N_13065);
or U14764 (N_14764,N_13246,N_13248);
or U14765 (N_14765,N_13734,N_13818);
or U14766 (N_14766,N_13772,N_13793);
nand U14767 (N_14767,N_13305,N_13138);
or U14768 (N_14768,N_13517,N_13802);
and U14769 (N_14769,N_13049,N_13617);
nor U14770 (N_14770,N_13157,N_13161);
xor U14771 (N_14771,N_13708,N_13631);
or U14772 (N_14772,N_13166,N_13616);
and U14773 (N_14773,N_13280,N_13143);
nor U14774 (N_14774,N_13317,N_13801);
nor U14775 (N_14775,N_13542,N_13870);
or U14776 (N_14776,N_13577,N_13614);
and U14777 (N_14777,N_13405,N_13269);
or U14778 (N_14778,N_13414,N_13576);
nor U14779 (N_14779,N_13442,N_13139);
or U14780 (N_14780,N_13643,N_13516);
nor U14781 (N_14781,N_13932,N_13173);
xnor U14782 (N_14782,N_13019,N_13825);
xor U14783 (N_14783,N_13679,N_13805);
and U14784 (N_14784,N_13924,N_13147);
nor U14785 (N_14785,N_13024,N_13462);
nand U14786 (N_14786,N_13609,N_13733);
or U14787 (N_14787,N_13631,N_13608);
or U14788 (N_14788,N_13501,N_13375);
nor U14789 (N_14789,N_13173,N_13767);
nand U14790 (N_14790,N_13871,N_13867);
nor U14791 (N_14791,N_13272,N_13919);
nor U14792 (N_14792,N_13217,N_13092);
nor U14793 (N_14793,N_13964,N_13804);
and U14794 (N_14794,N_13193,N_13624);
and U14795 (N_14795,N_13456,N_13316);
nand U14796 (N_14796,N_13050,N_13098);
nor U14797 (N_14797,N_13006,N_13515);
nand U14798 (N_14798,N_13714,N_13567);
and U14799 (N_14799,N_13800,N_13540);
nand U14800 (N_14800,N_13750,N_13313);
or U14801 (N_14801,N_13620,N_13614);
nor U14802 (N_14802,N_13304,N_13944);
or U14803 (N_14803,N_13533,N_13943);
and U14804 (N_14804,N_13094,N_13620);
and U14805 (N_14805,N_13640,N_13567);
nor U14806 (N_14806,N_13703,N_13059);
and U14807 (N_14807,N_13073,N_13606);
and U14808 (N_14808,N_13040,N_13203);
nand U14809 (N_14809,N_13894,N_13178);
or U14810 (N_14810,N_13897,N_13327);
nor U14811 (N_14811,N_13443,N_13481);
nand U14812 (N_14812,N_13767,N_13204);
nor U14813 (N_14813,N_13974,N_13578);
nor U14814 (N_14814,N_13866,N_13827);
xnor U14815 (N_14815,N_13641,N_13694);
nand U14816 (N_14816,N_13912,N_13636);
xnor U14817 (N_14817,N_13213,N_13773);
nand U14818 (N_14818,N_13870,N_13710);
and U14819 (N_14819,N_13281,N_13011);
nor U14820 (N_14820,N_13640,N_13362);
nor U14821 (N_14821,N_13483,N_13185);
nor U14822 (N_14822,N_13031,N_13194);
or U14823 (N_14823,N_13157,N_13681);
and U14824 (N_14824,N_13392,N_13560);
and U14825 (N_14825,N_13560,N_13217);
or U14826 (N_14826,N_13735,N_13054);
nand U14827 (N_14827,N_13211,N_13542);
nand U14828 (N_14828,N_13053,N_13734);
xnor U14829 (N_14829,N_13271,N_13131);
and U14830 (N_14830,N_13572,N_13691);
xor U14831 (N_14831,N_13621,N_13149);
xor U14832 (N_14832,N_13546,N_13137);
xnor U14833 (N_14833,N_13323,N_13225);
xnor U14834 (N_14834,N_13518,N_13372);
and U14835 (N_14835,N_13915,N_13737);
nand U14836 (N_14836,N_13063,N_13591);
nand U14837 (N_14837,N_13068,N_13573);
and U14838 (N_14838,N_13734,N_13824);
nand U14839 (N_14839,N_13859,N_13780);
nand U14840 (N_14840,N_13463,N_13674);
xor U14841 (N_14841,N_13014,N_13648);
nor U14842 (N_14842,N_13082,N_13523);
nor U14843 (N_14843,N_13324,N_13367);
and U14844 (N_14844,N_13645,N_13493);
or U14845 (N_14845,N_13514,N_13808);
xor U14846 (N_14846,N_13296,N_13525);
nand U14847 (N_14847,N_13969,N_13882);
and U14848 (N_14848,N_13982,N_13698);
xor U14849 (N_14849,N_13553,N_13724);
xnor U14850 (N_14850,N_13858,N_13331);
nand U14851 (N_14851,N_13481,N_13145);
and U14852 (N_14852,N_13798,N_13591);
nor U14853 (N_14853,N_13764,N_13996);
and U14854 (N_14854,N_13498,N_13137);
nand U14855 (N_14855,N_13418,N_13355);
and U14856 (N_14856,N_13153,N_13744);
nor U14857 (N_14857,N_13745,N_13550);
and U14858 (N_14858,N_13316,N_13069);
nand U14859 (N_14859,N_13733,N_13337);
or U14860 (N_14860,N_13438,N_13166);
nor U14861 (N_14861,N_13061,N_13394);
nor U14862 (N_14862,N_13044,N_13742);
or U14863 (N_14863,N_13916,N_13341);
and U14864 (N_14864,N_13664,N_13200);
xor U14865 (N_14865,N_13744,N_13803);
nor U14866 (N_14866,N_13543,N_13672);
nand U14867 (N_14867,N_13630,N_13245);
nand U14868 (N_14868,N_13385,N_13574);
and U14869 (N_14869,N_13382,N_13098);
nand U14870 (N_14870,N_13295,N_13026);
or U14871 (N_14871,N_13470,N_13587);
and U14872 (N_14872,N_13996,N_13399);
and U14873 (N_14873,N_13669,N_13433);
and U14874 (N_14874,N_13282,N_13999);
xor U14875 (N_14875,N_13406,N_13451);
and U14876 (N_14876,N_13833,N_13720);
xnor U14877 (N_14877,N_13510,N_13101);
xor U14878 (N_14878,N_13298,N_13819);
or U14879 (N_14879,N_13958,N_13766);
xor U14880 (N_14880,N_13847,N_13893);
nor U14881 (N_14881,N_13397,N_13288);
nor U14882 (N_14882,N_13459,N_13830);
and U14883 (N_14883,N_13373,N_13871);
and U14884 (N_14884,N_13187,N_13920);
or U14885 (N_14885,N_13734,N_13857);
nor U14886 (N_14886,N_13225,N_13579);
xnor U14887 (N_14887,N_13487,N_13822);
nor U14888 (N_14888,N_13274,N_13200);
nand U14889 (N_14889,N_13158,N_13726);
nor U14890 (N_14890,N_13725,N_13122);
xor U14891 (N_14891,N_13160,N_13415);
and U14892 (N_14892,N_13216,N_13254);
xnor U14893 (N_14893,N_13848,N_13818);
xor U14894 (N_14894,N_13625,N_13767);
and U14895 (N_14895,N_13699,N_13072);
xnor U14896 (N_14896,N_13508,N_13403);
and U14897 (N_14897,N_13235,N_13822);
nor U14898 (N_14898,N_13972,N_13386);
xor U14899 (N_14899,N_13073,N_13040);
and U14900 (N_14900,N_13124,N_13643);
nand U14901 (N_14901,N_13726,N_13386);
and U14902 (N_14902,N_13010,N_13007);
and U14903 (N_14903,N_13946,N_13602);
or U14904 (N_14904,N_13905,N_13984);
xnor U14905 (N_14905,N_13252,N_13376);
and U14906 (N_14906,N_13284,N_13173);
nand U14907 (N_14907,N_13947,N_13796);
xor U14908 (N_14908,N_13910,N_13621);
xor U14909 (N_14909,N_13408,N_13168);
xnor U14910 (N_14910,N_13502,N_13877);
xnor U14911 (N_14911,N_13341,N_13377);
nand U14912 (N_14912,N_13878,N_13038);
nand U14913 (N_14913,N_13780,N_13144);
xor U14914 (N_14914,N_13604,N_13208);
xnor U14915 (N_14915,N_13877,N_13773);
nand U14916 (N_14916,N_13828,N_13448);
xor U14917 (N_14917,N_13748,N_13114);
nand U14918 (N_14918,N_13093,N_13280);
nor U14919 (N_14919,N_13694,N_13791);
xnor U14920 (N_14920,N_13887,N_13709);
or U14921 (N_14921,N_13387,N_13103);
or U14922 (N_14922,N_13407,N_13649);
or U14923 (N_14923,N_13613,N_13981);
and U14924 (N_14924,N_13028,N_13125);
nand U14925 (N_14925,N_13813,N_13243);
nor U14926 (N_14926,N_13044,N_13706);
nand U14927 (N_14927,N_13296,N_13826);
xnor U14928 (N_14928,N_13890,N_13423);
nand U14929 (N_14929,N_13574,N_13458);
or U14930 (N_14930,N_13688,N_13917);
xnor U14931 (N_14931,N_13204,N_13448);
nor U14932 (N_14932,N_13876,N_13996);
or U14933 (N_14933,N_13918,N_13066);
xor U14934 (N_14934,N_13192,N_13043);
and U14935 (N_14935,N_13728,N_13493);
or U14936 (N_14936,N_13857,N_13668);
and U14937 (N_14937,N_13409,N_13576);
nor U14938 (N_14938,N_13407,N_13876);
xnor U14939 (N_14939,N_13968,N_13193);
and U14940 (N_14940,N_13376,N_13221);
nand U14941 (N_14941,N_13944,N_13025);
nor U14942 (N_14942,N_13784,N_13614);
nand U14943 (N_14943,N_13621,N_13250);
or U14944 (N_14944,N_13459,N_13080);
nand U14945 (N_14945,N_13272,N_13960);
and U14946 (N_14946,N_13621,N_13459);
nand U14947 (N_14947,N_13130,N_13028);
nand U14948 (N_14948,N_13680,N_13528);
and U14949 (N_14949,N_13671,N_13811);
nand U14950 (N_14950,N_13310,N_13370);
nand U14951 (N_14951,N_13973,N_13919);
xor U14952 (N_14952,N_13583,N_13673);
xnor U14953 (N_14953,N_13384,N_13528);
nand U14954 (N_14954,N_13797,N_13672);
and U14955 (N_14955,N_13465,N_13505);
xnor U14956 (N_14956,N_13987,N_13481);
or U14957 (N_14957,N_13566,N_13519);
xnor U14958 (N_14958,N_13997,N_13028);
or U14959 (N_14959,N_13223,N_13450);
nor U14960 (N_14960,N_13637,N_13853);
nand U14961 (N_14961,N_13127,N_13618);
xnor U14962 (N_14962,N_13511,N_13931);
nor U14963 (N_14963,N_13452,N_13736);
nand U14964 (N_14964,N_13905,N_13928);
nor U14965 (N_14965,N_13672,N_13166);
nor U14966 (N_14966,N_13704,N_13494);
nor U14967 (N_14967,N_13218,N_13599);
xnor U14968 (N_14968,N_13989,N_13751);
nand U14969 (N_14969,N_13943,N_13332);
nor U14970 (N_14970,N_13974,N_13088);
nand U14971 (N_14971,N_13890,N_13275);
and U14972 (N_14972,N_13623,N_13486);
nor U14973 (N_14973,N_13428,N_13910);
xor U14974 (N_14974,N_13742,N_13683);
or U14975 (N_14975,N_13789,N_13971);
xor U14976 (N_14976,N_13706,N_13643);
xor U14977 (N_14977,N_13012,N_13260);
nor U14978 (N_14978,N_13537,N_13850);
xor U14979 (N_14979,N_13594,N_13832);
and U14980 (N_14980,N_13897,N_13445);
nor U14981 (N_14981,N_13653,N_13421);
nand U14982 (N_14982,N_13716,N_13330);
and U14983 (N_14983,N_13777,N_13823);
xor U14984 (N_14984,N_13699,N_13635);
nand U14985 (N_14985,N_13405,N_13948);
nand U14986 (N_14986,N_13604,N_13426);
xor U14987 (N_14987,N_13709,N_13361);
and U14988 (N_14988,N_13161,N_13212);
nor U14989 (N_14989,N_13141,N_13020);
nor U14990 (N_14990,N_13150,N_13404);
nor U14991 (N_14991,N_13001,N_13581);
nand U14992 (N_14992,N_13197,N_13297);
or U14993 (N_14993,N_13212,N_13330);
nor U14994 (N_14994,N_13751,N_13089);
or U14995 (N_14995,N_13207,N_13391);
xnor U14996 (N_14996,N_13926,N_13046);
xor U14997 (N_14997,N_13040,N_13272);
nand U14998 (N_14998,N_13470,N_13823);
nand U14999 (N_14999,N_13574,N_13654);
nor U15000 (N_15000,N_14631,N_14742);
nor U15001 (N_15001,N_14174,N_14836);
nor U15002 (N_15002,N_14261,N_14472);
and U15003 (N_15003,N_14210,N_14438);
nand U15004 (N_15004,N_14092,N_14659);
and U15005 (N_15005,N_14349,N_14905);
or U15006 (N_15006,N_14143,N_14051);
nand U15007 (N_15007,N_14373,N_14673);
nor U15008 (N_15008,N_14094,N_14990);
xor U15009 (N_15009,N_14778,N_14952);
xor U15010 (N_15010,N_14095,N_14079);
or U15011 (N_15011,N_14755,N_14813);
or U15012 (N_15012,N_14661,N_14628);
and U15013 (N_15013,N_14885,N_14965);
and U15014 (N_15014,N_14535,N_14356);
nor U15015 (N_15015,N_14933,N_14522);
or U15016 (N_15016,N_14328,N_14130);
xnor U15017 (N_15017,N_14000,N_14162);
nand U15018 (N_15018,N_14649,N_14001);
nor U15019 (N_15019,N_14276,N_14856);
nand U15020 (N_15020,N_14724,N_14519);
xor U15021 (N_15021,N_14539,N_14053);
xor U15022 (N_15022,N_14196,N_14288);
or U15023 (N_15023,N_14082,N_14037);
or U15024 (N_15024,N_14721,N_14940);
or U15025 (N_15025,N_14528,N_14131);
nand U15026 (N_15026,N_14573,N_14675);
and U15027 (N_15027,N_14518,N_14733);
xor U15028 (N_15028,N_14224,N_14616);
or U15029 (N_15029,N_14478,N_14071);
nand U15030 (N_15030,N_14794,N_14188);
and U15031 (N_15031,N_14284,N_14064);
and U15032 (N_15032,N_14756,N_14278);
and U15033 (N_15033,N_14789,N_14170);
nand U15034 (N_15034,N_14916,N_14760);
xor U15035 (N_15035,N_14708,N_14643);
nand U15036 (N_15036,N_14250,N_14561);
nor U15037 (N_15037,N_14049,N_14784);
nand U15038 (N_15038,N_14936,N_14425);
and U15039 (N_15039,N_14371,N_14372);
nor U15040 (N_15040,N_14879,N_14259);
and U15041 (N_15041,N_14927,N_14719);
nand U15042 (N_15042,N_14776,N_14321);
and U15043 (N_15043,N_14818,N_14011);
nand U15044 (N_15044,N_14791,N_14099);
nor U15045 (N_15045,N_14112,N_14903);
or U15046 (N_15046,N_14468,N_14597);
nor U15047 (N_15047,N_14388,N_14139);
xor U15048 (N_15048,N_14298,N_14422);
nand U15049 (N_15049,N_14848,N_14795);
nor U15050 (N_15050,N_14516,N_14601);
nand U15051 (N_15051,N_14446,N_14638);
and U15052 (N_15052,N_14774,N_14378);
nor U15053 (N_15053,N_14912,N_14462);
and U15054 (N_15054,N_14687,N_14979);
xnor U15055 (N_15055,N_14360,N_14351);
and U15056 (N_15056,N_14752,N_14065);
or U15057 (N_15057,N_14758,N_14456);
nor U15058 (N_15058,N_14431,N_14014);
or U15059 (N_15059,N_14269,N_14466);
nor U15060 (N_15060,N_14861,N_14796);
and U15061 (N_15061,N_14963,N_14052);
and U15062 (N_15062,N_14394,N_14692);
or U15063 (N_15063,N_14024,N_14364);
xnor U15064 (N_15064,N_14995,N_14206);
xnor U15065 (N_15065,N_14840,N_14013);
nand U15066 (N_15066,N_14954,N_14391);
nor U15067 (N_15067,N_14853,N_14017);
nor U15068 (N_15068,N_14006,N_14635);
xnor U15069 (N_15069,N_14902,N_14824);
xnor U15070 (N_15070,N_14549,N_14567);
xnor U15071 (N_15071,N_14487,N_14076);
nand U15072 (N_15072,N_14666,N_14312);
and U15073 (N_15073,N_14846,N_14681);
and U15074 (N_15074,N_14827,N_14622);
nand U15075 (N_15075,N_14226,N_14403);
xor U15076 (N_15076,N_14587,N_14350);
and U15077 (N_15077,N_14343,N_14073);
and U15078 (N_15078,N_14458,N_14173);
and U15079 (N_15079,N_14639,N_14480);
nor U15080 (N_15080,N_14797,N_14738);
or U15081 (N_15081,N_14720,N_14397);
xor U15082 (N_15082,N_14301,N_14385);
xor U15083 (N_15083,N_14189,N_14991);
nor U15084 (N_15084,N_14485,N_14685);
xor U15085 (N_15085,N_14010,N_14124);
and U15086 (N_15086,N_14823,N_14652);
nor U15087 (N_15087,N_14283,N_14999);
and U15088 (N_15088,N_14988,N_14566);
or U15089 (N_15089,N_14324,N_14946);
xor U15090 (N_15090,N_14727,N_14303);
nor U15091 (N_15091,N_14159,N_14163);
and U15092 (N_15092,N_14676,N_14955);
nor U15093 (N_15093,N_14662,N_14589);
nor U15094 (N_15094,N_14297,N_14571);
nor U15095 (N_15095,N_14435,N_14832);
nor U15096 (N_15096,N_14494,N_14200);
nor U15097 (N_15097,N_14503,N_14945);
xnor U15098 (N_15098,N_14078,N_14097);
nand U15099 (N_15099,N_14490,N_14187);
nand U15100 (N_15100,N_14627,N_14347);
and U15101 (N_15101,N_14938,N_14722);
nor U15102 (N_15102,N_14232,N_14004);
nand U15103 (N_15103,N_14619,N_14151);
nand U15104 (N_15104,N_14906,N_14207);
nor U15105 (N_15105,N_14266,N_14254);
or U15106 (N_15106,N_14514,N_14704);
and U15107 (N_15107,N_14591,N_14811);
and U15108 (N_15108,N_14670,N_14409);
and U15109 (N_15109,N_14067,N_14396);
nand U15110 (N_15110,N_14041,N_14858);
nor U15111 (N_15111,N_14251,N_14421);
or U15112 (N_15112,N_14033,N_14888);
and U15113 (N_15113,N_14181,N_14081);
nor U15114 (N_15114,N_14809,N_14960);
or U15115 (N_15115,N_14678,N_14376);
xor U15116 (N_15116,N_14291,N_14793);
or U15117 (N_15117,N_14723,N_14949);
xnor U15118 (N_15118,N_14197,N_14896);
nand U15119 (N_15119,N_14969,N_14660);
xnor U15120 (N_15120,N_14294,N_14444);
and U15121 (N_15121,N_14241,N_14536);
nor U15122 (N_15122,N_14602,N_14633);
and U15123 (N_15123,N_14498,N_14021);
or U15124 (N_15124,N_14019,N_14304);
xor U15125 (N_15125,N_14452,N_14154);
or U15126 (N_15126,N_14728,N_14679);
and U15127 (N_15127,N_14016,N_14672);
or U15128 (N_15128,N_14667,N_14871);
nor U15129 (N_15129,N_14557,N_14594);
or U15130 (N_15130,N_14816,N_14997);
nor U15131 (N_15131,N_14677,N_14632);
nor U15132 (N_15132,N_14127,N_14100);
and U15133 (N_15133,N_14798,N_14491);
nand U15134 (N_15134,N_14517,N_14167);
nand U15135 (N_15135,N_14015,N_14607);
nor U15136 (N_15136,N_14803,N_14160);
xor U15137 (N_15137,N_14346,N_14499);
nand U15138 (N_15138,N_14157,N_14085);
or U15139 (N_15139,N_14511,N_14406);
xor U15140 (N_15140,N_14886,N_14866);
nand U15141 (N_15141,N_14384,N_14031);
and U15142 (N_15142,N_14552,N_14904);
or U15143 (N_15143,N_14176,N_14715);
xor U15144 (N_15144,N_14762,N_14548);
and U15145 (N_15145,N_14982,N_14883);
or U15146 (N_15146,N_14482,N_14749);
nand U15147 (N_15147,N_14357,N_14786);
and U15148 (N_15148,N_14111,N_14495);
xor U15149 (N_15149,N_14575,N_14265);
or U15150 (N_15150,N_14621,N_14348);
nand U15151 (N_15151,N_14048,N_14640);
nand U15152 (N_15152,N_14747,N_14586);
and U15153 (N_15153,N_14763,N_14086);
nor U15154 (N_15154,N_14529,N_14464);
or U15155 (N_15155,N_14802,N_14822);
or U15156 (N_15156,N_14964,N_14109);
nand U15157 (N_15157,N_14600,N_14253);
and U15158 (N_15158,N_14113,N_14493);
nor U15159 (N_15159,N_14231,N_14668);
nand U15160 (N_15160,N_14674,N_14923);
xnor U15161 (N_15161,N_14381,N_14941);
or U15162 (N_15162,N_14230,N_14996);
nor U15163 (N_15163,N_14759,N_14702);
and U15164 (N_15164,N_14551,N_14931);
or U15165 (N_15165,N_14576,N_14863);
or U15166 (N_15166,N_14026,N_14433);
or U15167 (N_15167,N_14027,N_14974);
or U15168 (N_15168,N_14987,N_14893);
and U15169 (N_15169,N_14243,N_14882);
nor U15170 (N_15170,N_14264,N_14689);
nor U15171 (N_15171,N_14018,N_14958);
nand U15172 (N_15172,N_14273,N_14046);
or U15173 (N_15173,N_14985,N_14845);
and U15174 (N_15174,N_14107,N_14544);
nand U15175 (N_15175,N_14408,N_14302);
and U15176 (N_15176,N_14116,N_14664);
or U15177 (N_15177,N_14465,N_14655);
or U15178 (N_15178,N_14367,N_14411);
nand U15179 (N_15179,N_14970,N_14383);
nand U15180 (N_15180,N_14305,N_14977);
or U15181 (N_15181,N_14153,N_14042);
nand U15182 (N_15182,N_14476,N_14834);
and U15183 (N_15183,N_14496,N_14398);
nor U15184 (N_15184,N_14208,N_14029);
nor U15185 (N_15185,N_14541,N_14775);
nand U15186 (N_15186,N_14935,N_14634);
xnor U15187 (N_15187,N_14274,N_14686);
nand U15188 (N_15188,N_14355,N_14325);
or U15189 (N_15189,N_14684,N_14369);
nor U15190 (N_15190,N_14864,N_14165);
nand U15191 (N_15191,N_14943,N_14047);
nand U15192 (N_15192,N_14924,N_14754);
xor U15193 (N_15193,N_14175,N_14336);
and U15194 (N_15194,N_14532,N_14387);
or U15195 (N_15195,N_14467,N_14331);
and U15196 (N_15196,N_14564,N_14258);
or U15197 (N_15197,N_14530,N_14642);
nor U15198 (N_15198,N_14698,N_14335);
or U15199 (N_15199,N_14671,N_14220);
nor U15200 (N_15200,N_14101,N_14972);
and U15201 (N_15201,N_14077,N_14645);
and U15202 (N_15202,N_14128,N_14966);
xnor U15203 (N_15203,N_14821,N_14202);
and U15204 (N_15204,N_14296,N_14432);
or U15205 (N_15205,N_14582,N_14569);
and U15206 (N_15206,N_14929,N_14777);
xnor U15207 (N_15207,N_14850,N_14365);
nor U15208 (N_15208,N_14537,N_14429);
and U15209 (N_15209,N_14590,N_14788);
and U15210 (N_15210,N_14473,N_14779);
and U15211 (N_15211,N_14819,N_14044);
or U15212 (N_15212,N_14504,N_14469);
nor U15213 (N_15213,N_14901,N_14837);
and U15214 (N_15214,N_14152,N_14734);
or U15215 (N_15215,N_14028,N_14359);
nor U15216 (N_15216,N_14857,N_14599);
nand U15217 (N_15217,N_14193,N_14579);
and U15218 (N_15218,N_14108,N_14038);
nand U15219 (N_15219,N_14096,N_14262);
nand U15220 (N_15220,N_14229,N_14329);
nand U15221 (N_15221,N_14417,N_14300);
nand U15222 (N_15222,N_14217,N_14072);
and U15223 (N_15223,N_14790,N_14177);
nand U15224 (N_15224,N_14316,N_14695);
xor U15225 (N_15225,N_14869,N_14158);
and U15226 (N_15226,N_14980,N_14757);
and U15227 (N_15227,N_14959,N_14275);
xor U15228 (N_15228,N_14618,N_14523);
xor U15229 (N_15229,N_14457,N_14764);
nand U15230 (N_15230,N_14613,N_14463);
xor U15231 (N_15231,N_14451,N_14867);
or U15232 (N_15232,N_14138,N_14132);
nor U15233 (N_15233,N_14327,N_14322);
xnor U15234 (N_15234,N_14088,N_14709);
and U15235 (N_15235,N_14743,N_14110);
nand U15236 (N_15236,N_14669,N_14654);
or U15237 (N_15237,N_14263,N_14502);
nand U15238 (N_15238,N_14105,N_14962);
nor U15239 (N_15239,N_14688,N_14693);
and U15240 (N_15240,N_14479,N_14892);
nor U15241 (N_15241,N_14257,N_14948);
xor U15242 (N_15242,N_14787,N_14937);
or U15243 (N_15243,N_14002,N_14062);
and U15244 (N_15244,N_14334,N_14104);
or U15245 (N_15245,N_14595,N_14184);
and U15246 (N_15246,N_14833,N_14855);
nand U15247 (N_15247,N_14615,N_14910);
nand U15248 (N_15248,N_14534,N_14550);
or U15249 (N_15249,N_14983,N_14792);
and U15250 (N_15250,N_14236,N_14123);
or U15251 (N_15251,N_14238,N_14087);
and U15252 (N_15252,N_14282,N_14286);
or U15253 (N_15253,N_14172,N_14363);
xnor U15254 (N_15254,N_14887,N_14326);
or U15255 (N_15255,N_14609,N_14290);
xor U15256 (N_15256,N_14390,N_14563);
or U15257 (N_15257,N_14361,N_14075);
xor U15258 (N_15258,N_14647,N_14370);
or U15259 (N_15259,N_14829,N_14293);
and U15260 (N_15260,N_14022,N_14070);
and U15261 (N_15261,N_14917,N_14828);
xnor U15262 (N_15262,N_14588,N_14691);
xor U15263 (N_15263,N_14145,N_14900);
nor U15264 (N_15264,N_14657,N_14930);
xor U15265 (N_15265,N_14374,N_14084);
nor U15266 (N_15266,N_14225,N_14714);
nand U15267 (N_15267,N_14129,N_14911);
xor U15268 (N_15268,N_14093,N_14428);
nor U15269 (N_15269,N_14651,N_14209);
and U15270 (N_15270,N_14656,N_14748);
nand U15271 (N_15271,N_14553,N_14546);
or U15272 (N_15272,N_14309,N_14913);
and U15273 (N_15273,N_14507,N_14993);
xnor U15274 (N_15274,N_14404,N_14914);
or U15275 (N_15275,N_14820,N_14603);
and U15276 (N_15276,N_14799,N_14289);
nor U15277 (N_15277,N_14596,N_14287);
or U15278 (N_15278,N_14877,N_14746);
xnor U15279 (N_15279,N_14148,N_14583);
nand U15280 (N_15280,N_14817,N_14835);
nand U15281 (N_15281,N_14868,N_14558);
or U15282 (N_15282,N_14069,N_14825);
nand U15283 (N_15283,N_14121,N_14474);
and U15284 (N_15284,N_14570,N_14399);
xor U15285 (N_15285,N_14847,N_14992);
and U15286 (N_15286,N_14068,N_14611);
and U15287 (N_15287,N_14909,N_14280);
nand U15288 (N_15288,N_14513,N_14898);
and U15289 (N_15289,N_14285,N_14292);
nor U15290 (N_15290,N_14354,N_14453);
and U15291 (N_15291,N_14765,N_14353);
nand U15292 (N_15292,N_14120,N_14716);
nand U15293 (N_15293,N_14707,N_14448);
nor U15294 (N_15294,N_14339,N_14612);
nor U15295 (N_15295,N_14826,N_14577);
nand U15296 (N_15296,N_14234,N_14862);
or U15297 (N_15297,N_14899,N_14838);
and U15298 (N_15298,N_14460,N_14711);
nand U15299 (N_15299,N_14227,N_14771);
or U15300 (N_15300,N_14808,N_14233);
nor U15301 (N_15301,N_14279,N_14731);
and U15302 (N_15302,N_14574,N_14418);
or U15303 (N_15303,N_14035,N_14812);
nand U15304 (N_15304,N_14956,N_14135);
and U15305 (N_15305,N_14277,N_14683);
and U15306 (N_15306,N_14423,N_14450);
and U15307 (N_15307,N_14098,N_14445);
or U15308 (N_15308,N_14141,N_14424);
and U15309 (N_15309,N_14800,N_14481);
nor U15310 (N_15310,N_14769,N_14091);
or U15311 (N_15311,N_14598,N_14745);
or U15312 (N_15312,N_14056,N_14003);
and U15313 (N_15313,N_14501,N_14020);
xor U15314 (N_15314,N_14981,N_14461);
xnor U15315 (N_15315,N_14247,N_14410);
or U15316 (N_15316,N_14168,N_14830);
or U15317 (N_15317,N_14256,N_14245);
or U15318 (N_15318,N_14620,N_14951);
nor U15319 (N_15319,N_14984,N_14801);
nor U15320 (N_15320,N_14106,N_14524);
nand U15321 (N_15321,N_14295,N_14308);
and U15322 (N_15322,N_14040,N_14565);
or U15323 (N_15323,N_14054,N_14060);
nor U15324 (N_15324,N_14039,N_14012);
and U15325 (N_15325,N_14216,N_14059);
or U15326 (N_15326,N_14271,N_14190);
nand U15327 (N_15327,N_14646,N_14630);
nor U15328 (N_15328,N_14314,N_14058);
nor U15329 (N_15329,N_14785,N_14415);
nor U15330 (N_15330,N_14147,N_14007);
and U15331 (N_15331,N_14712,N_14194);
or U15332 (N_15332,N_14875,N_14696);
or U15333 (N_15333,N_14894,N_14119);
or U15334 (N_15334,N_14851,N_14810);
xnor U15335 (N_15335,N_14500,N_14865);
or U15336 (N_15336,N_14736,N_14890);
and U15337 (N_15337,N_14344,N_14509);
nand U15338 (N_15338,N_14136,N_14045);
or U15339 (N_15339,N_14626,N_14585);
or U15340 (N_15340,N_14515,N_14961);
or U15341 (N_15341,N_14780,N_14986);
or U15342 (N_15342,N_14260,N_14400);
and U15343 (N_15343,N_14114,N_14214);
nor U15344 (N_15344,N_14741,N_14430);
xor U15345 (N_15345,N_14213,N_14606);
nor U15346 (N_15346,N_14806,N_14538);
xor U15347 (N_15347,N_14436,N_14614);
and U15348 (N_15348,N_14455,N_14957);
nor U15349 (N_15349,N_14608,N_14183);
nor U15350 (N_15350,N_14126,N_14486);
or U15351 (N_15351,N_14807,N_14204);
xor U15352 (N_15352,N_14268,N_14252);
and U15353 (N_15353,N_14919,N_14117);
or U15354 (N_15354,N_14080,N_14392);
and U15355 (N_15355,N_14781,N_14380);
xnor U15356 (N_15356,N_14375,N_14454);
and U15357 (N_15357,N_14362,N_14248);
nor U15358 (N_15358,N_14842,N_14717);
or U15359 (N_15359,N_14860,N_14699);
xor U15360 (N_15360,N_14744,N_14125);
nand U15361 (N_15361,N_14377,N_14648);
nand U15362 (N_15362,N_14533,N_14783);
xor U15363 (N_15363,N_14706,N_14506);
nor U15364 (N_15364,N_14680,N_14944);
and U15365 (N_15365,N_14407,N_14306);
nand U15366 (N_15366,N_14973,N_14934);
or U15367 (N_15367,N_14313,N_14215);
and U15368 (N_15368,N_14761,N_14235);
or U15369 (N_15369,N_14249,N_14008);
nand U15370 (N_15370,N_14443,N_14531);
and U15371 (N_15371,N_14427,N_14604);
xor U15372 (N_15372,N_14508,N_14891);
and U15373 (N_15373,N_14337,N_14636);
nand U15374 (N_15374,N_14118,N_14488);
and U15375 (N_15375,N_14697,N_14218);
and U15376 (N_15376,N_14897,N_14185);
or U15377 (N_15377,N_14426,N_14700);
or U15378 (N_15378,N_14804,N_14239);
xnor U15379 (N_15379,N_14317,N_14179);
and U15380 (N_15380,N_14849,N_14839);
or U15381 (N_15381,N_14971,N_14873);
nand U15382 (N_15382,N_14772,N_14342);
and U15383 (N_15383,N_14525,N_14144);
and U15384 (N_15384,N_14246,N_14171);
nor U15385 (N_15385,N_14156,N_14178);
nand U15386 (N_15386,N_14405,N_14512);
and U15387 (N_15387,N_14942,N_14057);
nor U15388 (N_15388,N_14023,N_14844);
and U15389 (N_15389,N_14718,N_14950);
nand U15390 (N_15390,N_14061,N_14470);
xor U15391 (N_15391,N_14975,N_14554);
or U15392 (N_15392,N_14782,N_14483);
xor U15393 (N_15393,N_14926,N_14730);
xnor U15394 (N_15394,N_14526,N_14939);
xnor U15395 (N_15395,N_14032,N_14694);
nand U15396 (N_15396,N_14442,N_14663);
or U15397 (N_15397,N_14164,N_14166);
nand U15398 (N_15398,N_14617,N_14439);
nor U15399 (N_15399,N_14644,N_14315);
xnor U15400 (N_15400,N_14102,N_14884);
nor U15401 (N_15401,N_14034,N_14416);
nor U15402 (N_15402,N_14547,N_14332);
xnor U15403 (N_15403,N_14637,N_14750);
or U15404 (N_15404,N_14272,N_14814);
and U15405 (N_15405,N_14815,N_14043);
nor U15406 (N_15406,N_14201,N_14767);
and U15407 (N_15407,N_14191,N_14228);
and U15408 (N_15408,N_14489,N_14368);
nand U15409 (N_15409,N_14701,N_14690);
nand U15410 (N_15410,N_14475,N_14149);
nor U15411 (N_15411,N_14922,N_14729);
nand U15412 (N_15412,N_14089,N_14976);
or U15413 (N_15413,N_14198,N_14221);
xor U15414 (N_15414,N_14137,N_14319);
or U15415 (N_15415,N_14841,N_14063);
nor U15416 (N_15416,N_14318,N_14036);
xor U15417 (N_15417,N_14270,N_14330);
nand U15418 (N_15418,N_14307,N_14255);
and U15419 (N_15419,N_14310,N_14665);
nor U15420 (N_15420,N_14843,N_14967);
or U15421 (N_15421,N_14419,N_14859);
or U15422 (N_15422,N_14978,N_14623);
nand U15423 (N_15423,N_14641,N_14593);
xor U15424 (N_15424,N_14740,N_14420);
nor U15425 (N_15425,N_14895,N_14401);
or U15426 (N_15426,N_14437,N_14341);
nand U15427 (N_15427,N_14323,N_14918);
xnor U15428 (N_15428,N_14751,N_14393);
and U15429 (N_15429,N_14055,N_14908);
and U15430 (N_15430,N_14989,N_14831);
or U15431 (N_15431,N_14212,N_14520);
and U15432 (N_15432,N_14345,N_14920);
or U15433 (N_15433,N_14876,N_14653);
and U15434 (N_15434,N_14770,N_14074);
or U15435 (N_15435,N_14223,N_14878);
and U15436 (N_15436,N_14705,N_14650);
and U15437 (N_15437,N_14471,N_14682);
xnor U15438 (N_15438,N_14872,N_14542);
nand U15439 (N_15439,N_14915,N_14998);
xnor U15440 (N_15440,N_14203,N_14497);
xnor U15441 (N_15441,N_14340,N_14555);
xnor U15442 (N_15442,N_14492,N_14739);
nor U15443 (N_15443,N_14805,N_14560);
nor U15444 (N_15444,N_14186,N_14115);
nor U15445 (N_15445,N_14580,N_14880);
or U15446 (N_15446,N_14870,N_14240);
nand U15447 (N_15447,N_14180,N_14169);
or U15448 (N_15448,N_14389,N_14103);
nor U15449 (N_15449,N_14994,N_14009);
or U15450 (N_15450,N_14205,N_14725);
xor U15451 (N_15451,N_14311,N_14703);
nand U15452 (N_15452,N_14559,N_14932);
xor U15453 (N_15453,N_14737,N_14625);
or U15454 (N_15454,N_14928,N_14182);
and U15455 (N_15455,N_14556,N_14581);
xor U15456 (N_15456,N_14584,N_14766);
nand U15457 (N_15457,N_14192,N_14545);
xor U15458 (N_15458,N_14505,N_14134);
or U15459 (N_15459,N_14414,N_14881);
nor U15460 (N_15460,N_14658,N_14366);
xor U15461 (N_15461,N_14773,N_14459);
nand U15462 (N_15462,N_14219,N_14768);
nand U15463 (N_15463,N_14449,N_14925);
nand U15464 (N_15464,N_14568,N_14338);
and U15465 (N_15465,N_14624,N_14379);
xor U15466 (N_15466,N_14484,N_14953);
and U15467 (N_15467,N_14382,N_14358);
and U15468 (N_15468,N_14402,N_14199);
nand U15469 (N_15469,N_14267,N_14050);
nand U15470 (N_15470,N_14090,N_14713);
nor U15471 (N_15471,N_14440,N_14510);
nor U15472 (N_15472,N_14578,N_14907);
nor U15473 (N_15473,N_14543,N_14710);
nand U15474 (N_15474,N_14413,N_14195);
and U15475 (N_15475,N_14150,N_14889);
or U15476 (N_15476,N_14244,N_14562);
xnor U15477 (N_15477,N_14083,N_14237);
and U15478 (N_15478,N_14155,N_14726);
nand U15479 (N_15479,N_14447,N_14605);
or U15480 (N_15480,N_14921,N_14477);
xnor U15481 (N_15481,N_14947,N_14299);
xor U15482 (N_15482,N_14592,N_14854);
nand U15483 (N_15483,N_14527,N_14753);
nand U15484 (N_15484,N_14386,N_14441);
or U15485 (N_15485,N_14540,N_14610);
nand U15486 (N_15486,N_14320,N_14434);
nand U15487 (N_15487,N_14133,N_14030);
nor U15488 (N_15488,N_14521,N_14281);
nand U15489 (N_15489,N_14629,N_14852);
nand U15490 (N_15490,N_14968,N_14352);
xnor U15491 (N_15491,N_14142,N_14211);
xor U15492 (N_15492,N_14066,N_14161);
nor U15493 (N_15493,N_14333,N_14395);
nor U15494 (N_15494,N_14735,N_14025);
and U15495 (N_15495,N_14140,N_14222);
xnor U15496 (N_15496,N_14412,N_14242);
or U15497 (N_15497,N_14572,N_14005);
xor U15498 (N_15498,N_14874,N_14732);
nor U15499 (N_15499,N_14122,N_14146);
xnor U15500 (N_15500,N_14527,N_14479);
nor U15501 (N_15501,N_14929,N_14727);
nor U15502 (N_15502,N_14323,N_14671);
nand U15503 (N_15503,N_14171,N_14976);
nand U15504 (N_15504,N_14556,N_14725);
xnor U15505 (N_15505,N_14019,N_14623);
and U15506 (N_15506,N_14373,N_14496);
and U15507 (N_15507,N_14975,N_14055);
nand U15508 (N_15508,N_14610,N_14510);
xnor U15509 (N_15509,N_14271,N_14362);
xnor U15510 (N_15510,N_14604,N_14994);
or U15511 (N_15511,N_14505,N_14003);
xnor U15512 (N_15512,N_14593,N_14723);
xor U15513 (N_15513,N_14243,N_14199);
nand U15514 (N_15514,N_14943,N_14860);
nand U15515 (N_15515,N_14798,N_14450);
nor U15516 (N_15516,N_14914,N_14320);
and U15517 (N_15517,N_14852,N_14872);
or U15518 (N_15518,N_14661,N_14152);
nor U15519 (N_15519,N_14730,N_14419);
and U15520 (N_15520,N_14563,N_14654);
or U15521 (N_15521,N_14594,N_14567);
and U15522 (N_15522,N_14209,N_14073);
and U15523 (N_15523,N_14347,N_14426);
and U15524 (N_15524,N_14885,N_14070);
nand U15525 (N_15525,N_14977,N_14444);
nor U15526 (N_15526,N_14910,N_14841);
nand U15527 (N_15527,N_14178,N_14353);
and U15528 (N_15528,N_14342,N_14850);
nand U15529 (N_15529,N_14660,N_14747);
xor U15530 (N_15530,N_14191,N_14975);
nor U15531 (N_15531,N_14884,N_14038);
xnor U15532 (N_15532,N_14156,N_14051);
nor U15533 (N_15533,N_14788,N_14975);
nor U15534 (N_15534,N_14665,N_14028);
xor U15535 (N_15535,N_14501,N_14844);
or U15536 (N_15536,N_14078,N_14974);
and U15537 (N_15537,N_14424,N_14364);
and U15538 (N_15538,N_14474,N_14337);
nor U15539 (N_15539,N_14123,N_14537);
and U15540 (N_15540,N_14619,N_14371);
xnor U15541 (N_15541,N_14170,N_14646);
nor U15542 (N_15542,N_14196,N_14738);
or U15543 (N_15543,N_14260,N_14213);
and U15544 (N_15544,N_14517,N_14479);
nor U15545 (N_15545,N_14865,N_14481);
nand U15546 (N_15546,N_14921,N_14530);
and U15547 (N_15547,N_14248,N_14025);
xor U15548 (N_15548,N_14371,N_14082);
and U15549 (N_15549,N_14904,N_14348);
or U15550 (N_15550,N_14154,N_14035);
and U15551 (N_15551,N_14147,N_14653);
nand U15552 (N_15552,N_14915,N_14997);
xor U15553 (N_15553,N_14782,N_14499);
nor U15554 (N_15554,N_14270,N_14387);
nor U15555 (N_15555,N_14829,N_14497);
nand U15556 (N_15556,N_14529,N_14641);
or U15557 (N_15557,N_14940,N_14288);
and U15558 (N_15558,N_14893,N_14394);
nor U15559 (N_15559,N_14701,N_14597);
or U15560 (N_15560,N_14447,N_14346);
nand U15561 (N_15561,N_14441,N_14240);
nor U15562 (N_15562,N_14426,N_14045);
nor U15563 (N_15563,N_14774,N_14370);
and U15564 (N_15564,N_14202,N_14295);
nor U15565 (N_15565,N_14996,N_14666);
and U15566 (N_15566,N_14584,N_14153);
or U15567 (N_15567,N_14040,N_14017);
xor U15568 (N_15568,N_14866,N_14682);
nand U15569 (N_15569,N_14748,N_14158);
or U15570 (N_15570,N_14154,N_14992);
nand U15571 (N_15571,N_14265,N_14475);
xor U15572 (N_15572,N_14634,N_14992);
xnor U15573 (N_15573,N_14194,N_14146);
nor U15574 (N_15574,N_14572,N_14409);
and U15575 (N_15575,N_14291,N_14036);
and U15576 (N_15576,N_14718,N_14120);
and U15577 (N_15577,N_14482,N_14823);
nand U15578 (N_15578,N_14379,N_14946);
or U15579 (N_15579,N_14403,N_14689);
and U15580 (N_15580,N_14563,N_14231);
nor U15581 (N_15581,N_14925,N_14528);
xor U15582 (N_15582,N_14791,N_14695);
nor U15583 (N_15583,N_14384,N_14480);
or U15584 (N_15584,N_14336,N_14779);
and U15585 (N_15585,N_14713,N_14610);
xor U15586 (N_15586,N_14239,N_14846);
nor U15587 (N_15587,N_14951,N_14405);
xnor U15588 (N_15588,N_14385,N_14858);
or U15589 (N_15589,N_14754,N_14084);
xnor U15590 (N_15590,N_14192,N_14594);
xnor U15591 (N_15591,N_14355,N_14247);
and U15592 (N_15592,N_14726,N_14412);
xor U15593 (N_15593,N_14201,N_14274);
nand U15594 (N_15594,N_14159,N_14737);
and U15595 (N_15595,N_14678,N_14091);
or U15596 (N_15596,N_14494,N_14298);
and U15597 (N_15597,N_14723,N_14916);
or U15598 (N_15598,N_14245,N_14697);
nor U15599 (N_15599,N_14827,N_14214);
xnor U15600 (N_15600,N_14899,N_14023);
nor U15601 (N_15601,N_14628,N_14046);
xnor U15602 (N_15602,N_14740,N_14037);
nor U15603 (N_15603,N_14567,N_14463);
nand U15604 (N_15604,N_14263,N_14324);
xor U15605 (N_15605,N_14599,N_14720);
and U15606 (N_15606,N_14473,N_14554);
and U15607 (N_15607,N_14089,N_14538);
nand U15608 (N_15608,N_14874,N_14616);
nand U15609 (N_15609,N_14333,N_14203);
and U15610 (N_15610,N_14472,N_14645);
and U15611 (N_15611,N_14574,N_14117);
and U15612 (N_15612,N_14914,N_14471);
or U15613 (N_15613,N_14429,N_14115);
or U15614 (N_15614,N_14025,N_14693);
nand U15615 (N_15615,N_14515,N_14308);
nor U15616 (N_15616,N_14977,N_14954);
nand U15617 (N_15617,N_14247,N_14902);
xnor U15618 (N_15618,N_14929,N_14691);
and U15619 (N_15619,N_14145,N_14092);
or U15620 (N_15620,N_14651,N_14155);
nor U15621 (N_15621,N_14310,N_14113);
or U15622 (N_15622,N_14770,N_14107);
nand U15623 (N_15623,N_14173,N_14291);
and U15624 (N_15624,N_14375,N_14715);
nor U15625 (N_15625,N_14002,N_14042);
nor U15626 (N_15626,N_14779,N_14521);
nor U15627 (N_15627,N_14982,N_14938);
and U15628 (N_15628,N_14472,N_14108);
xnor U15629 (N_15629,N_14099,N_14596);
nand U15630 (N_15630,N_14756,N_14764);
nand U15631 (N_15631,N_14877,N_14834);
xnor U15632 (N_15632,N_14473,N_14243);
nor U15633 (N_15633,N_14910,N_14493);
or U15634 (N_15634,N_14503,N_14478);
and U15635 (N_15635,N_14292,N_14499);
or U15636 (N_15636,N_14137,N_14974);
xor U15637 (N_15637,N_14110,N_14064);
nand U15638 (N_15638,N_14497,N_14333);
and U15639 (N_15639,N_14378,N_14376);
nand U15640 (N_15640,N_14090,N_14037);
xor U15641 (N_15641,N_14101,N_14445);
xor U15642 (N_15642,N_14057,N_14913);
nand U15643 (N_15643,N_14456,N_14385);
and U15644 (N_15644,N_14862,N_14388);
nand U15645 (N_15645,N_14270,N_14099);
xnor U15646 (N_15646,N_14191,N_14557);
nand U15647 (N_15647,N_14440,N_14923);
nor U15648 (N_15648,N_14727,N_14576);
or U15649 (N_15649,N_14649,N_14330);
nand U15650 (N_15650,N_14269,N_14868);
xnor U15651 (N_15651,N_14977,N_14708);
or U15652 (N_15652,N_14260,N_14548);
nand U15653 (N_15653,N_14431,N_14408);
nor U15654 (N_15654,N_14220,N_14791);
nand U15655 (N_15655,N_14538,N_14303);
nand U15656 (N_15656,N_14035,N_14712);
xnor U15657 (N_15657,N_14657,N_14177);
nor U15658 (N_15658,N_14083,N_14510);
xnor U15659 (N_15659,N_14669,N_14221);
and U15660 (N_15660,N_14418,N_14800);
xor U15661 (N_15661,N_14831,N_14982);
and U15662 (N_15662,N_14027,N_14142);
xor U15663 (N_15663,N_14319,N_14191);
or U15664 (N_15664,N_14917,N_14699);
xor U15665 (N_15665,N_14273,N_14845);
xor U15666 (N_15666,N_14113,N_14919);
or U15667 (N_15667,N_14489,N_14137);
and U15668 (N_15668,N_14708,N_14978);
xnor U15669 (N_15669,N_14435,N_14284);
xor U15670 (N_15670,N_14472,N_14128);
or U15671 (N_15671,N_14485,N_14138);
nand U15672 (N_15672,N_14640,N_14489);
xor U15673 (N_15673,N_14710,N_14465);
nand U15674 (N_15674,N_14372,N_14163);
xor U15675 (N_15675,N_14400,N_14664);
or U15676 (N_15676,N_14046,N_14131);
or U15677 (N_15677,N_14405,N_14309);
xor U15678 (N_15678,N_14144,N_14919);
xnor U15679 (N_15679,N_14865,N_14101);
nor U15680 (N_15680,N_14737,N_14121);
nand U15681 (N_15681,N_14969,N_14233);
or U15682 (N_15682,N_14401,N_14385);
and U15683 (N_15683,N_14204,N_14707);
xnor U15684 (N_15684,N_14392,N_14094);
nand U15685 (N_15685,N_14903,N_14972);
nand U15686 (N_15686,N_14235,N_14587);
or U15687 (N_15687,N_14391,N_14339);
nor U15688 (N_15688,N_14783,N_14666);
nand U15689 (N_15689,N_14941,N_14212);
nand U15690 (N_15690,N_14464,N_14840);
nand U15691 (N_15691,N_14989,N_14819);
or U15692 (N_15692,N_14273,N_14259);
nor U15693 (N_15693,N_14268,N_14829);
or U15694 (N_15694,N_14866,N_14089);
nand U15695 (N_15695,N_14726,N_14309);
or U15696 (N_15696,N_14299,N_14713);
and U15697 (N_15697,N_14483,N_14647);
and U15698 (N_15698,N_14950,N_14128);
or U15699 (N_15699,N_14822,N_14383);
nor U15700 (N_15700,N_14045,N_14252);
nor U15701 (N_15701,N_14026,N_14322);
and U15702 (N_15702,N_14442,N_14771);
nand U15703 (N_15703,N_14789,N_14346);
nand U15704 (N_15704,N_14823,N_14832);
nand U15705 (N_15705,N_14700,N_14901);
nand U15706 (N_15706,N_14719,N_14202);
and U15707 (N_15707,N_14060,N_14946);
and U15708 (N_15708,N_14834,N_14452);
nand U15709 (N_15709,N_14971,N_14481);
nor U15710 (N_15710,N_14052,N_14587);
and U15711 (N_15711,N_14437,N_14636);
or U15712 (N_15712,N_14831,N_14496);
nor U15713 (N_15713,N_14212,N_14194);
nor U15714 (N_15714,N_14863,N_14145);
xor U15715 (N_15715,N_14485,N_14797);
or U15716 (N_15716,N_14091,N_14713);
nand U15717 (N_15717,N_14003,N_14404);
nand U15718 (N_15718,N_14109,N_14737);
nand U15719 (N_15719,N_14404,N_14919);
nor U15720 (N_15720,N_14735,N_14601);
nor U15721 (N_15721,N_14130,N_14402);
nand U15722 (N_15722,N_14739,N_14793);
and U15723 (N_15723,N_14655,N_14466);
and U15724 (N_15724,N_14989,N_14601);
nand U15725 (N_15725,N_14467,N_14359);
or U15726 (N_15726,N_14472,N_14501);
or U15727 (N_15727,N_14504,N_14779);
or U15728 (N_15728,N_14363,N_14271);
and U15729 (N_15729,N_14803,N_14017);
nor U15730 (N_15730,N_14784,N_14510);
nand U15731 (N_15731,N_14174,N_14926);
xor U15732 (N_15732,N_14487,N_14868);
nor U15733 (N_15733,N_14392,N_14835);
or U15734 (N_15734,N_14803,N_14701);
and U15735 (N_15735,N_14968,N_14955);
xnor U15736 (N_15736,N_14697,N_14451);
nand U15737 (N_15737,N_14196,N_14320);
xnor U15738 (N_15738,N_14603,N_14295);
and U15739 (N_15739,N_14073,N_14425);
or U15740 (N_15740,N_14297,N_14230);
xor U15741 (N_15741,N_14318,N_14460);
and U15742 (N_15742,N_14889,N_14003);
xor U15743 (N_15743,N_14809,N_14708);
nor U15744 (N_15744,N_14176,N_14961);
and U15745 (N_15745,N_14411,N_14738);
or U15746 (N_15746,N_14554,N_14991);
and U15747 (N_15747,N_14134,N_14630);
or U15748 (N_15748,N_14081,N_14339);
or U15749 (N_15749,N_14457,N_14383);
nor U15750 (N_15750,N_14740,N_14441);
nand U15751 (N_15751,N_14214,N_14602);
and U15752 (N_15752,N_14466,N_14180);
or U15753 (N_15753,N_14187,N_14532);
and U15754 (N_15754,N_14375,N_14467);
nor U15755 (N_15755,N_14332,N_14578);
nor U15756 (N_15756,N_14805,N_14400);
or U15757 (N_15757,N_14177,N_14069);
or U15758 (N_15758,N_14377,N_14812);
or U15759 (N_15759,N_14972,N_14631);
nor U15760 (N_15760,N_14130,N_14832);
xor U15761 (N_15761,N_14871,N_14311);
nor U15762 (N_15762,N_14029,N_14940);
nand U15763 (N_15763,N_14134,N_14104);
or U15764 (N_15764,N_14393,N_14146);
or U15765 (N_15765,N_14215,N_14344);
nor U15766 (N_15766,N_14128,N_14199);
or U15767 (N_15767,N_14377,N_14393);
and U15768 (N_15768,N_14012,N_14602);
nand U15769 (N_15769,N_14622,N_14591);
and U15770 (N_15770,N_14674,N_14704);
or U15771 (N_15771,N_14603,N_14565);
or U15772 (N_15772,N_14272,N_14471);
nor U15773 (N_15773,N_14115,N_14314);
nor U15774 (N_15774,N_14557,N_14444);
or U15775 (N_15775,N_14227,N_14554);
or U15776 (N_15776,N_14011,N_14821);
or U15777 (N_15777,N_14766,N_14778);
and U15778 (N_15778,N_14622,N_14000);
xnor U15779 (N_15779,N_14346,N_14215);
nand U15780 (N_15780,N_14869,N_14421);
and U15781 (N_15781,N_14176,N_14051);
and U15782 (N_15782,N_14362,N_14914);
and U15783 (N_15783,N_14038,N_14851);
or U15784 (N_15784,N_14944,N_14939);
nor U15785 (N_15785,N_14633,N_14711);
or U15786 (N_15786,N_14899,N_14258);
nor U15787 (N_15787,N_14114,N_14383);
and U15788 (N_15788,N_14506,N_14827);
or U15789 (N_15789,N_14369,N_14349);
nand U15790 (N_15790,N_14200,N_14340);
nand U15791 (N_15791,N_14207,N_14883);
and U15792 (N_15792,N_14190,N_14030);
or U15793 (N_15793,N_14672,N_14080);
and U15794 (N_15794,N_14668,N_14634);
nand U15795 (N_15795,N_14792,N_14979);
nor U15796 (N_15796,N_14447,N_14966);
xnor U15797 (N_15797,N_14513,N_14720);
xnor U15798 (N_15798,N_14983,N_14558);
and U15799 (N_15799,N_14444,N_14140);
or U15800 (N_15800,N_14751,N_14863);
or U15801 (N_15801,N_14284,N_14552);
and U15802 (N_15802,N_14108,N_14670);
xnor U15803 (N_15803,N_14803,N_14774);
nor U15804 (N_15804,N_14485,N_14171);
and U15805 (N_15805,N_14010,N_14759);
and U15806 (N_15806,N_14669,N_14409);
and U15807 (N_15807,N_14890,N_14943);
nand U15808 (N_15808,N_14253,N_14266);
xnor U15809 (N_15809,N_14840,N_14540);
or U15810 (N_15810,N_14305,N_14056);
nand U15811 (N_15811,N_14690,N_14284);
nand U15812 (N_15812,N_14058,N_14261);
nor U15813 (N_15813,N_14467,N_14300);
or U15814 (N_15814,N_14902,N_14509);
and U15815 (N_15815,N_14385,N_14053);
nor U15816 (N_15816,N_14494,N_14299);
or U15817 (N_15817,N_14690,N_14614);
nor U15818 (N_15818,N_14505,N_14535);
and U15819 (N_15819,N_14335,N_14230);
xnor U15820 (N_15820,N_14406,N_14686);
nand U15821 (N_15821,N_14675,N_14083);
nor U15822 (N_15822,N_14000,N_14104);
xor U15823 (N_15823,N_14524,N_14503);
nor U15824 (N_15824,N_14517,N_14031);
xnor U15825 (N_15825,N_14485,N_14764);
nand U15826 (N_15826,N_14115,N_14368);
and U15827 (N_15827,N_14462,N_14405);
nand U15828 (N_15828,N_14721,N_14060);
nor U15829 (N_15829,N_14711,N_14662);
or U15830 (N_15830,N_14407,N_14408);
and U15831 (N_15831,N_14085,N_14514);
nand U15832 (N_15832,N_14529,N_14916);
nand U15833 (N_15833,N_14895,N_14803);
nor U15834 (N_15834,N_14843,N_14412);
and U15835 (N_15835,N_14922,N_14616);
xnor U15836 (N_15836,N_14168,N_14245);
xor U15837 (N_15837,N_14620,N_14832);
and U15838 (N_15838,N_14570,N_14501);
nor U15839 (N_15839,N_14869,N_14986);
and U15840 (N_15840,N_14990,N_14013);
and U15841 (N_15841,N_14396,N_14506);
nor U15842 (N_15842,N_14112,N_14235);
nand U15843 (N_15843,N_14917,N_14435);
nand U15844 (N_15844,N_14448,N_14502);
or U15845 (N_15845,N_14430,N_14472);
or U15846 (N_15846,N_14264,N_14746);
nor U15847 (N_15847,N_14662,N_14970);
and U15848 (N_15848,N_14222,N_14560);
or U15849 (N_15849,N_14590,N_14396);
nand U15850 (N_15850,N_14048,N_14343);
nor U15851 (N_15851,N_14517,N_14805);
nor U15852 (N_15852,N_14012,N_14199);
or U15853 (N_15853,N_14103,N_14789);
nand U15854 (N_15854,N_14939,N_14672);
and U15855 (N_15855,N_14010,N_14739);
nand U15856 (N_15856,N_14545,N_14087);
nor U15857 (N_15857,N_14754,N_14621);
and U15858 (N_15858,N_14841,N_14967);
nand U15859 (N_15859,N_14934,N_14637);
xor U15860 (N_15860,N_14557,N_14232);
or U15861 (N_15861,N_14620,N_14616);
or U15862 (N_15862,N_14574,N_14672);
and U15863 (N_15863,N_14473,N_14557);
nand U15864 (N_15864,N_14624,N_14363);
nand U15865 (N_15865,N_14304,N_14969);
xnor U15866 (N_15866,N_14319,N_14688);
nor U15867 (N_15867,N_14441,N_14582);
and U15868 (N_15868,N_14268,N_14349);
nor U15869 (N_15869,N_14843,N_14704);
xor U15870 (N_15870,N_14433,N_14993);
and U15871 (N_15871,N_14614,N_14251);
and U15872 (N_15872,N_14130,N_14013);
nor U15873 (N_15873,N_14877,N_14664);
or U15874 (N_15874,N_14313,N_14823);
nor U15875 (N_15875,N_14628,N_14451);
xor U15876 (N_15876,N_14018,N_14641);
xor U15877 (N_15877,N_14153,N_14409);
nand U15878 (N_15878,N_14973,N_14048);
or U15879 (N_15879,N_14889,N_14287);
xnor U15880 (N_15880,N_14088,N_14003);
nor U15881 (N_15881,N_14322,N_14470);
and U15882 (N_15882,N_14243,N_14032);
xor U15883 (N_15883,N_14506,N_14877);
xor U15884 (N_15884,N_14243,N_14011);
and U15885 (N_15885,N_14003,N_14139);
nor U15886 (N_15886,N_14111,N_14584);
nor U15887 (N_15887,N_14339,N_14976);
or U15888 (N_15888,N_14019,N_14175);
nand U15889 (N_15889,N_14980,N_14840);
nor U15890 (N_15890,N_14376,N_14732);
xnor U15891 (N_15891,N_14694,N_14046);
xnor U15892 (N_15892,N_14477,N_14453);
nor U15893 (N_15893,N_14227,N_14739);
or U15894 (N_15894,N_14092,N_14835);
nor U15895 (N_15895,N_14731,N_14213);
xnor U15896 (N_15896,N_14354,N_14381);
and U15897 (N_15897,N_14704,N_14474);
xor U15898 (N_15898,N_14618,N_14640);
and U15899 (N_15899,N_14186,N_14331);
xnor U15900 (N_15900,N_14874,N_14543);
or U15901 (N_15901,N_14974,N_14594);
and U15902 (N_15902,N_14481,N_14052);
and U15903 (N_15903,N_14202,N_14333);
xor U15904 (N_15904,N_14817,N_14603);
nand U15905 (N_15905,N_14783,N_14376);
or U15906 (N_15906,N_14238,N_14346);
nor U15907 (N_15907,N_14799,N_14428);
xnor U15908 (N_15908,N_14181,N_14372);
nand U15909 (N_15909,N_14546,N_14720);
xor U15910 (N_15910,N_14191,N_14001);
nor U15911 (N_15911,N_14397,N_14363);
nor U15912 (N_15912,N_14760,N_14002);
nor U15913 (N_15913,N_14547,N_14885);
and U15914 (N_15914,N_14701,N_14717);
or U15915 (N_15915,N_14220,N_14862);
nor U15916 (N_15916,N_14191,N_14938);
nor U15917 (N_15917,N_14027,N_14099);
and U15918 (N_15918,N_14725,N_14242);
nand U15919 (N_15919,N_14704,N_14373);
and U15920 (N_15920,N_14290,N_14553);
xor U15921 (N_15921,N_14169,N_14835);
nor U15922 (N_15922,N_14503,N_14359);
and U15923 (N_15923,N_14034,N_14861);
nor U15924 (N_15924,N_14870,N_14339);
nand U15925 (N_15925,N_14350,N_14483);
nand U15926 (N_15926,N_14746,N_14841);
nand U15927 (N_15927,N_14821,N_14003);
or U15928 (N_15928,N_14406,N_14278);
nand U15929 (N_15929,N_14540,N_14206);
and U15930 (N_15930,N_14397,N_14104);
nor U15931 (N_15931,N_14533,N_14522);
and U15932 (N_15932,N_14617,N_14192);
nor U15933 (N_15933,N_14221,N_14929);
nand U15934 (N_15934,N_14255,N_14696);
or U15935 (N_15935,N_14764,N_14777);
xor U15936 (N_15936,N_14916,N_14670);
or U15937 (N_15937,N_14378,N_14762);
xor U15938 (N_15938,N_14481,N_14492);
nand U15939 (N_15939,N_14915,N_14042);
xor U15940 (N_15940,N_14084,N_14443);
or U15941 (N_15941,N_14865,N_14062);
and U15942 (N_15942,N_14020,N_14347);
and U15943 (N_15943,N_14100,N_14606);
xnor U15944 (N_15944,N_14085,N_14614);
xnor U15945 (N_15945,N_14170,N_14261);
and U15946 (N_15946,N_14375,N_14427);
or U15947 (N_15947,N_14263,N_14384);
xor U15948 (N_15948,N_14324,N_14693);
xor U15949 (N_15949,N_14561,N_14088);
xnor U15950 (N_15950,N_14867,N_14808);
and U15951 (N_15951,N_14960,N_14856);
or U15952 (N_15952,N_14788,N_14477);
xor U15953 (N_15953,N_14512,N_14742);
xnor U15954 (N_15954,N_14366,N_14306);
or U15955 (N_15955,N_14481,N_14868);
and U15956 (N_15956,N_14102,N_14470);
xnor U15957 (N_15957,N_14873,N_14471);
or U15958 (N_15958,N_14146,N_14574);
nor U15959 (N_15959,N_14219,N_14359);
or U15960 (N_15960,N_14990,N_14895);
nand U15961 (N_15961,N_14009,N_14894);
xnor U15962 (N_15962,N_14797,N_14026);
nor U15963 (N_15963,N_14992,N_14109);
and U15964 (N_15964,N_14072,N_14794);
or U15965 (N_15965,N_14193,N_14638);
or U15966 (N_15966,N_14825,N_14703);
or U15967 (N_15967,N_14274,N_14909);
xnor U15968 (N_15968,N_14276,N_14176);
and U15969 (N_15969,N_14257,N_14330);
nand U15970 (N_15970,N_14156,N_14033);
or U15971 (N_15971,N_14137,N_14523);
nand U15972 (N_15972,N_14895,N_14874);
nor U15973 (N_15973,N_14474,N_14297);
nor U15974 (N_15974,N_14516,N_14277);
and U15975 (N_15975,N_14380,N_14589);
xnor U15976 (N_15976,N_14478,N_14727);
and U15977 (N_15977,N_14356,N_14501);
nand U15978 (N_15978,N_14395,N_14135);
nor U15979 (N_15979,N_14842,N_14261);
and U15980 (N_15980,N_14690,N_14080);
xor U15981 (N_15981,N_14983,N_14267);
or U15982 (N_15982,N_14618,N_14338);
nand U15983 (N_15983,N_14770,N_14577);
nor U15984 (N_15984,N_14909,N_14397);
nand U15985 (N_15985,N_14212,N_14546);
and U15986 (N_15986,N_14401,N_14296);
nand U15987 (N_15987,N_14435,N_14371);
nor U15988 (N_15988,N_14616,N_14044);
or U15989 (N_15989,N_14534,N_14377);
and U15990 (N_15990,N_14367,N_14001);
nand U15991 (N_15991,N_14284,N_14574);
and U15992 (N_15992,N_14601,N_14689);
nand U15993 (N_15993,N_14434,N_14670);
nor U15994 (N_15994,N_14002,N_14281);
xor U15995 (N_15995,N_14852,N_14876);
xor U15996 (N_15996,N_14176,N_14865);
nor U15997 (N_15997,N_14391,N_14472);
xnor U15998 (N_15998,N_14807,N_14780);
xnor U15999 (N_15999,N_14048,N_14784);
nor U16000 (N_16000,N_15856,N_15333);
nor U16001 (N_16001,N_15782,N_15969);
nand U16002 (N_16002,N_15269,N_15009);
nand U16003 (N_16003,N_15613,N_15200);
nor U16004 (N_16004,N_15444,N_15805);
and U16005 (N_16005,N_15278,N_15676);
and U16006 (N_16006,N_15165,N_15799);
or U16007 (N_16007,N_15489,N_15937);
and U16008 (N_16008,N_15452,N_15152);
nor U16009 (N_16009,N_15946,N_15218);
or U16010 (N_16010,N_15540,N_15596);
or U16011 (N_16011,N_15216,N_15705);
nand U16012 (N_16012,N_15783,N_15350);
xnor U16013 (N_16013,N_15589,N_15629);
or U16014 (N_16014,N_15945,N_15881);
xor U16015 (N_16015,N_15495,N_15276);
and U16016 (N_16016,N_15742,N_15592);
or U16017 (N_16017,N_15459,N_15259);
and U16018 (N_16018,N_15307,N_15264);
or U16019 (N_16019,N_15911,N_15939);
and U16020 (N_16020,N_15361,N_15751);
xnor U16021 (N_16021,N_15882,N_15857);
nor U16022 (N_16022,N_15367,N_15222);
and U16023 (N_16023,N_15324,N_15951);
nor U16024 (N_16024,N_15295,N_15957);
nor U16025 (N_16025,N_15959,N_15153);
xor U16026 (N_16026,N_15767,N_15312);
and U16027 (N_16027,N_15518,N_15718);
nor U16028 (N_16028,N_15373,N_15673);
xnor U16029 (N_16029,N_15864,N_15173);
nor U16030 (N_16030,N_15344,N_15995);
or U16031 (N_16031,N_15168,N_15570);
and U16032 (N_16032,N_15482,N_15615);
and U16033 (N_16033,N_15042,N_15651);
nand U16034 (N_16034,N_15710,N_15377);
xor U16035 (N_16035,N_15897,N_15722);
nor U16036 (N_16036,N_15178,N_15720);
or U16037 (N_16037,N_15028,N_15401);
nand U16038 (N_16038,N_15733,N_15352);
nor U16039 (N_16039,N_15019,N_15744);
nor U16040 (N_16040,N_15950,N_15662);
nor U16041 (N_16041,N_15023,N_15885);
or U16042 (N_16042,N_15268,N_15300);
or U16043 (N_16043,N_15156,N_15895);
and U16044 (N_16044,N_15031,N_15790);
nor U16045 (N_16045,N_15977,N_15090);
nand U16046 (N_16046,N_15699,N_15020);
nor U16047 (N_16047,N_15354,N_15494);
nand U16048 (N_16048,N_15996,N_15119);
or U16049 (N_16049,N_15768,N_15924);
and U16050 (N_16050,N_15228,N_15618);
nor U16051 (N_16051,N_15891,N_15774);
and U16052 (N_16052,N_15828,N_15778);
and U16053 (N_16053,N_15785,N_15519);
or U16054 (N_16054,N_15807,N_15320);
or U16055 (N_16055,N_15385,N_15638);
nand U16056 (N_16056,N_15772,N_15780);
xor U16057 (N_16057,N_15998,N_15148);
nand U16058 (N_16058,N_15674,N_15823);
nor U16059 (N_16059,N_15628,N_15552);
or U16060 (N_16060,N_15314,N_15713);
xor U16061 (N_16061,N_15260,N_15183);
nand U16062 (N_16062,N_15441,N_15964);
nand U16063 (N_16063,N_15787,N_15773);
xnor U16064 (N_16064,N_15563,N_15625);
and U16065 (N_16065,N_15703,N_15928);
xor U16066 (N_16066,N_15319,N_15079);
nand U16067 (N_16067,N_15983,N_15282);
nand U16068 (N_16068,N_15830,N_15867);
nand U16069 (N_16069,N_15397,N_15739);
nand U16070 (N_16070,N_15726,N_15762);
nor U16071 (N_16071,N_15682,N_15191);
xor U16072 (N_16072,N_15932,N_15217);
xor U16073 (N_16073,N_15449,N_15186);
or U16074 (N_16074,N_15632,N_15698);
or U16075 (N_16075,N_15484,N_15973);
nand U16076 (N_16076,N_15701,N_15914);
or U16077 (N_16077,N_15415,N_15815);
nand U16078 (N_16078,N_15360,N_15275);
or U16079 (N_16079,N_15004,N_15039);
and U16080 (N_16080,N_15128,N_15547);
nor U16081 (N_16081,N_15340,N_15729);
and U16082 (N_16082,N_15188,N_15109);
nor U16083 (N_16083,N_15985,N_15080);
nor U16084 (N_16084,N_15305,N_15487);
xnor U16085 (N_16085,N_15796,N_15808);
and U16086 (N_16086,N_15992,N_15043);
nor U16087 (N_16087,N_15606,N_15302);
xor U16088 (N_16088,N_15229,N_15378);
nand U16089 (N_16089,N_15577,N_15212);
and U16090 (N_16090,N_15686,N_15126);
xnor U16091 (N_16091,N_15149,N_15303);
nand U16092 (N_16092,N_15110,N_15163);
nor U16093 (N_16093,N_15952,N_15409);
nand U16094 (N_16094,N_15477,N_15053);
xnor U16095 (N_16095,N_15461,N_15037);
or U16096 (N_16096,N_15918,N_15193);
nor U16097 (N_16097,N_15752,N_15100);
and U16098 (N_16098,N_15383,N_15021);
xnor U16099 (N_16099,N_15266,N_15876);
xor U16100 (N_16100,N_15763,N_15531);
and U16101 (N_16101,N_15557,N_15386);
nor U16102 (N_16102,N_15586,N_15058);
or U16103 (N_16103,N_15051,N_15408);
nand U16104 (N_16104,N_15491,N_15761);
nand U16105 (N_16105,N_15697,N_15886);
nand U16106 (N_16106,N_15201,N_15658);
xor U16107 (N_16107,N_15463,N_15961);
or U16108 (N_16108,N_15930,N_15137);
and U16109 (N_16109,N_15167,N_15829);
nor U16110 (N_16110,N_15299,N_15421);
or U16111 (N_16111,N_15479,N_15061);
and U16112 (N_16112,N_15716,N_15448);
nand U16113 (N_16113,N_15908,N_15439);
and U16114 (N_16114,N_15108,N_15369);
nor U16115 (N_16115,N_15555,N_15187);
nand U16116 (N_16116,N_15712,N_15453);
xnor U16117 (N_16117,N_15363,N_15791);
xnor U16118 (N_16118,N_15388,N_15970);
nor U16119 (N_16119,N_15888,N_15656);
and U16120 (N_16120,N_15211,N_15226);
xor U16121 (N_16121,N_15664,N_15696);
and U16122 (N_16122,N_15633,N_15814);
and U16123 (N_16123,N_15113,N_15162);
xnor U16124 (N_16124,N_15347,N_15542);
nand U16125 (N_16125,N_15237,N_15393);
nand U16126 (N_16126,N_15953,N_15827);
nand U16127 (N_16127,N_15887,N_15512);
nand U16128 (N_16128,N_15581,N_15590);
nand U16129 (N_16129,N_15223,N_15166);
nand U16130 (N_16130,N_15313,N_15835);
nor U16131 (N_16131,N_15256,N_15436);
or U16132 (N_16132,N_15685,N_15261);
and U16133 (N_16133,N_15455,N_15084);
and U16134 (N_16134,N_15670,N_15405);
xnor U16135 (N_16135,N_15483,N_15943);
and U16136 (N_16136,N_15342,N_15708);
or U16137 (N_16137,N_15464,N_15690);
nand U16138 (N_16138,N_15598,N_15280);
nand U16139 (N_16139,N_15277,N_15567);
and U16140 (N_16140,N_15136,N_15879);
nand U16141 (N_16141,N_15068,N_15225);
xor U16142 (N_16142,N_15896,N_15248);
or U16143 (N_16143,N_15515,N_15721);
nand U16144 (N_16144,N_15125,N_15094);
xnor U16145 (N_16145,N_15734,N_15454);
xnor U16146 (N_16146,N_15677,N_15991);
nand U16147 (N_16147,N_15873,N_15883);
xor U16148 (N_16148,N_15473,N_15714);
or U16149 (N_16149,N_15366,N_15003);
nor U16150 (N_16150,N_15420,N_15472);
xnor U16151 (N_16151,N_15346,N_15660);
xor U16152 (N_16152,N_15258,N_15535);
xnor U16153 (N_16153,N_15919,N_15204);
xor U16154 (N_16154,N_15528,N_15921);
nor U16155 (N_16155,N_15654,N_15077);
nor U16156 (N_16156,N_15445,N_15396);
nor U16157 (N_16157,N_15859,N_15101);
nand U16158 (N_16158,N_15643,N_15612);
or U16159 (N_16159,N_15521,N_15982);
nand U16160 (N_16160,N_15574,N_15076);
nor U16161 (N_16161,N_15853,N_15786);
and U16162 (N_16162,N_15206,N_15600);
or U16163 (N_16163,N_15154,N_15368);
xor U16164 (N_16164,N_15728,N_15182);
and U16165 (N_16165,N_15012,N_15760);
and U16166 (N_16166,N_15064,N_15757);
and U16167 (N_16167,N_15349,N_15532);
or U16168 (N_16168,N_15511,N_15289);
nor U16169 (N_16169,N_15948,N_15017);
nor U16170 (N_16170,N_15678,N_15839);
nor U16171 (N_16171,N_15146,N_15000);
and U16172 (N_16172,N_15120,N_15184);
nand U16173 (N_16173,N_15245,N_15550);
or U16174 (N_16174,N_15435,N_15817);
or U16175 (N_16175,N_15706,N_15724);
nor U16176 (N_16176,N_15123,N_15838);
nand U16177 (N_16177,N_15675,N_15679);
xnor U16178 (N_16178,N_15416,N_15232);
and U16179 (N_16179,N_15040,N_15174);
xor U16180 (N_16180,N_15339,N_15680);
and U16181 (N_16181,N_15938,N_15322);
or U16182 (N_16182,N_15516,N_15608);
xnor U16183 (N_16183,N_15129,N_15981);
or U16184 (N_16184,N_15980,N_15711);
or U16185 (N_16185,N_15603,N_15164);
nor U16186 (N_16186,N_15024,N_15356);
nand U16187 (N_16187,N_15854,N_15103);
nand U16188 (N_16188,N_15907,N_15649);
nor U16189 (N_16189,N_15593,N_15317);
and U16190 (N_16190,N_15104,N_15587);
nor U16191 (N_16191,N_15849,N_15741);
nand U16192 (N_16192,N_15655,N_15890);
xor U16193 (N_16193,N_15358,N_15374);
or U16194 (N_16194,N_15826,N_15781);
or U16195 (N_16195,N_15355,N_15580);
and U16196 (N_16196,N_15311,N_15536);
xor U16197 (N_16197,N_15426,N_15884);
nand U16198 (N_16198,N_15509,N_15803);
or U16199 (N_16199,N_15816,N_15442);
and U16200 (N_16200,N_15810,N_15855);
xnor U16201 (N_16201,N_15318,N_15548);
xor U16202 (N_16202,N_15749,N_15387);
xor U16203 (N_16203,N_15062,N_15576);
nand U16204 (N_16204,N_15530,N_15868);
and U16205 (N_16205,N_15236,N_15789);
nor U16206 (N_16206,N_15290,N_15195);
or U16207 (N_16207,N_15496,N_15267);
nor U16208 (N_16208,N_15912,N_15138);
or U16209 (N_16209,N_15418,N_15870);
xor U16210 (N_16210,N_15372,N_15234);
nor U16211 (N_16211,N_15848,N_15041);
and U16212 (N_16212,N_15990,N_15106);
or U16213 (N_16213,N_15811,N_15272);
and U16214 (N_16214,N_15994,N_15913);
nand U16215 (N_16215,N_15866,N_15537);
and U16216 (N_16216,N_15797,N_15145);
or U16217 (N_16217,N_15327,N_15978);
and U16218 (N_16218,N_15582,N_15779);
or U16219 (N_16219,N_15055,N_15700);
or U16220 (N_16220,N_15784,N_15291);
or U16221 (N_16221,N_15652,N_15429);
nand U16222 (N_16222,N_15860,N_15018);
xor U16223 (N_16223,N_15695,N_15813);
nand U16224 (N_16224,N_15247,N_15428);
xnor U16225 (N_16225,N_15645,N_15499);
and U16226 (N_16226,N_15958,N_15309);
nor U16227 (N_16227,N_15093,N_15620);
and U16228 (N_16228,N_15871,N_15433);
and U16229 (N_16229,N_15792,N_15765);
nand U16230 (N_16230,N_15279,N_15920);
nor U16231 (N_16231,N_15427,N_15623);
and U16232 (N_16232,N_15395,N_15007);
xnor U16233 (N_16233,N_15931,N_15975);
xnor U16234 (N_16234,N_15553,N_15476);
nor U16235 (N_16235,N_15458,N_15666);
nand U16236 (N_16236,N_15124,N_15610);
nor U16237 (N_16237,N_15379,N_15987);
xnor U16238 (N_16238,N_15692,N_15524);
or U16239 (N_16239,N_15648,N_15157);
xor U16240 (N_16240,N_15822,N_15392);
xor U16241 (N_16241,N_15889,N_15262);
nand U16242 (N_16242,N_15529,N_15723);
nor U16243 (N_16243,N_15402,N_15766);
nor U16244 (N_16244,N_15155,N_15844);
or U16245 (N_16245,N_15497,N_15292);
nand U16246 (N_16246,N_15467,N_15617);
xor U16247 (N_16247,N_15667,N_15335);
or U16248 (N_16248,N_15926,N_15231);
nor U16249 (N_16249,N_15597,N_15503);
nor U16250 (N_16250,N_15066,N_15099);
and U16251 (N_16251,N_15240,N_15894);
nor U16252 (N_16252,N_15558,N_15900);
and U16253 (N_16253,N_15254,N_15862);
nor U16254 (N_16254,N_15451,N_15381);
xnor U16255 (N_16255,N_15665,N_15604);
or U16256 (N_16256,N_15285,N_15414);
and U16257 (N_16257,N_15045,N_15955);
and U16258 (N_16258,N_15422,N_15177);
xor U16259 (N_16259,N_15922,N_15502);
and U16260 (N_16260,N_15539,N_15127);
xnor U16261 (N_16261,N_15036,N_15565);
xor U16262 (N_16262,N_15821,N_15989);
and U16263 (N_16263,N_15874,N_15669);
nand U16264 (N_16264,N_15475,N_15044);
xnor U16265 (N_16265,N_15083,N_15820);
nor U16266 (N_16266,N_15709,N_15770);
or U16267 (N_16267,N_15091,N_15514);
nand U16268 (N_16268,N_15286,N_15326);
nor U16269 (N_16269,N_15480,N_15022);
nor U16270 (N_16270,N_15988,N_15646);
nor U16271 (N_16271,N_15263,N_15909);
or U16272 (N_16272,N_15960,N_15601);
and U16273 (N_16273,N_15176,N_15046);
and U16274 (N_16274,N_15025,N_15121);
nand U16275 (N_16275,N_15910,N_15825);
and U16276 (N_16276,N_15147,N_15543);
xor U16277 (N_16277,N_15224,N_15923);
nand U16278 (N_16278,N_15450,N_15198);
xnor U16279 (N_16279,N_15583,N_15430);
or U16280 (N_16280,N_15172,N_15134);
or U16281 (N_16281,N_15438,N_15556);
or U16282 (N_16282,N_15190,N_15230);
and U16283 (N_16283,N_15798,N_15845);
nor U16284 (N_16284,N_15836,N_15659);
xnor U16285 (N_16285,N_15050,N_15671);
nand U16286 (N_16286,N_15490,N_15424);
xnor U16287 (N_16287,N_15351,N_15199);
nor U16288 (N_16288,N_15566,N_15133);
nor U16289 (N_16289,N_15621,N_15688);
nand U16290 (N_16290,N_15965,N_15049);
or U16291 (N_16291,N_15437,N_15933);
nand U16292 (N_16292,N_15026,N_15691);
and U16293 (N_16293,N_15082,N_15488);
and U16294 (N_16294,N_15942,N_15595);
and U16295 (N_16295,N_15070,N_15241);
nand U16296 (N_16296,N_15689,N_15971);
nor U16297 (N_16297,N_15384,N_15010);
or U16298 (N_16298,N_15641,N_15534);
nand U16299 (N_16299,N_15525,N_15607);
and U16300 (N_16300,N_15298,N_15533);
or U16301 (N_16301,N_15239,N_15214);
or U16302 (N_16302,N_15905,N_15086);
and U16303 (N_16303,N_15215,N_15657);
or U16304 (N_16304,N_15257,N_15034);
nand U16305 (N_16305,N_15391,N_15081);
or U16306 (N_16306,N_15337,N_15668);
nand U16307 (N_16307,N_15578,N_15892);
nor U16308 (N_16308,N_15635,N_15095);
xor U16309 (N_16309,N_15376,N_15842);
nor U16310 (N_16310,N_15717,N_15325);
and U16311 (N_16311,N_15114,N_15793);
nand U16312 (N_16312,N_15935,N_15976);
nand U16313 (N_16313,N_15619,N_15863);
or U16314 (N_16314,N_15501,N_15411);
xnor U16315 (N_16315,N_15069,N_15902);
xor U16316 (N_16316,N_15343,N_15795);
xnor U16317 (N_16317,N_15903,N_15456);
nand U16318 (N_16318,N_15348,N_15967);
nor U16319 (N_16319,N_15161,N_15181);
and U16320 (N_16320,N_15747,N_15560);
nand U16321 (N_16321,N_15468,N_15060);
nand U16322 (N_16322,N_15627,N_15549);
and U16323 (N_16323,N_15308,N_15750);
nor U16324 (N_16324,N_15471,N_15545);
nor U16325 (N_16325,N_15107,N_15624);
and U16326 (N_16326,N_15085,N_15251);
or U16327 (N_16327,N_15088,N_15893);
and U16328 (N_16328,N_15192,N_15802);
nand U16329 (N_16329,N_15571,N_15554);
xor U16330 (N_16330,N_15636,N_15956);
or U16331 (N_16331,N_15252,N_15375);
xor U16332 (N_16332,N_15404,N_15640);
nor U16333 (N_16333,N_15731,N_15197);
xor U16334 (N_16334,N_15869,N_15273);
and U16335 (N_16335,N_15008,N_15014);
and U16336 (N_16336,N_15599,N_15440);
nand U16337 (N_16337,N_15297,N_15141);
xor U16338 (N_16338,N_15283,N_15131);
and U16339 (N_16339,N_15917,N_15653);
nand U16340 (N_16340,N_15073,N_15833);
and U16341 (N_16341,N_15160,N_15075);
or U16342 (N_16342,N_15227,N_15929);
or U16343 (N_16343,N_15746,N_15562);
nor U16344 (N_16344,N_15219,N_15837);
and U16345 (N_16345,N_15611,N_15171);
nor U16346 (N_16346,N_15336,N_15067);
xnor U16347 (N_16347,N_15622,N_15736);
nand U16348 (N_16348,N_15389,N_15210);
nand U16349 (N_16349,N_15238,N_15831);
nand U16350 (N_16350,N_15614,N_15647);
nor U16351 (N_16351,N_15399,N_15116);
xor U16352 (N_16352,N_15737,N_15875);
nor U16353 (N_16353,N_15898,N_15777);
and U16354 (N_16354,N_15927,N_15105);
and U16355 (N_16355,N_15293,N_15115);
nor U16356 (N_16356,N_15840,N_15602);
xnor U16357 (N_16357,N_15208,N_15800);
nor U16358 (N_16358,N_15804,N_15097);
nand U16359 (N_16359,N_15253,N_15071);
xnor U16360 (N_16360,N_15730,N_15288);
xnor U16361 (N_16361,N_15812,N_15052);
xnor U16362 (N_16362,N_15801,N_15609);
and U16363 (N_16363,N_15818,N_15915);
or U16364 (N_16364,N_15693,N_15203);
or U16365 (N_16365,N_15189,N_15330);
nand U16366 (N_16366,N_15423,N_15754);
nor U16367 (N_16367,N_15304,N_15447);
nor U16368 (N_16368,N_15359,N_15522);
nand U16369 (N_16369,N_15513,N_15568);
or U16370 (N_16370,N_15999,N_15132);
xnor U16371 (N_16371,N_15353,N_15013);
xor U16372 (N_16372,N_15794,N_15296);
or U16373 (N_16373,N_15112,N_15498);
nand U16374 (N_16374,N_15431,N_15150);
xnor U16375 (N_16375,N_15029,N_15748);
nand U16376 (N_16376,N_15087,N_15630);
nand U16377 (N_16377,N_15650,N_15281);
or U16378 (N_16378,N_15158,N_15370);
or U16379 (N_16379,N_15434,N_15469);
or U16380 (N_16380,N_15944,N_15033);
or U16381 (N_16381,N_15851,N_15274);
nand U16382 (N_16382,N_15541,N_15002);
xnor U16383 (N_16383,N_15332,N_15984);
nor U16384 (N_16384,N_15235,N_15588);
nand U16385 (N_16385,N_15771,N_15398);
or U16386 (N_16386,N_15758,N_15221);
nor U16387 (N_16387,N_15968,N_15143);
and U16388 (N_16388,N_15047,N_15694);
or U16389 (N_16389,N_15481,N_15294);
or U16390 (N_16390,N_15966,N_15834);
xor U16391 (N_16391,N_15284,N_15507);
and U16392 (N_16392,N_15687,N_15179);
or U16393 (N_16393,N_15520,N_15546);
nand U16394 (N_16394,N_15380,N_15287);
nand U16395 (N_16395,N_15997,N_15663);
and U16396 (N_16396,N_15707,N_15819);
nand U16397 (N_16397,N_15631,N_15074);
xor U16398 (N_16398,N_15725,N_15341);
or U16399 (N_16399,N_15465,N_15048);
nor U16400 (N_16400,N_15059,N_15704);
nor U16401 (N_16401,N_15032,N_15057);
or U16402 (N_16402,N_15270,N_15642);
nor U16403 (N_16403,N_15637,N_15403);
and U16404 (N_16404,N_15139,N_15310);
or U16405 (N_16405,N_15585,N_15575);
and U16406 (N_16406,N_15243,N_15196);
or U16407 (N_16407,N_15974,N_15569);
xor U16408 (N_16408,N_15419,N_15365);
and U16409 (N_16409,N_15135,N_15170);
xnor U16410 (N_16410,N_15702,N_15321);
nand U16411 (N_16411,N_15878,N_15412);
xnor U16412 (N_16412,N_15719,N_15756);
nand U16413 (N_16413,N_15551,N_15806);
and U16414 (N_16414,N_15925,N_15011);
and U16415 (N_16415,N_15005,N_15364);
nand U16416 (N_16416,N_15413,N_15544);
nand U16417 (N_16417,N_15843,N_15233);
nand U16418 (N_16418,N_15858,N_15035);
or U16419 (N_16419,N_15824,N_15329);
or U16420 (N_16420,N_15250,N_15432);
nor U16421 (N_16421,N_15151,N_15072);
nor U16422 (N_16422,N_15425,N_15916);
xnor U16423 (N_16423,N_15510,N_15338);
and U16424 (N_16424,N_15159,N_15872);
xnor U16425 (N_16425,N_15205,N_15255);
and U16426 (N_16426,N_15407,N_15092);
nand U16427 (N_16427,N_15056,N_15140);
xor U16428 (N_16428,N_15220,N_15847);
and U16429 (N_16429,N_15775,N_15316);
nor U16430 (N_16430,N_15605,N_15030);
nand U16431 (N_16431,N_15331,N_15271);
nand U16432 (N_16432,N_15523,N_15394);
and U16433 (N_16433,N_15334,N_15443);
or U16434 (N_16434,N_15776,N_15584);
nor U16435 (N_16435,N_15462,N_15941);
nor U16436 (N_16436,N_15323,N_15579);
nor U16437 (N_16437,N_15400,N_15493);
xnor U16438 (N_16438,N_15972,N_15144);
or U16439 (N_16439,N_15213,N_15063);
nand U16440 (N_16440,N_15315,N_15979);
nand U16441 (N_16441,N_15460,N_15573);
nor U16442 (N_16442,N_15591,N_15526);
nand U16443 (N_16443,N_15306,N_15947);
nand U16444 (N_16444,N_15616,N_15561);
or U16445 (N_16445,N_15169,N_15117);
xor U16446 (N_16446,N_15572,N_15390);
xnor U16447 (N_16447,N_15901,N_15672);
and U16448 (N_16448,N_15371,N_15993);
nand U16449 (N_16449,N_15743,N_15745);
xor U16450 (N_16450,N_15759,N_15446);
xnor U16451 (N_16451,N_15684,N_15506);
nor U16452 (N_16452,N_15417,N_15001);
nor U16453 (N_16453,N_15207,N_15505);
or U16454 (N_16454,N_15644,N_15301);
nor U16455 (N_16455,N_15936,N_15492);
and U16456 (N_16456,N_15406,N_15715);
nor U16457 (N_16457,N_15328,N_15118);
nor U16458 (N_16458,N_15244,N_15357);
and U16459 (N_16459,N_15559,N_15594);
xor U16460 (N_16460,N_15098,N_15769);
or U16461 (N_16461,N_15962,N_15934);
and U16462 (N_16462,N_15486,N_15016);
xor U16463 (N_16463,N_15732,N_15850);
xor U16464 (N_16464,N_15111,N_15661);
nor U16465 (N_16465,N_15410,N_15809);
and U16466 (N_16466,N_15906,N_15841);
xor U16467 (N_16467,N_15527,N_15142);
or U16468 (N_16468,N_15564,N_15102);
and U16469 (N_16469,N_15089,N_15639);
nand U16470 (N_16470,N_15194,N_15904);
or U16471 (N_16471,N_15735,N_15852);
or U16472 (N_16472,N_15517,N_15634);
xor U16473 (N_16473,N_15202,N_15209);
xor U16474 (N_16474,N_15949,N_15899);
nand U16475 (N_16475,N_15242,N_15500);
and U16476 (N_16476,N_15065,N_15078);
nand U16477 (N_16477,N_15006,N_15175);
or U16478 (N_16478,N_15986,N_15508);
nand U16479 (N_16479,N_15681,N_15683);
xnor U16480 (N_16480,N_15130,N_15861);
nand U16481 (N_16481,N_15832,N_15738);
and U16482 (N_16482,N_15954,N_15457);
nand U16483 (N_16483,N_15466,N_15485);
nor U16484 (N_16484,N_15362,N_15470);
xnor U16485 (N_16485,N_15474,N_15865);
or U16486 (N_16486,N_15345,N_15180);
nand U16487 (N_16487,N_15880,N_15963);
nor U16488 (N_16488,N_15504,N_15846);
and U16489 (N_16489,N_15015,N_15382);
nor U16490 (N_16490,N_15054,N_15246);
xnor U16491 (N_16491,N_15096,N_15265);
nor U16492 (N_16492,N_15185,N_15764);
nand U16493 (N_16493,N_15753,N_15877);
xnor U16494 (N_16494,N_15249,N_15478);
nor U16495 (N_16495,N_15755,N_15740);
nand U16496 (N_16496,N_15940,N_15038);
or U16497 (N_16497,N_15788,N_15538);
nor U16498 (N_16498,N_15626,N_15027);
and U16499 (N_16499,N_15727,N_15122);
or U16500 (N_16500,N_15551,N_15469);
xnor U16501 (N_16501,N_15201,N_15441);
nor U16502 (N_16502,N_15060,N_15398);
xnor U16503 (N_16503,N_15857,N_15792);
xor U16504 (N_16504,N_15380,N_15992);
or U16505 (N_16505,N_15920,N_15191);
nand U16506 (N_16506,N_15817,N_15970);
nor U16507 (N_16507,N_15041,N_15115);
nor U16508 (N_16508,N_15801,N_15304);
and U16509 (N_16509,N_15797,N_15189);
nand U16510 (N_16510,N_15403,N_15082);
or U16511 (N_16511,N_15461,N_15759);
and U16512 (N_16512,N_15135,N_15540);
nand U16513 (N_16513,N_15565,N_15370);
xnor U16514 (N_16514,N_15278,N_15339);
nand U16515 (N_16515,N_15167,N_15914);
or U16516 (N_16516,N_15892,N_15663);
xor U16517 (N_16517,N_15274,N_15087);
nand U16518 (N_16518,N_15620,N_15157);
or U16519 (N_16519,N_15793,N_15261);
nand U16520 (N_16520,N_15024,N_15539);
and U16521 (N_16521,N_15160,N_15099);
nand U16522 (N_16522,N_15929,N_15344);
or U16523 (N_16523,N_15167,N_15720);
nand U16524 (N_16524,N_15147,N_15612);
or U16525 (N_16525,N_15924,N_15584);
and U16526 (N_16526,N_15883,N_15743);
and U16527 (N_16527,N_15531,N_15254);
nand U16528 (N_16528,N_15427,N_15224);
nor U16529 (N_16529,N_15931,N_15841);
or U16530 (N_16530,N_15998,N_15310);
nor U16531 (N_16531,N_15766,N_15972);
xor U16532 (N_16532,N_15353,N_15106);
or U16533 (N_16533,N_15522,N_15040);
nor U16534 (N_16534,N_15901,N_15148);
or U16535 (N_16535,N_15724,N_15895);
nor U16536 (N_16536,N_15848,N_15292);
and U16537 (N_16537,N_15339,N_15204);
nor U16538 (N_16538,N_15399,N_15623);
or U16539 (N_16539,N_15457,N_15902);
xor U16540 (N_16540,N_15529,N_15758);
xor U16541 (N_16541,N_15336,N_15297);
or U16542 (N_16542,N_15919,N_15318);
and U16543 (N_16543,N_15841,N_15240);
or U16544 (N_16544,N_15362,N_15740);
or U16545 (N_16545,N_15254,N_15955);
xor U16546 (N_16546,N_15473,N_15382);
xor U16547 (N_16547,N_15417,N_15524);
xnor U16548 (N_16548,N_15507,N_15093);
nor U16549 (N_16549,N_15932,N_15733);
nand U16550 (N_16550,N_15113,N_15056);
nand U16551 (N_16551,N_15505,N_15609);
xor U16552 (N_16552,N_15514,N_15995);
and U16553 (N_16553,N_15604,N_15508);
nand U16554 (N_16554,N_15267,N_15792);
nand U16555 (N_16555,N_15367,N_15196);
or U16556 (N_16556,N_15199,N_15780);
and U16557 (N_16557,N_15247,N_15574);
or U16558 (N_16558,N_15273,N_15523);
nand U16559 (N_16559,N_15861,N_15463);
nor U16560 (N_16560,N_15048,N_15203);
or U16561 (N_16561,N_15267,N_15154);
xnor U16562 (N_16562,N_15768,N_15065);
nand U16563 (N_16563,N_15335,N_15232);
and U16564 (N_16564,N_15936,N_15673);
nand U16565 (N_16565,N_15118,N_15138);
or U16566 (N_16566,N_15614,N_15851);
nor U16567 (N_16567,N_15079,N_15276);
nor U16568 (N_16568,N_15996,N_15885);
and U16569 (N_16569,N_15449,N_15094);
nand U16570 (N_16570,N_15676,N_15794);
nor U16571 (N_16571,N_15823,N_15847);
or U16572 (N_16572,N_15495,N_15144);
nor U16573 (N_16573,N_15761,N_15840);
xnor U16574 (N_16574,N_15354,N_15382);
nor U16575 (N_16575,N_15630,N_15126);
or U16576 (N_16576,N_15090,N_15379);
and U16577 (N_16577,N_15737,N_15087);
or U16578 (N_16578,N_15666,N_15906);
and U16579 (N_16579,N_15328,N_15917);
xnor U16580 (N_16580,N_15279,N_15542);
xor U16581 (N_16581,N_15316,N_15764);
or U16582 (N_16582,N_15198,N_15281);
and U16583 (N_16583,N_15300,N_15876);
nand U16584 (N_16584,N_15745,N_15961);
and U16585 (N_16585,N_15600,N_15756);
or U16586 (N_16586,N_15022,N_15019);
and U16587 (N_16587,N_15444,N_15202);
xor U16588 (N_16588,N_15248,N_15336);
nand U16589 (N_16589,N_15989,N_15721);
or U16590 (N_16590,N_15408,N_15862);
nor U16591 (N_16591,N_15429,N_15162);
nor U16592 (N_16592,N_15728,N_15918);
and U16593 (N_16593,N_15251,N_15132);
or U16594 (N_16594,N_15773,N_15271);
nor U16595 (N_16595,N_15476,N_15357);
nand U16596 (N_16596,N_15894,N_15689);
and U16597 (N_16597,N_15521,N_15967);
nand U16598 (N_16598,N_15640,N_15397);
or U16599 (N_16599,N_15011,N_15289);
nand U16600 (N_16600,N_15023,N_15671);
or U16601 (N_16601,N_15900,N_15064);
xor U16602 (N_16602,N_15146,N_15548);
xor U16603 (N_16603,N_15989,N_15564);
and U16604 (N_16604,N_15893,N_15699);
nor U16605 (N_16605,N_15192,N_15997);
and U16606 (N_16606,N_15821,N_15741);
and U16607 (N_16607,N_15395,N_15954);
or U16608 (N_16608,N_15360,N_15201);
xnor U16609 (N_16609,N_15956,N_15030);
nand U16610 (N_16610,N_15051,N_15519);
or U16611 (N_16611,N_15386,N_15368);
or U16612 (N_16612,N_15550,N_15585);
and U16613 (N_16613,N_15912,N_15734);
xor U16614 (N_16614,N_15677,N_15283);
nor U16615 (N_16615,N_15401,N_15550);
nand U16616 (N_16616,N_15718,N_15895);
nor U16617 (N_16617,N_15670,N_15553);
nor U16618 (N_16618,N_15237,N_15359);
and U16619 (N_16619,N_15969,N_15513);
nand U16620 (N_16620,N_15891,N_15477);
nand U16621 (N_16621,N_15642,N_15851);
nand U16622 (N_16622,N_15721,N_15944);
nor U16623 (N_16623,N_15759,N_15331);
nand U16624 (N_16624,N_15954,N_15003);
or U16625 (N_16625,N_15454,N_15076);
nand U16626 (N_16626,N_15388,N_15474);
nand U16627 (N_16627,N_15209,N_15996);
or U16628 (N_16628,N_15372,N_15076);
xor U16629 (N_16629,N_15550,N_15744);
nand U16630 (N_16630,N_15695,N_15483);
xor U16631 (N_16631,N_15130,N_15441);
xor U16632 (N_16632,N_15755,N_15108);
and U16633 (N_16633,N_15813,N_15410);
nor U16634 (N_16634,N_15776,N_15092);
and U16635 (N_16635,N_15986,N_15627);
nor U16636 (N_16636,N_15156,N_15519);
nor U16637 (N_16637,N_15591,N_15862);
and U16638 (N_16638,N_15300,N_15499);
or U16639 (N_16639,N_15703,N_15643);
xor U16640 (N_16640,N_15854,N_15266);
xor U16641 (N_16641,N_15248,N_15109);
and U16642 (N_16642,N_15043,N_15698);
and U16643 (N_16643,N_15644,N_15237);
nor U16644 (N_16644,N_15723,N_15881);
nand U16645 (N_16645,N_15022,N_15656);
nor U16646 (N_16646,N_15381,N_15823);
or U16647 (N_16647,N_15834,N_15015);
nand U16648 (N_16648,N_15042,N_15674);
or U16649 (N_16649,N_15853,N_15167);
nor U16650 (N_16650,N_15303,N_15518);
xor U16651 (N_16651,N_15449,N_15459);
nor U16652 (N_16652,N_15694,N_15674);
nand U16653 (N_16653,N_15527,N_15710);
or U16654 (N_16654,N_15770,N_15780);
xnor U16655 (N_16655,N_15164,N_15452);
and U16656 (N_16656,N_15632,N_15474);
nor U16657 (N_16657,N_15399,N_15379);
xor U16658 (N_16658,N_15162,N_15763);
xnor U16659 (N_16659,N_15617,N_15143);
nand U16660 (N_16660,N_15266,N_15431);
or U16661 (N_16661,N_15548,N_15035);
nand U16662 (N_16662,N_15101,N_15637);
and U16663 (N_16663,N_15885,N_15028);
xor U16664 (N_16664,N_15702,N_15172);
xor U16665 (N_16665,N_15445,N_15792);
nand U16666 (N_16666,N_15969,N_15022);
nand U16667 (N_16667,N_15864,N_15458);
nor U16668 (N_16668,N_15448,N_15808);
nor U16669 (N_16669,N_15255,N_15072);
nand U16670 (N_16670,N_15323,N_15960);
nand U16671 (N_16671,N_15048,N_15552);
or U16672 (N_16672,N_15611,N_15473);
nor U16673 (N_16673,N_15744,N_15268);
xnor U16674 (N_16674,N_15721,N_15786);
or U16675 (N_16675,N_15710,N_15700);
and U16676 (N_16676,N_15334,N_15414);
or U16677 (N_16677,N_15758,N_15690);
or U16678 (N_16678,N_15487,N_15599);
nor U16679 (N_16679,N_15377,N_15555);
xnor U16680 (N_16680,N_15959,N_15111);
nand U16681 (N_16681,N_15840,N_15131);
nor U16682 (N_16682,N_15502,N_15078);
and U16683 (N_16683,N_15195,N_15836);
nand U16684 (N_16684,N_15807,N_15271);
nand U16685 (N_16685,N_15326,N_15299);
xor U16686 (N_16686,N_15364,N_15726);
and U16687 (N_16687,N_15275,N_15878);
or U16688 (N_16688,N_15686,N_15207);
or U16689 (N_16689,N_15075,N_15622);
or U16690 (N_16690,N_15467,N_15364);
nand U16691 (N_16691,N_15840,N_15802);
xnor U16692 (N_16692,N_15890,N_15755);
nand U16693 (N_16693,N_15520,N_15899);
or U16694 (N_16694,N_15971,N_15434);
nor U16695 (N_16695,N_15627,N_15681);
and U16696 (N_16696,N_15628,N_15357);
nand U16697 (N_16697,N_15617,N_15068);
nand U16698 (N_16698,N_15489,N_15110);
or U16699 (N_16699,N_15442,N_15681);
xor U16700 (N_16700,N_15121,N_15366);
and U16701 (N_16701,N_15705,N_15956);
nor U16702 (N_16702,N_15761,N_15694);
and U16703 (N_16703,N_15578,N_15979);
xor U16704 (N_16704,N_15652,N_15540);
xor U16705 (N_16705,N_15970,N_15455);
or U16706 (N_16706,N_15266,N_15880);
nand U16707 (N_16707,N_15952,N_15219);
or U16708 (N_16708,N_15430,N_15275);
nand U16709 (N_16709,N_15540,N_15036);
xor U16710 (N_16710,N_15418,N_15438);
nor U16711 (N_16711,N_15896,N_15253);
or U16712 (N_16712,N_15374,N_15902);
xor U16713 (N_16713,N_15341,N_15644);
xor U16714 (N_16714,N_15509,N_15436);
and U16715 (N_16715,N_15861,N_15969);
nor U16716 (N_16716,N_15041,N_15130);
nand U16717 (N_16717,N_15358,N_15609);
xnor U16718 (N_16718,N_15543,N_15716);
or U16719 (N_16719,N_15762,N_15278);
and U16720 (N_16720,N_15220,N_15035);
or U16721 (N_16721,N_15015,N_15259);
nand U16722 (N_16722,N_15996,N_15526);
nand U16723 (N_16723,N_15064,N_15754);
and U16724 (N_16724,N_15554,N_15238);
xnor U16725 (N_16725,N_15793,N_15766);
xor U16726 (N_16726,N_15976,N_15737);
nor U16727 (N_16727,N_15638,N_15619);
nor U16728 (N_16728,N_15983,N_15445);
nand U16729 (N_16729,N_15325,N_15338);
and U16730 (N_16730,N_15526,N_15565);
xor U16731 (N_16731,N_15528,N_15460);
and U16732 (N_16732,N_15793,N_15181);
and U16733 (N_16733,N_15678,N_15599);
xnor U16734 (N_16734,N_15699,N_15318);
and U16735 (N_16735,N_15530,N_15460);
or U16736 (N_16736,N_15587,N_15166);
or U16737 (N_16737,N_15804,N_15811);
nor U16738 (N_16738,N_15649,N_15552);
xor U16739 (N_16739,N_15624,N_15778);
nor U16740 (N_16740,N_15642,N_15886);
xor U16741 (N_16741,N_15815,N_15210);
or U16742 (N_16742,N_15739,N_15963);
nand U16743 (N_16743,N_15281,N_15372);
and U16744 (N_16744,N_15071,N_15860);
nand U16745 (N_16745,N_15610,N_15465);
xnor U16746 (N_16746,N_15574,N_15146);
nor U16747 (N_16747,N_15897,N_15796);
or U16748 (N_16748,N_15759,N_15631);
or U16749 (N_16749,N_15685,N_15200);
or U16750 (N_16750,N_15836,N_15486);
and U16751 (N_16751,N_15538,N_15077);
nand U16752 (N_16752,N_15980,N_15680);
nand U16753 (N_16753,N_15126,N_15508);
or U16754 (N_16754,N_15385,N_15883);
and U16755 (N_16755,N_15292,N_15231);
nand U16756 (N_16756,N_15904,N_15350);
and U16757 (N_16757,N_15915,N_15430);
xor U16758 (N_16758,N_15302,N_15812);
xor U16759 (N_16759,N_15420,N_15462);
and U16760 (N_16760,N_15779,N_15610);
nand U16761 (N_16761,N_15922,N_15129);
nor U16762 (N_16762,N_15738,N_15051);
xnor U16763 (N_16763,N_15427,N_15378);
nor U16764 (N_16764,N_15893,N_15792);
xnor U16765 (N_16765,N_15179,N_15051);
nor U16766 (N_16766,N_15225,N_15954);
or U16767 (N_16767,N_15110,N_15239);
xnor U16768 (N_16768,N_15598,N_15518);
or U16769 (N_16769,N_15533,N_15423);
and U16770 (N_16770,N_15311,N_15231);
nand U16771 (N_16771,N_15727,N_15650);
nor U16772 (N_16772,N_15588,N_15360);
and U16773 (N_16773,N_15943,N_15860);
xnor U16774 (N_16774,N_15997,N_15495);
xor U16775 (N_16775,N_15670,N_15918);
nand U16776 (N_16776,N_15612,N_15542);
xnor U16777 (N_16777,N_15123,N_15665);
nor U16778 (N_16778,N_15990,N_15441);
nor U16779 (N_16779,N_15534,N_15214);
nor U16780 (N_16780,N_15416,N_15820);
and U16781 (N_16781,N_15966,N_15301);
and U16782 (N_16782,N_15625,N_15247);
nand U16783 (N_16783,N_15098,N_15644);
nand U16784 (N_16784,N_15195,N_15345);
or U16785 (N_16785,N_15001,N_15464);
and U16786 (N_16786,N_15516,N_15554);
and U16787 (N_16787,N_15389,N_15066);
nand U16788 (N_16788,N_15725,N_15102);
and U16789 (N_16789,N_15645,N_15141);
xnor U16790 (N_16790,N_15531,N_15985);
or U16791 (N_16791,N_15117,N_15687);
nand U16792 (N_16792,N_15700,N_15569);
xnor U16793 (N_16793,N_15822,N_15222);
xnor U16794 (N_16794,N_15589,N_15309);
xnor U16795 (N_16795,N_15351,N_15764);
xor U16796 (N_16796,N_15650,N_15062);
nand U16797 (N_16797,N_15137,N_15465);
nor U16798 (N_16798,N_15464,N_15688);
nor U16799 (N_16799,N_15650,N_15477);
nand U16800 (N_16800,N_15808,N_15480);
nor U16801 (N_16801,N_15336,N_15892);
nor U16802 (N_16802,N_15936,N_15546);
xnor U16803 (N_16803,N_15470,N_15012);
nor U16804 (N_16804,N_15088,N_15913);
nand U16805 (N_16805,N_15675,N_15559);
and U16806 (N_16806,N_15915,N_15681);
or U16807 (N_16807,N_15441,N_15044);
or U16808 (N_16808,N_15179,N_15437);
nand U16809 (N_16809,N_15119,N_15514);
or U16810 (N_16810,N_15989,N_15192);
and U16811 (N_16811,N_15959,N_15945);
or U16812 (N_16812,N_15136,N_15552);
nor U16813 (N_16813,N_15634,N_15289);
and U16814 (N_16814,N_15038,N_15377);
nor U16815 (N_16815,N_15609,N_15159);
xnor U16816 (N_16816,N_15029,N_15355);
nand U16817 (N_16817,N_15764,N_15278);
nand U16818 (N_16818,N_15862,N_15661);
nand U16819 (N_16819,N_15517,N_15478);
and U16820 (N_16820,N_15809,N_15591);
nand U16821 (N_16821,N_15375,N_15795);
xor U16822 (N_16822,N_15683,N_15739);
and U16823 (N_16823,N_15761,N_15220);
xnor U16824 (N_16824,N_15624,N_15348);
nor U16825 (N_16825,N_15512,N_15587);
and U16826 (N_16826,N_15199,N_15137);
nand U16827 (N_16827,N_15668,N_15587);
or U16828 (N_16828,N_15765,N_15362);
and U16829 (N_16829,N_15826,N_15824);
and U16830 (N_16830,N_15026,N_15308);
nor U16831 (N_16831,N_15493,N_15971);
xor U16832 (N_16832,N_15871,N_15582);
nand U16833 (N_16833,N_15284,N_15626);
and U16834 (N_16834,N_15963,N_15961);
nor U16835 (N_16835,N_15286,N_15053);
and U16836 (N_16836,N_15693,N_15732);
nor U16837 (N_16837,N_15125,N_15239);
xnor U16838 (N_16838,N_15933,N_15569);
nand U16839 (N_16839,N_15418,N_15217);
nor U16840 (N_16840,N_15482,N_15188);
nor U16841 (N_16841,N_15200,N_15765);
nor U16842 (N_16842,N_15514,N_15460);
nand U16843 (N_16843,N_15915,N_15814);
and U16844 (N_16844,N_15263,N_15303);
xor U16845 (N_16845,N_15619,N_15414);
or U16846 (N_16846,N_15782,N_15806);
xnor U16847 (N_16847,N_15385,N_15499);
nor U16848 (N_16848,N_15643,N_15324);
and U16849 (N_16849,N_15015,N_15345);
xnor U16850 (N_16850,N_15487,N_15139);
or U16851 (N_16851,N_15280,N_15063);
nor U16852 (N_16852,N_15381,N_15610);
and U16853 (N_16853,N_15894,N_15191);
nand U16854 (N_16854,N_15847,N_15398);
xor U16855 (N_16855,N_15537,N_15097);
or U16856 (N_16856,N_15733,N_15034);
xor U16857 (N_16857,N_15553,N_15396);
and U16858 (N_16858,N_15961,N_15181);
xor U16859 (N_16859,N_15405,N_15465);
xor U16860 (N_16860,N_15364,N_15553);
nand U16861 (N_16861,N_15061,N_15468);
nor U16862 (N_16862,N_15149,N_15583);
xnor U16863 (N_16863,N_15450,N_15961);
or U16864 (N_16864,N_15447,N_15272);
and U16865 (N_16865,N_15722,N_15915);
nor U16866 (N_16866,N_15519,N_15749);
nor U16867 (N_16867,N_15738,N_15112);
xnor U16868 (N_16868,N_15835,N_15472);
and U16869 (N_16869,N_15905,N_15108);
nand U16870 (N_16870,N_15816,N_15334);
and U16871 (N_16871,N_15128,N_15553);
nand U16872 (N_16872,N_15065,N_15412);
nor U16873 (N_16873,N_15207,N_15020);
xor U16874 (N_16874,N_15967,N_15487);
nand U16875 (N_16875,N_15010,N_15336);
nand U16876 (N_16876,N_15563,N_15668);
nand U16877 (N_16877,N_15553,N_15654);
or U16878 (N_16878,N_15203,N_15313);
or U16879 (N_16879,N_15166,N_15296);
xnor U16880 (N_16880,N_15471,N_15954);
and U16881 (N_16881,N_15616,N_15231);
nor U16882 (N_16882,N_15308,N_15511);
xnor U16883 (N_16883,N_15413,N_15324);
and U16884 (N_16884,N_15296,N_15127);
or U16885 (N_16885,N_15039,N_15720);
xor U16886 (N_16886,N_15705,N_15927);
and U16887 (N_16887,N_15540,N_15446);
xor U16888 (N_16888,N_15666,N_15199);
nand U16889 (N_16889,N_15895,N_15814);
nand U16890 (N_16890,N_15377,N_15950);
xnor U16891 (N_16891,N_15873,N_15213);
and U16892 (N_16892,N_15871,N_15149);
nor U16893 (N_16893,N_15815,N_15080);
nor U16894 (N_16894,N_15934,N_15158);
or U16895 (N_16895,N_15526,N_15615);
xnor U16896 (N_16896,N_15791,N_15610);
and U16897 (N_16897,N_15989,N_15410);
xor U16898 (N_16898,N_15596,N_15814);
and U16899 (N_16899,N_15758,N_15391);
or U16900 (N_16900,N_15878,N_15235);
xnor U16901 (N_16901,N_15395,N_15964);
xor U16902 (N_16902,N_15905,N_15466);
and U16903 (N_16903,N_15551,N_15430);
or U16904 (N_16904,N_15069,N_15638);
and U16905 (N_16905,N_15900,N_15041);
nand U16906 (N_16906,N_15413,N_15046);
or U16907 (N_16907,N_15890,N_15634);
nor U16908 (N_16908,N_15372,N_15486);
xnor U16909 (N_16909,N_15014,N_15217);
nand U16910 (N_16910,N_15283,N_15756);
nand U16911 (N_16911,N_15441,N_15868);
or U16912 (N_16912,N_15315,N_15227);
xor U16913 (N_16913,N_15135,N_15647);
nand U16914 (N_16914,N_15777,N_15642);
and U16915 (N_16915,N_15151,N_15006);
nand U16916 (N_16916,N_15935,N_15389);
or U16917 (N_16917,N_15808,N_15012);
nor U16918 (N_16918,N_15940,N_15049);
nand U16919 (N_16919,N_15452,N_15444);
and U16920 (N_16920,N_15380,N_15770);
nor U16921 (N_16921,N_15355,N_15843);
nor U16922 (N_16922,N_15132,N_15342);
nand U16923 (N_16923,N_15331,N_15857);
and U16924 (N_16924,N_15066,N_15803);
or U16925 (N_16925,N_15313,N_15592);
nor U16926 (N_16926,N_15070,N_15596);
or U16927 (N_16927,N_15881,N_15454);
xnor U16928 (N_16928,N_15825,N_15258);
xor U16929 (N_16929,N_15345,N_15119);
nand U16930 (N_16930,N_15104,N_15224);
xnor U16931 (N_16931,N_15817,N_15743);
nand U16932 (N_16932,N_15968,N_15014);
xor U16933 (N_16933,N_15137,N_15698);
xnor U16934 (N_16934,N_15730,N_15951);
nand U16935 (N_16935,N_15873,N_15740);
or U16936 (N_16936,N_15978,N_15996);
nand U16937 (N_16937,N_15659,N_15739);
nor U16938 (N_16938,N_15857,N_15407);
xnor U16939 (N_16939,N_15549,N_15528);
or U16940 (N_16940,N_15444,N_15107);
or U16941 (N_16941,N_15781,N_15432);
and U16942 (N_16942,N_15585,N_15031);
xnor U16943 (N_16943,N_15299,N_15613);
nor U16944 (N_16944,N_15730,N_15729);
and U16945 (N_16945,N_15104,N_15769);
xnor U16946 (N_16946,N_15204,N_15764);
and U16947 (N_16947,N_15891,N_15886);
xnor U16948 (N_16948,N_15814,N_15795);
nand U16949 (N_16949,N_15224,N_15378);
nor U16950 (N_16950,N_15734,N_15271);
nand U16951 (N_16951,N_15164,N_15324);
nand U16952 (N_16952,N_15558,N_15609);
and U16953 (N_16953,N_15607,N_15674);
nor U16954 (N_16954,N_15109,N_15439);
xor U16955 (N_16955,N_15276,N_15128);
nor U16956 (N_16956,N_15431,N_15924);
or U16957 (N_16957,N_15213,N_15658);
nor U16958 (N_16958,N_15162,N_15732);
or U16959 (N_16959,N_15578,N_15349);
nand U16960 (N_16960,N_15839,N_15408);
nand U16961 (N_16961,N_15087,N_15122);
xor U16962 (N_16962,N_15201,N_15489);
and U16963 (N_16963,N_15852,N_15630);
nor U16964 (N_16964,N_15682,N_15522);
nand U16965 (N_16965,N_15081,N_15567);
nor U16966 (N_16966,N_15896,N_15039);
nor U16967 (N_16967,N_15178,N_15403);
and U16968 (N_16968,N_15809,N_15781);
and U16969 (N_16969,N_15308,N_15881);
or U16970 (N_16970,N_15326,N_15029);
nor U16971 (N_16971,N_15433,N_15617);
xnor U16972 (N_16972,N_15083,N_15214);
or U16973 (N_16973,N_15171,N_15185);
and U16974 (N_16974,N_15714,N_15622);
and U16975 (N_16975,N_15329,N_15797);
and U16976 (N_16976,N_15373,N_15211);
nor U16977 (N_16977,N_15087,N_15524);
or U16978 (N_16978,N_15314,N_15069);
xor U16979 (N_16979,N_15328,N_15620);
nor U16980 (N_16980,N_15407,N_15915);
or U16981 (N_16981,N_15263,N_15433);
nand U16982 (N_16982,N_15382,N_15541);
xor U16983 (N_16983,N_15169,N_15970);
nor U16984 (N_16984,N_15022,N_15221);
and U16985 (N_16985,N_15758,N_15537);
nand U16986 (N_16986,N_15470,N_15408);
nand U16987 (N_16987,N_15797,N_15806);
nor U16988 (N_16988,N_15293,N_15492);
and U16989 (N_16989,N_15667,N_15370);
nand U16990 (N_16990,N_15747,N_15389);
nand U16991 (N_16991,N_15103,N_15678);
nand U16992 (N_16992,N_15666,N_15962);
nand U16993 (N_16993,N_15959,N_15755);
nor U16994 (N_16994,N_15742,N_15925);
or U16995 (N_16995,N_15300,N_15097);
nor U16996 (N_16996,N_15026,N_15905);
nor U16997 (N_16997,N_15297,N_15819);
nor U16998 (N_16998,N_15961,N_15643);
or U16999 (N_16999,N_15856,N_15249);
nor U17000 (N_17000,N_16648,N_16344);
or U17001 (N_17001,N_16674,N_16859);
nand U17002 (N_17002,N_16407,N_16329);
nand U17003 (N_17003,N_16378,N_16755);
nor U17004 (N_17004,N_16541,N_16372);
nor U17005 (N_17005,N_16932,N_16895);
nand U17006 (N_17006,N_16984,N_16621);
or U17007 (N_17007,N_16906,N_16682);
nand U17008 (N_17008,N_16708,N_16321);
xnor U17009 (N_17009,N_16221,N_16093);
nand U17010 (N_17010,N_16518,N_16588);
nand U17011 (N_17011,N_16752,N_16606);
or U17012 (N_17012,N_16560,N_16150);
nand U17013 (N_17013,N_16454,N_16696);
and U17014 (N_17014,N_16631,N_16624);
nor U17015 (N_17015,N_16191,N_16431);
nor U17016 (N_17016,N_16449,N_16699);
nand U17017 (N_17017,N_16297,N_16470);
xnor U17018 (N_17018,N_16172,N_16780);
nor U17019 (N_17019,N_16576,N_16641);
xor U17020 (N_17020,N_16957,N_16205);
nor U17021 (N_17021,N_16281,N_16626);
nand U17022 (N_17022,N_16800,N_16178);
nor U17023 (N_17023,N_16254,N_16760);
or U17024 (N_17024,N_16818,N_16291);
xnor U17025 (N_17025,N_16202,N_16968);
xor U17026 (N_17026,N_16990,N_16060);
nand U17027 (N_17027,N_16869,N_16052);
xnor U17028 (N_17028,N_16128,N_16652);
and U17029 (N_17029,N_16843,N_16704);
nor U17030 (N_17030,N_16724,N_16815);
or U17031 (N_17031,N_16305,N_16979);
nor U17032 (N_17032,N_16424,N_16328);
nand U17033 (N_17033,N_16034,N_16529);
nor U17034 (N_17034,N_16551,N_16428);
nand U17035 (N_17035,N_16583,N_16725);
nor U17036 (N_17036,N_16850,N_16183);
nand U17037 (N_17037,N_16473,N_16582);
xnor U17038 (N_17038,N_16914,N_16059);
nor U17039 (N_17039,N_16065,N_16834);
and U17040 (N_17040,N_16103,N_16279);
nor U17041 (N_17041,N_16090,N_16591);
xor U17042 (N_17042,N_16601,N_16115);
xor U17043 (N_17043,N_16675,N_16379);
or U17044 (N_17044,N_16846,N_16743);
xnor U17045 (N_17045,N_16444,N_16534);
nand U17046 (N_17046,N_16478,N_16862);
nor U17047 (N_17047,N_16233,N_16505);
nor U17048 (N_17048,N_16463,N_16326);
xor U17049 (N_17049,N_16717,N_16796);
or U17050 (N_17050,N_16058,N_16822);
nor U17051 (N_17051,N_16738,N_16828);
or U17052 (N_17052,N_16075,N_16167);
xor U17053 (N_17053,N_16019,N_16426);
and U17054 (N_17054,N_16746,N_16298);
nor U17055 (N_17055,N_16734,N_16711);
and U17056 (N_17056,N_16294,N_16779);
nor U17057 (N_17057,N_16055,N_16563);
or U17058 (N_17058,N_16113,N_16035);
xor U17059 (N_17059,N_16311,N_16559);
and U17060 (N_17060,N_16083,N_16340);
nor U17061 (N_17061,N_16067,N_16215);
nor U17062 (N_17062,N_16510,N_16129);
nor U17063 (N_17063,N_16912,N_16749);
and U17064 (N_17064,N_16471,N_16047);
nor U17065 (N_17065,N_16741,N_16369);
or U17066 (N_17066,N_16848,N_16185);
or U17067 (N_17067,N_16812,N_16341);
or U17068 (N_17068,N_16985,N_16343);
xor U17069 (N_17069,N_16893,N_16229);
or U17070 (N_17070,N_16509,N_16671);
and U17071 (N_17071,N_16520,N_16657);
nor U17072 (N_17072,N_16439,N_16013);
nor U17073 (N_17073,N_16995,N_16706);
nand U17074 (N_17074,N_16683,N_16147);
xor U17075 (N_17075,N_16345,N_16765);
and U17076 (N_17076,N_16646,N_16920);
and U17077 (N_17077,N_16049,N_16645);
and U17078 (N_17078,N_16468,N_16080);
or U17079 (N_17079,N_16698,N_16756);
nor U17080 (N_17080,N_16353,N_16038);
nor U17081 (N_17081,N_16293,N_16209);
or U17082 (N_17082,N_16567,N_16351);
and U17083 (N_17083,N_16266,N_16697);
xnor U17084 (N_17084,N_16947,N_16940);
and U17085 (N_17085,N_16029,N_16085);
nand U17086 (N_17086,N_16982,N_16346);
nand U17087 (N_17087,N_16225,N_16307);
xor U17088 (N_17088,N_16974,N_16339);
xnor U17089 (N_17089,N_16836,N_16377);
and U17090 (N_17090,N_16247,N_16519);
or U17091 (N_17091,N_16732,N_16548);
and U17092 (N_17092,N_16317,N_16420);
nand U17093 (N_17093,N_16173,N_16913);
and U17094 (N_17094,N_16039,N_16584);
xnor U17095 (N_17095,N_16903,N_16292);
and U17096 (N_17096,N_16479,N_16056);
xnor U17097 (N_17097,N_16829,N_16003);
nor U17098 (N_17098,N_16441,N_16145);
xor U17099 (N_17099,N_16821,N_16376);
or U17100 (N_17100,N_16112,N_16282);
nor U17101 (N_17101,N_16252,N_16168);
and U17102 (N_17102,N_16174,N_16265);
and U17103 (N_17103,N_16495,N_16415);
nor U17104 (N_17104,N_16585,N_16285);
and U17105 (N_17105,N_16587,N_16599);
or U17106 (N_17106,N_16797,N_16676);
xnor U17107 (N_17107,N_16180,N_16772);
xor U17108 (N_17108,N_16110,N_16048);
and U17109 (N_17109,N_16164,N_16702);
or U17110 (N_17110,N_16506,N_16322);
nand U17111 (N_17111,N_16273,N_16062);
nand U17112 (N_17112,N_16745,N_16199);
and U17113 (N_17113,N_16936,N_16169);
and U17114 (N_17114,N_16161,N_16320);
or U17115 (N_17115,N_16600,N_16270);
and U17116 (N_17116,N_16735,N_16907);
nand U17117 (N_17117,N_16046,N_16027);
nand U17118 (N_17118,N_16958,N_16006);
or U17119 (N_17119,N_16962,N_16955);
or U17120 (N_17120,N_16158,N_16234);
nor U17121 (N_17121,N_16334,N_16627);
xor U17122 (N_17122,N_16018,N_16536);
or U17123 (N_17123,N_16368,N_16805);
nor U17124 (N_17124,N_16200,N_16824);
and U17125 (N_17125,N_16782,N_16988);
xor U17126 (N_17126,N_16036,N_16204);
nor U17127 (N_17127,N_16492,N_16747);
and U17128 (N_17128,N_16261,N_16280);
or U17129 (N_17129,N_16792,N_16950);
and U17130 (N_17130,N_16148,N_16884);
xnor U17131 (N_17131,N_16243,N_16616);
or U17132 (N_17132,N_16357,N_16214);
xnor U17133 (N_17133,N_16461,N_16485);
nand U17134 (N_17134,N_16195,N_16232);
xor U17135 (N_17135,N_16902,N_16935);
nor U17136 (N_17136,N_16143,N_16386);
nor U17137 (N_17137,N_16781,N_16136);
and U17138 (N_17138,N_16690,N_16991);
xnor U17139 (N_17139,N_16121,N_16422);
nand U17140 (N_17140,N_16695,N_16748);
nor U17141 (N_17141,N_16921,N_16020);
or U17142 (N_17142,N_16951,N_16635);
or U17143 (N_17143,N_16486,N_16669);
or U17144 (N_17144,N_16009,N_16632);
nor U17145 (N_17145,N_16474,N_16678);
nand U17146 (N_17146,N_16803,N_16375);
and U17147 (N_17147,N_16452,N_16637);
and U17148 (N_17148,N_16011,N_16758);
nand U17149 (N_17149,N_16533,N_16179);
or U17150 (N_17150,N_16289,N_16466);
or U17151 (N_17151,N_16070,N_16394);
or U17152 (N_17152,N_16728,N_16041);
nand U17153 (N_17153,N_16142,N_16414);
nor U17154 (N_17154,N_16367,N_16566);
or U17155 (N_17155,N_16689,N_16064);
xor U17156 (N_17156,N_16082,N_16686);
and U17157 (N_17157,N_16392,N_16393);
xor U17158 (N_17158,N_16245,N_16944);
xnor U17159 (N_17159,N_16638,N_16483);
or U17160 (N_17160,N_16419,N_16237);
or U17161 (N_17161,N_16881,N_16491);
and U17162 (N_17162,N_16433,N_16457);
or U17163 (N_17163,N_16937,N_16050);
nand U17164 (N_17164,N_16855,N_16943);
nor U17165 (N_17165,N_16998,N_16885);
xnor U17166 (N_17166,N_16839,N_16448);
and U17167 (N_17167,N_16876,N_16999);
nor U17168 (N_17168,N_16889,N_16552);
and U17169 (N_17169,N_16097,N_16840);
nand U17170 (N_17170,N_16010,N_16549);
or U17171 (N_17171,N_16131,N_16666);
and U17172 (N_17172,N_16612,N_16973);
nand U17173 (N_17173,N_16374,N_16092);
or U17174 (N_17174,N_16253,N_16107);
nor U17175 (N_17175,N_16622,N_16832);
nor U17176 (N_17176,N_16417,N_16489);
and U17177 (N_17177,N_16787,N_16198);
or U17178 (N_17178,N_16068,N_16865);
or U17179 (N_17179,N_16916,N_16355);
or U17180 (N_17180,N_16108,N_16714);
and U17181 (N_17181,N_16878,N_16927);
nand U17182 (N_17182,N_16274,N_16146);
nor U17183 (N_17183,N_16399,N_16771);
xnor U17184 (N_17184,N_16924,N_16134);
and U17185 (N_17185,N_16596,N_16182);
nor U17186 (N_17186,N_16153,N_16138);
xnor U17187 (N_17187,N_16565,N_16939);
xnor U17188 (N_17188,N_16459,N_16574);
nor U17189 (N_17189,N_16996,N_16084);
xnor U17190 (N_17190,N_16240,N_16685);
and U17191 (N_17191,N_16740,N_16380);
xor U17192 (N_17192,N_16628,N_16061);
xnor U17193 (N_17193,N_16926,N_16284);
nand U17194 (N_17194,N_16391,N_16443);
xnor U17195 (N_17195,N_16593,N_16469);
nand U17196 (N_17196,N_16531,N_16137);
nand U17197 (N_17197,N_16618,N_16501);
nor U17198 (N_17198,N_16480,N_16201);
nand U17199 (N_17199,N_16109,N_16838);
and U17200 (N_17200,N_16693,N_16316);
nand U17201 (N_17201,N_16929,N_16810);
nand U17202 (N_17202,N_16365,N_16502);
or U17203 (N_17203,N_16928,N_16976);
or U17204 (N_17204,N_16511,N_16946);
xor U17205 (N_17205,N_16713,N_16484);
nand U17206 (N_17206,N_16833,N_16844);
nand U17207 (N_17207,N_16715,N_16421);
and U17208 (N_17208,N_16649,N_16527);
or U17209 (N_17209,N_16120,N_16668);
xor U17210 (N_17210,N_16324,N_16258);
or U17211 (N_17211,N_16409,N_16338);
nand U17212 (N_17212,N_16144,N_16342);
and U17213 (N_17213,N_16362,N_16619);
or U17214 (N_17214,N_16608,N_16319);
or U17215 (N_17215,N_16595,N_16450);
nor U17216 (N_17216,N_16364,N_16660);
xnor U17217 (N_17217,N_16166,N_16387);
or U17218 (N_17218,N_16037,N_16931);
nor U17219 (N_17219,N_16945,N_16042);
and U17220 (N_17220,N_16954,N_16813);
xor U17221 (N_17221,N_16460,N_16707);
and U17222 (N_17222,N_16630,N_16401);
nand U17223 (N_17223,N_16874,N_16575);
xnor U17224 (N_17224,N_16766,N_16425);
xor U17225 (N_17225,N_16301,N_16602);
nor U17226 (N_17226,N_16482,N_16709);
nand U17227 (N_17227,N_16845,N_16790);
or U17228 (N_17228,N_16352,N_16744);
nor U17229 (N_17229,N_16476,N_16272);
nor U17230 (N_17230,N_16323,N_16442);
xnor U17231 (N_17231,N_16858,N_16910);
nor U17232 (N_17232,N_16804,N_16694);
xor U17233 (N_17233,N_16278,N_16639);
xor U17234 (N_17234,N_16408,N_16400);
xnor U17235 (N_17235,N_16592,N_16122);
or U17236 (N_17236,N_16287,N_16680);
or U17237 (N_17237,N_16830,N_16909);
nor U17238 (N_17238,N_16403,N_16523);
xnor U17239 (N_17239,N_16163,N_16700);
and U17240 (N_17240,N_16133,N_16564);
nand U17241 (N_17241,N_16535,N_16462);
xnor U17242 (N_17242,N_16308,N_16892);
nand U17243 (N_17243,N_16262,N_16868);
nand U17244 (N_17244,N_16949,N_16397);
nor U17245 (N_17245,N_16111,N_16794);
nand U17246 (N_17246,N_16942,N_16769);
xor U17247 (N_17247,N_16091,N_16494);
xnor U17248 (N_17248,N_16188,N_16318);
xor U17249 (N_17249,N_16983,N_16647);
nor U17250 (N_17250,N_16739,N_16959);
xor U17251 (N_17251,N_16481,N_16808);
xnor U17252 (N_17252,N_16314,N_16192);
and U17253 (N_17253,N_16132,N_16263);
or U17254 (N_17254,N_16312,N_16860);
or U17255 (N_17255,N_16371,N_16089);
nor U17256 (N_17256,N_16719,N_16900);
or U17257 (N_17257,N_16206,N_16388);
and U17258 (N_17258,N_16327,N_16569);
and U17259 (N_17259,N_16017,N_16687);
nor U17260 (N_17260,N_16662,N_16762);
nand U17261 (N_17261,N_16472,N_16643);
nor U17262 (N_17262,N_16212,N_16795);
xor U17263 (N_17263,N_16250,N_16823);
xor U17264 (N_17264,N_16521,N_16537);
nor U17265 (N_17265,N_16451,N_16992);
and U17266 (N_17266,N_16544,N_16223);
or U17267 (N_17267,N_16898,N_16157);
and U17268 (N_17268,N_16348,N_16905);
or U17269 (N_17269,N_16577,N_16960);
or U17270 (N_17270,N_16500,N_16964);
or U17271 (N_17271,N_16594,N_16970);
nand U17272 (N_17272,N_16000,N_16788);
and U17273 (N_17273,N_16241,N_16498);
or U17274 (N_17274,N_16149,N_16736);
nor U17275 (N_17275,N_16499,N_16785);
and U17276 (N_17276,N_16605,N_16727);
or U17277 (N_17277,N_16337,N_16891);
xnor U17278 (N_17278,N_16508,N_16249);
nor U17279 (N_17279,N_16542,N_16159);
nand U17280 (N_17280,N_16679,N_16774);
nor U17281 (N_17281,N_16802,N_16268);
nand U17282 (N_17282,N_16044,N_16071);
nand U17283 (N_17283,N_16886,N_16246);
or U17284 (N_17284,N_16546,N_16135);
or U17285 (N_17285,N_16731,N_16852);
or U17286 (N_17286,N_16586,N_16691);
nor U17287 (N_17287,N_16809,N_16434);
and U17288 (N_17288,N_16525,N_16644);
nor U17289 (N_17289,N_16402,N_16222);
nor U17290 (N_17290,N_16854,N_16636);
xor U17291 (N_17291,N_16730,N_16130);
and U17292 (N_17292,N_16496,N_16969);
nor U17293 (N_17293,N_16640,N_16776);
xnor U17294 (N_17294,N_16922,N_16773);
and U17295 (N_17295,N_16656,N_16888);
nor U17296 (N_17296,N_16015,N_16141);
xor U17297 (N_17297,N_16579,N_16218);
and U17298 (N_17298,N_16742,N_16978);
xnor U17299 (N_17299,N_16681,N_16032);
or U17300 (N_17300,N_16455,N_16894);
nor U17301 (N_17301,N_16966,N_16875);
xor U17302 (N_17302,N_16589,N_16081);
nand U17303 (N_17303,N_16102,N_16242);
xor U17304 (N_17304,N_16310,N_16313);
or U17305 (N_17305,N_16786,N_16770);
nor U17306 (N_17306,N_16623,N_16677);
nand U17307 (N_17307,N_16490,N_16238);
xnor U17308 (N_17308,N_16975,N_16165);
nand U17309 (N_17309,N_16827,N_16295);
xor U17310 (N_17310,N_16290,N_16361);
or U17311 (N_17311,N_16175,N_16177);
or U17312 (N_17312,N_16556,N_16751);
or U17313 (N_17313,N_16404,N_16581);
nor U17314 (N_17314,N_16349,N_16077);
xor U17315 (N_17315,N_16007,N_16562);
nor U17316 (N_17316,N_16555,N_16550);
nand U17317 (N_17317,N_16512,N_16436);
xnor U17318 (N_17318,N_16775,N_16354);
nand U17319 (N_17319,N_16106,N_16418);
and U17320 (N_17320,N_16477,N_16497);
nand U17321 (N_17321,N_16186,N_16688);
nand U17322 (N_17322,N_16754,N_16098);
and U17323 (N_17323,N_16720,N_16919);
xor U17324 (N_17324,N_16887,N_16033);
and U17325 (N_17325,N_16072,N_16692);
nand U17326 (N_17326,N_16503,N_16664);
and U17327 (N_17327,N_16088,N_16941);
xor U17328 (N_17328,N_16151,N_16557);
or U17329 (N_17329,N_16430,N_16021);
or U17330 (N_17330,N_16456,N_16373);
and U17331 (N_17331,N_16737,N_16458);
nor U17332 (N_17332,N_16008,N_16235);
and U17333 (N_17333,N_16767,N_16358);
or U17334 (N_17334,N_16437,N_16267);
and U17335 (N_17335,N_16890,N_16897);
and U17336 (N_17336,N_16315,N_16406);
nand U17337 (N_17337,N_16799,N_16634);
and U17338 (N_17338,N_16571,N_16880);
nand U17339 (N_17339,N_16972,N_16100);
and U17340 (N_17340,N_16866,N_16123);
and U17341 (N_17341,N_16573,N_16789);
nor U17342 (N_17342,N_16286,N_16127);
nand U17343 (N_17343,N_16930,N_16659);
xnor U17344 (N_17344,N_16723,N_16410);
nor U17345 (N_17345,N_16203,N_16296);
xor U17346 (N_17346,N_16851,N_16210);
xor U17347 (N_17347,N_16069,N_16872);
or U17348 (N_17348,N_16005,N_16395);
xnor U17349 (N_17349,N_16896,N_16915);
nor U17350 (N_17350,N_16952,N_16761);
nand U17351 (N_17351,N_16051,N_16208);
nand U17352 (N_17352,N_16837,N_16918);
xnor U17353 (N_17353,N_16467,N_16873);
xor U17354 (N_17354,N_16543,N_16863);
or U17355 (N_17355,N_16820,N_16096);
and U17356 (N_17356,N_16590,N_16625);
or U17357 (N_17357,N_16074,N_16488);
xor U17358 (N_17358,N_16184,N_16193);
nand U17359 (N_17359,N_16211,N_16302);
nor U17360 (N_17360,N_16412,N_16516);
nor U17361 (N_17361,N_16194,N_16239);
and U17362 (N_17362,N_16244,N_16763);
nand U17363 (N_17363,N_16445,N_16269);
and U17364 (N_17364,N_16615,N_16784);
xnor U17365 (N_17365,N_16189,N_16597);
xor U17366 (N_17366,N_16712,N_16216);
and U17367 (N_17367,N_16396,N_16086);
and U17368 (N_17368,N_16528,N_16908);
and U17369 (N_17369,N_16768,N_16911);
or U17370 (N_17370,N_16028,N_16227);
xor U17371 (N_17371,N_16025,N_16538);
or U17372 (N_17372,N_16152,N_16335);
xor U17373 (N_17373,N_16197,N_16139);
and U17374 (N_17374,N_16553,N_16066);
and U17375 (N_17375,N_16118,N_16814);
nor U17376 (N_17376,N_16938,N_16793);
or U17377 (N_17377,N_16578,N_16798);
xor U17378 (N_17378,N_16934,N_16381);
and U17379 (N_17379,N_16332,N_16217);
nand U17380 (N_17380,N_16043,N_16653);
xor U17381 (N_17381,N_16611,N_16603);
nor U17382 (N_17382,N_16288,N_16791);
nand U17383 (N_17383,N_16405,N_16002);
xnor U17384 (N_17384,N_16435,N_16001);
and U17385 (N_17385,N_16016,N_16811);
nand U17386 (N_17386,N_16155,N_16099);
nor U17387 (N_17387,N_16119,N_16617);
nor U17388 (N_17388,N_16980,N_16213);
nor U17389 (N_17389,N_16904,N_16642);
or U17390 (N_17390,N_16514,N_16331);
or U17391 (N_17391,N_16259,N_16716);
and U17392 (N_17392,N_16023,N_16271);
or U17393 (N_17393,N_16105,N_16350);
xor U17394 (N_17394,N_16826,N_16987);
nor U17395 (N_17395,N_16162,N_16299);
nor U17396 (N_17396,N_16094,N_16385);
nor U17397 (N_17397,N_16513,N_16264);
nand U17398 (N_17398,N_16580,N_16012);
and U17399 (N_17399,N_16963,N_16994);
and U17400 (N_17400,N_16124,N_16398);
nor U17401 (N_17401,N_16650,N_16382);
nand U17402 (N_17402,N_16026,N_16275);
or U17403 (N_17403,N_16718,N_16359);
xnor U17404 (N_17404,N_16883,N_16078);
and U17405 (N_17405,N_16515,N_16306);
xnor U17406 (N_17406,N_16778,N_16114);
nor U17407 (N_17407,N_16857,N_16076);
xnor U17408 (N_17408,N_16879,N_16087);
nor U17409 (N_17409,N_16721,N_16524);
xnor U17410 (N_17410,N_16733,N_16140);
nand U17411 (N_17411,N_16607,N_16663);
nor U17412 (N_17412,N_16554,N_16613);
and U17413 (N_17413,N_16722,N_16030);
xnor U17414 (N_17414,N_16568,N_16750);
nand U17415 (N_17415,N_16757,N_16672);
and U17416 (N_17416,N_16370,N_16953);
nand U17417 (N_17417,N_16079,N_16610);
xnor U17418 (N_17418,N_16236,N_16801);
nor U17419 (N_17419,N_16423,N_16842);
or U17420 (N_17420,N_16224,N_16665);
or U17421 (N_17421,N_16276,N_16125);
and U17422 (N_17422,N_16004,N_16429);
and U17423 (N_17423,N_16759,N_16220);
or U17424 (N_17424,N_16899,N_16117);
and U17425 (N_17425,N_16849,N_16095);
or U17426 (N_17426,N_16545,N_16255);
or U17427 (N_17427,N_16446,N_16325);
and U17428 (N_17428,N_16753,N_16684);
and U17429 (N_17429,N_16230,N_16877);
nor U17430 (N_17430,N_16104,N_16304);
and U17431 (N_17431,N_16231,N_16882);
and U17432 (N_17432,N_16160,N_16336);
nand U17433 (N_17433,N_16522,N_16226);
nand U17434 (N_17434,N_16925,N_16257);
nor U17435 (N_17435,N_16710,N_16126);
and U17436 (N_17436,N_16867,N_16532);
or U17437 (N_17437,N_16933,N_16360);
nand U17438 (N_17438,N_16053,N_16453);
or U17439 (N_17439,N_16819,N_16620);
nand U17440 (N_17440,N_16277,N_16447);
or U17441 (N_17441,N_16228,N_16871);
or U17442 (N_17442,N_16835,N_16256);
or U17443 (N_17443,N_16063,N_16540);
nor U17444 (N_17444,N_16726,N_16967);
or U17445 (N_17445,N_16923,N_16864);
and U17446 (N_17446,N_16629,N_16363);
nor U17447 (N_17447,N_16427,N_16154);
and U17448 (N_17448,N_16190,N_16411);
xor U17449 (N_17449,N_16777,N_16570);
and U17450 (N_17450,N_16604,N_16847);
and U17451 (N_17451,N_16300,N_16661);
xnor U17452 (N_17452,N_16993,N_16633);
xnor U17453 (N_17453,N_16917,N_16817);
xor U17454 (N_17454,N_16283,N_16156);
or U17455 (N_17455,N_16670,N_16654);
nor U17456 (N_17456,N_16171,N_16539);
nand U17457 (N_17457,N_16413,N_16651);
xnor U17458 (N_17458,N_16219,N_16667);
xor U17459 (N_17459,N_16701,N_16330);
and U17460 (N_17460,N_16438,N_16530);
xor U17461 (N_17461,N_16416,N_16825);
nor U17462 (N_17462,N_16807,N_16116);
xor U17463 (N_17463,N_16598,N_16031);
nor U17464 (N_17464,N_16389,N_16870);
nor U17465 (N_17465,N_16432,N_16504);
nor U17466 (N_17466,N_16806,N_16073);
xor U17467 (N_17467,N_16956,N_16054);
xor U17468 (N_17468,N_16764,N_16609);
nand U17469 (N_17469,N_16986,N_16366);
nand U17470 (N_17470,N_16572,N_16507);
xor U17471 (N_17471,N_16853,N_16655);
xnor U17472 (N_17472,N_16705,N_16383);
nand U17473 (N_17473,N_16526,N_16176);
nand U17474 (N_17474,N_16465,N_16040);
nor U17475 (N_17475,N_16356,N_16517);
xor U17476 (N_17476,N_16057,N_16971);
nand U17477 (N_17477,N_16207,N_16022);
or U17478 (N_17478,N_16558,N_16347);
and U17479 (N_17479,N_16561,N_16333);
nand U17480 (N_17480,N_16309,N_16464);
nor U17481 (N_17481,N_16831,N_16989);
nor U17482 (N_17482,N_16614,N_16856);
xnor U17483 (N_17483,N_16303,N_16948);
nand U17484 (N_17484,N_16196,N_16816);
or U17485 (N_17485,N_16251,N_16170);
nand U17486 (N_17486,N_16181,N_16475);
xnor U17487 (N_17487,N_16658,N_16045);
or U17488 (N_17488,N_16783,N_16997);
xor U17489 (N_17489,N_16248,N_16101);
or U17490 (N_17490,N_16547,N_16861);
nor U17491 (N_17491,N_16673,N_16977);
or U17492 (N_17492,N_16841,N_16965);
nor U17493 (N_17493,N_16487,N_16961);
or U17494 (N_17494,N_16440,N_16187);
or U17495 (N_17495,N_16260,N_16901);
or U17496 (N_17496,N_16390,N_16493);
or U17497 (N_17497,N_16729,N_16703);
or U17498 (N_17498,N_16384,N_16981);
nor U17499 (N_17499,N_16014,N_16024);
and U17500 (N_17500,N_16047,N_16964);
nand U17501 (N_17501,N_16706,N_16265);
or U17502 (N_17502,N_16821,N_16391);
nand U17503 (N_17503,N_16115,N_16420);
nor U17504 (N_17504,N_16507,N_16191);
and U17505 (N_17505,N_16590,N_16637);
nor U17506 (N_17506,N_16364,N_16416);
and U17507 (N_17507,N_16215,N_16087);
nand U17508 (N_17508,N_16268,N_16535);
and U17509 (N_17509,N_16385,N_16947);
and U17510 (N_17510,N_16344,N_16835);
or U17511 (N_17511,N_16946,N_16796);
nand U17512 (N_17512,N_16311,N_16249);
or U17513 (N_17513,N_16004,N_16912);
xnor U17514 (N_17514,N_16321,N_16977);
or U17515 (N_17515,N_16246,N_16311);
nand U17516 (N_17516,N_16966,N_16448);
or U17517 (N_17517,N_16932,N_16230);
and U17518 (N_17518,N_16040,N_16323);
nor U17519 (N_17519,N_16420,N_16501);
xnor U17520 (N_17520,N_16568,N_16033);
and U17521 (N_17521,N_16316,N_16856);
nor U17522 (N_17522,N_16665,N_16604);
xnor U17523 (N_17523,N_16675,N_16202);
or U17524 (N_17524,N_16369,N_16562);
nor U17525 (N_17525,N_16116,N_16218);
nand U17526 (N_17526,N_16687,N_16397);
nor U17527 (N_17527,N_16516,N_16376);
nand U17528 (N_17528,N_16081,N_16473);
and U17529 (N_17529,N_16770,N_16620);
nor U17530 (N_17530,N_16825,N_16133);
and U17531 (N_17531,N_16065,N_16006);
xor U17532 (N_17532,N_16427,N_16179);
or U17533 (N_17533,N_16654,N_16882);
nor U17534 (N_17534,N_16858,N_16608);
nand U17535 (N_17535,N_16407,N_16450);
and U17536 (N_17536,N_16784,N_16600);
xnor U17537 (N_17537,N_16932,N_16274);
or U17538 (N_17538,N_16218,N_16727);
xnor U17539 (N_17539,N_16721,N_16257);
xnor U17540 (N_17540,N_16324,N_16818);
nand U17541 (N_17541,N_16807,N_16297);
and U17542 (N_17542,N_16755,N_16339);
or U17543 (N_17543,N_16197,N_16797);
and U17544 (N_17544,N_16011,N_16784);
nor U17545 (N_17545,N_16950,N_16012);
nor U17546 (N_17546,N_16400,N_16430);
nor U17547 (N_17547,N_16052,N_16578);
nand U17548 (N_17548,N_16741,N_16817);
or U17549 (N_17549,N_16931,N_16187);
and U17550 (N_17550,N_16221,N_16455);
and U17551 (N_17551,N_16712,N_16948);
or U17552 (N_17552,N_16181,N_16876);
nand U17553 (N_17553,N_16503,N_16254);
or U17554 (N_17554,N_16604,N_16689);
nor U17555 (N_17555,N_16968,N_16603);
or U17556 (N_17556,N_16103,N_16467);
nand U17557 (N_17557,N_16461,N_16454);
nor U17558 (N_17558,N_16653,N_16262);
xor U17559 (N_17559,N_16199,N_16477);
and U17560 (N_17560,N_16773,N_16674);
nor U17561 (N_17561,N_16704,N_16168);
nor U17562 (N_17562,N_16647,N_16308);
and U17563 (N_17563,N_16974,N_16303);
and U17564 (N_17564,N_16118,N_16736);
and U17565 (N_17565,N_16510,N_16026);
or U17566 (N_17566,N_16115,N_16606);
and U17567 (N_17567,N_16234,N_16534);
and U17568 (N_17568,N_16671,N_16041);
nor U17569 (N_17569,N_16419,N_16342);
or U17570 (N_17570,N_16365,N_16450);
nand U17571 (N_17571,N_16514,N_16210);
nand U17572 (N_17572,N_16633,N_16658);
nor U17573 (N_17573,N_16711,N_16180);
and U17574 (N_17574,N_16959,N_16960);
and U17575 (N_17575,N_16636,N_16449);
nand U17576 (N_17576,N_16855,N_16827);
xnor U17577 (N_17577,N_16428,N_16241);
and U17578 (N_17578,N_16259,N_16781);
xor U17579 (N_17579,N_16563,N_16313);
nand U17580 (N_17580,N_16287,N_16369);
and U17581 (N_17581,N_16753,N_16852);
or U17582 (N_17582,N_16002,N_16437);
nor U17583 (N_17583,N_16200,N_16316);
nand U17584 (N_17584,N_16848,N_16351);
xnor U17585 (N_17585,N_16281,N_16272);
and U17586 (N_17586,N_16853,N_16693);
nand U17587 (N_17587,N_16895,N_16223);
and U17588 (N_17588,N_16987,N_16290);
and U17589 (N_17589,N_16486,N_16419);
nor U17590 (N_17590,N_16897,N_16977);
xnor U17591 (N_17591,N_16310,N_16998);
and U17592 (N_17592,N_16694,N_16203);
xor U17593 (N_17593,N_16646,N_16725);
or U17594 (N_17594,N_16628,N_16804);
or U17595 (N_17595,N_16179,N_16301);
xnor U17596 (N_17596,N_16745,N_16338);
or U17597 (N_17597,N_16256,N_16881);
nor U17598 (N_17598,N_16012,N_16186);
xnor U17599 (N_17599,N_16076,N_16386);
xnor U17600 (N_17600,N_16973,N_16757);
nand U17601 (N_17601,N_16093,N_16867);
and U17602 (N_17602,N_16077,N_16435);
xnor U17603 (N_17603,N_16897,N_16654);
xnor U17604 (N_17604,N_16517,N_16602);
or U17605 (N_17605,N_16665,N_16021);
and U17606 (N_17606,N_16155,N_16273);
nand U17607 (N_17607,N_16942,N_16083);
nor U17608 (N_17608,N_16867,N_16785);
or U17609 (N_17609,N_16985,N_16762);
and U17610 (N_17610,N_16149,N_16486);
nand U17611 (N_17611,N_16302,N_16748);
and U17612 (N_17612,N_16725,N_16674);
nor U17613 (N_17613,N_16482,N_16136);
nand U17614 (N_17614,N_16523,N_16715);
and U17615 (N_17615,N_16155,N_16950);
nor U17616 (N_17616,N_16460,N_16575);
xor U17617 (N_17617,N_16964,N_16562);
nand U17618 (N_17618,N_16014,N_16754);
and U17619 (N_17619,N_16030,N_16444);
nor U17620 (N_17620,N_16602,N_16700);
nor U17621 (N_17621,N_16519,N_16961);
nor U17622 (N_17622,N_16484,N_16133);
or U17623 (N_17623,N_16727,N_16638);
nand U17624 (N_17624,N_16192,N_16351);
xnor U17625 (N_17625,N_16136,N_16706);
xor U17626 (N_17626,N_16134,N_16599);
nand U17627 (N_17627,N_16952,N_16189);
nand U17628 (N_17628,N_16900,N_16559);
or U17629 (N_17629,N_16497,N_16857);
nand U17630 (N_17630,N_16479,N_16159);
nor U17631 (N_17631,N_16491,N_16765);
nor U17632 (N_17632,N_16432,N_16309);
or U17633 (N_17633,N_16715,N_16732);
and U17634 (N_17634,N_16954,N_16185);
xor U17635 (N_17635,N_16502,N_16370);
nand U17636 (N_17636,N_16247,N_16005);
nor U17637 (N_17637,N_16271,N_16727);
nor U17638 (N_17638,N_16004,N_16778);
or U17639 (N_17639,N_16025,N_16568);
xor U17640 (N_17640,N_16450,N_16210);
nor U17641 (N_17641,N_16967,N_16786);
xnor U17642 (N_17642,N_16950,N_16476);
nand U17643 (N_17643,N_16191,N_16406);
nand U17644 (N_17644,N_16283,N_16770);
and U17645 (N_17645,N_16300,N_16623);
and U17646 (N_17646,N_16535,N_16431);
and U17647 (N_17647,N_16694,N_16351);
or U17648 (N_17648,N_16603,N_16019);
and U17649 (N_17649,N_16138,N_16023);
nor U17650 (N_17650,N_16097,N_16892);
xor U17651 (N_17651,N_16154,N_16679);
nand U17652 (N_17652,N_16715,N_16624);
xor U17653 (N_17653,N_16074,N_16955);
xnor U17654 (N_17654,N_16662,N_16219);
or U17655 (N_17655,N_16419,N_16059);
xor U17656 (N_17656,N_16218,N_16383);
or U17657 (N_17657,N_16180,N_16155);
or U17658 (N_17658,N_16767,N_16059);
nor U17659 (N_17659,N_16219,N_16926);
xor U17660 (N_17660,N_16127,N_16437);
nand U17661 (N_17661,N_16730,N_16761);
or U17662 (N_17662,N_16145,N_16318);
xnor U17663 (N_17663,N_16426,N_16779);
xnor U17664 (N_17664,N_16832,N_16814);
xor U17665 (N_17665,N_16187,N_16293);
nand U17666 (N_17666,N_16325,N_16303);
and U17667 (N_17667,N_16229,N_16581);
xor U17668 (N_17668,N_16955,N_16245);
nor U17669 (N_17669,N_16702,N_16226);
nand U17670 (N_17670,N_16350,N_16575);
nand U17671 (N_17671,N_16891,N_16276);
and U17672 (N_17672,N_16504,N_16204);
nor U17673 (N_17673,N_16471,N_16415);
and U17674 (N_17674,N_16062,N_16276);
and U17675 (N_17675,N_16824,N_16022);
nor U17676 (N_17676,N_16236,N_16972);
nor U17677 (N_17677,N_16306,N_16709);
nor U17678 (N_17678,N_16580,N_16797);
or U17679 (N_17679,N_16694,N_16440);
and U17680 (N_17680,N_16318,N_16532);
and U17681 (N_17681,N_16809,N_16739);
or U17682 (N_17682,N_16872,N_16112);
xor U17683 (N_17683,N_16613,N_16324);
xnor U17684 (N_17684,N_16810,N_16584);
nand U17685 (N_17685,N_16231,N_16349);
and U17686 (N_17686,N_16235,N_16153);
nand U17687 (N_17687,N_16127,N_16362);
nor U17688 (N_17688,N_16747,N_16160);
and U17689 (N_17689,N_16920,N_16304);
nor U17690 (N_17690,N_16189,N_16031);
or U17691 (N_17691,N_16114,N_16171);
nand U17692 (N_17692,N_16453,N_16121);
nor U17693 (N_17693,N_16371,N_16657);
and U17694 (N_17694,N_16067,N_16589);
or U17695 (N_17695,N_16451,N_16840);
xor U17696 (N_17696,N_16609,N_16386);
and U17697 (N_17697,N_16147,N_16976);
and U17698 (N_17698,N_16093,N_16680);
nor U17699 (N_17699,N_16467,N_16768);
xnor U17700 (N_17700,N_16650,N_16155);
or U17701 (N_17701,N_16086,N_16775);
xnor U17702 (N_17702,N_16896,N_16904);
and U17703 (N_17703,N_16150,N_16219);
or U17704 (N_17704,N_16569,N_16177);
nor U17705 (N_17705,N_16071,N_16876);
or U17706 (N_17706,N_16497,N_16827);
or U17707 (N_17707,N_16145,N_16402);
and U17708 (N_17708,N_16723,N_16936);
or U17709 (N_17709,N_16814,N_16442);
or U17710 (N_17710,N_16174,N_16326);
or U17711 (N_17711,N_16063,N_16827);
nor U17712 (N_17712,N_16308,N_16573);
and U17713 (N_17713,N_16507,N_16349);
nand U17714 (N_17714,N_16027,N_16817);
nand U17715 (N_17715,N_16392,N_16261);
and U17716 (N_17716,N_16123,N_16331);
and U17717 (N_17717,N_16071,N_16843);
xnor U17718 (N_17718,N_16682,N_16843);
and U17719 (N_17719,N_16298,N_16890);
and U17720 (N_17720,N_16352,N_16980);
xor U17721 (N_17721,N_16130,N_16004);
xor U17722 (N_17722,N_16301,N_16048);
nand U17723 (N_17723,N_16082,N_16689);
xnor U17724 (N_17724,N_16391,N_16697);
xnor U17725 (N_17725,N_16988,N_16187);
nand U17726 (N_17726,N_16139,N_16259);
xor U17727 (N_17727,N_16713,N_16543);
xnor U17728 (N_17728,N_16623,N_16617);
nand U17729 (N_17729,N_16536,N_16486);
nand U17730 (N_17730,N_16812,N_16199);
xor U17731 (N_17731,N_16274,N_16540);
or U17732 (N_17732,N_16038,N_16341);
nor U17733 (N_17733,N_16847,N_16162);
or U17734 (N_17734,N_16793,N_16313);
xnor U17735 (N_17735,N_16649,N_16062);
nor U17736 (N_17736,N_16170,N_16031);
nor U17737 (N_17737,N_16663,N_16727);
nor U17738 (N_17738,N_16198,N_16438);
nand U17739 (N_17739,N_16468,N_16109);
and U17740 (N_17740,N_16050,N_16545);
or U17741 (N_17741,N_16643,N_16334);
nor U17742 (N_17742,N_16442,N_16911);
nand U17743 (N_17743,N_16391,N_16439);
xnor U17744 (N_17744,N_16066,N_16983);
and U17745 (N_17745,N_16847,N_16614);
and U17746 (N_17746,N_16678,N_16496);
xnor U17747 (N_17747,N_16966,N_16243);
xor U17748 (N_17748,N_16977,N_16117);
and U17749 (N_17749,N_16625,N_16546);
nor U17750 (N_17750,N_16293,N_16784);
nor U17751 (N_17751,N_16629,N_16763);
nor U17752 (N_17752,N_16798,N_16779);
and U17753 (N_17753,N_16681,N_16328);
xor U17754 (N_17754,N_16199,N_16226);
nand U17755 (N_17755,N_16520,N_16455);
nor U17756 (N_17756,N_16161,N_16552);
xor U17757 (N_17757,N_16680,N_16061);
or U17758 (N_17758,N_16477,N_16336);
xnor U17759 (N_17759,N_16271,N_16096);
and U17760 (N_17760,N_16327,N_16643);
and U17761 (N_17761,N_16732,N_16432);
xnor U17762 (N_17762,N_16586,N_16861);
or U17763 (N_17763,N_16929,N_16946);
nor U17764 (N_17764,N_16049,N_16754);
xnor U17765 (N_17765,N_16499,N_16648);
or U17766 (N_17766,N_16036,N_16258);
xnor U17767 (N_17767,N_16584,N_16946);
nor U17768 (N_17768,N_16008,N_16993);
nand U17769 (N_17769,N_16890,N_16218);
or U17770 (N_17770,N_16766,N_16119);
and U17771 (N_17771,N_16878,N_16308);
nand U17772 (N_17772,N_16571,N_16997);
or U17773 (N_17773,N_16303,N_16644);
xnor U17774 (N_17774,N_16729,N_16001);
nor U17775 (N_17775,N_16699,N_16341);
or U17776 (N_17776,N_16827,N_16528);
xor U17777 (N_17777,N_16996,N_16869);
or U17778 (N_17778,N_16554,N_16970);
and U17779 (N_17779,N_16441,N_16935);
or U17780 (N_17780,N_16591,N_16486);
and U17781 (N_17781,N_16095,N_16226);
nand U17782 (N_17782,N_16578,N_16178);
nor U17783 (N_17783,N_16950,N_16152);
nor U17784 (N_17784,N_16955,N_16674);
and U17785 (N_17785,N_16021,N_16831);
or U17786 (N_17786,N_16390,N_16003);
and U17787 (N_17787,N_16441,N_16967);
nor U17788 (N_17788,N_16725,N_16994);
nand U17789 (N_17789,N_16546,N_16027);
or U17790 (N_17790,N_16806,N_16045);
nand U17791 (N_17791,N_16546,N_16488);
xor U17792 (N_17792,N_16244,N_16938);
nand U17793 (N_17793,N_16465,N_16755);
nor U17794 (N_17794,N_16607,N_16317);
and U17795 (N_17795,N_16721,N_16629);
nand U17796 (N_17796,N_16543,N_16963);
nor U17797 (N_17797,N_16880,N_16096);
and U17798 (N_17798,N_16712,N_16908);
xnor U17799 (N_17799,N_16696,N_16259);
nor U17800 (N_17800,N_16876,N_16800);
and U17801 (N_17801,N_16342,N_16734);
and U17802 (N_17802,N_16742,N_16088);
nand U17803 (N_17803,N_16537,N_16710);
and U17804 (N_17804,N_16779,N_16410);
nand U17805 (N_17805,N_16976,N_16241);
xor U17806 (N_17806,N_16320,N_16899);
nand U17807 (N_17807,N_16973,N_16321);
nand U17808 (N_17808,N_16322,N_16331);
or U17809 (N_17809,N_16759,N_16437);
or U17810 (N_17810,N_16593,N_16185);
and U17811 (N_17811,N_16330,N_16210);
xor U17812 (N_17812,N_16927,N_16176);
xor U17813 (N_17813,N_16666,N_16562);
and U17814 (N_17814,N_16718,N_16371);
and U17815 (N_17815,N_16898,N_16160);
nor U17816 (N_17816,N_16682,N_16130);
or U17817 (N_17817,N_16619,N_16189);
or U17818 (N_17818,N_16247,N_16346);
nand U17819 (N_17819,N_16857,N_16678);
nand U17820 (N_17820,N_16397,N_16768);
nor U17821 (N_17821,N_16503,N_16316);
nand U17822 (N_17822,N_16738,N_16514);
and U17823 (N_17823,N_16931,N_16606);
and U17824 (N_17824,N_16395,N_16364);
nand U17825 (N_17825,N_16680,N_16183);
xnor U17826 (N_17826,N_16007,N_16611);
and U17827 (N_17827,N_16105,N_16000);
nor U17828 (N_17828,N_16308,N_16336);
nor U17829 (N_17829,N_16645,N_16740);
xor U17830 (N_17830,N_16254,N_16788);
xor U17831 (N_17831,N_16973,N_16056);
nand U17832 (N_17832,N_16792,N_16837);
and U17833 (N_17833,N_16252,N_16196);
or U17834 (N_17834,N_16166,N_16874);
and U17835 (N_17835,N_16812,N_16698);
nor U17836 (N_17836,N_16303,N_16552);
xnor U17837 (N_17837,N_16418,N_16416);
nor U17838 (N_17838,N_16500,N_16958);
xnor U17839 (N_17839,N_16956,N_16024);
nor U17840 (N_17840,N_16047,N_16990);
and U17841 (N_17841,N_16957,N_16037);
xor U17842 (N_17842,N_16854,N_16236);
and U17843 (N_17843,N_16379,N_16540);
nand U17844 (N_17844,N_16652,N_16813);
and U17845 (N_17845,N_16796,N_16199);
xnor U17846 (N_17846,N_16241,N_16728);
or U17847 (N_17847,N_16019,N_16911);
nor U17848 (N_17848,N_16638,N_16656);
or U17849 (N_17849,N_16837,N_16461);
xor U17850 (N_17850,N_16699,N_16701);
nand U17851 (N_17851,N_16388,N_16168);
xnor U17852 (N_17852,N_16941,N_16484);
nand U17853 (N_17853,N_16363,N_16355);
and U17854 (N_17854,N_16517,N_16665);
nor U17855 (N_17855,N_16700,N_16568);
nor U17856 (N_17856,N_16591,N_16916);
and U17857 (N_17857,N_16919,N_16534);
xor U17858 (N_17858,N_16323,N_16592);
and U17859 (N_17859,N_16020,N_16763);
or U17860 (N_17860,N_16213,N_16412);
or U17861 (N_17861,N_16696,N_16124);
and U17862 (N_17862,N_16824,N_16436);
or U17863 (N_17863,N_16825,N_16236);
and U17864 (N_17864,N_16713,N_16201);
or U17865 (N_17865,N_16759,N_16853);
or U17866 (N_17866,N_16533,N_16925);
nand U17867 (N_17867,N_16566,N_16269);
nor U17868 (N_17868,N_16769,N_16966);
xnor U17869 (N_17869,N_16571,N_16916);
nor U17870 (N_17870,N_16241,N_16448);
or U17871 (N_17871,N_16173,N_16289);
and U17872 (N_17872,N_16031,N_16382);
xnor U17873 (N_17873,N_16981,N_16650);
nand U17874 (N_17874,N_16558,N_16197);
and U17875 (N_17875,N_16450,N_16161);
and U17876 (N_17876,N_16542,N_16193);
or U17877 (N_17877,N_16573,N_16377);
nor U17878 (N_17878,N_16636,N_16204);
and U17879 (N_17879,N_16407,N_16879);
nand U17880 (N_17880,N_16863,N_16817);
nor U17881 (N_17881,N_16065,N_16132);
or U17882 (N_17882,N_16696,N_16163);
or U17883 (N_17883,N_16136,N_16073);
xor U17884 (N_17884,N_16404,N_16183);
nor U17885 (N_17885,N_16276,N_16380);
and U17886 (N_17886,N_16036,N_16926);
xor U17887 (N_17887,N_16000,N_16655);
or U17888 (N_17888,N_16503,N_16598);
nor U17889 (N_17889,N_16177,N_16304);
or U17890 (N_17890,N_16142,N_16202);
or U17891 (N_17891,N_16770,N_16551);
xor U17892 (N_17892,N_16594,N_16959);
nand U17893 (N_17893,N_16815,N_16358);
or U17894 (N_17894,N_16478,N_16073);
nand U17895 (N_17895,N_16164,N_16890);
nand U17896 (N_17896,N_16543,N_16748);
or U17897 (N_17897,N_16119,N_16435);
or U17898 (N_17898,N_16270,N_16026);
xor U17899 (N_17899,N_16022,N_16394);
xor U17900 (N_17900,N_16632,N_16467);
or U17901 (N_17901,N_16564,N_16217);
nor U17902 (N_17902,N_16844,N_16417);
and U17903 (N_17903,N_16759,N_16186);
nand U17904 (N_17904,N_16910,N_16471);
nand U17905 (N_17905,N_16723,N_16010);
xor U17906 (N_17906,N_16280,N_16334);
or U17907 (N_17907,N_16812,N_16445);
xor U17908 (N_17908,N_16653,N_16346);
nor U17909 (N_17909,N_16587,N_16236);
xor U17910 (N_17910,N_16738,N_16208);
nor U17911 (N_17911,N_16761,N_16728);
nor U17912 (N_17912,N_16981,N_16799);
nand U17913 (N_17913,N_16022,N_16836);
nor U17914 (N_17914,N_16462,N_16551);
or U17915 (N_17915,N_16178,N_16918);
nand U17916 (N_17916,N_16881,N_16165);
and U17917 (N_17917,N_16941,N_16657);
nor U17918 (N_17918,N_16874,N_16003);
nand U17919 (N_17919,N_16843,N_16100);
and U17920 (N_17920,N_16925,N_16787);
or U17921 (N_17921,N_16163,N_16572);
nor U17922 (N_17922,N_16992,N_16444);
or U17923 (N_17923,N_16272,N_16560);
and U17924 (N_17924,N_16745,N_16690);
nor U17925 (N_17925,N_16308,N_16637);
or U17926 (N_17926,N_16332,N_16492);
nand U17927 (N_17927,N_16171,N_16061);
nor U17928 (N_17928,N_16203,N_16576);
or U17929 (N_17929,N_16781,N_16748);
nor U17930 (N_17930,N_16865,N_16207);
nand U17931 (N_17931,N_16291,N_16623);
xnor U17932 (N_17932,N_16307,N_16476);
nand U17933 (N_17933,N_16200,N_16800);
and U17934 (N_17934,N_16322,N_16884);
or U17935 (N_17935,N_16574,N_16306);
nor U17936 (N_17936,N_16056,N_16142);
nor U17937 (N_17937,N_16609,N_16781);
or U17938 (N_17938,N_16702,N_16727);
nor U17939 (N_17939,N_16115,N_16464);
nand U17940 (N_17940,N_16638,N_16213);
and U17941 (N_17941,N_16040,N_16887);
or U17942 (N_17942,N_16007,N_16982);
and U17943 (N_17943,N_16959,N_16461);
nor U17944 (N_17944,N_16976,N_16354);
xor U17945 (N_17945,N_16817,N_16226);
nand U17946 (N_17946,N_16806,N_16564);
and U17947 (N_17947,N_16814,N_16502);
xnor U17948 (N_17948,N_16846,N_16035);
or U17949 (N_17949,N_16928,N_16634);
and U17950 (N_17950,N_16224,N_16670);
nor U17951 (N_17951,N_16165,N_16475);
and U17952 (N_17952,N_16265,N_16677);
and U17953 (N_17953,N_16769,N_16346);
nor U17954 (N_17954,N_16843,N_16752);
and U17955 (N_17955,N_16816,N_16571);
or U17956 (N_17956,N_16075,N_16479);
nand U17957 (N_17957,N_16795,N_16179);
or U17958 (N_17958,N_16699,N_16320);
nand U17959 (N_17959,N_16344,N_16440);
and U17960 (N_17960,N_16486,N_16053);
or U17961 (N_17961,N_16915,N_16626);
xnor U17962 (N_17962,N_16333,N_16570);
or U17963 (N_17963,N_16112,N_16167);
nand U17964 (N_17964,N_16670,N_16990);
or U17965 (N_17965,N_16110,N_16806);
or U17966 (N_17966,N_16421,N_16234);
or U17967 (N_17967,N_16765,N_16749);
or U17968 (N_17968,N_16768,N_16159);
or U17969 (N_17969,N_16648,N_16704);
xnor U17970 (N_17970,N_16369,N_16607);
and U17971 (N_17971,N_16139,N_16880);
and U17972 (N_17972,N_16796,N_16735);
or U17973 (N_17973,N_16987,N_16208);
nand U17974 (N_17974,N_16335,N_16291);
xnor U17975 (N_17975,N_16205,N_16860);
nand U17976 (N_17976,N_16480,N_16946);
xor U17977 (N_17977,N_16412,N_16900);
nor U17978 (N_17978,N_16042,N_16952);
nand U17979 (N_17979,N_16224,N_16646);
xor U17980 (N_17980,N_16580,N_16767);
nor U17981 (N_17981,N_16051,N_16744);
nand U17982 (N_17982,N_16767,N_16016);
and U17983 (N_17983,N_16805,N_16900);
nor U17984 (N_17984,N_16435,N_16393);
nand U17985 (N_17985,N_16668,N_16644);
and U17986 (N_17986,N_16042,N_16423);
or U17987 (N_17987,N_16744,N_16328);
and U17988 (N_17988,N_16721,N_16728);
xor U17989 (N_17989,N_16597,N_16747);
or U17990 (N_17990,N_16471,N_16845);
nor U17991 (N_17991,N_16991,N_16453);
xnor U17992 (N_17992,N_16583,N_16754);
and U17993 (N_17993,N_16825,N_16918);
or U17994 (N_17994,N_16373,N_16881);
or U17995 (N_17995,N_16847,N_16942);
or U17996 (N_17996,N_16587,N_16079);
nor U17997 (N_17997,N_16469,N_16026);
and U17998 (N_17998,N_16811,N_16444);
and U17999 (N_17999,N_16603,N_16701);
and U18000 (N_18000,N_17325,N_17338);
nor U18001 (N_18001,N_17679,N_17908);
and U18002 (N_18002,N_17083,N_17410);
nor U18003 (N_18003,N_17375,N_17824);
xnor U18004 (N_18004,N_17466,N_17765);
and U18005 (N_18005,N_17712,N_17825);
and U18006 (N_18006,N_17512,N_17427);
or U18007 (N_18007,N_17799,N_17472);
nor U18008 (N_18008,N_17389,N_17626);
nor U18009 (N_18009,N_17571,N_17729);
xor U18010 (N_18010,N_17659,N_17148);
or U18011 (N_18011,N_17110,N_17182);
nor U18012 (N_18012,N_17502,N_17282);
nor U18013 (N_18013,N_17412,N_17280);
nor U18014 (N_18014,N_17175,N_17085);
or U18015 (N_18015,N_17969,N_17257);
nand U18016 (N_18016,N_17040,N_17095);
or U18017 (N_18017,N_17009,N_17832);
and U18018 (N_18018,N_17483,N_17658);
xor U18019 (N_18019,N_17887,N_17865);
or U18020 (N_18020,N_17408,N_17178);
nand U18021 (N_18021,N_17437,N_17365);
nand U18022 (N_18022,N_17344,N_17761);
nor U18023 (N_18023,N_17164,N_17743);
and U18024 (N_18024,N_17407,N_17147);
and U18025 (N_18025,N_17060,N_17414);
and U18026 (N_18026,N_17478,N_17168);
or U18027 (N_18027,N_17254,N_17318);
or U18028 (N_18028,N_17284,N_17634);
and U18029 (N_18029,N_17620,N_17805);
or U18030 (N_18030,N_17114,N_17721);
or U18031 (N_18031,N_17666,N_17103);
xor U18032 (N_18032,N_17736,N_17686);
or U18033 (N_18033,N_17079,N_17874);
nor U18034 (N_18034,N_17584,N_17443);
or U18035 (N_18035,N_17004,N_17102);
xnor U18036 (N_18036,N_17923,N_17803);
and U18037 (N_18037,N_17812,N_17193);
nand U18038 (N_18038,N_17610,N_17156);
or U18039 (N_18039,N_17189,N_17059);
or U18040 (N_18040,N_17081,N_17920);
nand U18041 (N_18041,N_17810,N_17546);
nand U18042 (N_18042,N_17678,N_17046);
and U18043 (N_18043,N_17248,N_17903);
nor U18044 (N_18044,N_17073,N_17696);
nand U18045 (N_18045,N_17202,N_17816);
and U18046 (N_18046,N_17861,N_17566);
nand U18047 (N_18047,N_17401,N_17646);
nor U18048 (N_18048,N_17235,N_17632);
nand U18049 (N_18049,N_17115,N_17575);
nor U18050 (N_18050,N_17195,N_17953);
or U18051 (N_18051,N_17654,N_17904);
and U18052 (N_18052,N_17531,N_17432);
or U18053 (N_18053,N_17460,N_17776);
xor U18054 (N_18054,N_17902,N_17053);
nor U18055 (N_18055,N_17197,N_17532);
xnor U18056 (N_18056,N_17932,N_17064);
nand U18057 (N_18057,N_17767,N_17315);
xnor U18058 (N_18058,N_17804,N_17356);
nand U18059 (N_18059,N_17017,N_17467);
nor U18060 (N_18060,N_17553,N_17304);
and U18061 (N_18061,N_17265,N_17368);
nor U18062 (N_18062,N_17281,N_17688);
nor U18063 (N_18063,N_17582,N_17151);
xor U18064 (N_18064,N_17405,N_17998);
nor U18065 (N_18065,N_17723,N_17455);
and U18066 (N_18066,N_17770,N_17070);
nor U18067 (N_18067,N_17409,N_17504);
nor U18068 (N_18068,N_17612,N_17627);
xnor U18069 (N_18069,N_17314,N_17153);
and U18070 (N_18070,N_17897,N_17594);
nand U18071 (N_18071,N_17676,N_17527);
nor U18072 (N_18072,N_17041,N_17087);
nand U18073 (N_18073,N_17837,N_17436);
and U18074 (N_18074,N_17888,N_17433);
or U18075 (N_18075,N_17749,N_17690);
and U18076 (N_18076,N_17541,N_17851);
or U18077 (N_18077,N_17668,N_17786);
xor U18078 (N_18078,N_17801,N_17977);
nor U18079 (N_18079,N_17909,N_17732);
xor U18080 (N_18080,N_17373,N_17342);
and U18081 (N_18081,N_17878,N_17753);
or U18082 (N_18082,N_17976,N_17458);
or U18083 (N_18083,N_17914,N_17072);
nor U18084 (N_18084,N_17973,N_17683);
or U18085 (N_18085,N_17277,N_17781);
or U18086 (N_18086,N_17317,N_17449);
nor U18087 (N_18087,N_17430,N_17827);
nand U18088 (N_18088,N_17341,N_17636);
nand U18089 (N_18089,N_17294,N_17003);
nand U18090 (N_18090,N_17336,N_17955);
nor U18091 (N_18091,N_17382,N_17497);
or U18092 (N_18092,N_17561,N_17345);
nand U18093 (N_18093,N_17881,N_17489);
xor U18094 (N_18094,N_17928,N_17623);
nand U18095 (N_18095,N_17031,N_17901);
xor U18096 (N_18096,N_17844,N_17350);
nand U18097 (N_18097,N_17943,N_17196);
nor U18098 (N_18098,N_17154,N_17563);
xor U18099 (N_18099,N_17963,N_17339);
and U18100 (N_18100,N_17689,N_17391);
nor U18101 (N_18101,N_17716,N_17989);
or U18102 (N_18102,N_17012,N_17983);
nand U18103 (N_18103,N_17351,N_17372);
nand U18104 (N_18104,N_17702,N_17127);
or U18105 (N_18105,N_17451,N_17573);
nand U18106 (N_18106,N_17875,N_17930);
nor U18107 (N_18107,N_17967,N_17867);
nor U18108 (N_18108,N_17899,N_17005);
or U18109 (N_18109,N_17773,N_17643);
or U18110 (N_18110,N_17250,N_17919);
nand U18111 (N_18111,N_17606,N_17353);
and U18112 (N_18112,N_17360,N_17921);
nand U18113 (N_18113,N_17354,N_17171);
nor U18114 (N_18114,N_17845,N_17379);
xnor U18115 (N_18115,N_17607,N_17077);
nand U18116 (N_18116,N_17130,N_17698);
nand U18117 (N_18117,N_17440,N_17048);
or U18118 (N_18118,N_17468,N_17424);
xor U18119 (N_18119,N_17183,N_17775);
or U18120 (N_18120,N_17649,N_17388);
and U18121 (N_18121,N_17213,N_17728);
or U18122 (N_18122,N_17714,N_17385);
nand U18123 (N_18123,N_17694,N_17695);
xnor U18124 (N_18124,N_17501,N_17752);
nor U18125 (N_18125,N_17105,N_17276);
xnor U18126 (N_18126,N_17768,N_17033);
nand U18127 (N_18127,N_17206,N_17956);
and U18128 (N_18128,N_17641,N_17199);
nand U18129 (N_18129,N_17305,N_17094);
nor U18130 (N_18130,N_17320,N_17045);
and U18131 (N_18131,N_17493,N_17057);
and U18132 (N_18132,N_17818,N_17751);
xor U18133 (N_18133,N_17605,N_17292);
xor U18134 (N_18134,N_17435,N_17230);
and U18135 (N_18135,N_17035,N_17335);
xnor U18136 (N_18136,N_17330,N_17507);
xor U18137 (N_18137,N_17913,N_17988);
nor U18138 (N_18138,N_17426,N_17101);
nand U18139 (N_18139,N_17950,N_17535);
xor U18140 (N_18140,N_17098,N_17603);
nor U18141 (N_18141,N_17122,N_17194);
and U18142 (N_18142,N_17415,N_17526);
xnor U18143 (N_18143,N_17664,N_17633);
or U18144 (N_18144,N_17790,N_17533);
nor U18145 (N_18145,N_17108,N_17028);
xnor U18146 (N_18146,N_17681,N_17298);
nor U18147 (N_18147,N_17422,N_17525);
xnor U18148 (N_18148,N_17660,N_17067);
nor U18149 (N_18149,N_17026,N_17759);
nor U18150 (N_18150,N_17974,N_17207);
and U18151 (N_18151,N_17833,N_17706);
nand U18152 (N_18152,N_17948,N_17043);
nand U18153 (N_18153,N_17369,N_17991);
xor U18154 (N_18154,N_17500,N_17715);
nand U18155 (N_18155,N_17866,N_17120);
nor U18156 (N_18156,N_17815,N_17144);
and U18157 (N_18157,N_17348,N_17251);
nor U18158 (N_18158,N_17279,N_17310);
xor U18159 (N_18159,N_17241,N_17647);
nand U18160 (N_18160,N_17718,N_17049);
xnor U18161 (N_18161,N_17037,N_17551);
nor U18162 (N_18162,N_17826,N_17585);
or U18163 (N_18163,N_17465,N_17029);
and U18164 (N_18164,N_17739,N_17879);
xnor U18165 (N_18165,N_17722,N_17789);
or U18166 (N_18166,N_17598,N_17161);
nand U18167 (N_18167,N_17784,N_17872);
or U18168 (N_18168,N_17644,N_17847);
xnor U18169 (N_18169,N_17568,N_17793);
xnor U18170 (N_18170,N_17530,N_17002);
or U18171 (N_18171,N_17180,N_17788);
nor U18172 (N_18172,N_17217,N_17682);
nand U18173 (N_18173,N_17985,N_17579);
nor U18174 (N_18174,N_17418,N_17289);
or U18175 (N_18175,N_17581,N_17665);
or U18176 (N_18176,N_17811,N_17225);
or U18177 (N_18177,N_17392,N_17078);
and U18178 (N_18178,N_17381,N_17562);
nor U18179 (N_18179,N_17515,N_17856);
nand U18180 (N_18180,N_17806,N_17733);
nor U18181 (N_18181,N_17510,N_17547);
and U18182 (N_18182,N_17475,N_17223);
or U18183 (N_18183,N_17125,N_17852);
and U18184 (N_18184,N_17982,N_17177);
xor U18185 (N_18185,N_17592,N_17454);
nand U18186 (N_18186,N_17513,N_17024);
nand U18187 (N_18187,N_17931,N_17726);
or U18188 (N_18188,N_17830,N_17889);
or U18189 (N_18189,N_17051,N_17179);
or U18190 (N_18190,N_17518,N_17687);
nand U18191 (N_18191,N_17295,N_17481);
nor U18192 (N_18192,N_17741,N_17758);
nand U18193 (N_18193,N_17222,N_17756);
nor U18194 (N_18194,N_17860,N_17308);
or U18195 (N_18195,N_17795,N_17554);
or U18196 (N_18196,N_17018,N_17020);
or U18197 (N_18197,N_17677,N_17819);
and U18198 (N_18198,N_17343,N_17326);
nand U18199 (N_18199,N_17229,N_17999);
xor U18200 (N_18200,N_17648,N_17302);
xor U18201 (N_18201,N_17524,N_17162);
nor U18202 (N_18202,N_17560,N_17742);
xor U18203 (N_18203,N_17590,N_17853);
xor U18204 (N_18204,N_17783,N_17538);
nor U18205 (N_18205,N_17673,N_17091);
nor U18206 (N_18206,N_17639,N_17270);
nand U18207 (N_18207,N_17132,N_17210);
xnor U18208 (N_18208,N_17763,N_17380);
and U18209 (N_18209,N_17534,N_17490);
and U18210 (N_18210,N_17447,N_17374);
nand U18211 (N_18211,N_17494,N_17692);
and U18212 (N_18212,N_17608,N_17635);
and U18213 (N_18213,N_17319,N_17915);
or U18214 (N_18214,N_17960,N_17086);
xnor U18215 (N_18215,N_17441,N_17700);
nor U18216 (N_18216,N_17572,N_17188);
nor U18217 (N_18217,N_17312,N_17972);
and U18218 (N_18218,N_17228,N_17710);
and U18219 (N_18219,N_17589,N_17755);
and U18220 (N_18220,N_17269,N_17614);
xnor U18221 (N_18221,N_17717,N_17129);
nor U18222 (N_18222,N_17656,N_17174);
and U18223 (N_18223,N_17448,N_17629);
or U18224 (N_18224,N_17946,N_17047);
and U18225 (N_18225,N_17271,N_17275);
xor U18226 (N_18226,N_17624,N_17640);
xnor U18227 (N_18227,N_17158,N_17119);
nor U18228 (N_18228,N_17013,N_17996);
nor U18229 (N_18229,N_17476,N_17044);
nor U18230 (N_18230,N_17015,N_17220);
xor U18231 (N_18231,N_17025,N_17394);
nand U18232 (N_18232,N_17400,N_17821);
xnor U18233 (N_18233,N_17034,N_17613);
or U18234 (N_18234,N_17906,N_17016);
or U18235 (N_18235,N_17027,N_17591);
xnor U18236 (N_18236,N_17685,N_17258);
xor U18237 (N_18237,N_17212,N_17705);
xnor U18238 (N_18238,N_17109,N_17157);
xor U18239 (N_18239,N_17508,N_17364);
xor U18240 (N_18240,N_17420,N_17621);
nor U18241 (N_18241,N_17693,N_17601);
nand U18242 (N_18242,N_17442,N_17911);
or U18243 (N_18243,N_17877,N_17285);
nor U18244 (N_18244,N_17630,N_17544);
nor U18245 (N_18245,N_17140,N_17464);
or U18246 (N_18246,N_17080,N_17181);
nand U18247 (N_18247,N_17128,N_17322);
xnor U18248 (N_18248,N_17557,N_17316);
xor U18249 (N_18249,N_17855,N_17617);
nor U18250 (N_18250,N_17042,N_17802);
and U18251 (N_18251,N_17709,N_17933);
nand U18252 (N_18252,N_17366,N_17227);
or U18253 (N_18253,N_17672,N_17263);
or U18254 (N_18254,N_17747,N_17779);
xor U18255 (N_18255,N_17347,N_17234);
or U18256 (N_18256,N_17987,N_17880);
and U18257 (N_18257,N_17615,N_17576);
or U18258 (N_18258,N_17349,N_17170);
xor U18259 (N_18259,N_17246,N_17910);
nor U18260 (N_18260,N_17434,N_17792);
or U18261 (N_18261,N_17934,N_17912);
or U18262 (N_18262,N_17517,N_17249);
nor U18263 (N_18263,N_17986,N_17300);
nand U18264 (N_18264,N_17404,N_17021);
nor U18265 (N_18265,N_17484,N_17262);
or U18266 (N_18266,N_17863,N_17307);
and U18267 (N_18267,N_17994,N_17564);
or U18268 (N_18268,N_17857,N_17187);
or U18269 (N_18269,N_17296,N_17425);
nand U18270 (N_18270,N_17291,N_17416);
nor U18271 (N_18271,N_17737,N_17586);
or U18272 (N_18272,N_17396,N_17201);
xnor U18273 (N_18273,N_17480,N_17399);
nand U18274 (N_18274,N_17650,N_17331);
nand U18275 (N_18275,N_17352,N_17965);
and U18276 (N_18276,N_17286,N_17746);
nand U18277 (N_18277,N_17618,N_17406);
and U18278 (N_18278,N_17456,N_17495);
nand U18279 (N_18279,N_17868,N_17940);
or U18280 (N_18280,N_17328,N_17839);
nand U18281 (N_18281,N_17727,N_17152);
xor U18282 (N_18282,N_17390,N_17071);
and U18283 (N_18283,N_17978,N_17927);
xor U18284 (N_18284,N_17864,N_17961);
nor U18285 (N_18285,N_17264,N_17657);
nand U18286 (N_18286,N_17093,N_17069);
or U18287 (N_18287,N_17503,N_17293);
nand U18288 (N_18288,N_17699,N_17762);
or U18289 (N_18289,N_17036,N_17951);
nor U18290 (N_18290,N_17890,N_17653);
nor U18291 (N_18291,N_17273,N_17421);
or U18292 (N_18292,N_17539,N_17469);
xnor U18293 (N_18293,N_17542,N_17578);
nand U18294 (N_18294,N_17886,N_17155);
nor U18295 (N_18295,N_17240,N_17457);
nand U18296 (N_18296,N_17964,N_17791);
nand U18297 (N_18297,N_17232,N_17894);
nor U18298 (N_18298,N_17859,N_17750);
nand U18299 (N_18299,N_17488,N_17007);
or U18300 (N_18300,N_17870,N_17124);
and U18301 (N_18301,N_17252,N_17173);
nor U18302 (N_18302,N_17509,N_17209);
or U18303 (N_18303,N_17216,N_17597);
nor U18304 (N_18304,N_17214,N_17907);
or U18305 (N_18305,N_17444,N_17023);
nand U18306 (N_18306,N_17938,N_17744);
or U18307 (N_18307,N_17567,N_17200);
nand U18308 (N_18308,N_17001,N_17580);
nor U18309 (N_18309,N_17704,N_17491);
and U18310 (N_18310,N_17735,N_17149);
xnor U18311 (N_18311,N_17334,N_17112);
nor U18312 (N_18312,N_17239,N_17817);
xnor U18313 (N_18313,N_17787,N_17287);
xor U18314 (N_18314,N_17014,N_17807);
and U18315 (N_18315,N_17439,N_17849);
nor U18316 (N_18316,N_17054,N_17492);
nand U18317 (N_18317,N_17935,N_17367);
nand U18318 (N_18318,N_17738,N_17203);
and U18319 (N_18319,N_17089,N_17011);
or U18320 (N_18320,N_17522,N_17099);
and U18321 (N_18321,N_17482,N_17126);
nand U18322 (N_18322,N_17370,N_17452);
or U18323 (N_18323,N_17226,N_17663);
and U18324 (N_18324,N_17268,N_17355);
or U18325 (N_18325,N_17713,N_17190);
nor U18326 (N_18326,N_17555,N_17117);
xor U18327 (N_18327,N_17981,N_17387);
nand U18328 (N_18328,N_17076,N_17486);
or U18329 (N_18329,N_17583,N_17949);
and U18330 (N_18330,N_17244,N_17595);
and U18331 (N_18331,N_17808,N_17383);
xnor U18332 (N_18332,N_17219,N_17511);
and U18333 (N_18333,N_17674,N_17652);
or U18334 (N_18334,N_17274,N_17896);
nor U18335 (N_18335,N_17947,N_17218);
and U18336 (N_18336,N_17655,N_17778);
xor U18337 (N_18337,N_17428,N_17602);
and U18338 (N_18338,N_17869,N_17184);
nand U18339 (N_18339,N_17552,N_17858);
and U18340 (N_18340,N_17836,N_17133);
and U18341 (N_18341,N_17850,N_17800);
nand U18342 (N_18342,N_17463,N_17167);
nor U18343 (N_18343,N_17609,N_17145);
xor U18344 (N_18344,N_17288,N_17204);
nand U18345 (N_18345,N_17523,N_17135);
or U18346 (N_18346,N_17697,N_17116);
xnor U18347 (N_18347,N_17008,N_17651);
xor U18348 (N_18348,N_17892,N_17010);
and U18349 (N_18349,N_17924,N_17980);
xnor U18350 (N_18350,N_17667,N_17160);
nor U18351 (N_18351,N_17905,N_17487);
nor U18352 (N_18352,N_17675,N_17088);
nand U18353 (N_18353,N_17055,N_17565);
or U18354 (N_18354,N_17703,N_17740);
and U18355 (N_18355,N_17701,N_17106);
or U18356 (N_18356,N_17211,N_17809);
and U18357 (N_18357,N_17306,N_17205);
and U18358 (N_18358,N_17473,N_17431);
xor U18359 (N_18359,N_17954,N_17942);
or U18360 (N_18360,N_17876,N_17842);
nor U18361 (N_18361,N_17402,N_17997);
or U18362 (N_18362,N_17131,N_17993);
nand U18363 (N_18363,N_17061,N_17096);
and U18364 (N_18364,N_17321,N_17680);
xnor U18365 (N_18365,N_17438,N_17691);
nor U18366 (N_18366,N_17537,N_17558);
xor U18367 (N_18367,N_17720,N_17900);
xnor U18368 (N_18368,N_17022,N_17327);
xor U18369 (N_18369,N_17032,N_17599);
xor U18370 (N_18370,N_17039,N_17358);
or U18371 (N_18371,N_17766,N_17984);
nor U18372 (N_18372,N_17313,N_17937);
xor U18373 (N_18373,N_17377,N_17670);
or U18374 (N_18374,N_17461,N_17479);
and U18375 (N_18375,N_17303,N_17172);
xor U18376 (N_18376,N_17134,N_17895);
nand U18377 (N_18377,N_17471,N_17242);
and U18378 (N_18378,N_17764,N_17176);
or U18379 (N_18379,N_17221,N_17519);
nand U18380 (N_18380,N_17662,N_17926);
xnor U18381 (N_18381,N_17333,N_17569);
or U18382 (N_18382,N_17062,N_17378);
or U18383 (N_18383,N_17311,N_17104);
xnor U18384 (N_18384,N_17959,N_17671);
nor U18385 (N_18385,N_17628,N_17528);
and U18386 (N_18386,N_17141,N_17556);
xor U18387 (N_18387,N_17782,N_17916);
nor U18388 (N_18388,N_17669,N_17499);
or U18389 (N_18389,N_17297,N_17843);
and U18390 (N_18390,N_17848,N_17068);
nor U18391 (N_18391,N_17841,N_17097);
xnor U18392 (N_18392,N_17090,N_17814);
xnor U18393 (N_18393,N_17403,N_17477);
or U18394 (N_18394,N_17893,N_17820);
or U18395 (N_18395,N_17604,N_17237);
nand U18396 (N_18396,N_17642,N_17118);
nor U18397 (N_18397,N_17329,N_17450);
or U18398 (N_18398,N_17970,N_17417);
xor U18399 (N_18399,N_17550,N_17266);
nand U18400 (N_18400,N_17245,N_17834);
nor U18401 (N_18401,N_17191,N_17540);
nand U18402 (N_18402,N_17952,N_17611);
nor U18403 (N_18403,N_17299,N_17243);
or U18404 (N_18404,N_17332,N_17975);
nor U18405 (N_18405,N_17038,N_17253);
or U18406 (N_18406,N_17185,N_17470);
nand U18407 (N_18407,N_17395,N_17957);
nor U18408 (N_18408,N_17357,N_17208);
nor U18409 (N_18409,N_17885,N_17769);
or U18410 (N_18410,N_17772,N_17146);
nand U18411 (N_18411,N_17163,N_17111);
nor U18412 (N_18412,N_17882,N_17918);
nand U18413 (N_18413,N_17346,N_17058);
nand U18414 (N_18414,N_17625,N_17521);
and U18415 (N_18415,N_17514,N_17459);
nor U18416 (N_18416,N_17883,N_17075);
nand U18417 (N_18417,N_17261,N_17577);
xor U18418 (N_18418,N_17267,N_17376);
or U18419 (N_18419,N_17917,N_17835);
nor U18420 (N_18420,N_17159,N_17884);
nand U18421 (N_18421,N_17797,N_17529);
nor U18422 (N_18422,N_17397,N_17247);
or U18423 (N_18423,N_17359,N_17588);
nor U18424 (N_18424,N_17719,N_17423);
nor U18425 (N_18425,N_17121,N_17255);
nor U18426 (N_18426,N_17944,N_17631);
nand U18427 (N_18427,N_17453,N_17574);
or U18428 (N_18428,N_17616,N_17559);
and U18429 (N_18429,N_17637,N_17259);
xnor U18430 (N_18430,N_17074,N_17192);
or U18431 (N_18431,N_17309,N_17798);
xor U18432 (N_18432,N_17731,N_17990);
or U18433 (N_18433,N_17337,N_17445);
nand U18434 (N_18434,N_17757,N_17186);
xnor U18435 (N_18435,N_17516,N_17169);
nand U18436 (N_18436,N_17139,N_17822);
or U18437 (N_18437,N_17543,N_17992);
nand U18438 (N_18438,N_17939,N_17256);
nor U18439 (N_18439,N_17138,N_17113);
or U18440 (N_18440,N_17622,N_17361);
nand U18441 (N_18441,N_17260,N_17813);
nand U18442 (N_18442,N_17323,N_17238);
and U18443 (N_18443,N_17941,N_17570);
nor U18444 (N_18444,N_17082,N_17000);
nor U18445 (N_18445,N_17596,N_17780);
xor U18446 (N_18446,N_17520,N_17945);
xnor U18447 (N_18447,N_17411,N_17063);
nor U18448 (N_18448,N_17362,N_17958);
nor U18449 (N_18449,N_17107,N_17371);
nor U18450 (N_18450,N_17050,N_17066);
and U18451 (N_18451,N_17873,N_17462);
and U18452 (N_18452,N_17363,N_17725);
xnor U18453 (N_18453,N_17748,N_17136);
or U18454 (N_18454,N_17587,N_17340);
xor U18455 (N_18455,N_17734,N_17829);
and U18456 (N_18456,N_17290,N_17966);
nand U18457 (N_18457,N_17084,N_17198);
nand U18458 (N_18458,N_17862,N_17898);
and U18459 (N_18459,N_17707,N_17231);
nor U18460 (N_18460,N_17549,N_17545);
and U18461 (N_18461,N_17962,N_17137);
nand U18462 (N_18462,N_17638,N_17708);
and U18463 (N_18463,N_17052,N_17536);
nand U18464 (N_18464,N_17925,N_17684);
and U18465 (N_18465,N_17661,N_17236);
nor U18466 (N_18466,N_17272,N_17474);
or U18467 (N_18467,N_17854,N_17840);
nand U18468 (N_18468,N_17142,N_17092);
and U18469 (N_18469,N_17498,N_17324);
xor U18470 (N_18470,N_17384,N_17030);
nor U18471 (N_18471,N_17754,N_17166);
or U18472 (N_18472,N_17165,N_17386);
or U18473 (N_18473,N_17446,N_17922);
nand U18474 (N_18474,N_17143,N_17823);
nor U18475 (N_18475,N_17301,N_17724);
nor U18476 (N_18476,N_17838,N_17600);
or U18477 (N_18477,N_17777,N_17760);
nand U18478 (N_18478,N_17006,N_17065);
and U18479 (N_18479,N_17774,N_17929);
or U18480 (N_18480,N_17745,N_17548);
xor U18481 (N_18481,N_17828,N_17278);
or U18482 (N_18482,N_17995,N_17831);
nor U18483 (N_18483,N_17496,N_17871);
and U18484 (N_18484,N_17393,N_17971);
xor U18485 (N_18485,N_17215,N_17019);
nand U18486 (N_18486,N_17785,N_17398);
xnor U18487 (N_18487,N_17413,N_17968);
nor U18488 (N_18488,N_17891,N_17645);
or U18489 (N_18489,N_17619,N_17233);
xnor U18490 (N_18490,N_17429,N_17100);
or U18491 (N_18491,N_17593,N_17283);
nor U18492 (N_18492,N_17794,N_17056);
or U18493 (N_18493,N_17796,N_17505);
and U18494 (N_18494,N_17150,N_17846);
nand U18495 (N_18495,N_17730,N_17419);
or U18496 (N_18496,N_17506,N_17224);
xor U18497 (N_18497,N_17771,N_17936);
nor U18498 (N_18498,N_17979,N_17711);
and U18499 (N_18499,N_17123,N_17485);
nand U18500 (N_18500,N_17717,N_17377);
nand U18501 (N_18501,N_17786,N_17081);
nor U18502 (N_18502,N_17717,N_17085);
nor U18503 (N_18503,N_17717,N_17957);
nand U18504 (N_18504,N_17011,N_17301);
nor U18505 (N_18505,N_17940,N_17709);
or U18506 (N_18506,N_17214,N_17141);
xnor U18507 (N_18507,N_17491,N_17682);
nand U18508 (N_18508,N_17816,N_17293);
nand U18509 (N_18509,N_17429,N_17064);
and U18510 (N_18510,N_17461,N_17480);
or U18511 (N_18511,N_17532,N_17827);
nand U18512 (N_18512,N_17250,N_17947);
xor U18513 (N_18513,N_17246,N_17695);
nand U18514 (N_18514,N_17723,N_17774);
and U18515 (N_18515,N_17298,N_17878);
nor U18516 (N_18516,N_17752,N_17308);
nand U18517 (N_18517,N_17497,N_17446);
nor U18518 (N_18518,N_17425,N_17886);
or U18519 (N_18519,N_17517,N_17497);
and U18520 (N_18520,N_17992,N_17228);
nor U18521 (N_18521,N_17969,N_17475);
nand U18522 (N_18522,N_17249,N_17150);
nor U18523 (N_18523,N_17629,N_17313);
nor U18524 (N_18524,N_17509,N_17314);
and U18525 (N_18525,N_17914,N_17724);
nand U18526 (N_18526,N_17981,N_17806);
nand U18527 (N_18527,N_17106,N_17193);
nand U18528 (N_18528,N_17007,N_17754);
nor U18529 (N_18529,N_17540,N_17282);
xor U18530 (N_18530,N_17399,N_17837);
xor U18531 (N_18531,N_17299,N_17829);
nand U18532 (N_18532,N_17968,N_17014);
nand U18533 (N_18533,N_17443,N_17887);
and U18534 (N_18534,N_17229,N_17883);
nor U18535 (N_18535,N_17656,N_17932);
xor U18536 (N_18536,N_17064,N_17172);
xor U18537 (N_18537,N_17883,N_17480);
xnor U18538 (N_18538,N_17650,N_17819);
nor U18539 (N_18539,N_17163,N_17918);
or U18540 (N_18540,N_17510,N_17339);
xor U18541 (N_18541,N_17082,N_17015);
or U18542 (N_18542,N_17125,N_17137);
and U18543 (N_18543,N_17110,N_17617);
nor U18544 (N_18544,N_17802,N_17294);
nand U18545 (N_18545,N_17046,N_17992);
nand U18546 (N_18546,N_17188,N_17330);
xnor U18547 (N_18547,N_17744,N_17524);
nand U18548 (N_18548,N_17808,N_17760);
nand U18549 (N_18549,N_17990,N_17186);
nor U18550 (N_18550,N_17244,N_17302);
nor U18551 (N_18551,N_17435,N_17042);
and U18552 (N_18552,N_17948,N_17653);
xor U18553 (N_18553,N_17351,N_17287);
nor U18554 (N_18554,N_17850,N_17243);
or U18555 (N_18555,N_17649,N_17895);
and U18556 (N_18556,N_17828,N_17640);
xor U18557 (N_18557,N_17739,N_17196);
and U18558 (N_18558,N_17349,N_17115);
nand U18559 (N_18559,N_17875,N_17331);
nor U18560 (N_18560,N_17944,N_17014);
xor U18561 (N_18561,N_17892,N_17511);
nor U18562 (N_18562,N_17519,N_17545);
nor U18563 (N_18563,N_17463,N_17350);
and U18564 (N_18564,N_17925,N_17650);
nand U18565 (N_18565,N_17986,N_17907);
nor U18566 (N_18566,N_17043,N_17328);
nand U18567 (N_18567,N_17835,N_17522);
and U18568 (N_18568,N_17393,N_17238);
nand U18569 (N_18569,N_17074,N_17373);
xor U18570 (N_18570,N_17654,N_17558);
xor U18571 (N_18571,N_17577,N_17403);
xnor U18572 (N_18572,N_17020,N_17315);
nand U18573 (N_18573,N_17664,N_17186);
and U18574 (N_18574,N_17389,N_17101);
nor U18575 (N_18575,N_17708,N_17050);
nor U18576 (N_18576,N_17824,N_17646);
nand U18577 (N_18577,N_17621,N_17162);
nand U18578 (N_18578,N_17466,N_17069);
and U18579 (N_18579,N_17963,N_17829);
and U18580 (N_18580,N_17416,N_17648);
or U18581 (N_18581,N_17574,N_17778);
xor U18582 (N_18582,N_17097,N_17750);
or U18583 (N_18583,N_17295,N_17077);
or U18584 (N_18584,N_17705,N_17241);
nor U18585 (N_18585,N_17303,N_17943);
nor U18586 (N_18586,N_17025,N_17166);
nor U18587 (N_18587,N_17076,N_17777);
nand U18588 (N_18588,N_17711,N_17030);
nor U18589 (N_18589,N_17931,N_17337);
xnor U18590 (N_18590,N_17595,N_17028);
or U18591 (N_18591,N_17268,N_17413);
and U18592 (N_18592,N_17929,N_17746);
nand U18593 (N_18593,N_17104,N_17019);
nand U18594 (N_18594,N_17080,N_17248);
and U18595 (N_18595,N_17732,N_17481);
and U18596 (N_18596,N_17444,N_17989);
or U18597 (N_18597,N_17724,N_17596);
xor U18598 (N_18598,N_17642,N_17459);
nor U18599 (N_18599,N_17199,N_17990);
nand U18600 (N_18600,N_17711,N_17370);
nand U18601 (N_18601,N_17885,N_17830);
and U18602 (N_18602,N_17783,N_17433);
and U18603 (N_18603,N_17670,N_17081);
xnor U18604 (N_18604,N_17046,N_17924);
or U18605 (N_18605,N_17897,N_17437);
nand U18606 (N_18606,N_17809,N_17138);
nor U18607 (N_18607,N_17900,N_17686);
xnor U18608 (N_18608,N_17100,N_17498);
nor U18609 (N_18609,N_17533,N_17519);
and U18610 (N_18610,N_17329,N_17925);
xor U18611 (N_18611,N_17495,N_17457);
nand U18612 (N_18612,N_17618,N_17238);
xor U18613 (N_18613,N_17635,N_17890);
nor U18614 (N_18614,N_17359,N_17141);
nor U18615 (N_18615,N_17198,N_17529);
or U18616 (N_18616,N_17587,N_17491);
nand U18617 (N_18617,N_17561,N_17790);
or U18618 (N_18618,N_17958,N_17188);
or U18619 (N_18619,N_17583,N_17899);
and U18620 (N_18620,N_17345,N_17370);
or U18621 (N_18621,N_17715,N_17328);
xnor U18622 (N_18622,N_17429,N_17442);
and U18623 (N_18623,N_17935,N_17184);
or U18624 (N_18624,N_17184,N_17202);
nand U18625 (N_18625,N_17334,N_17391);
xnor U18626 (N_18626,N_17400,N_17231);
or U18627 (N_18627,N_17858,N_17401);
and U18628 (N_18628,N_17993,N_17146);
and U18629 (N_18629,N_17539,N_17263);
nor U18630 (N_18630,N_17527,N_17516);
or U18631 (N_18631,N_17202,N_17665);
or U18632 (N_18632,N_17486,N_17814);
nor U18633 (N_18633,N_17838,N_17615);
nand U18634 (N_18634,N_17861,N_17027);
and U18635 (N_18635,N_17131,N_17783);
xnor U18636 (N_18636,N_17895,N_17680);
or U18637 (N_18637,N_17511,N_17866);
xor U18638 (N_18638,N_17359,N_17155);
nor U18639 (N_18639,N_17697,N_17434);
or U18640 (N_18640,N_17237,N_17550);
nor U18641 (N_18641,N_17723,N_17837);
nor U18642 (N_18642,N_17312,N_17687);
or U18643 (N_18643,N_17796,N_17826);
nor U18644 (N_18644,N_17839,N_17184);
xor U18645 (N_18645,N_17918,N_17060);
nor U18646 (N_18646,N_17621,N_17883);
and U18647 (N_18647,N_17227,N_17709);
nand U18648 (N_18648,N_17881,N_17364);
nand U18649 (N_18649,N_17608,N_17801);
xnor U18650 (N_18650,N_17554,N_17020);
nand U18651 (N_18651,N_17930,N_17402);
xnor U18652 (N_18652,N_17798,N_17543);
xor U18653 (N_18653,N_17024,N_17863);
nor U18654 (N_18654,N_17327,N_17157);
and U18655 (N_18655,N_17926,N_17375);
nand U18656 (N_18656,N_17278,N_17611);
nand U18657 (N_18657,N_17004,N_17043);
and U18658 (N_18658,N_17814,N_17854);
or U18659 (N_18659,N_17598,N_17496);
and U18660 (N_18660,N_17514,N_17928);
xor U18661 (N_18661,N_17023,N_17624);
and U18662 (N_18662,N_17358,N_17587);
nand U18663 (N_18663,N_17346,N_17525);
or U18664 (N_18664,N_17969,N_17911);
or U18665 (N_18665,N_17495,N_17189);
and U18666 (N_18666,N_17490,N_17162);
nand U18667 (N_18667,N_17284,N_17458);
xnor U18668 (N_18668,N_17252,N_17395);
or U18669 (N_18669,N_17430,N_17059);
or U18670 (N_18670,N_17946,N_17989);
xor U18671 (N_18671,N_17345,N_17127);
nor U18672 (N_18672,N_17256,N_17429);
nor U18673 (N_18673,N_17056,N_17116);
or U18674 (N_18674,N_17825,N_17209);
xor U18675 (N_18675,N_17118,N_17440);
and U18676 (N_18676,N_17767,N_17335);
nand U18677 (N_18677,N_17893,N_17343);
or U18678 (N_18678,N_17919,N_17265);
xnor U18679 (N_18679,N_17287,N_17291);
xor U18680 (N_18680,N_17278,N_17961);
nand U18681 (N_18681,N_17334,N_17770);
nand U18682 (N_18682,N_17048,N_17390);
xnor U18683 (N_18683,N_17792,N_17243);
nor U18684 (N_18684,N_17427,N_17159);
xor U18685 (N_18685,N_17264,N_17319);
xnor U18686 (N_18686,N_17407,N_17734);
nor U18687 (N_18687,N_17357,N_17148);
nor U18688 (N_18688,N_17379,N_17749);
nand U18689 (N_18689,N_17982,N_17145);
nor U18690 (N_18690,N_17686,N_17370);
nor U18691 (N_18691,N_17537,N_17148);
and U18692 (N_18692,N_17012,N_17170);
nand U18693 (N_18693,N_17002,N_17504);
or U18694 (N_18694,N_17154,N_17038);
nor U18695 (N_18695,N_17229,N_17317);
and U18696 (N_18696,N_17859,N_17572);
nor U18697 (N_18697,N_17240,N_17366);
or U18698 (N_18698,N_17295,N_17950);
or U18699 (N_18699,N_17136,N_17897);
or U18700 (N_18700,N_17062,N_17004);
and U18701 (N_18701,N_17890,N_17274);
nand U18702 (N_18702,N_17566,N_17374);
or U18703 (N_18703,N_17240,N_17981);
or U18704 (N_18704,N_17856,N_17750);
or U18705 (N_18705,N_17244,N_17406);
and U18706 (N_18706,N_17226,N_17939);
xor U18707 (N_18707,N_17577,N_17021);
or U18708 (N_18708,N_17959,N_17168);
and U18709 (N_18709,N_17984,N_17702);
nand U18710 (N_18710,N_17840,N_17051);
nand U18711 (N_18711,N_17355,N_17682);
xor U18712 (N_18712,N_17439,N_17435);
nor U18713 (N_18713,N_17851,N_17950);
and U18714 (N_18714,N_17894,N_17383);
and U18715 (N_18715,N_17982,N_17231);
or U18716 (N_18716,N_17689,N_17902);
and U18717 (N_18717,N_17471,N_17582);
and U18718 (N_18718,N_17047,N_17013);
nand U18719 (N_18719,N_17101,N_17652);
nand U18720 (N_18720,N_17187,N_17585);
xor U18721 (N_18721,N_17998,N_17379);
nand U18722 (N_18722,N_17301,N_17923);
nor U18723 (N_18723,N_17087,N_17129);
or U18724 (N_18724,N_17638,N_17129);
nor U18725 (N_18725,N_17254,N_17971);
or U18726 (N_18726,N_17714,N_17502);
and U18727 (N_18727,N_17493,N_17990);
and U18728 (N_18728,N_17254,N_17925);
nor U18729 (N_18729,N_17435,N_17926);
and U18730 (N_18730,N_17900,N_17805);
xnor U18731 (N_18731,N_17699,N_17127);
or U18732 (N_18732,N_17673,N_17463);
or U18733 (N_18733,N_17955,N_17099);
xnor U18734 (N_18734,N_17503,N_17319);
and U18735 (N_18735,N_17665,N_17340);
nor U18736 (N_18736,N_17484,N_17339);
and U18737 (N_18737,N_17723,N_17140);
xor U18738 (N_18738,N_17238,N_17817);
xor U18739 (N_18739,N_17524,N_17399);
xnor U18740 (N_18740,N_17523,N_17735);
and U18741 (N_18741,N_17843,N_17774);
nand U18742 (N_18742,N_17264,N_17123);
nor U18743 (N_18743,N_17813,N_17434);
xnor U18744 (N_18744,N_17137,N_17017);
xor U18745 (N_18745,N_17265,N_17484);
nand U18746 (N_18746,N_17178,N_17504);
nand U18747 (N_18747,N_17080,N_17830);
and U18748 (N_18748,N_17152,N_17416);
nor U18749 (N_18749,N_17813,N_17367);
or U18750 (N_18750,N_17524,N_17552);
xor U18751 (N_18751,N_17198,N_17262);
and U18752 (N_18752,N_17206,N_17545);
nand U18753 (N_18753,N_17545,N_17862);
or U18754 (N_18754,N_17434,N_17659);
or U18755 (N_18755,N_17868,N_17930);
or U18756 (N_18756,N_17353,N_17519);
xnor U18757 (N_18757,N_17128,N_17281);
and U18758 (N_18758,N_17683,N_17136);
nand U18759 (N_18759,N_17111,N_17579);
nand U18760 (N_18760,N_17557,N_17586);
nor U18761 (N_18761,N_17196,N_17980);
and U18762 (N_18762,N_17557,N_17416);
or U18763 (N_18763,N_17402,N_17574);
and U18764 (N_18764,N_17251,N_17572);
xor U18765 (N_18765,N_17233,N_17713);
nand U18766 (N_18766,N_17815,N_17758);
nand U18767 (N_18767,N_17617,N_17642);
nor U18768 (N_18768,N_17836,N_17008);
xnor U18769 (N_18769,N_17824,N_17201);
nor U18770 (N_18770,N_17967,N_17901);
nor U18771 (N_18771,N_17389,N_17917);
xor U18772 (N_18772,N_17069,N_17563);
nand U18773 (N_18773,N_17447,N_17498);
and U18774 (N_18774,N_17750,N_17473);
nand U18775 (N_18775,N_17947,N_17051);
nor U18776 (N_18776,N_17183,N_17611);
nand U18777 (N_18777,N_17568,N_17678);
nand U18778 (N_18778,N_17827,N_17678);
and U18779 (N_18779,N_17989,N_17955);
nor U18780 (N_18780,N_17590,N_17624);
nor U18781 (N_18781,N_17061,N_17071);
or U18782 (N_18782,N_17895,N_17212);
and U18783 (N_18783,N_17452,N_17831);
nor U18784 (N_18784,N_17210,N_17854);
and U18785 (N_18785,N_17714,N_17445);
xor U18786 (N_18786,N_17874,N_17702);
or U18787 (N_18787,N_17141,N_17613);
and U18788 (N_18788,N_17405,N_17981);
or U18789 (N_18789,N_17655,N_17908);
nand U18790 (N_18790,N_17387,N_17060);
nand U18791 (N_18791,N_17873,N_17321);
or U18792 (N_18792,N_17750,N_17659);
nand U18793 (N_18793,N_17908,N_17269);
or U18794 (N_18794,N_17481,N_17453);
nor U18795 (N_18795,N_17629,N_17722);
nand U18796 (N_18796,N_17099,N_17442);
or U18797 (N_18797,N_17995,N_17465);
xnor U18798 (N_18798,N_17422,N_17657);
nor U18799 (N_18799,N_17710,N_17560);
or U18800 (N_18800,N_17001,N_17682);
xnor U18801 (N_18801,N_17607,N_17354);
nand U18802 (N_18802,N_17092,N_17147);
and U18803 (N_18803,N_17573,N_17870);
and U18804 (N_18804,N_17663,N_17693);
nand U18805 (N_18805,N_17870,N_17841);
or U18806 (N_18806,N_17659,N_17646);
and U18807 (N_18807,N_17144,N_17203);
nand U18808 (N_18808,N_17560,N_17153);
xnor U18809 (N_18809,N_17972,N_17975);
nor U18810 (N_18810,N_17209,N_17703);
nor U18811 (N_18811,N_17674,N_17147);
and U18812 (N_18812,N_17722,N_17316);
nand U18813 (N_18813,N_17764,N_17543);
or U18814 (N_18814,N_17169,N_17419);
or U18815 (N_18815,N_17010,N_17798);
or U18816 (N_18816,N_17105,N_17172);
and U18817 (N_18817,N_17717,N_17099);
nand U18818 (N_18818,N_17854,N_17434);
or U18819 (N_18819,N_17193,N_17729);
and U18820 (N_18820,N_17081,N_17590);
nor U18821 (N_18821,N_17761,N_17141);
or U18822 (N_18822,N_17121,N_17001);
nor U18823 (N_18823,N_17955,N_17430);
xnor U18824 (N_18824,N_17836,N_17240);
or U18825 (N_18825,N_17253,N_17107);
or U18826 (N_18826,N_17709,N_17850);
nor U18827 (N_18827,N_17268,N_17983);
nand U18828 (N_18828,N_17546,N_17248);
xor U18829 (N_18829,N_17317,N_17786);
nor U18830 (N_18830,N_17026,N_17601);
nor U18831 (N_18831,N_17569,N_17383);
or U18832 (N_18832,N_17894,N_17562);
or U18833 (N_18833,N_17325,N_17958);
or U18834 (N_18834,N_17725,N_17494);
and U18835 (N_18835,N_17630,N_17900);
and U18836 (N_18836,N_17492,N_17951);
or U18837 (N_18837,N_17827,N_17078);
and U18838 (N_18838,N_17132,N_17573);
xnor U18839 (N_18839,N_17122,N_17953);
and U18840 (N_18840,N_17149,N_17340);
or U18841 (N_18841,N_17590,N_17831);
xor U18842 (N_18842,N_17817,N_17709);
and U18843 (N_18843,N_17487,N_17402);
nor U18844 (N_18844,N_17682,N_17698);
xor U18845 (N_18845,N_17032,N_17305);
and U18846 (N_18846,N_17501,N_17848);
and U18847 (N_18847,N_17401,N_17443);
xnor U18848 (N_18848,N_17917,N_17291);
xnor U18849 (N_18849,N_17908,N_17401);
or U18850 (N_18850,N_17906,N_17368);
nor U18851 (N_18851,N_17267,N_17453);
nand U18852 (N_18852,N_17975,N_17364);
nand U18853 (N_18853,N_17103,N_17367);
or U18854 (N_18854,N_17858,N_17644);
xor U18855 (N_18855,N_17136,N_17605);
xnor U18856 (N_18856,N_17145,N_17967);
nand U18857 (N_18857,N_17296,N_17255);
xor U18858 (N_18858,N_17587,N_17646);
nor U18859 (N_18859,N_17250,N_17986);
nor U18860 (N_18860,N_17767,N_17548);
xor U18861 (N_18861,N_17088,N_17845);
and U18862 (N_18862,N_17758,N_17570);
nor U18863 (N_18863,N_17251,N_17088);
and U18864 (N_18864,N_17623,N_17919);
and U18865 (N_18865,N_17659,N_17135);
nor U18866 (N_18866,N_17206,N_17768);
xnor U18867 (N_18867,N_17799,N_17430);
xor U18868 (N_18868,N_17882,N_17526);
or U18869 (N_18869,N_17426,N_17305);
nor U18870 (N_18870,N_17753,N_17722);
or U18871 (N_18871,N_17804,N_17706);
and U18872 (N_18872,N_17943,N_17586);
or U18873 (N_18873,N_17069,N_17755);
xor U18874 (N_18874,N_17758,N_17829);
nand U18875 (N_18875,N_17383,N_17278);
nand U18876 (N_18876,N_17336,N_17864);
nor U18877 (N_18877,N_17050,N_17154);
or U18878 (N_18878,N_17947,N_17858);
nand U18879 (N_18879,N_17178,N_17511);
or U18880 (N_18880,N_17168,N_17104);
and U18881 (N_18881,N_17329,N_17297);
xnor U18882 (N_18882,N_17182,N_17581);
and U18883 (N_18883,N_17385,N_17802);
or U18884 (N_18884,N_17024,N_17605);
nand U18885 (N_18885,N_17840,N_17103);
or U18886 (N_18886,N_17002,N_17871);
nand U18887 (N_18887,N_17058,N_17266);
and U18888 (N_18888,N_17812,N_17255);
nand U18889 (N_18889,N_17662,N_17442);
nand U18890 (N_18890,N_17015,N_17023);
xor U18891 (N_18891,N_17345,N_17447);
nor U18892 (N_18892,N_17628,N_17659);
and U18893 (N_18893,N_17803,N_17780);
xnor U18894 (N_18894,N_17850,N_17961);
nand U18895 (N_18895,N_17858,N_17888);
nor U18896 (N_18896,N_17837,N_17792);
and U18897 (N_18897,N_17415,N_17811);
and U18898 (N_18898,N_17201,N_17377);
and U18899 (N_18899,N_17351,N_17152);
nor U18900 (N_18900,N_17037,N_17598);
xnor U18901 (N_18901,N_17375,N_17100);
and U18902 (N_18902,N_17037,N_17909);
xor U18903 (N_18903,N_17800,N_17629);
or U18904 (N_18904,N_17156,N_17190);
nor U18905 (N_18905,N_17276,N_17442);
and U18906 (N_18906,N_17128,N_17454);
nand U18907 (N_18907,N_17248,N_17698);
xor U18908 (N_18908,N_17269,N_17070);
nor U18909 (N_18909,N_17664,N_17718);
xnor U18910 (N_18910,N_17278,N_17701);
xnor U18911 (N_18911,N_17676,N_17843);
and U18912 (N_18912,N_17567,N_17292);
and U18913 (N_18913,N_17102,N_17637);
and U18914 (N_18914,N_17901,N_17471);
or U18915 (N_18915,N_17758,N_17415);
xor U18916 (N_18916,N_17354,N_17190);
nand U18917 (N_18917,N_17754,N_17462);
xor U18918 (N_18918,N_17808,N_17065);
and U18919 (N_18919,N_17712,N_17062);
xor U18920 (N_18920,N_17778,N_17151);
nand U18921 (N_18921,N_17697,N_17828);
and U18922 (N_18922,N_17228,N_17601);
nand U18923 (N_18923,N_17287,N_17190);
nor U18924 (N_18924,N_17308,N_17022);
xor U18925 (N_18925,N_17874,N_17594);
nand U18926 (N_18926,N_17518,N_17289);
xor U18927 (N_18927,N_17070,N_17555);
xnor U18928 (N_18928,N_17566,N_17313);
nand U18929 (N_18929,N_17784,N_17260);
or U18930 (N_18930,N_17857,N_17760);
and U18931 (N_18931,N_17428,N_17225);
or U18932 (N_18932,N_17835,N_17123);
and U18933 (N_18933,N_17779,N_17986);
nor U18934 (N_18934,N_17072,N_17282);
and U18935 (N_18935,N_17146,N_17385);
xnor U18936 (N_18936,N_17923,N_17428);
nand U18937 (N_18937,N_17516,N_17553);
and U18938 (N_18938,N_17596,N_17010);
nand U18939 (N_18939,N_17048,N_17170);
nand U18940 (N_18940,N_17642,N_17170);
or U18941 (N_18941,N_17069,N_17770);
nor U18942 (N_18942,N_17826,N_17267);
or U18943 (N_18943,N_17578,N_17306);
or U18944 (N_18944,N_17180,N_17083);
and U18945 (N_18945,N_17523,N_17188);
or U18946 (N_18946,N_17109,N_17519);
xor U18947 (N_18947,N_17436,N_17064);
or U18948 (N_18948,N_17855,N_17647);
nand U18949 (N_18949,N_17515,N_17818);
nand U18950 (N_18950,N_17074,N_17525);
xnor U18951 (N_18951,N_17421,N_17460);
or U18952 (N_18952,N_17054,N_17511);
nand U18953 (N_18953,N_17318,N_17880);
nand U18954 (N_18954,N_17623,N_17812);
nand U18955 (N_18955,N_17938,N_17625);
xor U18956 (N_18956,N_17159,N_17880);
and U18957 (N_18957,N_17694,N_17394);
xor U18958 (N_18958,N_17099,N_17516);
xor U18959 (N_18959,N_17595,N_17466);
nand U18960 (N_18960,N_17471,N_17116);
and U18961 (N_18961,N_17328,N_17879);
nor U18962 (N_18962,N_17361,N_17350);
nand U18963 (N_18963,N_17110,N_17165);
or U18964 (N_18964,N_17067,N_17729);
nor U18965 (N_18965,N_17686,N_17877);
or U18966 (N_18966,N_17045,N_17731);
xor U18967 (N_18967,N_17091,N_17237);
and U18968 (N_18968,N_17971,N_17144);
nor U18969 (N_18969,N_17913,N_17886);
nor U18970 (N_18970,N_17313,N_17677);
and U18971 (N_18971,N_17957,N_17482);
and U18972 (N_18972,N_17580,N_17525);
xor U18973 (N_18973,N_17274,N_17469);
nand U18974 (N_18974,N_17242,N_17713);
nand U18975 (N_18975,N_17372,N_17314);
nand U18976 (N_18976,N_17003,N_17835);
xnor U18977 (N_18977,N_17359,N_17322);
nor U18978 (N_18978,N_17152,N_17089);
nor U18979 (N_18979,N_17272,N_17457);
nor U18980 (N_18980,N_17203,N_17406);
xnor U18981 (N_18981,N_17028,N_17869);
xor U18982 (N_18982,N_17013,N_17526);
nand U18983 (N_18983,N_17991,N_17390);
xnor U18984 (N_18984,N_17110,N_17347);
nor U18985 (N_18985,N_17620,N_17484);
and U18986 (N_18986,N_17844,N_17816);
nand U18987 (N_18987,N_17741,N_17977);
nor U18988 (N_18988,N_17297,N_17385);
nor U18989 (N_18989,N_17664,N_17505);
nor U18990 (N_18990,N_17211,N_17993);
or U18991 (N_18991,N_17200,N_17893);
and U18992 (N_18992,N_17379,N_17042);
xor U18993 (N_18993,N_17711,N_17179);
nor U18994 (N_18994,N_17598,N_17955);
and U18995 (N_18995,N_17503,N_17518);
nor U18996 (N_18996,N_17725,N_17160);
nor U18997 (N_18997,N_17899,N_17368);
nand U18998 (N_18998,N_17855,N_17457);
nand U18999 (N_18999,N_17907,N_17530);
xnor U19000 (N_19000,N_18056,N_18771);
xnor U19001 (N_19001,N_18029,N_18570);
and U19002 (N_19002,N_18469,N_18114);
nand U19003 (N_19003,N_18211,N_18822);
and U19004 (N_19004,N_18895,N_18388);
xor U19005 (N_19005,N_18195,N_18662);
or U19006 (N_19006,N_18117,N_18521);
nor U19007 (N_19007,N_18476,N_18333);
nor U19008 (N_19008,N_18269,N_18849);
nand U19009 (N_19009,N_18463,N_18228);
nand U19010 (N_19010,N_18216,N_18322);
or U19011 (N_19011,N_18430,N_18580);
xnor U19012 (N_19012,N_18185,N_18670);
xnor U19013 (N_19013,N_18827,N_18561);
or U19014 (N_19014,N_18278,N_18740);
nor U19015 (N_19015,N_18683,N_18960);
xnor U19016 (N_19016,N_18551,N_18439);
nor U19017 (N_19017,N_18001,N_18470);
nand U19018 (N_19018,N_18595,N_18692);
nand U19019 (N_19019,N_18268,N_18896);
nand U19020 (N_19020,N_18499,N_18651);
nand U19021 (N_19021,N_18397,N_18594);
xnor U19022 (N_19022,N_18673,N_18980);
or U19023 (N_19023,N_18017,N_18680);
or U19024 (N_19024,N_18031,N_18631);
nand U19025 (N_19025,N_18274,N_18254);
nand U19026 (N_19026,N_18644,N_18073);
xor U19027 (N_19027,N_18838,N_18824);
and U19028 (N_19028,N_18335,N_18128);
xnor U19029 (N_19029,N_18305,N_18668);
nor U19030 (N_19030,N_18474,N_18492);
and U19031 (N_19031,N_18303,N_18759);
xor U19032 (N_19032,N_18801,N_18317);
xor U19033 (N_19033,N_18091,N_18732);
nand U19034 (N_19034,N_18893,N_18377);
xnor U19035 (N_19035,N_18458,N_18378);
nor U19036 (N_19036,N_18196,N_18347);
xnor U19037 (N_19037,N_18675,N_18637);
or U19038 (N_19038,N_18601,N_18559);
or U19039 (N_19039,N_18634,N_18413);
nand U19040 (N_19040,N_18574,N_18910);
nor U19041 (N_19041,N_18197,N_18447);
nor U19042 (N_19042,N_18816,N_18194);
and U19043 (N_19043,N_18183,N_18524);
or U19044 (N_19044,N_18516,N_18190);
xnor U19045 (N_19045,N_18178,N_18563);
nor U19046 (N_19046,N_18703,N_18804);
xnor U19047 (N_19047,N_18622,N_18156);
and U19048 (N_19048,N_18267,N_18300);
and U19049 (N_19049,N_18752,N_18812);
nand U19050 (N_19050,N_18270,N_18766);
nor U19051 (N_19051,N_18215,N_18945);
xnor U19052 (N_19052,N_18768,N_18681);
or U19053 (N_19053,N_18359,N_18348);
and U19054 (N_19054,N_18172,N_18965);
nor U19055 (N_19055,N_18022,N_18481);
nor U19056 (N_19056,N_18493,N_18281);
nand U19057 (N_19057,N_18057,N_18297);
nand U19058 (N_19058,N_18449,N_18018);
nor U19059 (N_19059,N_18466,N_18315);
xnor U19060 (N_19060,N_18165,N_18402);
xor U19061 (N_19061,N_18072,N_18109);
and U19062 (N_19062,N_18730,N_18888);
nand U19063 (N_19063,N_18659,N_18951);
or U19064 (N_19064,N_18336,N_18189);
and U19065 (N_19065,N_18743,N_18598);
or U19066 (N_19066,N_18999,N_18608);
or U19067 (N_19067,N_18203,N_18296);
nor U19068 (N_19068,N_18357,N_18859);
nand U19069 (N_19069,N_18411,N_18177);
xor U19070 (N_19070,N_18238,N_18867);
and U19071 (N_19071,N_18519,N_18817);
nand U19072 (N_19072,N_18232,N_18331);
nand U19073 (N_19073,N_18913,N_18636);
nand U19074 (N_19074,N_18915,N_18009);
nand U19075 (N_19075,N_18299,N_18145);
nand U19076 (N_19076,N_18410,N_18632);
xor U19077 (N_19077,N_18095,N_18166);
or U19078 (N_19078,N_18955,N_18863);
xnor U19079 (N_19079,N_18635,N_18967);
nor U19080 (N_19080,N_18934,N_18656);
nand U19081 (N_19081,N_18080,N_18004);
xnor U19082 (N_19082,N_18369,N_18991);
or U19083 (N_19083,N_18019,N_18905);
nor U19084 (N_19084,N_18546,N_18865);
nor U19085 (N_19085,N_18749,N_18383);
xor U19086 (N_19086,N_18892,N_18465);
nand U19087 (N_19087,N_18415,N_18414);
or U19088 (N_19088,N_18682,N_18510);
nand U19089 (N_19089,N_18836,N_18878);
or U19090 (N_19090,N_18412,N_18974);
and U19091 (N_19091,N_18207,N_18167);
nand U19092 (N_19092,N_18605,N_18065);
nand U19093 (N_19093,N_18401,N_18987);
or U19094 (N_19094,N_18904,N_18082);
or U19095 (N_19095,N_18319,N_18107);
nor U19096 (N_19096,N_18294,N_18797);
nand U19097 (N_19097,N_18051,N_18445);
nand U19098 (N_19098,N_18421,N_18728);
nand U19099 (N_19099,N_18649,N_18747);
nand U19100 (N_19100,N_18814,N_18802);
nor U19101 (N_19101,N_18837,N_18137);
xnor U19102 (N_19102,N_18577,N_18223);
nand U19103 (N_19103,N_18852,N_18717);
xnor U19104 (N_19104,N_18220,N_18597);
and U19105 (N_19105,N_18125,N_18856);
nand U19106 (N_19106,N_18119,N_18028);
and U19107 (N_19107,N_18993,N_18919);
xnor U19108 (N_19108,N_18272,N_18337);
xor U19109 (N_19109,N_18209,N_18462);
nand U19110 (N_19110,N_18933,N_18809);
nor U19111 (N_19111,N_18526,N_18174);
nor U19112 (N_19112,N_18158,N_18050);
xor U19113 (N_19113,N_18777,N_18136);
nand U19114 (N_19114,N_18655,N_18338);
nand U19115 (N_19115,N_18456,N_18020);
nand U19116 (N_19116,N_18188,N_18826);
nor U19117 (N_19117,N_18611,N_18155);
nor U19118 (N_19118,N_18719,N_18342);
nor U19119 (N_19119,N_18503,N_18937);
xnor U19120 (N_19120,N_18828,N_18699);
xnor U19121 (N_19121,N_18427,N_18565);
nor U19122 (N_19122,N_18688,N_18164);
and U19123 (N_19123,N_18970,N_18061);
xor U19124 (N_19124,N_18154,N_18906);
or U19125 (N_19125,N_18021,N_18201);
xor U19126 (N_19126,N_18053,N_18286);
xor U19127 (N_19127,N_18063,N_18173);
xor U19128 (N_19128,N_18064,N_18600);
nor U19129 (N_19129,N_18576,N_18376);
or U19130 (N_19130,N_18442,N_18518);
xor U19131 (N_19131,N_18231,N_18494);
or U19132 (N_19132,N_18758,N_18697);
and U19133 (N_19133,N_18725,N_18566);
and U19134 (N_19134,N_18162,N_18111);
xor U19135 (N_19135,N_18657,N_18276);
xnor U19136 (N_19136,N_18473,N_18508);
nand U19137 (N_19137,N_18047,N_18149);
nor U19138 (N_19138,N_18938,N_18567);
nand U19139 (N_19139,N_18589,N_18040);
and U19140 (N_19140,N_18006,N_18762);
nand U19141 (N_19141,N_18687,N_18433);
nor U19142 (N_19142,N_18161,N_18460);
xnor U19143 (N_19143,N_18243,N_18710);
xor U19144 (N_19144,N_18448,N_18964);
nand U19145 (N_19145,N_18874,N_18182);
nor U19146 (N_19146,N_18988,N_18479);
or U19147 (N_19147,N_18030,N_18568);
nand U19148 (N_19148,N_18606,N_18897);
nand U19149 (N_19149,N_18490,N_18695);
or U19150 (N_19150,N_18391,N_18792);
and U19151 (N_19151,N_18429,N_18841);
nor U19152 (N_19152,N_18723,N_18943);
and U19153 (N_19153,N_18741,N_18092);
xor U19154 (N_19154,N_18144,N_18264);
xor U19155 (N_19155,N_18123,N_18693);
nor U19156 (N_19156,N_18779,N_18864);
and U19157 (N_19157,N_18418,N_18204);
or U19158 (N_19158,N_18776,N_18721);
or U19159 (N_19159,N_18773,N_18328);
and U19160 (N_19160,N_18187,N_18640);
xnor U19161 (N_19161,N_18461,N_18715);
nand U19162 (N_19162,N_18179,N_18074);
nand U19163 (N_19163,N_18726,N_18210);
and U19164 (N_19164,N_18525,N_18389);
or U19165 (N_19165,N_18579,N_18130);
xor U19166 (N_19166,N_18706,N_18014);
and U19167 (N_19167,N_18101,N_18782);
nand U19168 (N_19168,N_18587,N_18532);
or U19169 (N_19169,N_18971,N_18373);
xor U19170 (N_19170,N_18821,N_18240);
xor U19171 (N_19171,N_18894,N_18135);
and U19172 (N_19172,N_18285,N_18646);
or U19173 (N_19173,N_18265,N_18311);
and U19174 (N_19174,N_18116,N_18055);
xnor U19175 (N_19175,N_18027,N_18332);
and U19176 (N_19176,N_18396,N_18557);
nor U19177 (N_19177,N_18142,N_18395);
nand U19178 (N_19178,N_18948,N_18590);
nand U19179 (N_19179,N_18581,N_18536);
xor U19180 (N_19180,N_18700,N_18720);
nand U19181 (N_19181,N_18630,N_18374);
nand U19182 (N_19182,N_18879,N_18090);
nor U19183 (N_19183,N_18186,N_18247);
or U19184 (N_19184,N_18972,N_18868);
xor U19185 (N_19185,N_18086,N_18298);
and U19186 (N_19186,N_18538,N_18037);
nand U19187 (N_19187,N_18244,N_18550);
and U19188 (N_19188,N_18039,N_18160);
xnor U19189 (N_19189,N_18750,N_18251);
nand U19190 (N_19190,N_18925,N_18236);
nor U19191 (N_19191,N_18392,N_18224);
xor U19192 (N_19192,N_18578,N_18486);
nor U19193 (N_19193,N_18446,N_18290);
xnor U19194 (N_19194,N_18941,N_18434);
nor U19195 (N_19195,N_18045,N_18033);
xor U19196 (N_19196,N_18513,N_18077);
nor U19197 (N_19197,N_18898,N_18151);
or U19198 (N_19198,N_18918,N_18834);
and U19199 (N_19199,N_18032,N_18150);
and U19200 (N_19200,N_18643,N_18483);
or U19201 (N_19201,N_18853,N_18572);
and U19202 (N_19202,N_18321,N_18769);
and U19203 (N_19203,N_18855,N_18059);
nor U19204 (N_19204,N_18757,N_18094);
nor U19205 (N_19205,N_18908,N_18025);
nor U19206 (N_19206,N_18341,N_18043);
nor U19207 (N_19207,N_18422,N_18148);
nand U19208 (N_19208,N_18308,N_18184);
nand U19209 (N_19209,N_18873,N_18582);
xor U19210 (N_19210,N_18529,N_18275);
nand U19211 (N_19211,N_18736,N_18984);
nor U19212 (N_19212,N_18259,N_18255);
nor U19213 (N_19213,N_18157,N_18093);
or U19214 (N_19214,N_18181,N_18962);
and U19215 (N_19215,N_18356,N_18237);
nor U19216 (N_19216,N_18097,N_18935);
or U19217 (N_19217,N_18534,N_18927);
xor U19218 (N_19218,N_18813,N_18803);
xor U19219 (N_19219,N_18253,N_18035);
or U19220 (N_19220,N_18753,N_18542);
and U19221 (N_19221,N_18441,N_18126);
nand U19222 (N_19222,N_18671,N_18372);
and U19223 (N_19223,N_18366,N_18891);
and U19224 (N_19224,N_18667,N_18903);
or U19225 (N_19225,N_18121,N_18531);
nand U19226 (N_19226,N_18129,N_18507);
and U19227 (N_19227,N_18686,N_18553);
or U19228 (N_19228,N_18044,N_18786);
xnor U19229 (N_19229,N_18626,N_18046);
or U19230 (N_19230,N_18423,N_18241);
nor U19231 (N_19231,N_18607,N_18731);
xnor U19232 (N_19232,N_18942,N_18751);
nor U19233 (N_19233,N_18641,N_18295);
nand U19234 (N_19234,N_18451,N_18248);
and U19235 (N_19235,N_18318,N_18760);
xnor U19236 (N_19236,N_18217,N_18957);
or U19237 (N_19237,N_18176,N_18953);
and U19238 (N_19238,N_18857,N_18191);
or U19239 (N_19239,N_18528,N_18475);
and U19240 (N_19240,N_18602,N_18684);
or U19241 (N_19241,N_18523,N_18497);
and U19242 (N_19242,N_18940,N_18573);
or U19243 (N_19243,N_18963,N_18609);
xor U19244 (N_19244,N_18810,N_18159);
nand U19245 (N_19245,N_18540,N_18781);
or U19246 (N_19246,N_18008,N_18271);
xor U19247 (N_19247,N_18599,N_18085);
nand U19248 (N_19248,N_18844,N_18242);
xor U19249 (N_19249,N_18845,N_18936);
or U19250 (N_19250,N_18950,N_18990);
or U19251 (N_19251,N_18301,N_18979);
or U19252 (N_19252,N_18661,N_18115);
xnor U19253 (N_19253,N_18102,N_18424);
or U19254 (N_19254,N_18010,N_18304);
and U19255 (N_19255,N_18917,N_18007);
or U19256 (N_19256,N_18515,N_18808);
and U19257 (N_19257,N_18478,N_18920);
nand U19258 (N_19258,N_18306,N_18440);
nor U19259 (N_19259,N_18929,N_18192);
xor U19260 (N_19260,N_18928,N_18882);
and U19261 (N_19261,N_18875,N_18454);
nand U19262 (N_19262,N_18283,N_18261);
nand U19263 (N_19263,N_18024,N_18527);
or U19264 (N_19264,N_18835,N_18501);
and U19265 (N_19265,N_18370,N_18737);
and U19266 (N_19266,N_18807,N_18084);
nor U19267 (N_19267,N_18952,N_18729);
nand U19268 (N_19268,N_18754,N_18900);
xnor U19269 (N_19269,N_18112,N_18793);
and U19270 (N_19270,N_18070,N_18833);
xor U19271 (N_19271,N_18060,N_18509);
nand U19272 (N_19272,N_18947,N_18062);
nor U19273 (N_19273,N_18282,N_18761);
nor U19274 (N_19274,N_18639,N_18805);
nand U19275 (N_19275,N_18124,N_18537);
xor U19276 (N_19276,N_18789,N_18548);
and U19277 (N_19277,N_18256,N_18795);
xor U19278 (N_19278,N_18036,N_18847);
xor U19279 (N_19279,N_18489,N_18076);
nor U19280 (N_19280,N_18380,N_18628);
nand U19281 (N_19281,N_18914,N_18885);
nand U19282 (N_19282,N_18081,N_18075);
and U19283 (N_19283,N_18830,N_18825);
nor U19284 (N_19284,N_18419,N_18616);
xor U19285 (N_19285,N_18484,N_18417);
nor U19286 (N_19286,N_18707,N_18664);
nand U19287 (N_19287,N_18648,N_18214);
nand U19288 (N_19288,N_18712,N_18949);
or U19289 (N_19289,N_18624,N_18390);
nand U19290 (N_19290,N_18405,N_18170);
and U19291 (N_19291,N_18502,N_18386);
nor U19292 (N_19292,N_18998,N_18617);
and U19293 (N_19293,N_18069,N_18504);
nand U19294 (N_19294,N_18742,N_18200);
xnor U19295 (N_19295,N_18213,N_18250);
xnor U19296 (N_19296,N_18312,N_18288);
or U19297 (N_19297,N_18778,N_18431);
or U19298 (N_19298,N_18575,N_18978);
or U19299 (N_19299,N_18477,N_18310);
xnor U19300 (N_19300,N_18926,N_18067);
xor U19301 (N_19301,N_18593,N_18564);
or U19302 (N_19302,N_18467,N_18280);
nand U19303 (N_19303,N_18485,N_18302);
nor U19304 (N_19304,N_18552,N_18716);
and U19305 (N_19305,N_18482,N_18514);
xor U19306 (N_19306,N_18708,N_18108);
and U19307 (N_19307,N_18432,N_18225);
nor U19308 (N_19308,N_18881,N_18541);
and U19309 (N_19309,N_18916,N_18691);
nor U19310 (N_19310,N_18175,N_18104);
xnor U19311 (N_19311,N_18398,N_18367);
nand U19312 (N_19312,N_18379,N_18235);
or U19313 (N_19313,N_18887,N_18351);
and U19314 (N_19314,N_18924,N_18698);
nor U19315 (N_19315,N_18153,N_18629);
and U19316 (N_19316,N_18132,N_18774);
nor U19317 (N_19317,N_18621,N_18694);
and U19318 (N_19318,N_18193,N_18921);
nor U19319 (N_19319,N_18293,N_18556);
xor U19320 (N_19320,N_18995,N_18083);
or U19321 (N_19321,N_18428,N_18480);
nand U19322 (N_19322,N_18842,N_18393);
nand U19323 (N_19323,N_18890,N_18973);
nor U19324 (N_19324,N_18724,N_18384);
nor U19325 (N_19325,N_18738,N_18861);
xor U19326 (N_19326,N_18784,N_18180);
and U19327 (N_19327,N_18586,N_18652);
or U19328 (N_19328,N_18669,N_18711);
xor U19329 (N_19329,N_18877,N_18562);
xor U19330 (N_19330,N_18831,N_18245);
nor U19331 (N_19331,N_18012,N_18403);
nand U19332 (N_19332,N_18491,N_18871);
nor U19333 (N_19333,N_18343,N_18958);
nor U19334 (N_19334,N_18038,N_18218);
xor U19335 (N_19335,N_18665,N_18246);
xnor U19336 (N_19336,N_18406,N_18324);
nand U19337 (N_19337,N_18986,N_18872);
or U19338 (N_19338,N_18696,N_18404);
nor U19339 (N_19339,N_18889,N_18498);
nand U19340 (N_19340,N_18992,N_18096);
nor U19341 (N_19341,N_18883,N_18443);
and U19342 (N_19342,N_18260,N_18098);
nor U19343 (N_19343,N_18353,N_18848);
nor U19344 (N_19344,N_18122,N_18105);
nand U19345 (N_19345,N_18326,N_18277);
or U19346 (N_19346,N_18545,N_18968);
nor U19347 (N_19347,N_18100,N_18547);
and U19348 (N_19348,N_18066,N_18798);
xnor U19349 (N_19349,N_18387,N_18287);
and U19350 (N_19350,N_18638,N_18912);
or U19351 (N_19351,N_18400,N_18820);
nor U19352 (N_19352,N_18876,N_18560);
xor U19353 (N_19353,N_18042,N_18131);
nand U19354 (N_19354,N_18511,N_18003);
nand U19355 (N_19355,N_18079,N_18292);
nand U19356 (N_19356,N_18767,N_18437);
xor U19357 (N_19357,N_18862,N_18262);
xnor U19358 (N_19358,N_18530,N_18487);
xor U19359 (N_19359,N_18596,N_18147);
xnor U19360 (N_19360,N_18152,N_18860);
and U19361 (N_19361,N_18832,N_18744);
nor U19362 (N_19362,N_18846,N_18705);
xor U19363 (N_19363,N_18613,N_18120);
xor U19364 (N_19364,N_18989,N_18394);
xnor U19365 (N_19365,N_18714,N_18199);
nor U19366 (N_19366,N_18505,N_18654);
nor U19367 (N_19367,N_18034,N_18869);
xor U19368 (N_19368,N_18625,N_18346);
and U19369 (N_19369,N_18959,N_18584);
nand U19370 (N_19370,N_18704,N_18226);
xor U19371 (N_19371,N_18977,N_18291);
xnor U19372 (N_19372,N_18266,N_18666);
nor U19373 (N_19373,N_18780,N_18202);
and U19374 (N_19374,N_18983,N_18932);
nand U19375 (N_19375,N_18840,N_18273);
nand U19376 (N_19376,N_18829,N_18138);
xor U19377 (N_19377,N_18089,N_18426);
nor U19378 (N_19378,N_18327,N_18171);
or U19379 (N_19379,N_18591,N_18169);
nand U19380 (N_19380,N_18823,N_18385);
or U19381 (N_19381,N_18015,N_18420);
nor U19382 (N_19382,N_18339,N_18365);
or U19383 (N_19383,N_18880,N_18994);
and U19384 (N_19384,N_18647,N_18763);
xor U19385 (N_19385,N_18775,N_18672);
xor U19386 (N_19386,N_18701,N_18450);
xnor U19387 (N_19387,N_18911,N_18361);
xor U19388 (N_19388,N_18309,N_18068);
nand U19389 (N_19389,N_18229,N_18764);
nand U19390 (N_19390,N_18127,N_18011);
and U19391 (N_19391,N_18330,N_18884);
nand U19392 (N_19392,N_18041,N_18650);
xnor U19393 (N_19393,N_18689,N_18364);
or U19394 (N_19394,N_18252,N_18555);
xnor U19395 (N_19395,N_18614,N_18642);
xor U19396 (N_19396,N_18263,N_18746);
and U19397 (N_19397,N_18206,N_18354);
nand U19398 (N_19398,N_18360,N_18850);
nand U19399 (N_19399,N_18645,N_18103);
or U19400 (N_19400,N_18790,N_18118);
nor U19401 (N_19401,N_18314,N_18002);
nand U19402 (N_19402,N_18212,N_18843);
nand U19403 (N_19403,N_18284,N_18819);
or U19404 (N_19404,N_18358,N_18633);
and U19405 (N_19405,N_18961,N_18785);
or U19406 (N_19406,N_18851,N_18619);
nor U19407 (N_19407,N_18222,N_18425);
xor U19408 (N_19408,N_18146,N_18054);
or U19409 (N_19409,N_18783,N_18071);
nand U19410 (N_19410,N_18946,N_18791);
or U19411 (N_19411,N_18583,N_18976);
or U19412 (N_19412,N_18755,N_18788);
or U19413 (N_19413,N_18678,N_18016);
nand U19414 (N_19414,N_18571,N_18713);
nand U19415 (N_19415,N_18543,N_18722);
or U19416 (N_19416,N_18539,N_18944);
nand U19417 (N_19417,N_18141,N_18013);
nor U19418 (N_19418,N_18230,N_18996);
xnor U19419 (N_19419,N_18163,N_18239);
or U19420 (N_19420,N_18615,N_18858);
nand U19421 (N_19421,N_18756,N_18676);
nand U19422 (N_19422,N_18409,N_18495);
or U19423 (N_19423,N_18168,N_18049);
and U19424 (N_19424,N_18899,N_18727);
nand U19425 (N_19425,N_18907,N_18316);
nor U19426 (N_19426,N_18258,N_18585);
and U19427 (N_19427,N_18679,N_18488);
and U19428 (N_19428,N_18966,N_18806);
or U19429 (N_19429,N_18923,N_18350);
nor U19430 (N_19430,N_18345,N_18005);
nand U19431 (N_19431,N_18770,N_18772);
and U19432 (N_19432,N_18416,N_18997);
nand U19433 (N_19433,N_18133,N_18496);
nand U19434 (N_19434,N_18355,N_18745);
nor U19435 (N_19435,N_18457,N_18208);
or U19436 (N_19436,N_18444,N_18023);
nor U19437 (N_19437,N_18592,N_18139);
xnor U19438 (N_19438,N_18436,N_18815);
nor U19439 (N_19439,N_18134,N_18099);
nand U19440 (N_19440,N_18058,N_18088);
or U19441 (N_19441,N_18969,N_18748);
nand U19442 (N_19442,N_18198,N_18623);
and U19443 (N_19443,N_18663,N_18610);
nor U19444 (N_19444,N_18982,N_18363);
xor U19445 (N_19445,N_18110,N_18257);
and U19446 (N_19446,N_18048,N_18718);
nor U19447 (N_19447,N_18739,N_18506);
xnor U19448 (N_19448,N_18459,N_18975);
nor U19449 (N_19449,N_18549,N_18901);
xnor U19450 (N_19450,N_18325,N_18733);
xor U19451 (N_19451,N_18381,N_18334);
and U19452 (N_19452,N_18472,N_18603);
or U19453 (N_19453,N_18787,N_18866);
nor U19454 (N_19454,N_18512,N_18765);
nand U19455 (N_19455,N_18794,N_18522);
xnor U19456 (N_19456,N_18811,N_18399);
and U19457 (N_19457,N_18939,N_18307);
nand U19458 (N_19458,N_18902,N_18249);
nand U19459 (N_19459,N_18452,N_18455);
or U19460 (N_19460,N_18620,N_18233);
nand U19461 (N_19461,N_18349,N_18627);
and U19462 (N_19462,N_18227,N_18981);
and U19463 (N_19463,N_18818,N_18221);
nand U19464 (N_19464,N_18554,N_18087);
and U19465 (N_19465,N_18677,N_18653);
and U19466 (N_19466,N_18922,N_18464);
or U19467 (N_19467,N_18886,N_18909);
or U19468 (N_19468,N_18735,N_18438);
nor U19469 (N_19469,N_18660,N_18796);
nand U19470 (N_19470,N_18734,N_18344);
and U19471 (N_19471,N_18362,N_18279);
or U19472 (N_19472,N_18140,N_18320);
xor U19473 (N_19473,N_18533,N_18435);
and U19474 (N_19474,N_18340,N_18371);
xnor U19475 (N_19475,N_18352,N_18368);
xor U19476 (N_19476,N_18453,N_18800);
xnor U19477 (N_19477,N_18500,N_18468);
or U19478 (N_19478,N_18323,N_18234);
nor U19479 (N_19479,N_18408,N_18674);
or U19480 (N_19480,N_18520,N_18078);
nor U19481 (N_19481,N_18931,N_18558);
nor U19482 (N_19482,N_18799,N_18113);
xnor U19483 (N_19483,N_18000,N_18685);
or U19484 (N_19484,N_18658,N_18106);
and U19485 (N_19485,N_18289,N_18930);
nor U19486 (N_19486,N_18870,N_18854);
nor U19487 (N_19487,N_18690,N_18026);
xnor U19488 (N_19488,N_18219,N_18329);
or U19489 (N_19489,N_18535,N_18143);
and U19490 (N_19490,N_18954,N_18375);
nor U19491 (N_19491,N_18956,N_18544);
and U19492 (N_19492,N_18517,N_18407);
nor U19493 (N_19493,N_18382,N_18709);
xnor U19494 (N_19494,N_18588,N_18471);
nand U19495 (N_19495,N_18612,N_18839);
nand U19496 (N_19496,N_18618,N_18604);
nand U19497 (N_19497,N_18569,N_18052);
nand U19498 (N_19498,N_18985,N_18205);
nor U19499 (N_19499,N_18313,N_18702);
or U19500 (N_19500,N_18448,N_18267);
and U19501 (N_19501,N_18363,N_18135);
or U19502 (N_19502,N_18549,N_18535);
or U19503 (N_19503,N_18015,N_18258);
and U19504 (N_19504,N_18754,N_18570);
or U19505 (N_19505,N_18966,N_18637);
nor U19506 (N_19506,N_18994,N_18323);
xor U19507 (N_19507,N_18734,N_18858);
and U19508 (N_19508,N_18442,N_18489);
and U19509 (N_19509,N_18849,N_18739);
nor U19510 (N_19510,N_18171,N_18724);
nor U19511 (N_19511,N_18289,N_18809);
nor U19512 (N_19512,N_18401,N_18386);
nand U19513 (N_19513,N_18737,N_18236);
nor U19514 (N_19514,N_18160,N_18709);
nor U19515 (N_19515,N_18591,N_18212);
nor U19516 (N_19516,N_18027,N_18937);
and U19517 (N_19517,N_18946,N_18535);
nor U19518 (N_19518,N_18901,N_18448);
nand U19519 (N_19519,N_18611,N_18185);
xor U19520 (N_19520,N_18236,N_18210);
nor U19521 (N_19521,N_18368,N_18451);
nand U19522 (N_19522,N_18329,N_18393);
xor U19523 (N_19523,N_18596,N_18968);
or U19524 (N_19524,N_18096,N_18259);
nand U19525 (N_19525,N_18751,N_18853);
xor U19526 (N_19526,N_18526,N_18734);
xor U19527 (N_19527,N_18877,N_18090);
nand U19528 (N_19528,N_18017,N_18782);
nand U19529 (N_19529,N_18247,N_18590);
nor U19530 (N_19530,N_18821,N_18500);
or U19531 (N_19531,N_18515,N_18307);
and U19532 (N_19532,N_18726,N_18730);
nand U19533 (N_19533,N_18412,N_18864);
xnor U19534 (N_19534,N_18814,N_18381);
nand U19535 (N_19535,N_18376,N_18704);
and U19536 (N_19536,N_18822,N_18455);
or U19537 (N_19537,N_18854,N_18218);
nand U19538 (N_19538,N_18460,N_18474);
nand U19539 (N_19539,N_18754,N_18372);
and U19540 (N_19540,N_18279,N_18648);
nor U19541 (N_19541,N_18296,N_18515);
and U19542 (N_19542,N_18242,N_18748);
nand U19543 (N_19543,N_18716,N_18638);
and U19544 (N_19544,N_18536,N_18546);
or U19545 (N_19545,N_18799,N_18207);
or U19546 (N_19546,N_18023,N_18647);
nand U19547 (N_19547,N_18175,N_18334);
xor U19548 (N_19548,N_18272,N_18035);
nand U19549 (N_19549,N_18139,N_18188);
and U19550 (N_19550,N_18631,N_18174);
xnor U19551 (N_19551,N_18913,N_18158);
nor U19552 (N_19552,N_18895,N_18102);
nand U19553 (N_19553,N_18903,N_18124);
or U19554 (N_19554,N_18512,N_18397);
and U19555 (N_19555,N_18679,N_18525);
xnor U19556 (N_19556,N_18710,N_18838);
nand U19557 (N_19557,N_18494,N_18136);
xnor U19558 (N_19558,N_18142,N_18573);
nor U19559 (N_19559,N_18428,N_18261);
nand U19560 (N_19560,N_18882,N_18455);
and U19561 (N_19561,N_18299,N_18321);
xor U19562 (N_19562,N_18572,N_18989);
xnor U19563 (N_19563,N_18878,N_18604);
xnor U19564 (N_19564,N_18641,N_18899);
nand U19565 (N_19565,N_18990,N_18128);
and U19566 (N_19566,N_18553,N_18555);
and U19567 (N_19567,N_18094,N_18962);
nand U19568 (N_19568,N_18868,N_18473);
nand U19569 (N_19569,N_18840,N_18006);
nand U19570 (N_19570,N_18055,N_18850);
nand U19571 (N_19571,N_18419,N_18735);
nand U19572 (N_19572,N_18111,N_18564);
nor U19573 (N_19573,N_18378,N_18554);
and U19574 (N_19574,N_18948,N_18857);
nor U19575 (N_19575,N_18368,N_18402);
and U19576 (N_19576,N_18836,N_18456);
xor U19577 (N_19577,N_18170,N_18459);
or U19578 (N_19578,N_18985,N_18750);
nor U19579 (N_19579,N_18612,N_18038);
nand U19580 (N_19580,N_18802,N_18245);
nor U19581 (N_19581,N_18390,N_18534);
nand U19582 (N_19582,N_18968,N_18347);
xnor U19583 (N_19583,N_18802,N_18058);
or U19584 (N_19584,N_18122,N_18417);
nor U19585 (N_19585,N_18606,N_18880);
or U19586 (N_19586,N_18532,N_18443);
nor U19587 (N_19587,N_18833,N_18072);
nand U19588 (N_19588,N_18589,N_18842);
nor U19589 (N_19589,N_18236,N_18086);
nand U19590 (N_19590,N_18079,N_18188);
nor U19591 (N_19591,N_18706,N_18554);
nand U19592 (N_19592,N_18027,N_18399);
or U19593 (N_19593,N_18615,N_18779);
and U19594 (N_19594,N_18228,N_18762);
or U19595 (N_19595,N_18347,N_18503);
xor U19596 (N_19596,N_18351,N_18916);
and U19597 (N_19597,N_18732,N_18115);
nor U19598 (N_19598,N_18908,N_18439);
nor U19599 (N_19599,N_18125,N_18680);
nand U19600 (N_19600,N_18052,N_18959);
or U19601 (N_19601,N_18333,N_18764);
xor U19602 (N_19602,N_18924,N_18070);
xor U19603 (N_19603,N_18771,N_18909);
or U19604 (N_19604,N_18498,N_18557);
and U19605 (N_19605,N_18218,N_18337);
nor U19606 (N_19606,N_18327,N_18095);
xnor U19607 (N_19607,N_18066,N_18122);
or U19608 (N_19608,N_18411,N_18497);
or U19609 (N_19609,N_18343,N_18642);
and U19610 (N_19610,N_18521,N_18500);
or U19611 (N_19611,N_18063,N_18463);
nor U19612 (N_19612,N_18345,N_18459);
nand U19613 (N_19613,N_18759,N_18444);
xnor U19614 (N_19614,N_18826,N_18746);
nand U19615 (N_19615,N_18869,N_18052);
or U19616 (N_19616,N_18772,N_18310);
or U19617 (N_19617,N_18631,N_18745);
or U19618 (N_19618,N_18431,N_18672);
nor U19619 (N_19619,N_18109,N_18478);
and U19620 (N_19620,N_18505,N_18587);
xnor U19621 (N_19621,N_18962,N_18252);
and U19622 (N_19622,N_18476,N_18580);
and U19623 (N_19623,N_18990,N_18505);
and U19624 (N_19624,N_18046,N_18424);
nor U19625 (N_19625,N_18734,N_18452);
or U19626 (N_19626,N_18429,N_18226);
and U19627 (N_19627,N_18950,N_18167);
nand U19628 (N_19628,N_18232,N_18142);
nor U19629 (N_19629,N_18290,N_18238);
and U19630 (N_19630,N_18747,N_18810);
xor U19631 (N_19631,N_18412,N_18029);
nand U19632 (N_19632,N_18648,N_18108);
or U19633 (N_19633,N_18828,N_18210);
nor U19634 (N_19634,N_18090,N_18268);
or U19635 (N_19635,N_18794,N_18031);
xnor U19636 (N_19636,N_18330,N_18416);
nor U19637 (N_19637,N_18520,N_18159);
xor U19638 (N_19638,N_18290,N_18555);
nand U19639 (N_19639,N_18660,N_18685);
xnor U19640 (N_19640,N_18993,N_18695);
and U19641 (N_19641,N_18093,N_18275);
xnor U19642 (N_19642,N_18265,N_18495);
and U19643 (N_19643,N_18641,N_18382);
xnor U19644 (N_19644,N_18591,N_18720);
and U19645 (N_19645,N_18646,N_18364);
and U19646 (N_19646,N_18988,N_18318);
and U19647 (N_19647,N_18186,N_18346);
nor U19648 (N_19648,N_18155,N_18449);
and U19649 (N_19649,N_18770,N_18882);
or U19650 (N_19650,N_18255,N_18713);
nand U19651 (N_19651,N_18440,N_18524);
nor U19652 (N_19652,N_18784,N_18271);
nand U19653 (N_19653,N_18147,N_18090);
or U19654 (N_19654,N_18079,N_18973);
or U19655 (N_19655,N_18136,N_18232);
nand U19656 (N_19656,N_18759,N_18770);
and U19657 (N_19657,N_18276,N_18382);
and U19658 (N_19658,N_18147,N_18468);
nand U19659 (N_19659,N_18351,N_18532);
xor U19660 (N_19660,N_18214,N_18662);
or U19661 (N_19661,N_18461,N_18027);
or U19662 (N_19662,N_18173,N_18790);
xor U19663 (N_19663,N_18077,N_18544);
nand U19664 (N_19664,N_18811,N_18845);
or U19665 (N_19665,N_18451,N_18138);
nor U19666 (N_19666,N_18492,N_18354);
nand U19667 (N_19667,N_18074,N_18374);
and U19668 (N_19668,N_18067,N_18724);
nor U19669 (N_19669,N_18935,N_18448);
or U19670 (N_19670,N_18166,N_18786);
xor U19671 (N_19671,N_18850,N_18147);
xor U19672 (N_19672,N_18706,N_18518);
nand U19673 (N_19673,N_18386,N_18468);
nor U19674 (N_19674,N_18878,N_18584);
nand U19675 (N_19675,N_18282,N_18934);
or U19676 (N_19676,N_18488,N_18729);
and U19677 (N_19677,N_18027,N_18872);
or U19678 (N_19678,N_18550,N_18760);
and U19679 (N_19679,N_18921,N_18876);
xor U19680 (N_19680,N_18377,N_18771);
xnor U19681 (N_19681,N_18467,N_18140);
or U19682 (N_19682,N_18105,N_18891);
nor U19683 (N_19683,N_18852,N_18425);
or U19684 (N_19684,N_18811,N_18269);
nor U19685 (N_19685,N_18442,N_18073);
or U19686 (N_19686,N_18230,N_18558);
or U19687 (N_19687,N_18769,N_18936);
and U19688 (N_19688,N_18625,N_18168);
nor U19689 (N_19689,N_18833,N_18061);
or U19690 (N_19690,N_18026,N_18201);
and U19691 (N_19691,N_18006,N_18090);
xnor U19692 (N_19692,N_18447,N_18181);
xor U19693 (N_19693,N_18118,N_18070);
or U19694 (N_19694,N_18916,N_18387);
xor U19695 (N_19695,N_18356,N_18537);
and U19696 (N_19696,N_18841,N_18084);
xor U19697 (N_19697,N_18505,N_18669);
nor U19698 (N_19698,N_18151,N_18366);
and U19699 (N_19699,N_18645,N_18660);
nor U19700 (N_19700,N_18456,N_18775);
and U19701 (N_19701,N_18116,N_18940);
or U19702 (N_19702,N_18361,N_18602);
or U19703 (N_19703,N_18117,N_18966);
xnor U19704 (N_19704,N_18023,N_18920);
nor U19705 (N_19705,N_18818,N_18176);
or U19706 (N_19706,N_18867,N_18963);
nand U19707 (N_19707,N_18413,N_18434);
nand U19708 (N_19708,N_18613,N_18867);
nor U19709 (N_19709,N_18164,N_18619);
nor U19710 (N_19710,N_18610,N_18175);
nor U19711 (N_19711,N_18066,N_18608);
and U19712 (N_19712,N_18474,N_18696);
and U19713 (N_19713,N_18912,N_18714);
or U19714 (N_19714,N_18944,N_18381);
and U19715 (N_19715,N_18068,N_18067);
nor U19716 (N_19716,N_18157,N_18143);
and U19717 (N_19717,N_18791,N_18248);
xor U19718 (N_19718,N_18223,N_18494);
xor U19719 (N_19719,N_18230,N_18138);
or U19720 (N_19720,N_18986,N_18326);
nand U19721 (N_19721,N_18630,N_18619);
nor U19722 (N_19722,N_18157,N_18378);
or U19723 (N_19723,N_18727,N_18654);
nand U19724 (N_19724,N_18304,N_18582);
nand U19725 (N_19725,N_18805,N_18797);
nand U19726 (N_19726,N_18632,N_18727);
nand U19727 (N_19727,N_18853,N_18363);
and U19728 (N_19728,N_18645,N_18860);
and U19729 (N_19729,N_18856,N_18994);
nor U19730 (N_19730,N_18857,N_18847);
nand U19731 (N_19731,N_18155,N_18139);
nor U19732 (N_19732,N_18816,N_18638);
and U19733 (N_19733,N_18315,N_18547);
nand U19734 (N_19734,N_18521,N_18558);
or U19735 (N_19735,N_18306,N_18265);
xnor U19736 (N_19736,N_18526,N_18920);
or U19737 (N_19737,N_18938,N_18454);
or U19738 (N_19738,N_18485,N_18626);
and U19739 (N_19739,N_18303,N_18444);
and U19740 (N_19740,N_18705,N_18618);
and U19741 (N_19741,N_18732,N_18683);
nor U19742 (N_19742,N_18674,N_18577);
and U19743 (N_19743,N_18036,N_18678);
and U19744 (N_19744,N_18922,N_18927);
and U19745 (N_19745,N_18825,N_18885);
and U19746 (N_19746,N_18042,N_18136);
or U19747 (N_19747,N_18332,N_18051);
xnor U19748 (N_19748,N_18966,N_18448);
nor U19749 (N_19749,N_18163,N_18484);
and U19750 (N_19750,N_18134,N_18914);
or U19751 (N_19751,N_18884,N_18418);
and U19752 (N_19752,N_18236,N_18828);
or U19753 (N_19753,N_18275,N_18060);
nor U19754 (N_19754,N_18863,N_18452);
nand U19755 (N_19755,N_18143,N_18932);
and U19756 (N_19756,N_18182,N_18897);
xnor U19757 (N_19757,N_18584,N_18557);
and U19758 (N_19758,N_18701,N_18648);
or U19759 (N_19759,N_18590,N_18388);
nand U19760 (N_19760,N_18328,N_18484);
xnor U19761 (N_19761,N_18204,N_18781);
nand U19762 (N_19762,N_18716,N_18762);
nand U19763 (N_19763,N_18702,N_18145);
and U19764 (N_19764,N_18568,N_18144);
xor U19765 (N_19765,N_18088,N_18533);
or U19766 (N_19766,N_18393,N_18820);
nor U19767 (N_19767,N_18057,N_18031);
nand U19768 (N_19768,N_18205,N_18125);
nand U19769 (N_19769,N_18366,N_18317);
or U19770 (N_19770,N_18482,N_18350);
and U19771 (N_19771,N_18185,N_18294);
and U19772 (N_19772,N_18450,N_18213);
xnor U19773 (N_19773,N_18915,N_18621);
xnor U19774 (N_19774,N_18457,N_18986);
nor U19775 (N_19775,N_18078,N_18721);
nor U19776 (N_19776,N_18064,N_18897);
nor U19777 (N_19777,N_18336,N_18261);
nor U19778 (N_19778,N_18988,N_18759);
and U19779 (N_19779,N_18188,N_18050);
nand U19780 (N_19780,N_18200,N_18161);
and U19781 (N_19781,N_18633,N_18385);
nand U19782 (N_19782,N_18484,N_18910);
nor U19783 (N_19783,N_18819,N_18026);
nand U19784 (N_19784,N_18140,N_18530);
nor U19785 (N_19785,N_18052,N_18058);
and U19786 (N_19786,N_18340,N_18708);
or U19787 (N_19787,N_18520,N_18614);
nand U19788 (N_19788,N_18336,N_18659);
nor U19789 (N_19789,N_18979,N_18487);
or U19790 (N_19790,N_18357,N_18977);
nor U19791 (N_19791,N_18190,N_18166);
xor U19792 (N_19792,N_18788,N_18838);
nand U19793 (N_19793,N_18909,N_18114);
and U19794 (N_19794,N_18435,N_18626);
nor U19795 (N_19795,N_18876,N_18472);
and U19796 (N_19796,N_18640,N_18635);
and U19797 (N_19797,N_18391,N_18790);
xnor U19798 (N_19798,N_18832,N_18988);
xor U19799 (N_19799,N_18426,N_18966);
and U19800 (N_19800,N_18899,N_18274);
xor U19801 (N_19801,N_18611,N_18670);
or U19802 (N_19802,N_18519,N_18122);
nand U19803 (N_19803,N_18205,N_18269);
xor U19804 (N_19804,N_18630,N_18213);
xor U19805 (N_19805,N_18741,N_18695);
nand U19806 (N_19806,N_18819,N_18987);
or U19807 (N_19807,N_18813,N_18090);
nand U19808 (N_19808,N_18877,N_18872);
nand U19809 (N_19809,N_18932,N_18785);
nor U19810 (N_19810,N_18419,N_18791);
and U19811 (N_19811,N_18418,N_18986);
or U19812 (N_19812,N_18367,N_18109);
and U19813 (N_19813,N_18722,N_18507);
xor U19814 (N_19814,N_18583,N_18688);
xor U19815 (N_19815,N_18714,N_18393);
nand U19816 (N_19816,N_18124,N_18797);
nand U19817 (N_19817,N_18085,N_18697);
or U19818 (N_19818,N_18620,N_18569);
and U19819 (N_19819,N_18691,N_18206);
nand U19820 (N_19820,N_18712,N_18668);
xnor U19821 (N_19821,N_18624,N_18459);
xnor U19822 (N_19822,N_18035,N_18770);
or U19823 (N_19823,N_18205,N_18560);
and U19824 (N_19824,N_18404,N_18623);
xor U19825 (N_19825,N_18311,N_18992);
nor U19826 (N_19826,N_18606,N_18618);
xnor U19827 (N_19827,N_18218,N_18871);
and U19828 (N_19828,N_18478,N_18305);
or U19829 (N_19829,N_18175,N_18785);
or U19830 (N_19830,N_18630,N_18880);
xnor U19831 (N_19831,N_18239,N_18994);
nand U19832 (N_19832,N_18677,N_18035);
nand U19833 (N_19833,N_18562,N_18535);
xor U19834 (N_19834,N_18228,N_18943);
xor U19835 (N_19835,N_18715,N_18156);
xnor U19836 (N_19836,N_18227,N_18718);
or U19837 (N_19837,N_18613,N_18955);
xnor U19838 (N_19838,N_18108,N_18150);
or U19839 (N_19839,N_18718,N_18824);
xnor U19840 (N_19840,N_18719,N_18066);
nand U19841 (N_19841,N_18287,N_18641);
or U19842 (N_19842,N_18965,N_18422);
and U19843 (N_19843,N_18964,N_18968);
or U19844 (N_19844,N_18228,N_18803);
and U19845 (N_19845,N_18062,N_18767);
and U19846 (N_19846,N_18064,N_18262);
nand U19847 (N_19847,N_18850,N_18437);
or U19848 (N_19848,N_18867,N_18115);
nand U19849 (N_19849,N_18745,N_18983);
xnor U19850 (N_19850,N_18349,N_18644);
xor U19851 (N_19851,N_18969,N_18371);
and U19852 (N_19852,N_18596,N_18935);
and U19853 (N_19853,N_18594,N_18798);
xnor U19854 (N_19854,N_18748,N_18186);
or U19855 (N_19855,N_18997,N_18074);
nor U19856 (N_19856,N_18739,N_18233);
or U19857 (N_19857,N_18230,N_18473);
nor U19858 (N_19858,N_18521,N_18051);
xor U19859 (N_19859,N_18582,N_18136);
nand U19860 (N_19860,N_18162,N_18196);
nand U19861 (N_19861,N_18407,N_18065);
and U19862 (N_19862,N_18654,N_18739);
or U19863 (N_19863,N_18852,N_18511);
nand U19864 (N_19864,N_18253,N_18510);
and U19865 (N_19865,N_18969,N_18352);
nand U19866 (N_19866,N_18458,N_18791);
nor U19867 (N_19867,N_18682,N_18444);
or U19868 (N_19868,N_18074,N_18127);
or U19869 (N_19869,N_18707,N_18146);
and U19870 (N_19870,N_18569,N_18049);
and U19871 (N_19871,N_18914,N_18236);
and U19872 (N_19872,N_18569,N_18629);
and U19873 (N_19873,N_18847,N_18235);
nor U19874 (N_19874,N_18362,N_18883);
xnor U19875 (N_19875,N_18733,N_18018);
nor U19876 (N_19876,N_18824,N_18116);
nand U19877 (N_19877,N_18670,N_18762);
nor U19878 (N_19878,N_18742,N_18188);
and U19879 (N_19879,N_18899,N_18843);
xor U19880 (N_19880,N_18662,N_18929);
and U19881 (N_19881,N_18185,N_18064);
or U19882 (N_19882,N_18703,N_18486);
and U19883 (N_19883,N_18131,N_18714);
xor U19884 (N_19884,N_18244,N_18831);
nand U19885 (N_19885,N_18678,N_18181);
nor U19886 (N_19886,N_18413,N_18347);
or U19887 (N_19887,N_18805,N_18403);
nor U19888 (N_19888,N_18603,N_18136);
nand U19889 (N_19889,N_18985,N_18805);
xnor U19890 (N_19890,N_18192,N_18298);
nor U19891 (N_19891,N_18079,N_18126);
nor U19892 (N_19892,N_18468,N_18501);
nor U19893 (N_19893,N_18384,N_18326);
nor U19894 (N_19894,N_18364,N_18136);
and U19895 (N_19895,N_18666,N_18417);
nor U19896 (N_19896,N_18846,N_18750);
or U19897 (N_19897,N_18707,N_18561);
xor U19898 (N_19898,N_18276,N_18022);
nand U19899 (N_19899,N_18388,N_18539);
nand U19900 (N_19900,N_18836,N_18294);
xor U19901 (N_19901,N_18617,N_18430);
nor U19902 (N_19902,N_18894,N_18034);
or U19903 (N_19903,N_18241,N_18534);
xor U19904 (N_19904,N_18963,N_18492);
xor U19905 (N_19905,N_18948,N_18716);
xnor U19906 (N_19906,N_18877,N_18328);
xnor U19907 (N_19907,N_18752,N_18100);
xnor U19908 (N_19908,N_18563,N_18289);
nor U19909 (N_19909,N_18527,N_18300);
xor U19910 (N_19910,N_18745,N_18350);
xnor U19911 (N_19911,N_18407,N_18040);
nor U19912 (N_19912,N_18689,N_18496);
nor U19913 (N_19913,N_18227,N_18338);
or U19914 (N_19914,N_18283,N_18441);
and U19915 (N_19915,N_18206,N_18922);
or U19916 (N_19916,N_18568,N_18267);
and U19917 (N_19917,N_18899,N_18278);
xnor U19918 (N_19918,N_18817,N_18905);
and U19919 (N_19919,N_18675,N_18474);
nor U19920 (N_19920,N_18253,N_18570);
xor U19921 (N_19921,N_18412,N_18333);
and U19922 (N_19922,N_18146,N_18831);
and U19923 (N_19923,N_18090,N_18063);
and U19924 (N_19924,N_18750,N_18004);
and U19925 (N_19925,N_18141,N_18627);
or U19926 (N_19926,N_18343,N_18415);
xnor U19927 (N_19927,N_18017,N_18616);
and U19928 (N_19928,N_18705,N_18802);
and U19929 (N_19929,N_18979,N_18363);
nand U19930 (N_19930,N_18435,N_18619);
and U19931 (N_19931,N_18045,N_18558);
or U19932 (N_19932,N_18953,N_18115);
and U19933 (N_19933,N_18022,N_18369);
xnor U19934 (N_19934,N_18830,N_18344);
nor U19935 (N_19935,N_18652,N_18566);
and U19936 (N_19936,N_18831,N_18110);
nand U19937 (N_19937,N_18172,N_18532);
and U19938 (N_19938,N_18835,N_18360);
xor U19939 (N_19939,N_18452,N_18266);
xor U19940 (N_19940,N_18913,N_18650);
or U19941 (N_19941,N_18180,N_18400);
or U19942 (N_19942,N_18388,N_18879);
and U19943 (N_19943,N_18637,N_18917);
nand U19944 (N_19944,N_18803,N_18367);
nor U19945 (N_19945,N_18107,N_18401);
and U19946 (N_19946,N_18509,N_18264);
and U19947 (N_19947,N_18798,N_18384);
nand U19948 (N_19948,N_18347,N_18564);
xor U19949 (N_19949,N_18065,N_18797);
or U19950 (N_19950,N_18335,N_18325);
nand U19951 (N_19951,N_18509,N_18098);
or U19952 (N_19952,N_18657,N_18010);
nand U19953 (N_19953,N_18348,N_18593);
or U19954 (N_19954,N_18772,N_18059);
nor U19955 (N_19955,N_18698,N_18057);
and U19956 (N_19956,N_18889,N_18693);
nand U19957 (N_19957,N_18155,N_18812);
nor U19958 (N_19958,N_18565,N_18064);
and U19959 (N_19959,N_18159,N_18010);
xnor U19960 (N_19960,N_18815,N_18615);
and U19961 (N_19961,N_18853,N_18356);
nor U19962 (N_19962,N_18601,N_18724);
or U19963 (N_19963,N_18832,N_18368);
nor U19964 (N_19964,N_18090,N_18012);
or U19965 (N_19965,N_18973,N_18907);
and U19966 (N_19966,N_18083,N_18414);
and U19967 (N_19967,N_18903,N_18358);
nor U19968 (N_19968,N_18072,N_18972);
xor U19969 (N_19969,N_18924,N_18430);
nor U19970 (N_19970,N_18685,N_18762);
xor U19971 (N_19971,N_18394,N_18914);
and U19972 (N_19972,N_18154,N_18839);
or U19973 (N_19973,N_18864,N_18031);
and U19974 (N_19974,N_18824,N_18996);
and U19975 (N_19975,N_18680,N_18144);
nor U19976 (N_19976,N_18279,N_18897);
and U19977 (N_19977,N_18624,N_18599);
xnor U19978 (N_19978,N_18842,N_18060);
nor U19979 (N_19979,N_18592,N_18246);
nand U19980 (N_19980,N_18153,N_18267);
nand U19981 (N_19981,N_18057,N_18916);
nor U19982 (N_19982,N_18913,N_18488);
and U19983 (N_19983,N_18510,N_18162);
nand U19984 (N_19984,N_18011,N_18000);
or U19985 (N_19985,N_18049,N_18947);
nor U19986 (N_19986,N_18682,N_18508);
or U19987 (N_19987,N_18055,N_18624);
xnor U19988 (N_19988,N_18809,N_18539);
xor U19989 (N_19989,N_18816,N_18064);
or U19990 (N_19990,N_18553,N_18160);
nor U19991 (N_19991,N_18917,N_18092);
nand U19992 (N_19992,N_18106,N_18260);
nor U19993 (N_19993,N_18455,N_18684);
nor U19994 (N_19994,N_18584,N_18271);
nor U19995 (N_19995,N_18557,N_18836);
nand U19996 (N_19996,N_18239,N_18609);
or U19997 (N_19997,N_18760,N_18394);
and U19998 (N_19998,N_18614,N_18454);
nand U19999 (N_19999,N_18824,N_18572);
or U20000 (N_20000,N_19588,N_19256);
xnor U20001 (N_20001,N_19883,N_19103);
and U20002 (N_20002,N_19468,N_19593);
and U20003 (N_20003,N_19381,N_19773);
or U20004 (N_20004,N_19957,N_19142);
nand U20005 (N_20005,N_19411,N_19535);
xor U20006 (N_20006,N_19393,N_19796);
or U20007 (N_20007,N_19286,N_19722);
xnor U20008 (N_20008,N_19960,N_19230);
nor U20009 (N_20009,N_19565,N_19191);
xor U20010 (N_20010,N_19457,N_19017);
or U20011 (N_20011,N_19463,N_19047);
nand U20012 (N_20012,N_19113,N_19741);
or U20013 (N_20013,N_19440,N_19476);
xor U20014 (N_20014,N_19136,N_19895);
and U20015 (N_20015,N_19231,N_19543);
nor U20016 (N_20016,N_19108,N_19707);
xor U20017 (N_20017,N_19687,N_19786);
and U20018 (N_20018,N_19644,N_19257);
or U20019 (N_20019,N_19331,N_19522);
and U20020 (N_20020,N_19268,N_19979);
nand U20021 (N_20021,N_19408,N_19653);
and U20022 (N_20022,N_19672,N_19985);
nand U20023 (N_20023,N_19812,N_19569);
and U20024 (N_20024,N_19594,N_19726);
and U20025 (N_20025,N_19209,N_19474);
nor U20026 (N_20026,N_19157,N_19838);
or U20027 (N_20027,N_19616,N_19458);
xor U20028 (N_20028,N_19785,N_19184);
or U20029 (N_20029,N_19928,N_19844);
xnor U20030 (N_20030,N_19898,N_19533);
xor U20031 (N_20031,N_19831,N_19098);
and U20032 (N_20032,N_19161,N_19443);
xor U20033 (N_20033,N_19480,N_19076);
xnor U20034 (N_20034,N_19878,N_19822);
nor U20035 (N_20035,N_19996,N_19348);
xor U20036 (N_20036,N_19228,N_19328);
and U20037 (N_20037,N_19704,N_19832);
and U20038 (N_20038,N_19819,N_19206);
nor U20039 (N_20039,N_19573,N_19825);
xnor U20040 (N_20040,N_19524,N_19399);
and U20041 (N_20041,N_19173,N_19225);
and U20042 (N_20042,N_19974,N_19767);
nand U20043 (N_20043,N_19969,N_19905);
and U20044 (N_20044,N_19506,N_19043);
and U20045 (N_20045,N_19787,N_19032);
or U20046 (N_20046,N_19788,N_19077);
and U20047 (N_20047,N_19038,N_19249);
and U20048 (N_20048,N_19770,N_19659);
xnor U20049 (N_20049,N_19083,N_19920);
nand U20050 (N_20050,N_19530,N_19336);
and U20051 (N_20051,N_19299,N_19681);
nand U20052 (N_20052,N_19536,N_19948);
and U20053 (N_20053,N_19337,N_19045);
and U20054 (N_20054,N_19246,N_19298);
or U20055 (N_20055,N_19149,N_19266);
xnor U20056 (N_20056,N_19833,N_19310);
or U20057 (N_20057,N_19454,N_19532);
nor U20058 (N_20058,N_19224,N_19664);
or U20059 (N_20059,N_19547,N_19714);
xor U20060 (N_20060,N_19194,N_19489);
xnor U20061 (N_20061,N_19860,N_19708);
nand U20062 (N_20062,N_19074,N_19188);
or U20063 (N_20063,N_19315,N_19226);
or U20064 (N_20064,N_19586,N_19003);
and U20065 (N_20065,N_19768,N_19596);
nor U20066 (N_20066,N_19159,N_19362);
and U20067 (N_20067,N_19564,N_19295);
nor U20068 (N_20068,N_19144,N_19733);
xor U20069 (N_20069,N_19061,N_19439);
nand U20070 (N_20070,N_19863,N_19452);
nand U20071 (N_20071,N_19575,N_19420);
nand U20072 (N_20072,N_19124,N_19134);
nor U20073 (N_20073,N_19202,N_19683);
nand U20074 (N_20074,N_19738,N_19684);
nor U20075 (N_20075,N_19650,N_19654);
nor U20076 (N_20076,N_19637,N_19732);
and U20077 (N_20077,N_19952,N_19875);
nand U20078 (N_20078,N_19538,N_19027);
xnor U20079 (N_20079,N_19438,N_19419);
nor U20080 (N_20080,N_19783,N_19235);
or U20081 (N_20081,N_19418,N_19303);
and U20082 (N_20082,N_19021,N_19668);
nand U20083 (N_20083,N_19401,N_19431);
or U20084 (N_20084,N_19484,N_19917);
nand U20085 (N_20085,N_19250,N_19006);
xor U20086 (N_20086,N_19599,N_19265);
nand U20087 (N_20087,N_19873,N_19175);
or U20088 (N_20088,N_19389,N_19070);
nand U20089 (N_20089,N_19504,N_19436);
or U20090 (N_20090,N_19065,N_19060);
or U20091 (N_20091,N_19936,N_19550);
and U20092 (N_20092,N_19571,N_19459);
nand U20093 (N_20093,N_19079,N_19828);
nand U20094 (N_20094,N_19754,N_19020);
xnor U20095 (N_20095,N_19433,N_19397);
nand U20096 (N_20096,N_19182,N_19180);
nor U20097 (N_20097,N_19485,N_19271);
nand U20098 (N_20098,N_19217,N_19035);
nor U20099 (N_20099,N_19329,N_19642);
xor U20100 (N_20100,N_19574,N_19585);
or U20101 (N_20101,N_19958,N_19730);
or U20102 (N_20102,N_19261,N_19369);
nor U20103 (N_20103,N_19667,N_19498);
xor U20104 (N_20104,N_19848,N_19041);
nor U20105 (N_20105,N_19053,N_19676);
nor U20106 (N_20106,N_19197,N_19992);
nand U20107 (N_20107,N_19198,N_19404);
or U20108 (N_20108,N_19717,N_19647);
or U20109 (N_20109,N_19201,N_19203);
xor U20110 (N_20110,N_19758,N_19744);
nor U20111 (N_20111,N_19379,N_19423);
xor U20112 (N_20112,N_19253,N_19497);
or U20113 (N_20113,N_19284,N_19777);
nand U20114 (N_20114,N_19410,N_19674);
and U20115 (N_20115,N_19008,N_19709);
and U20116 (N_20116,N_19264,N_19131);
and U20117 (N_20117,N_19950,N_19772);
and U20118 (N_20118,N_19229,N_19115);
or U20119 (N_20119,N_19743,N_19220);
and U20120 (N_20120,N_19304,N_19472);
nand U20121 (N_20121,N_19534,N_19449);
xor U20122 (N_20122,N_19340,N_19789);
nand U20123 (N_20123,N_19267,N_19486);
and U20124 (N_20124,N_19057,N_19857);
nor U20125 (N_20125,N_19673,N_19806);
nand U20126 (N_20126,N_19523,N_19214);
or U20127 (N_20127,N_19631,N_19495);
nor U20128 (N_20128,N_19697,N_19502);
and U20129 (N_20129,N_19364,N_19002);
and U20130 (N_20130,N_19211,N_19291);
nand U20131 (N_20131,N_19482,N_19924);
nand U20132 (N_20132,N_19123,N_19510);
and U20133 (N_20133,N_19769,N_19207);
nor U20134 (N_20134,N_19196,N_19890);
or U20135 (N_20135,N_19091,N_19368);
and U20136 (N_20136,N_19398,N_19749);
or U20137 (N_20137,N_19839,N_19519);
or U20138 (N_20138,N_19849,N_19407);
nor U20139 (N_20139,N_19488,N_19039);
and U20140 (N_20140,N_19973,N_19372);
xnor U20141 (N_20141,N_19375,N_19186);
nor U20142 (N_20142,N_19395,N_19911);
or U20143 (N_20143,N_19162,N_19881);
nor U20144 (N_20144,N_19814,N_19701);
nor U20145 (N_20145,N_19613,N_19170);
or U20146 (N_20146,N_19311,N_19174);
nand U20147 (N_20147,N_19711,N_19560);
nor U20148 (N_20148,N_19199,N_19932);
nor U20149 (N_20149,N_19894,N_19269);
and U20150 (N_20150,N_19169,N_19827);
and U20151 (N_20151,N_19645,N_19023);
and U20152 (N_20152,N_19998,N_19804);
nor U20153 (N_20153,N_19809,N_19470);
or U20154 (N_20154,N_19102,N_19260);
and U20155 (N_20155,N_19568,N_19289);
nor U20156 (N_20156,N_19651,N_19349);
nand U20157 (N_20157,N_19048,N_19661);
xnor U20158 (N_20158,N_19556,N_19791);
and U20159 (N_20159,N_19344,N_19602);
or U20160 (N_20160,N_19273,N_19515);
and U20161 (N_20161,N_19778,N_19137);
nor U20162 (N_20162,N_19902,N_19012);
xnor U20163 (N_20163,N_19988,N_19578);
or U20164 (N_20164,N_19652,N_19429);
xor U20165 (N_20165,N_19354,N_19852);
nand U20166 (N_20166,N_19531,N_19109);
xnor U20167 (N_20167,N_19447,N_19846);
nor U20168 (N_20168,N_19824,N_19409);
and U20169 (N_20169,N_19633,N_19384);
nor U20170 (N_20170,N_19031,N_19628);
and U20171 (N_20171,N_19634,N_19858);
and U20172 (N_20172,N_19346,N_19305);
xor U20173 (N_20173,N_19500,N_19587);
xnor U20174 (N_20174,N_19887,N_19183);
nand U20175 (N_20175,N_19855,N_19294);
and U20176 (N_20176,N_19723,N_19323);
nand U20177 (N_20177,N_19830,N_19318);
or U20178 (N_20178,N_19623,N_19870);
and U20179 (N_20179,N_19528,N_19636);
nand U20180 (N_20180,N_19278,N_19581);
or U20181 (N_20181,N_19916,N_19949);
xor U20182 (N_20182,N_19927,N_19914);
xor U20183 (N_20183,N_19835,N_19425);
and U20184 (N_20184,N_19312,N_19945);
xnor U20185 (N_20185,N_19513,N_19105);
nand U20186 (N_20186,N_19682,N_19826);
xnor U20187 (N_20187,N_19559,N_19876);
nand U20188 (N_20188,N_19234,N_19277);
or U20189 (N_20189,N_19984,N_19189);
or U20190 (N_20190,N_19866,N_19096);
xor U20191 (N_20191,N_19242,N_19583);
nand U20192 (N_20192,N_19748,N_19499);
or U20193 (N_20193,N_19141,N_19370);
nand U20194 (N_20194,N_19288,N_19233);
and U20195 (N_20195,N_19491,N_19241);
nor U20196 (N_20196,N_19387,N_19243);
xnor U20197 (N_20197,N_19615,N_19118);
xor U20198 (N_20198,N_19412,N_19545);
and U20199 (N_20199,N_19516,N_19563);
nor U20200 (N_20200,N_19200,N_19094);
or U20201 (N_20201,N_19837,N_19308);
and U20202 (N_20202,N_19662,N_19084);
nand U20203 (N_20203,N_19448,N_19656);
nor U20204 (N_20204,N_19475,N_19823);
or U20205 (N_20205,N_19710,N_19301);
xnor U20206 (N_20206,N_19821,N_19549);
nor U20207 (N_20207,N_19293,N_19872);
or U20208 (N_20208,N_19167,N_19403);
xnor U20209 (N_20209,N_19817,N_19861);
nor U20210 (N_20210,N_19319,N_19970);
and U20211 (N_20211,N_19841,N_19867);
xnor U20212 (N_20212,N_19630,N_19981);
xnor U20213 (N_20213,N_19376,N_19263);
and U20214 (N_20214,N_19363,N_19120);
nor U20215 (N_20215,N_19158,N_19781);
nor U20216 (N_20216,N_19054,N_19068);
or U20217 (N_20217,N_19238,N_19993);
or U20218 (N_20218,N_19223,N_19465);
and U20219 (N_20219,N_19392,N_19051);
nand U20220 (N_20220,N_19147,N_19705);
or U20221 (N_20221,N_19956,N_19089);
or U20222 (N_20222,N_19320,N_19925);
or U20223 (N_20223,N_19192,N_19893);
nand U20224 (N_20224,N_19753,N_19582);
nand U20225 (N_20225,N_19334,N_19601);
xor U20226 (N_20226,N_19739,N_19978);
nor U20227 (N_20227,N_19737,N_19059);
nand U20228 (N_20228,N_19111,N_19171);
nor U20229 (N_20229,N_19024,N_19605);
xor U20230 (N_20230,N_19736,N_19450);
nand U20231 (N_20231,N_19889,N_19001);
nand U20232 (N_20232,N_19390,N_19374);
xnor U20233 (N_20233,N_19731,N_19658);
or U20234 (N_20234,N_19212,N_19544);
or U20235 (N_20235,N_19942,N_19641);
nor U20236 (N_20236,N_19521,N_19721);
nand U20237 (N_20237,N_19897,N_19750);
and U20238 (N_20238,N_19280,N_19620);
or U20239 (N_20239,N_19155,N_19501);
nand U20240 (N_20240,N_19900,N_19481);
and U20241 (N_20241,N_19466,N_19845);
or U20242 (N_20242,N_19116,N_19324);
nand U20243 (N_20243,N_19671,N_19555);
and U20244 (N_20244,N_19944,N_19316);
or U20245 (N_20245,N_19720,N_19082);
nor U20246 (N_20246,N_19446,N_19614);
nor U20247 (N_20247,N_19918,N_19529);
and U20248 (N_20248,N_19135,N_19326);
nand U20249 (N_20249,N_19665,N_19509);
nand U20250 (N_20250,N_19980,N_19908);
nor U20251 (N_20251,N_19891,N_19526);
xnor U20252 (N_20252,N_19332,N_19871);
nor U20253 (N_20253,N_19757,N_19240);
or U20254 (N_20254,N_19907,N_19762);
nor U20255 (N_20255,N_19455,N_19740);
xor U20256 (N_20256,N_19570,N_19025);
or U20257 (N_20257,N_19385,N_19239);
or U20258 (N_20258,N_19805,N_19081);
nor U20259 (N_20259,N_19297,N_19760);
xor U20260 (N_20260,N_19343,N_19690);
and U20261 (N_20261,N_19540,N_19358);
or U20262 (N_20262,N_19371,N_19551);
nor U20263 (N_20263,N_19909,N_19702);
xor U20264 (N_20264,N_19735,N_19270);
and U20265 (N_20265,N_19745,N_19910);
and U20266 (N_20266,N_19421,N_19706);
xor U20267 (N_20267,N_19546,N_19864);
nand U20268 (N_20268,N_19983,N_19276);
and U20269 (N_20269,N_19355,N_19365);
xor U20270 (N_20270,N_19215,N_19462);
or U20271 (N_20271,N_19935,N_19700);
xor U20272 (N_20272,N_19929,N_19179);
xnor U20273 (N_20273,N_19037,N_19727);
and U20274 (N_20274,N_19107,N_19255);
nand U20275 (N_20275,N_19367,N_19566);
xnor U20276 (N_20276,N_19353,N_19473);
nand U20277 (N_20277,N_19680,N_19085);
or U20278 (N_20278,N_19177,N_19520);
or U20279 (N_20279,N_19989,N_19906);
or U20280 (N_20280,N_19606,N_19595);
nor U20281 (N_20281,N_19558,N_19675);
or U20282 (N_20282,N_19285,N_19766);
nand U20283 (N_20283,N_19213,N_19759);
nand U20284 (N_20284,N_19281,N_19442);
or U20285 (N_20285,N_19487,N_19210);
or U20286 (N_20286,N_19921,N_19496);
xor U20287 (N_20287,N_19232,N_19087);
nand U20288 (N_20288,N_19029,N_19287);
nand U20289 (N_20289,N_19435,N_19150);
nor U20290 (N_20290,N_19193,N_19525);
and U20291 (N_20291,N_19703,N_19933);
or U20292 (N_20292,N_19884,N_19148);
nor U20293 (N_20293,N_19512,N_19597);
and U20294 (N_20294,N_19152,N_19899);
xor U20295 (N_20295,N_19959,N_19800);
nand U20296 (N_20296,N_19306,N_19430);
and U20297 (N_20297,N_19548,N_19943);
and U20298 (N_20298,N_19880,N_19040);
or U20299 (N_20299,N_19274,N_19632);
and U20300 (N_20300,N_19492,N_19716);
or U20301 (N_20301,N_19811,N_19694);
and U20302 (N_20302,N_19790,N_19624);
or U20303 (N_20303,N_19460,N_19869);
and U20304 (N_20304,N_19483,N_19112);
and U20305 (N_20305,N_19254,N_19129);
and U20306 (N_20306,N_19154,N_19046);
nor U20307 (N_20307,N_19127,N_19009);
and U20308 (N_20308,N_19090,N_19792);
or U20309 (N_20309,N_19527,N_19874);
and U20310 (N_20310,N_19479,N_19850);
or U20311 (N_20311,N_19577,N_19356);
nand U20312 (N_20312,N_19780,N_19128);
and U20313 (N_20313,N_19341,N_19836);
nand U20314 (N_20314,N_19954,N_19840);
nand U20315 (N_20315,N_19508,N_19114);
or U20316 (N_20316,N_19181,N_19396);
and U20317 (N_20317,N_19033,N_19865);
nor U20318 (N_20318,N_19699,N_19885);
and U20319 (N_20319,N_19245,N_19445);
nor U20320 (N_20320,N_19622,N_19794);
or U20321 (N_20321,N_19752,N_19366);
nand U20322 (N_20322,N_19604,N_19388);
and U20323 (N_20323,N_19797,N_19557);
or U20324 (N_20324,N_19607,N_19903);
nand U20325 (N_20325,N_19494,N_19882);
nor U20326 (N_20326,N_19088,N_19097);
nor U20327 (N_20327,N_19221,N_19005);
xnor U20328 (N_20328,N_19946,N_19205);
nor U20329 (N_20329,N_19746,N_19886);
and U20330 (N_20330,N_19937,N_19859);
nand U20331 (N_20331,N_19456,N_19086);
or U20332 (N_20332,N_19351,N_19888);
nor U20333 (N_20333,N_19939,N_19638);
and U20334 (N_20334,N_19262,N_19856);
or U20335 (N_20335,N_19755,N_19471);
and U20336 (N_20336,N_19073,N_19133);
or U20337 (N_20337,N_19879,N_19685);
nor U20338 (N_20338,N_19991,N_19938);
nand U20339 (N_20339,N_19649,N_19007);
nor U20340 (N_20340,N_19793,N_19414);
xnor U20341 (N_20341,N_19330,N_19539);
xnor U20342 (N_20342,N_19693,N_19314);
or U20343 (N_20343,N_19934,N_19842);
nand U20344 (N_20344,N_19300,N_19307);
or U20345 (N_20345,N_19541,N_19776);
nor U20346 (N_20346,N_19764,N_19734);
and U20347 (N_20347,N_19063,N_19567);
nor U20348 (N_20348,N_19052,N_19627);
xor U20349 (N_20349,N_19434,N_19064);
nor U20350 (N_20350,N_19117,N_19854);
or U20351 (N_20351,N_19119,N_19771);
nor U20352 (N_20352,N_19507,N_19056);
xor U20353 (N_20353,N_19325,N_19756);
or U20354 (N_20354,N_19208,N_19156);
nand U20355 (N_20355,N_19919,N_19345);
or U20356 (N_20356,N_19987,N_19818);
xor U20357 (N_20357,N_19218,N_19335);
nand U20358 (N_20358,N_19576,N_19069);
nand U20359 (N_20359,N_19994,N_19347);
or U20360 (N_20360,N_19093,N_19400);
nor U20361 (N_20361,N_19947,N_19322);
nand U20362 (N_20362,N_19010,N_19621);
nand U20363 (N_20363,N_19603,N_19967);
xnor U20364 (N_20364,N_19640,N_19629);
nor U20365 (N_20365,N_19561,N_19961);
nor U20366 (N_20366,N_19784,N_19013);
and U20367 (N_20367,N_19378,N_19417);
nor U20368 (N_20368,N_19258,N_19075);
nor U20369 (N_20369,N_19626,N_19067);
xnor U20370 (N_20370,N_19643,N_19477);
or U20371 (N_20371,N_19413,N_19724);
xor U20372 (N_20372,N_19813,N_19282);
nor U20373 (N_20373,N_19453,N_19584);
nor U20374 (N_20374,N_19913,N_19049);
xor U20375 (N_20375,N_19660,N_19729);
and U20376 (N_20376,N_19930,N_19923);
nand U20377 (N_20377,N_19505,N_19517);
nor U20378 (N_20378,N_19405,N_19416);
xnor U20379 (N_20379,N_19321,N_19380);
or U20380 (N_20380,N_19437,N_19333);
and U20381 (N_20381,N_19553,N_19600);
xnor U20382 (N_20382,N_19428,N_19511);
nand U20383 (N_20383,N_19503,N_19377);
and U20384 (N_20384,N_19514,N_19000);
or U20385 (N_20385,N_19247,N_19971);
and U20386 (N_20386,N_19763,N_19713);
nor U20387 (N_20387,N_19359,N_19327);
xor U20388 (N_20388,N_19868,N_19296);
nand U20389 (N_20389,N_19892,N_19972);
xnor U20390 (N_20390,N_19691,N_19696);
xor U20391 (N_20391,N_19272,N_19617);
nand U20392 (N_20392,N_19619,N_19195);
or U20393 (N_20393,N_19187,N_19782);
nand U20394 (N_20394,N_19490,N_19386);
nand U20395 (N_20395,N_19926,N_19648);
or U20396 (N_20396,N_19391,N_19901);
nand U20397 (N_20397,N_19080,N_19799);
xor U20398 (N_20398,N_19598,N_19761);
xor U20399 (N_20399,N_19066,N_19999);
nand U20400 (N_20400,N_19044,N_19055);
and U20401 (N_20401,N_19016,N_19815);
or U20402 (N_20402,N_19982,N_19802);
nor U20403 (N_20403,N_19252,N_19432);
nor U20404 (N_20404,N_19580,N_19165);
nand U20405 (N_20405,N_19132,N_19145);
and U20406 (N_20406,N_19178,N_19011);
or U20407 (N_20407,N_19122,N_19072);
xor U20408 (N_20408,N_19406,N_19227);
xor U20409 (N_20409,N_19725,N_19779);
nand U20410 (N_20410,N_19309,N_19222);
nand U20411 (N_20411,N_19966,N_19719);
or U20412 (N_20412,N_19689,N_19244);
nor U20413 (N_20413,N_19589,N_19042);
and U20414 (N_20414,N_19663,N_19775);
xor U20415 (N_20415,N_19100,N_19237);
or U20416 (N_20416,N_19807,N_19669);
or U20417 (N_20417,N_19185,N_19951);
nor U20418 (N_20418,N_19216,N_19339);
and U20419 (N_20419,N_19030,N_19130);
nor U20420 (N_20420,N_19610,N_19975);
and U20421 (N_20421,N_19915,N_19106);
xor U20422 (N_20422,N_19751,N_19976);
nor U20423 (N_20423,N_19292,N_19283);
xnor U20424 (N_20424,N_19138,N_19896);
xnor U20425 (N_20425,N_19121,N_19034);
xnor U20426 (N_20426,N_19591,N_19451);
or U20427 (N_20427,N_19140,N_19092);
and U20428 (N_20428,N_19712,N_19742);
nand U20429 (N_20429,N_19026,N_19931);
and U20430 (N_20430,N_19373,N_19078);
or U20431 (N_20431,N_19518,N_19313);
nor U20432 (N_20432,N_19028,N_19810);
or U20433 (N_20433,N_19904,N_19014);
or U20434 (N_20434,N_19164,N_19678);
and U20435 (N_20435,N_19383,N_19166);
or U20436 (N_20436,N_19427,N_19698);
nor U20437 (N_20437,N_19562,N_19611);
xor U20438 (N_20438,N_19146,N_19099);
nand U20439 (N_20439,N_19572,N_19402);
nor U20440 (N_20440,N_19747,N_19441);
nor U20441 (N_20441,N_19965,N_19964);
nand U20442 (N_20442,N_19139,N_19338);
nor U20443 (N_20443,N_19426,N_19677);
xnor U20444 (N_20444,N_19110,N_19382);
nand U20445 (N_20445,N_19554,N_19843);
or U20446 (N_20446,N_19968,N_19478);
nand U20447 (N_20447,N_19248,N_19774);
xor U20448 (N_20448,N_19143,N_19579);
nand U20449 (N_20449,N_19424,N_19666);
nand U20450 (N_20450,N_19646,N_19352);
nand U20451 (N_20451,N_19655,N_19126);
nor U20452 (N_20452,N_19350,N_19963);
nand U20453 (N_20453,N_19877,N_19618);
nor U20454 (N_20454,N_19259,N_19829);
and U20455 (N_20455,N_19692,N_19467);
and U20456 (N_20456,N_19394,N_19803);
and U20457 (N_20457,N_19962,N_19153);
nand U20458 (N_20458,N_19695,N_19986);
nand U20459 (N_20459,N_19022,N_19019);
nor U20460 (N_20460,N_19361,N_19104);
nor U20461 (N_20461,N_19612,N_19058);
or U20462 (N_20462,N_19728,N_19415);
nand U20463 (N_20463,N_19190,N_19912);
or U20464 (N_20464,N_19101,N_19552);
or U20465 (N_20465,N_19290,N_19977);
xnor U20466 (N_20466,N_19816,N_19635);
xnor U20467 (N_20467,N_19820,N_19657);
xor U20468 (N_20468,N_19342,N_19590);
nand U20469 (N_20469,N_19493,N_19464);
xnor U20470 (N_20470,N_19004,N_19095);
nor U20471 (N_20471,N_19422,N_19219);
or U20472 (N_20472,N_19922,N_19151);
or U20473 (N_20473,N_19036,N_19251);
or U20474 (N_20474,N_19163,N_19940);
nor U20475 (N_20475,N_19204,N_19125);
or U20476 (N_20476,N_19469,N_19862);
xnor U20477 (N_20477,N_19071,N_19997);
xnor U20478 (N_20478,N_19808,N_19715);
and U20479 (N_20479,N_19625,N_19461);
xnor U20480 (N_20480,N_19686,N_19176);
or U20481 (N_20481,N_19718,N_19302);
nor U20482 (N_20482,N_19592,N_19639);
nand U20483 (N_20483,N_19851,N_19542);
nand U20484 (N_20484,N_19834,N_19941);
or U20485 (N_20485,N_19801,N_19798);
or U20486 (N_20486,N_19847,N_19160);
and U20487 (N_20487,N_19050,N_19279);
nor U20488 (N_20488,N_19853,N_19444);
or U20489 (N_20489,N_19018,N_19795);
or U20490 (N_20490,N_19015,N_19317);
or U20491 (N_20491,N_19168,N_19172);
and U20492 (N_20492,N_19953,N_19537);
nand U20493 (N_20493,N_19236,N_19995);
or U20494 (N_20494,N_19062,N_19357);
xnor U20495 (N_20495,N_19688,N_19679);
nor U20496 (N_20496,N_19765,N_19609);
xnor U20497 (N_20497,N_19955,N_19990);
and U20498 (N_20498,N_19670,N_19608);
or U20499 (N_20499,N_19360,N_19275);
or U20500 (N_20500,N_19317,N_19122);
xnor U20501 (N_20501,N_19904,N_19882);
or U20502 (N_20502,N_19387,N_19875);
and U20503 (N_20503,N_19999,N_19501);
and U20504 (N_20504,N_19163,N_19890);
nand U20505 (N_20505,N_19685,N_19232);
xor U20506 (N_20506,N_19212,N_19114);
xor U20507 (N_20507,N_19586,N_19164);
xor U20508 (N_20508,N_19868,N_19850);
or U20509 (N_20509,N_19952,N_19839);
nor U20510 (N_20510,N_19969,N_19057);
or U20511 (N_20511,N_19634,N_19990);
nor U20512 (N_20512,N_19231,N_19200);
xnor U20513 (N_20513,N_19842,N_19893);
or U20514 (N_20514,N_19624,N_19116);
or U20515 (N_20515,N_19653,N_19300);
xor U20516 (N_20516,N_19330,N_19854);
xor U20517 (N_20517,N_19768,N_19580);
xor U20518 (N_20518,N_19101,N_19765);
and U20519 (N_20519,N_19295,N_19929);
nor U20520 (N_20520,N_19057,N_19951);
or U20521 (N_20521,N_19502,N_19250);
xor U20522 (N_20522,N_19379,N_19554);
nand U20523 (N_20523,N_19031,N_19376);
and U20524 (N_20524,N_19717,N_19075);
and U20525 (N_20525,N_19899,N_19053);
or U20526 (N_20526,N_19074,N_19988);
nand U20527 (N_20527,N_19341,N_19710);
and U20528 (N_20528,N_19840,N_19286);
xnor U20529 (N_20529,N_19431,N_19323);
nor U20530 (N_20530,N_19953,N_19732);
nor U20531 (N_20531,N_19519,N_19987);
and U20532 (N_20532,N_19428,N_19925);
and U20533 (N_20533,N_19543,N_19400);
nand U20534 (N_20534,N_19414,N_19288);
and U20535 (N_20535,N_19987,N_19061);
nor U20536 (N_20536,N_19586,N_19546);
or U20537 (N_20537,N_19687,N_19420);
xor U20538 (N_20538,N_19439,N_19389);
nand U20539 (N_20539,N_19798,N_19279);
or U20540 (N_20540,N_19542,N_19420);
and U20541 (N_20541,N_19859,N_19498);
nor U20542 (N_20542,N_19913,N_19353);
nand U20543 (N_20543,N_19741,N_19079);
xor U20544 (N_20544,N_19031,N_19311);
or U20545 (N_20545,N_19139,N_19495);
nand U20546 (N_20546,N_19228,N_19719);
and U20547 (N_20547,N_19768,N_19553);
nand U20548 (N_20548,N_19480,N_19071);
nor U20549 (N_20549,N_19236,N_19527);
xor U20550 (N_20550,N_19877,N_19944);
and U20551 (N_20551,N_19783,N_19454);
nor U20552 (N_20552,N_19383,N_19796);
nand U20553 (N_20553,N_19906,N_19261);
and U20554 (N_20554,N_19400,N_19297);
nand U20555 (N_20555,N_19303,N_19148);
and U20556 (N_20556,N_19282,N_19719);
or U20557 (N_20557,N_19970,N_19755);
nor U20558 (N_20558,N_19458,N_19920);
nand U20559 (N_20559,N_19204,N_19389);
nand U20560 (N_20560,N_19773,N_19187);
xnor U20561 (N_20561,N_19381,N_19920);
nand U20562 (N_20562,N_19934,N_19966);
nand U20563 (N_20563,N_19679,N_19693);
and U20564 (N_20564,N_19481,N_19024);
xnor U20565 (N_20565,N_19449,N_19345);
nand U20566 (N_20566,N_19324,N_19645);
or U20567 (N_20567,N_19461,N_19571);
and U20568 (N_20568,N_19900,N_19473);
nor U20569 (N_20569,N_19208,N_19984);
or U20570 (N_20570,N_19861,N_19322);
nand U20571 (N_20571,N_19532,N_19174);
nor U20572 (N_20572,N_19054,N_19013);
or U20573 (N_20573,N_19112,N_19117);
xnor U20574 (N_20574,N_19899,N_19145);
or U20575 (N_20575,N_19549,N_19174);
and U20576 (N_20576,N_19007,N_19028);
or U20577 (N_20577,N_19117,N_19846);
and U20578 (N_20578,N_19516,N_19366);
nor U20579 (N_20579,N_19762,N_19071);
xnor U20580 (N_20580,N_19481,N_19074);
nor U20581 (N_20581,N_19123,N_19663);
or U20582 (N_20582,N_19130,N_19872);
xor U20583 (N_20583,N_19694,N_19832);
nand U20584 (N_20584,N_19857,N_19192);
nor U20585 (N_20585,N_19887,N_19665);
nor U20586 (N_20586,N_19855,N_19033);
and U20587 (N_20587,N_19471,N_19576);
and U20588 (N_20588,N_19355,N_19263);
nor U20589 (N_20589,N_19655,N_19835);
xnor U20590 (N_20590,N_19988,N_19754);
nor U20591 (N_20591,N_19397,N_19420);
nand U20592 (N_20592,N_19323,N_19838);
nor U20593 (N_20593,N_19336,N_19743);
and U20594 (N_20594,N_19759,N_19881);
or U20595 (N_20595,N_19385,N_19562);
and U20596 (N_20596,N_19935,N_19832);
xor U20597 (N_20597,N_19556,N_19205);
nor U20598 (N_20598,N_19209,N_19381);
xnor U20599 (N_20599,N_19235,N_19751);
and U20600 (N_20600,N_19116,N_19604);
nor U20601 (N_20601,N_19861,N_19541);
and U20602 (N_20602,N_19399,N_19034);
nor U20603 (N_20603,N_19631,N_19736);
xnor U20604 (N_20604,N_19869,N_19682);
nand U20605 (N_20605,N_19908,N_19830);
or U20606 (N_20606,N_19358,N_19053);
and U20607 (N_20607,N_19737,N_19202);
xnor U20608 (N_20608,N_19241,N_19267);
or U20609 (N_20609,N_19619,N_19689);
nand U20610 (N_20610,N_19933,N_19103);
nor U20611 (N_20611,N_19633,N_19046);
nand U20612 (N_20612,N_19985,N_19229);
nor U20613 (N_20613,N_19228,N_19793);
nand U20614 (N_20614,N_19649,N_19781);
xnor U20615 (N_20615,N_19742,N_19454);
xnor U20616 (N_20616,N_19016,N_19976);
and U20617 (N_20617,N_19620,N_19092);
xor U20618 (N_20618,N_19147,N_19294);
nor U20619 (N_20619,N_19151,N_19133);
xnor U20620 (N_20620,N_19621,N_19952);
xnor U20621 (N_20621,N_19317,N_19147);
nor U20622 (N_20622,N_19927,N_19584);
and U20623 (N_20623,N_19413,N_19609);
or U20624 (N_20624,N_19451,N_19624);
or U20625 (N_20625,N_19254,N_19952);
or U20626 (N_20626,N_19503,N_19204);
xnor U20627 (N_20627,N_19300,N_19607);
and U20628 (N_20628,N_19542,N_19262);
and U20629 (N_20629,N_19699,N_19230);
and U20630 (N_20630,N_19396,N_19114);
xor U20631 (N_20631,N_19905,N_19158);
and U20632 (N_20632,N_19621,N_19279);
and U20633 (N_20633,N_19037,N_19423);
or U20634 (N_20634,N_19482,N_19831);
nand U20635 (N_20635,N_19603,N_19099);
xnor U20636 (N_20636,N_19250,N_19303);
or U20637 (N_20637,N_19213,N_19308);
xnor U20638 (N_20638,N_19455,N_19586);
or U20639 (N_20639,N_19597,N_19971);
or U20640 (N_20640,N_19223,N_19489);
nor U20641 (N_20641,N_19536,N_19847);
or U20642 (N_20642,N_19359,N_19860);
or U20643 (N_20643,N_19677,N_19279);
and U20644 (N_20644,N_19772,N_19280);
or U20645 (N_20645,N_19947,N_19422);
or U20646 (N_20646,N_19596,N_19718);
nor U20647 (N_20647,N_19539,N_19244);
or U20648 (N_20648,N_19960,N_19009);
xor U20649 (N_20649,N_19748,N_19592);
or U20650 (N_20650,N_19940,N_19461);
nand U20651 (N_20651,N_19917,N_19446);
xor U20652 (N_20652,N_19688,N_19998);
nand U20653 (N_20653,N_19619,N_19155);
xnor U20654 (N_20654,N_19508,N_19373);
nand U20655 (N_20655,N_19159,N_19605);
and U20656 (N_20656,N_19642,N_19778);
nand U20657 (N_20657,N_19874,N_19847);
nor U20658 (N_20658,N_19763,N_19719);
nand U20659 (N_20659,N_19945,N_19405);
and U20660 (N_20660,N_19253,N_19400);
xnor U20661 (N_20661,N_19679,N_19887);
nor U20662 (N_20662,N_19693,N_19495);
nand U20663 (N_20663,N_19014,N_19433);
xor U20664 (N_20664,N_19820,N_19112);
and U20665 (N_20665,N_19003,N_19642);
and U20666 (N_20666,N_19225,N_19424);
nand U20667 (N_20667,N_19604,N_19510);
nand U20668 (N_20668,N_19553,N_19685);
or U20669 (N_20669,N_19733,N_19651);
or U20670 (N_20670,N_19936,N_19382);
nand U20671 (N_20671,N_19301,N_19651);
xor U20672 (N_20672,N_19789,N_19538);
and U20673 (N_20673,N_19370,N_19112);
or U20674 (N_20674,N_19456,N_19024);
xnor U20675 (N_20675,N_19799,N_19905);
and U20676 (N_20676,N_19014,N_19829);
or U20677 (N_20677,N_19633,N_19655);
nor U20678 (N_20678,N_19394,N_19124);
xor U20679 (N_20679,N_19616,N_19486);
and U20680 (N_20680,N_19807,N_19601);
nand U20681 (N_20681,N_19037,N_19496);
and U20682 (N_20682,N_19275,N_19666);
nor U20683 (N_20683,N_19416,N_19031);
xor U20684 (N_20684,N_19511,N_19673);
nor U20685 (N_20685,N_19147,N_19116);
nor U20686 (N_20686,N_19035,N_19061);
xor U20687 (N_20687,N_19804,N_19058);
nor U20688 (N_20688,N_19935,N_19406);
and U20689 (N_20689,N_19880,N_19404);
nand U20690 (N_20690,N_19358,N_19817);
nor U20691 (N_20691,N_19024,N_19947);
or U20692 (N_20692,N_19223,N_19283);
or U20693 (N_20693,N_19656,N_19621);
nand U20694 (N_20694,N_19033,N_19631);
and U20695 (N_20695,N_19986,N_19353);
nor U20696 (N_20696,N_19577,N_19804);
and U20697 (N_20697,N_19163,N_19267);
nand U20698 (N_20698,N_19466,N_19205);
and U20699 (N_20699,N_19137,N_19979);
and U20700 (N_20700,N_19642,N_19379);
nor U20701 (N_20701,N_19314,N_19755);
and U20702 (N_20702,N_19559,N_19587);
nor U20703 (N_20703,N_19264,N_19575);
nand U20704 (N_20704,N_19937,N_19267);
or U20705 (N_20705,N_19539,N_19567);
xor U20706 (N_20706,N_19377,N_19713);
nor U20707 (N_20707,N_19411,N_19374);
or U20708 (N_20708,N_19857,N_19798);
or U20709 (N_20709,N_19830,N_19639);
nor U20710 (N_20710,N_19961,N_19426);
xor U20711 (N_20711,N_19103,N_19919);
nor U20712 (N_20712,N_19859,N_19395);
nand U20713 (N_20713,N_19604,N_19324);
nand U20714 (N_20714,N_19084,N_19320);
and U20715 (N_20715,N_19559,N_19809);
and U20716 (N_20716,N_19664,N_19436);
or U20717 (N_20717,N_19844,N_19892);
xor U20718 (N_20718,N_19425,N_19255);
nor U20719 (N_20719,N_19643,N_19571);
xor U20720 (N_20720,N_19542,N_19334);
xnor U20721 (N_20721,N_19194,N_19922);
nor U20722 (N_20722,N_19467,N_19619);
and U20723 (N_20723,N_19684,N_19627);
xnor U20724 (N_20724,N_19511,N_19540);
nand U20725 (N_20725,N_19018,N_19568);
or U20726 (N_20726,N_19242,N_19958);
xor U20727 (N_20727,N_19848,N_19636);
nor U20728 (N_20728,N_19746,N_19961);
nand U20729 (N_20729,N_19844,N_19275);
nor U20730 (N_20730,N_19136,N_19438);
nand U20731 (N_20731,N_19832,N_19519);
or U20732 (N_20732,N_19416,N_19486);
xor U20733 (N_20733,N_19305,N_19661);
and U20734 (N_20734,N_19743,N_19700);
and U20735 (N_20735,N_19345,N_19532);
nor U20736 (N_20736,N_19023,N_19141);
nor U20737 (N_20737,N_19857,N_19080);
nor U20738 (N_20738,N_19532,N_19642);
nor U20739 (N_20739,N_19161,N_19580);
or U20740 (N_20740,N_19556,N_19007);
nand U20741 (N_20741,N_19768,N_19997);
or U20742 (N_20742,N_19374,N_19196);
or U20743 (N_20743,N_19296,N_19375);
nor U20744 (N_20744,N_19668,N_19060);
or U20745 (N_20745,N_19731,N_19017);
nand U20746 (N_20746,N_19588,N_19671);
or U20747 (N_20747,N_19480,N_19821);
and U20748 (N_20748,N_19047,N_19962);
nand U20749 (N_20749,N_19117,N_19328);
nor U20750 (N_20750,N_19585,N_19065);
nand U20751 (N_20751,N_19058,N_19438);
nand U20752 (N_20752,N_19519,N_19910);
nand U20753 (N_20753,N_19469,N_19606);
xnor U20754 (N_20754,N_19951,N_19555);
nand U20755 (N_20755,N_19404,N_19388);
or U20756 (N_20756,N_19783,N_19476);
nor U20757 (N_20757,N_19809,N_19679);
nand U20758 (N_20758,N_19362,N_19295);
nor U20759 (N_20759,N_19890,N_19495);
nand U20760 (N_20760,N_19128,N_19567);
xnor U20761 (N_20761,N_19595,N_19618);
or U20762 (N_20762,N_19328,N_19928);
and U20763 (N_20763,N_19289,N_19586);
or U20764 (N_20764,N_19551,N_19975);
xnor U20765 (N_20765,N_19807,N_19805);
nor U20766 (N_20766,N_19639,N_19145);
or U20767 (N_20767,N_19594,N_19823);
and U20768 (N_20768,N_19334,N_19607);
xnor U20769 (N_20769,N_19860,N_19192);
nand U20770 (N_20770,N_19782,N_19518);
and U20771 (N_20771,N_19186,N_19751);
and U20772 (N_20772,N_19547,N_19806);
and U20773 (N_20773,N_19426,N_19531);
xnor U20774 (N_20774,N_19309,N_19467);
xnor U20775 (N_20775,N_19768,N_19089);
nand U20776 (N_20776,N_19719,N_19967);
or U20777 (N_20777,N_19319,N_19625);
nor U20778 (N_20778,N_19201,N_19314);
nand U20779 (N_20779,N_19941,N_19056);
xnor U20780 (N_20780,N_19418,N_19142);
nor U20781 (N_20781,N_19329,N_19413);
nand U20782 (N_20782,N_19458,N_19251);
nand U20783 (N_20783,N_19894,N_19188);
or U20784 (N_20784,N_19227,N_19305);
xnor U20785 (N_20785,N_19478,N_19860);
xnor U20786 (N_20786,N_19734,N_19924);
or U20787 (N_20787,N_19736,N_19830);
or U20788 (N_20788,N_19605,N_19557);
or U20789 (N_20789,N_19408,N_19299);
xnor U20790 (N_20790,N_19542,N_19438);
xnor U20791 (N_20791,N_19833,N_19076);
nor U20792 (N_20792,N_19624,N_19314);
nand U20793 (N_20793,N_19566,N_19948);
nor U20794 (N_20794,N_19363,N_19171);
xor U20795 (N_20795,N_19022,N_19962);
nand U20796 (N_20796,N_19515,N_19308);
nand U20797 (N_20797,N_19862,N_19963);
nand U20798 (N_20798,N_19234,N_19885);
nor U20799 (N_20799,N_19413,N_19575);
nand U20800 (N_20800,N_19531,N_19216);
xor U20801 (N_20801,N_19383,N_19126);
and U20802 (N_20802,N_19214,N_19856);
and U20803 (N_20803,N_19395,N_19393);
nand U20804 (N_20804,N_19849,N_19323);
or U20805 (N_20805,N_19232,N_19725);
or U20806 (N_20806,N_19771,N_19806);
or U20807 (N_20807,N_19508,N_19119);
xor U20808 (N_20808,N_19654,N_19165);
or U20809 (N_20809,N_19167,N_19651);
nor U20810 (N_20810,N_19683,N_19377);
nand U20811 (N_20811,N_19674,N_19456);
or U20812 (N_20812,N_19969,N_19416);
nand U20813 (N_20813,N_19454,N_19112);
nor U20814 (N_20814,N_19516,N_19758);
or U20815 (N_20815,N_19427,N_19184);
xnor U20816 (N_20816,N_19720,N_19535);
or U20817 (N_20817,N_19661,N_19849);
nor U20818 (N_20818,N_19129,N_19448);
nor U20819 (N_20819,N_19817,N_19286);
nor U20820 (N_20820,N_19434,N_19110);
nand U20821 (N_20821,N_19226,N_19302);
nor U20822 (N_20822,N_19612,N_19450);
and U20823 (N_20823,N_19654,N_19066);
or U20824 (N_20824,N_19038,N_19801);
xor U20825 (N_20825,N_19351,N_19781);
nand U20826 (N_20826,N_19764,N_19831);
and U20827 (N_20827,N_19161,N_19251);
and U20828 (N_20828,N_19795,N_19533);
nand U20829 (N_20829,N_19022,N_19561);
and U20830 (N_20830,N_19555,N_19199);
or U20831 (N_20831,N_19318,N_19978);
nor U20832 (N_20832,N_19698,N_19852);
xnor U20833 (N_20833,N_19921,N_19150);
and U20834 (N_20834,N_19632,N_19686);
nand U20835 (N_20835,N_19529,N_19309);
xor U20836 (N_20836,N_19719,N_19316);
nand U20837 (N_20837,N_19547,N_19962);
xor U20838 (N_20838,N_19624,N_19246);
nor U20839 (N_20839,N_19517,N_19334);
and U20840 (N_20840,N_19484,N_19676);
or U20841 (N_20841,N_19742,N_19013);
or U20842 (N_20842,N_19036,N_19716);
and U20843 (N_20843,N_19381,N_19236);
nand U20844 (N_20844,N_19337,N_19322);
or U20845 (N_20845,N_19008,N_19738);
nand U20846 (N_20846,N_19916,N_19268);
or U20847 (N_20847,N_19687,N_19446);
and U20848 (N_20848,N_19620,N_19879);
xnor U20849 (N_20849,N_19977,N_19537);
and U20850 (N_20850,N_19683,N_19631);
xor U20851 (N_20851,N_19191,N_19716);
nor U20852 (N_20852,N_19742,N_19178);
and U20853 (N_20853,N_19900,N_19625);
nand U20854 (N_20854,N_19657,N_19707);
and U20855 (N_20855,N_19244,N_19235);
nand U20856 (N_20856,N_19369,N_19607);
nand U20857 (N_20857,N_19920,N_19425);
and U20858 (N_20858,N_19780,N_19327);
or U20859 (N_20859,N_19158,N_19417);
xor U20860 (N_20860,N_19224,N_19210);
nand U20861 (N_20861,N_19660,N_19344);
xor U20862 (N_20862,N_19952,N_19043);
xor U20863 (N_20863,N_19521,N_19327);
nor U20864 (N_20864,N_19034,N_19518);
nand U20865 (N_20865,N_19941,N_19805);
xor U20866 (N_20866,N_19252,N_19208);
xor U20867 (N_20867,N_19614,N_19514);
nor U20868 (N_20868,N_19135,N_19052);
and U20869 (N_20869,N_19466,N_19409);
or U20870 (N_20870,N_19061,N_19106);
nand U20871 (N_20871,N_19840,N_19340);
or U20872 (N_20872,N_19135,N_19378);
nand U20873 (N_20873,N_19406,N_19099);
nor U20874 (N_20874,N_19465,N_19004);
and U20875 (N_20875,N_19841,N_19238);
or U20876 (N_20876,N_19565,N_19053);
nor U20877 (N_20877,N_19325,N_19925);
xnor U20878 (N_20878,N_19677,N_19112);
xnor U20879 (N_20879,N_19361,N_19241);
and U20880 (N_20880,N_19686,N_19436);
nor U20881 (N_20881,N_19970,N_19523);
nor U20882 (N_20882,N_19388,N_19187);
nand U20883 (N_20883,N_19459,N_19624);
and U20884 (N_20884,N_19383,N_19043);
nand U20885 (N_20885,N_19986,N_19283);
and U20886 (N_20886,N_19132,N_19071);
nand U20887 (N_20887,N_19878,N_19562);
nor U20888 (N_20888,N_19687,N_19594);
or U20889 (N_20889,N_19021,N_19619);
nor U20890 (N_20890,N_19695,N_19255);
and U20891 (N_20891,N_19729,N_19981);
nor U20892 (N_20892,N_19698,N_19610);
and U20893 (N_20893,N_19357,N_19340);
nand U20894 (N_20894,N_19202,N_19330);
or U20895 (N_20895,N_19336,N_19354);
nand U20896 (N_20896,N_19481,N_19853);
nor U20897 (N_20897,N_19549,N_19319);
or U20898 (N_20898,N_19997,N_19740);
xnor U20899 (N_20899,N_19465,N_19352);
nand U20900 (N_20900,N_19897,N_19155);
nor U20901 (N_20901,N_19323,N_19360);
nand U20902 (N_20902,N_19253,N_19603);
xor U20903 (N_20903,N_19148,N_19622);
nor U20904 (N_20904,N_19651,N_19603);
or U20905 (N_20905,N_19210,N_19070);
and U20906 (N_20906,N_19533,N_19315);
and U20907 (N_20907,N_19015,N_19739);
or U20908 (N_20908,N_19163,N_19457);
and U20909 (N_20909,N_19438,N_19382);
nand U20910 (N_20910,N_19969,N_19494);
or U20911 (N_20911,N_19135,N_19054);
and U20912 (N_20912,N_19506,N_19201);
or U20913 (N_20913,N_19043,N_19388);
and U20914 (N_20914,N_19045,N_19984);
and U20915 (N_20915,N_19448,N_19733);
nand U20916 (N_20916,N_19546,N_19467);
nor U20917 (N_20917,N_19438,N_19402);
xnor U20918 (N_20918,N_19046,N_19129);
xor U20919 (N_20919,N_19030,N_19964);
xnor U20920 (N_20920,N_19521,N_19929);
and U20921 (N_20921,N_19748,N_19528);
and U20922 (N_20922,N_19237,N_19136);
or U20923 (N_20923,N_19165,N_19884);
and U20924 (N_20924,N_19468,N_19666);
nor U20925 (N_20925,N_19112,N_19256);
or U20926 (N_20926,N_19704,N_19779);
or U20927 (N_20927,N_19615,N_19239);
nand U20928 (N_20928,N_19905,N_19703);
nand U20929 (N_20929,N_19031,N_19717);
and U20930 (N_20930,N_19352,N_19738);
or U20931 (N_20931,N_19614,N_19523);
nor U20932 (N_20932,N_19551,N_19740);
nand U20933 (N_20933,N_19515,N_19259);
nor U20934 (N_20934,N_19592,N_19705);
nor U20935 (N_20935,N_19716,N_19846);
xor U20936 (N_20936,N_19202,N_19716);
and U20937 (N_20937,N_19518,N_19996);
xnor U20938 (N_20938,N_19119,N_19260);
nor U20939 (N_20939,N_19102,N_19663);
or U20940 (N_20940,N_19636,N_19282);
nor U20941 (N_20941,N_19204,N_19328);
or U20942 (N_20942,N_19884,N_19106);
or U20943 (N_20943,N_19344,N_19377);
xor U20944 (N_20944,N_19398,N_19228);
or U20945 (N_20945,N_19337,N_19265);
or U20946 (N_20946,N_19127,N_19949);
and U20947 (N_20947,N_19153,N_19616);
or U20948 (N_20948,N_19830,N_19722);
xor U20949 (N_20949,N_19668,N_19382);
and U20950 (N_20950,N_19608,N_19594);
and U20951 (N_20951,N_19393,N_19878);
nor U20952 (N_20952,N_19868,N_19743);
xor U20953 (N_20953,N_19902,N_19536);
nand U20954 (N_20954,N_19195,N_19779);
and U20955 (N_20955,N_19326,N_19056);
or U20956 (N_20956,N_19552,N_19511);
or U20957 (N_20957,N_19620,N_19860);
nand U20958 (N_20958,N_19355,N_19775);
xor U20959 (N_20959,N_19440,N_19329);
nor U20960 (N_20960,N_19297,N_19564);
xnor U20961 (N_20961,N_19885,N_19900);
or U20962 (N_20962,N_19417,N_19582);
xnor U20963 (N_20963,N_19426,N_19756);
xnor U20964 (N_20964,N_19192,N_19028);
nand U20965 (N_20965,N_19267,N_19191);
nand U20966 (N_20966,N_19644,N_19436);
or U20967 (N_20967,N_19027,N_19837);
and U20968 (N_20968,N_19814,N_19598);
nor U20969 (N_20969,N_19948,N_19982);
or U20970 (N_20970,N_19372,N_19746);
or U20971 (N_20971,N_19996,N_19386);
or U20972 (N_20972,N_19706,N_19211);
nor U20973 (N_20973,N_19600,N_19820);
xor U20974 (N_20974,N_19542,N_19209);
and U20975 (N_20975,N_19696,N_19179);
or U20976 (N_20976,N_19363,N_19748);
nor U20977 (N_20977,N_19655,N_19153);
nand U20978 (N_20978,N_19507,N_19122);
nand U20979 (N_20979,N_19096,N_19936);
and U20980 (N_20980,N_19481,N_19301);
nand U20981 (N_20981,N_19073,N_19176);
and U20982 (N_20982,N_19021,N_19078);
nand U20983 (N_20983,N_19687,N_19603);
xor U20984 (N_20984,N_19951,N_19223);
or U20985 (N_20985,N_19242,N_19300);
or U20986 (N_20986,N_19615,N_19934);
or U20987 (N_20987,N_19848,N_19874);
nand U20988 (N_20988,N_19649,N_19101);
nor U20989 (N_20989,N_19672,N_19160);
nand U20990 (N_20990,N_19732,N_19943);
nand U20991 (N_20991,N_19914,N_19231);
nand U20992 (N_20992,N_19123,N_19070);
nand U20993 (N_20993,N_19410,N_19034);
nand U20994 (N_20994,N_19026,N_19991);
xnor U20995 (N_20995,N_19982,N_19111);
nand U20996 (N_20996,N_19009,N_19400);
and U20997 (N_20997,N_19313,N_19935);
or U20998 (N_20998,N_19202,N_19169);
nand U20999 (N_20999,N_19248,N_19392);
xor U21000 (N_21000,N_20977,N_20023);
or U21001 (N_21001,N_20301,N_20249);
nand U21002 (N_21002,N_20118,N_20745);
xnor U21003 (N_21003,N_20610,N_20324);
nand U21004 (N_21004,N_20241,N_20509);
nor U21005 (N_21005,N_20450,N_20021);
nand U21006 (N_21006,N_20197,N_20674);
xor U21007 (N_21007,N_20128,N_20865);
or U21008 (N_21008,N_20753,N_20972);
xnor U21009 (N_21009,N_20133,N_20199);
and U21010 (N_21010,N_20067,N_20104);
nand U21011 (N_21011,N_20729,N_20086);
nand U21012 (N_21012,N_20093,N_20192);
or U21013 (N_21013,N_20231,N_20982);
nand U21014 (N_21014,N_20766,N_20054);
nand U21015 (N_21015,N_20285,N_20860);
nand U21016 (N_21016,N_20418,N_20845);
nor U21017 (N_21017,N_20015,N_20205);
nand U21018 (N_21018,N_20648,N_20840);
or U21019 (N_21019,N_20469,N_20783);
nand U21020 (N_21020,N_20772,N_20874);
nand U21021 (N_21021,N_20835,N_20373);
nand U21022 (N_21022,N_20536,N_20432);
or U21023 (N_21023,N_20375,N_20158);
or U21024 (N_21024,N_20593,N_20777);
and U21025 (N_21025,N_20555,N_20893);
or U21026 (N_21026,N_20239,N_20687);
xnor U21027 (N_21027,N_20020,N_20750);
and U21028 (N_21028,N_20743,N_20725);
nand U21029 (N_21029,N_20526,N_20665);
and U21030 (N_21030,N_20580,N_20075);
or U21031 (N_21031,N_20853,N_20083);
or U21032 (N_21032,N_20574,N_20191);
and U21033 (N_21033,N_20833,N_20468);
nand U21034 (N_21034,N_20990,N_20952);
nand U21035 (N_21035,N_20973,N_20639);
or U21036 (N_21036,N_20919,N_20867);
nand U21037 (N_21037,N_20483,N_20635);
and U21038 (N_21038,N_20559,N_20905);
or U21039 (N_21039,N_20993,N_20364);
or U21040 (N_21040,N_20332,N_20415);
xor U21041 (N_21041,N_20934,N_20516);
or U21042 (N_21042,N_20140,N_20568);
xor U21043 (N_21043,N_20855,N_20683);
or U21044 (N_21044,N_20802,N_20524);
or U21045 (N_21045,N_20870,N_20727);
nor U21046 (N_21046,N_20137,N_20314);
xnor U21047 (N_21047,N_20566,N_20911);
or U21048 (N_21048,N_20269,N_20286);
xor U21049 (N_21049,N_20031,N_20082);
nor U21050 (N_21050,N_20071,N_20436);
or U21051 (N_21051,N_20931,N_20254);
xor U21052 (N_21052,N_20986,N_20357);
or U21053 (N_21053,N_20120,N_20393);
xor U21054 (N_21054,N_20955,N_20603);
and U21055 (N_21055,N_20848,N_20511);
xor U21056 (N_21056,N_20821,N_20504);
nand U21057 (N_21057,N_20278,N_20922);
or U21058 (N_21058,N_20562,N_20527);
and U21059 (N_21059,N_20116,N_20452);
and U21060 (N_21060,N_20765,N_20784);
or U21061 (N_21061,N_20569,N_20200);
xnor U21062 (N_21062,N_20421,N_20994);
or U21063 (N_21063,N_20878,N_20155);
xnor U21064 (N_21064,N_20045,N_20275);
or U21065 (N_21065,N_20781,N_20462);
or U21066 (N_21066,N_20726,N_20447);
nand U21067 (N_21067,N_20429,N_20607);
nor U21068 (N_21068,N_20970,N_20394);
nor U21069 (N_21069,N_20696,N_20228);
or U21070 (N_21070,N_20299,N_20715);
and U21071 (N_21071,N_20804,N_20805);
xnor U21072 (N_21072,N_20287,N_20974);
xor U21073 (N_21073,N_20573,N_20721);
or U21074 (N_21074,N_20068,N_20327);
xnor U21075 (N_21075,N_20737,N_20789);
xor U21076 (N_21076,N_20401,N_20303);
nor U21077 (N_21077,N_20502,N_20288);
and U21078 (N_21078,N_20242,N_20954);
nand U21079 (N_21079,N_20708,N_20035);
xor U21080 (N_21080,N_20260,N_20608);
xnor U21081 (N_21081,N_20733,N_20591);
nor U21082 (N_21082,N_20551,N_20300);
xnor U21083 (N_21083,N_20222,N_20305);
nor U21084 (N_21084,N_20512,N_20077);
and U21085 (N_21085,N_20882,N_20255);
nand U21086 (N_21086,N_20538,N_20666);
nor U21087 (N_21087,N_20486,N_20995);
nor U21088 (N_21088,N_20892,N_20353);
or U21089 (N_21089,N_20969,N_20206);
nand U21090 (N_21090,N_20383,N_20984);
xor U21091 (N_21091,N_20700,N_20331);
nand U21092 (N_21092,N_20194,N_20474);
nor U21093 (N_21093,N_20355,N_20791);
or U21094 (N_21094,N_20265,N_20003);
nand U21095 (N_21095,N_20460,N_20564);
xor U21096 (N_21096,N_20038,N_20283);
and U21097 (N_21097,N_20245,N_20862);
and U21098 (N_21098,N_20746,N_20382);
and U21099 (N_21099,N_20144,N_20647);
and U21100 (N_21100,N_20032,N_20742);
nand U21101 (N_21101,N_20686,N_20177);
xor U21102 (N_21102,N_20461,N_20230);
nand U21103 (N_21103,N_20004,N_20018);
nor U21104 (N_21104,N_20800,N_20274);
nor U21105 (N_21105,N_20810,N_20291);
or U21106 (N_21106,N_20413,N_20496);
and U21107 (N_21107,N_20698,N_20653);
and U21108 (N_21108,N_20361,N_20497);
xor U21109 (N_21109,N_20170,N_20136);
nor U21110 (N_21110,N_20614,N_20220);
nand U21111 (N_21111,N_20159,N_20214);
nor U21112 (N_21112,N_20836,N_20762);
or U21113 (N_21113,N_20384,N_20325);
or U21114 (N_21114,N_20088,N_20704);
or U21115 (N_21115,N_20780,N_20962);
xnor U21116 (N_21116,N_20050,N_20362);
xor U21117 (N_21117,N_20433,N_20290);
or U21118 (N_21118,N_20978,N_20112);
nand U21119 (N_21119,N_20216,N_20585);
nor U21120 (N_21120,N_20404,N_20545);
xnor U21121 (N_21121,N_20042,N_20084);
xnor U21122 (N_21122,N_20289,N_20351);
and U21123 (N_21123,N_20567,N_20051);
xor U21124 (N_21124,N_20929,N_20473);
nor U21125 (N_21125,N_20861,N_20349);
xnor U21126 (N_21126,N_20012,N_20902);
and U21127 (N_21127,N_20329,N_20221);
nor U21128 (N_21128,N_20487,N_20797);
or U21129 (N_21129,N_20025,N_20940);
xor U21130 (N_21130,N_20823,N_20831);
xnor U21131 (N_21131,N_20198,N_20918);
nand U21132 (N_21132,N_20690,N_20506);
and U21133 (N_21133,N_20407,N_20234);
xor U21134 (N_21134,N_20352,N_20033);
and U21135 (N_21135,N_20061,N_20759);
nor U21136 (N_21136,N_20310,N_20098);
nor U21137 (N_21137,N_20963,N_20103);
and U21138 (N_21138,N_20028,N_20097);
nor U21139 (N_21139,N_20901,N_20139);
nor U21140 (N_21140,N_20296,N_20992);
nand U21141 (N_21141,N_20711,N_20204);
or U21142 (N_21142,N_20839,N_20634);
xor U21143 (N_21143,N_20034,N_20798);
nand U21144 (N_21144,N_20667,N_20793);
or U21145 (N_21145,N_20572,N_20047);
nand U21146 (N_21146,N_20040,N_20253);
nor U21147 (N_21147,N_20838,N_20672);
nand U21148 (N_21148,N_20420,N_20514);
or U21149 (N_21149,N_20760,N_20812);
or U21150 (N_21150,N_20212,N_20517);
nand U21151 (N_21151,N_20428,N_20942);
nand U21152 (N_21152,N_20157,N_20163);
and U21153 (N_21153,N_20115,N_20423);
nand U21154 (N_21154,N_20425,N_20550);
xnor U21155 (N_21155,N_20341,N_20751);
and U21156 (N_21156,N_20145,N_20196);
nor U21157 (N_21157,N_20825,N_20964);
nand U21158 (N_21158,N_20074,N_20907);
nand U21159 (N_21159,N_20149,N_20662);
nor U21160 (N_21160,N_20691,N_20722);
nand U21161 (N_21161,N_20164,N_20135);
and U21162 (N_21162,N_20642,N_20264);
or U21163 (N_21163,N_20092,N_20431);
and U21164 (N_21164,N_20859,N_20561);
or U21165 (N_21165,N_20215,N_20632);
xnor U21166 (N_21166,N_20426,N_20008);
nand U21167 (N_21167,N_20530,N_20081);
nand U21168 (N_21168,N_20367,N_20251);
xor U21169 (N_21169,N_20983,N_20724);
nand U21170 (N_21170,N_20770,N_20270);
nor U21171 (N_21171,N_20630,N_20225);
and U21172 (N_21172,N_20832,N_20454);
xnor U21173 (N_21173,N_20085,N_20043);
nand U21174 (N_21174,N_20078,N_20069);
nor U21175 (N_21175,N_20592,N_20606);
and U21176 (N_21176,N_20763,N_20186);
and U21177 (N_21177,N_20363,N_20224);
nand U21178 (N_21178,N_20250,N_20443);
and U21179 (N_21179,N_20890,N_20340);
and U21180 (N_21180,N_20856,N_20651);
nor U21181 (N_21181,N_20076,N_20702);
nand U21182 (N_21182,N_20879,N_20001);
and U21183 (N_21183,N_20619,N_20485);
nor U21184 (N_21184,N_20943,N_20307);
xor U21185 (N_21185,N_20609,N_20761);
and U21186 (N_21186,N_20888,N_20132);
and U21187 (N_21187,N_20440,N_20152);
and U21188 (N_21188,N_20312,N_20178);
xor U21189 (N_21189,N_20261,N_20827);
xor U21190 (N_21190,N_20828,N_20446);
or U21191 (N_21191,N_20933,N_20876);
or U21192 (N_21192,N_20681,N_20563);
nor U21193 (N_21193,N_20937,N_20409);
or U21194 (N_21194,N_20884,N_20162);
or U21195 (N_21195,N_20895,N_20676);
nor U21196 (N_21196,N_20900,N_20801);
nor U21197 (N_21197,N_20985,N_20655);
nor U21198 (N_21198,N_20424,N_20165);
and U21199 (N_21199,N_20237,N_20660);
nor U21200 (N_21200,N_20803,N_20932);
nor U21201 (N_21201,N_20011,N_20786);
xnor U21202 (N_21202,N_20673,N_20022);
and U21203 (N_21203,N_20476,N_20101);
or U21204 (N_21204,N_20013,N_20598);
or U21205 (N_21205,N_20965,N_20953);
or U21206 (N_21206,N_20557,N_20734);
and U21207 (N_21207,N_20534,N_20176);
xnor U21208 (N_21208,N_20909,N_20481);
nand U21209 (N_21209,N_20489,N_20259);
xnor U21210 (N_21210,N_20295,N_20604);
nor U21211 (N_21211,N_20981,N_20492);
nand U21212 (N_21212,N_20350,N_20546);
and U21213 (N_21213,N_20376,N_20749);
nand U21214 (N_21214,N_20731,N_20099);
and U21215 (N_21215,N_20449,N_20682);
or U21216 (N_21216,N_20988,N_20208);
and U21217 (N_21217,N_20202,N_20358);
nand U21218 (N_21218,N_20684,N_20185);
xnor U21219 (N_21219,N_20999,N_20380);
or U21220 (N_21220,N_20153,N_20671);
and U21221 (N_21221,N_20243,N_20044);
or U21222 (N_21222,N_20834,N_20638);
xor U21223 (N_21223,N_20218,N_20629);
or U21224 (N_21224,N_20055,N_20588);
xnor U21225 (N_21225,N_20595,N_20997);
nand U21226 (N_21226,N_20656,N_20000);
nor U21227 (N_21227,N_20612,N_20755);
or U21228 (N_21228,N_20586,N_20589);
or U21229 (N_21229,N_20464,N_20266);
and U21230 (N_21230,N_20842,N_20774);
or U21231 (N_21231,N_20806,N_20778);
or U21232 (N_21232,N_20887,N_20430);
and U21233 (N_21233,N_20542,N_20372);
and U21234 (N_21234,N_20499,N_20847);
or U21235 (N_21235,N_20663,N_20070);
nor U21236 (N_21236,N_20475,N_20959);
nand U21237 (N_21237,N_20529,N_20851);
xor U21238 (N_21238,N_20718,N_20544);
and U21239 (N_21239,N_20906,N_20613);
xor U21240 (N_21240,N_20408,N_20921);
and U21241 (N_21241,N_20392,N_20650);
nand U21242 (N_21242,N_20026,N_20720);
nor U21243 (N_21243,N_20773,N_20455);
or U21244 (N_21244,N_20438,N_20041);
nor U21245 (N_21245,N_20414,N_20936);
and U21246 (N_21246,N_20688,N_20172);
nand U21247 (N_21247,N_20841,N_20824);
xnor U21248 (N_21248,N_20935,N_20180);
nor U21249 (N_21249,N_20583,N_20769);
and U21250 (N_21250,N_20058,N_20628);
and U21251 (N_21251,N_20480,N_20063);
nand U21252 (N_21252,N_20693,N_20668);
nand U21253 (N_21253,N_20495,N_20880);
nor U21254 (N_21254,N_20252,N_20435);
xor U21255 (N_21255,N_20866,N_20680);
xnor U21256 (N_21256,N_20723,N_20796);
nor U21257 (N_21257,N_20397,N_20419);
nor U21258 (N_21258,N_20263,N_20543);
nor U21259 (N_21259,N_20601,N_20819);
and U21260 (N_21260,N_20597,N_20620);
xor U21261 (N_21261,N_20284,N_20016);
or U21262 (N_21262,N_20121,N_20811);
and U21263 (N_21263,N_20881,N_20297);
or U21264 (N_21264,N_20279,N_20633);
or U21265 (N_21265,N_20968,N_20179);
xnor U21266 (N_21266,N_20169,N_20826);
or U21267 (N_21267,N_20123,N_20926);
nor U21268 (N_21268,N_20677,N_20049);
xor U21269 (N_21269,N_20110,N_20226);
and U21270 (N_21270,N_20411,N_20294);
or U21271 (N_21271,N_20491,N_20850);
nand U21272 (N_21272,N_20590,N_20657);
nor U21273 (N_21273,N_20171,N_20471);
nand U21274 (N_21274,N_20066,N_20948);
or U21275 (N_21275,N_20852,N_20211);
nor U21276 (N_21276,N_20330,N_20658);
nor U21277 (N_21277,N_20019,N_20479);
nor U21278 (N_21278,N_20600,N_20571);
or U21279 (N_21279,N_20477,N_20405);
nor U21280 (N_21280,N_20360,N_20445);
nor U21281 (N_21281,N_20302,N_20422);
xor U21282 (N_21282,N_20125,N_20377);
nor U21283 (N_21283,N_20369,N_20427);
nand U21284 (N_21284,N_20280,N_20441);
nand U21285 (N_21285,N_20519,N_20980);
or U21286 (N_21286,N_20090,N_20966);
nor U21287 (N_21287,N_20320,N_20809);
or U21288 (N_21288,N_20175,N_20442);
or U21289 (N_21289,N_20466,N_20412);
nor U21290 (N_21290,N_20244,N_20508);
and U21291 (N_21291,N_20549,N_20318);
nand U21292 (N_21292,N_20605,N_20960);
nand U21293 (N_21293,N_20209,N_20713);
xor U21294 (N_21294,N_20553,N_20515);
and U21295 (N_21295,N_20822,N_20740);
nor U21296 (N_21296,N_20877,N_20379);
nand U21297 (N_21297,N_20036,N_20057);
and U21298 (N_21298,N_20467,N_20448);
nor U21299 (N_21299,N_20304,N_20281);
nand U21300 (N_21300,N_20872,N_20277);
nand U21301 (N_21301,N_20336,N_20525);
or U21302 (N_21302,N_20712,N_20354);
xnor U21303 (N_21303,N_20520,N_20347);
nand U21304 (N_21304,N_20368,N_20685);
xnor U21305 (N_21305,N_20089,N_20256);
and U21306 (N_21306,N_20857,N_20146);
and U21307 (N_21307,N_20105,N_20183);
and U21308 (N_21308,N_20343,N_20150);
nand U21309 (N_21309,N_20359,N_20518);
nor U21310 (N_21310,N_20174,N_20095);
or U21311 (N_21311,N_20795,N_20659);
nand U21312 (N_21312,N_20410,N_20378);
nor U21313 (N_21313,N_20143,N_20151);
and U21314 (N_21314,N_20548,N_20989);
xor U21315 (N_21315,N_20581,N_20637);
and U21316 (N_21316,N_20941,N_20732);
nor U21317 (N_21317,N_20315,N_20602);
nand U21318 (N_21318,N_20465,N_20864);
xor U21319 (N_21319,N_20913,N_20385);
nor U21320 (N_21320,N_20670,N_20843);
or U21321 (N_21321,N_20108,N_20463);
nor U21322 (N_21322,N_20898,N_20193);
or U21323 (N_21323,N_20064,N_20370);
or U21324 (N_21324,N_20552,N_20262);
nand U21325 (N_21325,N_20883,N_20160);
nor U21326 (N_21326,N_20947,N_20168);
nor U21327 (N_21327,N_20617,N_20182);
or U21328 (N_21328,N_20903,N_20556);
and U21329 (N_21329,N_20818,N_20868);
or U21330 (N_21330,N_20537,N_20024);
nand U21331 (N_21331,N_20958,N_20579);
or U21332 (N_21332,N_20894,N_20345);
and U21333 (N_21333,N_20794,N_20494);
and U21334 (N_21334,N_20748,N_20338);
xor U21335 (N_21335,N_20166,N_20488);
xor U21336 (N_21336,N_20346,N_20808);
and U21337 (N_21337,N_20920,N_20998);
or U21338 (N_21338,N_20500,N_20788);
xnor U21339 (N_21339,N_20871,N_20560);
and U21340 (N_21340,N_20457,N_20652);
and U21341 (N_21341,N_20594,N_20714);
and U21342 (N_21342,N_20006,N_20621);
xor U21343 (N_21343,N_20037,N_20799);
nand U21344 (N_21344,N_20365,N_20271);
xor U21345 (N_21345,N_20694,N_20699);
or U21346 (N_21346,N_20048,N_20535);
nor U21347 (N_21347,N_20062,N_20891);
nand U21348 (N_21348,N_20439,N_20775);
or U21349 (N_21349,N_20388,N_20203);
or U21350 (N_21350,N_20317,N_20060);
nor U21351 (N_21351,N_20776,N_20645);
or U21352 (N_21352,N_20366,N_20273);
or U21353 (N_21353,N_20889,N_20946);
xor U21354 (N_21354,N_20106,N_20623);
and U21355 (N_21355,N_20173,N_20923);
nand U21356 (N_21356,N_20744,N_20858);
xor U21357 (N_21357,N_20323,N_20232);
and U21358 (N_21358,N_20507,N_20678);
xor U21359 (N_21359,N_20402,N_20939);
xor U21360 (N_21360,N_20912,N_20956);
and U21361 (N_21361,N_20771,N_20710);
xnor U21362 (N_21362,N_20820,N_20342);
nand U21363 (N_21363,N_20626,N_20844);
nand U21364 (N_21364,N_20719,N_20052);
xnor U21365 (N_21365,N_20622,N_20124);
nand U21366 (N_21366,N_20741,N_20578);
nor U21367 (N_21367,N_20830,N_20949);
or U21368 (N_21368,N_20107,N_20235);
nor U21369 (N_21369,N_20053,N_20417);
nor U21370 (N_21370,N_20961,N_20126);
xor U21371 (N_21371,N_20371,N_20854);
nand U21372 (N_21372,N_20885,N_20308);
nand U21373 (N_21373,N_20532,N_20505);
or U21374 (N_21374,N_20928,N_20849);
or U21375 (N_21375,N_20736,N_20756);
nor U21376 (N_21376,N_20470,N_20576);
xor U21377 (N_21377,N_20391,N_20625);
or U21378 (N_21378,N_20190,N_20967);
xor U21379 (N_21379,N_20403,N_20498);
nor U21380 (N_21380,N_20484,N_20916);
xnor U21381 (N_21381,N_20181,N_20971);
or U21382 (N_21382,N_20258,N_20437);
or U21383 (N_21383,N_20207,N_20127);
or U21384 (N_21384,N_20213,N_20636);
nand U21385 (N_21385,N_20925,N_20975);
xnor U21386 (N_21386,N_20017,N_20787);
xor U21387 (N_21387,N_20386,N_20908);
or U21388 (N_21388,N_20005,N_20754);
or U21389 (N_21389,N_20339,N_20709);
nand U21390 (N_21390,N_20779,N_20240);
or U21391 (N_21391,N_20458,N_20079);
or U21392 (N_21392,N_20521,N_20896);
and U21393 (N_21393,N_20189,N_20117);
nor U21394 (N_21394,N_20344,N_20661);
nand U21395 (N_21395,N_20914,N_20434);
nand U21396 (N_21396,N_20927,N_20113);
nand U21397 (N_21397,N_20390,N_20570);
and U21398 (N_21398,N_20316,N_20531);
or U21399 (N_21399,N_20875,N_20416);
nand U21400 (N_21400,N_20991,N_20236);
xor U21401 (N_21401,N_20523,N_20616);
and U21402 (N_21402,N_20453,N_20247);
nor U21403 (N_21403,N_20669,N_20142);
xnor U21404 (N_21404,N_20558,N_20009);
and U21405 (N_21405,N_20807,N_20829);
xor U21406 (N_21406,N_20930,N_20703);
xor U21407 (N_21407,N_20272,N_20631);
nand U21408 (N_21408,N_20080,N_20813);
nor U21409 (N_21409,N_20072,N_20114);
or U21410 (N_21410,N_20134,N_20785);
or U21411 (N_21411,N_20309,N_20768);
or U21412 (N_21412,N_20007,N_20326);
nand U21413 (N_21413,N_20904,N_20782);
and U21414 (N_21414,N_20910,N_20705);
nand U21415 (N_21415,N_20223,N_20679);
nand U21416 (N_21416,N_20689,N_20298);
xnor U21417 (N_21417,N_20161,N_20094);
or U21418 (N_21418,N_20387,N_20167);
and U21419 (N_21419,N_20790,N_20147);
and U21420 (N_21420,N_20188,N_20522);
nor U21421 (N_21421,N_20611,N_20381);
nand U21422 (N_21422,N_20792,N_20701);
nor U21423 (N_21423,N_20587,N_20335);
nor U21424 (N_21424,N_20141,N_20027);
nand U21425 (N_21425,N_20915,N_20644);
nand U21426 (N_21426,N_20675,N_20282);
nor U21427 (N_21427,N_20615,N_20472);
nand U21428 (N_21428,N_20267,N_20201);
and U21429 (N_21429,N_20238,N_20451);
and U21430 (N_21430,N_20533,N_20950);
xnor U21431 (N_21431,N_20087,N_20643);
nand U21432 (N_21432,N_20730,N_20654);
nor U21433 (N_21433,N_20131,N_20501);
and U21434 (N_21434,N_20029,N_20091);
nor U21435 (N_21435,N_20697,N_20707);
xor U21436 (N_21436,N_20109,N_20119);
nand U21437 (N_21437,N_20195,N_20513);
nand U21438 (N_21438,N_20356,N_20596);
nor U21439 (N_21439,N_20398,N_20739);
nand U21440 (N_21440,N_20348,N_20624);
nand U21441 (N_21441,N_20406,N_20002);
or U21442 (N_21442,N_20747,N_20333);
nor U21443 (N_21443,N_20627,N_20306);
xor U21444 (N_21444,N_20400,N_20456);
nand U21445 (N_21445,N_20395,N_20319);
nor U21446 (N_21446,N_20577,N_20046);
xor U21447 (N_21447,N_20917,N_20837);
nand U21448 (N_21448,N_20539,N_20944);
nand U21449 (N_21449,N_20374,N_20010);
nor U21450 (N_21450,N_20257,N_20056);
nand U21451 (N_21451,N_20030,N_20510);
or U21452 (N_21452,N_20399,N_20328);
and U21453 (N_21453,N_20246,N_20292);
nor U21454 (N_21454,N_20459,N_20184);
nand U21455 (N_21455,N_20478,N_20863);
or U21456 (N_21456,N_20695,N_20482);
and U21457 (N_21457,N_20976,N_20716);
nand U21458 (N_21458,N_20065,N_20664);
nor U21459 (N_21459,N_20951,N_20814);
nand U21460 (N_21460,N_20311,N_20444);
nand U21461 (N_21461,N_20584,N_20957);
and U21462 (N_21462,N_20268,N_20122);
or U21463 (N_21463,N_20641,N_20728);
and U21464 (N_21464,N_20389,N_20210);
xnor U21465 (N_21465,N_20987,N_20129);
and U21466 (N_21466,N_20565,N_20248);
xnor U21467 (N_21467,N_20293,N_20575);
xnor U21468 (N_21468,N_20767,N_20014);
xor U21469 (N_21469,N_20738,N_20706);
xnor U21470 (N_21470,N_20490,N_20111);
nand U21471 (N_21471,N_20337,N_20547);
nand U21472 (N_21472,N_20899,N_20100);
nand U21473 (N_21473,N_20554,N_20752);
and U21474 (N_21474,N_20735,N_20322);
nand U21475 (N_21475,N_20528,N_20846);
nand U21476 (N_21476,N_20540,N_20817);
nor U21477 (N_21477,N_20227,N_20276);
nand U21478 (N_21478,N_20073,N_20873);
nand U21479 (N_21479,N_20154,N_20102);
nor U21480 (N_21480,N_20924,N_20979);
or U21481 (N_21481,N_20187,N_20640);
xor U21482 (N_21482,N_20599,N_20897);
and U21483 (N_21483,N_20541,N_20334);
xor U21484 (N_21484,N_20649,N_20130);
nor U21485 (N_21485,N_20758,N_20815);
xor U21486 (N_21486,N_20148,N_20692);
or U21487 (N_21487,N_20217,N_20618);
xnor U21488 (N_21488,N_20219,N_20996);
nand U21489 (N_21489,N_20321,N_20493);
xor U21490 (N_21490,N_20816,N_20229);
nand U21491 (N_21491,N_20156,N_20039);
and U21492 (N_21492,N_20313,N_20945);
nand U21493 (N_21493,N_20938,N_20886);
xnor U21494 (N_21494,N_20096,N_20138);
and U21495 (N_21495,N_20582,N_20396);
or U21496 (N_21496,N_20764,N_20869);
nand U21497 (N_21497,N_20757,N_20059);
nand U21498 (N_21498,N_20717,N_20233);
nor U21499 (N_21499,N_20646,N_20503);
or U21500 (N_21500,N_20870,N_20788);
xnor U21501 (N_21501,N_20604,N_20822);
nor U21502 (N_21502,N_20908,N_20002);
or U21503 (N_21503,N_20727,N_20402);
xor U21504 (N_21504,N_20696,N_20024);
nor U21505 (N_21505,N_20401,N_20013);
xnor U21506 (N_21506,N_20501,N_20123);
xnor U21507 (N_21507,N_20607,N_20495);
or U21508 (N_21508,N_20183,N_20755);
or U21509 (N_21509,N_20794,N_20027);
nor U21510 (N_21510,N_20342,N_20948);
or U21511 (N_21511,N_20669,N_20040);
nor U21512 (N_21512,N_20578,N_20150);
xor U21513 (N_21513,N_20241,N_20635);
nor U21514 (N_21514,N_20301,N_20435);
and U21515 (N_21515,N_20504,N_20103);
nand U21516 (N_21516,N_20001,N_20709);
nand U21517 (N_21517,N_20992,N_20388);
or U21518 (N_21518,N_20414,N_20240);
and U21519 (N_21519,N_20497,N_20580);
nand U21520 (N_21520,N_20191,N_20909);
nand U21521 (N_21521,N_20567,N_20018);
xnor U21522 (N_21522,N_20496,N_20487);
nor U21523 (N_21523,N_20715,N_20993);
or U21524 (N_21524,N_20637,N_20622);
nor U21525 (N_21525,N_20852,N_20677);
and U21526 (N_21526,N_20991,N_20961);
and U21527 (N_21527,N_20307,N_20866);
nor U21528 (N_21528,N_20198,N_20279);
nor U21529 (N_21529,N_20680,N_20286);
and U21530 (N_21530,N_20125,N_20209);
xor U21531 (N_21531,N_20135,N_20803);
nand U21532 (N_21532,N_20516,N_20932);
or U21533 (N_21533,N_20523,N_20197);
or U21534 (N_21534,N_20258,N_20462);
and U21535 (N_21535,N_20687,N_20443);
and U21536 (N_21536,N_20517,N_20398);
nor U21537 (N_21537,N_20878,N_20833);
or U21538 (N_21538,N_20016,N_20811);
xor U21539 (N_21539,N_20916,N_20286);
or U21540 (N_21540,N_20554,N_20529);
or U21541 (N_21541,N_20264,N_20215);
nand U21542 (N_21542,N_20497,N_20768);
or U21543 (N_21543,N_20869,N_20249);
nor U21544 (N_21544,N_20851,N_20034);
and U21545 (N_21545,N_20057,N_20154);
nor U21546 (N_21546,N_20030,N_20623);
xnor U21547 (N_21547,N_20471,N_20373);
xnor U21548 (N_21548,N_20630,N_20623);
nor U21549 (N_21549,N_20460,N_20571);
xor U21550 (N_21550,N_20413,N_20173);
xor U21551 (N_21551,N_20748,N_20833);
and U21552 (N_21552,N_20280,N_20468);
nand U21553 (N_21553,N_20053,N_20717);
nand U21554 (N_21554,N_20264,N_20624);
or U21555 (N_21555,N_20655,N_20716);
or U21556 (N_21556,N_20834,N_20040);
and U21557 (N_21557,N_20294,N_20782);
nor U21558 (N_21558,N_20162,N_20146);
or U21559 (N_21559,N_20883,N_20290);
and U21560 (N_21560,N_20925,N_20301);
xnor U21561 (N_21561,N_20231,N_20201);
nand U21562 (N_21562,N_20571,N_20014);
nor U21563 (N_21563,N_20161,N_20148);
and U21564 (N_21564,N_20883,N_20645);
xnor U21565 (N_21565,N_20506,N_20717);
or U21566 (N_21566,N_20726,N_20566);
and U21567 (N_21567,N_20276,N_20485);
or U21568 (N_21568,N_20868,N_20008);
and U21569 (N_21569,N_20601,N_20046);
or U21570 (N_21570,N_20556,N_20033);
nand U21571 (N_21571,N_20510,N_20933);
or U21572 (N_21572,N_20180,N_20947);
nor U21573 (N_21573,N_20054,N_20412);
and U21574 (N_21574,N_20226,N_20172);
xor U21575 (N_21575,N_20063,N_20768);
nand U21576 (N_21576,N_20476,N_20163);
nor U21577 (N_21577,N_20151,N_20492);
or U21578 (N_21578,N_20911,N_20619);
nor U21579 (N_21579,N_20178,N_20845);
xnor U21580 (N_21580,N_20218,N_20361);
or U21581 (N_21581,N_20219,N_20497);
xor U21582 (N_21582,N_20837,N_20367);
or U21583 (N_21583,N_20811,N_20328);
nor U21584 (N_21584,N_20639,N_20459);
and U21585 (N_21585,N_20320,N_20547);
or U21586 (N_21586,N_20596,N_20035);
nand U21587 (N_21587,N_20483,N_20968);
nand U21588 (N_21588,N_20378,N_20402);
and U21589 (N_21589,N_20462,N_20330);
xor U21590 (N_21590,N_20301,N_20681);
or U21591 (N_21591,N_20256,N_20924);
nor U21592 (N_21592,N_20184,N_20813);
nor U21593 (N_21593,N_20520,N_20079);
nor U21594 (N_21594,N_20169,N_20847);
nor U21595 (N_21595,N_20926,N_20639);
xor U21596 (N_21596,N_20231,N_20247);
and U21597 (N_21597,N_20655,N_20888);
or U21598 (N_21598,N_20431,N_20062);
or U21599 (N_21599,N_20608,N_20984);
or U21600 (N_21600,N_20278,N_20520);
or U21601 (N_21601,N_20498,N_20981);
or U21602 (N_21602,N_20515,N_20110);
and U21603 (N_21603,N_20432,N_20416);
xnor U21604 (N_21604,N_20943,N_20364);
or U21605 (N_21605,N_20292,N_20751);
nand U21606 (N_21606,N_20079,N_20946);
and U21607 (N_21607,N_20742,N_20014);
xor U21608 (N_21608,N_20825,N_20385);
and U21609 (N_21609,N_20632,N_20541);
and U21610 (N_21610,N_20549,N_20365);
and U21611 (N_21611,N_20842,N_20195);
xor U21612 (N_21612,N_20616,N_20036);
and U21613 (N_21613,N_20946,N_20552);
xor U21614 (N_21614,N_20162,N_20860);
xnor U21615 (N_21615,N_20287,N_20608);
xnor U21616 (N_21616,N_20723,N_20560);
and U21617 (N_21617,N_20038,N_20107);
and U21618 (N_21618,N_20770,N_20182);
nand U21619 (N_21619,N_20870,N_20909);
xor U21620 (N_21620,N_20467,N_20580);
and U21621 (N_21621,N_20013,N_20667);
nand U21622 (N_21622,N_20740,N_20023);
nor U21623 (N_21623,N_20726,N_20138);
nor U21624 (N_21624,N_20629,N_20219);
or U21625 (N_21625,N_20173,N_20340);
and U21626 (N_21626,N_20130,N_20337);
xor U21627 (N_21627,N_20808,N_20583);
xor U21628 (N_21628,N_20111,N_20343);
nand U21629 (N_21629,N_20850,N_20770);
xnor U21630 (N_21630,N_20232,N_20643);
nor U21631 (N_21631,N_20514,N_20466);
nand U21632 (N_21632,N_20772,N_20795);
nor U21633 (N_21633,N_20323,N_20683);
nor U21634 (N_21634,N_20382,N_20607);
xor U21635 (N_21635,N_20025,N_20200);
or U21636 (N_21636,N_20690,N_20086);
nor U21637 (N_21637,N_20924,N_20986);
xnor U21638 (N_21638,N_20346,N_20689);
nor U21639 (N_21639,N_20912,N_20043);
or U21640 (N_21640,N_20914,N_20123);
nor U21641 (N_21641,N_20296,N_20757);
nand U21642 (N_21642,N_20845,N_20991);
or U21643 (N_21643,N_20476,N_20060);
nor U21644 (N_21644,N_20129,N_20198);
nand U21645 (N_21645,N_20078,N_20505);
and U21646 (N_21646,N_20888,N_20855);
nor U21647 (N_21647,N_20253,N_20260);
and U21648 (N_21648,N_20352,N_20509);
xnor U21649 (N_21649,N_20517,N_20239);
and U21650 (N_21650,N_20055,N_20051);
nor U21651 (N_21651,N_20210,N_20567);
nor U21652 (N_21652,N_20838,N_20569);
nand U21653 (N_21653,N_20255,N_20545);
and U21654 (N_21654,N_20909,N_20453);
nor U21655 (N_21655,N_20390,N_20561);
xnor U21656 (N_21656,N_20509,N_20478);
or U21657 (N_21657,N_20803,N_20310);
nand U21658 (N_21658,N_20882,N_20459);
or U21659 (N_21659,N_20297,N_20634);
and U21660 (N_21660,N_20294,N_20945);
or U21661 (N_21661,N_20562,N_20146);
nor U21662 (N_21662,N_20820,N_20494);
and U21663 (N_21663,N_20755,N_20187);
nand U21664 (N_21664,N_20094,N_20611);
xor U21665 (N_21665,N_20965,N_20449);
xnor U21666 (N_21666,N_20020,N_20695);
nand U21667 (N_21667,N_20417,N_20390);
or U21668 (N_21668,N_20828,N_20431);
xnor U21669 (N_21669,N_20759,N_20104);
nor U21670 (N_21670,N_20149,N_20300);
or U21671 (N_21671,N_20388,N_20969);
or U21672 (N_21672,N_20463,N_20265);
nor U21673 (N_21673,N_20301,N_20401);
nand U21674 (N_21674,N_20964,N_20149);
xor U21675 (N_21675,N_20474,N_20307);
and U21676 (N_21676,N_20817,N_20580);
nor U21677 (N_21677,N_20539,N_20292);
nor U21678 (N_21678,N_20519,N_20981);
and U21679 (N_21679,N_20037,N_20409);
xnor U21680 (N_21680,N_20972,N_20839);
and U21681 (N_21681,N_20190,N_20714);
nand U21682 (N_21682,N_20537,N_20205);
nand U21683 (N_21683,N_20478,N_20041);
or U21684 (N_21684,N_20267,N_20116);
or U21685 (N_21685,N_20902,N_20140);
and U21686 (N_21686,N_20310,N_20314);
nand U21687 (N_21687,N_20238,N_20974);
xor U21688 (N_21688,N_20235,N_20403);
and U21689 (N_21689,N_20220,N_20890);
nand U21690 (N_21690,N_20827,N_20079);
and U21691 (N_21691,N_20666,N_20191);
and U21692 (N_21692,N_20874,N_20734);
nor U21693 (N_21693,N_20871,N_20954);
and U21694 (N_21694,N_20538,N_20466);
or U21695 (N_21695,N_20942,N_20400);
xnor U21696 (N_21696,N_20920,N_20865);
xnor U21697 (N_21697,N_20305,N_20321);
nor U21698 (N_21698,N_20340,N_20332);
and U21699 (N_21699,N_20157,N_20418);
nand U21700 (N_21700,N_20268,N_20086);
and U21701 (N_21701,N_20176,N_20154);
or U21702 (N_21702,N_20374,N_20953);
xor U21703 (N_21703,N_20467,N_20672);
and U21704 (N_21704,N_20996,N_20005);
and U21705 (N_21705,N_20975,N_20998);
and U21706 (N_21706,N_20962,N_20305);
xnor U21707 (N_21707,N_20602,N_20034);
nand U21708 (N_21708,N_20837,N_20968);
nand U21709 (N_21709,N_20448,N_20343);
nand U21710 (N_21710,N_20045,N_20851);
xnor U21711 (N_21711,N_20053,N_20729);
xnor U21712 (N_21712,N_20263,N_20347);
or U21713 (N_21713,N_20860,N_20689);
xnor U21714 (N_21714,N_20742,N_20186);
xnor U21715 (N_21715,N_20182,N_20847);
nand U21716 (N_21716,N_20672,N_20327);
or U21717 (N_21717,N_20671,N_20695);
nor U21718 (N_21718,N_20585,N_20264);
or U21719 (N_21719,N_20955,N_20252);
xnor U21720 (N_21720,N_20585,N_20135);
and U21721 (N_21721,N_20921,N_20919);
xor U21722 (N_21722,N_20173,N_20812);
xor U21723 (N_21723,N_20613,N_20581);
and U21724 (N_21724,N_20354,N_20895);
or U21725 (N_21725,N_20521,N_20716);
and U21726 (N_21726,N_20705,N_20950);
nor U21727 (N_21727,N_20048,N_20406);
or U21728 (N_21728,N_20935,N_20883);
nor U21729 (N_21729,N_20428,N_20890);
or U21730 (N_21730,N_20242,N_20568);
or U21731 (N_21731,N_20975,N_20954);
and U21732 (N_21732,N_20171,N_20607);
xnor U21733 (N_21733,N_20300,N_20609);
and U21734 (N_21734,N_20485,N_20649);
xor U21735 (N_21735,N_20286,N_20010);
nor U21736 (N_21736,N_20574,N_20340);
or U21737 (N_21737,N_20114,N_20386);
and U21738 (N_21738,N_20116,N_20438);
nor U21739 (N_21739,N_20745,N_20351);
nand U21740 (N_21740,N_20391,N_20898);
and U21741 (N_21741,N_20667,N_20946);
nor U21742 (N_21742,N_20967,N_20571);
xor U21743 (N_21743,N_20294,N_20535);
or U21744 (N_21744,N_20699,N_20339);
and U21745 (N_21745,N_20047,N_20098);
xor U21746 (N_21746,N_20255,N_20015);
and U21747 (N_21747,N_20649,N_20607);
or U21748 (N_21748,N_20704,N_20590);
nand U21749 (N_21749,N_20456,N_20225);
nor U21750 (N_21750,N_20849,N_20518);
and U21751 (N_21751,N_20908,N_20173);
nand U21752 (N_21752,N_20129,N_20727);
xor U21753 (N_21753,N_20720,N_20377);
and U21754 (N_21754,N_20391,N_20852);
nand U21755 (N_21755,N_20428,N_20165);
nor U21756 (N_21756,N_20404,N_20288);
nor U21757 (N_21757,N_20783,N_20277);
and U21758 (N_21758,N_20231,N_20281);
or U21759 (N_21759,N_20348,N_20921);
xor U21760 (N_21760,N_20592,N_20855);
and U21761 (N_21761,N_20296,N_20286);
xnor U21762 (N_21762,N_20138,N_20415);
nand U21763 (N_21763,N_20325,N_20216);
nor U21764 (N_21764,N_20844,N_20695);
or U21765 (N_21765,N_20458,N_20897);
xnor U21766 (N_21766,N_20637,N_20714);
nor U21767 (N_21767,N_20768,N_20574);
nand U21768 (N_21768,N_20223,N_20113);
nor U21769 (N_21769,N_20162,N_20153);
xnor U21770 (N_21770,N_20161,N_20181);
nor U21771 (N_21771,N_20504,N_20769);
nor U21772 (N_21772,N_20739,N_20024);
nand U21773 (N_21773,N_20596,N_20105);
or U21774 (N_21774,N_20979,N_20563);
xnor U21775 (N_21775,N_20321,N_20475);
xnor U21776 (N_21776,N_20829,N_20828);
nor U21777 (N_21777,N_20512,N_20687);
nor U21778 (N_21778,N_20920,N_20569);
or U21779 (N_21779,N_20622,N_20446);
xnor U21780 (N_21780,N_20539,N_20044);
nand U21781 (N_21781,N_20464,N_20468);
nor U21782 (N_21782,N_20753,N_20207);
or U21783 (N_21783,N_20546,N_20699);
or U21784 (N_21784,N_20413,N_20447);
or U21785 (N_21785,N_20657,N_20768);
or U21786 (N_21786,N_20516,N_20501);
and U21787 (N_21787,N_20047,N_20559);
and U21788 (N_21788,N_20997,N_20934);
nor U21789 (N_21789,N_20045,N_20899);
xor U21790 (N_21790,N_20827,N_20584);
xor U21791 (N_21791,N_20955,N_20664);
nand U21792 (N_21792,N_20296,N_20032);
nor U21793 (N_21793,N_20133,N_20916);
or U21794 (N_21794,N_20394,N_20190);
nand U21795 (N_21795,N_20323,N_20817);
nand U21796 (N_21796,N_20575,N_20827);
nor U21797 (N_21797,N_20466,N_20499);
and U21798 (N_21798,N_20094,N_20384);
xnor U21799 (N_21799,N_20215,N_20893);
xor U21800 (N_21800,N_20707,N_20603);
nand U21801 (N_21801,N_20101,N_20236);
xor U21802 (N_21802,N_20168,N_20435);
or U21803 (N_21803,N_20067,N_20422);
or U21804 (N_21804,N_20815,N_20637);
and U21805 (N_21805,N_20385,N_20716);
or U21806 (N_21806,N_20251,N_20753);
or U21807 (N_21807,N_20666,N_20453);
nand U21808 (N_21808,N_20068,N_20637);
nand U21809 (N_21809,N_20443,N_20485);
nor U21810 (N_21810,N_20231,N_20751);
and U21811 (N_21811,N_20272,N_20765);
or U21812 (N_21812,N_20711,N_20785);
xor U21813 (N_21813,N_20657,N_20436);
or U21814 (N_21814,N_20113,N_20331);
xor U21815 (N_21815,N_20698,N_20240);
nor U21816 (N_21816,N_20148,N_20600);
nor U21817 (N_21817,N_20192,N_20814);
or U21818 (N_21818,N_20011,N_20139);
xnor U21819 (N_21819,N_20533,N_20494);
nand U21820 (N_21820,N_20100,N_20432);
nor U21821 (N_21821,N_20576,N_20861);
xor U21822 (N_21822,N_20539,N_20482);
xnor U21823 (N_21823,N_20706,N_20283);
or U21824 (N_21824,N_20895,N_20139);
nand U21825 (N_21825,N_20875,N_20058);
nand U21826 (N_21826,N_20294,N_20179);
or U21827 (N_21827,N_20378,N_20569);
xor U21828 (N_21828,N_20692,N_20843);
xnor U21829 (N_21829,N_20269,N_20287);
nor U21830 (N_21830,N_20226,N_20626);
and U21831 (N_21831,N_20508,N_20646);
and U21832 (N_21832,N_20448,N_20457);
or U21833 (N_21833,N_20596,N_20895);
nand U21834 (N_21834,N_20101,N_20749);
nor U21835 (N_21835,N_20288,N_20075);
nand U21836 (N_21836,N_20624,N_20391);
nand U21837 (N_21837,N_20705,N_20389);
or U21838 (N_21838,N_20572,N_20323);
or U21839 (N_21839,N_20009,N_20944);
nor U21840 (N_21840,N_20586,N_20311);
nand U21841 (N_21841,N_20926,N_20490);
xnor U21842 (N_21842,N_20735,N_20328);
nor U21843 (N_21843,N_20942,N_20063);
nor U21844 (N_21844,N_20094,N_20766);
nor U21845 (N_21845,N_20224,N_20005);
and U21846 (N_21846,N_20868,N_20120);
or U21847 (N_21847,N_20989,N_20096);
xor U21848 (N_21848,N_20616,N_20679);
xor U21849 (N_21849,N_20781,N_20084);
nand U21850 (N_21850,N_20497,N_20201);
and U21851 (N_21851,N_20029,N_20517);
xnor U21852 (N_21852,N_20991,N_20704);
xnor U21853 (N_21853,N_20068,N_20699);
nand U21854 (N_21854,N_20136,N_20220);
and U21855 (N_21855,N_20531,N_20890);
nor U21856 (N_21856,N_20283,N_20843);
and U21857 (N_21857,N_20346,N_20565);
xor U21858 (N_21858,N_20136,N_20570);
or U21859 (N_21859,N_20240,N_20152);
and U21860 (N_21860,N_20024,N_20646);
and U21861 (N_21861,N_20325,N_20338);
or U21862 (N_21862,N_20398,N_20922);
or U21863 (N_21863,N_20343,N_20134);
or U21864 (N_21864,N_20052,N_20717);
xor U21865 (N_21865,N_20965,N_20575);
xor U21866 (N_21866,N_20765,N_20321);
xnor U21867 (N_21867,N_20772,N_20147);
nand U21868 (N_21868,N_20324,N_20483);
nand U21869 (N_21869,N_20912,N_20838);
or U21870 (N_21870,N_20322,N_20512);
or U21871 (N_21871,N_20429,N_20135);
or U21872 (N_21872,N_20433,N_20708);
nand U21873 (N_21873,N_20535,N_20129);
and U21874 (N_21874,N_20162,N_20529);
nand U21875 (N_21875,N_20905,N_20578);
nand U21876 (N_21876,N_20844,N_20484);
xor U21877 (N_21877,N_20033,N_20375);
or U21878 (N_21878,N_20639,N_20199);
nor U21879 (N_21879,N_20610,N_20113);
nand U21880 (N_21880,N_20043,N_20513);
and U21881 (N_21881,N_20396,N_20977);
nand U21882 (N_21882,N_20914,N_20992);
nor U21883 (N_21883,N_20830,N_20093);
nor U21884 (N_21884,N_20303,N_20216);
xnor U21885 (N_21885,N_20682,N_20272);
or U21886 (N_21886,N_20958,N_20823);
and U21887 (N_21887,N_20229,N_20381);
or U21888 (N_21888,N_20749,N_20744);
nor U21889 (N_21889,N_20245,N_20232);
nor U21890 (N_21890,N_20764,N_20099);
or U21891 (N_21891,N_20091,N_20323);
nand U21892 (N_21892,N_20150,N_20883);
or U21893 (N_21893,N_20414,N_20883);
nand U21894 (N_21894,N_20475,N_20602);
nor U21895 (N_21895,N_20881,N_20252);
nor U21896 (N_21896,N_20701,N_20365);
and U21897 (N_21897,N_20492,N_20617);
and U21898 (N_21898,N_20776,N_20168);
or U21899 (N_21899,N_20635,N_20055);
xor U21900 (N_21900,N_20007,N_20459);
or U21901 (N_21901,N_20066,N_20751);
xnor U21902 (N_21902,N_20510,N_20081);
xor U21903 (N_21903,N_20426,N_20051);
or U21904 (N_21904,N_20316,N_20911);
or U21905 (N_21905,N_20139,N_20198);
nor U21906 (N_21906,N_20957,N_20780);
xnor U21907 (N_21907,N_20973,N_20070);
nor U21908 (N_21908,N_20853,N_20103);
or U21909 (N_21909,N_20449,N_20151);
xnor U21910 (N_21910,N_20195,N_20514);
nand U21911 (N_21911,N_20449,N_20126);
nand U21912 (N_21912,N_20362,N_20415);
xnor U21913 (N_21913,N_20004,N_20140);
nor U21914 (N_21914,N_20216,N_20914);
and U21915 (N_21915,N_20253,N_20011);
nand U21916 (N_21916,N_20596,N_20539);
nor U21917 (N_21917,N_20233,N_20893);
and U21918 (N_21918,N_20340,N_20076);
or U21919 (N_21919,N_20999,N_20560);
xor U21920 (N_21920,N_20767,N_20594);
or U21921 (N_21921,N_20849,N_20390);
and U21922 (N_21922,N_20275,N_20805);
nor U21923 (N_21923,N_20440,N_20652);
and U21924 (N_21924,N_20041,N_20174);
or U21925 (N_21925,N_20934,N_20437);
or U21926 (N_21926,N_20238,N_20093);
xor U21927 (N_21927,N_20436,N_20246);
or U21928 (N_21928,N_20973,N_20691);
and U21929 (N_21929,N_20295,N_20430);
nor U21930 (N_21930,N_20878,N_20210);
or U21931 (N_21931,N_20147,N_20737);
nand U21932 (N_21932,N_20519,N_20544);
xnor U21933 (N_21933,N_20958,N_20556);
xor U21934 (N_21934,N_20776,N_20047);
nand U21935 (N_21935,N_20127,N_20060);
nor U21936 (N_21936,N_20099,N_20651);
or U21937 (N_21937,N_20985,N_20247);
and U21938 (N_21938,N_20156,N_20953);
xor U21939 (N_21939,N_20877,N_20609);
and U21940 (N_21940,N_20212,N_20325);
and U21941 (N_21941,N_20112,N_20891);
xor U21942 (N_21942,N_20034,N_20248);
nand U21943 (N_21943,N_20606,N_20365);
or U21944 (N_21944,N_20730,N_20954);
nand U21945 (N_21945,N_20908,N_20103);
or U21946 (N_21946,N_20172,N_20573);
nor U21947 (N_21947,N_20933,N_20107);
or U21948 (N_21948,N_20787,N_20845);
nand U21949 (N_21949,N_20386,N_20290);
and U21950 (N_21950,N_20503,N_20112);
and U21951 (N_21951,N_20881,N_20934);
xnor U21952 (N_21952,N_20091,N_20808);
nor U21953 (N_21953,N_20528,N_20540);
nor U21954 (N_21954,N_20489,N_20465);
and U21955 (N_21955,N_20262,N_20829);
and U21956 (N_21956,N_20639,N_20381);
or U21957 (N_21957,N_20284,N_20107);
or U21958 (N_21958,N_20489,N_20241);
nand U21959 (N_21959,N_20618,N_20264);
and U21960 (N_21960,N_20961,N_20248);
xnor U21961 (N_21961,N_20928,N_20130);
nor U21962 (N_21962,N_20905,N_20389);
nor U21963 (N_21963,N_20095,N_20970);
or U21964 (N_21964,N_20801,N_20120);
xnor U21965 (N_21965,N_20201,N_20380);
nand U21966 (N_21966,N_20128,N_20164);
nand U21967 (N_21967,N_20286,N_20712);
xor U21968 (N_21968,N_20213,N_20261);
and U21969 (N_21969,N_20607,N_20465);
nand U21970 (N_21970,N_20691,N_20906);
nor U21971 (N_21971,N_20256,N_20729);
nor U21972 (N_21972,N_20176,N_20387);
or U21973 (N_21973,N_20841,N_20557);
nand U21974 (N_21974,N_20758,N_20217);
or U21975 (N_21975,N_20169,N_20994);
or U21976 (N_21976,N_20568,N_20803);
nand U21977 (N_21977,N_20037,N_20461);
or U21978 (N_21978,N_20925,N_20867);
nand U21979 (N_21979,N_20032,N_20198);
and U21980 (N_21980,N_20884,N_20347);
nor U21981 (N_21981,N_20998,N_20644);
xnor U21982 (N_21982,N_20896,N_20550);
nand U21983 (N_21983,N_20941,N_20283);
nor U21984 (N_21984,N_20141,N_20532);
and U21985 (N_21985,N_20295,N_20452);
nand U21986 (N_21986,N_20201,N_20224);
and U21987 (N_21987,N_20136,N_20573);
and U21988 (N_21988,N_20212,N_20985);
nand U21989 (N_21989,N_20639,N_20947);
nor U21990 (N_21990,N_20948,N_20431);
or U21991 (N_21991,N_20043,N_20468);
nand U21992 (N_21992,N_20468,N_20188);
and U21993 (N_21993,N_20475,N_20119);
xnor U21994 (N_21994,N_20745,N_20176);
xnor U21995 (N_21995,N_20340,N_20380);
nand U21996 (N_21996,N_20464,N_20010);
xor U21997 (N_21997,N_20353,N_20842);
and U21998 (N_21998,N_20322,N_20495);
nor U21999 (N_21999,N_20897,N_20983);
nand U22000 (N_22000,N_21914,N_21773);
xnor U22001 (N_22001,N_21912,N_21780);
nand U22002 (N_22002,N_21365,N_21558);
and U22003 (N_22003,N_21438,N_21772);
xor U22004 (N_22004,N_21147,N_21280);
nor U22005 (N_22005,N_21846,N_21844);
xnor U22006 (N_22006,N_21199,N_21384);
xnor U22007 (N_22007,N_21598,N_21310);
nor U22008 (N_22008,N_21276,N_21983);
nand U22009 (N_22009,N_21560,N_21335);
or U22010 (N_22010,N_21795,N_21273);
nor U22011 (N_22011,N_21179,N_21877);
nand U22012 (N_22012,N_21151,N_21244);
nand U22013 (N_22013,N_21858,N_21981);
nor U22014 (N_22014,N_21348,N_21111);
and U22015 (N_22015,N_21107,N_21488);
nand U22016 (N_22016,N_21727,N_21045);
or U22017 (N_22017,N_21189,N_21415);
or U22018 (N_22018,N_21880,N_21638);
nor U22019 (N_22019,N_21440,N_21177);
xor U22020 (N_22020,N_21832,N_21411);
nand U22021 (N_22021,N_21817,N_21630);
nand U22022 (N_22022,N_21715,N_21896);
nor U22023 (N_22023,N_21661,N_21609);
and U22024 (N_22024,N_21614,N_21432);
xnor U22025 (N_22025,N_21927,N_21682);
nor U22026 (N_22026,N_21929,N_21875);
xor U22027 (N_22027,N_21746,N_21815);
xnor U22028 (N_22028,N_21294,N_21262);
nor U22029 (N_22029,N_21659,N_21651);
nand U22030 (N_22030,N_21302,N_21963);
nor U22031 (N_22031,N_21602,N_21745);
or U22032 (N_22032,N_21368,N_21391);
nand U22033 (N_22033,N_21988,N_21706);
nand U22034 (N_22034,N_21517,N_21737);
nor U22035 (N_22035,N_21545,N_21057);
nand U22036 (N_22036,N_21504,N_21980);
and U22037 (N_22037,N_21325,N_21126);
and U22038 (N_22038,N_21283,N_21489);
xor U22039 (N_22039,N_21864,N_21272);
nor U22040 (N_22040,N_21578,N_21006);
nand U22041 (N_22041,N_21032,N_21627);
or U22042 (N_22042,N_21305,N_21655);
or U22043 (N_22043,N_21732,N_21175);
nor U22044 (N_22044,N_21190,N_21704);
nor U22045 (N_22045,N_21364,N_21689);
or U22046 (N_22046,N_21378,N_21756);
nor U22047 (N_22047,N_21721,N_21758);
xnor U22048 (N_22048,N_21700,N_21785);
or U22049 (N_22049,N_21579,N_21446);
nor U22050 (N_22050,N_21142,N_21643);
and U22051 (N_22051,N_21781,N_21889);
or U22052 (N_22052,N_21991,N_21020);
xor U22053 (N_22053,N_21080,N_21270);
nand U22054 (N_22054,N_21928,N_21100);
xnor U22055 (N_22055,N_21634,N_21185);
or U22056 (N_22056,N_21881,N_21744);
or U22057 (N_22057,N_21334,N_21261);
nand U22058 (N_22058,N_21118,N_21413);
or U22059 (N_22059,N_21347,N_21218);
or U22060 (N_22060,N_21121,N_21385);
and U22061 (N_22061,N_21601,N_21926);
nor U22062 (N_22062,N_21134,N_21469);
xor U22063 (N_22063,N_21580,N_21913);
xnor U22064 (N_22064,N_21074,N_21358);
xnor U22065 (N_22065,N_21725,N_21559);
and U22066 (N_22066,N_21344,N_21550);
nand U22067 (N_22067,N_21998,N_21482);
and U22068 (N_22068,N_21242,N_21122);
nand U22069 (N_22069,N_21872,N_21752);
or U22070 (N_22070,N_21328,N_21128);
or U22071 (N_22071,N_21642,N_21805);
nor U22072 (N_22072,N_21381,N_21342);
and U22073 (N_22073,N_21716,N_21596);
and U22074 (N_22074,N_21571,N_21603);
nor U22075 (N_22075,N_21527,N_21748);
xor U22076 (N_22076,N_21743,N_21339);
or U22077 (N_22077,N_21985,N_21709);
xnor U22078 (N_22078,N_21007,N_21231);
xnor U22079 (N_22079,N_21870,N_21241);
nor U22080 (N_22080,N_21026,N_21309);
xor U22081 (N_22081,N_21388,N_21585);
xor U22082 (N_22082,N_21292,N_21480);
xnor U22083 (N_22083,N_21290,N_21588);
xor U22084 (N_22084,N_21131,N_21996);
xor U22085 (N_22085,N_21589,N_21931);
or U22086 (N_22086,N_21407,N_21546);
and U22087 (N_22087,N_21911,N_21736);
nand U22088 (N_22088,N_21628,N_21573);
xnor U22089 (N_22089,N_21256,N_21897);
xor U22090 (N_22090,N_21572,N_21994);
or U22091 (N_22091,N_21888,N_21629);
or U22092 (N_22092,N_21060,N_21209);
nor U22093 (N_22093,N_21239,N_21949);
and U22094 (N_22094,N_21740,N_21169);
nand U22095 (N_22095,N_21922,N_21769);
or U22096 (N_22096,N_21867,N_21883);
nand U22097 (N_22097,N_21719,N_21813);
and U22098 (N_22098,N_21197,N_21027);
and U22099 (N_22099,N_21308,N_21569);
nor U22100 (N_22100,N_21974,N_21451);
nand U22101 (N_22101,N_21120,N_21022);
and U22102 (N_22102,N_21321,N_21925);
xor U22103 (N_22103,N_21798,N_21252);
nor U22104 (N_22104,N_21072,N_21427);
xor U22105 (N_22105,N_21275,N_21034);
nor U22106 (N_22106,N_21606,N_21054);
or U22107 (N_22107,N_21437,N_21291);
nor U22108 (N_22108,N_21965,N_21257);
xor U22109 (N_22109,N_21729,N_21136);
nor U22110 (N_22110,N_21787,N_21069);
xnor U22111 (N_22111,N_21472,N_21314);
nand U22112 (N_22112,N_21425,N_21238);
and U22113 (N_22113,N_21954,N_21894);
xor U22114 (N_22114,N_21491,N_21502);
or U22115 (N_22115,N_21140,N_21818);
or U22116 (N_22116,N_21675,N_21028);
and U22117 (N_22117,N_21397,N_21948);
or U22118 (N_22118,N_21277,N_21049);
and U22119 (N_22119,N_21935,N_21555);
or U22120 (N_22120,N_21133,N_21821);
and U22121 (N_22121,N_21374,N_21953);
and U22122 (N_22122,N_21899,N_21694);
nor U22123 (N_22123,N_21492,N_21456);
xnor U22124 (N_22124,N_21982,N_21459);
and U22125 (N_22125,N_21208,N_21731);
nor U22126 (N_22126,N_21833,N_21530);
nor U22127 (N_22127,N_21116,N_21848);
nand U22128 (N_22128,N_21874,N_21454);
and U22129 (N_22129,N_21195,N_21157);
and U22130 (N_22130,N_21794,N_21561);
xnor U22131 (N_22131,N_21944,N_21783);
nor U22132 (N_22132,N_21767,N_21916);
xnor U22133 (N_22133,N_21450,N_21264);
or U22134 (N_22134,N_21724,N_21686);
and U22135 (N_22135,N_21387,N_21850);
xor U22136 (N_22136,N_21093,N_21708);
xor U22137 (N_22137,N_21095,N_21105);
nand U22138 (N_22138,N_21876,N_21205);
nand U22139 (N_22139,N_21807,N_21950);
or U22140 (N_22140,N_21905,N_21676);
xor U22141 (N_22141,N_21211,N_21206);
and U22142 (N_22142,N_21350,N_21720);
and U22143 (N_22143,N_21320,N_21371);
nor U22144 (N_22144,N_21849,N_21330);
or U22145 (N_22145,N_21409,N_21011);
nand U22146 (N_22146,N_21673,N_21599);
nor U22147 (N_22147,N_21934,N_21200);
and U22148 (N_22148,N_21019,N_21379);
and U22149 (N_22149,N_21553,N_21827);
nand U22150 (N_22150,N_21386,N_21424);
nor U22151 (N_22151,N_21863,N_21015);
nand U22152 (N_22152,N_21043,N_21376);
and U22153 (N_22153,N_21898,N_21871);
or U22154 (N_22154,N_21298,N_21669);
xnor U22155 (N_22155,N_21021,N_21778);
or U22156 (N_22156,N_21574,N_21796);
nand U22157 (N_22157,N_21741,N_21164);
nor U22158 (N_22158,N_21331,N_21824);
and U22159 (N_22159,N_21056,N_21220);
nand U22160 (N_22160,N_21524,N_21036);
and U22161 (N_22161,N_21969,N_21453);
xor U22162 (N_22162,N_21235,N_21764);
nand U22163 (N_22163,N_21044,N_21367);
and U22164 (N_22164,N_21906,N_21804);
nand U22165 (N_22165,N_21541,N_21964);
or U22166 (N_22166,N_21608,N_21547);
and U22167 (N_22167,N_21542,N_21712);
or U22168 (N_22168,N_21445,N_21611);
xnor U22169 (N_22169,N_21652,N_21198);
nand U22170 (N_22170,N_21016,N_21345);
nor U22171 (N_22171,N_21885,N_21004);
xor U22172 (N_22172,N_21154,N_21228);
and U22173 (N_22173,N_21483,N_21452);
nand U22174 (N_22174,N_21711,N_21058);
nor U22175 (N_22175,N_21507,N_21124);
nor U22176 (N_22176,N_21610,N_21930);
xor U22177 (N_22177,N_21307,N_21890);
nor U22178 (N_22178,N_21259,N_21887);
and U22179 (N_22179,N_21624,N_21570);
xor U22180 (N_22180,N_21755,N_21869);
or U22181 (N_22181,N_21039,N_21420);
nand U22182 (N_22182,N_21514,N_21830);
nand U22183 (N_22183,N_21551,N_21428);
and U22184 (N_22184,N_21650,N_21597);
nand U22185 (N_22185,N_21078,N_21496);
nor U22186 (N_22186,N_21053,N_21088);
or U22187 (N_22187,N_21390,N_21616);
nand U22188 (N_22188,N_21217,N_21506);
and U22189 (N_22189,N_21089,N_21666);
xor U22190 (N_22190,N_21742,N_21343);
xnor U22191 (N_22191,N_21082,N_21993);
xor U22192 (N_22192,N_21470,N_21417);
xnor U22193 (N_22193,N_21865,N_21523);
xor U22194 (N_22194,N_21618,N_21995);
and U22195 (N_22195,N_21907,N_21696);
xor U22196 (N_22196,N_21775,N_21522);
and U22197 (N_22197,N_21679,N_21735);
nand U22198 (N_22198,N_21108,N_21722);
nor U22199 (N_22199,N_21498,N_21800);
nor U22200 (N_22200,N_21751,N_21494);
nand U22201 (N_22201,N_21315,N_21677);
and U22202 (N_22202,N_21831,N_21271);
and U22203 (N_22203,N_21699,N_21337);
and U22204 (N_22204,N_21174,N_21695);
nor U22205 (N_22205,N_21915,N_21859);
nor U22206 (N_22206,N_21158,N_21029);
nand U22207 (N_22207,N_21941,N_21959);
nand U22208 (N_22208,N_21464,N_21490);
nand U22209 (N_22209,N_21620,N_21789);
and U22210 (N_22210,N_21046,N_21267);
xor U22211 (N_22211,N_21000,N_21641);
xor U22212 (N_22212,N_21683,N_21648);
and U22213 (N_22213,N_21803,N_21975);
or U22214 (N_22214,N_21441,N_21346);
xnor U22215 (N_22215,N_21843,N_21510);
nor U22216 (N_22216,N_21565,N_21663);
nor U22217 (N_22217,N_21229,N_21626);
and U22218 (N_22218,N_21484,N_21811);
or U22219 (N_22219,N_21508,N_21923);
or U22220 (N_22220,N_21279,N_21685);
or U22221 (N_22221,N_21063,N_21566);
and U22222 (N_22222,N_21486,N_21989);
nand U22223 (N_22223,N_21639,N_21123);
nor U22224 (N_22224,N_21443,N_21525);
nand U22225 (N_22225,N_21012,N_21442);
and U22226 (N_22226,N_21265,N_21129);
nor U22227 (N_22227,N_21976,N_21536);
and U22228 (N_22228,N_21224,N_21127);
and U22229 (N_22229,N_21726,N_21528);
nand U22230 (N_22230,N_21543,N_21115);
or U22231 (N_22231,N_21644,N_21968);
and U22232 (N_22232,N_21003,N_21145);
xor U22233 (N_22233,N_21924,N_21230);
nand U22234 (N_22234,N_21750,N_21770);
nand U22235 (N_22235,N_21637,N_21526);
or U22236 (N_22236,N_21225,N_21050);
xnor U22237 (N_22237,N_21853,N_21847);
nand U22238 (N_22238,N_21816,N_21477);
or U22239 (N_22239,N_21356,N_21101);
or U22240 (N_22240,N_21248,N_21263);
xor U22241 (N_22241,N_21014,N_21734);
xnor U22242 (N_22242,N_21563,N_21943);
and U22243 (N_22243,N_21799,N_21165);
and U22244 (N_22244,N_21067,N_21061);
nor U22245 (N_22245,N_21444,N_21967);
and U22246 (N_22246,N_21808,N_21852);
nand U22247 (N_22247,N_21372,N_21202);
xor U22248 (N_22248,N_21768,N_21581);
or U22249 (N_22249,N_21667,N_21473);
or U22250 (N_22250,N_21904,N_21670);
xor U22251 (N_22251,N_21357,N_21892);
nor U22252 (N_22252,N_21901,N_21654);
nand U22253 (N_22253,N_21268,N_21146);
xnor U22254 (N_22254,N_21426,N_21434);
nand U22255 (N_22255,N_21668,N_21448);
nor U22256 (N_22256,N_21033,N_21373);
nand U22257 (N_22257,N_21187,N_21084);
nor U22258 (N_22258,N_21921,N_21349);
and U22259 (N_22259,N_21132,N_21835);
and U22260 (N_22260,N_21405,N_21879);
nand U22261 (N_22261,N_21868,N_21592);
and U22262 (N_22262,N_21041,N_21085);
and U22263 (N_22263,N_21845,N_21946);
nand U22264 (N_22264,N_21354,N_21180);
xor U22265 (N_22265,N_21857,N_21529);
nor U22266 (N_22266,N_21293,N_21087);
xor U22267 (N_22267,N_21260,N_21854);
or U22268 (N_22268,N_21207,N_21355);
or U22269 (N_22269,N_21287,N_21094);
or U22270 (N_22270,N_21567,N_21604);
or U22271 (N_22271,N_21837,N_21693);
nand U22272 (N_22272,N_21839,N_21900);
or U22273 (N_22273,N_21144,N_21336);
and U22274 (N_22274,N_21814,N_21250);
nand U22275 (N_22275,N_21184,N_21856);
and U22276 (N_22276,N_21851,N_21018);
xor U22277 (N_22277,N_21499,N_21430);
and U22278 (N_22278,N_21102,N_21421);
nor U22279 (N_22279,N_21825,N_21083);
and U22280 (N_22280,N_21243,N_21801);
and U22281 (N_22281,N_21812,N_21152);
and U22282 (N_22282,N_21777,N_21657);
or U22283 (N_22283,N_21590,N_21753);
and U22284 (N_22284,N_21173,N_21861);
or U22285 (N_22285,N_21797,N_21392);
or U22286 (N_22286,N_21191,N_21977);
xor U22287 (N_22287,N_21568,N_21163);
and U22288 (N_22288,N_21586,N_21575);
nor U22289 (N_22289,N_21192,N_21073);
nor U22290 (N_22290,N_21463,N_21024);
nand U22291 (N_22291,N_21516,N_21707);
xor U22292 (N_22292,N_21705,N_21840);
nor U22293 (N_22293,N_21493,N_21792);
and U22294 (N_22294,N_21710,N_21380);
or U22295 (N_22295,N_21471,N_21377);
nor U22296 (N_22296,N_21210,N_21961);
nand U22297 (N_22297,N_21790,N_21918);
nor U22298 (N_22298,N_21125,N_21402);
or U22299 (N_22299,N_21703,N_21802);
or U22300 (N_22300,N_21957,N_21204);
nand U22301 (N_22301,N_21393,N_21782);
nor U22302 (N_22302,N_21647,N_21149);
xor U22303 (N_22303,N_21017,N_21401);
xor U22304 (N_22304,N_21316,N_21625);
xor U22305 (N_22305,N_21564,N_21360);
and U22306 (N_22306,N_21064,N_21739);
xor U22307 (N_22307,N_21282,N_21117);
nor U22308 (N_22308,N_21640,N_21671);
xnor U22309 (N_22309,N_21979,N_21070);
and U22310 (N_22310,N_21951,N_21829);
nand U22311 (N_22311,N_21886,N_21786);
xor U22312 (N_22312,N_21497,N_21423);
nand U22313 (N_22313,N_21148,N_21322);
xnor U22314 (N_22314,N_21382,N_21457);
and U22315 (N_22315,N_21791,N_21828);
nor U22316 (N_22316,N_21509,N_21607);
and U22317 (N_22317,N_21340,N_21687);
or U22318 (N_22318,N_21237,N_21103);
xor U22319 (N_22319,N_21664,N_21366);
or U22320 (N_22320,N_21077,N_21159);
xnor U22321 (N_22321,N_21665,N_21245);
or U22322 (N_22322,N_21160,N_21219);
nor U22323 (N_22323,N_21702,N_21826);
xor U22324 (N_22324,N_21836,N_21819);
nor U22325 (N_22325,N_21433,N_21619);
xor U22326 (N_22326,N_21774,N_21986);
xnor U22327 (N_22327,N_21549,N_21232);
xnor U22328 (N_22328,N_21414,N_21531);
or U22329 (N_22329,N_21327,N_21138);
or U22330 (N_22330,N_21577,N_21038);
nand U22331 (N_22331,N_21503,N_21987);
or U22332 (N_22332,N_21168,N_21690);
or U22333 (N_22333,N_21701,N_21051);
or U22334 (N_22334,N_21447,N_21406);
nor U22335 (N_22335,N_21416,N_21945);
nor U22336 (N_22336,N_21593,N_21806);
or U22337 (N_22337,N_21674,N_21251);
nor U22338 (N_22338,N_21515,N_21984);
nor U22339 (N_22339,N_21688,N_21059);
or U22340 (N_22340,N_21461,N_21698);
xor U22341 (N_22341,N_21540,N_21296);
and U22342 (N_22342,N_21458,N_21418);
or U22343 (N_22343,N_21730,N_21227);
or U22344 (N_22344,N_21884,N_21375);
nor U22345 (N_22345,N_21071,N_21042);
nor U22346 (N_22346,N_21784,N_21025);
nand U22347 (N_22347,N_21485,N_21254);
nor U22348 (N_22348,N_21762,N_21035);
xor U22349 (N_22349,N_21919,N_21505);
xnor U22350 (N_22350,N_21476,N_21646);
or U22351 (N_22351,N_21249,N_21917);
and U22352 (N_22352,N_21324,N_21212);
and U22353 (N_22353,N_21188,N_21130);
nand U22354 (N_22354,N_21970,N_21662);
nor U22355 (N_22355,N_21594,N_21351);
xnor U22356 (N_22356,N_21001,N_21958);
xor U22357 (N_22357,N_21398,N_21222);
or U22358 (N_22358,N_21400,N_21891);
nor U22359 (N_22359,N_21009,N_21623);
or U22360 (N_22360,N_21181,N_21600);
and U22361 (N_22361,N_21023,N_21533);
nor U22362 (N_22362,N_21408,N_21738);
and U22363 (N_22363,N_21359,N_21311);
and U22364 (N_22364,N_21672,N_21266);
nor U22365 (N_22365,N_21234,N_21369);
nor U22366 (N_22366,N_21040,N_21660);
or U22367 (N_22367,N_21952,N_21820);
nor U22368 (N_22368,N_21500,N_21288);
nor U22369 (N_22369,N_21465,N_21155);
and U22370 (N_22370,N_21656,N_21902);
xnor U22371 (N_22371,N_21304,N_21584);
and U22372 (N_22372,N_21936,N_21394);
or U22373 (N_22373,N_21692,N_21633);
nor U22374 (N_22374,N_21862,N_21990);
nand U22375 (N_22375,N_21285,N_21535);
or U22376 (N_22376,N_21055,N_21513);
or U22377 (N_22377,N_21246,N_21363);
and U22378 (N_22378,N_21595,N_21554);
nand U22379 (N_22379,N_21226,N_21395);
or U22380 (N_22380,N_21462,N_21841);
and U22381 (N_22381,N_21299,N_21697);
nor U22382 (N_22382,N_21475,N_21086);
or U22383 (N_22383,N_21537,N_21431);
or U22384 (N_22384,N_21466,N_21326);
or U22385 (N_22385,N_21396,N_21338);
nand U22386 (N_22386,N_21763,N_21460);
xnor U22387 (N_22387,N_21713,N_21882);
xnor U22388 (N_22388,N_21632,N_21313);
and U22389 (N_22389,N_21538,N_21081);
xor U22390 (N_22390,N_21539,N_21183);
nand U22391 (N_22391,N_21178,N_21135);
nand U22392 (N_22392,N_21215,N_21370);
xnor U22393 (N_22393,N_21194,N_21300);
xor U22394 (N_22394,N_21939,N_21793);
nor U22395 (N_22395,N_21532,N_21903);
or U22396 (N_22396,N_21878,N_21947);
and U22397 (N_22397,N_21992,N_21008);
nand U22398 (N_22398,N_21749,N_21429);
or U22399 (N_22399,N_21435,N_21978);
or U22400 (N_22400,N_21353,N_21119);
and U22401 (N_22401,N_21048,N_21842);
xor U22402 (N_22402,N_21201,N_21112);
or U22403 (N_22403,N_21855,N_21153);
nand U22404 (N_22404,N_21362,N_21822);
nor U22405 (N_22405,N_21612,N_21582);
xnor U22406 (N_22406,N_21779,N_21520);
or U22407 (N_22407,N_21942,N_21319);
nor U22408 (N_22408,N_21823,N_21519);
xnor U22409 (N_22409,N_21167,N_21332);
nor U22410 (N_22410,N_21973,N_21240);
nor U22411 (N_22411,N_21455,N_21247);
nor U22412 (N_22412,N_21809,N_21718);
nor U22413 (N_22413,N_21765,N_21098);
or U22414 (N_22414,N_21909,N_21838);
and U22415 (N_22415,N_21478,N_21312);
nor U22416 (N_22416,N_21002,N_21196);
and U22417 (N_22417,N_21562,N_21511);
nand U22418 (N_22418,N_21317,N_21557);
and U22419 (N_22419,N_21236,N_21333);
nand U22420 (N_22420,N_21096,N_21306);
xor U22421 (N_22421,N_21269,N_21481);
nand U22422 (N_22422,N_21962,N_21439);
xor U22423 (N_22423,N_21161,N_21213);
or U22424 (N_22424,N_21047,N_21295);
xor U22425 (N_22425,N_21092,N_21079);
nand U22426 (N_22426,N_21893,N_21113);
nand U22427 (N_22427,N_21274,N_21728);
xor U22428 (N_22428,N_21932,N_21436);
and U22429 (N_22429,N_21352,N_21341);
and U22430 (N_22430,N_21895,N_21583);
nand U22431 (N_22431,N_21920,N_21631);
nor U22432 (N_22432,N_21810,N_21605);
or U22433 (N_22433,N_21216,N_21621);
nor U22434 (N_22434,N_21170,N_21591);
nor U22435 (N_22435,N_21615,N_21005);
or U22436 (N_22436,N_21065,N_21114);
and U22437 (N_22437,N_21099,N_21281);
nand U22438 (N_22438,N_21141,N_21091);
nand U22439 (N_22439,N_21691,N_21495);
and U22440 (N_22440,N_21076,N_21090);
nand U22441 (N_22441,N_21278,N_21106);
nor U22442 (N_22442,N_21171,N_21097);
nor U22443 (N_22443,N_21031,N_21449);
nand U22444 (N_22444,N_21361,N_21908);
and U22445 (N_22445,N_21714,N_21972);
xor U22446 (N_22446,N_21955,N_21757);
or U22447 (N_22447,N_21766,N_21754);
and U22448 (N_22448,N_21318,N_21389);
nand U22449 (N_22449,N_21617,N_21971);
xor U22450 (N_22450,N_21297,N_21622);
nor U22451 (N_22451,N_21501,N_21649);
nor U22452 (N_22452,N_21329,N_21176);
or U22453 (N_22453,N_21474,N_21062);
and U22454 (N_22454,N_21110,N_21010);
xor U22455 (N_22455,N_21576,N_21253);
nor U22456 (N_22456,N_21518,N_21037);
nand U22457 (N_22457,N_21717,N_21521);
nor U22458 (N_22458,N_21487,N_21645);
xnor U22459 (N_22459,N_21162,N_21534);
and U22460 (N_22460,N_21156,N_21653);
or U22461 (N_22461,N_21860,N_21468);
nor U22462 (N_22462,N_21422,N_21233);
and U22463 (N_22463,N_21143,N_21137);
nand U22464 (N_22464,N_21771,N_21933);
nand U22465 (N_22465,N_21479,N_21166);
nor U22466 (N_22466,N_21289,N_21587);
nand U22467 (N_22467,N_21636,N_21301);
and U22468 (N_22468,N_21214,N_21068);
nand U22469 (N_22469,N_21258,N_21383);
and U22470 (N_22470,N_21221,N_21172);
nand U22471 (N_22471,N_21556,N_21544);
nand U22472 (N_22472,N_21419,N_21303);
nand U22473 (N_22473,N_21404,N_21075);
nand U22474 (N_22474,N_21776,N_21966);
xnor U22475 (N_22475,N_21186,N_21203);
xnor U22476 (N_22476,N_21323,N_21938);
and U22477 (N_22477,N_21193,N_21613);
and U22478 (N_22478,N_21723,N_21410);
and U22479 (N_22479,N_21873,N_21910);
nand U22480 (N_22480,N_21052,N_21759);
nor U22481 (N_22481,N_21866,N_21412);
or U22482 (N_22482,N_21940,N_21680);
and U22483 (N_22483,N_21999,N_21552);
xor U22484 (N_22484,N_21678,N_21760);
nor U22485 (N_22485,N_21467,N_21182);
or U22486 (N_22486,N_21512,N_21150);
and U22487 (N_22487,N_21747,N_21761);
xnor U22488 (N_22488,N_21223,N_21733);
nor U22489 (N_22489,N_21139,N_21109);
nor U22490 (N_22490,N_21960,N_21284);
nor U22491 (N_22491,N_21834,N_21255);
nor U22492 (N_22492,N_21013,N_21937);
xor U22493 (N_22493,N_21104,N_21684);
nand U22494 (N_22494,N_21788,N_21681);
nor U22495 (N_22495,N_21658,N_21548);
or U22496 (N_22496,N_21635,N_21066);
nor U22497 (N_22497,N_21403,N_21286);
nand U22498 (N_22498,N_21030,N_21956);
xnor U22499 (N_22499,N_21399,N_21997);
and U22500 (N_22500,N_21356,N_21838);
or U22501 (N_22501,N_21561,N_21606);
nor U22502 (N_22502,N_21758,N_21823);
and U22503 (N_22503,N_21227,N_21530);
and U22504 (N_22504,N_21117,N_21071);
xnor U22505 (N_22505,N_21964,N_21209);
and U22506 (N_22506,N_21499,N_21432);
or U22507 (N_22507,N_21836,N_21326);
or U22508 (N_22508,N_21238,N_21251);
nor U22509 (N_22509,N_21546,N_21132);
nand U22510 (N_22510,N_21260,N_21444);
and U22511 (N_22511,N_21316,N_21171);
xor U22512 (N_22512,N_21431,N_21235);
nand U22513 (N_22513,N_21658,N_21065);
and U22514 (N_22514,N_21698,N_21658);
nor U22515 (N_22515,N_21216,N_21817);
and U22516 (N_22516,N_21208,N_21508);
nor U22517 (N_22517,N_21592,N_21919);
or U22518 (N_22518,N_21440,N_21167);
and U22519 (N_22519,N_21390,N_21386);
xor U22520 (N_22520,N_21907,N_21108);
nand U22521 (N_22521,N_21005,N_21555);
or U22522 (N_22522,N_21115,N_21569);
or U22523 (N_22523,N_21074,N_21374);
nor U22524 (N_22524,N_21110,N_21174);
or U22525 (N_22525,N_21335,N_21117);
xnor U22526 (N_22526,N_21206,N_21862);
and U22527 (N_22527,N_21307,N_21600);
nor U22528 (N_22528,N_21493,N_21426);
xor U22529 (N_22529,N_21614,N_21030);
or U22530 (N_22530,N_21883,N_21330);
or U22531 (N_22531,N_21158,N_21269);
nor U22532 (N_22532,N_21392,N_21399);
and U22533 (N_22533,N_21995,N_21699);
xnor U22534 (N_22534,N_21962,N_21648);
nand U22535 (N_22535,N_21141,N_21943);
and U22536 (N_22536,N_21989,N_21847);
or U22537 (N_22537,N_21236,N_21984);
or U22538 (N_22538,N_21668,N_21269);
nand U22539 (N_22539,N_21712,N_21738);
nor U22540 (N_22540,N_21783,N_21798);
nor U22541 (N_22541,N_21346,N_21726);
nand U22542 (N_22542,N_21493,N_21938);
or U22543 (N_22543,N_21329,N_21109);
or U22544 (N_22544,N_21175,N_21008);
or U22545 (N_22545,N_21760,N_21964);
or U22546 (N_22546,N_21939,N_21783);
nor U22547 (N_22547,N_21655,N_21230);
xnor U22548 (N_22548,N_21031,N_21222);
nor U22549 (N_22549,N_21936,N_21173);
nor U22550 (N_22550,N_21336,N_21739);
nand U22551 (N_22551,N_21913,N_21198);
nand U22552 (N_22552,N_21277,N_21494);
xnor U22553 (N_22553,N_21083,N_21654);
nor U22554 (N_22554,N_21748,N_21287);
xor U22555 (N_22555,N_21302,N_21727);
xnor U22556 (N_22556,N_21430,N_21768);
xor U22557 (N_22557,N_21768,N_21851);
xor U22558 (N_22558,N_21960,N_21177);
and U22559 (N_22559,N_21616,N_21636);
xor U22560 (N_22560,N_21817,N_21283);
nor U22561 (N_22561,N_21001,N_21564);
nand U22562 (N_22562,N_21022,N_21174);
xnor U22563 (N_22563,N_21813,N_21034);
xnor U22564 (N_22564,N_21980,N_21513);
nor U22565 (N_22565,N_21852,N_21941);
xnor U22566 (N_22566,N_21249,N_21823);
xnor U22567 (N_22567,N_21009,N_21539);
nand U22568 (N_22568,N_21791,N_21107);
and U22569 (N_22569,N_21701,N_21231);
or U22570 (N_22570,N_21936,N_21404);
or U22571 (N_22571,N_21081,N_21902);
and U22572 (N_22572,N_21051,N_21261);
nand U22573 (N_22573,N_21728,N_21030);
or U22574 (N_22574,N_21993,N_21622);
xor U22575 (N_22575,N_21445,N_21306);
xnor U22576 (N_22576,N_21612,N_21630);
xnor U22577 (N_22577,N_21931,N_21446);
or U22578 (N_22578,N_21218,N_21657);
xor U22579 (N_22579,N_21389,N_21586);
xor U22580 (N_22580,N_21313,N_21875);
or U22581 (N_22581,N_21708,N_21768);
or U22582 (N_22582,N_21429,N_21643);
or U22583 (N_22583,N_21452,N_21387);
nand U22584 (N_22584,N_21564,N_21812);
nand U22585 (N_22585,N_21538,N_21657);
and U22586 (N_22586,N_21897,N_21209);
nand U22587 (N_22587,N_21062,N_21875);
or U22588 (N_22588,N_21331,N_21975);
nand U22589 (N_22589,N_21353,N_21400);
and U22590 (N_22590,N_21487,N_21620);
nand U22591 (N_22591,N_21846,N_21360);
or U22592 (N_22592,N_21042,N_21084);
or U22593 (N_22593,N_21364,N_21077);
nand U22594 (N_22594,N_21203,N_21574);
xnor U22595 (N_22595,N_21256,N_21153);
and U22596 (N_22596,N_21416,N_21862);
xnor U22597 (N_22597,N_21519,N_21146);
nand U22598 (N_22598,N_21362,N_21986);
xor U22599 (N_22599,N_21136,N_21156);
or U22600 (N_22600,N_21188,N_21682);
or U22601 (N_22601,N_21678,N_21237);
xor U22602 (N_22602,N_21870,N_21170);
xnor U22603 (N_22603,N_21228,N_21718);
nand U22604 (N_22604,N_21130,N_21244);
nor U22605 (N_22605,N_21350,N_21367);
nand U22606 (N_22606,N_21090,N_21430);
xnor U22607 (N_22607,N_21209,N_21670);
or U22608 (N_22608,N_21378,N_21916);
or U22609 (N_22609,N_21477,N_21327);
or U22610 (N_22610,N_21413,N_21561);
xnor U22611 (N_22611,N_21335,N_21279);
or U22612 (N_22612,N_21465,N_21081);
xnor U22613 (N_22613,N_21163,N_21246);
nand U22614 (N_22614,N_21203,N_21589);
xnor U22615 (N_22615,N_21723,N_21146);
and U22616 (N_22616,N_21740,N_21581);
nor U22617 (N_22617,N_21702,N_21421);
nor U22618 (N_22618,N_21763,N_21244);
nor U22619 (N_22619,N_21281,N_21775);
or U22620 (N_22620,N_21055,N_21037);
and U22621 (N_22621,N_21266,N_21420);
and U22622 (N_22622,N_21355,N_21642);
nand U22623 (N_22623,N_21797,N_21953);
or U22624 (N_22624,N_21323,N_21646);
xnor U22625 (N_22625,N_21014,N_21919);
nand U22626 (N_22626,N_21264,N_21702);
nor U22627 (N_22627,N_21620,N_21781);
and U22628 (N_22628,N_21338,N_21949);
and U22629 (N_22629,N_21185,N_21789);
nand U22630 (N_22630,N_21296,N_21822);
and U22631 (N_22631,N_21325,N_21360);
nor U22632 (N_22632,N_21352,N_21858);
xor U22633 (N_22633,N_21782,N_21959);
or U22634 (N_22634,N_21346,N_21305);
nand U22635 (N_22635,N_21937,N_21675);
nand U22636 (N_22636,N_21492,N_21861);
nor U22637 (N_22637,N_21029,N_21336);
nand U22638 (N_22638,N_21104,N_21900);
and U22639 (N_22639,N_21235,N_21802);
nand U22640 (N_22640,N_21654,N_21520);
nor U22641 (N_22641,N_21280,N_21411);
nor U22642 (N_22642,N_21820,N_21887);
nor U22643 (N_22643,N_21799,N_21397);
xnor U22644 (N_22644,N_21278,N_21732);
nor U22645 (N_22645,N_21860,N_21331);
or U22646 (N_22646,N_21930,N_21950);
and U22647 (N_22647,N_21749,N_21075);
nand U22648 (N_22648,N_21579,N_21744);
and U22649 (N_22649,N_21571,N_21308);
or U22650 (N_22650,N_21820,N_21596);
xor U22651 (N_22651,N_21552,N_21638);
nand U22652 (N_22652,N_21638,N_21152);
nand U22653 (N_22653,N_21683,N_21930);
nand U22654 (N_22654,N_21307,N_21553);
and U22655 (N_22655,N_21434,N_21805);
and U22656 (N_22656,N_21236,N_21507);
nor U22657 (N_22657,N_21465,N_21901);
nor U22658 (N_22658,N_21894,N_21008);
nand U22659 (N_22659,N_21511,N_21196);
nor U22660 (N_22660,N_21072,N_21552);
xnor U22661 (N_22661,N_21641,N_21252);
nor U22662 (N_22662,N_21246,N_21336);
nand U22663 (N_22663,N_21850,N_21462);
nand U22664 (N_22664,N_21576,N_21821);
nor U22665 (N_22665,N_21148,N_21773);
nand U22666 (N_22666,N_21587,N_21334);
nand U22667 (N_22667,N_21322,N_21981);
or U22668 (N_22668,N_21407,N_21176);
and U22669 (N_22669,N_21464,N_21920);
nand U22670 (N_22670,N_21960,N_21463);
nand U22671 (N_22671,N_21339,N_21482);
nor U22672 (N_22672,N_21321,N_21708);
xor U22673 (N_22673,N_21153,N_21980);
and U22674 (N_22674,N_21128,N_21867);
and U22675 (N_22675,N_21962,N_21613);
and U22676 (N_22676,N_21626,N_21688);
and U22677 (N_22677,N_21214,N_21035);
nor U22678 (N_22678,N_21683,N_21611);
xor U22679 (N_22679,N_21541,N_21567);
xnor U22680 (N_22680,N_21853,N_21935);
or U22681 (N_22681,N_21214,N_21447);
and U22682 (N_22682,N_21678,N_21831);
xor U22683 (N_22683,N_21881,N_21593);
or U22684 (N_22684,N_21652,N_21218);
nor U22685 (N_22685,N_21210,N_21212);
or U22686 (N_22686,N_21274,N_21531);
xnor U22687 (N_22687,N_21400,N_21582);
or U22688 (N_22688,N_21463,N_21906);
nand U22689 (N_22689,N_21817,N_21592);
and U22690 (N_22690,N_21233,N_21369);
nor U22691 (N_22691,N_21666,N_21015);
xor U22692 (N_22692,N_21725,N_21860);
or U22693 (N_22693,N_21634,N_21747);
or U22694 (N_22694,N_21946,N_21639);
nor U22695 (N_22695,N_21289,N_21917);
and U22696 (N_22696,N_21593,N_21940);
nand U22697 (N_22697,N_21528,N_21305);
nor U22698 (N_22698,N_21674,N_21352);
xor U22699 (N_22699,N_21699,N_21762);
nand U22700 (N_22700,N_21521,N_21067);
nor U22701 (N_22701,N_21993,N_21240);
or U22702 (N_22702,N_21439,N_21444);
nand U22703 (N_22703,N_21285,N_21101);
or U22704 (N_22704,N_21029,N_21091);
xnor U22705 (N_22705,N_21442,N_21639);
or U22706 (N_22706,N_21160,N_21353);
and U22707 (N_22707,N_21992,N_21062);
nand U22708 (N_22708,N_21690,N_21643);
nor U22709 (N_22709,N_21515,N_21563);
and U22710 (N_22710,N_21368,N_21748);
nor U22711 (N_22711,N_21390,N_21146);
nand U22712 (N_22712,N_21026,N_21658);
nand U22713 (N_22713,N_21577,N_21065);
or U22714 (N_22714,N_21225,N_21309);
nor U22715 (N_22715,N_21633,N_21532);
xor U22716 (N_22716,N_21171,N_21366);
or U22717 (N_22717,N_21407,N_21788);
and U22718 (N_22718,N_21220,N_21032);
and U22719 (N_22719,N_21399,N_21855);
and U22720 (N_22720,N_21170,N_21751);
or U22721 (N_22721,N_21757,N_21434);
and U22722 (N_22722,N_21579,N_21076);
nor U22723 (N_22723,N_21317,N_21461);
or U22724 (N_22724,N_21388,N_21139);
nor U22725 (N_22725,N_21640,N_21133);
nand U22726 (N_22726,N_21776,N_21291);
xnor U22727 (N_22727,N_21637,N_21004);
or U22728 (N_22728,N_21979,N_21117);
xnor U22729 (N_22729,N_21631,N_21533);
and U22730 (N_22730,N_21809,N_21902);
nand U22731 (N_22731,N_21677,N_21803);
and U22732 (N_22732,N_21493,N_21199);
or U22733 (N_22733,N_21644,N_21352);
nor U22734 (N_22734,N_21397,N_21167);
nor U22735 (N_22735,N_21340,N_21520);
xnor U22736 (N_22736,N_21168,N_21610);
nor U22737 (N_22737,N_21419,N_21759);
nor U22738 (N_22738,N_21865,N_21471);
and U22739 (N_22739,N_21018,N_21940);
nand U22740 (N_22740,N_21257,N_21736);
nor U22741 (N_22741,N_21893,N_21258);
xnor U22742 (N_22742,N_21381,N_21275);
nor U22743 (N_22743,N_21419,N_21935);
nand U22744 (N_22744,N_21694,N_21916);
or U22745 (N_22745,N_21112,N_21948);
nor U22746 (N_22746,N_21388,N_21774);
and U22747 (N_22747,N_21712,N_21624);
and U22748 (N_22748,N_21366,N_21035);
xnor U22749 (N_22749,N_21404,N_21498);
and U22750 (N_22750,N_21907,N_21982);
xnor U22751 (N_22751,N_21141,N_21717);
nand U22752 (N_22752,N_21022,N_21561);
nor U22753 (N_22753,N_21885,N_21819);
and U22754 (N_22754,N_21754,N_21982);
nor U22755 (N_22755,N_21126,N_21566);
and U22756 (N_22756,N_21746,N_21791);
nor U22757 (N_22757,N_21094,N_21733);
and U22758 (N_22758,N_21577,N_21649);
nand U22759 (N_22759,N_21203,N_21210);
nor U22760 (N_22760,N_21059,N_21032);
and U22761 (N_22761,N_21614,N_21107);
and U22762 (N_22762,N_21244,N_21026);
and U22763 (N_22763,N_21288,N_21567);
or U22764 (N_22764,N_21774,N_21882);
or U22765 (N_22765,N_21624,N_21500);
nor U22766 (N_22766,N_21465,N_21572);
and U22767 (N_22767,N_21831,N_21886);
nand U22768 (N_22768,N_21800,N_21099);
xnor U22769 (N_22769,N_21053,N_21910);
and U22770 (N_22770,N_21079,N_21615);
nand U22771 (N_22771,N_21565,N_21629);
xor U22772 (N_22772,N_21788,N_21129);
or U22773 (N_22773,N_21658,N_21200);
xnor U22774 (N_22774,N_21842,N_21711);
nor U22775 (N_22775,N_21309,N_21076);
and U22776 (N_22776,N_21999,N_21969);
or U22777 (N_22777,N_21483,N_21670);
nor U22778 (N_22778,N_21908,N_21673);
nand U22779 (N_22779,N_21687,N_21668);
nand U22780 (N_22780,N_21979,N_21090);
nor U22781 (N_22781,N_21396,N_21908);
or U22782 (N_22782,N_21087,N_21954);
xor U22783 (N_22783,N_21625,N_21791);
nand U22784 (N_22784,N_21249,N_21505);
and U22785 (N_22785,N_21154,N_21191);
nor U22786 (N_22786,N_21489,N_21472);
xnor U22787 (N_22787,N_21362,N_21127);
and U22788 (N_22788,N_21719,N_21896);
nand U22789 (N_22789,N_21830,N_21999);
nor U22790 (N_22790,N_21050,N_21284);
nand U22791 (N_22791,N_21865,N_21952);
nand U22792 (N_22792,N_21705,N_21981);
and U22793 (N_22793,N_21946,N_21858);
nor U22794 (N_22794,N_21311,N_21143);
or U22795 (N_22795,N_21086,N_21255);
nor U22796 (N_22796,N_21371,N_21615);
nand U22797 (N_22797,N_21470,N_21213);
nor U22798 (N_22798,N_21654,N_21102);
and U22799 (N_22799,N_21688,N_21695);
xor U22800 (N_22800,N_21068,N_21384);
and U22801 (N_22801,N_21611,N_21753);
nor U22802 (N_22802,N_21334,N_21820);
or U22803 (N_22803,N_21868,N_21724);
nor U22804 (N_22804,N_21888,N_21381);
and U22805 (N_22805,N_21722,N_21074);
nand U22806 (N_22806,N_21130,N_21556);
and U22807 (N_22807,N_21880,N_21208);
xor U22808 (N_22808,N_21598,N_21295);
and U22809 (N_22809,N_21989,N_21544);
or U22810 (N_22810,N_21223,N_21142);
and U22811 (N_22811,N_21060,N_21948);
nor U22812 (N_22812,N_21234,N_21325);
xnor U22813 (N_22813,N_21947,N_21834);
xor U22814 (N_22814,N_21707,N_21560);
nand U22815 (N_22815,N_21065,N_21842);
nor U22816 (N_22816,N_21273,N_21211);
or U22817 (N_22817,N_21546,N_21594);
and U22818 (N_22818,N_21347,N_21698);
nand U22819 (N_22819,N_21777,N_21625);
and U22820 (N_22820,N_21070,N_21240);
xnor U22821 (N_22821,N_21390,N_21452);
nand U22822 (N_22822,N_21048,N_21145);
nand U22823 (N_22823,N_21372,N_21077);
nand U22824 (N_22824,N_21550,N_21796);
nor U22825 (N_22825,N_21108,N_21184);
xor U22826 (N_22826,N_21106,N_21840);
nand U22827 (N_22827,N_21660,N_21295);
or U22828 (N_22828,N_21576,N_21998);
or U22829 (N_22829,N_21516,N_21749);
or U22830 (N_22830,N_21905,N_21970);
nor U22831 (N_22831,N_21971,N_21116);
and U22832 (N_22832,N_21736,N_21926);
and U22833 (N_22833,N_21640,N_21507);
nand U22834 (N_22834,N_21856,N_21398);
and U22835 (N_22835,N_21396,N_21542);
nor U22836 (N_22836,N_21315,N_21634);
nand U22837 (N_22837,N_21871,N_21916);
nor U22838 (N_22838,N_21447,N_21767);
nand U22839 (N_22839,N_21408,N_21272);
nor U22840 (N_22840,N_21333,N_21946);
xor U22841 (N_22841,N_21614,N_21215);
nand U22842 (N_22842,N_21227,N_21053);
and U22843 (N_22843,N_21792,N_21447);
xor U22844 (N_22844,N_21051,N_21370);
nand U22845 (N_22845,N_21929,N_21243);
nor U22846 (N_22846,N_21349,N_21613);
or U22847 (N_22847,N_21311,N_21390);
and U22848 (N_22848,N_21252,N_21369);
nor U22849 (N_22849,N_21363,N_21020);
and U22850 (N_22850,N_21747,N_21438);
xnor U22851 (N_22851,N_21451,N_21399);
xnor U22852 (N_22852,N_21901,N_21614);
or U22853 (N_22853,N_21345,N_21307);
nand U22854 (N_22854,N_21404,N_21359);
xor U22855 (N_22855,N_21257,N_21907);
and U22856 (N_22856,N_21041,N_21956);
or U22857 (N_22857,N_21126,N_21567);
or U22858 (N_22858,N_21874,N_21992);
xor U22859 (N_22859,N_21265,N_21415);
nand U22860 (N_22860,N_21457,N_21726);
xnor U22861 (N_22861,N_21538,N_21000);
nor U22862 (N_22862,N_21068,N_21983);
nand U22863 (N_22863,N_21301,N_21308);
nand U22864 (N_22864,N_21111,N_21680);
or U22865 (N_22865,N_21196,N_21085);
xor U22866 (N_22866,N_21756,N_21784);
and U22867 (N_22867,N_21418,N_21663);
and U22868 (N_22868,N_21292,N_21006);
nor U22869 (N_22869,N_21921,N_21072);
xnor U22870 (N_22870,N_21757,N_21540);
and U22871 (N_22871,N_21225,N_21949);
nor U22872 (N_22872,N_21586,N_21157);
and U22873 (N_22873,N_21143,N_21970);
and U22874 (N_22874,N_21316,N_21646);
xor U22875 (N_22875,N_21705,N_21066);
and U22876 (N_22876,N_21959,N_21390);
and U22877 (N_22877,N_21240,N_21061);
nor U22878 (N_22878,N_21163,N_21493);
xor U22879 (N_22879,N_21140,N_21001);
or U22880 (N_22880,N_21523,N_21546);
or U22881 (N_22881,N_21199,N_21516);
nor U22882 (N_22882,N_21369,N_21188);
xor U22883 (N_22883,N_21334,N_21136);
nand U22884 (N_22884,N_21174,N_21915);
xnor U22885 (N_22885,N_21524,N_21404);
or U22886 (N_22886,N_21930,N_21516);
and U22887 (N_22887,N_21291,N_21833);
and U22888 (N_22888,N_21790,N_21239);
xnor U22889 (N_22889,N_21539,N_21394);
nand U22890 (N_22890,N_21847,N_21337);
xnor U22891 (N_22891,N_21011,N_21531);
or U22892 (N_22892,N_21607,N_21948);
or U22893 (N_22893,N_21994,N_21270);
nor U22894 (N_22894,N_21218,N_21658);
xor U22895 (N_22895,N_21895,N_21237);
nor U22896 (N_22896,N_21996,N_21959);
or U22897 (N_22897,N_21908,N_21676);
xnor U22898 (N_22898,N_21408,N_21976);
or U22899 (N_22899,N_21545,N_21201);
or U22900 (N_22900,N_21791,N_21614);
and U22901 (N_22901,N_21861,N_21731);
nor U22902 (N_22902,N_21319,N_21651);
and U22903 (N_22903,N_21117,N_21057);
nor U22904 (N_22904,N_21279,N_21372);
nand U22905 (N_22905,N_21444,N_21588);
or U22906 (N_22906,N_21334,N_21908);
and U22907 (N_22907,N_21477,N_21576);
nor U22908 (N_22908,N_21950,N_21749);
nor U22909 (N_22909,N_21181,N_21632);
xnor U22910 (N_22910,N_21687,N_21045);
nor U22911 (N_22911,N_21384,N_21113);
and U22912 (N_22912,N_21360,N_21664);
or U22913 (N_22913,N_21270,N_21620);
and U22914 (N_22914,N_21907,N_21003);
and U22915 (N_22915,N_21634,N_21531);
nor U22916 (N_22916,N_21317,N_21756);
xnor U22917 (N_22917,N_21854,N_21358);
nand U22918 (N_22918,N_21034,N_21719);
or U22919 (N_22919,N_21453,N_21421);
nand U22920 (N_22920,N_21758,N_21163);
nand U22921 (N_22921,N_21553,N_21394);
nor U22922 (N_22922,N_21037,N_21284);
nand U22923 (N_22923,N_21774,N_21694);
or U22924 (N_22924,N_21919,N_21499);
or U22925 (N_22925,N_21252,N_21287);
nand U22926 (N_22926,N_21408,N_21715);
xnor U22927 (N_22927,N_21507,N_21982);
xnor U22928 (N_22928,N_21624,N_21345);
xnor U22929 (N_22929,N_21900,N_21011);
nor U22930 (N_22930,N_21100,N_21252);
xor U22931 (N_22931,N_21739,N_21396);
nor U22932 (N_22932,N_21772,N_21161);
nor U22933 (N_22933,N_21732,N_21458);
xnor U22934 (N_22934,N_21813,N_21826);
or U22935 (N_22935,N_21713,N_21517);
nand U22936 (N_22936,N_21678,N_21935);
xnor U22937 (N_22937,N_21910,N_21555);
nor U22938 (N_22938,N_21065,N_21079);
nand U22939 (N_22939,N_21766,N_21402);
xor U22940 (N_22940,N_21836,N_21988);
or U22941 (N_22941,N_21180,N_21912);
nor U22942 (N_22942,N_21969,N_21072);
xnor U22943 (N_22943,N_21325,N_21308);
nor U22944 (N_22944,N_21381,N_21411);
nor U22945 (N_22945,N_21120,N_21581);
and U22946 (N_22946,N_21963,N_21688);
or U22947 (N_22947,N_21440,N_21646);
nor U22948 (N_22948,N_21361,N_21923);
nand U22949 (N_22949,N_21970,N_21491);
nand U22950 (N_22950,N_21848,N_21146);
nand U22951 (N_22951,N_21923,N_21240);
xor U22952 (N_22952,N_21778,N_21053);
nand U22953 (N_22953,N_21437,N_21223);
nor U22954 (N_22954,N_21291,N_21540);
and U22955 (N_22955,N_21110,N_21497);
nand U22956 (N_22956,N_21643,N_21729);
xor U22957 (N_22957,N_21391,N_21432);
xor U22958 (N_22958,N_21809,N_21771);
nand U22959 (N_22959,N_21934,N_21896);
nor U22960 (N_22960,N_21161,N_21112);
or U22961 (N_22961,N_21473,N_21023);
nand U22962 (N_22962,N_21148,N_21494);
nand U22963 (N_22963,N_21661,N_21276);
and U22964 (N_22964,N_21066,N_21883);
nor U22965 (N_22965,N_21818,N_21051);
nor U22966 (N_22966,N_21139,N_21081);
nand U22967 (N_22967,N_21219,N_21282);
and U22968 (N_22968,N_21731,N_21877);
or U22969 (N_22969,N_21457,N_21157);
and U22970 (N_22970,N_21525,N_21086);
and U22971 (N_22971,N_21907,N_21522);
nand U22972 (N_22972,N_21786,N_21995);
and U22973 (N_22973,N_21439,N_21043);
nand U22974 (N_22974,N_21126,N_21156);
nor U22975 (N_22975,N_21396,N_21645);
nand U22976 (N_22976,N_21758,N_21351);
nor U22977 (N_22977,N_21093,N_21183);
nor U22978 (N_22978,N_21573,N_21167);
or U22979 (N_22979,N_21314,N_21502);
nor U22980 (N_22980,N_21651,N_21907);
xnor U22981 (N_22981,N_21072,N_21449);
xor U22982 (N_22982,N_21806,N_21958);
xor U22983 (N_22983,N_21709,N_21884);
nand U22984 (N_22984,N_21183,N_21004);
and U22985 (N_22985,N_21814,N_21314);
nand U22986 (N_22986,N_21855,N_21779);
and U22987 (N_22987,N_21714,N_21512);
and U22988 (N_22988,N_21997,N_21915);
nand U22989 (N_22989,N_21434,N_21383);
nand U22990 (N_22990,N_21858,N_21030);
nand U22991 (N_22991,N_21317,N_21155);
or U22992 (N_22992,N_21899,N_21827);
nor U22993 (N_22993,N_21497,N_21217);
nand U22994 (N_22994,N_21763,N_21254);
or U22995 (N_22995,N_21511,N_21096);
and U22996 (N_22996,N_21908,N_21305);
xor U22997 (N_22997,N_21275,N_21043);
and U22998 (N_22998,N_21340,N_21436);
and U22999 (N_22999,N_21622,N_21170);
nand U23000 (N_23000,N_22917,N_22079);
xor U23001 (N_23001,N_22329,N_22179);
and U23002 (N_23002,N_22235,N_22066);
and U23003 (N_23003,N_22971,N_22171);
nor U23004 (N_23004,N_22626,N_22904);
or U23005 (N_23005,N_22906,N_22839);
xor U23006 (N_23006,N_22552,N_22475);
nand U23007 (N_23007,N_22806,N_22283);
and U23008 (N_23008,N_22916,N_22631);
or U23009 (N_23009,N_22429,N_22222);
nand U23010 (N_23010,N_22820,N_22989);
and U23011 (N_23011,N_22950,N_22697);
nor U23012 (N_23012,N_22870,N_22221);
nand U23013 (N_23013,N_22943,N_22751);
xnor U23014 (N_23014,N_22273,N_22008);
and U23015 (N_23015,N_22567,N_22117);
and U23016 (N_23016,N_22483,N_22979);
or U23017 (N_23017,N_22951,N_22776);
xnor U23018 (N_23018,N_22534,N_22188);
and U23019 (N_23019,N_22494,N_22175);
and U23020 (N_23020,N_22912,N_22669);
xor U23021 (N_23021,N_22443,N_22309);
nand U23022 (N_23022,N_22793,N_22985);
nor U23023 (N_23023,N_22553,N_22696);
xnor U23024 (N_23024,N_22208,N_22190);
nor U23025 (N_23025,N_22770,N_22430);
and U23026 (N_23026,N_22377,N_22275);
xor U23027 (N_23027,N_22047,N_22815);
xor U23028 (N_23028,N_22667,N_22423);
or U23029 (N_23029,N_22063,N_22603);
nand U23030 (N_23030,N_22942,N_22587);
xor U23031 (N_23031,N_22241,N_22525);
nor U23032 (N_23032,N_22217,N_22010);
nand U23033 (N_23033,N_22670,N_22480);
xor U23034 (N_23034,N_22037,N_22516);
nor U23035 (N_23035,N_22167,N_22386);
and U23036 (N_23036,N_22666,N_22141);
and U23037 (N_23037,N_22324,N_22156);
nand U23038 (N_23038,N_22163,N_22816);
and U23039 (N_23039,N_22784,N_22238);
and U23040 (N_23040,N_22144,N_22284);
or U23041 (N_23041,N_22592,N_22093);
nand U23042 (N_23042,N_22419,N_22286);
nand U23043 (N_23043,N_22433,N_22285);
nand U23044 (N_23044,N_22654,N_22691);
or U23045 (N_23045,N_22558,N_22456);
and U23046 (N_23046,N_22340,N_22426);
nor U23047 (N_23047,N_22395,N_22864);
or U23048 (N_23048,N_22024,N_22062);
or U23049 (N_23049,N_22360,N_22783);
xor U23050 (N_23050,N_22131,N_22116);
nand U23051 (N_23051,N_22227,N_22434);
nand U23052 (N_23052,N_22759,N_22688);
nand U23053 (N_23053,N_22245,N_22299);
or U23054 (N_23054,N_22956,N_22503);
nor U23055 (N_23055,N_22978,N_22708);
and U23056 (N_23056,N_22851,N_22214);
nor U23057 (N_23057,N_22780,N_22763);
nand U23058 (N_23058,N_22658,N_22936);
nor U23059 (N_23059,N_22575,N_22849);
xnor U23060 (N_23060,N_22888,N_22501);
xor U23061 (N_23061,N_22844,N_22479);
or U23062 (N_23062,N_22510,N_22898);
nor U23063 (N_23063,N_22316,N_22987);
nand U23064 (N_23064,N_22113,N_22502);
or U23065 (N_23065,N_22346,N_22665);
nor U23066 (N_23066,N_22098,N_22745);
nor U23067 (N_23067,N_22353,N_22524);
and U23068 (N_23068,N_22440,N_22327);
nor U23069 (N_23069,N_22647,N_22741);
and U23070 (N_23070,N_22859,N_22335);
nor U23071 (N_23071,N_22915,N_22519);
nand U23072 (N_23072,N_22084,N_22385);
nand U23073 (N_23073,N_22409,N_22656);
and U23074 (N_23074,N_22274,N_22952);
and U23075 (N_23075,N_22835,N_22879);
nand U23076 (N_23076,N_22657,N_22919);
and U23077 (N_23077,N_22493,N_22684);
or U23078 (N_23078,N_22344,N_22056);
and U23079 (N_23079,N_22400,N_22321);
or U23080 (N_23080,N_22536,N_22709);
or U23081 (N_23081,N_22143,N_22339);
xor U23082 (N_23082,N_22035,N_22837);
xnor U23083 (N_23083,N_22925,N_22805);
and U23084 (N_23084,N_22584,N_22396);
nor U23085 (N_23085,N_22108,N_22933);
xnor U23086 (N_23086,N_22506,N_22091);
xor U23087 (N_23087,N_22498,N_22875);
and U23088 (N_23088,N_22249,N_22313);
xnor U23089 (N_23089,N_22075,N_22205);
xnor U23090 (N_23090,N_22633,N_22161);
and U23091 (N_23091,N_22251,N_22099);
nor U23092 (N_23092,N_22325,N_22187);
and U23093 (N_23093,N_22865,N_22823);
xor U23094 (N_23094,N_22458,N_22383);
nand U23095 (N_23095,N_22550,N_22361);
nand U23096 (N_23096,N_22638,N_22444);
and U23097 (N_23097,N_22761,N_22323);
or U23098 (N_23098,N_22659,N_22546);
nor U23099 (N_23099,N_22090,N_22949);
nand U23100 (N_23100,N_22371,N_22388);
or U23101 (N_23101,N_22632,N_22146);
or U23102 (N_23102,N_22862,N_22442);
nor U23103 (N_23103,N_22269,N_22932);
xnor U23104 (N_23104,N_22046,N_22723);
nor U23105 (N_23105,N_22198,N_22454);
or U23106 (N_23106,N_22508,N_22120);
nor U23107 (N_23107,N_22636,N_22449);
nor U23108 (N_23108,N_22045,N_22769);
or U23109 (N_23109,N_22651,N_22474);
and U23110 (N_23110,N_22927,N_22122);
and U23111 (N_23111,N_22964,N_22164);
and U23112 (N_23112,N_22529,N_22314);
and U23113 (N_23113,N_22678,N_22293);
xnor U23114 (N_23114,N_22643,N_22893);
xor U23115 (N_23115,N_22840,N_22679);
nand U23116 (N_23116,N_22850,N_22350);
nand U23117 (N_23117,N_22112,N_22760);
nor U23118 (N_23118,N_22995,N_22027);
nand U23119 (N_23119,N_22310,N_22562);
and U23120 (N_23120,N_22941,N_22559);
nand U23121 (N_23121,N_22206,N_22089);
and U23122 (N_23122,N_22954,N_22040);
nand U23123 (N_23123,N_22076,N_22485);
or U23124 (N_23124,N_22965,N_22347);
nand U23125 (N_23125,N_22739,N_22722);
or U23126 (N_23126,N_22903,N_22064);
xor U23127 (N_23127,N_22137,N_22422);
and U23128 (N_23128,N_22911,N_22184);
and U23129 (N_23129,N_22367,N_22311);
or U23130 (N_23130,N_22374,N_22702);
xor U23131 (N_23131,N_22348,N_22604);
xor U23132 (N_23132,N_22734,N_22100);
nor U23133 (N_23133,N_22980,N_22052);
and U23134 (N_23134,N_22757,N_22407);
nor U23135 (N_23135,N_22960,N_22042);
nor U23136 (N_23136,N_22154,N_22414);
and U23137 (N_23137,N_22565,N_22594);
nand U23138 (N_23138,N_22629,N_22050);
nor U23139 (N_23139,N_22012,N_22884);
nor U23140 (N_23140,N_22548,N_22982);
nand U23141 (N_23141,N_22504,N_22455);
or U23142 (N_23142,N_22652,N_22107);
and U23143 (N_23143,N_22031,N_22991);
or U23144 (N_23144,N_22261,N_22464);
xor U23145 (N_23145,N_22677,N_22788);
nand U23146 (N_23146,N_22142,N_22532);
and U23147 (N_23147,N_22615,N_22599);
or U23148 (N_23148,N_22526,N_22557);
xnor U23149 (N_23149,N_22445,N_22145);
nand U23150 (N_23150,N_22945,N_22219);
nand U23151 (N_23151,N_22814,N_22686);
nor U23152 (N_23152,N_22857,N_22459);
and U23153 (N_23153,N_22280,N_22488);
and U23154 (N_23154,N_22999,N_22004);
nor U23155 (N_23155,N_22590,N_22034);
xnor U23156 (N_23156,N_22572,N_22399);
nor U23157 (N_23157,N_22614,N_22799);
nand U23158 (N_23158,N_22025,N_22938);
nor U23159 (N_23159,N_22975,N_22185);
nor U23160 (N_23160,N_22586,N_22929);
xnor U23161 (N_23161,N_22319,N_22298);
and U23162 (N_23162,N_22264,N_22181);
nand U23163 (N_23163,N_22258,N_22650);
or U23164 (N_23164,N_22551,N_22817);
xnor U23165 (N_23165,N_22994,N_22133);
nor U23166 (N_23166,N_22556,N_22866);
nand U23167 (N_23167,N_22831,N_22055);
or U23168 (N_23168,N_22662,N_22176);
xnor U23169 (N_23169,N_22289,N_22372);
xor U23170 (N_23170,N_22417,N_22002);
nand U23171 (N_23171,N_22860,N_22051);
and U23172 (N_23172,N_22721,N_22822);
xor U23173 (N_23173,N_22356,N_22328);
nor U23174 (N_23174,N_22425,N_22856);
or U23175 (N_23175,N_22438,N_22140);
xor U23176 (N_23176,N_22109,N_22819);
nand U23177 (N_23177,N_22343,N_22946);
nor U23178 (N_23178,N_22082,N_22048);
or U23179 (N_23179,N_22973,N_22096);
nand U23180 (N_23180,N_22305,N_22021);
nand U23181 (N_23181,N_22779,N_22229);
and U23182 (N_23182,N_22880,N_22663);
nand U23183 (N_23183,N_22207,N_22922);
and U23184 (N_23184,N_22993,N_22097);
or U23185 (N_23185,N_22029,N_22829);
xnor U23186 (N_23186,N_22637,N_22341);
nand U23187 (N_23187,N_22451,N_22810);
or U23188 (N_23188,N_22078,N_22500);
xor U23189 (N_23189,N_22660,N_22265);
nand U23190 (N_23190,N_22130,N_22716);
nor U23191 (N_23191,N_22259,N_22996);
and U23192 (N_23192,N_22674,N_22931);
or U23193 (N_23193,N_22199,N_22103);
and U23194 (N_23194,N_22373,N_22162);
or U23195 (N_23195,N_22026,N_22706);
or U23196 (N_23196,N_22640,N_22364);
nor U23197 (N_23197,N_22191,N_22410);
nand U23198 (N_23198,N_22088,N_22135);
xnor U23199 (N_23199,N_22539,N_22635);
xnor U23200 (N_23200,N_22366,N_22907);
and U23201 (N_23201,N_22481,N_22520);
and U23202 (N_23202,N_22809,N_22153);
nor U23203 (N_23203,N_22899,N_22067);
nor U23204 (N_23204,N_22527,N_22201);
and U23205 (N_23205,N_22778,N_22606);
nand U23206 (N_23206,N_22731,N_22482);
xnor U23207 (N_23207,N_22699,N_22969);
and U23208 (N_23208,N_22254,N_22389);
nor U23209 (N_23209,N_22472,N_22782);
nor U23210 (N_23210,N_22391,N_22795);
nand U23211 (N_23211,N_22266,N_22873);
and U23212 (N_23212,N_22682,N_22974);
xnor U23213 (N_23213,N_22023,N_22457);
or U23214 (N_23214,N_22649,N_22297);
or U23215 (N_23215,N_22150,N_22095);
xnor U23216 (N_23216,N_22123,N_22641);
or U23217 (N_23217,N_22215,N_22607);
nor U23218 (N_23218,N_22852,N_22484);
xnor U23219 (N_23219,N_22009,N_22126);
or U23220 (N_23220,N_22984,N_22826);
or U23221 (N_23221,N_22178,N_22495);
nand U23222 (N_23222,N_22762,N_22883);
nor U23223 (N_23223,N_22111,N_22256);
xor U23224 (N_23224,N_22303,N_22735);
xor U23225 (N_23225,N_22593,N_22541);
xor U23226 (N_23226,N_22773,N_22489);
nor U23227 (N_23227,N_22448,N_22465);
xor U23228 (N_23228,N_22671,N_22128);
and U23229 (N_23229,N_22715,N_22896);
xor U23230 (N_23230,N_22777,N_22953);
nand U23231 (N_23231,N_22262,N_22807);
and U23232 (N_23232,N_22071,N_22247);
and U23233 (N_23233,N_22753,N_22825);
xor U23234 (N_23234,N_22402,N_22039);
and U23235 (N_23235,N_22194,N_22081);
or U23236 (N_23236,N_22939,N_22596);
nor U23237 (N_23237,N_22756,N_22959);
xnor U23238 (N_23238,N_22487,N_22882);
xor U23239 (N_23239,N_22804,N_22874);
nand U23240 (N_23240,N_22522,N_22446);
xnor U23241 (N_23241,N_22909,N_22664);
or U23242 (N_23242,N_22743,N_22710);
xor U23243 (N_23243,N_22591,N_22694);
nand U23244 (N_23244,N_22692,N_22384);
and U23245 (N_23245,N_22749,N_22058);
nand U23246 (N_23246,N_22910,N_22742);
xnor U23247 (N_23247,N_22848,N_22398);
or U23248 (N_23248,N_22174,N_22582);
nand U23249 (N_23249,N_22608,N_22014);
nand U23250 (N_23250,N_22846,N_22411);
xnor U23251 (N_23251,N_22585,N_22155);
and U23252 (N_23252,N_22152,N_22216);
nand U23253 (N_23253,N_22855,N_22533);
nand U23254 (N_23254,N_22292,N_22543);
nand U23255 (N_23255,N_22331,N_22424);
nor U23256 (N_23256,N_22701,N_22203);
nand U23257 (N_23257,N_22560,N_22774);
or U23258 (N_23258,N_22237,N_22041);
nand U23259 (N_23259,N_22166,N_22988);
nor U23260 (N_23260,N_22032,N_22690);
or U23261 (N_23261,N_22787,N_22797);
nand U23262 (N_23262,N_22106,N_22955);
and U23263 (N_23263,N_22513,N_22581);
and U23264 (N_23264,N_22499,N_22887);
or U23265 (N_23265,N_22278,N_22876);
nand U23266 (N_23266,N_22054,N_22255);
or U23267 (N_23267,N_22785,N_22792);
nand U23268 (N_23268,N_22461,N_22600);
or U23269 (N_23269,N_22228,N_22644);
nand U23270 (N_23270,N_22634,N_22765);
xnor U23271 (N_23271,N_22720,N_22653);
nor U23272 (N_23272,N_22713,N_22272);
and U23273 (N_23273,N_22281,N_22333);
or U23274 (N_23274,N_22905,N_22382);
nor U23275 (N_23275,N_22200,N_22867);
nor U23276 (N_23276,N_22732,N_22704);
and U23277 (N_23277,N_22589,N_22576);
xor U23278 (N_23278,N_22376,N_22030);
nor U23279 (N_23279,N_22204,N_22342);
nor U23280 (N_23280,N_22068,N_22291);
nand U23281 (N_23281,N_22623,N_22101);
or U23282 (N_23282,N_22436,N_22157);
nor U23283 (N_23283,N_22754,N_22295);
nor U23284 (N_23284,N_22966,N_22843);
xnor U23285 (N_23285,N_22028,N_22791);
nand U23286 (N_23286,N_22935,N_22698);
xor U23287 (N_23287,N_22061,N_22220);
and U23288 (N_23288,N_22033,N_22416);
or U23289 (N_23289,N_22147,N_22290);
or U23290 (N_23290,N_22452,N_22225);
and U23291 (N_23291,N_22365,N_22110);
or U23292 (N_23292,N_22940,N_22270);
and U23293 (N_23293,N_22515,N_22802);
nor U23294 (N_23294,N_22038,N_22612);
nand U23295 (N_23295,N_22944,N_22209);
nor U23296 (N_23296,N_22926,N_22013);
nor U23297 (N_23297,N_22744,N_22958);
nand U23298 (N_23298,N_22948,N_22714);
or U23299 (N_23299,N_22854,N_22233);
xnor U23300 (N_23300,N_22136,N_22467);
nor U23301 (N_23301,N_22397,N_22359);
nor U23302 (N_23302,N_22719,N_22183);
or U23303 (N_23303,N_22730,N_22177);
and U23304 (N_23304,N_22072,N_22517);
and U23305 (N_23305,N_22841,N_22937);
nand U23306 (N_23306,N_22655,N_22394);
and U23307 (N_23307,N_22967,N_22300);
or U23308 (N_23308,N_22404,N_22628);
or U23309 (N_23309,N_22053,N_22127);
xor U23310 (N_23310,N_22357,N_22583);
nand U23311 (N_23311,N_22900,N_22412);
xnor U23312 (N_23312,N_22405,N_22354);
xor U23313 (N_23313,N_22330,N_22748);
and U23314 (N_23314,N_22571,N_22363);
nor U23315 (N_23315,N_22923,N_22868);
xor U23316 (N_23316,N_22003,N_22712);
nand U23317 (N_23317,N_22320,N_22160);
xnor U23318 (N_23318,N_22977,N_22711);
nor U23319 (N_23319,N_22891,N_22798);
xor U23320 (N_23320,N_22470,N_22326);
nand U23321 (N_23321,N_22733,N_22523);
or U23322 (N_23322,N_22118,N_22134);
nand U23323 (N_23323,N_22312,N_22598);
nand U23324 (N_23324,N_22447,N_22332);
or U23325 (N_23325,N_22928,N_22378);
or U23326 (N_23326,N_22195,N_22192);
xnor U23327 (N_23327,N_22717,N_22561);
xnor U23328 (N_23328,N_22369,N_22390);
nor U23329 (N_23329,N_22695,N_22420);
and U23330 (N_23330,N_22758,N_22511);
nor U23331 (N_23331,N_22252,N_22775);
xnor U23332 (N_23332,N_22648,N_22125);
and U23333 (N_23333,N_22828,N_22387);
nand U23334 (N_23334,N_22639,N_22193);
nand U23335 (N_23335,N_22740,N_22007);
and U23336 (N_23336,N_22083,N_22355);
or U23337 (N_23337,N_22727,N_22535);
and U23338 (N_23338,N_22248,N_22036);
and U23339 (N_23339,N_22240,N_22681);
nor U23340 (N_23340,N_22976,N_22808);
and U23341 (N_23341,N_22920,N_22537);
and U23342 (N_23342,N_22250,N_22947);
xor U23343 (N_23343,N_22092,N_22158);
nor U23344 (N_23344,N_22213,N_22005);
nor U23345 (N_23345,N_22886,N_22796);
nor U23346 (N_23346,N_22646,N_22086);
xnor U23347 (N_23347,N_22022,N_22263);
nor U23348 (N_23348,N_22579,N_22403);
and U23349 (N_23349,N_22318,N_22415);
or U23350 (N_23350,N_22705,N_22491);
and U23351 (N_23351,N_22441,N_22771);
nand U23352 (N_23352,N_22000,N_22963);
xor U23353 (N_23353,N_22672,N_22102);
or U23354 (N_23354,N_22673,N_22268);
nand U23355 (N_23355,N_22838,N_22683);
nand U23356 (N_23356,N_22555,N_22957);
xor U23357 (N_23357,N_22435,N_22149);
xnor U23358 (N_23358,N_22577,N_22017);
or U23359 (N_23359,N_22317,N_22800);
nand U23360 (N_23360,N_22352,N_22921);
nand U23361 (N_23361,N_22642,N_22223);
or U23362 (N_23362,N_22276,N_22094);
nor U23363 (N_23363,N_22863,N_22685);
nor U23364 (N_23364,N_22902,N_22821);
nor U23365 (N_23365,N_22858,N_22728);
xnor U23366 (N_23366,N_22794,N_22124);
nand U23367 (N_23367,N_22138,N_22401);
or U23368 (N_23368,N_22738,N_22689);
xor U23369 (N_23369,N_22392,N_22468);
nor U23370 (N_23370,N_22197,N_22497);
nand U23371 (N_23371,N_22218,N_22080);
and U23372 (N_23372,N_22990,N_22148);
nor U23373 (N_23373,N_22306,N_22169);
xnor U23374 (N_23374,N_22507,N_22224);
and U23375 (N_23375,N_22119,N_22530);
and U23376 (N_23376,N_22512,N_22408);
and U23377 (N_23377,N_22847,N_22267);
nor U23378 (N_23378,N_22613,N_22358);
or U23379 (N_23379,N_22542,N_22609);
and U23380 (N_23380,N_22746,N_22381);
or U23381 (N_23381,N_22226,N_22842);
xor U23382 (N_23382,N_22832,N_22496);
nand U23383 (N_23383,N_22246,N_22833);
nor U23384 (N_23384,N_22845,N_22315);
nand U23385 (N_23385,N_22619,N_22294);
or U23386 (N_23386,N_22540,N_22244);
and U23387 (N_23387,N_22172,N_22492);
nand U23388 (N_23388,N_22563,N_22789);
nand U23389 (N_23389,N_22307,N_22878);
nand U23390 (N_23390,N_22752,N_22432);
nor U23391 (N_23391,N_22531,N_22627);
or U23392 (N_23392,N_22074,N_22308);
nor U23393 (N_23393,N_22869,N_22700);
xnor U23394 (N_23394,N_22620,N_22296);
nand U23395 (N_23395,N_22718,N_22580);
nand U23396 (N_23396,N_22380,N_22070);
xor U23397 (N_23397,N_22618,N_22564);
nand U23398 (N_23398,N_22057,N_22243);
xor U23399 (N_23399,N_22545,N_22375);
and U23400 (N_23400,N_22345,N_22755);
nor U23401 (N_23401,N_22073,N_22992);
or U23402 (N_23402,N_22790,N_22729);
nand U23403 (N_23403,N_22818,N_22894);
xor U23404 (N_23404,N_22231,N_22824);
nor U23405 (N_23405,N_22439,N_22334);
nand U23406 (N_23406,N_22211,N_22336);
and U23407 (N_23407,N_22132,N_22624);
nor U23408 (N_23408,N_22602,N_22277);
nor U23409 (N_23409,N_22597,N_22834);
nor U23410 (N_23410,N_22930,N_22578);
and U23411 (N_23411,N_22772,N_22983);
and U23412 (N_23412,N_22767,N_22180);
or U23413 (N_23413,N_22693,N_22006);
nand U23414 (N_23414,N_22707,N_22087);
and U23415 (N_23415,N_22528,N_22018);
or U23416 (N_23416,N_22737,N_22924);
nor U23417 (N_23417,N_22505,N_22114);
nand U23418 (N_23418,N_22463,N_22961);
nand U23419 (N_23419,N_22889,N_22020);
and U23420 (N_23420,N_22901,N_22370);
and U23421 (N_23421,N_22962,N_22170);
nand U23422 (N_23422,N_22768,N_22288);
nand U23423 (N_23423,N_22750,N_22338);
xnor U23424 (N_23424,N_22595,N_22431);
and U23425 (N_23425,N_22812,N_22913);
nand U23426 (N_23426,N_22060,N_22115);
or U23427 (N_23427,N_22478,N_22453);
nor U23428 (N_23428,N_22680,N_22630);
and U23429 (N_23429,N_22044,N_22853);
and U23430 (N_23430,N_22885,N_22813);
or U23431 (N_23431,N_22016,N_22895);
xor U23432 (N_23432,N_22049,N_22766);
nor U23433 (N_23433,N_22239,N_22043);
nor U23434 (N_23434,N_22803,N_22476);
xor U23435 (N_23435,N_22568,N_22668);
nand U23436 (N_23436,N_22968,N_22349);
nor U23437 (N_23437,N_22544,N_22986);
xnor U23438 (N_23438,N_22981,N_22890);
and U23439 (N_23439,N_22521,N_22617);
nand U23440 (N_23440,N_22362,N_22918);
or U23441 (N_23441,N_22625,N_22574);
or U23442 (N_23442,N_22892,N_22085);
nand U23443 (N_23443,N_22159,N_22605);
nor U23444 (N_23444,N_22260,N_22687);
nor U23445 (N_23445,N_22588,N_22724);
nor U23446 (N_23446,N_22418,N_22427);
xor U23447 (N_23447,N_22872,N_22151);
and U23448 (N_23448,N_22279,N_22379);
nor U23449 (N_23449,N_22703,N_22059);
nor U23450 (N_23450,N_22271,N_22322);
nor U23451 (N_23451,N_22351,N_22621);
xor U23452 (N_23452,N_22549,N_22182);
xor U23453 (N_23453,N_22764,N_22105);
nor U23454 (N_23454,N_22547,N_22747);
or U23455 (N_23455,N_22861,N_22236);
nor U23456 (N_23456,N_22566,N_22509);
and U23457 (N_23457,N_22473,N_22573);
or U23458 (N_23458,N_22077,N_22570);
and U23459 (N_23459,N_22477,N_22611);
or U23460 (N_23460,N_22877,N_22302);
and U23461 (N_23461,N_22428,N_22908);
xor U23462 (N_23462,N_22230,N_22301);
nor U23463 (N_23463,N_22786,N_22304);
and U23464 (N_23464,N_22337,N_22736);
and U23465 (N_23465,N_22486,N_22676);
nand U23466 (N_23466,N_22196,N_22393);
nor U23467 (N_23467,N_22368,N_22811);
or U23468 (N_23468,N_22569,N_22253);
xor U23469 (N_23469,N_22998,N_22514);
nor U23470 (N_23470,N_22001,N_22554);
xor U23471 (N_23471,N_22069,N_22616);
xor U23472 (N_23472,N_22421,N_22406);
nor U23473 (N_23473,N_22645,N_22019);
nand U23474 (N_23474,N_22830,N_22801);
xor U23475 (N_23475,N_22997,N_22469);
nand U23476 (N_23476,N_22972,N_22437);
nor U23477 (N_23477,N_22871,N_22011);
nor U23478 (N_23478,N_22518,N_22827);
nor U23479 (N_23479,N_22173,N_22490);
nor U23480 (N_23480,N_22610,N_22897);
nand U23481 (N_23481,N_22538,N_22168);
nor U23482 (N_23482,N_22675,N_22601);
or U23483 (N_23483,N_22726,N_22413);
nand U23484 (N_23484,N_22661,N_22212);
nand U23485 (N_23485,N_22460,N_22471);
and U23486 (N_23486,N_22104,N_22242);
nor U23487 (N_23487,N_22282,N_22934);
or U23488 (N_23488,N_22065,N_22202);
or U23489 (N_23489,N_22165,N_22970);
and U23490 (N_23490,N_22781,N_22287);
nor U23491 (N_23491,N_22466,N_22622);
and U23492 (N_23492,N_22914,N_22210);
nand U23493 (N_23493,N_22462,N_22186);
or U23494 (N_23494,N_22234,N_22257);
nand U23495 (N_23495,N_22121,N_22232);
nor U23496 (N_23496,N_22450,N_22881);
and U23497 (N_23497,N_22189,N_22129);
or U23498 (N_23498,N_22725,N_22836);
xnor U23499 (N_23499,N_22139,N_22015);
and U23500 (N_23500,N_22127,N_22924);
nor U23501 (N_23501,N_22417,N_22868);
nand U23502 (N_23502,N_22367,N_22658);
xnor U23503 (N_23503,N_22330,N_22432);
xor U23504 (N_23504,N_22004,N_22215);
and U23505 (N_23505,N_22764,N_22881);
or U23506 (N_23506,N_22993,N_22084);
or U23507 (N_23507,N_22161,N_22387);
nor U23508 (N_23508,N_22508,N_22043);
nor U23509 (N_23509,N_22805,N_22701);
or U23510 (N_23510,N_22449,N_22098);
nand U23511 (N_23511,N_22638,N_22107);
nand U23512 (N_23512,N_22171,N_22982);
and U23513 (N_23513,N_22377,N_22070);
xnor U23514 (N_23514,N_22320,N_22131);
xnor U23515 (N_23515,N_22538,N_22115);
xnor U23516 (N_23516,N_22107,N_22643);
xnor U23517 (N_23517,N_22173,N_22713);
nand U23518 (N_23518,N_22015,N_22041);
or U23519 (N_23519,N_22811,N_22967);
and U23520 (N_23520,N_22253,N_22839);
nand U23521 (N_23521,N_22491,N_22112);
nand U23522 (N_23522,N_22497,N_22776);
nor U23523 (N_23523,N_22173,N_22904);
xor U23524 (N_23524,N_22211,N_22539);
nor U23525 (N_23525,N_22255,N_22237);
nand U23526 (N_23526,N_22142,N_22779);
or U23527 (N_23527,N_22902,N_22663);
and U23528 (N_23528,N_22487,N_22379);
nor U23529 (N_23529,N_22521,N_22413);
nand U23530 (N_23530,N_22724,N_22214);
nand U23531 (N_23531,N_22345,N_22855);
xnor U23532 (N_23532,N_22533,N_22919);
nor U23533 (N_23533,N_22719,N_22963);
xor U23534 (N_23534,N_22066,N_22010);
xor U23535 (N_23535,N_22722,N_22478);
or U23536 (N_23536,N_22311,N_22737);
or U23537 (N_23537,N_22136,N_22250);
nand U23538 (N_23538,N_22560,N_22108);
nand U23539 (N_23539,N_22685,N_22731);
nor U23540 (N_23540,N_22909,N_22106);
nand U23541 (N_23541,N_22220,N_22980);
nand U23542 (N_23542,N_22988,N_22306);
nor U23543 (N_23543,N_22995,N_22956);
nor U23544 (N_23544,N_22024,N_22299);
or U23545 (N_23545,N_22662,N_22573);
and U23546 (N_23546,N_22158,N_22816);
and U23547 (N_23547,N_22220,N_22716);
and U23548 (N_23548,N_22735,N_22562);
or U23549 (N_23549,N_22139,N_22377);
xor U23550 (N_23550,N_22189,N_22283);
and U23551 (N_23551,N_22094,N_22452);
nor U23552 (N_23552,N_22604,N_22513);
xnor U23553 (N_23553,N_22833,N_22257);
and U23554 (N_23554,N_22771,N_22423);
nor U23555 (N_23555,N_22681,N_22361);
xnor U23556 (N_23556,N_22050,N_22525);
or U23557 (N_23557,N_22842,N_22719);
or U23558 (N_23558,N_22593,N_22576);
or U23559 (N_23559,N_22200,N_22520);
or U23560 (N_23560,N_22892,N_22380);
xnor U23561 (N_23561,N_22644,N_22356);
xnor U23562 (N_23562,N_22570,N_22880);
or U23563 (N_23563,N_22422,N_22233);
nor U23564 (N_23564,N_22701,N_22876);
xnor U23565 (N_23565,N_22629,N_22815);
and U23566 (N_23566,N_22267,N_22536);
nand U23567 (N_23567,N_22980,N_22640);
or U23568 (N_23568,N_22626,N_22725);
or U23569 (N_23569,N_22546,N_22818);
or U23570 (N_23570,N_22737,N_22879);
or U23571 (N_23571,N_22198,N_22097);
or U23572 (N_23572,N_22681,N_22504);
and U23573 (N_23573,N_22048,N_22002);
and U23574 (N_23574,N_22005,N_22956);
or U23575 (N_23575,N_22196,N_22628);
nand U23576 (N_23576,N_22216,N_22468);
xnor U23577 (N_23577,N_22708,N_22121);
nor U23578 (N_23578,N_22070,N_22433);
nand U23579 (N_23579,N_22218,N_22833);
and U23580 (N_23580,N_22459,N_22508);
nand U23581 (N_23581,N_22967,N_22243);
and U23582 (N_23582,N_22211,N_22072);
nor U23583 (N_23583,N_22425,N_22643);
and U23584 (N_23584,N_22839,N_22591);
nand U23585 (N_23585,N_22334,N_22981);
and U23586 (N_23586,N_22727,N_22074);
and U23587 (N_23587,N_22939,N_22392);
nor U23588 (N_23588,N_22680,N_22419);
or U23589 (N_23589,N_22225,N_22041);
nor U23590 (N_23590,N_22520,N_22105);
and U23591 (N_23591,N_22739,N_22222);
nor U23592 (N_23592,N_22673,N_22392);
or U23593 (N_23593,N_22625,N_22402);
and U23594 (N_23594,N_22429,N_22208);
or U23595 (N_23595,N_22052,N_22860);
or U23596 (N_23596,N_22624,N_22695);
nor U23597 (N_23597,N_22547,N_22651);
nor U23598 (N_23598,N_22290,N_22495);
xnor U23599 (N_23599,N_22011,N_22428);
xnor U23600 (N_23600,N_22636,N_22172);
nor U23601 (N_23601,N_22563,N_22139);
or U23602 (N_23602,N_22485,N_22494);
nor U23603 (N_23603,N_22749,N_22109);
and U23604 (N_23604,N_22637,N_22027);
and U23605 (N_23605,N_22348,N_22629);
or U23606 (N_23606,N_22442,N_22515);
and U23607 (N_23607,N_22316,N_22222);
nor U23608 (N_23608,N_22789,N_22336);
xor U23609 (N_23609,N_22560,N_22922);
nor U23610 (N_23610,N_22550,N_22254);
and U23611 (N_23611,N_22709,N_22356);
or U23612 (N_23612,N_22905,N_22766);
and U23613 (N_23613,N_22874,N_22374);
and U23614 (N_23614,N_22190,N_22155);
xnor U23615 (N_23615,N_22475,N_22691);
xnor U23616 (N_23616,N_22067,N_22341);
and U23617 (N_23617,N_22115,N_22931);
nand U23618 (N_23618,N_22597,N_22091);
nor U23619 (N_23619,N_22125,N_22381);
nand U23620 (N_23620,N_22276,N_22638);
nor U23621 (N_23621,N_22726,N_22422);
and U23622 (N_23622,N_22785,N_22178);
or U23623 (N_23623,N_22248,N_22839);
or U23624 (N_23624,N_22288,N_22717);
xor U23625 (N_23625,N_22149,N_22534);
nor U23626 (N_23626,N_22288,N_22747);
nor U23627 (N_23627,N_22639,N_22641);
nand U23628 (N_23628,N_22669,N_22709);
nand U23629 (N_23629,N_22447,N_22930);
and U23630 (N_23630,N_22090,N_22741);
or U23631 (N_23631,N_22871,N_22680);
and U23632 (N_23632,N_22764,N_22852);
nand U23633 (N_23633,N_22157,N_22474);
nor U23634 (N_23634,N_22025,N_22498);
nand U23635 (N_23635,N_22384,N_22584);
nand U23636 (N_23636,N_22777,N_22053);
xnor U23637 (N_23637,N_22023,N_22720);
and U23638 (N_23638,N_22188,N_22007);
or U23639 (N_23639,N_22462,N_22572);
and U23640 (N_23640,N_22627,N_22662);
or U23641 (N_23641,N_22535,N_22084);
and U23642 (N_23642,N_22659,N_22007);
nand U23643 (N_23643,N_22901,N_22286);
nand U23644 (N_23644,N_22061,N_22178);
xor U23645 (N_23645,N_22031,N_22084);
or U23646 (N_23646,N_22182,N_22880);
nand U23647 (N_23647,N_22237,N_22889);
nor U23648 (N_23648,N_22334,N_22252);
xor U23649 (N_23649,N_22438,N_22528);
nor U23650 (N_23650,N_22138,N_22147);
nor U23651 (N_23651,N_22287,N_22176);
or U23652 (N_23652,N_22600,N_22555);
and U23653 (N_23653,N_22452,N_22224);
xnor U23654 (N_23654,N_22849,N_22944);
nor U23655 (N_23655,N_22683,N_22291);
or U23656 (N_23656,N_22974,N_22168);
nor U23657 (N_23657,N_22147,N_22346);
or U23658 (N_23658,N_22988,N_22948);
or U23659 (N_23659,N_22720,N_22621);
nand U23660 (N_23660,N_22480,N_22836);
and U23661 (N_23661,N_22986,N_22817);
nor U23662 (N_23662,N_22595,N_22071);
or U23663 (N_23663,N_22353,N_22181);
and U23664 (N_23664,N_22473,N_22690);
or U23665 (N_23665,N_22191,N_22442);
nor U23666 (N_23666,N_22288,N_22648);
and U23667 (N_23667,N_22285,N_22691);
nor U23668 (N_23668,N_22273,N_22689);
nand U23669 (N_23669,N_22718,N_22115);
and U23670 (N_23670,N_22315,N_22240);
xor U23671 (N_23671,N_22306,N_22026);
nor U23672 (N_23672,N_22257,N_22538);
or U23673 (N_23673,N_22992,N_22828);
nand U23674 (N_23674,N_22961,N_22365);
or U23675 (N_23675,N_22674,N_22155);
xor U23676 (N_23676,N_22229,N_22667);
and U23677 (N_23677,N_22161,N_22510);
xnor U23678 (N_23678,N_22541,N_22761);
xor U23679 (N_23679,N_22447,N_22981);
or U23680 (N_23680,N_22724,N_22141);
or U23681 (N_23681,N_22914,N_22796);
and U23682 (N_23682,N_22827,N_22068);
and U23683 (N_23683,N_22073,N_22195);
or U23684 (N_23684,N_22677,N_22914);
xnor U23685 (N_23685,N_22978,N_22530);
nand U23686 (N_23686,N_22845,N_22587);
and U23687 (N_23687,N_22819,N_22142);
nand U23688 (N_23688,N_22358,N_22164);
nand U23689 (N_23689,N_22347,N_22764);
and U23690 (N_23690,N_22137,N_22980);
nand U23691 (N_23691,N_22624,N_22437);
nor U23692 (N_23692,N_22565,N_22190);
and U23693 (N_23693,N_22876,N_22854);
and U23694 (N_23694,N_22557,N_22307);
xnor U23695 (N_23695,N_22480,N_22744);
and U23696 (N_23696,N_22358,N_22968);
and U23697 (N_23697,N_22613,N_22566);
nor U23698 (N_23698,N_22566,N_22453);
nand U23699 (N_23699,N_22570,N_22922);
or U23700 (N_23700,N_22073,N_22346);
xnor U23701 (N_23701,N_22311,N_22179);
nor U23702 (N_23702,N_22107,N_22783);
or U23703 (N_23703,N_22512,N_22734);
and U23704 (N_23704,N_22361,N_22179);
nor U23705 (N_23705,N_22194,N_22264);
nor U23706 (N_23706,N_22990,N_22307);
or U23707 (N_23707,N_22322,N_22895);
xor U23708 (N_23708,N_22685,N_22418);
nand U23709 (N_23709,N_22887,N_22075);
or U23710 (N_23710,N_22356,N_22244);
and U23711 (N_23711,N_22391,N_22603);
xnor U23712 (N_23712,N_22127,N_22054);
xnor U23713 (N_23713,N_22765,N_22366);
nand U23714 (N_23714,N_22230,N_22744);
or U23715 (N_23715,N_22831,N_22584);
nand U23716 (N_23716,N_22618,N_22209);
and U23717 (N_23717,N_22659,N_22406);
xnor U23718 (N_23718,N_22191,N_22088);
nand U23719 (N_23719,N_22673,N_22980);
or U23720 (N_23720,N_22173,N_22666);
and U23721 (N_23721,N_22091,N_22971);
and U23722 (N_23722,N_22281,N_22197);
or U23723 (N_23723,N_22250,N_22429);
and U23724 (N_23724,N_22761,N_22380);
nand U23725 (N_23725,N_22318,N_22582);
xor U23726 (N_23726,N_22014,N_22065);
nor U23727 (N_23727,N_22450,N_22584);
nor U23728 (N_23728,N_22748,N_22446);
nor U23729 (N_23729,N_22416,N_22119);
or U23730 (N_23730,N_22859,N_22782);
nor U23731 (N_23731,N_22694,N_22702);
and U23732 (N_23732,N_22194,N_22492);
nor U23733 (N_23733,N_22796,N_22007);
nor U23734 (N_23734,N_22077,N_22735);
nor U23735 (N_23735,N_22832,N_22215);
or U23736 (N_23736,N_22503,N_22642);
nand U23737 (N_23737,N_22646,N_22346);
and U23738 (N_23738,N_22973,N_22203);
and U23739 (N_23739,N_22549,N_22238);
nand U23740 (N_23740,N_22687,N_22143);
nand U23741 (N_23741,N_22953,N_22442);
nand U23742 (N_23742,N_22589,N_22411);
nor U23743 (N_23743,N_22366,N_22324);
or U23744 (N_23744,N_22635,N_22575);
or U23745 (N_23745,N_22411,N_22148);
and U23746 (N_23746,N_22010,N_22408);
xor U23747 (N_23747,N_22311,N_22854);
xnor U23748 (N_23748,N_22875,N_22069);
and U23749 (N_23749,N_22959,N_22201);
or U23750 (N_23750,N_22680,N_22778);
xor U23751 (N_23751,N_22233,N_22680);
or U23752 (N_23752,N_22164,N_22980);
or U23753 (N_23753,N_22841,N_22512);
nand U23754 (N_23754,N_22301,N_22583);
or U23755 (N_23755,N_22831,N_22267);
nand U23756 (N_23756,N_22171,N_22248);
and U23757 (N_23757,N_22787,N_22633);
xor U23758 (N_23758,N_22987,N_22856);
nor U23759 (N_23759,N_22289,N_22574);
xnor U23760 (N_23760,N_22933,N_22193);
or U23761 (N_23761,N_22660,N_22180);
nor U23762 (N_23762,N_22235,N_22406);
xor U23763 (N_23763,N_22802,N_22916);
and U23764 (N_23764,N_22132,N_22041);
and U23765 (N_23765,N_22364,N_22418);
and U23766 (N_23766,N_22956,N_22212);
and U23767 (N_23767,N_22396,N_22450);
xnor U23768 (N_23768,N_22065,N_22618);
xnor U23769 (N_23769,N_22337,N_22466);
and U23770 (N_23770,N_22670,N_22820);
or U23771 (N_23771,N_22553,N_22704);
nand U23772 (N_23772,N_22747,N_22274);
or U23773 (N_23773,N_22075,N_22769);
nand U23774 (N_23774,N_22719,N_22422);
and U23775 (N_23775,N_22025,N_22671);
and U23776 (N_23776,N_22350,N_22077);
nand U23777 (N_23777,N_22401,N_22432);
or U23778 (N_23778,N_22714,N_22329);
xor U23779 (N_23779,N_22219,N_22350);
or U23780 (N_23780,N_22269,N_22398);
or U23781 (N_23781,N_22510,N_22756);
nand U23782 (N_23782,N_22566,N_22792);
and U23783 (N_23783,N_22119,N_22591);
and U23784 (N_23784,N_22923,N_22563);
xor U23785 (N_23785,N_22109,N_22172);
and U23786 (N_23786,N_22386,N_22445);
and U23787 (N_23787,N_22886,N_22389);
and U23788 (N_23788,N_22476,N_22447);
or U23789 (N_23789,N_22334,N_22403);
nor U23790 (N_23790,N_22279,N_22545);
and U23791 (N_23791,N_22812,N_22471);
nand U23792 (N_23792,N_22630,N_22475);
nor U23793 (N_23793,N_22061,N_22032);
nor U23794 (N_23794,N_22627,N_22796);
nor U23795 (N_23795,N_22584,N_22758);
or U23796 (N_23796,N_22938,N_22143);
xor U23797 (N_23797,N_22362,N_22521);
xor U23798 (N_23798,N_22803,N_22459);
or U23799 (N_23799,N_22417,N_22502);
xnor U23800 (N_23800,N_22377,N_22459);
and U23801 (N_23801,N_22996,N_22245);
nand U23802 (N_23802,N_22310,N_22432);
nand U23803 (N_23803,N_22638,N_22855);
xnor U23804 (N_23804,N_22832,N_22356);
or U23805 (N_23805,N_22166,N_22864);
nand U23806 (N_23806,N_22620,N_22556);
or U23807 (N_23807,N_22298,N_22269);
nor U23808 (N_23808,N_22857,N_22256);
or U23809 (N_23809,N_22566,N_22647);
xor U23810 (N_23810,N_22352,N_22861);
xor U23811 (N_23811,N_22813,N_22568);
nand U23812 (N_23812,N_22704,N_22184);
nand U23813 (N_23813,N_22230,N_22040);
nor U23814 (N_23814,N_22931,N_22989);
xor U23815 (N_23815,N_22229,N_22756);
and U23816 (N_23816,N_22272,N_22523);
nand U23817 (N_23817,N_22319,N_22890);
xor U23818 (N_23818,N_22324,N_22321);
nor U23819 (N_23819,N_22205,N_22208);
xnor U23820 (N_23820,N_22207,N_22186);
and U23821 (N_23821,N_22657,N_22766);
and U23822 (N_23822,N_22454,N_22228);
nor U23823 (N_23823,N_22366,N_22186);
or U23824 (N_23824,N_22886,N_22497);
xnor U23825 (N_23825,N_22223,N_22847);
or U23826 (N_23826,N_22584,N_22820);
and U23827 (N_23827,N_22062,N_22981);
and U23828 (N_23828,N_22613,N_22837);
and U23829 (N_23829,N_22358,N_22917);
nand U23830 (N_23830,N_22298,N_22944);
or U23831 (N_23831,N_22061,N_22014);
or U23832 (N_23832,N_22965,N_22387);
or U23833 (N_23833,N_22597,N_22728);
xnor U23834 (N_23834,N_22470,N_22044);
or U23835 (N_23835,N_22937,N_22688);
xor U23836 (N_23836,N_22257,N_22354);
xnor U23837 (N_23837,N_22798,N_22325);
or U23838 (N_23838,N_22138,N_22277);
or U23839 (N_23839,N_22036,N_22478);
nor U23840 (N_23840,N_22418,N_22833);
or U23841 (N_23841,N_22617,N_22507);
and U23842 (N_23842,N_22763,N_22925);
or U23843 (N_23843,N_22861,N_22382);
or U23844 (N_23844,N_22135,N_22242);
or U23845 (N_23845,N_22667,N_22179);
or U23846 (N_23846,N_22451,N_22872);
and U23847 (N_23847,N_22661,N_22072);
xnor U23848 (N_23848,N_22151,N_22767);
nand U23849 (N_23849,N_22728,N_22093);
xnor U23850 (N_23850,N_22652,N_22880);
nor U23851 (N_23851,N_22720,N_22684);
nand U23852 (N_23852,N_22573,N_22918);
xnor U23853 (N_23853,N_22624,N_22843);
nor U23854 (N_23854,N_22895,N_22335);
nor U23855 (N_23855,N_22828,N_22583);
or U23856 (N_23856,N_22129,N_22581);
or U23857 (N_23857,N_22515,N_22209);
and U23858 (N_23858,N_22454,N_22579);
nor U23859 (N_23859,N_22996,N_22887);
nand U23860 (N_23860,N_22868,N_22009);
and U23861 (N_23861,N_22305,N_22545);
nor U23862 (N_23862,N_22824,N_22878);
nand U23863 (N_23863,N_22326,N_22245);
nand U23864 (N_23864,N_22857,N_22618);
nor U23865 (N_23865,N_22776,N_22641);
or U23866 (N_23866,N_22381,N_22764);
and U23867 (N_23867,N_22098,N_22891);
xor U23868 (N_23868,N_22699,N_22318);
xnor U23869 (N_23869,N_22377,N_22367);
or U23870 (N_23870,N_22936,N_22052);
or U23871 (N_23871,N_22267,N_22293);
xor U23872 (N_23872,N_22497,N_22621);
xnor U23873 (N_23873,N_22663,N_22426);
xor U23874 (N_23874,N_22260,N_22288);
or U23875 (N_23875,N_22899,N_22139);
nor U23876 (N_23876,N_22869,N_22717);
and U23877 (N_23877,N_22067,N_22651);
nor U23878 (N_23878,N_22346,N_22100);
nand U23879 (N_23879,N_22401,N_22953);
or U23880 (N_23880,N_22794,N_22669);
and U23881 (N_23881,N_22315,N_22377);
nand U23882 (N_23882,N_22570,N_22915);
nand U23883 (N_23883,N_22425,N_22491);
xor U23884 (N_23884,N_22947,N_22375);
xor U23885 (N_23885,N_22848,N_22381);
and U23886 (N_23886,N_22703,N_22567);
or U23887 (N_23887,N_22929,N_22082);
nand U23888 (N_23888,N_22405,N_22237);
nor U23889 (N_23889,N_22518,N_22145);
xor U23890 (N_23890,N_22659,N_22367);
nand U23891 (N_23891,N_22499,N_22430);
or U23892 (N_23892,N_22990,N_22186);
xor U23893 (N_23893,N_22780,N_22857);
nor U23894 (N_23894,N_22725,N_22814);
xnor U23895 (N_23895,N_22140,N_22406);
or U23896 (N_23896,N_22913,N_22200);
nand U23897 (N_23897,N_22264,N_22614);
nor U23898 (N_23898,N_22629,N_22321);
xor U23899 (N_23899,N_22652,N_22606);
nand U23900 (N_23900,N_22369,N_22291);
nor U23901 (N_23901,N_22459,N_22859);
nor U23902 (N_23902,N_22876,N_22864);
or U23903 (N_23903,N_22436,N_22433);
or U23904 (N_23904,N_22644,N_22492);
xor U23905 (N_23905,N_22672,N_22662);
or U23906 (N_23906,N_22385,N_22468);
xnor U23907 (N_23907,N_22318,N_22761);
nand U23908 (N_23908,N_22734,N_22737);
nor U23909 (N_23909,N_22969,N_22707);
nand U23910 (N_23910,N_22032,N_22940);
or U23911 (N_23911,N_22293,N_22774);
or U23912 (N_23912,N_22694,N_22766);
and U23913 (N_23913,N_22755,N_22169);
xnor U23914 (N_23914,N_22843,N_22003);
or U23915 (N_23915,N_22240,N_22850);
nor U23916 (N_23916,N_22389,N_22093);
and U23917 (N_23917,N_22228,N_22586);
nor U23918 (N_23918,N_22117,N_22254);
and U23919 (N_23919,N_22731,N_22077);
or U23920 (N_23920,N_22924,N_22894);
and U23921 (N_23921,N_22802,N_22738);
or U23922 (N_23922,N_22787,N_22306);
nor U23923 (N_23923,N_22743,N_22367);
and U23924 (N_23924,N_22767,N_22025);
nand U23925 (N_23925,N_22234,N_22349);
and U23926 (N_23926,N_22033,N_22751);
and U23927 (N_23927,N_22021,N_22897);
or U23928 (N_23928,N_22569,N_22986);
or U23929 (N_23929,N_22696,N_22199);
nor U23930 (N_23930,N_22749,N_22793);
and U23931 (N_23931,N_22215,N_22881);
or U23932 (N_23932,N_22393,N_22928);
and U23933 (N_23933,N_22703,N_22287);
or U23934 (N_23934,N_22109,N_22313);
nand U23935 (N_23935,N_22648,N_22797);
xor U23936 (N_23936,N_22325,N_22692);
nor U23937 (N_23937,N_22090,N_22765);
nor U23938 (N_23938,N_22349,N_22073);
or U23939 (N_23939,N_22025,N_22121);
xnor U23940 (N_23940,N_22059,N_22050);
and U23941 (N_23941,N_22462,N_22182);
nand U23942 (N_23942,N_22720,N_22826);
nor U23943 (N_23943,N_22627,N_22706);
or U23944 (N_23944,N_22421,N_22198);
or U23945 (N_23945,N_22860,N_22594);
or U23946 (N_23946,N_22256,N_22657);
or U23947 (N_23947,N_22602,N_22333);
xor U23948 (N_23948,N_22537,N_22751);
xnor U23949 (N_23949,N_22189,N_22461);
nor U23950 (N_23950,N_22234,N_22351);
xnor U23951 (N_23951,N_22761,N_22243);
or U23952 (N_23952,N_22512,N_22349);
nand U23953 (N_23953,N_22299,N_22642);
xnor U23954 (N_23954,N_22099,N_22060);
and U23955 (N_23955,N_22086,N_22104);
or U23956 (N_23956,N_22545,N_22755);
or U23957 (N_23957,N_22725,N_22654);
nand U23958 (N_23958,N_22662,N_22847);
and U23959 (N_23959,N_22338,N_22822);
xnor U23960 (N_23960,N_22382,N_22213);
or U23961 (N_23961,N_22462,N_22768);
and U23962 (N_23962,N_22827,N_22215);
nand U23963 (N_23963,N_22289,N_22063);
xor U23964 (N_23964,N_22791,N_22475);
nor U23965 (N_23965,N_22942,N_22070);
and U23966 (N_23966,N_22149,N_22761);
nand U23967 (N_23967,N_22162,N_22376);
or U23968 (N_23968,N_22306,N_22005);
xor U23969 (N_23969,N_22225,N_22678);
nand U23970 (N_23970,N_22397,N_22676);
or U23971 (N_23971,N_22417,N_22184);
and U23972 (N_23972,N_22163,N_22817);
or U23973 (N_23973,N_22825,N_22624);
and U23974 (N_23974,N_22558,N_22819);
nand U23975 (N_23975,N_22552,N_22467);
or U23976 (N_23976,N_22662,N_22722);
or U23977 (N_23977,N_22705,N_22654);
and U23978 (N_23978,N_22665,N_22270);
nor U23979 (N_23979,N_22503,N_22119);
xor U23980 (N_23980,N_22054,N_22890);
nand U23981 (N_23981,N_22698,N_22541);
nor U23982 (N_23982,N_22452,N_22534);
nand U23983 (N_23983,N_22429,N_22865);
and U23984 (N_23984,N_22880,N_22897);
nand U23985 (N_23985,N_22400,N_22429);
nor U23986 (N_23986,N_22116,N_22870);
and U23987 (N_23987,N_22236,N_22136);
xor U23988 (N_23988,N_22831,N_22281);
and U23989 (N_23989,N_22474,N_22258);
or U23990 (N_23990,N_22776,N_22034);
nor U23991 (N_23991,N_22368,N_22882);
nand U23992 (N_23992,N_22065,N_22550);
xor U23993 (N_23993,N_22218,N_22303);
and U23994 (N_23994,N_22564,N_22906);
and U23995 (N_23995,N_22455,N_22770);
and U23996 (N_23996,N_22778,N_22906);
nor U23997 (N_23997,N_22200,N_22762);
nor U23998 (N_23998,N_22068,N_22752);
nor U23999 (N_23999,N_22100,N_22241);
xnor U24000 (N_24000,N_23066,N_23906);
and U24001 (N_24001,N_23028,N_23851);
nand U24002 (N_24002,N_23325,N_23804);
xnor U24003 (N_24003,N_23393,N_23562);
or U24004 (N_24004,N_23553,N_23782);
xor U24005 (N_24005,N_23526,N_23963);
or U24006 (N_24006,N_23874,N_23311);
or U24007 (N_24007,N_23012,N_23558);
and U24008 (N_24008,N_23069,N_23828);
and U24009 (N_24009,N_23456,N_23151);
xor U24010 (N_24010,N_23376,N_23822);
nor U24011 (N_24011,N_23612,N_23208);
or U24012 (N_24012,N_23459,N_23572);
nand U24013 (N_24013,N_23132,N_23330);
nand U24014 (N_24014,N_23267,N_23165);
nor U24015 (N_24015,N_23847,N_23682);
or U24016 (N_24016,N_23735,N_23549);
xnor U24017 (N_24017,N_23001,N_23273);
nand U24018 (N_24018,N_23889,N_23450);
nand U24019 (N_24019,N_23105,N_23808);
nand U24020 (N_24020,N_23952,N_23888);
or U24021 (N_24021,N_23202,N_23849);
or U24022 (N_24022,N_23248,N_23207);
nor U24023 (N_24023,N_23044,N_23719);
or U24024 (N_24024,N_23995,N_23865);
nor U24025 (N_24025,N_23726,N_23184);
nor U24026 (N_24026,N_23984,N_23446);
and U24027 (N_24027,N_23848,N_23884);
nand U24028 (N_24028,N_23877,N_23366);
or U24029 (N_24029,N_23518,N_23217);
nand U24030 (N_24030,N_23815,N_23029);
xor U24031 (N_24031,N_23644,N_23814);
nand U24032 (N_24032,N_23126,N_23466);
nand U24033 (N_24033,N_23098,N_23896);
nor U24034 (N_24034,N_23994,N_23654);
or U24035 (N_24035,N_23762,N_23320);
xnor U24036 (N_24036,N_23975,N_23234);
or U24037 (N_24037,N_23426,N_23103);
nand U24038 (N_24038,N_23667,N_23869);
nor U24039 (N_24039,N_23580,N_23809);
nor U24040 (N_24040,N_23844,N_23390);
nor U24041 (N_24041,N_23062,N_23628);
or U24042 (N_24042,N_23964,N_23065);
and U24043 (N_24043,N_23806,N_23635);
and U24044 (N_24044,N_23759,N_23693);
or U24045 (N_24045,N_23647,N_23858);
xor U24046 (N_24046,N_23510,N_23625);
or U24047 (N_24047,N_23435,N_23344);
nor U24048 (N_24048,N_23381,N_23528);
nor U24049 (N_24049,N_23919,N_23680);
nand U24050 (N_24050,N_23880,N_23597);
or U24051 (N_24051,N_23198,N_23465);
nand U24052 (N_24052,N_23798,N_23479);
nor U24053 (N_24053,N_23675,N_23214);
xor U24054 (N_24054,N_23700,N_23595);
and U24055 (N_24055,N_23041,N_23441);
nor U24056 (N_24056,N_23371,N_23986);
or U24057 (N_24057,N_23536,N_23057);
nor U24058 (N_24058,N_23111,N_23965);
nor U24059 (N_24059,N_23474,N_23616);
and U24060 (N_24060,N_23006,N_23548);
or U24061 (N_24061,N_23070,N_23818);
and U24062 (N_24062,N_23911,N_23302);
nor U24063 (N_24063,N_23710,N_23801);
and U24064 (N_24064,N_23331,N_23615);
xnor U24065 (N_24065,N_23568,N_23530);
or U24066 (N_24066,N_23347,N_23707);
nor U24067 (N_24067,N_23564,N_23251);
nand U24068 (N_24068,N_23443,N_23221);
and U24069 (N_24069,N_23715,N_23797);
or U24070 (N_24070,N_23477,N_23457);
xnor U24071 (N_24071,N_23133,N_23689);
nand U24072 (N_24072,N_23772,N_23928);
and U24073 (N_24073,N_23945,N_23183);
xnor U24074 (N_24074,N_23543,N_23698);
nor U24075 (N_24075,N_23600,N_23577);
nor U24076 (N_24076,N_23396,N_23739);
and U24077 (N_24077,N_23895,N_23876);
and U24078 (N_24078,N_23279,N_23054);
and U24079 (N_24079,N_23145,N_23898);
nand U24080 (N_24080,N_23736,N_23345);
or U24081 (N_24081,N_23607,N_23665);
nand U24082 (N_24082,N_23645,N_23020);
nor U24083 (N_24083,N_23867,N_23387);
and U24084 (N_24084,N_23051,N_23516);
or U24085 (N_24085,N_23500,N_23959);
or U24086 (N_24086,N_23451,N_23432);
xnor U24087 (N_24087,N_23398,N_23533);
and U24088 (N_24088,N_23829,N_23250);
or U24089 (N_24089,N_23610,N_23901);
xor U24090 (N_24090,N_23786,N_23493);
or U24091 (N_24091,N_23596,N_23282);
and U24092 (N_24092,N_23671,N_23196);
and U24093 (N_24093,N_23714,N_23497);
and U24094 (N_24094,N_23767,N_23777);
nand U24095 (N_24095,N_23143,N_23318);
xor U24096 (N_24096,N_23556,N_23378);
nand U24097 (N_24097,N_23269,N_23550);
xor U24098 (N_24098,N_23840,N_23966);
and U24099 (N_24099,N_23873,N_23990);
nand U24100 (N_24100,N_23447,N_23420);
nor U24101 (N_24101,N_23134,N_23476);
nor U24102 (N_24102,N_23584,N_23704);
nor U24103 (N_24103,N_23690,N_23899);
and U24104 (N_24104,N_23579,N_23983);
nor U24105 (N_24105,N_23440,N_23352);
and U24106 (N_24106,N_23604,N_23365);
nand U24107 (N_24107,N_23931,N_23399);
and U24108 (N_24108,N_23483,N_23316);
xor U24109 (N_24109,N_23425,N_23769);
nor U24110 (N_24110,N_23537,N_23571);
nand U24111 (N_24111,N_23047,N_23169);
nand U24112 (N_24112,N_23587,N_23846);
or U24113 (N_24113,N_23638,N_23758);
xnor U24114 (N_24114,N_23663,N_23108);
xor U24115 (N_24115,N_23172,N_23890);
nand U24116 (N_24116,N_23669,N_23512);
and U24117 (N_24117,N_23223,N_23744);
xor U24118 (N_24118,N_23032,N_23683);
nand U24119 (N_24119,N_23130,N_23583);
nand U24120 (N_24120,N_23127,N_23629);
or U24121 (N_24121,N_23545,N_23664);
nor U24122 (N_24122,N_23490,N_23712);
or U24123 (N_24123,N_23229,N_23329);
and U24124 (N_24124,N_23115,N_23787);
xor U24125 (N_24125,N_23862,N_23951);
nand U24126 (N_24126,N_23323,N_23010);
xnor U24127 (N_24127,N_23071,N_23845);
nand U24128 (N_24128,N_23831,N_23188);
nand U24129 (N_24129,N_23158,N_23546);
xnor U24130 (N_24130,N_23042,N_23552);
and U24131 (N_24131,N_23886,N_23651);
nor U24132 (N_24132,N_23695,N_23096);
xnor U24133 (N_24133,N_23921,N_23298);
or U24134 (N_24134,N_23296,N_23303);
nand U24135 (N_24135,N_23839,N_23072);
or U24136 (N_24136,N_23637,N_23007);
nor U24137 (N_24137,N_23531,N_23887);
and U24138 (N_24138,N_23283,N_23468);
xor U24139 (N_24139,N_23720,N_23464);
nand U24140 (N_24140,N_23023,N_23471);
nor U24141 (N_24141,N_23294,N_23780);
or U24142 (N_24142,N_23292,N_23394);
nor U24143 (N_24143,N_23227,N_23509);
or U24144 (N_24144,N_23308,N_23264);
xor U24145 (N_24145,N_23192,N_23403);
nand U24146 (N_24146,N_23110,N_23702);
and U24147 (N_24147,N_23993,N_23241);
and U24148 (N_24148,N_23025,N_23833);
nand U24149 (N_24149,N_23709,N_23412);
and U24150 (N_24150,N_23494,N_23971);
and U24151 (N_24151,N_23670,N_23148);
xor U24152 (N_24152,N_23073,N_23788);
and U24153 (N_24153,N_23703,N_23730);
xor U24154 (N_24154,N_23406,N_23045);
xnor U24155 (N_24155,N_23961,N_23355);
or U24156 (N_24156,N_23827,N_23137);
nor U24157 (N_24157,N_23035,N_23729);
xor U24158 (N_24158,N_23778,N_23245);
and U24159 (N_24159,N_23742,N_23409);
nor U24160 (N_24160,N_23688,N_23418);
nand U24161 (N_24161,N_23560,N_23244);
and U24162 (N_24162,N_23978,N_23757);
nand U24163 (N_24163,N_23713,N_23908);
xor U24164 (N_24164,N_23470,N_23799);
xor U24165 (N_24165,N_23519,N_23673);
nor U24166 (N_24166,N_23124,N_23834);
nand U24167 (N_24167,N_23350,N_23734);
nor U24168 (N_24168,N_23106,N_23046);
nand U24169 (N_24169,N_23307,N_23861);
nor U24170 (N_24170,N_23542,N_23222);
and U24171 (N_24171,N_23383,N_23014);
nor U24172 (N_24172,N_23754,N_23237);
nor U24173 (N_24173,N_23349,N_23236);
nand U24174 (N_24174,N_23495,N_23104);
and U24175 (N_24175,N_23375,N_23226);
or U24176 (N_24176,N_23745,N_23201);
and U24177 (N_24177,N_23946,N_23872);
nor U24178 (N_24178,N_23085,N_23036);
nor U24179 (N_24179,N_23751,N_23776);
nand U24180 (N_24180,N_23287,N_23860);
and U24181 (N_24181,N_23416,N_23179);
and U24182 (N_24182,N_23838,N_23415);
and U24183 (N_24183,N_23711,N_23753);
nor U24184 (N_24184,N_23074,N_23534);
or U24185 (N_24185,N_23231,N_23960);
xnor U24186 (N_24186,N_23684,N_23659);
and U24187 (N_24187,N_23974,N_23033);
or U24188 (N_24188,N_23826,N_23634);
and U24189 (N_24189,N_23436,N_23168);
nand U24190 (N_24190,N_23167,N_23400);
nand U24191 (N_24191,N_23121,N_23590);
or U24192 (N_24192,N_23166,N_23621);
xnor U24193 (N_24193,N_23706,N_23206);
or U24194 (N_24194,N_23322,N_23658);
xnor U24195 (N_24195,N_23181,N_23177);
xor U24196 (N_24196,N_23360,N_23334);
and U24197 (N_24197,N_23864,N_23339);
xor U24198 (N_24198,N_23902,N_23107);
nand U24199 (N_24199,N_23609,N_23136);
and U24200 (N_24200,N_23953,N_23968);
or U24201 (N_24201,N_23270,N_23541);
nand U24202 (N_24202,N_23927,N_23271);
or U24203 (N_24203,N_23100,N_23048);
nand U24204 (N_24204,N_23011,N_23170);
xnor U24205 (N_24205,N_23699,N_23980);
nand U24206 (N_24206,N_23795,N_23348);
nor U24207 (N_24207,N_23082,N_23727);
xnor U24208 (N_24208,N_23022,N_23280);
xor U24209 (N_24209,N_23925,N_23557);
xor U24210 (N_24210,N_23544,N_23337);
and U24211 (N_24211,N_23697,N_23923);
xnor U24212 (N_24212,N_23414,N_23487);
xnor U24213 (N_24213,N_23262,N_23314);
or U24214 (N_24214,N_23841,N_23402);
and U24215 (N_24215,N_23084,N_23146);
or U24216 (N_24216,N_23149,N_23305);
and U24217 (N_24217,N_23195,N_23508);
xnor U24218 (N_24218,N_23038,N_23737);
and U24219 (N_24219,N_23527,N_23892);
nand U24220 (N_24220,N_23775,N_23463);
nor U24221 (N_24221,N_23164,N_23934);
nor U24222 (N_24222,N_23328,N_23218);
or U24223 (N_24223,N_23407,N_23233);
and U24224 (N_24224,N_23653,N_23224);
and U24225 (N_24225,N_23336,N_23897);
and U24226 (N_24226,N_23306,N_23160);
nor U24227 (N_24227,N_23920,N_23173);
nor U24228 (N_24228,N_23948,N_23228);
xnor U24229 (N_24229,N_23354,N_23086);
nand U24230 (N_24230,N_23346,N_23362);
or U24231 (N_24231,N_23091,N_23353);
or U24232 (N_24232,N_23657,N_23943);
or U24233 (N_24233,N_23662,N_23434);
or U24234 (N_24234,N_23685,N_23599);
and U24235 (N_24235,N_23204,N_23554);
and U24236 (N_24236,N_23112,N_23586);
nor U24237 (N_24237,N_23504,N_23640);
nor U24238 (N_24238,N_23191,N_23099);
and U24239 (N_24239,N_23410,N_23589);
nand U24240 (N_24240,N_23243,N_23197);
or U24241 (N_24241,N_23981,N_23515);
and U24242 (N_24242,N_23220,N_23796);
nand U24243 (N_24243,N_23142,N_23750);
nand U24244 (N_24244,N_23593,N_23225);
and U24245 (N_24245,N_23812,N_23304);
and U24246 (N_24246,N_23211,N_23430);
nor U24247 (N_24247,N_23120,N_23836);
and U24248 (N_24248,N_23982,N_23524);
xnor U24249 (N_24249,N_23823,N_23574);
nor U24250 (N_24250,N_23652,N_23962);
and U24251 (N_24251,N_23448,N_23004);
and U24252 (N_24252,N_23239,N_23914);
xnor U24253 (N_24253,N_23924,N_23342);
and U24254 (N_24254,N_23760,N_23768);
nor U24255 (N_24255,N_23295,N_23521);
or U24256 (N_24256,N_23335,N_23947);
nand U24257 (N_24257,N_23404,N_23602);
xnor U24258 (N_24258,N_23681,N_23077);
and U24259 (N_24259,N_23940,N_23816);
nand U24260 (N_24260,N_23930,N_23361);
and U24261 (N_24261,N_23128,N_23857);
xnor U24262 (N_24262,N_23079,N_23255);
or U24263 (N_24263,N_23254,N_23891);
nand U24264 (N_24264,N_23547,N_23591);
and U24265 (N_24265,N_23868,N_23391);
or U24266 (N_24266,N_23900,N_23395);
nand U24267 (N_24267,N_23819,N_23087);
nand U24268 (N_24268,N_23655,N_23193);
nand U24269 (N_24269,N_23850,N_23722);
xor U24270 (N_24270,N_23357,N_23122);
xnor U24271 (N_24271,N_23053,N_23917);
xnor U24272 (N_24272,N_23405,N_23453);
nand U24273 (N_24273,N_23408,N_23388);
or U24274 (N_24274,N_23871,N_23427);
nor U24275 (N_24275,N_23219,N_23150);
nor U24276 (N_24276,N_23529,N_23257);
nand U24277 (N_24277,N_23429,N_23469);
xnor U24278 (N_24278,N_23461,N_23532);
nand U24279 (N_24279,N_23310,N_23364);
and U24280 (N_24280,N_23538,N_23437);
nand U24281 (N_24281,N_23419,N_23300);
and U24282 (N_24282,N_23489,N_23368);
nor U24283 (N_24283,N_23505,N_23094);
nor U24284 (N_24284,N_23771,N_23731);
or U24285 (N_24285,N_23958,N_23049);
xnor U24286 (N_24286,N_23370,N_23392);
xnor U24287 (N_24287,N_23648,N_23904);
nor U24288 (N_24288,N_23747,N_23830);
or U24289 (N_24289,N_23118,N_23213);
nor U24290 (N_24290,N_23268,N_23639);
or U24291 (N_24291,N_23905,N_23341);
nand U24292 (N_24292,N_23601,N_23043);
or U24293 (N_24293,N_23358,N_23472);
and U24294 (N_24294,N_23676,N_23356);
xor U24295 (N_24295,N_23761,N_23691);
and U24296 (N_24296,N_23422,N_23794);
nor U24297 (N_24297,N_23379,N_23999);
nand U24298 (N_24298,N_23878,N_23240);
or U24299 (N_24299,N_23256,N_23040);
xnor U24300 (N_24300,N_23588,N_23511);
nor U24301 (N_24301,N_23613,N_23611);
and U24302 (N_24302,N_23113,N_23467);
and U24303 (N_24303,N_23277,N_23642);
nor U24304 (N_24304,N_23929,N_23825);
nor U24305 (N_24305,N_23748,N_23752);
and U24306 (N_24306,N_23992,N_23774);
and U24307 (N_24307,N_23954,N_23926);
xnor U24308 (N_24308,N_23176,N_23116);
nand U24309 (N_24309,N_23632,N_23566);
nand U24310 (N_24310,N_23154,N_23125);
and U24311 (N_24311,N_23174,N_23253);
or U24312 (N_24312,N_23162,N_23017);
nand U24313 (N_24313,N_23977,N_23030);
and U24314 (N_24314,N_23175,N_23488);
or U24315 (N_24315,N_23083,N_23090);
nor U24316 (N_24316,N_23272,N_23484);
nand U24317 (N_24317,N_23031,N_23458);
nor U24318 (N_24318,N_23944,N_23517);
or U24319 (N_24319,N_23081,N_23016);
nor U24320 (N_24320,N_23369,N_23247);
or U24321 (N_24321,N_23097,N_23856);
and U24322 (N_24322,N_23837,N_23563);
nand U24323 (N_24323,N_23626,N_23442);
or U24324 (N_24324,N_23882,N_23144);
xnor U24325 (N_24325,N_23721,N_23514);
nor U24326 (N_24326,N_23058,N_23499);
xor U24327 (N_24327,N_23486,N_23382);
nor U24328 (N_24328,N_23766,N_23285);
nor U24329 (N_24329,N_23912,N_23485);
nand U24330 (N_24330,N_23991,N_23153);
xnor U24331 (N_24331,N_23506,N_23424);
and U24332 (N_24332,N_23672,N_23525);
or U24333 (N_24333,N_23582,N_23743);
and U24334 (N_24334,N_23377,N_23941);
xor U24335 (N_24335,N_23646,N_23749);
xor U24336 (N_24336,N_23520,N_23343);
and U24337 (N_24337,N_23385,N_23018);
nor U24338 (N_24338,N_23853,N_23988);
nor U24339 (N_24339,N_23363,N_23955);
and U24340 (N_24340,N_23449,N_23810);
nand U24341 (N_24341,N_23265,N_23199);
nand U24342 (N_24342,N_23324,N_23050);
xnor U24343 (N_24343,N_23679,N_23705);
nand U24344 (N_24344,N_23903,N_23608);
xor U24345 (N_24345,N_23970,N_23894);
xor U24346 (N_24346,N_23092,N_23428);
or U24347 (N_24347,N_23985,N_23078);
nor U24348 (N_24348,N_23821,N_23575);
or U24349 (N_24349,N_23026,N_23327);
and U24350 (N_24350,N_23694,N_23956);
xnor U24351 (N_24351,N_23843,N_23119);
nor U24352 (N_24352,N_23692,N_23592);
or U24353 (N_24353,N_23678,N_23246);
or U24354 (N_24354,N_23570,N_23718);
and U24355 (N_24355,N_23938,N_23002);
and U24356 (N_24356,N_23624,N_23275);
nand U24357 (N_24357,N_23101,N_23949);
nor U24358 (N_24358,N_23359,N_23171);
and U24359 (N_24359,N_23501,N_23156);
xnor U24360 (N_24360,N_23332,N_23622);
and U24361 (N_24361,N_23650,N_23024);
nor U24362 (N_24362,N_23910,N_23109);
nor U24363 (N_24363,N_23288,N_23242);
nand U24364 (N_24364,N_23061,N_23820);
nand U24365 (N_24365,N_23666,N_23475);
or U24366 (N_24366,N_23312,N_23135);
nand U24367 (N_24367,N_23454,N_23139);
nand U24368 (N_24368,N_23942,N_23005);
nor U24369 (N_24369,N_23384,N_23194);
nand U24370 (N_24370,N_23792,N_23067);
or U24371 (N_24371,N_23800,N_23000);
xnor U24372 (N_24372,N_23423,N_23123);
nand U24373 (N_24373,N_23832,N_23732);
nand U24374 (N_24374,N_23781,N_23617);
nor U24375 (N_24375,N_23452,N_23063);
nor U24376 (N_24376,N_23015,N_23835);
and U24377 (N_24377,N_23802,N_23870);
nand U24378 (N_24378,N_23631,N_23445);
and U24379 (N_24379,N_23034,N_23674);
and U24380 (N_24380,N_23998,N_23738);
or U24381 (N_24381,N_23301,N_23696);
and U24382 (N_24382,N_23481,N_23950);
xor U24383 (N_24383,N_23784,N_23997);
and U24384 (N_24384,N_23261,N_23351);
nor U24385 (N_24385,N_23129,N_23717);
or U24386 (N_24386,N_23907,N_23212);
nor U24387 (N_24387,N_23540,N_23284);
xnor U24388 (N_24388,N_23444,N_23817);
and U24389 (N_24389,N_23716,N_23996);
xnor U24390 (N_24390,N_23783,N_23186);
xnor U24391 (N_24391,N_23003,N_23523);
nor U24392 (N_24392,N_23421,N_23299);
xor U24393 (N_24393,N_23478,N_23064);
xnor U24394 (N_24394,N_23027,N_23462);
nor U24395 (N_24395,N_23076,N_23319);
nand U24396 (N_24396,N_23989,N_23633);
or U24397 (N_24397,N_23052,N_23913);
xnor U24398 (N_24398,N_23263,N_23668);
nand U24399 (N_24399,N_23230,N_23155);
and U24400 (N_24400,N_23138,N_23630);
xor U24401 (N_24401,N_23502,N_23503);
nor U24402 (N_24402,N_23259,N_23933);
nand U24403 (N_24403,N_23649,N_23496);
and U24404 (N_24404,N_23863,N_23763);
xor U24405 (N_24405,N_23431,N_23756);
xnor U24406 (N_24406,N_23535,N_23641);
nand U24407 (N_24407,N_23585,N_23551);
nor U24408 (N_24408,N_23102,N_23374);
and U24409 (N_24409,N_23367,N_23438);
or U24410 (N_24410,N_23576,N_23232);
xnor U24411 (N_24411,N_23513,N_23159);
nor U24412 (N_24412,N_23859,N_23764);
xor U24413 (N_24413,N_23972,N_23411);
xnor U24414 (N_24414,N_23918,N_23725);
nor U24415 (N_24415,N_23482,N_23187);
xnor U24416 (N_24416,N_23973,N_23340);
or U24417 (N_24417,N_23238,N_23937);
or U24418 (N_24418,N_23915,N_23555);
or U24419 (N_24419,N_23161,N_23687);
xor U24420 (N_24420,N_23728,N_23755);
and U24421 (N_24421,N_23297,N_23701);
nor U24422 (N_24422,N_23785,N_23627);
xnor U24423 (N_24423,N_23893,N_23203);
xnor U24424 (N_24424,N_23578,N_23807);
nor U24425 (N_24425,N_23854,N_23885);
and U24426 (N_24426,N_23498,N_23189);
nand U24427 (N_24427,N_23088,N_23075);
nor U24428 (N_24428,N_23656,N_23152);
nand U24429 (N_24429,N_23455,N_23724);
and U24430 (N_24430,N_23190,N_23559);
xor U24431 (N_24431,N_23258,N_23561);
nand U24432 (N_24432,N_23293,N_23290);
nor U24433 (N_24433,N_23274,N_23141);
and U24434 (N_24434,N_23317,N_23935);
and U24435 (N_24435,N_23235,N_23793);
or U24436 (N_24436,N_23740,N_23661);
xor U24437 (N_24437,N_23569,N_23773);
nor U24438 (N_24438,N_23039,N_23413);
nor U24439 (N_24439,N_23037,N_23492);
nor U24440 (N_24440,N_23200,N_23117);
and U24441 (N_24441,N_23338,N_23824);
xnor U24442 (N_24442,N_23842,N_23276);
or U24443 (N_24443,N_23916,N_23205);
nand U24444 (N_24444,N_23581,N_23278);
nand U24445 (N_24445,N_23185,N_23770);
xnor U24446 (N_24446,N_23068,N_23056);
or U24447 (N_24447,N_23723,N_23875);
xnor U24448 (N_24448,N_23987,N_23620);
nand U24449 (N_24449,N_23979,N_23879);
nor U24450 (N_24450,N_23686,N_23095);
nor U24451 (N_24451,N_23281,N_23636);
xnor U24452 (N_24452,N_23326,N_23803);
nor U24453 (N_24453,N_23008,N_23677);
xor U24454 (N_24454,N_23019,N_23321);
xnor U24455 (N_24455,N_23210,N_23417);
and U24456 (N_24456,N_23401,N_23114);
and U24457 (N_24457,N_23573,N_23507);
or U24458 (N_24458,N_23060,N_23178);
nor U24459 (N_24459,N_23813,N_23598);
and U24460 (N_24460,N_23055,N_23936);
xnor U24461 (N_24461,N_23614,N_23286);
nor U24462 (N_24462,N_23215,N_23791);
or U24463 (N_24463,N_23976,N_23618);
nor U24464 (N_24464,N_23539,N_23147);
xnor U24465 (N_24465,N_23089,N_23855);
nor U24466 (N_24466,N_23881,N_23252);
xor U24467 (N_24467,N_23140,N_23957);
or U24468 (N_24468,N_23059,N_23397);
nand U24469 (N_24469,N_23790,N_23805);
or U24470 (N_24470,N_23733,N_23373);
nand U24471 (N_24471,N_23741,N_23779);
and U24472 (N_24472,N_23309,N_23013);
nand U24473 (N_24473,N_23922,N_23266);
xnor U24474 (N_24474,N_23093,N_23883);
nor U24475 (N_24475,N_23932,N_23708);
and U24476 (N_24476,N_23386,N_23372);
and U24477 (N_24477,N_23643,N_23460);
or U24478 (N_24478,N_23811,N_23789);
nor U24479 (N_24479,N_23315,N_23605);
nand U24480 (N_24480,N_23249,N_23606);
or U24481 (N_24481,N_23289,N_23594);
or U24482 (N_24482,N_23209,N_23567);
and U24483 (N_24483,N_23565,N_23491);
or U24484 (N_24484,N_23021,N_23765);
nor U24485 (N_24485,N_23623,N_23433);
xnor U24486 (N_24486,N_23852,N_23216);
or U24487 (N_24487,N_23660,N_23291);
nor U24488 (N_24488,N_23909,N_23080);
nand U24489 (N_24489,N_23389,N_23619);
or U24490 (N_24490,N_23380,N_23969);
xor U24491 (N_24491,N_23009,N_23522);
nand U24492 (N_24492,N_23182,N_23131);
nor U24493 (N_24493,N_23439,N_23967);
or U24494 (N_24494,N_23473,N_23603);
and U24495 (N_24495,N_23180,N_23163);
and U24496 (N_24496,N_23260,N_23866);
and U24497 (N_24497,N_23333,N_23746);
or U24498 (N_24498,N_23313,N_23480);
nand U24499 (N_24499,N_23939,N_23157);
xnor U24500 (N_24500,N_23414,N_23590);
or U24501 (N_24501,N_23420,N_23917);
nor U24502 (N_24502,N_23192,N_23412);
nor U24503 (N_24503,N_23246,N_23504);
and U24504 (N_24504,N_23763,N_23794);
or U24505 (N_24505,N_23503,N_23216);
and U24506 (N_24506,N_23643,N_23583);
or U24507 (N_24507,N_23536,N_23100);
or U24508 (N_24508,N_23379,N_23554);
nor U24509 (N_24509,N_23271,N_23284);
nand U24510 (N_24510,N_23005,N_23411);
or U24511 (N_24511,N_23166,N_23827);
nor U24512 (N_24512,N_23381,N_23796);
nor U24513 (N_24513,N_23929,N_23150);
xor U24514 (N_24514,N_23335,N_23782);
and U24515 (N_24515,N_23332,N_23570);
nor U24516 (N_24516,N_23915,N_23095);
or U24517 (N_24517,N_23660,N_23511);
xnor U24518 (N_24518,N_23288,N_23812);
xnor U24519 (N_24519,N_23561,N_23962);
nand U24520 (N_24520,N_23557,N_23159);
and U24521 (N_24521,N_23869,N_23538);
nor U24522 (N_24522,N_23886,N_23999);
and U24523 (N_24523,N_23623,N_23501);
nor U24524 (N_24524,N_23809,N_23860);
nand U24525 (N_24525,N_23137,N_23253);
and U24526 (N_24526,N_23205,N_23130);
nand U24527 (N_24527,N_23095,N_23877);
and U24528 (N_24528,N_23278,N_23292);
and U24529 (N_24529,N_23934,N_23897);
nor U24530 (N_24530,N_23483,N_23623);
xnor U24531 (N_24531,N_23984,N_23333);
nor U24532 (N_24532,N_23762,N_23978);
nor U24533 (N_24533,N_23682,N_23840);
nand U24534 (N_24534,N_23627,N_23747);
nor U24535 (N_24535,N_23055,N_23501);
xor U24536 (N_24536,N_23821,N_23740);
nor U24537 (N_24537,N_23629,N_23542);
nand U24538 (N_24538,N_23122,N_23910);
and U24539 (N_24539,N_23053,N_23582);
and U24540 (N_24540,N_23912,N_23795);
xnor U24541 (N_24541,N_23793,N_23126);
nor U24542 (N_24542,N_23781,N_23704);
and U24543 (N_24543,N_23041,N_23761);
nand U24544 (N_24544,N_23944,N_23347);
xnor U24545 (N_24545,N_23531,N_23724);
or U24546 (N_24546,N_23771,N_23065);
xnor U24547 (N_24547,N_23025,N_23323);
xnor U24548 (N_24548,N_23732,N_23659);
and U24549 (N_24549,N_23914,N_23455);
nor U24550 (N_24550,N_23928,N_23905);
and U24551 (N_24551,N_23198,N_23815);
nand U24552 (N_24552,N_23341,N_23552);
nor U24553 (N_24553,N_23299,N_23389);
and U24554 (N_24554,N_23057,N_23657);
or U24555 (N_24555,N_23866,N_23658);
nor U24556 (N_24556,N_23788,N_23220);
or U24557 (N_24557,N_23754,N_23227);
and U24558 (N_24558,N_23867,N_23308);
or U24559 (N_24559,N_23411,N_23598);
xnor U24560 (N_24560,N_23425,N_23191);
and U24561 (N_24561,N_23426,N_23130);
nor U24562 (N_24562,N_23723,N_23678);
xnor U24563 (N_24563,N_23178,N_23763);
or U24564 (N_24564,N_23374,N_23578);
or U24565 (N_24565,N_23756,N_23196);
or U24566 (N_24566,N_23856,N_23871);
or U24567 (N_24567,N_23878,N_23121);
xnor U24568 (N_24568,N_23440,N_23636);
or U24569 (N_24569,N_23640,N_23208);
or U24570 (N_24570,N_23500,N_23482);
or U24571 (N_24571,N_23381,N_23773);
or U24572 (N_24572,N_23367,N_23389);
or U24573 (N_24573,N_23607,N_23549);
and U24574 (N_24574,N_23523,N_23042);
nor U24575 (N_24575,N_23429,N_23872);
nand U24576 (N_24576,N_23926,N_23757);
or U24577 (N_24577,N_23056,N_23565);
nor U24578 (N_24578,N_23387,N_23328);
and U24579 (N_24579,N_23867,N_23638);
and U24580 (N_24580,N_23002,N_23129);
nand U24581 (N_24581,N_23734,N_23965);
and U24582 (N_24582,N_23223,N_23529);
or U24583 (N_24583,N_23486,N_23936);
xor U24584 (N_24584,N_23717,N_23454);
nor U24585 (N_24585,N_23204,N_23279);
or U24586 (N_24586,N_23587,N_23965);
or U24587 (N_24587,N_23269,N_23601);
xnor U24588 (N_24588,N_23914,N_23079);
nor U24589 (N_24589,N_23902,N_23021);
xor U24590 (N_24590,N_23182,N_23328);
or U24591 (N_24591,N_23931,N_23079);
xnor U24592 (N_24592,N_23864,N_23621);
nand U24593 (N_24593,N_23441,N_23833);
and U24594 (N_24594,N_23319,N_23103);
xnor U24595 (N_24595,N_23213,N_23355);
xor U24596 (N_24596,N_23095,N_23068);
nor U24597 (N_24597,N_23310,N_23767);
nand U24598 (N_24598,N_23773,N_23533);
or U24599 (N_24599,N_23858,N_23473);
xnor U24600 (N_24600,N_23844,N_23027);
nor U24601 (N_24601,N_23843,N_23116);
nor U24602 (N_24602,N_23519,N_23258);
nor U24603 (N_24603,N_23223,N_23820);
xnor U24604 (N_24604,N_23308,N_23219);
xnor U24605 (N_24605,N_23878,N_23744);
and U24606 (N_24606,N_23889,N_23457);
nand U24607 (N_24607,N_23348,N_23047);
and U24608 (N_24608,N_23690,N_23199);
nand U24609 (N_24609,N_23623,N_23218);
nand U24610 (N_24610,N_23817,N_23743);
xor U24611 (N_24611,N_23340,N_23061);
xnor U24612 (N_24612,N_23814,N_23483);
xor U24613 (N_24613,N_23370,N_23021);
and U24614 (N_24614,N_23192,N_23779);
or U24615 (N_24615,N_23627,N_23435);
xnor U24616 (N_24616,N_23088,N_23264);
nand U24617 (N_24617,N_23338,N_23654);
or U24618 (N_24618,N_23106,N_23066);
and U24619 (N_24619,N_23094,N_23768);
nor U24620 (N_24620,N_23199,N_23018);
and U24621 (N_24621,N_23803,N_23989);
and U24622 (N_24622,N_23354,N_23888);
nor U24623 (N_24623,N_23432,N_23153);
nor U24624 (N_24624,N_23794,N_23589);
and U24625 (N_24625,N_23362,N_23767);
nor U24626 (N_24626,N_23245,N_23145);
nand U24627 (N_24627,N_23909,N_23952);
xnor U24628 (N_24628,N_23890,N_23979);
and U24629 (N_24629,N_23054,N_23931);
and U24630 (N_24630,N_23820,N_23084);
nor U24631 (N_24631,N_23785,N_23447);
or U24632 (N_24632,N_23408,N_23560);
nand U24633 (N_24633,N_23740,N_23308);
nand U24634 (N_24634,N_23405,N_23455);
or U24635 (N_24635,N_23544,N_23847);
xor U24636 (N_24636,N_23640,N_23844);
and U24637 (N_24637,N_23268,N_23885);
nand U24638 (N_24638,N_23724,N_23454);
nor U24639 (N_24639,N_23170,N_23733);
nand U24640 (N_24640,N_23864,N_23387);
and U24641 (N_24641,N_23610,N_23739);
or U24642 (N_24642,N_23805,N_23195);
or U24643 (N_24643,N_23422,N_23548);
nor U24644 (N_24644,N_23219,N_23451);
nor U24645 (N_24645,N_23230,N_23658);
or U24646 (N_24646,N_23905,N_23768);
and U24647 (N_24647,N_23492,N_23204);
nor U24648 (N_24648,N_23139,N_23655);
nor U24649 (N_24649,N_23531,N_23403);
and U24650 (N_24650,N_23114,N_23157);
or U24651 (N_24651,N_23444,N_23795);
and U24652 (N_24652,N_23366,N_23932);
xnor U24653 (N_24653,N_23266,N_23421);
nor U24654 (N_24654,N_23620,N_23938);
xor U24655 (N_24655,N_23701,N_23840);
and U24656 (N_24656,N_23208,N_23770);
and U24657 (N_24657,N_23232,N_23205);
nor U24658 (N_24658,N_23880,N_23093);
and U24659 (N_24659,N_23412,N_23557);
xor U24660 (N_24660,N_23861,N_23059);
or U24661 (N_24661,N_23314,N_23498);
and U24662 (N_24662,N_23032,N_23965);
xor U24663 (N_24663,N_23045,N_23415);
xnor U24664 (N_24664,N_23716,N_23052);
and U24665 (N_24665,N_23912,N_23448);
and U24666 (N_24666,N_23325,N_23318);
or U24667 (N_24667,N_23275,N_23106);
and U24668 (N_24668,N_23883,N_23349);
and U24669 (N_24669,N_23930,N_23634);
nand U24670 (N_24670,N_23533,N_23264);
and U24671 (N_24671,N_23019,N_23096);
nor U24672 (N_24672,N_23922,N_23459);
nor U24673 (N_24673,N_23678,N_23150);
and U24674 (N_24674,N_23324,N_23586);
or U24675 (N_24675,N_23147,N_23376);
or U24676 (N_24676,N_23061,N_23830);
and U24677 (N_24677,N_23667,N_23122);
nor U24678 (N_24678,N_23553,N_23152);
nand U24679 (N_24679,N_23659,N_23252);
nand U24680 (N_24680,N_23056,N_23122);
xor U24681 (N_24681,N_23515,N_23499);
and U24682 (N_24682,N_23662,N_23067);
nor U24683 (N_24683,N_23344,N_23022);
nor U24684 (N_24684,N_23063,N_23620);
or U24685 (N_24685,N_23606,N_23388);
and U24686 (N_24686,N_23119,N_23852);
nor U24687 (N_24687,N_23932,N_23827);
xnor U24688 (N_24688,N_23947,N_23042);
and U24689 (N_24689,N_23169,N_23401);
and U24690 (N_24690,N_23212,N_23548);
nand U24691 (N_24691,N_23459,N_23399);
or U24692 (N_24692,N_23573,N_23784);
and U24693 (N_24693,N_23080,N_23081);
nand U24694 (N_24694,N_23231,N_23258);
nand U24695 (N_24695,N_23660,N_23004);
xnor U24696 (N_24696,N_23378,N_23544);
or U24697 (N_24697,N_23406,N_23921);
and U24698 (N_24698,N_23139,N_23147);
nor U24699 (N_24699,N_23921,N_23206);
and U24700 (N_24700,N_23196,N_23010);
and U24701 (N_24701,N_23684,N_23831);
or U24702 (N_24702,N_23915,N_23216);
and U24703 (N_24703,N_23870,N_23711);
or U24704 (N_24704,N_23039,N_23405);
or U24705 (N_24705,N_23934,N_23660);
xor U24706 (N_24706,N_23738,N_23804);
nor U24707 (N_24707,N_23556,N_23540);
and U24708 (N_24708,N_23077,N_23911);
and U24709 (N_24709,N_23629,N_23221);
xnor U24710 (N_24710,N_23008,N_23669);
and U24711 (N_24711,N_23360,N_23114);
nand U24712 (N_24712,N_23817,N_23372);
and U24713 (N_24713,N_23618,N_23603);
nor U24714 (N_24714,N_23284,N_23639);
nor U24715 (N_24715,N_23996,N_23267);
and U24716 (N_24716,N_23397,N_23234);
and U24717 (N_24717,N_23210,N_23401);
nor U24718 (N_24718,N_23010,N_23530);
xor U24719 (N_24719,N_23838,N_23356);
xor U24720 (N_24720,N_23658,N_23273);
xor U24721 (N_24721,N_23952,N_23785);
or U24722 (N_24722,N_23945,N_23457);
and U24723 (N_24723,N_23747,N_23515);
xnor U24724 (N_24724,N_23236,N_23428);
and U24725 (N_24725,N_23108,N_23435);
nand U24726 (N_24726,N_23608,N_23140);
and U24727 (N_24727,N_23658,N_23577);
nor U24728 (N_24728,N_23906,N_23152);
nor U24729 (N_24729,N_23938,N_23690);
and U24730 (N_24730,N_23984,N_23824);
and U24731 (N_24731,N_23142,N_23290);
or U24732 (N_24732,N_23455,N_23260);
and U24733 (N_24733,N_23356,N_23765);
and U24734 (N_24734,N_23003,N_23720);
xnor U24735 (N_24735,N_23059,N_23313);
nand U24736 (N_24736,N_23952,N_23111);
xnor U24737 (N_24737,N_23595,N_23443);
or U24738 (N_24738,N_23189,N_23726);
or U24739 (N_24739,N_23670,N_23242);
and U24740 (N_24740,N_23139,N_23278);
xor U24741 (N_24741,N_23827,N_23815);
nor U24742 (N_24742,N_23099,N_23592);
xor U24743 (N_24743,N_23619,N_23777);
or U24744 (N_24744,N_23187,N_23284);
and U24745 (N_24745,N_23056,N_23871);
xor U24746 (N_24746,N_23222,N_23398);
or U24747 (N_24747,N_23032,N_23625);
xnor U24748 (N_24748,N_23217,N_23769);
nand U24749 (N_24749,N_23847,N_23852);
nand U24750 (N_24750,N_23787,N_23895);
xor U24751 (N_24751,N_23364,N_23623);
and U24752 (N_24752,N_23307,N_23282);
or U24753 (N_24753,N_23018,N_23258);
xor U24754 (N_24754,N_23897,N_23649);
and U24755 (N_24755,N_23205,N_23002);
xnor U24756 (N_24756,N_23490,N_23630);
nand U24757 (N_24757,N_23969,N_23960);
nor U24758 (N_24758,N_23386,N_23815);
xor U24759 (N_24759,N_23201,N_23214);
nor U24760 (N_24760,N_23221,N_23771);
xor U24761 (N_24761,N_23791,N_23870);
and U24762 (N_24762,N_23995,N_23655);
xor U24763 (N_24763,N_23030,N_23568);
or U24764 (N_24764,N_23151,N_23479);
and U24765 (N_24765,N_23333,N_23684);
nor U24766 (N_24766,N_23690,N_23300);
or U24767 (N_24767,N_23585,N_23162);
xor U24768 (N_24768,N_23996,N_23395);
nor U24769 (N_24769,N_23079,N_23924);
xnor U24770 (N_24770,N_23505,N_23445);
nor U24771 (N_24771,N_23359,N_23063);
nand U24772 (N_24772,N_23620,N_23246);
nand U24773 (N_24773,N_23396,N_23067);
and U24774 (N_24774,N_23989,N_23284);
xor U24775 (N_24775,N_23956,N_23356);
nand U24776 (N_24776,N_23795,N_23662);
nand U24777 (N_24777,N_23440,N_23591);
xnor U24778 (N_24778,N_23099,N_23330);
nand U24779 (N_24779,N_23994,N_23316);
or U24780 (N_24780,N_23908,N_23857);
or U24781 (N_24781,N_23902,N_23729);
xnor U24782 (N_24782,N_23389,N_23518);
nor U24783 (N_24783,N_23633,N_23276);
xor U24784 (N_24784,N_23572,N_23121);
or U24785 (N_24785,N_23774,N_23855);
nand U24786 (N_24786,N_23302,N_23074);
nand U24787 (N_24787,N_23640,N_23380);
nand U24788 (N_24788,N_23796,N_23618);
and U24789 (N_24789,N_23773,N_23927);
nand U24790 (N_24790,N_23195,N_23207);
xnor U24791 (N_24791,N_23999,N_23097);
nor U24792 (N_24792,N_23947,N_23843);
xnor U24793 (N_24793,N_23621,N_23055);
nor U24794 (N_24794,N_23942,N_23887);
xnor U24795 (N_24795,N_23967,N_23407);
xnor U24796 (N_24796,N_23652,N_23255);
nor U24797 (N_24797,N_23786,N_23268);
nand U24798 (N_24798,N_23457,N_23350);
or U24799 (N_24799,N_23863,N_23128);
nand U24800 (N_24800,N_23788,N_23957);
and U24801 (N_24801,N_23029,N_23893);
and U24802 (N_24802,N_23530,N_23494);
or U24803 (N_24803,N_23726,N_23802);
or U24804 (N_24804,N_23992,N_23693);
or U24805 (N_24805,N_23290,N_23639);
and U24806 (N_24806,N_23320,N_23217);
nor U24807 (N_24807,N_23747,N_23287);
or U24808 (N_24808,N_23274,N_23113);
xor U24809 (N_24809,N_23920,N_23030);
and U24810 (N_24810,N_23484,N_23343);
or U24811 (N_24811,N_23819,N_23897);
and U24812 (N_24812,N_23552,N_23170);
or U24813 (N_24813,N_23025,N_23582);
nand U24814 (N_24814,N_23729,N_23504);
and U24815 (N_24815,N_23933,N_23247);
nand U24816 (N_24816,N_23913,N_23329);
and U24817 (N_24817,N_23223,N_23768);
and U24818 (N_24818,N_23216,N_23702);
xor U24819 (N_24819,N_23228,N_23190);
or U24820 (N_24820,N_23444,N_23899);
or U24821 (N_24821,N_23315,N_23695);
nor U24822 (N_24822,N_23171,N_23179);
nand U24823 (N_24823,N_23260,N_23229);
nor U24824 (N_24824,N_23589,N_23266);
nor U24825 (N_24825,N_23432,N_23075);
nand U24826 (N_24826,N_23556,N_23755);
or U24827 (N_24827,N_23848,N_23337);
nand U24828 (N_24828,N_23845,N_23172);
nand U24829 (N_24829,N_23092,N_23797);
nor U24830 (N_24830,N_23116,N_23633);
xor U24831 (N_24831,N_23245,N_23502);
or U24832 (N_24832,N_23980,N_23107);
xor U24833 (N_24833,N_23921,N_23201);
nor U24834 (N_24834,N_23261,N_23693);
or U24835 (N_24835,N_23581,N_23692);
or U24836 (N_24836,N_23736,N_23788);
or U24837 (N_24837,N_23256,N_23950);
xnor U24838 (N_24838,N_23616,N_23612);
and U24839 (N_24839,N_23502,N_23694);
nand U24840 (N_24840,N_23582,N_23992);
nand U24841 (N_24841,N_23487,N_23116);
xor U24842 (N_24842,N_23929,N_23831);
nand U24843 (N_24843,N_23002,N_23737);
or U24844 (N_24844,N_23944,N_23642);
xnor U24845 (N_24845,N_23267,N_23501);
xor U24846 (N_24846,N_23121,N_23481);
xnor U24847 (N_24847,N_23064,N_23132);
or U24848 (N_24848,N_23160,N_23077);
and U24849 (N_24849,N_23786,N_23924);
or U24850 (N_24850,N_23848,N_23462);
or U24851 (N_24851,N_23066,N_23922);
or U24852 (N_24852,N_23423,N_23136);
or U24853 (N_24853,N_23304,N_23234);
nor U24854 (N_24854,N_23661,N_23043);
xor U24855 (N_24855,N_23270,N_23585);
and U24856 (N_24856,N_23239,N_23242);
or U24857 (N_24857,N_23653,N_23832);
xnor U24858 (N_24858,N_23728,N_23889);
xor U24859 (N_24859,N_23496,N_23967);
and U24860 (N_24860,N_23323,N_23998);
nor U24861 (N_24861,N_23622,N_23133);
xor U24862 (N_24862,N_23216,N_23807);
nand U24863 (N_24863,N_23246,N_23964);
xnor U24864 (N_24864,N_23770,N_23545);
xnor U24865 (N_24865,N_23314,N_23082);
and U24866 (N_24866,N_23241,N_23453);
nor U24867 (N_24867,N_23784,N_23888);
xnor U24868 (N_24868,N_23558,N_23059);
xor U24869 (N_24869,N_23850,N_23047);
and U24870 (N_24870,N_23789,N_23093);
and U24871 (N_24871,N_23830,N_23010);
and U24872 (N_24872,N_23523,N_23598);
xor U24873 (N_24873,N_23999,N_23380);
and U24874 (N_24874,N_23046,N_23854);
or U24875 (N_24875,N_23784,N_23425);
and U24876 (N_24876,N_23525,N_23835);
nor U24877 (N_24877,N_23674,N_23914);
xnor U24878 (N_24878,N_23002,N_23356);
nor U24879 (N_24879,N_23158,N_23053);
xor U24880 (N_24880,N_23906,N_23122);
and U24881 (N_24881,N_23227,N_23930);
xnor U24882 (N_24882,N_23916,N_23060);
nor U24883 (N_24883,N_23242,N_23171);
nor U24884 (N_24884,N_23532,N_23629);
nand U24885 (N_24885,N_23996,N_23215);
nand U24886 (N_24886,N_23151,N_23640);
xnor U24887 (N_24887,N_23757,N_23114);
or U24888 (N_24888,N_23244,N_23460);
or U24889 (N_24889,N_23149,N_23770);
nand U24890 (N_24890,N_23500,N_23704);
nor U24891 (N_24891,N_23546,N_23384);
xor U24892 (N_24892,N_23795,N_23052);
nor U24893 (N_24893,N_23511,N_23991);
nand U24894 (N_24894,N_23783,N_23899);
nand U24895 (N_24895,N_23881,N_23706);
nor U24896 (N_24896,N_23481,N_23980);
or U24897 (N_24897,N_23920,N_23432);
and U24898 (N_24898,N_23347,N_23660);
nand U24899 (N_24899,N_23072,N_23175);
nor U24900 (N_24900,N_23756,N_23107);
nor U24901 (N_24901,N_23159,N_23283);
nor U24902 (N_24902,N_23172,N_23431);
nor U24903 (N_24903,N_23276,N_23525);
and U24904 (N_24904,N_23737,N_23444);
or U24905 (N_24905,N_23550,N_23666);
or U24906 (N_24906,N_23752,N_23387);
xor U24907 (N_24907,N_23621,N_23631);
xor U24908 (N_24908,N_23336,N_23937);
and U24909 (N_24909,N_23156,N_23831);
or U24910 (N_24910,N_23458,N_23202);
or U24911 (N_24911,N_23595,N_23546);
xor U24912 (N_24912,N_23042,N_23757);
or U24913 (N_24913,N_23513,N_23183);
and U24914 (N_24914,N_23368,N_23454);
or U24915 (N_24915,N_23603,N_23392);
and U24916 (N_24916,N_23822,N_23091);
or U24917 (N_24917,N_23960,N_23459);
or U24918 (N_24918,N_23427,N_23318);
xor U24919 (N_24919,N_23212,N_23350);
and U24920 (N_24920,N_23130,N_23868);
or U24921 (N_24921,N_23337,N_23140);
and U24922 (N_24922,N_23068,N_23579);
nor U24923 (N_24923,N_23056,N_23364);
nor U24924 (N_24924,N_23561,N_23139);
nor U24925 (N_24925,N_23666,N_23694);
nor U24926 (N_24926,N_23690,N_23375);
and U24927 (N_24927,N_23018,N_23379);
and U24928 (N_24928,N_23867,N_23385);
nand U24929 (N_24929,N_23319,N_23800);
or U24930 (N_24930,N_23671,N_23427);
nor U24931 (N_24931,N_23502,N_23306);
xnor U24932 (N_24932,N_23343,N_23726);
nor U24933 (N_24933,N_23764,N_23730);
nor U24934 (N_24934,N_23291,N_23918);
nor U24935 (N_24935,N_23170,N_23324);
nor U24936 (N_24936,N_23301,N_23258);
nor U24937 (N_24937,N_23335,N_23579);
and U24938 (N_24938,N_23329,N_23809);
nor U24939 (N_24939,N_23254,N_23257);
or U24940 (N_24940,N_23223,N_23832);
or U24941 (N_24941,N_23458,N_23521);
nor U24942 (N_24942,N_23604,N_23038);
nor U24943 (N_24943,N_23259,N_23276);
nor U24944 (N_24944,N_23910,N_23280);
xor U24945 (N_24945,N_23820,N_23770);
and U24946 (N_24946,N_23558,N_23068);
nor U24947 (N_24947,N_23947,N_23432);
or U24948 (N_24948,N_23581,N_23922);
xor U24949 (N_24949,N_23622,N_23560);
nand U24950 (N_24950,N_23347,N_23029);
or U24951 (N_24951,N_23847,N_23395);
and U24952 (N_24952,N_23617,N_23419);
xor U24953 (N_24953,N_23727,N_23331);
nand U24954 (N_24954,N_23530,N_23423);
nand U24955 (N_24955,N_23615,N_23324);
xnor U24956 (N_24956,N_23883,N_23936);
nor U24957 (N_24957,N_23449,N_23567);
nand U24958 (N_24958,N_23577,N_23092);
nor U24959 (N_24959,N_23684,N_23577);
nor U24960 (N_24960,N_23641,N_23943);
nand U24961 (N_24961,N_23766,N_23704);
nand U24962 (N_24962,N_23731,N_23512);
xor U24963 (N_24963,N_23418,N_23906);
nand U24964 (N_24964,N_23172,N_23604);
nor U24965 (N_24965,N_23790,N_23464);
or U24966 (N_24966,N_23403,N_23902);
and U24967 (N_24967,N_23789,N_23706);
nor U24968 (N_24968,N_23569,N_23291);
or U24969 (N_24969,N_23431,N_23072);
and U24970 (N_24970,N_23992,N_23129);
or U24971 (N_24971,N_23644,N_23226);
and U24972 (N_24972,N_23745,N_23799);
and U24973 (N_24973,N_23703,N_23449);
nand U24974 (N_24974,N_23889,N_23577);
or U24975 (N_24975,N_23225,N_23656);
nor U24976 (N_24976,N_23790,N_23456);
nor U24977 (N_24977,N_23292,N_23922);
nor U24978 (N_24978,N_23816,N_23710);
nand U24979 (N_24979,N_23485,N_23851);
xnor U24980 (N_24980,N_23459,N_23110);
or U24981 (N_24981,N_23212,N_23867);
or U24982 (N_24982,N_23811,N_23134);
nor U24983 (N_24983,N_23653,N_23105);
nor U24984 (N_24984,N_23432,N_23373);
or U24985 (N_24985,N_23741,N_23368);
and U24986 (N_24986,N_23573,N_23073);
xnor U24987 (N_24987,N_23546,N_23317);
and U24988 (N_24988,N_23302,N_23098);
xor U24989 (N_24989,N_23063,N_23180);
xnor U24990 (N_24990,N_23179,N_23046);
nor U24991 (N_24991,N_23544,N_23111);
or U24992 (N_24992,N_23906,N_23330);
and U24993 (N_24993,N_23801,N_23538);
xor U24994 (N_24994,N_23017,N_23054);
and U24995 (N_24995,N_23063,N_23374);
nor U24996 (N_24996,N_23581,N_23782);
xnor U24997 (N_24997,N_23451,N_23130);
and U24998 (N_24998,N_23388,N_23948);
or U24999 (N_24999,N_23093,N_23151);
nor U25000 (N_25000,N_24727,N_24324);
xor U25001 (N_25001,N_24182,N_24776);
or U25002 (N_25002,N_24077,N_24397);
nand U25003 (N_25003,N_24508,N_24961);
nor U25004 (N_25004,N_24822,N_24940);
nor U25005 (N_25005,N_24827,N_24695);
nand U25006 (N_25006,N_24749,N_24837);
nor U25007 (N_25007,N_24434,N_24932);
and U25008 (N_25008,N_24585,N_24645);
and U25009 (N_25009,N_24462,N_24995);
nand U25010 (N_25010,N_24240,N_24733);
nor U25011 (N_25011,N_24890,N_24163);
nor U25012 (N_25012,N_24422,N_24730);
xnor U25013 (N_25013,N_24797,N_24748);
and U25014 (N_25014,N_24832,N_24202);
and U25015 (N_25015,N_24994,N_24945);
nor U25016 (N_25016,N_24878,N_24907);
nand U25017 (N_25017,N_24988,N_24195);
nand U25018 (N_25018,N_24157,N_24257);
or U25019 (N_25019,N_24281,N_24102);
xnor U25020 (N_25020,N_24357,N_24551);
and U25021 (N_25021,N_24902,N_24633);
nor U25022 (N_25022,N_24449,N_24471);
and U25023 (N_25023,N_24252,N_24181);
or U25024 (N_25024,N_24796,N_24675);
or U25025 (N_25025,N_24828,N_24680);
nand U25026 (N_25026,N_24308,N_24008);
nor U25027 (N_25027,N_24885,N_24371);
and U25028 (N_25028,N_24817,N_24520);
or U25029 (N_25029,N_24975,N_24858);
or U25030 (N_25030,N_24128,N_24039);
nor U25031 (N_25031,N_24140,N_24139);
nor U25032 (N_25032,N_24459,N_24944);
nand U25033 (N_25033,N_24581,N_24844);
nand U25034 (N_25034,N_24222,N_24093);
nor U25035 (N_25035,N_24385,N_24638);
or U25036 (N_25036,N_24887,N_24531);
and U25037 (N_25037,N_24103,N_24653);
and U25038 (N_25038,N_24414,N_24958);
nand U25039 (N_25039,N_24408,N_24435);
nor U25040 (N_25040,N_24491,N_24386);
xor U25041 (N_25041,N_24334,N_24665);
xnor U25042 (N_25042,N_24041,N_24873);
xor U25043 (N_25043,N_24819,N_24399);
and U25044 (N_25044,N_24861,N_24468);
nand U25045 (N_25045,N_24361,N_24369);
nand U25046 (N_25046,N_24319,N_24510);
nor U25047 (N_25047,N_24566,N_24348);
nand U25048 (N_25048,N_24007,N_24610);
nand U25049 (N_25049,N_24613,N_24609);
or U25050 (N_25050,N_24820,N_24081);
and U25051 (N_25051,N_24521,N_24575);
nor U25052 (N_25052,N_24302,N_24935);
or U25053 (N_25053,N_24325,N_24637);
and U25054 (N_25054,N_24923,N_24684);
nand U25055 (N_25055,N_24888,N_24719);
nor U25056 (N_25056,N_24326,N_24423);
or U25057 (N_25057,N_24495,N_24659);
xnor U25058 (N_25058,N_24078,N_24132);
nor U25059 (N_25059,N_24478,N_24260);
nand U25060 (N_25060,N_24560,N_24790);
xnor U25061 (N_25061,N_24118,N_24972);
nand U25062 (N_25062,N_24269,N_24073);
and U25063 (N_25063,N_24466,N_24528);
nand U25064 (N_25064,N_24607,N_24335);
and U25065 (N_25065,N_24753,N_24329);
nand U25066 (N_25066,N_24856,N_24722);
nand U25067 (N_25067,N_24838,N_24496);
xor U25068 (N_25068,N_24784,N_24745);
nor U25069 (N_25069,N_24494,N_24526);
nor U25070 (N_25070,N_24075,N_24293);
nor U25071 (N_25071,N_24500,N_24038);
nand U25072 (N_25072,N_24903,N_24952);
xnor U25073 (N_25073,N_24050,N_24999);
nand U25074 (N_25074,N_24470,N_24446);
xnor U25075 (N_25075,N_24666,N_24062);
or U25076 (N_25076,N_24063,N_24877);
and U25077 (N_25077,N_24064,N_24512);
or U25078 (N_25078,N_24806,N_24811);
nand U25079 (N_25079,N_24677,N_24321);
xnor U25080 (N_25080,N_24987,N_24897);
and U25081 (N_25081,N_24809,N_24271);
nand U25082 (N_25082,N_24804,N_24567);
xor U25083 (N_25083,N_24270,N_24892);
and U25084 (N_25084,N_24805,N_24908);
nor U25085 (N_25085,N_24869,N_24068);
and U25086 (N_25086,N_24590,N_24866);
nand U25087 (N_25087,N_24752,N_24682);
or U25088 (N_25088,N_24099,N_24712);
nand U25089 (N_25089,N_24403,N_24593);
xor U25090 (N_25090,N_24002,N_24652);
xnor U25091 (N_25091,N_24772,N_24009);
xnor U25092 (N_25092,N_24410,N_24830);
or U25093 (N_25093,N_24158,N_24261);
and U25094 (N_25094,N_24225,N_24026);
xor U25095 (N_25095,N_24555,N_24100);
nor U25096 (N_25096,N_24554,N_24913);
or U25097 (N_25097,N_24983,N_24189);
or U25098 (N_25098,N_24562,N_24358);
nand U25099 (N_25099,N_24649,N_24953);
or U25100 (N_25100,N_24455,N_24618);
and U25101 (N_25101,N_24254,N_24247);
nor U25102 (N_25102,N_24199,N_24979);
and U25103 (N_25103,N_24662,N_24272);
xnor U25104 (N_25104,N_24351,N_24810);
xor U25105 (N_25105,N_24742,N_24595);
nor U25106 (N_25106,N_24981,N_24829);
xnor U25107 (N_25107,N_24732,N_24962);
and U25108 (N_25108,N_24119,N_24125);
nor U25109 (N_25109,N_24905,N_24200);
nor U25110 (N_25110,N_24288,N_24214);
nor U25111 (N_25111,N_24264,N_24493);
nand U25112 (N_25112,N_24492,N_24028);
or U25113 (N_25113,N_24502,N_24543);
nand U25114 (N_25114,N_24396,N_24825);
xnor U25115 (N_25115,N_24540,N_24911);
or U25116 (N_25116,N_24497,N_24279);
nor U25117 (N_25117,N_24792,N_24721);
xnor U25118 (N_25118,N_24661,N_24051);
xor U25119 (N_25119,N_24926,N_24770);
nand U25120 (N_25120,N_24463,N_24815);
and U25121 (N_25121,N_24851,N_24854);
and U25122 (N_25122,N_24292,N_24924);
xor U25123 (N_25123,N_24121,N_24611);
or U25124 (N_25124,N_24341,N_24679);
xor U25125 (N_25125,N_24203,N_24299);
and U25126 (N_25126,N_24010,N_24453);
nor U25127 (N_25127,N_24527,N_24161);
and U25128 (N_25128,N_24920,N_24807);
xor U25129 (N_25129,N_24714,N_24978);
xor U25130 (N_25130,N_24579,N_24801);
and U25131 (N_25131,N_24516,N_24720);
and U25132 (N_25132,N_24131,N_24204);
nor U25133 (N_25133,N_24160,N_24896);
or U25134 (N_25134,N_24333,N_24065);
and U25135 (N_25135,N_24223,N_24461);
and U25136 (N_25136,N_24098,N_24197);
xor U25137 (N_25137,N_24879,N_24320);
nor U25138 (N_25138,N_24697,N_24359);
nand U25139 (N_25139,N_24794,N_24951);
nor U25140 (N_25140,N_24212,N_24416);
and U25141 (N_25141,N_24146,N_24744);
or U25142 (N_25142,N_24640,N_24407);
nand U25143 (N_25143,N_24172,N_24159);
nor U25144 (N_25144,N_24032,N_24968);
or U25145 (N_25145,N_24339,N_24621);
and U25146 (N_25146,N_24362,N_24893);
nand U25147 (N_25147,N_24238,N_24600);
nand U25148 (N_25148,N_24969,N_24221);
nand U25149 (N_25149,N_24654,N_24305);
xor U25150 (N_25150,N_24473,N_24355);
nand U25151 (N_25151,N_24789,N_24249);
xnor U25152 (N_25152,N_24835,N_24875);
or U25153 (N_25153,N_24715,N_24283);
nor U25154 (N_25154,N_24291,N_24660);
and U25155 (N_25155,N_24232,N_24523);
xor U25156 (N_25156,N_24601,N_24843);
nand U25157 (N_25157,N_24939,N_24303);
xor U25158 (N_25158,N_24925,N_24013);
nand U25159 (N_25159,N_24023,N_24708);
or U25160 (N_25160,N_24855,N_24900);
and U25161 (N_25161,N_24419,N_24760);
xor U25162 (N_25162,N_24569,N_24895);
nand U25163 (N_25163,N_24703,N_24056);
and U25164 (N_25164,N_24184,N_24090);
nor U25165 (N_25165,N_24821,N_24375);
xnor U25166 (N_25166,N_24284,N_24176);
xor U25167 (N_25167,N_24052,N_24982);
xor U25168 (N_25168,N_24716,N_24522);
nand U25169 (N_25169,N_24239,N_24685);
nor U25170 (N_25170,N_24676,N_24244);
nor U25171 (N_25171,N_24365,N_24381);
nor U25172 (N_25172,N_24899,N_24812);
or U25173 (N_25173,N_24398,N_24533);
nor U25174 (N_25174,N_24559,N_24083);
nor U25175 (N_25175,N_24667,N_24231);
nand U25176 (N_25176,N_24834,N_24404);
nor U25177 (N_25177,N_24154,N_24725);
xor U25178 (N_25178,N_24227,N_24054);
nor U25179 (N_25179,N_24210,N_24848);
nor U25180 (N_25180,N_24229,N_24771);
nand U25181 (N_25181,N_24519,N_24430);
xor U25182 (N_25182,N_24113,N_24450);
xnor U25183 (N_25183,N_24743,N_24352);
or U25184 (N_25184,N_24144,N_24287);
or U25185 (N_25185,N_24641,N_24778);
xor U25186 (N_25186,N_24390,N_24942);
nand U25187 (N_25187,N_24779,N_24415);
and U25188 (N_25188,N_24738,N_24448);
xnor U25189 (N_25189,N_24631,N_24069);
nand U25190 (N_25190,N_24630,N_24773);
nor U25191 (N_25191,N_24524,N_24699);
nor U25192 (N_25192,N_24454,N_24717);
and U25193 (N_25193,N_24443,N_24027);
nor U25194 (N_25194,N_24927,N_24187);
and U25195 (N_25195,N_24646,N_24606);
or U25196 (N_25196,N_24731,N_24997);
xor U25197 (N_25197,N_24583,N_24273);
or U25198 (N_25198,N_24833,N_24483);
nand U25199 (N_25199,N_24766,N_24024);
nor U25200 (N_25200,N_24433,N_24263);
xor U25201 (N_25201,N_24992,N_24758);
xor U25202 (N_25202,N_24447,N_24763);
or U25203 (N_25203,N_24506,N_24356);
and U25204 (N_25204,N_24445,N_24599);
xnor U25205 (N_25205,N_24740,N_24694);
nor U25206 (N_25206,N_24162,N_24802);
or U25207 (N_25207,N_24363,N_24503);
xnor U25208 (N_25208,N_24373,N_24438);
or U25209 (N_25209,N_24209,N_24765);
nand U25210 (N_25210,N_24036,N_24929);
xnor U25211 (N_25211,N_24071,N_24253);
and U25212 (N_25212,N_24741,N_24173);
nand U25213 (N_25213,N_24636,N_24850);
xnor U25214 (N_25214,N_24267,N_24541);
or U25215 (N_25215,N_24127,N_24469);
and U25216 (N_25216,N_24309,N_24803);
or U25217 (N_25217,N_24233,N_24328);
nand U25218 (N_25218,N_24307,N_24984);
or U25219 (N_25219,N_24775,N_24624);
nand U25220 (N_25220,N_24530,N_24354);
or U25221 (N_25221,N_24620,N_24689);
xor U25222 (N_25222,N_24639,N_24781);
nand U25223 (N_25223,N_24910,N_24317);
xnor U25224 (N_25224,N_24870,N_24019);
or U25225 (N_25225,N_24735,N_24370);
xnor U25226 (N_25226,N_24564,N_24021);
nand U25227 (N_25227,N_24648,N_24933);
or U25228 (N_25228,N_24919,N_24346);
nor U25229 (N_25229,N_24529,N_24025);
nand U25230 (N_25230,N_24256,N_24669);
nand U25231 (N_25231,N_24191,N_24602);
or U25232 (N_25232,N_24691,N_24644);
or U25233 (N_25233,N_24109,N_24175);
and U25234 (N_25234,N_24536,N_24241);
and U25235 (N_25235,N_24723,N_24364);
and U25236 (N_25236,N_24693,N_24005);
nand U25237 (N_25237,N_24265,N_24420);
nor U25238 (N_25238,N_24067,N_24576);
xnor U25239 (N_25239,N_24499,N_24477);
nor U25240 (N_25240,N_24647,N_24045);
or U25241 (N_25241,N_24553,N_24996);
nand U25242 (N_25242,N_24836,N_24084);
nor U25243 (N_25243,N_24974,N_24993);
nand U25244 (N_25244,N_24156,N_24718);
or U25245 (N_25245,N_24035,N_24605);
nand U25246 (N_25246,N_24816,N_24846);
or U25247 (N_25247,N_24349,N_24300);
nand U25248 (N_25248,N_24580,N_24608);
xor U25249 (N_25249,N_24928,N_24702);
nor U25250 (N_25250,N_24436,N_24387);
nor U25251 (N_25251,N_24289,N_24245);
nand U25252 (N_25252,N_24990,N_24322);
nor U25253 (N_25253,N_24757,N_24114);
and U25254 (N_25254,N_24486,N_24168);
or U25255 (N_25255,N_24000,N_24936);
nand U25256 (N_25256,N_24101,N_24234);
nand U25257 (N_25257,N_24393,N_24343);
or U25258 (N_25258,N_24894,N_24220);
xnor U25259 (N_25259,N_24860,N_24490);
xor U25260 (N_25260,N_24550,N_24310);
or U25261 (N_25261,N_24006,N_24082);
xnor U25262 (N_25262,N_24561,N_24658);
and U25263 (N_25263,N_24947,N_24525);
nand U25264 (N_25264,N_24614,N_24571);
or U25265 (N_25265,N_24034,N_24484);
and U25266 (N_25266,N_24479,N_24603);
and U25267 (N_25267,N_24547,N_24055);
nor U25268 (N_25268,N_24331,N_24700);
xor U25269 (N_25269,N_24228,N_24970);
nand U25270 (N_25270,N_24642,N_24439);
xor U25271 (N_25271,N_24115,N_24474);
nor U25272 (N_25272,N_24251,N_24143);
xor U25273 (N_25273,N_24754,N_24736);
xor U25274 (N_25274,N_24788,N_24087);
nor U25275 (N_25275,N_24863,N_24169);
or U25276 (N_25276,N_24739,N_24872);
or U25277 (N_25277,N_24767,N_24934);
or U25278 (N_25278,N_24596,N_24344);
nor U25279 (N_25279,N_24441,N_24865);
nand U25280 (N_25280,N_24998,N_24237);
and U25281 (N_25281,N_24960,N_24504);
xnor U25282 (N_25282,N_24117,N_24138);
and U25283 (N_25283,N_24931,N_24015);
nor U25284 (N_25284,N_24318,N_24155);
nor U25285 (N_25285,N_24777,N_24342);
nor U25286 (N_25286,N_24456,N_24337);
nor U25287 (N_25287,N_24762,N_24625);
nand U25288 (N_25288,N_24148,N_24656);
xor U25289 (N_25289,N_24280,N_24350);
or U25290 (N_25290,N_24881,N_24565);
nand U25291 (N_25291,N_24769,N_24017);
or U25292 (N_25292,N_24437,N_24205);
nand U25293 (N_25293,N_24889,N_24482);
nor U25294 (N_25294,N_24574,N_24515);
or U25295 (N_25295,N_24088,N_24876);
xnor U25296 (N_25296,N_24498,N_24692);
nand U25297 (N_25297,N_24710,N_24388);
or U25298 (N_25298,N_24427,N_24224);
nor U25299 (N_25299,N_24517,N_24629);
or U25300 (N_25300,N_24120,N_24030);
and U25301 (N_25301,N_24316,N_24432);
or U25302 (N_25302,N_24460,N_24243);
or U25303 (N_25303,N_24250,N_24587);
and U25304 (N_25304,N_24313,N_24882);
or U25305 (N_25305,N_24966,N_24230);
nand U25306 (N_25306,N_24475,N_24130);
and U25307 (N_25307,N_24304,N_24518);
and U25308 (N_25308,N_24886,N_24042);
nand U25309 (N_25309,N_24626,N_24391);
xor U25310 (N_25310,N_24374,N_24110);
nand U25311 (N_25311,N_24840,N_24384);
nor U25312 (N_25312,N_24094,N_24290);
nor U25313 (N_25313,N_24294,N_24201);
nor U25314 (N_25314,N_24297,N_24734);
and U25315 (N_25315,N_24336,N_24409);
or U25316 (N_25316,N_24061,N_24395);
nand U25317 (N_25317,N_24800,N_24198);
and U25318 (N_25318,N_24458,N_24977);
nor U25319 (N_25319,N_24573,N_24729);
nor U25320 (N_25320,N_24548,N_24826);
nand U25321 (N_25321,N_24058,N_24582);
nor U25322 (N_25322,N_24557,N_24123);
nand U25323 (N_25323,N_24808,N_24246);
and U25324 (N_25324,N_24338,N_24372);
and U25325 (N_25325,N_24164,N_24783);
xnor U25326 (N_25326,N_24864,N_24105);
nand U25327 (N_25327,N_24696,N_24376);
or U25328 (N_25328,N_24286,N_24628);
xor U25329 (N_25329,N_24180,N_24853);
xnor U25330 (N_25330,N_24049,N_24793);
xnor U25331 (N_25331,N_24552,N_24142);
or U25332 (N_25332,N_24989,N_24429);
xor U25333 (N_25333,N_24406,N_24001);
or U25334 (N_25334,N_24428,N_24276);
nand U25335 (N_25335,N_24563,N_24186);
and U25336 (N_25336,N_24537,N_24884);
nor U25337 (N_25337,N_24086,N_24314);
nand U25338 (N_25338,N_24192,N_24586);
or U25339 (N_25339,N_24713,N_24029);
and U25340 (N_25340,N_24578,N_24688);
nor U25341 (N_25341,N_24122,N_24047);
nor U25342 (N_25342,N_24921,N_24133);
or U25343 (N_25343,N_24031,N_24444);
and U25344 (N_25344,N_24020,N_24871);
nor U25345 (N_25345,N_24672,N_24724);
nor U25346 (N_25346,N_24170,N_24405);
nor U25347 (N_25347,N_24033,N_24501);
nand U25348 (N_25348,N_24177,N_24687);
xor U25349 (N_25349,N_24467,N_24986);
nor U25350 (N_25350,N_24549,N_24706);
and U25351 (N_25351,N_24711,N_24780);
and U25352 (N_25352,N_24412,N_24219);
nor U25353 (N_25353,N_24671,N_24912);
nor U25354 (N_25354,N_24818,N_24141);
xor U25355 (N_25355,N_24037,N_24259);
nand U25356 (N_25356,N_24096,N_24558);
or U25357 (N_25357,N_24798,N_24768);
or U25358 (N_25358,N_24323,N_24060);
or U25359 (N_25359,N_24867,N_24965);
and U25360 (N_25360,N_24916,N_24898);
or U25361 (N_25361,N_24511,N_24298);
nor U25362 (N_25362,N_24532,N_24681);
nand U25363 (N_25363,N_24275,N_24213);
nand U25364 (N_25364,N_24592,N_24401);
and U25365 (N_25365,N_24904,N_24673);
nor U25366 (N_25366,N_24664,N_24040);
nor U25367 (N_25367,N_24849,N_24046);
nor U25368 (N_25368,N_24206,N_24003);
xor U25369 (N_25369,N_24179,N_24941);
xor U25370 (N_25370,N_24615,N_24755);
nand U25371 (N_25371,N_24092,N_24330);
xnor U25372 (N_25372,N_24591,N_24347);
and U25373 (N_25373,N_24786,N_24874);
xor U25374 (N_25374,N_24594,N_24909);
or U25375 (N_25375,N_24612,N_24380);
nand U25376 (N_25376,N_24489,N_24218);
xnor U25377 (N_25377,N_24868,N_24814);
xnor U25378 (N_25378,N_24340,N_24839);
xnor U25379 (N_25379,N_24426,N_24857);
xnor U25380 (N_25380,N_24514,N_24248);
or U25381 (N_25381,N_24085,N_24598);
or U25382 (N_25382,N_24080,N_24556);
or U25383 (N_25383,N_24306,N_24236);
nand U25384 (N_25384,N_24147,N_24535);
or U25385 (N_25385,N_24208,N_24413);
or U25386 (N_25386,N_24418,N_24417);
and U25387 (N_25387,N_24973,N_24847);
xnor U25388 (N_25388,N_24799,N_24570);
nor U25389 (N_25389,N_24568,N_24076);
nor U25390 (N_25390,N_24938,N_24185);
and U25391 (N_25391,N_24589,N_24481);
and U25392 (N_25392,N_24759,N_24278);
or U25393 (N_25393,N_24619,N_24627);
nand U25394 (N_25394,N_24930,N_24505);
xnor U25395 (N_25395,N_24971,N_24211);
or U25396 (N_25396,N_24967,N_24577);
nor U25397 (N_25397,N_24686,N_24883);
or U25398 (N_25398,N_24813,N_24622);
nor U25399 (N_25399,N_24487,N_24862);
nor U25400 (N_25400,N_24296,N_24043);
or U25401 (N_25401,N_24746,N_24137);
xor U25402 (N_25402,N_24980,N_24635);
and U25403 (N_25403,N_24472,N_24831);
or U25404 (N_25404,N_24091,N_24016);
or U25405 (N_25405,N_24507,N_24301);
xnor U25406 (N_25406,N_24787,N_24457);
nor U25407 (N_25407,N_24539,N_24650);
xnor U25408 (N_25408,N_24795,N_24976);
nand U25409 (N_25409,N_24957,N_24136);
nor U25410 (N_25410,N_24190,N_24216);
xor U25411 (N_25411,N_24891,N_24616);
nand U25412 (N_25412,N_24751,N_24345);
nand U25413 (N_25413,N_24150,N_24207);
xnor U25414 (N_25414,N_24985,N_24785);
xor U25415 (N_25415,N_24954,N_24285);
or U25416 (N_25416,N_24074,N_24152);
and U25417 (N_25417,N_24465,N_24488);
or U25418 (N_25418,N_24378,N_24106);
nor U25419 (N_25419,N_24111,N_24950);
xor U25420 (N_25420,N_24353,N_24424);
xor U25421 (N_25421,N_24668,N_24728);
nand U25422 (N_25422,N_24914,N_24072);
nand U25423 (N_25423,N_24657,N_24705);
xor U25424 (N_25424,N_24906,N_24171);
and U25425 (N_25425,N_24116,N_24922);
and U25426 (N_25426,N_24379,N_24709);
or U25427 (N_25427,N_24651,N_24044);
nand U25428 (N_25428,N_24774,N_24707);
xor U25429 (N_25429,N_24604,N_24623);
xnor U25430 (N_25430,N_24509,N_24217);
and U25431 (N_25431,N_24011,N_24066);
or U25432 (N_25432,N_24726,N_24262);
and U25433 (N_25433,N_24451,N_24949);
xnor U25434 (N_25434,N_24167,N_24242);
nor U25435 (N_25435,N_24126,N_24464);
or U25436 (N_25436,N_24617,N_24149);
xor U25437 (N_25437,N_24332,N_24674);
nand U25438 (N_25438,N_24698,N_24070);
nand U25439 (N_25439,N_24135,N_24761);
and U25440 (N_25440,N_24678,N_24166);
nand U25441 (N_25441,N_24004,N_24095);
nor U25442 (N_25442,N_24107,N_24655);
nor U25443 (N_25443,N_24315,N_24823);
nor U25444 (N_25444,N_24964,N_24112);
or U25445 (N_25445,N_24295,N_24480);
xnor U25446 (N_25446,N_24274,N_24268);
xor U25447 (N_25447,N_24383,N_24194);
or U25448 (N_25448,N_24670,N_24946);
and U25449 (N_25449,N_24476,N_24513);
and U25450 (N_25450,N_24012,N_24859);
and U25451 (N_25451,N_24151,N_24048);
nand U25452 (N_25452,N_24235,N_24991);
xor U25453 (N_25453,N_24632,N_24959);
or U25454 (N_25454,N_24057,N_24937);
or U25455 (N_25455,N_24394,N_24584);
xnor U25456 (N_25456,N_24282,N_24327);
nand U25457 (N_25457,N_24764,N_24108);
and U25458 (N_25458,N_24193,N_24485);
or U25459 (N_25459,N_24022,N_24421);
xor U25460 (N_25460,N_24842,N_24737);
nor U25461 (N_25461,N_24956,N_24588);
xnor U25462 (N_25462,N_24963,N_24145);
xor U25463 (N_25463,N_24377,N_24258);
nor U25464 (N_25464,N_24104,N_24367);
nand U25465 (N_25465,N_24188,N_24079);
or U25466 (N_25466,N_24690,N_24129);
xnor U25467 (N_25467,N_24845,N_24683);
xor U25468 (N_25468,N_24014,N_24841);
or U25469 (N_25469,N_24538,N_24901);
xor U25470 (N_25470,N_24634,N_24880);
or U25471 (N_25471,N_24442,N_24311);
xor U25472 (N_25472,N_24701,N_24542);
xor U25473 (N_25473,N_24183,N_24402);
nand U25474 (N_25474,N_24059,N_24425);
xor U25475 (N_25475,N_24178,N_24266);
xor U25476 (N_25476,N_24366,N_24534);
or U25477 (N_25477,N_24852,N_24704);
xor U25478 (N_25478,N_24165,N_24411);
or U25479 (N_25479,N_24918,N_24089);
nor U25480 (N_25480,N_24597,N_24948);
nor U25481 (N_25481,N_24153,N_24389);
nand U25482 (N_25482,N_24053,N_24643);
nor U25483 (N_25483,N_24226,N_24544);
or U25484 (N_25484,N_24134,N_24546);
or U25485 (N_25485,N_24452,N_24124);
nand U25486 (N_25486,N_24572,N_24782);
nand U25487 (N_25487,N_24368,N_24431);
nor U25488 (N_25488,N_24915,N_24917);
xor U25489 (N_25489,N_24392,N_24382);
xor U25490 (N_25490,N_24750,N_24747);
nor U25491 (N_25491,N_24400,N_24545);
nand U25492 (N_25492,N_24955,N_24097);
nor U25493 (N_25493,N_24943,N_24824);
and U25494 (N_25494,N_24360,N_24756);
or U25495 (N_25495,N_24196,N_24440);
nand U25496 (N_25496,N_24018,N_24312);
or U25497 (N_25497,N_24791,N_24663);
or U25498 (N_25498,N_24255,N_24215);
nor U25499 (N_25499,N_24277,N_24174);
xnor U25500 (N_25500,N_24474,N_24876);
xor U25501 (N_25501,N_24221,N_24447);
nor U25502 (N_25502,N_24866,N_24414);
nand U25503 (N_25503,N_24275,N_24840);
nor U25504 (N_25504,N_24821,N_24741);
and U25505 (N_25505,N_24995,N_24839);
or U25506 (N_25506,N_24169,N_24240);
and U25507 (N_25507,N_24163,N_24455);
nand U25508 (N_25508,N_24299,N_24394);
and U25509 (N_25509,N_24847,N_24290);
xor U25510 (N_25510,N_24005,N_24225);
or U25511 (N_25511,N_24086,N_24063);
xnor U25512 (N_25512,N_24034,N_24712);
nand U25513 (N_25513,N_24004,N_24661);
or U25514 (N_25514,N_24638,N_24254);
xnor U25515 (N_25515,N_24941,N_24912);
or U25516 (N_25516,N_24086,N_24493);
nor U25517 (N_25517,N_24878,N_24278);
nand U25518 (N_25518,N_24348,N_24556);
or U25519 (N_25519,N_24984,N_24306);
xnor U25520 (N_25520,N_24523,N_24651);
xnor U25521 (N_25521,N_24161,N_24143);
nand U25522 (N_25522,N_24055,N_24232);
or U25523 (N_25523,N_24029,N_24740);
xor U25524 (N_25524,N_24180,N_24800);
xor U25525 (N_25525,N_24498,N_24251);
nand U25526 (N_25526,N_24851,N_24947);
and U25527 (N_25527,N_24363,N_24041);
and U25528 (N_25528,N_24360,N_24396);
nand U25529 (N_25529,N_24834,N_24050);
nor U25530 (N_25530,N_24026,N_24262);
nor U25531 (N_25531,N_24054,N_24194);
nand U25532 (N_25532,N_24631,N_24048);
nand U25533 (N_25533,N_24496,N_24052);
and U25534 (N_25534,N_24017,N_24635);
or U25535 (N_25535,N_24440,N_24295);
or U25536 (N_25536,N_24213,N_24743);
nor U25537 (N_25537,N_24762,N_24824);
and U25538 (N_25538,N_24468,N_24152);
nand U25539 (N_25539,N_24786,N_24037);
or U25540 (N_25540,N_24688,N_24581);
and U25541 (N_25541,N_24311,N_24190);
nor U25542 (N_25542,N_24180,N_24612);
or U25543 (N_25543,N_24774,N_24608);
or U25544 (N_25544,N_24695,N_24775);
or U25545 (N_25545,N_24953,N_24156);
or U25546 (N_25546,N_24888,N_24246);
nand U25547 (N_25547,N_24792,N_24629);
xor U25548 (N_25548,N_24523,N_24383);
xor U25549 (N_25549,N_24337,N_24133);
nor U25550 (N_25550,N_24394,N_24558);
and U25551 (N_25551,N_24231,N_24183);
nand U25552 (N_25552,N_24604,N_24644);
xnor U25553 (N_25553,N_24918,N_24368);
or U25554 (N_25554,N_24387,N_24333);
and U25555 (N_25555,N_24910,N_24451);
nor U25556 (N_25556,N_24827,N_24663);
or U25557 (N_25557,N_24776,N_24190);
or U25558 (N_25558,N_24257,N_24602);
nand U25559 (N_25559,N_24344,N_24547);
and U25560 (N_25560,N_24505,N_24284);
nor U25561 (N_25561,N_24467,N_24773);
nand U25562 (N_25562,N_24609,N_24517);
or U25563 (N_25563,N_24749,N_24590);
and U25564 (N_25564,N_24085,N_24646);
or U25565 (N_25565,N_24573,N_24339);
xnor U25566 (N_25566,N_24290,N_24855);
nor U25567 (N_25567,N_24182,N_24534);
or U25568 (N_25568,N_24637,N_24869);
nor U25569 (N_25569,N_24670,N_24469);
nor U25570 (N_25570,N_24445,N_24614);
or U25571 (N_25571,N_24358,N_24592);
xor U25572 (N_25572,N_24767,N_24337);
xor U25573 (N_25573,N_24183,N_24199);
nor U25574 (N_25574,N_24345,N_24423);
nor U25575 (N_25575,N_24046,N_24347);
nor U25576 (N_25576,N_24352,N_24388);
xnor U25577 (N_25577,N_24815,N_24923);
nor U25578 (N_25578,N_24939,N_24198);
xor U25579 (N_25579,N_24476,N_24488);
and U25580 (N_25580,N_24540,N_24714);
nor U25581 (N_25581,N_24365,N_24356);
and U25582 (N_25582,N_24854,N_24883);
xnor U25583 (N_25583,N_24384,N_24858);
or U25584 (N_25584,N_24480,N_24420);
or U25585 (N_25585,N_24474,N_24460);
nand U25586 (N_25586,N_24627,N_24718);
and U25587 (N_25587,N_24291,N_24289);
nand U25588 (N_25588,N_24468,N_24073);
and U25589 (N_25589,N_24086,N_24883);
or U25590 (N_25590,N_24637,N_24287);
nand U25591 (N_25591,N_24384,N_24063);
and U25592 (N_25592,N_24339,N_24591);
nand U25593 (N_25593,N_24474,N_24959);
and U25594 (N_25594,N_24952,N_24490);
or U25595 (N_25595,N_24688,N_24211);
xnor U25596 (N_25596,N_24179,N_24520);
or U25597 (N_25597,N_24654,N_24207);
nor U25598 (N_25598,N_24658,N_24645);
nand U25599 (N_25599,N_24035,N_24431);
nor U25600 (N_25600,N_24330,N_24950);
xnor U25601 (N_25601,N_24496,N_24403);
xor U25602 (N_25602,N_24052,N_24199);
or U25603 (N_25603,N_24979,N_24026);
and U25604 (N_25604,N_24907,N_24880);
nand U25605 (N_25605,N_24119,N_24243);
nand U25606 (N_25606,N_24962,N_24819);
and U25607 (N_25607,N_24912,N_24106);
or U25608 (N_25608,N_24169,N_24256);
xor U25609 (N_25609,N_24856,N_24519);
nor U25610 (N_25610,N_24734,N_24013);
nor U25611 (N_25611,N_24511,N_24876);
or U25612 (N_25612,N_24063,N_24762);
nor U25613 (N_25613,N_24487,N_24452);
or U25614 (N_25614,N_24440,N_24471);
and U25615 (N_25615,N_24586,N_24109);
and U25616 (N_25616,N_24268,N_24401);
nor U25617 (N_25617,N_24729,N_24363);
or U25618 (N_25618,N_24858,N_24595);
nor U25619 (N_25619,N_24694,N_24874);
nor U25620 (N_25620,N_24510,N_24429);
nand U25621 (N_25621,N_24411,N_24420);
and U25622 (N_25622,N_24365,N_24562);
nand U25623 (N_25623,N_24991,N_24076);
and U25624 (N_25624,N_24249,N_24600);
and U25625 (N_25625,N_24544,N_24397);
nand U25626 (N_25626,N_24144,N_24614);
or U25627 (N_25627,N_24827,N_24015);
xor U25628 (N_25628,N_24968,N_24459);
or U25629 (N_25629,N_24105,N_24905);
and U25630 (N_25630,N_24307,N_24348);
nand U25631 (N_25631,N_24523,N_24874);
or U25632 (N_25632,N_24607,N_24471);
nor U25633 (N_25633,N_24106,N_24040);
xor U25634 (N_25634,N_24195,N_24936);
nand U25635 (N_25635,N_24007,N_24244);
or U25636 (N_25636,N_24933,N_24536);
or U25637 (N_25637,N_24213,N_24561);
nand U25638 (N_25638,N_24346,N_24830);
or U25639 (N_25639,N_24780,N_24140);
and U25640 (N_25640,N_24015,N_24150);
xnor U25641 (N_25641,N_24524,N_24762);
nand U25642 (N_25642,N_24681,N_24704);
or U25643 (N_25643,N_24599,N_24283);
and U25644 (N_25644,N_24167,N_24711);
or U25645 (N_25645,N_24683,N_24940);
or U25646 (N_25646,N_24451,N_24287);
xor U25647 (N_25647,N_24365,N_24136);
nor U25648 (N_25648,N_24685,N_24269);
and U25649 (N_25649,N_24805,N_24716);
xnor U25650 (N_25650,N_24907,N_24482);
and U25651 (N_25651,N_24878,N_24586);
or U25652 (N_25652,N_24277,N_24722);
nand U25653 (N_25653,N_24378,N_24863);
or U25654 (N_25654,N_24449,N_24663);
and U25655 (N_25655,N_24328,N_24445);
or U25656 (N_25656,N_24948,N_24829);
nor U25657 (N_25657,N_24086,N_24975);
nor U25658 (N_25658,N_24766,N_24005);
and U25659 (N_25659,N_24806,N_24877);
nor U25660 (N_25660,N_24515,N_24057);
nor U25661 (N_25661,N_24486,N_24182);
or U25662 (N_25662,N_24646,N_24390);
and U25663 (N_25663,N_24798,N_24351);
xnor U25664 (N_25664,N_24095,N_24631);
and U25665 (N_25665,N_24104,N_24125);
and U25666 (N_25666,N_24021,N_24610);
or U25667 (N_25667,N_24100,N_24081);
and U25668 (N_25668,N_24027,N_24168);
nand U25669 (N_25669,N_24241,N_24760);
nor U25670 (N_25670,N_24634,N_24853);
nand U25671 (N_25671,N_24391,N_24876);
and U25672 (N_25672,N_24453,N_24067);
xor U25673 (N_25673,N_24481,N_24602);
xnor U25674 (N_25674,N_24165,N_24895);
nor U25675 (N_25675,N_24126,N_24601);
or U25676 (N_25676,N_24198,N_24958);
xnor U25677 (N_25677,N_24458,N_24308);
xnor U25678 (N_25678,N_24443,N_24109);
and U25679 (N_25679,N_24442,N_24238);
nand U25680 (N_25680,N_24787,N_24602);
and U25681 (N_25681,N_24031,N_24496);
xnor U25682 (N_25682,N_24205,N_24814);
and U25683 (N_25683,N_24275,N_24039);
nand U25684 (N_25684,N_24215,N_24707);
xor U25685 (N_25685,N_24587,N_24772);
and U25686 (N_25686,N_24048,N_24300);
nand U25687 (N_25687,N_24682,N_24206);
or U25688 (N_25688,N_24116,N_24444);
or U25689 (N_25689,N_24351,N_24647);
xor U25690 (N_25690,N_24282,N_24189);
and U25691 (N_25691,N_24687,N_24509);
nand U25692 (N_25692,N_24827,N_24304);
and U25693 (N_25693,N_24387,N_24835);
and U25694 (N_25694,N_24386,N_24439);
and U25695 (N_25695,N_24684,N_24413);
and U25696 (N_25696,N_24202,N_24635);
or U25697 (N_25697,N_24258,N_24481);
xnor U25698 (N_25698,N_24375,N_24262);
or U25699 (N_25699,N_24506,N_24968);
nand U25700 (N_25700,N_24176,N_24102);
xor U25701 (N_25701,N_24579,N_24335);
or U25702 (N_25702,N_24628,N_24980);
xor U25703 (N_25703,N_24628,N_24019);
nand U25704 (N_25704,N_24045,N_24666);
and U25705 (N_25705,N_24563,N_24244);
xnor U25706 (N_25706,N_24994,N_24129);
nor U25707 (N_25707,N_24557,N_24039);
nand U25708 (N_25708,N_24556,N_24431);
and U25709 (N_25709,N_24307,N_24852);
nor U25710 (N_25710,N_24145,N_24647);
nor U25711 (N_25711,N_24245,N_24010);
xor U25712 (N_25712,N_24231,N_24032);
nor U25713 (N_25713,N_24886,N_24301);
nor U25714 (N_25714,N_24910,N_24049);
or U25715 (N_25715,N_24628,N_24839);
nor U25716 (N_25716,N_24066,N_24648);
nand U25717 (N_25717,N_24550,N_24635);
nor U25718 (N_25718,N_24294,N_24343);
or U25719 (N_25719,N_24682,N_24037);
or U25720 (N_25720,N_24375,N_24178);
nor U25721 (N_25721,N_24028,N_24167);
or U25722 (N_25722,N_24108,N_24153);
or U25723 (N_25723,N_24234,N_24563);
nor U25724 (N_25724,N_24129,N_24851);
or U25725 (N_25725,N_24399,N_24026);
nand U25726 (N_25726,N_24859,N_24839);
and U25727 (N_25727,N_24725,N_24671);
or U25728 (N_25728,N_24115,N_24864);
xnor U25729 (N_25729,N_24017,N_24895);
nand U25730 (N_25730,N_24008,N_24688);
xor U25731 (N_25731,N_24818,N_24150);
nand U25732 (N_25732,N_24316,N_24138);
nor U25733 (N_25733,N_24330,N_24380);
nand U25734 (N_25734,N_24384,N_24134);
and U25735 (N_25735,N_24841,N_24139);
nand U25736 (N_25736,N_24950,N_24365);
and U25737 (N_25737,N_24109,N_24504);
or U25738 (N_25738,N_24937,N_24186);
and U25739 (N_25739,N_24826,N_24342);
nor U25740 (N_25740,N_24437,N_24338);
nor U25741 (N_25741,N_24865,N_24644);
and U25742 (N_25742,N_24998,N_24474);
or U25743 (N_25743,N_24425,N_24283);
nor U25744 (N_25744,N_24169,N_24679);
nor U25745 (N_25745,N_24849,N_24043);
nand U25746 (N_25746,N_24596,N_24968);
nor U25747 (N_25747,N_24747,N_24325);
xor U25748 (N_25748,N_24868,N_24391);
nor U25749 (N_25749,N_24186,N_24052);
nor U25750 (N_25750,N_24009,N_24763);
xor U25751 (N_25751,N_24883,N_24885);
or U25752 (N_25752,N_24201,N_24908);
or U25753 (N_25753,N_24738,N_24156);
nor U25754 (N_25754,N_24640,N_24799);
and U25755 (N_25755,N_24000,N_24586);
or U25756 (N_25756,N_24127,N_24096);
nor U25757 (N_25757,N_24244,N_24210);
nand U25758 (N_25758,N_24293,N_24922);
xor U25759 (N_25759,N_24190,N_24154);
nor U25760 (N_25760,N_24969,N_24313);
nand U25761 (N_25761,N_24652,N_24538);
nand U25762 (N_25762,N_24206,N_24356);
and U25763 (N_25763,N_24817,N_24210);
and U25764 (N_25764,N_24932,N_24369);
nand U25765 (N_25765,N_24922,N_24666);
and U25766 (N_25766,N_24733,N_24349);
nor U25767 (N_25767,N_24512,N_24295);
nand U25768 (N_25768,N_24602,N_24683);
and U25769 (N_25769,N_24731,N_24872);
and U25770 (N_25770,N_24694,N_24369);
or U25771 (N_25771,N_24347,N_24779);
xnor U25772 (N_25772,N_24367,N_24686);
and U25773 (N_25773,N_24182,N_24338);
and U25774 (N_25774,N_24780,N_24803);
or U25775 (N_25775,N_24770,N_24217);
nand U25776 (N_25776,N_24680,N_24738);
nand U25777 (N_25777,N_24024,N_24422);
nand U25778 (N_25778,N_24763,N_24794);
nand U25779 (N_25779,N_24605,N_24898);
xor U25780 (N_25780,N_24847,N_24942);
nand U25781 (N_25781,N_24191,N_24638);
nand U25782 (N_25782,N_24839,N_24427);
xor U25783 (N_25783,N_24043,N_24866);
or U25784 (N_25784,N_24990,N_24468);
and U25785 (N_25785,N_24272,N_24690);
and U25786 (N_25786,N_24791,N_24096);
xnor U25787 (N_25787,N_24671,N_24770);
xnor U25788 (N_25788,N_24138,N_24001);
and U25789 (N_25789,N_24278,N_24571);
and U25790 (N_25790,N_24673,N_24569);
xor U25791 (N_25791,N_24321,N_24477);
nand U25792 (N_25792,N_24218,N_24674);
nor U25793 (N_25793,N_24855,N_24737);
nor U25794 (N_25794,N_24315,N_24087);
nor U25795 (N_25795,N_24587,N_24573);
and U25796 (N_25796,N_24835,N_24778);
nand U25797 (N_25797,N_24809,N_24190);
nand U25798 (N_25798,N_24660,N_24403);
nor U25799 (N_25799,N_24692,N_24094);
nor U25800 (N_25800,N_24575,N_24032);
xnor U25801 (N_25801,N_24061,N_24049);
nor U25802 (N_25802,N_24794,N_24515);
xnor U25803 (N_25803,N_24360,N_24048);
and U25804 (N_25804,N_24378,N_24020);
and U25805 (N_25805,N_24415,N_24287);
nor U25806 (N_25806,N_24098,N_24891);
and U25807 (N_25807,N_24299,N_24906);
xnor U25808 (N_25808,N_24704,N_24004);
nand U25809 (N_25809,N_24133,N_24925);
and U25810 (N_25810,N_24844,N_24015);
or U25811 (N_25811,N_24105,N_24487);
or U25812 (N_25812,N_24051,N_24959);
or U25813 (N_25813,N_24493,N_24758);
or U25814 (N_25814,N_24560,N_24291);
xnor U25815 (N_25815,N_24037,N_24705);
and U25816 (N_25816,N_24302,N_24932);
xor U25817 (N_25817,N_24597,N_24483);
nor U25818 (N_25818,N_24178,N_24115);
nand U25819 (N_25819,N_24544,N_24826);
xnor U25820 (N_25820,N_24526,N_24035);
or U25821 (N_25821,N_24398,N_24600);
xnor U25822 (N_25822,N_24824,N_24765);
nor U25823 (N_25823,N_24760,N_24398);
nand U25824 (N_25824,N_24425,N_24400);
nor U25825 (N_25825,N_24687,N_24237);
nand U25826 (N_25826,N_24935,N_24593);
nor U25827 (N_25827,N_24885,N_24133);
nand U25828 (N_25828,N_24867,N_24692);
and U25829 (N_25829,N_24004,N_24008);
and U25830 (N_25830,N_24851,N_24300);
or U25831 (N_25831,N_24691,N_24470);
and U25832 (N_25832,N_24856,N_24026);
xnor U25833 (N_25833,N_24133,N_24701);
xnor U25834 (N_25834,N_24853,N_24468);
xor U25835 (N_25835,N_24109,N_24194);
or U25836 (N_25836,N_24103,N_24436);
nor U25837 (N_25837,N_24695,N_24831);
xnor U25838 (N_25838,N_24732,N_24662);
and U25839 (N_25839,N_24666,N_24774);
nand U25840 (N_25840,N_24783,N_24324);
and U25841 (N_25841,N_24328,N_24299);
nor U25842 (N_25842,N_24356,N_24996);
or U25843 (N_25843,N_24765,N_24477);
and U25844 (N_25844,N_24326,N_24378);
nor U25845 (N_25845,N_24135,N_24923);
and U25846 (N_25846,N_24315,N_24767);
xnor U25847 (N_25847,N_24216,N_24064);
or U25848 (N_25848,N_24311,N_24711);
or U25849 (N_25849,N_24581,N_24536);
nand U25850 (N_25850,N_24567,N_24307);
nor U25851 (N_25851,N_24857,N_24469);
nand U25852 (N_25852,N_24988,N_24583);
or U25853 (N_25853,N_24283,N_24422);
nand U25854 (N_25854,N_24187,N_24499);
and U25855 (N_25855,N_24300,N_24628);
nor U25856 (N_25856,N_24180,N_24126);
xnor U25857 (N_25857,N_24578,N_24677);
and U25858 (N_25858,N_24538,N_24713);
xor U25859 (N_25859,N_24752,N_24930);
and U25860 (N_25860,N_24663,N_24670);
and U25861 (N_25861,N_24105,N_24583);
or U25862 (N_25862,N_24218,N_24867);
and U25863 (N_25863,N_24757,N_24522);
or U25864 (N_25864,N_24838,N_24157);
nor U25865 (N_25865,N_24154,N_24376);
or U25866 (N_25866,N_24631,N_24186);
nor U25867 (N_25867,N_24465,N_24910);
or U25868 (N_25868,N_24006,N_24073);
xnor U25869 (N_25869,N_24945,N_24871);
nor U25870 (N_25870,N_24680,N_24124);
xnor U25871 (N_25871,N_24805,N_24609);
xnor U25872 (N_25872,N_24704,N_24030);
or U25873 (N_25873,N_24190,N_24066);
xnor U25874 (N_25874,N_24897,N_24385);
and U25875 (N_25875,N_24689,N_24537);
nor U25876 (N_25876,N_24661,N_24705);
nand U25877 (N_25877,N_24668,N_24761);
nor U25878 (N_25878,N_24965,N_24485);
and U25879 (N_25879,N_24154,N_24694);
and U25880 (N_25880,N_24243,N_24141);
xnor U25881 (N_25881,N_24928,N_24762);
xor U25882 (N_25882,N_24626,N_24993);
nor U25883 (N_25883,N_24867,N_24841);
nor U25884 (N_25884,N_24779,N_24477);
nor U25885 (N_25885,N_24156,N_24803);
xnor U25886 (N_25886,N_24832,N_24188);
nor U25887 (N_25887,N_24236,N_24052);
and U25888 (N_25888,N_24561,N_24931);
nand U25889 (N_25889,N_24097,N_24041);
nand U25890 (N_25890,N_24565,N_24334);
or U25891 (N_25891,N_24876,N_24302);
nor U25892 (N_25892,N_24494,N_24566);
nand U25893 (N_25893,N_24640,N_24284);
xnor U25894 (N_25894,N_24308,N_24806);
xnor U25895 (N_25895,N_24044,N_24780);
and U25896 (N_25896,N_24875,N_24003);
or U25897 (N_25897,N_24176,N_24416);
and U25898 (N_25898,N_24475,N_24349);
or U25899 (N_25899,N_24496,N_24272);
nand U25900 (N_25900,N_24966,N_24999);
nand U25901 (N_25901,N_24308,N_24041);
or U25902 (N_25902,N_24856,N_24692);
nand U25903 (N_25903,N_24429,N_24593);
and U25904 (N_25904,N_24991,N_24764);
or U25905 (N_25905,N_24528,N_24697);
nand U25906 (N_25906,N_24117,N_24144);
nor U25907 (N_25907,N_24469,N_24928);
and U25908 (N_25908,N_24081,N_24355);
or U25909 (N_25909,N_24699,N_24164);
nor U25910 (N_25910,N_24467,N_24714);
nand U25911 (N_25911,N_24341,N_24261);
nor U25912 (N_25912,N_24217,N_24557);
nand U25913 (N_25913,N_24413,N_24946);
xor U25914 (N_25914,N_24144,N_24942);
nand U25915 (N_25915,N_24585,N_24694);
xnor U25916 (N_25916,N_24381,N_24017);
nor U25917 (N_25917,N_24985,N_24452);
nand U25918 (N_25918,N_24356,N_24827);
nor U25919 (N_25919,N_24170,N_24275);
xnor U25920 (N_25920,N_24801,N_24205);
or U25921 (N_25921,N_24981,N_24130);
and U25922 (N_25922,N_24114,N_24054);
nor U25923 (N_25923,N_24547,N_24389);
or U25924 (N_25924,N_24558,N_24503);
nor U25925 (N_25925,N_24184,N_24448);
nor U25926 (N_25926,N_24863,N_24039);
nand U25927 (N_25927,N_24674,N_24836);
or U25928 (N_25928,N_24365,N_24702);
and U25929 (N_25929,N_24629,N_24921);
and U25930 (N_25930,N_24289,N_24749);
nor U25931 (N_25931,N_24917,N_24982);
xnor U25932 (N_25932,N_24928,N_24504);
nor U25933 (N_25933,N_24124,N_24283);
or U25934 (N_25934,N_24816,N_24073);
xnor U25935 (N_25935,N_24161,N_24254);
xor U25936 (N_25936,N_24689,N_24180);
and U25937 (N_25937,N_24893,N_24171);
or U25938 (N_25938,N_24967,N_24472);
and U25939 (N_25939,N_24692,N_24672);
nand U25940 (N_25940,N_24510,N_24685);
xor U25941 (N_25941,N_24266,N_24718);
and U25942 (N_25942,N_24385,N_24765);
or U25943 (N_25943,N_24280,N_24749);
nor U25944 (N_25944,N_24231,N_24798);
nor U25945 (N_25945,N_24763,N_24274);
or U25946 (N_25946,N_24813,N_24607);
xor U25947 (N_25947,N_24555,N_24477);
nand U25948 (N_25948,N_24564,N_24281);
nor U25949 (N_25949,N_24648,N_24195);
nand U25950 (N_25950,N_24049,N_24423);
nand U25951 (N_25951,N_24509,N_24585);
nand U25952 (N_25952,N_24230,N_24925);
nor U25953 (N_25953,N_24302,N_24943);
nand U25954 (N_25954,N_24281,N_24955);
xnor U25955 (N_25955,N_24189,N_24509);
nand U25956 (N_25956,N_24050,N_24813);
xnor U25957 (N_25957,N_24148,N_24120);
or U25958 (N_25958,N_24891,N_24907);
xor U25959 (N_25959,N_24906,N_24109);
nand U25960 (N_25960,N_24074,N_24937);
or U25961 (N_25961,N_24722,N_24118);
xnor U25962 (N_25962,N_24411,N_24007);
nor U25963 (N_25963,N_24332,N_24669);
and U25964 (N_25964,N_24757,N_24116);
or U25965 (N_25965,N_24817,N_24924);
xnor U25966 (N_25966,N_24561,N_24300);
nor U25967 (N_25967,N_24676,N_24607);
and U25968 (N_25968,N_24009,N_24898);
xor U25969 (N_25969,N_24468,N_24225);
nand U25970 (N_25970,N_24005,N_24819);
xor U25971 (N_25971,N_24004,N_24322);
xor U25972 (N_25972,N_24081,N_24800);
nor U25973 (N_25973,N_24565,N_24969);
and U25974 (N_25974,N_24262,N_24244);
nand U25975 (N_25975,N_24088,N_24512);
xor U25976 (N_25976,N_24681,N_24829);
and U25977 (N_25977,N_24550,N_24519);
and U25978 (N_25978,N_24460,N_24788);
or U25979 (N_25979,N_24846,N_24225);
xor U25980 (N_25980,N_24982,N_24198);
xor U25981 (N_25981,N_24284,N_24144);
nor U25982 (N_25982,N_24025,N_24654);
xnor U25983 (N_25983,N_24487,N_24882);
nand U25984 (N_25984,N_24969,N_24439);
xnor U25985 (N_25985,N_24371,N_24444);
nand U25986 (N_25986,N_24402,N_24791);
xnor U25987 (N_25987,N_24400,N_24010);
nor U25988 (N_25988,N_24734,N_24206);
or U25989 (N_25989,N_24592,N_24986);
and U25990 (N_25990,N_24543,N_24415);
nand U25991 (N_25991,N_24571,N_24420);
and U25992 (N_25992,N_24813,N_24443);
xor U25993 (N_25993,N_24964,N_24268);
nor U25994 (N_25994,N_24856,N_24744);
and U25995 (N_25995,N_24179,N_24448);
nor U25996 (N_25996,N_24270,N_24954);
or U25997 (N_25997,N_24546,N_24716);
or U25998 (N_25998,N_24678,N_24816);
or U25999 (N_25999,N_24718,N_24407);
and U26000 (N_26000,N_25487,N_25877);
and U26001 (N_26001,N_25394,N_25233);
or U26002 (N_26002,N_25020,N_25288);
nor U26003 (N_26003,N_25389,N_25718);
xnor U26004 (N_26004,N_25384,N_25728);
nor U26005 (N_26005,N_25403,N_25033);
nand U26006 (N_26006,N_25558,N_25580);
nor U26007 (N_26007,N_25362,N_25939);
nor U26008 (N_26008,N_25331,N_25002);
and U26009 (N_26009,N_25620,N_25097);
nor U26010 (N_26010,N_25643,N_25459);
nand U26011 (N_26011,N_25817,N_25099);
and U26012 (N_26012,N_25985,N_25875);
and U26013 (N_26013,N_25352,N_25215);
and U26014 (N_26014,N_25096,N_25696);
or U26015 (N_26015,N_25294,N_25552);
nor U26016 (N_26016,N_25010,N_25964);
xor U26017 (N_26017,N_25351,N_25053);
and U26018 (N_26018,N_25113,N_25779);
nand U26019 (N_26019,N_25130,N_25955);
and U26020 (N_26020,N_25810,N_25448);
nand U26021 (N_26021,N_25514,N_25619);
nand U26022 (N_26022,N_25324,N_25885);
nor U26023 (N_26023,N_25135,N_25292);
and U26024 (N_26024,N_25952,N_25686);
nand U26025 (N_26025,N_25189,N_25860);
nand U26026 (N_26026,N_25128,N_25409);
or U26027 (N_26027,N_25105,N_25769);
nand U26028 (N_26028,N_25585,N_25417);
or U26029 (N_26029,N_25123,N_25469);
xnor U26030 (N_26030,N_25782,N_25344);
and U26031 (N_26031,N_25594,N_25063);
or U26032 (N_26032,N_25757,N_25239);
or U26033 (N_26033,N_25383,N_25311);
nand U26034 (N_26034,N_25687,N_25562);
and U26035 (N_26035,N_25160,N_25768);
or U26036 (N_26036,N_25517,N_25214);
xnor U26037 (N_26037,N_25369,N_25829);
xnor U26038 (N_26038,N_25826,N_25240);
and U26039 (N_26039,N_25200,N_25715);
nand U26040 (N_26040,N_25533,N_25906);
or U26041 (N_26041,N_25849,N_25868);
xnor U26042 (N_26042,N_25152,N_25059);
nor U26043 (N_26043,N_25651,N_25887);
nand U26044 (N_26044,N_25248,N_25554);
nand U26045 (N_26045,N_25088,N_25881);
nand U26046 (N_26046,N_25227,N_25583);
and U26047 (N_26047,N_25929,N_25336);
xnor U26048 (N_26048,N_25853,N_25867);
nor U26049 (N_26049,N_25541,N_25077);
nor U26050 (N_26050,N_25539,N_25150);
and U26051 (N_26051,N_25157,N_25988);
or U26052 (N_26052,N_25951,N_25682);
nor U26053 (N_26053,N_25180,N_25064);
nor U26054 (N_26054,N_25028,N_25357);
nor U26055 (N_26055,N_25425,N_25984);
xor U26056 (N_26056,N_25366,N_25264);
nor U26057 (N_26057,N_25149,N_25634);
or U26058 (N_26058,N_25041,N_25355);
or U26059 (N_26059,N_25298,N_25285);
nor U26060 (N_26060,N_25522,N_25304);
nand U26061 (N_26061,N_25612,N_25804);
xnor U26062 (N_26062,N_25386,N_25124);
nand U26063 (N_26063,N_25801,N_25173);
or U26064 (N_26064,N_25636,N_25231);
and U26065 (N_26065,N_25252,N_25865);
xor U26066 (N_26066,N_25121,N_25778);
nand U26067 (N_26067,N_25183,N_25969);
nand U26068 (N_26068,N_25812,N_25884);
xor U26069 (N_26069,N_25091,N_25481);
xnor U26070 (N_26070,N_25205,N_25914);
xnor U26071 (N_26071,N_25843,N_25850);
xnor U26072 (N_26072,N_25491,N_25246);
and U26073 (N_26073,N_25134,N_25996);
and U26074 (N_26074,N_25106,N_25748);
or U26075 (N_26075,N_25960,N_25238);
or U26076 (N_26076,N_25716,N_25673);
and U26077 (N_26077,N_25893,N_25090);
and U26078 (N_26078,N_25861,N_25464);
xnor U26079 (N_26079,N_25726,N_25460);
nor U26080 (N_26080,N_25838,N_25485);
nor U26081 (N_26081,N_25661,N_25856);
nor U26082 (N_26082,N_25222,N_25212);
and U26083 (N_26083,N_25642,N_25334);
xor U26084 (N_26084,N_25949,N_25257);
nand U26085 (N_26085,N_25669,N_25831);
and U26086 (N_26086,N_25618,N_25100);
and U26087 (N_26087,N_25819,N_25026);
nand U26088 (N_26088,N_25519,N_25511);
or U26089 (N_26089,N_25821,N_25407);
or U26090 (N_26090,N_25596,N_25019);
nand U26091 (N_26091,N_25083,N_25874);
xor U26092 (N_26092,N_25229,N_25547);
xnor U26093 (N_26093,N_25065,N_25270);
nor U26094 (N_26094,N_25493,N_25315);
and U26095 (N_26095,N_25319,N_25422);
nor U26096 (N_26096,N_25808,N_25740);
xnor U26097 (N_26097,N_25540,N_25898);
or U26098 (N_26098,N_25567,N_25080);
nor U26099 (N_26099,N_25873,N_25910);
nor U26100 (N_26100,N_25404,N_25937);
or U26101 (N_26101,N_25889,N_25604);
or U26102 (N_26102,N_25704,N_25746);
nand U26103 (N_26103,N_25926,N_25220);
or U26104 (N_26104,N_25377,N_25922);
or U26105 (N_26105,N_25117,N_25833);
nor U26106 (N_26106,N_25684,N_25842);
and U26107 (N_26107,N_25273,N_25378);
nor U26108 (N_26108,N_25530,N_25958);
xnor U26109 (N_26109,N_25442,N_25198);
xor U26110 (N_26110,N_25265,N_25145);
and U26111 (N_26111,N_25609,N_25399);
or U26112 (N_26112,N_25859,N_25216);
and U26113 (N_26113,N_25745,N_25249);
nand U26114 (N_26114,N_25471,N_25784);
and U26115 (N_26115,N_25155,N_25532);
xor U26116 (N_26116,N_25392,N_25272);
nor U26117 (N_26117,N_25602,N_25296);
and U26118 (N_26118,N_25089,N_25470);
and U26119 (N_26119,N_25341,N_25744);
nand U26120 (N_26120,N_25133,N_25866);
or U26121 (N_26121,N_25597,N_25503);
nand U26122 (N_26122,N_25360,N_25714);
xor U26123 (N_26123,N_25045,N_25649);
and U26124 (N_26124,N_25590,N_25423);
or U26125 (N_26125,N_25158,N_25827);
nor U26126 (N_26126,N_25933,N_25453);
or U26127 (N_26127,N_25251,N_25032);
and U26128 (N_26128,N_25375,N_25553);
or U26129 (N_26129,N_25162,N_25250);
nand U26130 (N_26130,N_25489,N_25892);
or U26131 (N_26131,N_25975,N_25830);
and U26132 (N_26132,N_25650,N_25538);
or U26133 (N_26133,N_25259,N_25452);
xor U26134 (N_26134,N_25862,N_25398);
and U26135 (N_26135,N_25616,N_25524);
xnor U26136 (N_26136,N_25879,N_25261);
nand U26137 (N_26137,N_25919,N_25428);
nor U26138 (N_26138,N_25593,N_25199);
xor U26139 (N_26139,N_25756,N_25408);
and U26140 (N_26140,N_25084,N_25675);
or U26141 (N_26141,N_25700,N_25773);
nor U26142 (N_26142,N_25112,N_25668);
nand U26143 (N_26143,N_25185,N_25092);
nand U26144 (N_26144,N_25380,N_25043);
nor U26145 (N_26145,N_25947,N_25531);
nand U26146 (N_26146,N_25815,N_25201);
nand U26147 (N_26147,N_25974,N_25681);
nor U26148 (N_26148,N_25477,N_25005);
or U26149 (N_26149,N_25094,N_25510);
or U26150 (N_26150,N_25965,N_25181);
and U26151 (N_26151,N_25820,N_25348);
xor U26152 (N_26152,N_25320,N_25750);
or U26153 (N_26153,N_25165,N_25052);
or U26154 (N_26154,N_25241,N_25391);
nand U26155 (N_26155,N_25855,N_25465);
nand U26156 (N_26156,N_25775,N_25709);
and U26157 (N_26157,N_25247,N_25372);
and U26158 (N_26158,N_25980,N_25601);
or U26159 (N_26159,N_25662,N_25701);
xor U26160 (N_26160,N_25115,N_25412);
xnor U26161 (N_26161,N_25328,N_25839);
nand U26162 (N_26162,N_25101,N_25577);
or U26163 (N_26163,N_25116,N_25466);
or U26164 (N_26164,N_25844,N_25799);
nand U26165 (N_26165,N_25835,N_25427);
xor U26166 (N_26166,N_25840,N_25790);
nand U26167 (N_26167,N_25615,N_25076);
and U26168 (N_26168,N_25488,N_25174);
or U26169 (N_26169,N_25918,N_25667);
and U26170 (N_26170,N_25513,N_25291);
nor U26171 (N_26171,N_25792,N_25689);
and U26172 (N_26172,N_25708,N_25195);
nand U26173 (N_26173,N_25379,N_25140);
nor U26174 (N_26174,N_25724,N_25103);
xor U26175 (N_26175,N_25752,N_25795);
nand U26176 (N_26176,N_25204,N_25758);
nor U26177 (N_26177,N_25573,N_25747);
or U26178 (N_26178,N_25230,N_25258);
and U26179 (N_26179,N_25764,N_25434);
xnor U26180 (N_26180,N_25303,N_25605);
or U26181 (N_26181,N_25433,N_25314);
and U26182 (N_26182,N_25930,N_25104);
and U26183 (N_26183,N_25382,N_25641);
xnor U26184 (N_26184,N_25279,N_25610);
nor U26185 (N_26185,N_25169,N_25313);
and U26186 (N_26186,N_25542,N_25927);
nand U26187 (N_26187,N_25447,N_25571);
and U26188 (N_26188,N_25537,N_25712);
xor U26189 (N_26189,N_25278,N_25621);
or U26190 (N_26190,N_25299,N_25413);
xor U26191 (N_26191,N_25339,N_25301);
nand U26192 (N_26192,N_25535,N_25648);
nand U26193 (N_26193,N_25907,N_25353);
xnor U26194 (N_26194,N_25986,N_25586);
or U26195 (N_26195,N_25559,N_25347);
nor U26196 (N_26196,N_25038,N_25759);
nand U26197 (N_26197,N_25056,N_25013);
or U26198 (N_26198,N_25373,N_25006);
xnor U26199 (N_26199,N_25846,N_25042);
and U26200 (N_26200,N_25994,N_25617);
and U26201 (N_26201,N_25972,N_25441);
or U26202 (N_26202,N_25191,N_25961);
or U26203 (N_26203,N_25289,N_25003);
xor U26204 (N_26204,N_25046,N_25405);
or U26205 (N_26205,N_25307,N_25455);
nor U26206 (N_26206,N_25979,N_25168);
and U26207 (N_26207,N_25126,N_25638);
nand U26208 (N_26208,N_25945,N_25589);
and U26209 (N_26209,N_25400,N_25934);
nor U26210 (N_26210,N_25818,N_25713);
and U26211 (N_26211,N_25946,N_25735);
or U26212 (N_26212,N_25060,N_25376);
or U26213 (N_26213,N_25526,N_25731);
xnor U26214 (N_26214,N_25219,N_25302);
xor U26215 (N_26215,N_25897,N_25645);
and U26216 (N_26216,N_25807,N_25802);
or U26217 (N_26217,N_25236,N_25991);
xor U26218 (N_26218,N_25880,N_25623);
nor U26219 (N_26219,N_25011,N_25190);
nand U26220 (N_26220,N_25385,N_25223);
nand U26221 (N_26221,N_25823,N_25450);
xnor U26222 (N_26222,N_25282,N_25057);
or U26223 (N_26223,N_25439,N_25139);
xor U26224 (N_26224,N_25674,N_25624);
nand U26225 (N_26225,N_25864,N_25549);
nand U26226 (N_26226,N_25837,N_25658);
and U26227 (N_26227,N_25388,N_25345);
and U26228 (N_26228,N_25119,N_25039);
nand U26229 (N_26229,N_25938,N_25652);
xnor U26230 (N_26230,N_25508,N_25018);
and U26231 (N_26231,N_25654,N_25671);
nor U26232 (N_26232,N_25297,N_25626);
and U26233 (N_26233,N_25131,N_25534);
or U26234 (N_26234,N_25141,N_25111);
and U26235 (N_26235,N_25677,N_25941);
or U26236 (N_26236,N_25401,N_25909);
nor U26237 (N_26237,N_25560,N_25209);
nand U26238 (N_26238,N_25579,N_25086);
or U26239 (N_26239,N_25551,N_25723);
and U26240 (N_26240,N_25688,N_25040);
xor U26241 (N_26241,N_25848,N_25482);
or U26242 (N_26242,N_25664,N_25698);
nor U26243 (N_26243,N_25473,N_25081);
xnor U26244 (N_26244,N_25911,N_25243);
or U26245 (N_26245,N_25281,N_25415);
or U26246 (N_26246,N_25772,N_25736);
and U26247 (N_26247,N_25672,N_25857);
or U26248 (N_26248,N_25515,N_25340);
xor U26249 (N_26249,N_25523,N_25587);
nand U26250 (N_26250,N_25520,N_25614);
or U26251 (N_26251,N_25406,N_25806);
and U26252 (N_26252,N_25738,N_25431);
xor U26253 (N_26253,N_25613,N_25147);
nor U26254 (N_26254,N_25498,N_25411);
nand U26255 (N_26255,N_25899,N_25557);
nand U26256 (N_26256,N_25923,N_25824);
nor U26257 (N_26257,N_25275,N_25068);
or U26258 (N_26258,N_25071,N_25981);
xor U26259 (N_26259,N_25765,N_25263);
or U26260 (N_26260,N_25916,N_25727);
and U26261 (N_26261,N_25917,N_25721);
and U26262 (N_26262,N_25931,N_25395);
or U26263 (N_26263,N_25500,N_25670);
or U26264 (N_26264,N_25639,N_25729);
and U26265 (N_26265,N_25496,N_25963);
xnor U26266 (N_26266,N_25635,N_25114);
and U26267 (N_26267,N_25228,N_25568);
and U26268 (N_26268,N_25543,N_25317);
xor U26269 (N_26269,N_25102,N_25581);
xor U26270 (N_26270,N_25970,N_25734);
nor U26271 (N_26271,N_25211,N_25333);
and U26272 (N_26272,N_25420,N_25170);
xnor U26273 (N_26273,N_25027,N_25332);
nand U26274 (N_26274,N_25108,N_25913);
nor U26275 (N_26275,N_25015,N_25628);
nor U26276 (N_26276,N_25944,N_25936);
nand U26277 (N_26277,N_25753,N_25786);
and U26278 (N_26278,N_25599,N_25956);
nor U26279 (N_26279,N_25679,N_25749);
xor U26280 (N_26280,N_25982,N_25739);
or U26281 (N_26281,N_25416,N_25107);
nor U26282 (N_26282,N_25995,N_25680);
or U26283 (N_26283,N_25132,N_25825);
nand U26284 (N_26284,N_25274,N_25009);
nand U26285 (N_26285,N_25284,N_25863);
and U26286 (N_26286,N_25188,N_25572);
nor U26287 (N_26287,N_25225,N_25025);
nor U26288 (N_26288,N_25777,N_25050);
xor U26289 (N_26289,N_25262,N_25555);
nor U26290 (N_26290,N_25235,N_25359);
nor U26291 (N_26291,N_25763,N_25280);
nor U26292 (N_26292,N_25021,N_25767);
xnor U26293 (N_26293,N_25475,N_25047);
or U26294 (N_26294,N_25566,N_25467);
or U26295 (N_26295,N_25563,N_25418);
and U26296 (N_26296,N_25363,N_25479);
xnor U26297 (N_26297,N_25544,N_25507);
nand U26298 (N_26298,N_25494,N_25891);
or U26299 (N_26299,N_25210,N_25125);
or U26300 (N_26300,N_25182,N_25954);
xor U26301 (N_26301,N_25998,N_25022);
xor U26302 (N_26302,N_25521,N_25276);
or U26303 (N_26303,N_25966,N_25267);
nor U26304 (N_26304,N_25213,N_25354);
and U26305 (N_26305,N_25871,N_25244);
or U26306 (N_26306,N_25999,N_25136);
nand U26307 (N_26307,N_25224,N_25424);
nor U26308 (N_26308,N_25561,N_25660);
xor U26309 (N_26309,N_25129,N_25781);
nand U26310 (N_26310,N_25869,N_25603);
xnor U26311 (N_26311,N_25148,N_25813);
nor U26312 (N_26312,N_25754,N_25226);
or U26313 (N_26313,N_25836,N_25968);
nand U26314 (N_26314,N_25785,N_25574);
nor U26315 (N_26315,N_25940,N_25527);
xor U26316 (N_26316,N_25419,N_25069);
nor U26317 (N_26317,N_25446,N_25054);
and U26318 (N_26318,N_25600,N_25548);
or U26319 (N_26319,N_25255,N_25845);
and U26320 (N_26320,N_25156,N_25034);
nand U26321 (N_26321,N_25512,N_25122);
or U26322 (N_26322,N_25942,N_25607);
and U26323 (N_26323,N_25458,N_25588);
nand U26324 (N_26324,N_25184,N_25269);
nor U26325 (N_26325,N_25364,N_25691);
and U26326 (N_26326,N_25449,N_25499);
nand U26327 (N_26327,N_25789,N_25166);
and U26328 (N_26328,N_25087,N_25797);
nand U26329 (N_26329,N_25438,N_25206);
xor U26330 (N_26330,N_25948,N_25349);
nor U26331 (N_26331,N_25565,N_25073);
xor U26332 (N_26332,N_25343,N_25232);
xnor U26333 (N_26333,N_25254,N_25397);
nor U26334 (N_26334,N_25787,N_25920);
nand U26335 (N_26335,N_25742,N_25720);
xnor U26336 (N_26336,N_25928,N_25900);
nand U26337 (N_26337,N_25330,N_25692);
nor U26338 (N_26338,N_25525,N_25242);
nor U26339 (N_26339,N_25075,N_25962);
and U26340 (N_26340,N_25161,N_25751);
or U26341 (N_26341,N_25367,N_25029);
or U26342 (N_26342,N_25598,N_25851);
nand U26343 (N_26343,N_25082,N_25872);
xor U26344 (N_26344,N_25575,N_25683);
nand U26345 (N_26345,N_25656,N_25396);
and U26346 (N_26346,N_25582,N_25444);
and U26347 (N_26347,N_25770,N_25888);
and U26348 (N_26348,N_25461,N_25932);
and U26349 (N_26349,N_25402,N_25834);
or U26350 (N_26350,N_25822,N_25159);
or U26351 (N_26351,N_25072,N_25295);
nor U26352 (N_26352,N_25591,N_25556);
nor U26353 (N_26353,N_25705,N_25172);
xnor U26354 (N_26354,N_25627,N_25058);
nand U26355 (N_26355,N_25305,N_25031);
nand U26356 (N_26356,N_25640,N_25067);
xor U26357 (N_26357,N_25545,N_25177);
xor U26358 (N_26358,N_25847,N_25832);
nor U26359 (N_26359,N_25480,N_25437);
nand U26360 (N_26360,N_25316,N_25653);
xor U26361 (N_26361,N_25908,N_25506);
nand U26362 (N_26362,N_25245,N_25894);
or U26363 (N_26363,N_25192,N_25287);
xor U26364 (N_26364,N_25576,N_25771);
xor U26365 (N_26365,N_25760,N_25904);
nor U26366 (N_26366,N_25761,N_25741);
and U26367 (N_26367,N_25608,N_25632);
xnor U26368 (N_26368,N_25693,N_25987);
nor U26369 (N_26369,N_25633,N_25007);
nand U26370 (N_26370,N_25967,N_25393);
nand U26371 (N_26371,N_25138,N_25803);
or U26372 (N_26372,N_25120,N_25990);
nor U26373 (N_26373,N_25895,N_25078);
nor U26374 (N_26374,N_25361,N_25203);
nor U26375 (N_26375,N_25666,N_25997);
or U26376 (N_26376,N_25992,N_25474);
xor U26377 (N_26377,N_25044,N_25008);
nand U26378 (N_26378,N_25410,N_25497);
and U26379 (N_26379,N_25085,N_25690);
xnor U26380 (N_26380,N_25783,N_25171);
nand U26381 (N_26381,N_25048,N_25983);
xnor U26382 (N_26382,N_25049,N_25164);
and U26383 (N_26383,N_25268,N_25733);
xnor U26384 (N_26384,N_25127,N_25989);
and U26385 (N_26385,N_25504,N_25959);
or U26386 (N_26386,N_25536,N_25828);
and U26387 (N_26387,N_25098,N_25023);
nor U26388 (N_26388,N_25426,N_25901);
or U26389 (N_26389,N_25374,N_25017);
and U26390 (N_26390,N_25358,N_25793);
nor U26391 (N_26391,N_25971,N_25143);
or U26392 (N_26392,N_25186,N_25208);
or U26393 (N_26393,N_25809,N_25478);
nor U26394 (N_26394,N_25154,N_25501);
xor U26395 (N_26395,N_25655,N_25676);
nand U26396 (N_26396,N_25516,N_25338);
xor U26397 (N_26397,N_25611,N_25454);
or U26398 (N_26398,N_25310,N_25657);
or U26399 (N_26399,N_25055,N_25776);
and U26400 (N_26400,N_25569,N_25915);
nand U26401 (N_26401,N_25732,N_25953);
xnor U26402 (N_26402,N_25462,N_25665);
nor U26403 (N_26403,N_25957,N_25429);
xnor U26404 (N_26404,N_25528,N_25518);
xnor U26405 (N_26405,N_25001,N_25421);
xor U26406 (N_26406,N_25993,N_25074);
and U26407 (N_26407,N_25346,N_25695);
or U26408 (N_26408,N_25630,N_25312);
or U26409 (N_26409,N_25490,N_25432);
and U26410 (N_26410,N_25890,N_25719);
nor U26411 (N_26411,N_25014,N_25622);
or U26412 (N_26412,N_25791,N_25024);
nand U26413 (N_26413,N_25277,N_25584);
or U26414 (N_26414,N_25925,N_25800);
or U26415 (N_26415,N_25436,N_25365);
or U26416 (N_26416,N_25631,N_25706);
nand U26417 (N_26417,N_25794,N_25202);
xor U26418 (N_26418,N_25703,N_25841);
nand U26419 (N_26419,N_25854,N_25435);
xor U26420 (N_26420,N_25722,N_25509);
xor U26421 (N_26421,N_25012,N_25144);
or U26422 (N_26422,N_25000,N_25730);
nand U26423 (N_26423,N_25179,N_25387);
or U26424 (N_26424,N_25702,N_25175);
or U26425 (N_26425,N_25858,N_25973);
nor U26426 (N_26426,N_25318,N_25896);
nand U26427 (N_26427,N_25079,N_25659);
nand U26428 (N_26428,N_25167,N_25443);
nand U26429 (N_26429,N_25327,N_25300);
or U26430 (N_26430,N_25286,N_25271);
or U26431 (N_26431,N_25468,N_25711);
xor U26432 (N_26432,N_25325,N_25350);
nand U26433 (N_26433,N_25570,N_25876);
nor U26434 (N_26434,N_25004,N_25606);
xnor U26435 (N_26435,N_25902,N_25356);
and U26436 (N_26436,N_25253,N_25737);
xnor U26437 (N_26437,N_25326,N_25066);
nor U26438 (N_26438,N_25492,N_25146);
or U26439 (N_26439,N_25805,N_25814);
and U26440 (N_26440,N_25451,N_25629);
or U26441 (N_26441,N_25811,N_25051);
nand U26442 (N_26442,N_25323,N_25153);
nor U26443 (N_26443,N_25882,N_25935);
xor U26444 (N_26444,N_25070,N_25883);
and U26445 (N_26445,N_25912,N_25109);
nor U26446 (N_26446,N_25976,N_25260);
nor U26447 (N_26447,N_25197,N_25062);
or U26448 (N_26448,N_25370,N_25163);
nor U26449 (N_26449,N_25256,N_25430);
or U26450 (N_26450,N_25550,N_25592);
nor U26451 (N_26451,N_25371,N_25266);
xor U26452 (N_26452,N_25564,N_25762);
xnor U26453 (N_26453,N_25694,N_25234);
nand U26454 (N_26454,N_25194,N_25093);
nor U26455 (N_26455,N_25546,N_25440);
and U26456 (N_26456,N_25176,N_25870);
or U26457 (N_26457,N_25414,N_25697);
nor U26458 (N_26458,N_25816,N_25486);
or U26459 (N_26459,N_25774,N_25886);
or U26460 (N_26460,N_25193,N_25529);
and U26461 (N_26461,N_25725,N_25381);
and U26462 (N_26462,N_25788,N_25678);
and U26463 (N_26463,N_25036,N_25625);
xor U26464 (N_26464,N_25780,N_25943);
nand U26465 (N_26465,N_25037,N_25142);
or U26466 (N_26466,N_25187,N_25978);
xnor U26467 (N_26467,N_25878,N_25921);
and U26468 (N_26468,N_25306,N_25637);
xor U26469 (N_26469,N_25217,N_25322);
xnor U26470 (N_26470,N_25924,N_25337);
nand U26471 (N_26471,N_25293,N_25110);
xnor U26472 (N_26472,N_25321,N_25644);
nand U26473 (N_26473,N_25905,N_25342);
or U26474 (N_26474,N_25237,N_25743);
nor U26475 (N_26475,N_25118,N_25309);
nor U26476 (N_26476,N_25977,N_25095);
or U26477 (N_26477,N_25456,N_25852);
or U26478 (N_26478,N_25218,N_25647);
nor U26479 (N_26479,N_25151,N_25196);
nor U26480 (N_26480,N_25329,N_25283);
nor U26481 (N_26481,N_25798,N_25710);
xor U26482 (N_26482,N_25335,N_25035);
and U26483 (N_26483,N_25950,N_25502);
xor U26484 (N_26484,N_25472,N_25207);
nor U26485 (N_26485,N_25476,N_25445);
and U26486 (N_26486,N_25903,N_25796);
xnor U26487 (N_26487,N_25221,N_25505);
xor U26488 (N_26488,N_25016,N_25483);
xor U26489 (N_26489,N_25368,N_25457);
nor U26490 (N_26490,N_25030,N_25178);
nor U26491 (N_26491,N_25390,N_25463);
nor U26492 (N_26492,N_25766,N_25707);
nand U26493 (N_26493,N_25308,N_25755);
and U26494 (N_26494,N_25290,N_25495);
nand U26495 (N_26495,N_25663,N_25717);
nand U26496 (N_26496,N_25699,N_25061);
or U26497 (N_26497,N_25484,N_25137);
xnor U26498 (N_26498,N_25685,N_25578);
or U26499 (N_26499,N_25646,N_25595);
nand U26500 (N_26500,N_25314,N_25108);
xor U26501 (N_26501,N_25882,N_25961);
nor U26502 (N_26502,N_25384,N_25161);
or U26503 (N_26503,N_25850,N_25678);
nand U26504 (N_26504,N_25018,N_25493);
nand U26505 (N_26505,N_25109,N_25627);
and U26506 (N_26506,N_25561,N_25825);
nand U26507 (N_26507,N_25514,N_25284);
and U26508 (N_26508,N_25823,N_25433);
or U26509 (N_26509,N_25407,N_25058);
or U26510 (N_26510,N_25580,N_25919);
and U26511 (N_26511,N_25802,N_25917);
nor U26512 (N_26512,N_25086,N_25134);
or U26513 (N_26513,N_25928,N_25585);
nand U26514 (N_26514,N_25276,N_25381);
or U26515 (N_26515,N_25528,N_25989);
nand U26516 (N_26516,N_25205,N_25588);
or U26517 (N_26517,N_25012,N_25820);
nand U26518 (N_26518,N_25310,N_25031);
nor U26519 (N_26519,N_25252,N_25992);
xor U26520 (N_26520,N_25416,N_25459);
xnor U26521 (N_26521,N_25006,N_25545);
and U26522 (N_26522,N_25615,N_25704);
or U26523 (N_26523,N_25839,N_25188);
nor U26524 (N_26524,N_25193,N_25437);
xor U26525 (N_26525,N_25244,N_25172);
nor U26526 (N_26526,N_25701,N_25782);
xor U26527 (N_26527,N_25079,N_25247);
xor U26528 (N_26528,N_25120,N_25959);
and U26529 (N_26529,N_25533,N_25977);
xor U26530 (N_26530,N_25244,N_25366);
or U26531 (N_26531,N_25572,N_25731);
and U26532 (N_26532,N_25035,N_25153);
and U26533 (N_26533,N_25369,N_25900);
and U26534 (N_26534,N_25564,N_25012);
xnor U26535 (N_26535,N_25512,N_25867);
nor U26536 (N_26536,N_25030,N_25541);
and U26537 (N_26537,N_25580,N_25384);
and U26538 (N_26538,N_25103,N_25320);
or U26539 (N_26539,N_25852,N_25873);
xor U26540 (N_26540,N_25565,N_25482);
or U26541 (N_26541,N_25087,N_25990);
or U26542 (N_26542,N_25631,N_25803);
nor U26543 (N_26543,N_25557,N_25346);
xor U26544 (N_26544,N_25835,N_25557);
nand U26545 (N_26545,N_25093,N_25649);
nand U26546 (N_26546,N_25000,N_25038);
and U26547 (N_26547,N_25683,N_25694);
or U26548 (N_26548,N_25090,N_25030);
xnor U26549 (N_26549,N_25678,N_25885);
xor U26550 (N_26550,N_25610,N_25997);
nor U26551 (N_26551,N_25227,N_25831);
and U26552 (N_26552,N_25334,N_25980);
nor U26553 (N_26553,N_25051,N_25302);
nand U26554 (N_26554,N_25520,N_25765);
nor U26555 (N_26555,N_25137,N_25122);
xor U26556 (N_26556,N_25651,N_25234);
or U26557 (N_26557,N_25292,N_25257);
xnor U26558 (N_26558,N_25905,N_25218);
xnor U26559 (N_26559,N_25509,N_25587);
xor U26560 (N_26560,N_25088,N_25424);
xor U26561 (N_26561,N_25630,N_25616);
or U26562 (N_26562,N_25252,N_25294);
or U26563 (N_26563,N_25441,N_25198);
nor U26564 (N_26564,N_25778,N_25095);
and U26565 (N_26565,N_25192,N_25450);
nor U26566 (N_26566,N_25734,N_25655);
nor U26567 (N_26567,N_25265,N_25890);
xnor U26568 (N_26568,N_25118,N_25881);
and U26569 (N_26569,N_25378,N_25770);
and U26570 (N_26570,N_25573,N_25183);
nand U26571 (N_26571,N_25218,N_25082);
nand U26572 (N_26572,N_25332,N_25031);
and U26573 (N_26573,N_25913,N_25529);
and U26574 (N_26574,N_25120,N_25279);
xnor U26575 (N_26575,N_25038,N_25594);
nor U26576 (N_26576,N_25310,N_25439);
nand U26577 (N_26577,N_25252,N_25325);
and U26578 (N_26578,N_25182,N_25030);
and U26579 (N_26579,N_25321,N_25855);
and U26580 (N_26580,N_25674,N_25669);
nand U26581 (N_26581,N_25199,N_25721);
nor U26582 (N_26582,N_25524,N_25719);
or U26583 (N_26583,N_25766,N_25792);
nor U26584 (N_26584,N_25010,N_25998);
xnor U26585 (N_26585,N_25772,N_25717);
xor U26586 (N_26586,N_25068,N_25463);
xnor U26587 (N_26587,N_25675,N_25842);
xnor U26588 (N_26588,N_25350,N_25717);
xnor U26589 (N_26589,N_25231,N_25673);
xor U26590 (N_26590,N_25847,N_25670);
nand U26591 (N_26591,N_25004,N_25150);
or U26592 (N_26592,N_25678,N_25642);
xor U26593 (N_26593,N_25063,N_25753);
nand U26594 (N_26594,N_25134,N_25610);
xnor U26595 (N_26595,N_25685,N_25658);
nor U26596 (N_26596,N_25605,N_25587);
or U26597 (N_26597,N_25749,N_25991);
or U26598 (N_26598,N_25427,N_25853);
or U26599 (N_26599,N_25508,N_25394);
or U26600 (N_26600,N_25756,N_25946);
and U26601 (N_26601,N_25690,N_25923);
nand U26602 (N_26602,N_25545,N_25990);
nand U26603 (N_26603,N_25043,N_25339);
xnor U26604 (N_26604,N_25057,N_25176);
nand U26605 (N_26605,N_25106,N_25338);
nand U26606 (N_26606,N_25468,N_25527);
nand U26607 (N_26607,N_25268,N_25108);
nor U26608 (N_26608,N_25209,N_25674);
nor U26609 (N_26609,N_25732,N_25271);
xnor U26610 (N_26610,N_25677,N_25705);
or U26611 (N_26611,N_25851,N_25729);
or U26612 (N_26612,N_25458,N_25919);
nand U26613 (N_26613,N_25702,N_25406);
xnor U26614 (N_26614,N_25808,N_25770);
xnor U26615 (N_26615,N_25682,N_25778);
nand U26616 (N_26616,N_25159,N_25804);
xor U26617 (N_26617,N_25374,N_25400);
or U26618 (N_26618,N_25894,N_25897);
nor U26619 (N_26619,N_25422,N_25902);
or U26620 (N_26620,N_25976,N_25596);
xnor U26621 (N_26621,N_25599,N_25172);
xnor U26622 (N_26622,N_25834,N_25025);
or U26623 (N_26623,N_25185,N_25033);
or U26624 (N_26624,N_25683,N_25344);
nor U26625 (N_26625,N_25448,N_25494);
xor U26626 (N_26626,N_25690,N_25408);
xnor U26627 (N_26627,N_25549,N_25442);
or U26628 (N_26628,N_25950,N_25690);
nand U26629 (N_26629,N_25909,N_25938);
and U26630 (N_26630,N_25901,N_25974);
or U26631 (N_26631,N_25474,N_25508);
xor U26632 (N_26632,N_25548,N_25518);
or U26633 (N_26633,N_25793,N_25493);
xor U26634 (N_26634,N_25093,N_25437);
nand U26635 (N_26635,N_25981,N_25729);
and U26636 (N_26636,N_25051,N_25748);
nand U26637 (N_26637,N_25920,N_25549);
or U26638 (N_26638,N_25240,N_25503);
nand U26639 (N_26639,N_25358,N_25461);
nand U26640 (N_26640,N_25903,N_25338);
nor U26641 (N_26641,N_25361,N_25352);
xnor U26642 (N_26642,N_25220,N_25706);
xor U26643 (N_26643,N_25521,N_25034);
and U26644 (N_26644,N_25316,N_25162);
nand U26645 (N_26645,N_25305,N_25863);
nand U26646 (N_26646,N_25805,N_25397);
xor U26647 (N_26647,N_25856,N_25210);
and U26648 (N_26648,N_25736,N_25863);
nand U26649 (N_26649,N_25324,N_25828);
nand U26650 (N_26650,N_25816,N_25318);
nor U26651 (N_26651,N_25799,N_25080);
or U26652 (N_26652,N_25297,N_25692);
xnor U26653 (N_26653,N_25316,N_25301);
xnor U26654 (N_26654,N_25420,N_25654);
nor U26655 (N_26655,N_25381,N_25416);
nand U26656 (N_26656,N_25764,N_25835);
xnor U26657 (N_26657,N_25716,N_25849);
nand U26658 (N_26658,N_25486,N_25449);
nand U26659 (N_26659,N_25896,N_25169);
nand U26660 (N_26660,N_25932,N_25924);
and U26661 (N_26661,N_25558,N_25404);
or U26662 (N_26662,N_25079,N_25160);
or U26663 (N_26663,N_25708,N_25331);
xor U26664 (N_26664,N_25910,N_25224);
nand U26665 (N_26665,N_25740,N_25453);
nor U26666 (N_26666,N_25100,N_25237);
and U26667 (N_26667,N_25208,N_25723);
nor U26668 (N_26668,N_25112,N_25430);
or U26669 (N_26669,N_25151,N_25270);
and U26670 (N_26670,N_25183,N_25194);
nor U26671 (N_26671,N_25192,N_25871);
or U26672 (N_26672,N_25288,N_25616);
nor U26673 (N_26673,N_25305,N_25784);
nand U26674 (N_26674,N_25382,N_25455);
xor U26675 (N_26675,N_25889,N_25939);
xnor U26676 (N_26676,N_25454,N_25809);
nand U26677 (N_26677,N_25798,N_25487);
nand U26678 (N_26678,N_25779,N_25567);
nor U26679 (N_26679,N_25402,N_25454);
or U26680 (N_26680,N_25937,N_25088);
and U26681 (N_26681,N_25079,N_25520);
or U26682 (N_26682,N_25504,N_25028);
or U26683 (N_26683,N_25341,N_25625);
and U26684 (N_26684,N_25648,N_25897);
xnor U26685 (N_26685,N_25690,N_25813);
nor U26686 (N_26686,N_25518,N_25272);
and U26687 (N_26687,N_25345,N_25591);
nor U26688 (N_26688,N_25512,N_25383);
xor U26689 (N_26689,N_25104,N_25849);
xor U26690 (N_26690,N_25327,N_25087);
xor U26691 (N_26691,N_25143,N_25427);
and U26692 (N_26692,N_25317,N_25061);
xnor U26693 (N_26693,N_25941,N_25066);
and U26694 (N_26694,N_25610,N_25623);
nor U26695 (N_26695,N_25155,N_25132);
xnor U26696 (N_26696,N_25279,N_25920);
nor U26697 (N_26697,N_25208,N_25045);
and U26698 (N_26698,N_25541,N_25579);
nand U26699 (N_26699,N_25014,N_25370);
nand U26700 (N_26700,N_25507,N_25612);
nor U26701 (N_26701,N_25731,N_25221);
or U26702 (N_26702,N_25389,N_25534);
xnor U26703 (N_26703,N_25624,N_25004);
or U26704 (N_26704,N_25194,N_25056);
or U26705 (N_26705,N_25688,N_25997);
nand U26706 (N_26706,N_25227,N_25623);
nor U26707 (N_26707,N_25988,N_25783);
nor U26708 (N_26708,N_25128,N_25487);
or U26709 (N_26709,N_25783,N_25955);
xor U26710 (N_26710,N_25939,N_25825);
xnor U26711 (N_26711,N_25293,N_25477);
and U26712 (N_26712,N_25000,N_25899);
nand U26713 (N_26713,N_25397,N_25905);
nand U26714 (N_26714,N_25674,N_25089);
nor U26715 (N_26715,N_25924,N_25773);
and U26716 (N_26716,N_25992,N_25436);
xnor U26717 (N_26717,N_25713,N_25551);
xor U26718 (N_26718,N_25905,N_25474);
nor U26719 (N_26719,N_25107,N_25520);
and U26720 (N_26720,N_25963,N_25707);
or U26721 (N_26721,N_25998,N_25650);
and U26722 (N_26722,N_25362,N_25551);
or U26723 (N_26723,N_25754,N_25016);
xnor U26724 (N_26724,N_25588,N_25477);
xor U26725 (N_26725,N_25458,N_25651);
nand U26726 (N_26726,N_25493,N_25103);
nor U26727 (N_26727,N_25755,N_25604);
or U26728 (N_26728,N_25727,N_25719);
nand U26729 (N_26729,N_25544,N_25983);
and U26730 (N_26730,N_25434,N_25852);
or U26731 (N_26731,N_25746,N_25615);
nand U26732 (N_26732,N_25737,N_25743);
xnor U26733 (N_26733,N_25722,N_25518);
nor U26734 (N_26734,N_25196,N_25984);
or U26735 (N_26735,N_25962,N_25972);
and U26736 (N_26736,N_25053,N_25223);
nor U26737 (N_26737,N_25991,N_25018);
xnor U26738 (N_26738,N_25672,N_25168);
and U26739 (N_26739,N_25086,N_25482);
xnor U26740 (N_26740,N_25107,N_25380);
nand U26741 (N_26741,N_25665,N_25500);
or U26742 (N_26742,N_25941,N_25180);
xnor U26743 (N_26743,N_25850,N_25738);
xor U26744 (N_26744,N_25153,N_25623);
or U26745 (N_26745,N_25258,N_25544);
and U26746 (N_26746,N_25088,N_25780);
or U26747 (N_26747,N_25914,N_25638);
or U26748 (N_26748,N_25109,N_25157);
xor U26749 (N_26749,N_25942,N_25707);
or U26750 (N_26750,N_25285,N_25745);
nand U26751 (N_26751,N_25922,N_25557);
nand U26752 (N_26752,N_25401,N_25319);
and U26753 (N_26753,N_25715,N_25340);
nand U26754 (N_26754,N_25656,N_25862);
nand U26755 (N_26755,N_25460,N_25076);
nand U26756 (N_26756,N_25616,N_25667);
or U26757 (N_26757,N_25203,N_25873);
and U26758 (N_26758,N_25450,N_25642);
nand U26759 (N_26759,N_25450,N_25624);
nor U26760 (N_26760,N_25059,N_25682);
xnor U26761 (N_26761,N_25112,N_25081);
xor U26762 (N_26762,N_25653,N_25691);
nand U26763 (N_26763,N_25410,N_25292);
or U26764 (N_26764,N_25564,N_25335);
or U26765 (N_26765,N_25134,N_25101);
nor U26766 (N_26766,N_25762,N_25730);
nand U26767 (N_26767,N_25126,N_25587);
and U26768 (N_26768,N_25313,N_25094);
xnor U26769 (N_26769,N_25232,N_25467);
or U26770 (N_26770,N_25841,N_25316);
or U26771 (N_26771,N_25838,N_25551);
xnor U26772 (N_26772,N_25363,N_25541);
and U26773 (N_26773,N_25243,N_25657);
nand U26774 (N_26774,N_25275,N_25274);
nand U26775 (N_26775,N_25706,N_25274);
nor U26776 (N_26776,N_25804,N_25652);
nor U26777 (N_26777,N_25335,N_25765);
and U26778 (N_26778,N_25108,N_25215);
nand U26779 (N_26779,N_25477,N_25652);
nand U26780 (N_26780,N_25371,N_25864);
nand U26781 (N_26781,N_25053,N_25761);
or U26782 (N_26782,N_25515,N_25638);
or U26783 (N_26783,N_25073,N_25966);
nand U26784 (N_26784,N_25085,N_25402);
or U26785 (N_26785,N_25726,N_25403);
or U26786 (N_26786,N_25435,N_25964);
and U26787 (N_26787,N_25804,N_25549);
or U26788 (N_26788,N_25252,N_25237);
nor U26789 (N_26789,N_25975,N_25105);
and U26790 (N_26790,N_25087,N_25295);
and U26791 (N_26791,N_25219,N_25113);
nor U26792 (N_26792,N_25871,N_25896);
or U26793 (N_26793,N_25356,N_25168);
nor U26794 (N_26794,N_25487,N_25810);
nor U26795 (N_26795,N_25680,N_25468);
or U26796 (N_26796,N_25976,N_25920);
nor U26797 (N_26797,N_25379,N_25760);
and U26798 (N_26798,N_25569,N_25805);
or U26799 (N_26799,N_25006,N_25756);
xnor U26800 (N_26800,N_25376,N_25327);
or U26801 (N_26801,N_25871,N_25680);
nor U26802 (N_26802,N_25815,N_25525);
or U26803 (N_26803,N_25123,N_25848);
nor U26804 (N_26804,N_25365,N_25557);
xnor U26805 (N_26805,N_25387,N_25359);
nor U26806 (N_26806,N_25693,N_25726);
or U26807 (N_26807,N_25597,N_25969);
nor U26808 (N_26808,N_25413,N_25687);
or U26809 (N_26809,N_25417,N_25077);
or U26810 (N_26810,N_25419,N_25081);
or U26811 (N_26811,N_25219,N_25991);
and U26812 (N_26812,N_25236,N_25708);
and U26813 (N_26813,N_25670,N_25864);
or U26814 (N_26814,N_25974,N_25273);
xnor U26815 (N_26815,N_25299,N_25185);
nand U26816 (N_26816,N_25200,N_25483);
xor U26817 (N_26817,N_25431,N_25600);
nor U26818 (N_26818,N_25839,N_25210);
nand U26819 (N_26819,N_25523,N_25524);
nor U26820 (N_26820,N_25928,N_25232);
nor U26821 (N_26821,N_25885,N_25574);
nand U26822 (N_26822,N_25388,N_25903);
xnor U26823 (N_26823,N_25067,N_25687);
or U26824 (N_26824,N_25611,N_25463);
xnor U26825 (N_26825,N_25359,N_25510);
nor U26826 (N_26826,N_25140,N_25033);
and U26827 (N_26827,N_25914,N_25637);
or U26828 (N_26828,N_25053,N_25939);
nor U26829 (N_26829,N_25977,N_25443);
nand U26830 (N_26830,N_25185,N_25868);
nand U26831 (N_26831,N_25403,N_25853);
nor U26832 (N_26832,N_25352,N_25875);
or U26833 (N_26833,N_25661,N_25270);
nand U26834 (N_26834,N_25678,N_25805);
xnor U26835 (N_26835,N_25378,N_25661);
nor U26836 (N_26836,N_25435,N_25001);
or U26837 (N_26837,N_25899,N_25886);
nor U26838 (N_26838,N_25238,N_25209);
or U26839 (N_26839,N_25461,N_25760);
or U26840 (N_26840,N_25728,N_25412);
and U26841 (N_26841,N_25926,N_25457);
or U26842 (N_26842,N_25968,N_25467);
nand U26843 (N_26843,N_25618,N_25697);
xor U26844 (N_26844,N_25158,N_25898);
nor U26845 (N_26845,N_25785,N_25150);
nand U26846 (N_26846,N_25220,N_25166);
and U26847 (N_26847,N_25622,N_25130);
or U26848 (N_26848,N_25793,N_25345);
or U26849 (N_26849,N_25043,N_25221);
nand U26850 (N_26850,N_25324,N_25305);
nor U26851 (N_26851,N_25431,N_25049);
nand U26852 (N_26852,N_25796,N_25705);
and U26853 (N_26853,N_25898,N_25068);
xnor U26854 (N_26854,N_25266,N_25022);
or U26855 (N_26855,N_25878,N_25362);
and U26856 (N_26856,N_25991,N_25722);
or U26857 (N_26857,N_25484,N_25331);
and U26858 (N_26858,N_25385,N_25808);
or U26859 (N_26859,N_25683,N_25989);
nor U26860 (N_26860,N_25092,N_25858);
xor U26861 (N_26861,N_25498,N_25419);
nand U26862 (N_26862,N_25962,N_25821);
nand U26863 (N_26863,N_25687,N_25915);
xor U26864 (N_26864,N_25673,N_25429);
nor U26865 (N_26865,N_25823,N_25797);
nand U26866 (N_26866,N_25759,N_25893);
and U26867 (N_26867,N_25524,N_25467);
xor U26868 (N_26868,N_25887,N_25354);
xor U26869 (N_26869,N_25537,N_25024);
nand U26870 (N_26870,N_25588,N_25675);
xnor U26871 (N_26871,N_25046,N_25519);
nor U26872 (N_26872,N_25521,N_25575);
nor U26873 (N_26873,N_25182,N_25844);
nand U26874 (N_26874,N_25600,N_25678);
nand U26875 (N_26875,N_25045,N_25573);
or U26876 (N_26876,N_25942,N_25377);
xor U26877 (N_26877,N_25551,N_25540);
nand U26878 (N_26878,N_25124,N_25022);
nand U26879 (N_26879,N_25100,N_25524);
nor U26880 (N_26880,N_25772,N_25043);
or U26881 (N_26881,N_25058,N_25498);
nand U26882 (N_26882,N_25982,N_25658);
xor U26883 (N_26883,N_25344,N_25452);
xnor U26884 (N_26884,N_25628,N_25149);
xnor U26885 (N_26885,N_25974,N_25663);
nand U26886 (N_26886,N_25234,N_25315);
xor U26887 (N_26887,N_25375,N_25119);
nor U26888 (N_26888,N_25333,N_25798);
nand U26889 (N_26889,N_25588,N_25840);
nand U26890 (N_26890,N_25508,N_25359);
or U26891 (N_26891,N_25354,N_25424);
nand U26892 (N_26892,N_25748,N_25185);
nor U26893 (N_26893,N_25861,N_25634);
and U26894 (N_26894,N_25423,N_25364);
nand U26895 (N_26895,N_25387,N_25366);
nor U26896 (N_26896,N_25502,N_25360);
or U26897 (N_26897,N_25109,N_25234);
nand U26898 (N_26898,N_25228,N_25847);
or U26899 (N_26899,N_25168,N_25935);
or U26900 (N_26900,N_25677,N_25910);
nor U26901 (N_26901,N_25162,N_25666);
xor U26902 (N_26902,N_25796,N_25870);
nand U26903 (N_26903,N_25534,N_25072);
nand U26904 (N_26904,N_25620,N_25092);
nor U26905 (N_26905,N_25826,N_25299);
and U26906 (N_26906,N_25854,N_25570);
xor U26907 (N_26907,N_25354,N_25116);
and U26908 (N_26908,N_25516,N_25059);
nor U26909 (N_26909,N_25187,N_25455);
or U26910 (N_26910,N_25989,N_25111);
nor U26911 (N_26911,N_25030,N_25164);
and U26912 (N_26912,N_25911,N_25011);
nor U26913 (N_26913,N_25654,N_25071);
nand U26914 (N_26914,N_25955,N_25284);
nand U26915 (N_26915,N_25117,N_25327);
nand U26916 (N_26916,N_25659,N_25636);
or U26917 (N_26917,N_25112,N_25315);
and U26918 (N_26918,N_25681,N_25743);
nand U26919 (N_26919,N_25866,N_25335);
nor U26920 (N_26920,N_25444,N_25242);
nand U26921 (N_26921,N_25810,N_25027);
and U26922 (N_26922,N_25758,N_25249);
and U26923 (N_26923,N_25425,N_25305);
nand U26924 (N_26924,N_25452,N_25262);
and U26925 (N_26925,N_25636,N_25913);
nand U26926 (N_26926,N_25869,N_25267);
nand U26927 (N_26927,N_25892,N_25707);
xor U26928 (N_26928,N_25897,N_25076);
and U26929 (N_26929,N_25818,N_25768);
xor U26930 (N_26930,N_25773,N_25155);
xnor U26931 (N_26931,N_25540,N_25653);
nand U26932 (N_26932,N_25125,N_25758);
and U26933 (N_26933,N_25204,N_25410);
nor U26934 (N_26934,N_25841,N_25512);
or U26935 (N_26935,N_25731,N_25948);
xor U26936 (N_26936,N_25201,N_25902);
nand U26937 (N_26937,N_25014,N_25325);
xor U26938 (N_26938,N_25316,N_25951);
or U26939 (N_26939,N_25966,N_25472);
nand U26940 (N_26940,N_25679,N_25802);
or U26941 (N_26941,N_25189,N_25116);
xnor U26942 (N_26942,N_25075,N_25776);
or U26943 (N_26943,N_25133,N_25053);
and U26944 (N_26944,N_25349,N_25242);
nor U26945 (N_26945,N_25290,N_25928);
nand U26946 (N_26946,N_25626,N_25406);
xor U26947 (N_26947,N_25379,N_25856);
nand U26948 (N_26948,N_25669,N_25491);
and U26949 (N_26949,N_25871,N_25806);
or U26950 (N_26950,N_25307,N_25168);
nor U26951 (N_26951,N_25083,N_25268);
or U26952 (N_26952,N_25182,N_25506);
nand U26953 (N_26953,N_25196,N_25449);
nor U26954 (N_26954,N_25651,N_25257);
or U26955 (N_26955,N_25217,N_25497);
nor U26956 (N_26956,N_25450,N_25898);
xnor U26957 (N_26957,N_25603,N_25660);
xnor U26958 (N_26958,N_25539,N_25250);
and U26959 (N_26959,N_25430,N_25957);
and U26960 (N_26960,N_25336,N_25722);
nand U26961 (N_26961,N_25651,N_25616);
nor U26962 (N_26962,N_25443,N_25060);
xnor U26963 (N_26963,N_25870,N_25977);
or U26964 (N_26964,N_25858,N_25424);
xor U26965 (N_26965,N_25789,N_25407);
xnor U26966 (N_26966,N_25908,N_25078);
xnor U26967 (N_26967,N_25973,N_25832);
and U26968 (N_26968,N_25819,N_25860);
nor U26969 (N_26969,N_25117,N_25128);
nor U26970 (N_26970,N_25907,N_25580);
nor U26971 (N_26971,N_25184,N_25607);
xor U26972 (N_26972,N_25655,N_25736);
nand U26973 (N_26973,N_25950,N_25184);
or U26974 (N_26974,N_25241,N_25845);
xor U26975 (N_26975,N_25703,N_25389);
and U26976 (N_26976,N_25813,N_25619);
nor U26977 (N_26977,N_25507,N_25566);
or U26978 (N_26978,N_25472,N_25943);
nor U26979 (N_26979,N_25932,N_25220);
xnor U26980 (N_26980,N_25330,N_25032);
and U26981 (N_26981,N_25078,N_25168);
or U26982 (N_26982,N_25710,N_25510);
nand U26983 (N_26983,N_25352,N_25075);
and U26984 (N_26984,N_25100,N_25060);
or U26985 (N_26985,N_25263,N_25673);
and U26986 (N_26986,N_25752,N_25970);
and U26987 (N_26987,N_25025,N_25229);
xor U26988 (N_26988,N_25538,N_25808);
or U26989 (N_26989,N_25006,N_25091);
xor U26990 (N_26990,N_25328,N_25332);
or U26991 (N_26991,N_25626,N_25176);
or U26992 (N_26992,N_25890,N_25743);
and U26993 (N_26993,N_25659,N_25150);
nand U26994 (N_26994,N_25885,N_25926);
nand U26995 (N_26995,N_25477,N_25206);
and U26996 (N_26996,N_25009,N_25155);
xnor U26997 (N_26997,N_25019,N_25384);
nor U26998 (N_26998,N_25376,N_25662);
and U26999 (N_26999,N_25053,N_25113);
or U27000 (N_27000,N_26851,N_26305);
xor U27001 (N_27001,N_26063,N_26831);
nor U27002 (N_27002,N_26370,N_26164);
nand U27003 (N_27003,N_26438,N_26419);
nand U27004 (N_27004,N_26790,N_26277);
nand U27005 (N_27005,N_26103,N_26604);
nand U27006 (N_27006,N_26367,N_26818);
or U27007 (N_27007,N_26060,N_26774);
or U27008 (N_27008,N_26251,N_26990);
xor U27009 (N_27009,N_26929,N_26308);
nand U27010 (N_27010,N_26866,N_26890);
xnor U27011 (N_27011,N_26746,N_26214);
and U27012 (N_27012,N_26054,N_26192);
xor U27013 (N_27013,N_26098,N_26382);
nand U27014 (N_27014,N_26613,N_26337);
and U27015 (N_27015,N_26801,N_26835);
and U27016 (N_27016,N_26872,N_26876);
xor U27017 (N_27017,N_26538,N_26348);
nand U27018 (N_27018,N_26915,N_26518);
or U27019 (N_27019,N_26920,N_26747);
and U27020 (N_27020,N_26887,N_26979);
or U27021 (N_27021,N_26927,N_26300);
or U27022 (N_27022,N_26510,N_26625);
nand U27023 (N_27023,N_26521,N_26474);
nor U27024 (N_27024,N_26936,N_26946);
or U27025 (N_27025,N_26499,N_26830);
nand U27026 (N_27026,N_26468,N_26579);
xor U27027 (N_27027,N_26183,N_26947);
or U27028 (N_27028,N_26800,N_26254);
nand U27029 (N_27029,N_26430,N_26738);
or U27030 (N_27030,N_26374,N_26140);
nand U27031 (N_27031,N_26914,N_26173);
and U27032 (N_27032,N_26490,N_26565);
and U27033 (N_27033,N_26100,N_26478);
nor U27034 (N_27034,N_26006,N_26061);
nor U27035 (N_27035,N_26597,N_26475);
and U27036 (N_27036,N_26689,N_26533);
or U27037 (N_27037,N_26058,N_26182);
nand U27038 (N_27038,N_26617,N_26664);
or U27039 (N_27039,N_26428,N_26281);
and U27040 (N_27040,N_26718,N_26812);
nor U27041 (N_27041,N_26796,N_26065);
or U27042 (N_27042,N_26825,N_26445);
and U27043 (N_27043,N_26697,N_26148);
or U27044 (N_27044,N_26519,N_26488);
nor U27045 (N_27045,N_26657,N_26442);
nor U27046 (N_27046,N_26024,N_26603);
and U27047 (N_27047,N_26807,N_26163);
or U27048 (N_27048,N_26449,N_26081);
nor U27049 (N_27049,N_26332,N_26663);
xnor U27050 (N_27050,N_26950,N_26751);
xor U27051 (N_27051,N_26549,N_26383);
nand U27052 (N_27052,N_26783,N_26471);
xor U27053 (N_27053,N_26693,N_26619);
nor U27054 (N_27054,N_26939,N_26373);
nor U27055 (N_27055,N_26126,N_26647);
nor U27056 (N_27056,N_26992,N_26109);
xnor U27057 (N_27057,N_26605,N_26757);
or U27058 (N_27058,N_26223,N_26028);
or U27059 (N_27059,N_26033,N_26396);
or U27060 (N_27060,N_26102,N_26494);
nand U27061 (N_27061,N_26491,N_26497);
xor U27062 (N_27062,N_26883,N_26320);
nor U27063 (N_27063,N_26969,N_26856);
or U27064 (N_27064,N_26484,N_26191);
and U27065 (N_27065,N_26411,N_26863);
xor U27066 (N_27066,N_26688,N_26362);
nor U27067 (N_27067,N_26021,N_26864);
nor U27068 (N_27068,N_26176,N_26687);
or U27069 (N_27069,N_26143,N_26379);
or U27070 (N_27070,N_26528,N_26514);
and U27071 (N_27071,N_26433,N_26234);
and U27072 (N_27072,N_26010,N_26014);
nor U27073 (N_27073,N_26788,N_26586);
nand U27074 (N_27074,N_26246,N_26261);
and U27075 (N_27075,N_26338,N_26561);
or U27076 (N_27076,N_26294,N_26712);
nor U27077 (N_27077,N_26541,N_26084);
or U27078 (N_27078,N_26543,N_26841);
or U27079 (N_27079,N_26628,N_26575);
nor U27080 (N_27080,N_26716,N_26053);
or U27081 (N_27081,N_26492,N_26509);
xor U27082 (N_27082,N_26624,N_26439);
xor U27083 (N_27083,N_26948,N_26553);
nand U27084 (N_27084,N_26525,N_26465);
nor U27085 (N_27085,N_26290,N_26850);
and U27086 (N_27086,N_26902,N_26544);
nand U27087 (N_27087,N_26934,N_26211);
or U27088 (N_27088,N_26982,N_26015);
and U27089 (N_27089,N_26766,N_26356);
or U27090 (N_27090,N_26827,N_26039);
and U27091 (N_27091,N_26202,N_26600);
xor U27092 (N_27092,N_26258,N_26517);
and U27093 (N_27093,N_26086,N_26804);
nand U27094 (N_27094,N_26001,N_26623);
and U27095 (N_27095,N_26498,N_26351);
and U27096 (N_27096,N_26302,N_26366);
nor U27097 (N_27097,N_26997,N_26740);
or U27098 (N_27098,N_26966,N_26298);
xnor U27099 (N_27099,N_26878,N_26069);
xor U27100 (N_27100,N_26570,N_26775);
nand U27101 (N_27101,N_26675,N_26314);
nor U27102 (N_27102,N_26273,N_26527);
nor U27103 (N_27103,N_26728,N_26177);
nor U27104 (N_27104,N_26481,N_26380);
xnor U27105 (N_27105,N_26736,N_26376);
nand U27106 (N_27106,N_26354,N_26545);
nand U27107 (N_27107,N_26059,N_26529);
and U27108 (N_27108,N_26161,N_26245);
xor U27109 (N_27109,N_26447,N_26304);
xor U27110 (N_27110,N_26452,N_26218);
xor U27111 (N_27111,N_26194,N_26897);
or U27112 (N_27112,N_26861,N_26330);
nand U27113 (N_27113,N_26477,N_26881);
or U27114 (N_27114,N_26486,N_26115);
xnor U27115 (N_27115,N_26555,N_26323);
nor U27116 (N_27116,N_26141,N_26653);
xnor U27117 (N_27117,N_26469,N_26507);
or U27118 (N_27118,N_26896,N_26369);
and U27119 (N_27119,N_26077,N_26965);
nor U27120 (N_27120,N_26765,N_26405);
nor U27121 (N_27121,N_26315,N_26023);
and U27122 (N_27122,N_26560,N_26834);
and U27123 (N_27123,N_26311,N_26096);
nand U27124 (N_27124,N_26386,N_26008);
xor U27125 (N_27125,N_26048,N_26973);
nor U27126 (N_27126,N_26794,N_26793);
nand U27127 (N_27127,N_26406,N_26641);
and U27128 (N_27128,N_26991,N_26677);
nand U27129 (N_27129,N_26836,N_26826);
nand U27130 (N_27130,N_26620,N_26900);
and U27131 (N_27131,N_26935,N_26892);
or U27132 (N_27132,N_26926,N_26847);
and U27133 (N_27133,N_26867,N_26003);
and U27134 (N_27134,N_26853,N_26811);
and U27135 (N_27135,N_26165,N_26952);
xor U27136 (N_27136,N_26903,N_26090);
xnor U27137 (N_27137,N_26108,N_26955);
and U27138 (N_27138,N_26172,N_26901);
or U27139 (N_27139,N_26359,N_26020);
nor U27140 (N_27140,N_26798,N_26113);
nand U27141 (N_27141,N_26989,N_26174);
nor U27142 (N_27142,N_26256,N_26993);
nand U27143 (N_27143,N_26389,N_26885);
and U27144 (N_27144,N_26000,N_26208);
nand U27145 (N_27145,N_26523,N_26542);
xnor U27146 (N_27146,N_26120,N_26707);
nand U27147 (N_27147,N_26678,N_26476);
or U27148 (N_27148,N_26440,N_26274);
and U27149 (N_27149,N_26050,N_26524);
and U27150 (N_27150,N_26012,N_26802);
nand U27151 (N_27151,N_26967,N_26135);
or U27152 (N_27152,N_26673,N_26668);
xnor U27153 (N_27153,N_26780,N_26363);
nor U27154 (N_27154,N_26995,N_26175);
xnor U27155 (N_27155,N_26004,N_26401);
and U27156 (N_27156,N_26513,N_26789);
nor U27157 (N_27157,N_26658,N_26124);
or U27158 (N_27158,N_26742,N_26041);
xnor U27159 (N_27159,N_26503,N_26791);
and U27160 (N_27160,N_26080,N_26075);
nand U27161 (N_27161,N_26564,N_26259);
nor U27162 (N_27162,N_26860,N_26840);
nor U27163 (N_27163,N_26680,N_26987);
and U27164 (N_27164,N_26988,N_26127);
xnor U27165 (N_27165,N_26640,N_26614);
or U27166 (N_27166,N_26422,N_26919);
nor U27167 (N_27167,N_26207,N_26588);
nand U27168 (N_27168,N_26416,N_26325);
nor U27169 (N_27169,N_26042,N_26350);
and U27170 (N_27170,N_26632,N_26312);
nor U27171 (N_27171,N_26587,N_26682);
or U27172 (N_27172,N_26621,N_26980);
xor U27173 (N_27173,N_26353,N_26996);
xnor U27174 (N_27174,N_26752,N_26489);
nor U27175 (N_27175,N_26040,N_26838);
or U27176 (N_27176,N_26009,N_26157);
xnor U27177 (N_27177,N_26378,N_26377);
nand U27178 (N_27178,N_26293,N_26870);
xor U27179 (N_27179,N_26267,N_26983);
nor U27180 (N_27180,N_26155,N_26949);
or U27181 (N_27181,N_26928,N_26436);
nand U27182 (N_27182,N_26782,N_26977);
nand U27183 (N_27183,N_26729,N_26816);
nand U27184 (N_27184,N_26122,N_26390);
and U27185 (N_27185,N_26925,N_26898);
or U27186 (N_27186,N_26909,N_26094);
xnor U27187 (N_27187,N_26643,N_26216);
or U27188 (N_27188,N_26723,N_26871);
or U27189 (N_27189,N_26891,N_26594);
nor U27190 (N_27190,N_26843,N_26413);
and U27191 (N_27191,N_26150,N_26288);
nor U27192 (N_27192,N_26038,N_26333);
xor U27193 (N_27193,N_26593,N_26691);
xnor U27194 (N_27194,N_26085,N_26758);
and U27195 (N_27195,N_26397,N_26777);
nor U27196 (N_27196,N_26147,N_26635);
and U27197 (N_27197,N_26726,N_26408);
nand U27198 (N_27198,N_26893,N_26701);
xnor U27199 (N_27199,N_26567,N_26372);
or U27200 (N_27200,N_26340,N_26692);
xor U27201 (N_27201,N_26101,N_26644);
nor U27202 (N_27202,N_26754,N_26868);
xor U27203 (N_27203,N_26733,N_26959);
nand U27204 (N_27204,N_26829,N_26392);
xnor U27205 (N_27205,N_26184,N_26321);
and U27206 (N_27206,N_26088,N_26210);
nand U27207 (N_27207,N_26125,N_26859);
nand U27208 (N_27208,N_26667,N_26307);
or U27209 (N_27209,N_26745,N_26698);
and U27210 (N_27210,N_26704,N_26232);
or U27211 (N_27211,N_26819,N_26722);
nand U27212 (N_27212,N_26067,N_26130);
nand U27213 (N_27213,N_26237,N_26717);
nand U27214 (N_27214,N_26889,N_26737);
xor U27215 (N_27215,N_26329,N_26485);
nand U27216 (N_27216,N_26646,N_26899);
or U27217 (N_27217,N_26224,N_26295);
xor U27218 (N_27218,N_26402,N_26665);
or U27219 (N_27219,N_26598,N_26072);
or U27220 (N_27220,N_26612,N_26091);
nor U27221 (N_27221,N_26070,N_26581);
or U27222 (N_27222,N_26546,N_26132);
nor U27223 (N_27223,N_26420,N_26683);
or U27224 (N_27224,N_26036,N_26963);
xnor U27225 (N_27225,N_26076,N_26622);
nand U27226 (N_27226,N_26534,N_26852);
nand U27227 (N_27227,N_26426,N_26137);
nor U27228 (N_27228,N_26355,N_26837);
nor U27229 (N_27229,N_26068,N_26240);
and U27230 (N_27230,N_26670,N_26958);
nand U27231 (N_27231,N_26539,N_26153);
nor U27232 (N_27232,N_26432,N_26154);
nor U27233 (N_27233,N_26626,N_26656);
and U27234 (N_27234,N_26134,N_26185);
and U27235 (N_27235,N_26264,N_26806);
or U27236 (N_27236,N_26779,N_26171);
nand U27237 (N_27237,N_26720,N_26417);
and U27238 (N_27238,N_26652,N_26703);
and U27239 (N_27239,N_26022,N_26199);
xor U27240 (N_27240,N_26654,N_26005);
xnor U27241 (N_27241,N_26971,N_26552);
nand U27242 (N_27242,N_26650,N_26713);
and U27243 (N_27243,N_26882,N_26287);
or U27244 (N_27244,N_26099,N_26708);
xnor U27245 (N_27245,N_26522,N_26299);
nor U27246 (N_27246,N_26444,N_26725);
nor U27247 (N_27247,N_26342,N_26945);
and U27248 (N_27248,N_26188,N_26272);
and U27249 (N_27249,N_26773,N_26795);
or U27250 (N_27250,N_26271,N_26152);
nor U27251 (N_27251,N_26985,N_26711);
xnor U27252 (N_27252,N_26110,N_26398);
or U27253 (N_27253,N_26998,N_26414);
or U27254 (N_27254,N_26778,N_26424);
or U27255 (N_27255,N_26505,N_26201);
nor U27256 (N_27256,N_26227,N_26249);
nor U27257 (N_27257,N_26292,N_26276);
xnor U27258 (N_27258,N_26467,N_26375);
nand U27259 (N_27259,N_26809,N_26384);
or U27260 (N_27260,N_26388,N_26285);
nand U27261 (N_27261,N_26423,N_26451);
xnor U27262 (N_27262,N_26862,N_26629);
xor U27263 (N_27263,N_26443,N_26255);
xnor U27264 (N_27264,N_26470,N_26573);
nand U27265 (N_27265,N_26975,N_26516);
or U27266 (N_27266,N_26031,N_26869);
nand U27267 (N_27267,N_26087,N_26219);
nor U27268 (N_27268,N_26360,N_26263);
and U27269 (N_27269,N_26336,N_26242);
nor U27270 (N_27270,N_26159,N_26345);
nor U27271 (N_27271,N_26911,N_26496);
xnor U27272 (N_27272,N_26933,N_26578);
nor U27273 (N_27273,N_26170,N_26093);
nor U27274 (N_27274,N_26418,N_26026);
nor U27275 (N_27275,N_26324,N_26705);
or U27276 (N_27276,N_26410,N_26787);
or U27277 (N_27277,N_26457,N_26195);
and U27278 (N_27278,N_26347,N_26762);
and U27279 (N_27279,N_26681,N_26116);
nor U27280 (N_27280,N_26590,N_26554);
or U27281 (N_27281,N_26262,N_26536);
or U27282 (N_27282,N_26974,N_26844);
nand U27283 (N_27283,N_26011,N_26639);
and U27284 (N_27284,N_26136,N_26349);
nand U27285 (N_27285,N_26574,N_26661);
nand U27286 (N_27286,N_26095,N_26669);
and U27287 (N_27287,N_26118,N_26453);
or U27288 (N_27288,N_26531,N_26943);
xnor U27289 (N_27289,N_26257,N_26556);
nor U27290 (N_27290,N_26049,N_26530);
nand U27291 (N_27291,N_26250,N_26894);
nor U27292 (N_27292,N_26149,N_26279);
nor U27293 (N_27293,N_26940,N_26540);
xor U27294 (N_27294,N_26352,N_26145);
xnor U27295 (N_27295,N_26695,N_26266);
nor U27296 (N_27296,N_26052,N_26608);
nand U27297 (N_27297,N_26606,N_26968);
and U27298 (N_27298,N_26303,N_26462);
nand U27299 (N_27299,N_26030,N_26180);
nand U27300 (N_27300,N_26228,N_26111);
nor U27301 (N_27301,N_26855,N_26615);
or U27302 (N_27302,N_26166,N_26078);
nand U27303 (N_27303,N_26627,N_26319);
xnor U27304 (N_27304,N_26699,N_26412);
or U27305 (N_27305,N_26584,N_26932);
and U27306 (N_27306,N_26601,N_26854);
or U27307 (N_27307,N_26365,N_26634);
xnor U27308 (N_27308,N_26181,N_26781);
or U27309 (N_27309,N_26391,N_26358);
and U27310 (N_27310,N_26649,N_26976);
xor U27311 (N_27311,N_26483,N_26585);
nand U27312 (N_27312,N_26511,N_26395);
and U27313 (N_27313,N_26637,N_26289);
or U27314 (N_27314,N_26415,N_26660);
and U27315 (N_27315,N_26225,N_26296);
nand U27316 (N_27316,N_26741,N_26364);
nand U27317 (N_27317,N_26270,N_26814);
nor U27318 (N_27318,N_26937,N_26595);
nor U27319 (N_27319,N_26361,N_26631);
and U27320 (N_27320,N_26760,N_26501);
or U27321 (N_27321,N_26709,N_26446);
xor U27322 (N_27322,N_26055,N_26727);
nand U27323 (N_27323,N_26633,N_26431);
nor U27324 (N_27324,N_26756,N_26112);
and U27325 (N_27325,N_26252,N_26648);
nor U27326 (N_27326,N_26269,N_26906);
nand U27327 (N_27327,N_26400,N_26032);
xnor U27328 (N_27328,N_26138,N_26817);
xnor U27329 (N_27329,N_26146,N_26198);
nand U27330 (N_27330,N_26822,N_26659);
nor U27331 (N_27331,N_26931,N_26387);
xor U27332 (N_27332,N_26128,N_26160);
nor U27333 (N_27333,N_26907,N_26815);
and U27334 (N_27334,N_26645,N_26941);
or U27335 (N_27335,N_26071,N_26810);
or U27336 (N_27336,N_26265,N_26761);
or U27337 (N_27337,N_26685,N_26073);
and U27338 (N_27338,N_26922,N_26743);
nand U27339 (N_27339,N_26089,N_26823);
and U27340 (N_27340,N_26301,N_26846);
or U27341 (N_27341,N_26248,N_26607);
nor U27342 (N_27342,N_26018,N_26755);
nor U27343 (N_27343,N_26924,N_26448);
xor U27344 (N_27344,N_26129,N_26082);
or U27345 (N_27345,N_26912,N_26616);
and U27346 (N_27346,N_26253,N_26849);
or U27347 (N_27347,N_26480,N_26178);
xnor U27348 (N_27348,N_26403,N_26306);
nor U27349 (N_27349,N_26557,N_26904);
and U27350 (N_27350,N_26425,N_26580);
nor U27351 (N_27351,N_26156,N_26611);
nor U27352 (N_27352,N_26334,N_26602);
nor U27353 (N_27353,N_26123,N_26651);
nand U27354 (N_27354,N_26526,N_26784);
nor U27355 (N_27355,N_26450,N_26763);
and U27356 (N_27356,N_26857,N_26551);
nor U27357 (N_27357,N_26236,N_26286);
and U27358 (N_27358,N_26599,N_26671);
nand U27359 (N_27359,N_26002,N_26437);
nand U27360 (N_27360,N_26828,N_26454);
xor U27361 (N_27361,N_26873,N_26189);
nor U27362 (N_27362,N_26502,N_26694);
nand U27363 (N_27363,N_26577,N_26335);
nor U27364 (N_27364,N_26618,N_26962);
nand U27365 (N_27365,N_26131,N_26385);
and U27366 (N_27366,N_26275,N_26917);
or U27367 (N_27367,N_26957,N_26535);
and U27368 (N_27368,N_26799,N_26092);
and U27369 (N_27369,N_26759,N_26994);
and U27370 (N_27370,N_26638,N_26187);
xnor U27371 (N_27371,N_26562,N_26047);
xor U27372 (N_27372,N_26179,N_26046);
and U27373 (N_27373,N_26074,N_26710);
and U27374 (N_27374,N_26767,N_26119);
nor U27375 (N_27375,N_26655,N_26220);
or U27376 (N_27376,N_26824,N_26676);
and U27377 (N_27377,N_26190,N_26700);
or U27378 (N_27378,N_26500,N_26504);
xor U27379 (N_27379,N_26913,N_26684);
xnor U27380 (N_27380,N_26461,N_26235);
or U27381 (N_27381,N_26596,N_26479);
nand U27382 (N_27382,N_26786,N_26686);
nor U27383 (N_27383,N_26435,N_26037);
nor U27384 (N_27384,N_26730,N_26884);
xor U27385 (N_27385,N_26547,N_26456);
and U27386 (N_27386,N_26203,N_26019);
and U27387 (N_27387,N_26404,N_26589);
nand U27388 (N_27388,N_26714,N_26317);
or U27389 (N_27389,N_26107,N_26548);
and U27390 (N_27390,N_26984,N_26785);
xnor U27391 (N_27391,N_26297,N_26144);
or U27392 (N_27392,N_26986,N_26609);
xor U27393 (N_27393,N_26916,N_26007);
nor U27394 (N_27394,N_26241,N_26744);
nor U27395 (N_27395,N_26520,N_26642);
xnor U27396 (N_27396,N_26283,N_26879);
xor U27397 (N_27397,N_26464,N_26865);
and U27398 (N_27398,N_26886,N_26895);
nand U27399 (N_27399,N_26630,N_26221);
and U27400 (N_27400,N_26572,N_26724);
and U27401 (N_27401,N_26662,N_26772);
or U27402 (N_27402,N_26169,N_26035);
or U27403 (N_27403,N_26013,N_26016);
xor U27404 (N_27404,N_26247,N_26243);
or U27405 (N_27405,N_26776,N_26960);
nand U27406 (N_27406,N_26749,N_26322);
xnor U27407 (N_27407,N_26381,N_26466);
nand U27408 (N_27408,N_26515,N_26908);
or U27409 (N_27409,N_26813,N_26158);
nor U27410 (N_27410,N_26506,N_26981);
xnor U27411 (N_27411,N_26291,N_26209);
nor U27412 (N_27412,N_26768,N_26399);
xor U27413 (N_27413,N_26197,N_26151);
nor U27414 (N_27414,N_26318,N_26953);
xor U27415 (N_27415,N_26346,N_26268);
nor U27416 (N_27416,N_26739,N_26942);
nand U27417 (N_27417,N_26139,N_26051);
or U27418 (N_27418,N_26167,N_26848);
nor U27419 (N_27419,N_26944,N_26532);
nor U27420 (N_27420,N_26674,N_26706);
and U27421 (N_27421,N_26029,N_26792);
nor U27422 (N_27422,N_26732,N_26582);
or U27423 (N_27423,N_26769,N_26905);
or U27424 (N_27424,N_26690,N_26217);
xor U27425 (N_27425,N_26910,N_26162);
and U27426 (N_27426,N_26239,N_26057);
or U27427 (N_27427,N_26079,N_26458);
or U27428 (N_27428,N_26874,N_26213);
nor U27429 (N_27429,N_26017,N_26244);
nand U27430 (N_27430,N_26429,N_26133);
or U27431 (N_27431,N_26226,N_26341);
or U27432 (N_27432,N_26064,N_26434);
or U27433 (N_27433,N_26820,N_26186);
xnor U27434 (N_27434,N_26563,N_26394);
and U27435 (N_27435,N_26284,N_26313);
or U27436 (N_27436,N_26231,N_26368);
nand U27437 (N_27437,N_26487,N_26702);
nor U27438 (N_27438,N_26459,N_26845);
xor U27439 (N_27439,N_26972,N_26566);
xnor U27440 (N_27440,N_26463,N_26238);
xor U27441 (N_27441,N_26328,N_26877);
nor U27442 (N_27442,N_26875,N_26105);
nor U27443 (N_27443,N_26044,N_26421);
nor U27444 (N_27444,N_26558,N_26576);
xnor U27445 (N_27445,N_26964,N_26316);
or U27446 (N_27446,N_26770,N_26821);
or U27447 (N_27447,N_26888,N_26260);
nor U27448 (N_27448,N_26025,N_26923);
nand U27449 (N_27449,N_26808,N_26951);
nand U27450 (N_27450,N_26339,N_26204);
nand U27451 (N_27451,N_26310,N_26482);
or U27452 (N_27452,N_26961,N_26493);
and U27453 (N_27453,N_26331,N_26921);
or U27454 (N_27454,N_26097,N_26066);
nand U27455 (N_27455,N_26956,N_26978);
xnor U27456 (N_27456,N_26679,N_26734);
nand U27457 (N_27457,N_26880,N_26610);
nand U27458 (N_27458,N_26230,N_26508);
nand U27459 (N_27459,N_26282,N_26833);
nand U27460 (N_27460,N_26027,N_26731);
and U27461 (N_27461,N_26999,N_26954);
nand U27462 (N_27462,N_26441,N_26193);
or U27463 (N_27463,N_26121,N_26344);
and U27464 (N_27464,N_26205,N_26559);
and U27465 (N_27465,N_26666,N_26056);
and U27466 (N_27466,N_26672,N_26721);
nor U27467 (N_27467,N_26764,N_26215);
nor U27468 (N_27468,N_26233,N_26719);
nand U27469 (N_27469,N_26858,N_26550);
xor U27470 (N_27470,N_26393,N_26326);
xnor U27471 (N_27471,N_26034,N_26280);
xor U27472 (N_27472,N_26309,N_26472);
nor U27473 (N_27473,N_26636,N_26455);
and U27474 (N_27474,N_26537,N_26473);
xor U27475 (N_27475,N_26083,N_26212);
nor U27476 (N_27476,N_26427,N_26460);
xnor U27477 (N_27477,N_26327,N_26771);
xnor U27478 (N_27478,N_26753,N_26045);
nand U27479 (N_27479,N_26591,N_26696);
nor U27480 (N_27480,N_26357,N_26748);
and U27481 (N_27481,N_26117,N_26206);
and U27482 (N_27482,N_26832,N_26930);
nor U27483 (N_27483,N_26106,N_26278);
nand U27484 (N_27484,N_26568,N_26142);
xnor U27485 (N_27485,N_26371,N_26750);
xor U27486 (N_27486,N_26803,N_26842);
or U27487 (N_27487,N_26114,N_26839);
or U27488 (N_27488,N_26918,N_26938);
xor U27489 (N_27489,N_26062,N_26797);
and U27490 (N_27490,N_26196,N_26495);
or U27491 (N_27491,N_26343,N_26043);
or U27492 (N_27492,N_26583,N_26407);
nor U27493 (N_27493,N_26512,N_26592);
and U27494 (N_27494,N_26222,N_26571);
xnor U27495 (N_27495,N_26569,N_26168);
and U27496 (N_27496,N_26200,N_26715);
nor U27497 (N_27497,N_26970,N_26229);
and U27498 (N_27498,N_26735,N_26805);
and U27499 (N_27499,N_26409,N_26104);
and U27500 (N_27500,N_26642,N_26004);
xor U27501 (N_27501,N_26966,N_26483);
nand U27502 (N_27502,N_26028,N_26915);
nor U27503 (N_27503,N_26698,N_26812);
and U27504 (N_27504,N_26958,N_26124);
xnor U27505 (N_27505,N_26036,N_26948);
nor U27506 (N_27506,N_26718,N_26743);
and U27507 (N_27507,N_26686,N_26721);
nand U27508 (N_27508,N_26194,N_26215);
nand U27509 (N_27509,N_26975,N_26024);
and U27510 (N_27510,N_26133,N_26027);
xnor U27511 (N_27511,N_26671,N_26888);
or U27512 (N_27512,N_26699,N_26747);
nor U27513 (N_27513,N_26994,N_26495);
nor U27514 (N_27514,N_26795,N_26213);
and U27515 (N_27515,N_26382,N_26306);
nand U27516 (N_27516,N_26093,N_26895);
xnor U27517 (N_27517,N_26221,N_26187);
and U27518 (N_27518,N_26945,N_26430);
or U27519 (N_27519,N_26556,N_26113);
or U27520 (N_27520,N_26706,N_26292);
and U27521 (N_27521,N_26264,N_26357);
nand U27522 (N_27522,N_26611,N_26992);
xnor U27523 (N_27523,N_26690,N_26745);
and U27524 (N_27524,N_26046,N_26504);
nor U27525 (N_27525,N_26297,N_26980);
or U27526 (N_27526,N_26150,N_26336);
nand U27527 (N_27527,N_26525,N_26795);
nor U27528 (N_27528,N_26194,N_26066);
or U27529 (N_27529,N_26090,N_26726);
xnor U27530 (N_27530,N_26672,N_26985);
and U27531 (N_27531,N_26451,N_26342);
xor U27532 (N_27532,N_26302,N_26089);
and U27533 (N_27533,N_26309,N_26918);
and U27534 (N_27534,N_26821,N_26749);
nand U27535 (N_27535,N_26488,N_26958);
nor U27536 (N_27536,N_26932,N_26590);
nand U27537 (N_27537,N_26838,N_26716);
nor U27538 (N_27538,N_26579,N_26045);
and U27539 (N_27539,N_26449,N_26787);
xnor U27540 (N_27540,N_26848,N_26165);
and U27541 (N_27541,N_26143,N_26510);
nand U27542 (N_27542,N_26832,N_26214);
nand U27543 (N_27543,N_26602,N_26847);
nand U27544 (N_27544,N_26673,N_26660);
nand U27545 (N_27545,N_26965,N_26150);
xor U27546 (N_27546,N_26186,N_26461);
nor U27547 (N_27547,N_26205,N_26646);
nand U27548 (N_27548,N_26968,N_26021);
xnor U27549 (N_27549,N_26544,N_26345);
nor U27550 (N_27550,N_26722,N_26006);
and U27551 (N_27551,N_26503,N_26061);
and U27552 (N_27552,N_26771,N_26755);
xor U27553 (N_27553,N_26018,N_26352);
or U27554 (N_27554,N_26872,N_26601);
xnor U27555 (N_27555,N_26544,N_26838);
and U27556 (N_27556,N_26777,N_26668);
nor U27557 (N_27557,N_26291,N_26543);
nand U27558 (N_27558,N_26972,N_26506);
and U27559 (N_27559,N_26721,N_26945);
or U27560 (N_27560,N_26680,N_26103);
nor U27561 (N_27561,N_26857,N_26416);
xor U27562 (N_27562,N_26668,N_26515);
xor U27563 (N_27563,N_26580,N_26510);
nand U27564 (N_27564,N_26831,N_26264);
or U27565 (N_27565,N_26236,N_26785);
nor U27566 (N_27566,N_26989,N_26326);
xnor U27567 (N_27567,N_26148,N_26719);
nand U27568 (N_27568,N_26766,N_26378);
xnor U27569 (N_27569,N_26072,N_26893);
xor U27570 (N_27570,N_26073,N_26275);
or U27571 (N_27571,N_26023,N_26909);
nand U27572 (N_27572,N_26530,N_26248);
nand U27573 (N_27573,N_26370,N_26285);
nand U27574 (N_27574,N_26906,N_26991);
xor U27575 (N_27575,N_26963,N_26669);
or U27576 (N_27576,N_26860,N_26530);
or U27577 (N_27577,N_26702,N_26619);
nand U27578 (N_27578,N_26950,N_26508);
xnor U27579 (N_27579,N_26423,N_26543);
xnor U27580 (N_27580,N_26395,N_26408);
xor U27581 (N_27581,N_26548,N_26070);
xor U27582 (N_27582,N_26946,N_26286);
nor U27583 (N_27583,N_26805,N_26031);
nand U27584 (N_27584,N_26867,N_26156);
and U27585 (N_27585,N_26901,N_26514);
and U27586 (N_27586,N_26890,N_26161);
or U27587 (N_27587,N_26485,N_26694);
nand U27588 (N_27588,N_26223,N_26986);
nor U27589 (N_27589,N_26579,N_26324);
nor U27590 (N_27590,N_26361,N_26851);
xnor U27591 (N_27591,N_26369,N_26543);
xor U27592 (N_27592,N_26624,N_26325);
nand U27593 (N_27593,N_26418,N_26976);
nand U27594 (N_27594,N_26770,N_26030);
and U27595 (N_27595,N_26098,N_26608);
nor U27596 (N_27596,N_26084,N_26163);
and U27597 (N_27597,N_26626,N_26967);
or U27598 (N_27598,N_26901,N_26742);
nand U27599 (N_27599,N_26265,N_26573);
xnor U27600 (N_27600,N_26875,N_26625);
or U27601 (N_27601,N_26598,N_26412);
and U27602 (N_27602,N_26560,N_26039);
or U27603 (N_27603,N_26985,N_26609);
xor U27604 (N_27604,N_26960,N_26540);
nor U27605 (N_27605,N_26841,N_26688);
and U27606 (N_27606,N_26782,N_26355);
xnor U27607 (N_27607,N_26390,N_26663);
nand U27608 (N_27608,N_26154,N_26797);
or U27609 (N_27609,N_26191,N_26927);
or U27610 (N_27610,N_26490,N_26189);
xor U27611 (N_27611,N_26648,N_26072);
nor U27612 (N_27612,N_26868,N_26561);
nand U27613 (N_27613,N_26273,N_26385);
nand U27614 (N_27614,N_26572,N_26050);
nand U27615 (N_27615,N_26004,N_26584);
nand U27616 (N_27616,N_26737,N_26891);
and U27617 (N_27617,N_26225,N_26586);
or U27618 (N_27618,N_26733,N_26730);
xnor U27619 (N_27619,N_26815,N_26970);
and U27620 (N_27620,N_26180,N_26333);
or U27621 (N_27621,N_26698,N_26620);
and U27622 (N_27622,N_26878,N_26667);
and U27623 (N_27623,N_26697,N_26789);
nor U27624 (N_27624,N_26381,N_26789);
xor U27625 (N_27625,N_26192,N_26419);
or U27626 (N_27626,N_26547,N_26687);
or U27627 (N_27627,N_26013,N_26464);
nor U27628 (N_27628,N_26258,N_26097);
nor U27629 (N_27629,N_26530,N_26362);
and U27630 (N_27630,N_26670,N_26299);
xnor U27631 (N_27631,N_26831,N_26693);
nand U27632 (N_27632,N_26189,N_26180);
nor U27633 (N_27633,N_26034,N_26650);
and U27634 (N_27634,N_26385,N_26142);
and U27635 (N_27635,N_26074,N_26783);
and U27636 (N_27636,N_26692,N_26944);
nand U27637 (N_27637,N_26895,N_26735);
nor U27638 (N_27638,N_26991,N_26709);
xor U27639 (N_27639,N_26806,N_26854);
and U27640 (N_27640,N_26692,N_26096);
and U27641 (N_27641,N_26858,N_26547);
nand U27642 (N_27642,N_26425,N_26405);
and U27643 (N_27643,N_26163,N_26065);
or U27644 (N_27644,N_26098,N_26698);
or U27645 (N_27645,N_26582,N_26516);
xnor U27646 (N_27646,N_26852,N_26601);
nor U27647 (N_27647,N_26961,N_26765);
xor U27648 (N_27648,N_26866,N_26168);
nand U27649 (N_27649,N_26174,N_26516);
or U27650 (N_27650,N_26661,N_26994);
and U27651 (N_27651,N_26648,N_26057);
or U27652 (N_27652,N_26157,N_26375);
nor U27653 (N_27653,N_26683,N_26815);
nor U27654 (N_27654,N_26223,N_26588);
or U27655 (N_27655,N_26176,N_26674);
xor U27656 (N_27656,N_26109,N_26481);
or U27657 (N_27657,N_26686,N_26189);
and U27658 (N_27658,N_26407,N_26381);
xor U27659 (N_27659,N_26915,N_26021);
xnor U27660 (N_27660,N_26859,N_26029);
and U27661 (N_27661,N_26080,N_26699);
nor U27662 (N_27662,N_26938,N_26414);
nand U27663 (N_27663,N_26134,N_26706);
or U27664 (N_27664,N_26028,N_26086);
nand U27665 (N_27665,N_26494,N_26146);
or U27666 (N_27666,N_26544,N_26606);
xnor U27667 (N_27667,N_26564,N_26129);
xnor U27668 (N_27668,N_26606,N_26608);
xnor U27669 (N_27669,N_26819,N_26853);
nor U27670 (N_27670,N_26579,N_26057);
nand U27671 (N_27671,N_26152,N_26900);
or U27672 (N_27672,N_26068,N_26495);
nor U27673 (N_27673,N_26362,N_26064);
nand U27674 (N_27674,N_26070,N_26980);
and U27675 (N_27675,N_26193,N_26445);
nand U27676 (N_27676,N_26120,N_26354);
or U27677 (N_27677,N_26287,N_26231);
nor U27678 (N_27678,N_26939,N_26613);
nand U27679 (N_27679,N_26282,N_26610);
xnor U27680 (N_27680,N_26976,N_26999);
nand U27681 (N_27681,N_26060,N_26930);
nor U27682 (N_27682,N_26099,N_26855);
nor U27683 (N_27683,N_26913,N_26041);
and U27684 (N_27684,N_26992,N_26954);
nand U27685 (N_27685,N_26384,N_26872);
nand U27686 (N_27686,N_26713,N_26332);
nor U27687 (N_27687,N_26616,N_26953);
nand U27688 (N_27688,N_26586,N_26053);
nor U27689 (N_27689,N_26898,N_26934);
or U27690 (N_27690,N_26356,N_26740);
and U27691 (N_27691,N_26180,N_26992);
nand U27692 (N_27692,N_26741,N_26205);
nand U27693 (N_27693,N_26474,N_26902);
xnor U27694 (N_27694,N_26327,N_26968);
and U27695 (N_27695,N_26070,N_26582);
xnor U27696 (N_27696,N_26918,N_26589);
xnor U27697 (N_27697,N_26465,N_26365);
nor U27698 (N_27698,N_26644,N_26359);
and U27699 (N_27699,N_26217,N_26540);
nor U27700 (N_27700,N_26373,N_26633);
or U27701 (N_27701,N_26647,N_26538);
xnor U27702 (N_27702,N_26071,N_26626);
nand U27703 (N_27703,N_26572,N_26033);
nand U27704 (N_27704,N_26849,N_26889);
nand U27705 (N_27705,N_26939,N_26031);
or U27706 (N_27706,N_26222,N_26446);
or U27707 (N_27707,N_26144,N_26199);
xor U27708 (N_27708,N_26446,N_26066);
and U27709 (N_27709,N_26766,N_26388);
xnor U27710 (N_27710,N_26224,N_26023);
nor U27711 (N_27711,N_26044,N_26028);
nor U27712 (N_27712,N_26141,N_26348);
nor U27713 (N_27713,N_26174,N_26177);
and U27714 (N_27714,N_26878,N_26177);
nand U27715 (N_27715,N_26983,N_26958);
xnor U27716 (N_27716,N_26582,N_26329);
or U27717 (N_27717,N_26335,N_26538);
xnor U27718 (N_27718,N_26476,N_26303);
and U27719 (N_27719,N_26619,N_26105);
and U27720 (N_27720,N_26660,N_26122);
or U27721 (N_27721,N_26569,N_26646);
xnor U27722 (N_27722,N_26885,N_26542);
nor U27723 (N_27723,N_26574,N_26181);
xor U27724 (N_27724,N_26517,N_26295);
xnor U27725 (N_27725,N_26288,N_26087);
and U27726 (N_27726,N_26601,N_26244);
nor U27727 (N_27727,N_26269,N_26300);
and U27728 (N_27728,N_26039,N_26202);
nor U27729 (N_27729,N_26400,N_26453);
or U27730 (N_27730,N_26451,N_26667);
and U27731 (N_27731,N_26912,N_26209);
xor U27732 (N_27732,N_26390,N_26169);
nor U27733 (N_27733,N_26824,N_26279);
nand U27734 (N_27734,N_26495,N_26437);
nand U27735 (N_27735,N_26106,N_26633);
nor U27736 (N_27736,N_26731,N_26945);
nor U27737 (N_27737,N_26305,N_26927);
or U27738 (N_27738,N_26875,N_26260);
nand U27739 (N_27739,N_26082,N_26034);
nand U27740 (N_27740,N_26243,N_26125);
nand U27741 (N_27741,N_26908,N_26711);
nand U27742 (N_27742,N_26150,N_26875);
xnor U27743 (N_27743,N_26800,N_26803);
and U27744 (N_27744,N_26379,N_26546);
and U27745 (N_27745,N_26282,N_26835);
nand U27746 (N_27746,N_26314,N_26827);
or U27747 (N_27747,N_26378,N_26480);
and U27748 (N_27748,N_26643,N_26836);
xnor U27749 (N_27749,N_26017,N_26185);
nand U27750 (N_27750,N_26851,N_26422);
nor U27751 (N_27751,N_26683,N_26338);
nand U27752 (N_27752,N_26291,N_26519);
or U27753 (N_27753,N_26910,N_26266);
or U27754 (N_27754,N_26312,N_26530);
nand U27755 (N_27755,N_26126,N_26138);
or U27756 (N_27756,N_26516,N_26711);
and U27757 (N_27757,N_26754,N_26538);
nor U27758 (N_27758,N_26395,N_26383);
xnor U27759 (N_27759,N_26226,N_26806);
or U27760 (N_27760,N_26555,N_26161);
xnor U27761 (N_27761,N_26594,N_26627);
nor U27762 (N_27762,N_26292,N_26561);
nor U27763 (N_27763,N_26040,N_26113);
nor U27764 (N_27764,N_26790,N_26434);
nand U27765 (N_27765,N_26496,N_26896);
and U27766 (N_27766,N_26238,N_26900);
nor U27767 (N_27767,N_26521,N_26139);
or U27768 (N_27768,N_26090,N_26466);
and U27769 (N_27769,N_26239,N_26260);
nand U27770 (N_27770,N_26221,N_26664);
and U27771 (N_27771,N_26942,N_26279);
nand U27772 (N_27772,N_26699,N_26748);
xnor U27773 (N_27773,N_26293,N_26775);
or U27774 (N_27774,N_26140,N_26845);
or U27775 (N_27775,N_26544,N_26770);
or U27776 (N_27776,N_26324,N_26361);
xor U27777 (N_27777,N_26506,N_26276);
nor U27778 (N_27778,N_26442,N_26087);
nor U27779 (N_27779,N_26402,N_26768);
xnor U27780 (N_27780,N_26583,N_26489);
nand U27781 (N_27781,N_26729,N_26727);
nand U27782 (N_27782,N_26402,N_26724);
nand U27783 (N_27783,N_26218,N_26732);
or U27784 (N_27784,N_26702,N_26016);
nor U27785 (N_27785,N_26584,N_26211);
or U27786 (N_27786,N_26484,N_26653);
and U27787 (N_27787,N_26210,N_26148);
or U27788 (N_27788,N_26209,N_26740);
nor U27789 (N_27789,N_26097,N_26570);
and U27790 (N_27790,N_26175,N_26901);
or U27791 (N_27791,N_26817,N_26705);
nor U27792 (N_27792,N_26608,N_26266);
xnor U27793 (N_27793,N_26410,N_26213);
nand U27794 (N_27794,N_26162,N_26588);
nand U27795 (N_27795,N_26393,N_26206);
nand U27796 (N_27796,N_26847,N_26712);
and U27797 (N_27797,N_26705,N_26209);
nor U27798 (N_27798,N_26116,N_26500);
and U27799 (N_27799,N_26277,N_26321);
and U27800 (N_27800,N_26987,N_26166);
or U27801 (N_27801,N_26062,N_26371);
xnor U27802 (N_27802,N_26868,N_26269);
xnor U27803 (N_27803,N_26820,N_26804);
nand U27804 (N_27804,N_26872,N_26011);
nor U27805 (N_27805,N_26773,N_26945);
xnor U27806 (N_27806,N_26287,N_26150);
and U27807 (N_27807,N_26895,N_26755);
nand U27808 (N_27808,N_26599,N_26912);
xnor U27809 (N_27809,N_26193,N_26645);
nand U27810 (N_27810,N_26713,N_26295);
nand U27811 (N_27811,N_26954,N_26016);
or U27812 (N_27812,N_26116,N_26689);
xnor U27813 (N_27813,N_26220,N_26688);
xor U27814 (N_27814,N_26420,N_26220);
nor U27815 (N_27815,N_26124,N_26483);
nand U27816 (N_27816,N_26632,N_26126);
nor U27817 (N_27817,N_26939,N_26953);
or U27818 (N_27818,N_26357,N_26467);
or U27819 (N_27819,N_26716,N_26300);
nor U27820 (N_27820,N_26198,N_26569);
and U27821 (N_27821,N_26740,N_26033);
xor U27822 (N_27822,N_26600,N_26261);
nor U27823 (N_27823,N_26222,N_26201);
nand U27824 (N_27824,N_26269,N_26018);
nor U27825 (N_27825,N_26235,N_26425);
xnor U27826 (N_27826,N_26735,N_26127);
nor U27827 (N_27827,N_26463,N_26110);
nand U27828 (N_27828,N_26595,N_26943);
nand U27829 (N_27829,N_26023,N_26163);
nor U27830 (N_27830,N_26250,N_26611);
nand U27831 (N_27831,N_26363,N_26152);
nor U27832 (N_27832,N_26211,N_26967);
xor U27833 (N_27833,N_26759,N_26537);
or U27834 (N_27834,N_26863,N_26919);
or U27835 (N_27835,N_26132,N_26026);
or U27836 (N_27836,N_26383,N_26284);
or U27837 (N_27837,N_26394,N_26727);
or U27838 (N_27838,N_26388,N_26713);
xnor U27839 (N_27839,N_26971,N_26430);
nand U27840 (N_27840,N_26868,N_26948);
nand U27841 (N_27841,N_26272,N_26334);
xnor U27842 (N_27842,N_26346,N_26456);
xor U27843 (N_27843,N_26674,N_26344);
and U27844 (N_27844,N_26966,N_26468);
xnor U27845 (N_27845,N_26889,N_26841);
xor U27846 (N_27846,N_26061,N_26551);
xnor U27847 (N_27847,N_26230,N_26759);
and U27848 (N_27848,N_26245,N_26270);
xnor U27849 (N_27849,N_26162,N_26750);
nor U27850 (N_27850,N_26971,N_26911);
nand U27851 (N_27851,N_26637,N_26827);
nand U27852 (N_27852,N_26442,N_26845);
xnor U27853 (N_27853,N_26138,N_26580);
nand U27854 (N_27854,N_26433,N_26152);
nand U27855 (N_27855,N_26126,N_26158);
nand U27856 (N_27856,N_26199,N_26642);
nand U27857 (N_27857,N_26848,N_26633);
xor U27858 (N_27858,N_26591,N_26230);
nand U27859 (N_27859,N_26510,N_26675);
and U27860 (N_27860,N_26121,N_26966);
nor U27861 (N_27861,N_26018,N_26430);
and U27862 (N_27862,N_26167,N_26911);
or U27863 (N_27863,N_26326,N_26079);
or U27864 (N_27864,N_26365,N_26575);
and U27865 (N_27865,N_26984,N_26359);
or U27866 (N_27866,N_26481,N_26980);
nand U27867 (N_27867,N_26903,N_26921);
nand U27868 (N_27868,N_26924,N_26722);
or U27869 (N_27869,N_26387,N_26982);
nand U27870 (N_27870,N_26569,N_26607);
nor U27871 (N_27871,N_26926,N_26340);
nand U27872 (N_27872,N_26838,N_26373);
nor U27873 (N_27873,N_26700,N_26534);
nand U27874 (N_27874,N_26271,N_26965);
nor U27875 (N_27875,N_26622,N_26695);
and U27876 (N_27876,N_26951,N_26408);
nand U27877 (N_27877,N_26041,N_26088);
xnor U27878 (N_27878,N_26475,N_26236);
nor U27879 (N_27879,N_26390,N_26738);
and U27880 (N_27880,N_26345,N_26837);
nand U27881 (N_27881,N_26278,N_26399);
nor U27882 (N_27882,N_26496,N_26261);
and U27883 (N_27883,N_26149,N_26232);
xor U27884 (N_27884,N_26774,N_26337);
and U27885 (N_27885,N_26546,N_26641);
nor U27886 (N_27886,N_26828,N_26995);
nand U27887 (N_27887,N_26423,N_26322);
and U27888 (N_27888,N_26633,N_26318);
nand U27889 (N_27889,N_26234,N_26568);
nand U27890 (N_27890,N_26108,N_26751);
nand U27891 (N_27891,N_26303,N_26360);
and U27892 (N_27892,N_26945,N_26509);
or U27893 (N_27893,N_26176,N_26115);
nor U27894 (N_27894,N_26095,N_26189);
nand U27895 (N_27895,N_26953,N_26810);
or U27896 (N_27896,N_26043,N_26568);
xor U27897 (N_27897,N_26577,N_26979);
nor U27898 (N_27898,N_26038,N_26411);
nand U27899 (N_27899,N_26354,N_26710);
or U27900 (N_27900,N_26135,N_26821);
nand U27901 (N_27901,N_26881,N_26256);
xnor U27902 (N_27902,N_26072,N_26192);
nor U27903 (N_27903,N_26976,N_26505);
nand U27904 (N_27904,N_26156,N_26821);
nor U27905 (N_27905,N_26211,N_26687);
and U27906 (N_27906,N_26758,N_26084);
and U27907 (N_27907,N_26870,N_26459);
or U27908 (N_27908,N_26321,N_26431);
nand U27909 (N_27909,N_26954,N_26672);
nor U27910 (N_27910,N_26566,N_26870);
nor U27911 (N_27911,N_26182,N_26790);
nor U27912 (N_27912,N_26087,N_26940);
xor U27913 (N_27913,N_26503,N_26052);
nor U27914 (N_27914,N_26526,N_26729);
xor U27915 (N_27915,N_26697,N_26163);
or U27916 (N_27916,N_26008,N_26865);
and U27917 (N_27917,N_26566,N_26638);
or U27918 (N_27918,N_26482,N_26723);
and U27919 (N_27919,N_26070,N_26880);
xnor U27920 (N_27920,N_26587,N_26432);
xor U27921 (N_27921,N_26078,N_26513);
and U27922 (N_27922,N_26544,N_26156);
or U27923 (N_27923,N_26374,N_26002);
or U27924 (N_27924,N_26706,N_26557);
and U27925 (N_27925,N_26703,N_26994);
or U27926 (N_27926,N_26599,N_26585);
and U27927 (N_27927,N_26091,N_26402);
or U27928 (N_27928,N_26277,N_26147);
nand U27929 (N_27929,N_26356,N_26388);
and U27930 (N_27930,N_26634,N_26904);
and U27931 (N_27931,N_26269,N_26065);
and U27932 (N_27932,N_26395,N_26058);
xnor U27933 (N_27933,N_26328,N_26041);
and U27934 (N_27934,N_26949,N_26570);
xor U27935 (N_27935,N_26359,N_26599);
xnor U27936 (N_27936,N_26395,N_26402);
xor U27937 (N_27937,N_26317,N_26167);
xnor U27938 (N_27938,N_26216,N_26459);
xor U27939 (N_27939,N_26063,N_26957);
nor U27940 (N_27940,N_26564,N_26819);
xor U27941 (N_27941,N_26153,N_26282);
nor U27942 (N_27942,N_26579,N_26601);
nand U27943 (N_27943,N_26360,N_26194);
or U27944 (N_27944,N_26553,N_26428);
nand U27945 (N_27945,N_26161,N_26534);
nor U27946 (N_27946,N_26253,N_26278);
nor U27947 (N_27947,N_26975,N_26959);
xor U27948 (N_27948,N_26413,N_26046);
nor U27949 (N_27949,N_26206,N_26561);
nand U27950 (N_27950,N_26781,N_26193);
xnor U27951 (N_27951,N_26998,N_26643);
xnor U27952 (N_27952,N_26715,N_26171);
nand U27953 (N_27953,N_26544,N_26191);
nand U27954 (N_27954,N_26020,N_26153);
nor U27955 (N_27955,N_26914,N_26617);
or U27956 (N_27956,N_26193,N_26261);
nor U27957 (N_27957,N_26535,N_26373);
nand U27958 (N_27958,N_26330,N_26426);
and U27959 (N_27959,N_26539,N_26547);
nor U27960 (N_27960,N_26954,N_26061);
nor U27961 (N_27961,N_26402,N_26908);
xnor U27962 (N_27962,N_26315,N_26341);
xnor U27963 (N_27963,N_26774,N_26415);
nand U27964 (N_27964,N_26960,N_26850);
or U27965 (N_27965,N_26714,N_26089);
or U27966 (N_27966,N_26460,N_26578);
nand U27967 (N_27967,N_26018,N_26543);
and U27968 (N_27968,N_26481,N_26818);
xnor U27969 (N_27969,N_26359,N_26686);
or U27970 (N_27970,N_26323,N_26766);
nand U27971 (N_27971,N_26864,N_26851);
nor U27972 (N_27972,N_26008,N_26097);
nand U27973 (N_27973,N_26682,N_26528);
or U27974 (N_27974,N_26446,N_26741);
or U27975 (N_27975,N_26060,N_26729);
and U27976 (N_27976,N_26098,N_26130);
or U27977 (N_27977,N_26076,N_26538);
and U27978 (N_27978,N_26755,N_26577);
nor U27979 (N_27979,N_26611,N_26725);
xnor U27980 (N_27980,N_26367,N_26985);
and U27981 (N_27981,N_26493,N_26694);
nor U27982 (N_27982,N_26920,N_26254);
and U27983 (N_27983,N_26256,N_26814);
xor U27984 (N_27984,N_26340,N_26739);
or U27985 (N_27985,N_26402,N_26569);
nand U27986 (N_27986,N_26456,N_26520);
nand U27987 (N_27987,N_26786,N_26151);
nand U27988 (N_27988,N_26485,N_26585);
and U27989 (N_27989,N_26271,N_26062);
or U27990 (N_27990,N_26525,N_26748);
nand U27991 (N_27991,N_26166,N_26991);
or U27992 (N_27992,N_26996,N_26400);
and U27993 (N_27993,N_26300,N_26818);
xnor U27994 (N_27994,N_26523,N_26000);
nor U27995 (N_27995,N_26035,N_26096);
and U27996 (N_27996,N_26115,N_26468);
and U27997 (N_27997,N_26284,N_26691);
and U27998 (N_27998,N_26955,N_26755);
xor U27999 (N_27999,N_26469,N_26131);
nor U28000 (N_28000,N_27665,N_27068);
nand U28001 (N_28001,N_27435,N_27641);
or U28002 (N_28002,N_27828,N_27941);
nor U28003 (N_28003,N_27553,N_27397);
nor U28004 (N_28004,N_27320,N_27996);
xnor U28005 (N_28005,N_27658,N_27004);
nand U28006 (N_28006,N_27655,N_27365);
xor U28007 (N_28007,N_27968,N_27548);
or U28008 (N_28008,N_27599,N_27637);
nand U28009 (N_28009,N_27503,N_27562);
and U28010 (N_28010,N_27438,N_27829);
or U28011 (N_28011,N_27416,N_27494);
or U28012 (N_28012,N_27674,N_27942);
nor U28013 (N_28013,N_27608,N_27887);
nor U28014 (N_28014,N_27404,N_27134);
nor U28015 (N_28015,N_27958,N_27045);
and U28016 (N_28016,N_27322,N_27496);
nand U28017 (N_28017,N_27116,N_27881);
and U28018 (N_28018,N_27596,N_27474);
and U28019 (N_28019,N_27077,N_27648);
nor U28020 (N_28020,N_27678,N_27780);
nand U28021 (N_28021,N_27291,N_27306);
and U28022 (N_28022,N_27594,N_27737);
or U28023 (N_28023,N_27650,N_27726);
and U28024 (N_28024,N_27471,N_27411);
nor U28025 (N_28025,N_27777,N_27634);
nand U28026 (N_28026,N_27927,N_27788);
nand U28027 (N_28027,N_27749,N_27135);
xor U28028 (N_28028,N_27247,N_27528);
and U28029 (N_28029,N_27569,N_27452);
or U28030 (N_28030,N_27835,N_27377);
nand U28031 (N_28031,N_27181,N_27522);
and U28032 (N_28032,N_27771,N_27506);
or U28033 (N_28033,N_27087,N_27701);
or U28034 (N_28034,N_27285,N_27172);
nand U28035 (N_28035,N_27038,N_27132);
and U28036 (N_28036,N_27673,N_27531);
nor U28037 (N_28037,N_27501,N_27344);
or U28038 (N_28038,N_27157,N_27883);
xor U28039 (N_28039,N_27081,N_27111);
or U28040 (N_28040,N_27629,N_27082);
xnor U28041 (N_28041,N_27241,N_27511);
nor U28042 (N_28042,N_27192,N_27744);
xor U28043 (N_28043,N_27717,N_27310);
or U28044 (N_28044,N_27453,N_27497);
or U28045 (N_28045,N_27603,N_27721);
nand U28046 (N_28046,N_27418,N_27309);
and U28047 (N_28047,N_27010,N_27393);
and U28048 (N_28048,N_27574,N_27284);
nor U28049 (N_28049,N_27083,N_27651);
xnor U28050 (N_28050,N_27867,N_27601);
or U28051 (N_28051,N_27822,N_27140);
and U28052 (N_28052,N_27832,N_27710);
or U28053 (N_28053,N_27598,N_27577);
nor U28054 (N_28054,N_27845,N_27993);
or U28055 (N_28055,N_27900,N_27451);
xnor U28056 (N_28056,N_27373,N_27049);
nor U28057 (N_28057,N_27858,N_27850);
or U28058 (N_28058,N_27493,N_27782);
nand U28059 (N_28059,N_27733,N_27508);
or U28060 (N_28060,N_27959,N_27789);
and U28061 (N_28061,N_27946,N_27565);
and U28062 (N_28062,N_27663,N_27035);
nor U28063 (N_28063,N_27849,N_27675);
or U28064 (N_28064,N_27619,N_27752);
or U28065 (N_28065,N_27666,N_27816);
or U28066 (N_28066,N_27950,N_27419);
or U28067 (N_28067,N_27412,N_27628);
nor U28068 (N_28068,N_27570,N_27218);
xnor U28069 (N_28069,N_27421,N_27933);
or U28070 (N_28070,N_27409,N_27088);
nand U28071 (N_28071,N_27903,N_27221);
nor U28072 (N_28072,N_27699,N_27462);
nand U28073 (N_28073,N_27052,N_27078);
nor U28074 (N_28074,N_27547,N_27815);
nand U28075 (N_28075,N_27269,N_27504);
and U28076 (N_28076,N_27544,N_27423);
xor U28077 (N_28077,N_27066,N_27892);
or U28078 (N_28078,N_27693,N_27575);
xnor U28079 (N_28079,N_27236,N_27338);
and U28080 (N_28080,N_27329,N_27841);
nand U28081 (N_28081,N_27473,N_27535);
xor U28082 (N_28082,N_27138,N_27399);
and U28083 (N_28083,N_27386,N_27872);
and U28084 (N_28084,N_27074,N_27298);
xnor U28085 (N_28085,N_27150,N_27530);
xnor U28086 (N_28086,N_27198,N_27489);
and U28087 (N_28087,N_27385,N_27659);
or U28088 (N_28088,N_27475,N_27359);
xor U28089 (N_28089,N_27302,N_27667);
or U28090 (N_28090,N_27913,N_27604);
nand U28091 (N_28091,N_27270,N_27184);
nand U28092 (N_28092,N_27387,N_27042);
or U28093 (N_28093,N_27804,N_27341);
nand U28094 (N_28094,N_27776,N_27722);
xor U28095 (N_28095,N_27334,N_27773);
nor U28096 (N_28096,N_27153,N_27937);
xor U28097 (N_28097,N_27264,N_27720);
or U28098 (N_28098,N_27700,N_27633);
nand U28099 (N_28099,N_27938,N_27444);
nor U28100 (N_28100,N_27591,N_27205);
or U28101 (N_28101,N_27612,N_27891);
and U28102 (N_28102,N_27561,N_27170);
and U28103 (N_28103,N_27449,N_27336);
or U28104 (N_28104,N_27799,N_27297);
or U28105 (N_28105,N_27164,N_27274);
and U28106 (N_28106,N_27551,N_27424);
or U28107 (N_28107,N_27037,N_27998);
or U28108 (N_28108,N_27517,N_27646);
nand U28109 (N_28109,N_27677,N_27963);
xor U28110 (N_28110,N_27206,N_27490);
xor U28111 (N_28111,N_27865,N_27689);
or U28112 (N_28112,N_27541,N_27193);
nand U28113 (N_28113,N_27803,N_27089);
nand U28114 (N_28114,N_27212,N_27163);
or U28115 (N_28115,N_27571,N_27048);
and U28116 (N_28116,N_27976,N_27566);
nor U28117 (N_28117,N_27560,N_27770);
nor U28118 (N_28118,N_27213,N_27145);
nand U28119 (N_28119,N_27239,N_27234);
nor U28120 (N_28120,N_27967,N_27639);
nand U28121 (N_28121,N_27820,N_27012);
nand U28122 (N_28122,N_27196,N_27645);
xor U28123 (N_28123,N_27115,N_27534);
xnor U28124 (N_28124,N_27039,N_27290);
and U28125 (N_28125,N_27031,N_27190);
nand U28126 (N_28126,N_27769,N_27786);
and U28127 (N_28127,N_27391,N_27884);
or U28128 (N_28128,N_27142,N_27846);
nor U28129 (N_28129,N_27252,N_27331);
nand U28130 (N_28130,N_27179,N_27249);
or U28131 (N_28131,N_27407,N_27388);
xnor U28132 (N_28132,N_27258,N_27956);
nand U28133 (N_28133,N_27590,N_27814);
nor U28134 (N_28134,N_27093,N_27901);
and U28135 (N_28135,N_27343,N_27169);
nand U28136 (N_28136,N_27311,N_27735);
xnor U28137 (N_28137,N_27706,N_27296);
xnor U28138 (N_28138,N_27127,N_27925);
or U28139 (N_28139,N_27580,N_27136);
xnor U28140 (N_28140,N_27791,N_27357);
xor U28141 (N_28141,N_27166,N_27800);
nand U28142 (N_28142,N_27632,N_27006);
xor U28143 (N_28143,N_27670,N_27630);
nor U28144 (N_28144,N_27669,N_27842);
or U28145 (N_28145,N_27191,N_27420);
and U28146 (N_28146,N_27469,N_27148);
and U28147 (N_28147,N_27918,N_27417);
xnor U28148 (N_28148,N_27027,N_27299);
or U28149 (N_28149,N_27360,N_27232);
nor U28150 (N_28150,N_27509,N_27464);
xor U28151 (N_28151,N_27873,N_27143);
xor U28152 (N_28152,N_27477,N_27347);
xnor U28153 (N_28153,N_27396,N_27986);
xor U28154 (N_28154,N_27739,N_27226);
nor U28155 (N_28155,N_27924,N_27358);
and U28156 (N_28156,N_27838,N_27466);
or U28157 (N_28157,N_27055,N_27459);
and U28158 (N_28158,N_27949,N_27716);
or U28159 (N_28159,N_27369,N_27970);
or U28160 (N_28160,N_27980,N_27684);
and U28161 (N_28161,N_27756,N_27500);
and U28162 (N_28162,N_27759,N_27026);
nand U28163 (N_28163,N_27187,N_27279);
and U28164 (N_28164,N_27428,N_27114);
nor U28165 (N_28165,N_27702,N_27810);
nor U28166 (N_28166,N_27581,N_27168);
or U28167 (N_28167,N_27040,N_27413);
nor U28168 (N_28168,N_27122,N_27723);
and U28169 (N_28169,N_27961,N_27613);
nor U28170 (N_28170,N_27476,N_27642);
and U28171 (N_28171,N_27130,N_27342);
xnor U28172 (N_28172,N_27392,N_27332);
xnor U28173 (N_28173,N_27217,N_27103);
or U28174 (N_28174,N_27817,N_27917);
nand U28175 (N_28175,N_27960,N_27194);
xnor U28176 (N_28176,N_27935,N_27394);
and U28177 (N_28177,N_27079,N_27415);
or U28178 (N_28178,N_27727,N_27618);
or U28179 (N_28179,N_27410,N_27044);
nand U28180 (N_28180,N_27932,N_27251);
and U28181 (N_28181,N_27660,N_27460);
xor U28182 (N_28182,N_27403,N_27615);
nand U28183 (N_28183,N_27273,N_27755);
and U28184 (N_28184,N_27705,N_27724);
and U28185 (N_28185,N_27875,N_27317);
nand U28186 (N_28186,N_27300,N_27758);
xor U28187 (N_28187,N_27906,N_27260);
xnor U28188 (N_28188,N_27091,N_27698);
xor U28189 (N_28189,N_27439,N_27313);
xnor U28190 (N_28190,N_27244,N_27871);
or U28191 (N_28191,N_27805,N_27003);
and U28192 (N_28192,N_27465,N_27186);
xor U28193 (N_28193,N_27761,N_27374);
xor U28194 (N_28194,N_27643,N_27209);
and U28195 (N_28195,N_27774,N_27515);
or U28196 (N_28196,N_27207,N_27866);
nor U28197 (N_28197,N_27876,N_27454);
and U28198 (N_28198,N_27537,N_27741);
or U28199 (N_28199,N_27679,N_27697);
nand U28200 (N_28200,N_27533,N_27909);
or U28201 (N_28201,N_27507,N_27118);
and U28202 (N_28202,N_27208,N_27216);
or U28203 (N_28203,N_27492,N_27408);
or U28204 (N_28204,N_27080,N_27324);
xor U28205 (N_28205,N_27100,N_27033);
or U28206 (N_28206,N_27458,N_27174);
xor U28207 (N_28207,N_27614,N_27071);
and U28208 (N_28208,N_27144,N_27231);
and U28209 (N_28209,N_27120,N_27000);
or U28210 (N_28210,N_27220,N_27808);
xor U28211 (N_28211,N_27141,N_27893);
nand U28212 (N_28212,N_27729,N_27943);
nand U28213 (N_28213,N_27671,N_27811);
nand U28214 (N_28214,N_27072,N_27362);
nand U28215 (N_28215,N_27050,N_27763);
xor U28216 (N_28216,N_27063,N_27018);
and U28217 (N_28217,N_27955,N_27856);
nor U28218 (N_28218,N_27885,N_27688);
nand U28219 (N_28219,N_27076,N_27227);
and U28220 (N_28220,N_27546,N_27105);
xnor U28221 (N_28221,N_27953,N_27984);
and U28222 (N_28222,N_27390,N_27339);
xnor U28223 (N_28223,N_27588,N_27266);
xor U28224 (N_28224,N_27243,N_27121);
nor U28225 (N_28225,N_27672,N_27096);
xor U28226 (N_28226,N_27538,N_27809);
nor U28227 (N_28227,N_27372,N_27529);
or U28228 (N_28228,N_27545,N_27847);
nand U28229 (N_28229,N_27276,N_27825);
nand U28230 (N_28230,N_27738,N_27095);
or U28231 (N_28231,N_27572,N_27032);
nand U28232 (N_28232,N_27487,N_27034);
xnor U28233 (N_28233,N_27526,N_27898);
xor U28234 (N_28234,N_27482,N_27330);
nor U28235 (N_28235,N_27664,N_27067);
nor U28236 (N_28236,N_27112,N_27165);
xor U28237 (N_28237,N_27092,N_27363);
and U28238 (N_28238,N_27951,N_27287);
and U28239 (N_28239,N_27557,N_27952);
xor U28240 (N_28240,N_27429,N_27889);
and U28241 (N_28241,N_27839,N_27223);
xor U28242 (N_28242,N_27499,N_27964);
xnor U28243 (N_28243,N_27802,N_27023);
nand U28244 (N_28244,N_27576,N_27395);
and U28245 (N_28245,N_27995,N_27008);
and U28246 (N_28246,N_27446,N_27430);
and U28247 (N_28247,N_27201,N_27286);
nand U28248 (N_28248,N_27292,N_27478);
or U28249 (N_28249,N_27694,N_27954);
xnor U28250 (N_28250,N_27676,N_27125);
xnor U28251 (N_28251,N_27860,N_27222);
nor U28252 (N_28252,N_27349,N_27367);
and U28253 (N_28253,N_27853,N_27886);
or U28254 (N_28254,N_27764,N_27868);
nor U28255 (N_28255,N_27389,N_27807);
nor U28256 (N_28256,N_27278,N_27238);
xnor U28257 (N_28257,N_27214,N_27237);
and U28258 (N_28258,N_27707,N_27215);
nor U28259 (N_28259,N_27277,N_27747);
xor U28260 (N_28260,N_27760,N_27161);
xnor U28261 (N_28261,N_27301,N_27861);
and U28262 (N_28262,N_27229,N_27472);
nor U28263 (N_28263,N_27975,N_27542);
and U28264 (N_28264,N_27611,N_27199);
xnor U28265 (N_28265,N_27793,N_27990);
or U28266 (N_28266,N_27991,N_27516);
nor U28267 (N_28267,N_27519,N_27987);
and U28268 (N_28268,N_27176,N_27874);
xor U28269 (N_28269,N_27593,N_27177);
nand U28270 (N_28270,N_27470,N_27532);
nor U28271 (N_28271,N_27896,N_27558);
and U28272 (N_28272,N_27307,N_27432);
xnor U28273 (N_28273,N_27109,N_27253);
nand U28274 (N_28274,N_27171,N_27731);
and U28275 (N_28275,N_27441,N_27514);
nor U28276 (N_28276,N_27275,N_27480);
xnor U28277 (N_28277,N_27704,N_27058);
and U28278 (N_28278,N_27921,N_27745);
and U28279 (N_28279,N_27978,N_27725);
and U28280 (N_28280,N_27728,N_27652);
nand U28281 (N_28281,N_27965,N_27864);
xor U28282 (N_28282,N_27246,N_27375);
and U28283 (N_28283,N_27353,N_27831);
or U28284 (N_28284,N_27834,N_27795);
or U28285 (N_28285,N_27308,N_27682);
and U28286 (N_28286,N_27895,N_27036);
nor U28287 (N_28287,N_27457,N_27314);
nand U28288 (N_28288,N_27543,N_27748);
xnor U28289 (N_28289,N_27054,N_27378);
or U28290 (N_28290,N_27491,N_27583);
xor U28291 (N_28291,N_27502,N_27319);
nor U28292 (N_28292,N_27564,N_27106);
nor U28293 (N_28293,N_27573,N_27303);
nand U28294 (N_28294,N_27992,N_27011);
nor U28295 (N_28295,N_27099,N_27321);
nor U28296 (N_28296,N_27379,N_27870);
or U28297 (N_28297,N_27597,N_27948);
nand U28298 (N_28298,N_27754,N_27592);
nand U28299 (N_28299,N_27610,N_27325);
or U28300 (N_28300,N_27090,N_27059);
nor U28301 (N_28301,N_27923,N_27129);
xor U28302 (N_28302,N_27732,N_27878);
nand U28303 (N_28303,N_27282,N_27073);
nand U28304 (N_28304,N_27128,N_27159);
nor U28305 (N_28305,N_27736,N_27155);
or U28306 (N_28306,N_27708,N_27440);
nor U28307 (N_28307,N_27488,N_27124);
nand U28308 (N_28308,N_27930,N_27204);
nor U28309 (N_28309,N_27843,N_27972);
nor U28310 (N_28310,N_27046,N_27765);
and U28311 (N_28311,N_27579,N_27711);
or U28312 (N_28312,N_27827,N_27233);
xnor U28313 (N_28313,N_27348,N_27346);
nand U28314 (N_28314,N_27550,N_27709);
and U28315 (N_28315,N_27981,N_27971);
nand U28316 (N_28316,N_27994,N_27219);
or U28317 (N_28317,N_27047,N_27695);
nand U28318 (N_28318,N_27848,N_27426);
xnor U28319 (N_28319,N_27173,N_27456);
xnor U28320 (N_28320,N_27484,N_27146);
and U28321 (N_28321,N_27656,N_27240);
nand U28322 (N_28322,N_27402,N_27351);
nor U28323 (N_28323,N_27520,N_27376);
or U28324 (N_28324,N_27180,N_27154);
and U28325 (N_28325,N_27915,N_27431);
nor U28326 (N_28326,N_27366,N_27830);
or U28327 (N_28327,N_27202,N_27826);
and U28328 (N_28328,N_27268,N_27340);
nand U28329 (N_28329,N_27119,N_27057);
or U28330 (N_28330,N_27719,N_27352);
nor U28331 (N_28331,N_27197,N_27328);
nand U28332 (N_28332,N_27203,N_27691);
or U28333 (N_28333,N_27785,N_27600);
nand U28334 (N_28334,N_27030,N_27380);
nand U28335 (N_28335,N_27294,N_27690);
xnor U28336 (N_28336,N_27017,N_27787);
xnor U28337 (N_28337,N_27433,N_27855);
nand U28338 (N_28338,N_27966,N_27242);
xnor U28339 (N_28339,N_27910,N_27609);
nor U28340 (N_28340,N_27595,N_27133);
and U28341 (N_28341,N_27772,N_27988);
and U28342 (N_28342,N_27383,N_27070);
and U28343 (N_28343,N_27920,N_27225);
nor U28344 (N_28344,N_27060,N_27200);
nand U28345 (N_28345,N_27002,N_27796);
and U28346 (N_28346,N_27685,N_27559);
nand U28347 (N_28347,N_27422,N_27683);
or U28348 (N_28348,N_27117,N_27162);
nand U28349 (N_28349,N_27696,N_27195);
and U28350 (N_28350,N_27427,N_27624);
and U28351 (N_28351,N_27160,N_27254);
xnor U28352 (N_28352,N_27897,N_27069);
nor U28353 (N_28353,N_27554,N_27405);
nand U28354 (N_28354,N_27350,N_27734);
nor U28355 (N_28355,N_27657,N_27781);
or U28356 (N_28356,N_27288,N_27644);
and U28357 (N_28357,N_27255,N_27944);
nand U28358 (N_28358,N_27053,N_27056);
or U28359 (N_28359,N_27108,N_27940);
and U28360 (N_28360,N_27468,N_27250);
xnor U28361 (N_28361,N_27936,N_27653);
nor U28362 (N_28362,N_27859,N_27043);
or U28363 (N_28363,N_27518,N_27625);
xnor U28364 (N_28364,N_27790,N_27649);
and U28365 (N_28365,N_27354,N_27863);
nand U28366 (N_28366,N_27962,N_27436);
and U28367 (N_28367,N_27263,N_27766);
or U28368 (N_28368,N_27483,N_27086);
nor U28369 (N_28369,N_27007,N_27510);
nand U28370 (N_28370,N_27293,N_27211);
or U28371 (N_28371,N_27448,N_27445);
nor U28372 (N_28372,N_27281,N_27261);
nor U28373 (N_28373,N_27447,N_27524);
and U28374 (N_28374,N_27730,N_27102);
nor U28375 (N_28375,N_27381,N_27167);
nand U28376 (N_28376,N_27271,N_27904);
nor U28377 (N_28377,N_27495,N_27686);
or U28378 (N_28378,N_27703,N_27064);
nand U28379 (N_28379,N_27742,N_27323);
xor U28380 (N_28380,N_27345,N_27461);
and U28381 (N_28381,N_27957,N_27585);
or U28382 (N_28382,N_27005,N_27015);
xnor U28383 (N_28383,N_27844,N_27152);
nor U28384 (N_28384,N_27455,N_27029);
xor U28385 (N_28385,N_27852,N_27467);
and U28386 (N_28386,N_27934,N_27327);
and U28387 (N_28387,N_27567,N_27806);
nor U28388 (N_28388,N_27914,N_27158);
and U28389 (N_28389,N_27009,N_27589);
and U28390 (N_28390,N_27563,N_27568);
nand U28391 (N_28391,N_27061,N_27794);
nand U28392 (N_28392,N_27540,N_27905);
nand U28393 (N_28393,N_27979,N_27587);
or U28394 (N_28394,N_27647,N_27051);
nand U28395 (N_28395,N_27549,N_27398);
or U28396 (N_28396,N_27224,N_27552);
and U28397 (N_28397,N_27210,N_27295);
nand U28398 (N_28398,N_27767,N_27779);
and U28399 (N_28399,N_27635,N_27084);
nor U28400 (N_28400,N_27370,N_27621);
nor U28401 (N_28401,N_27792,N_27123);
nand U28402 (N_28402,N_27337,N_27680);
or U28403 (N_28403,N_27974,N_27437);
nor U28404 (N_28404,N_27662,N_27620);
nand U28405 (N_28405,N_27361,N_27434);
xor U28406 (N_28406,N_27326,N_27718);
and U28407 (N_28407,N_27304,N_27692);
xnor U28408 (N_28408,N_27182,N_27021);
nand U28409 (N_28409,N_27740,N_27983);
nand U28410 (N_28410,N_27185,N_27024);
or U28411 (N_28411,N_27485,N_27753);
and U28412 (N_28412,N_27539,N_27025);
or U28413 (N_28413,N_27401,N_27661);
and U28414 (N_28414,N_27183,N_27265);
or U28415 (N_28415,N_27259,N_27775);
nor U28416 (N_28416,N_27305,N_27312);
or U28417 (N_28417,N_27836,N_27235);
nor U28418 (N_28418,N_27368,N_27486);
xor U28419 (N_28419,N_27584,N_27916);
xor U28420 (N_28420,N_27527,N_27926);
nand U28421 (N_28421,N_27819,N_27578);
nand U28422 (N_28422,N_27712,N_27245);
xor U28423 (N_28423,N_27824,N_27840);
or U28424 (N_28424,N_27149,N_27617);
nand U28425 (N_28425,N_27463,N_27912);
xor U28426 (N_28426,N_27098,N_27188);
or U28427 (N_28427,N_27681,N_27907);
or U28428 (N_28428,N_27801,N_27945);
nor U28429 (N_28429,N_27513,N_27022);
xor U28430 (N_28430,N_27999,N_27316);
nor U28431 (N_28431,N_27020,N_27147);
or U28432 (N_28432,N_27355,N_27890);
and U28433 (N_28433,N_27028,N_27762);
nor U28434 (N_28434,N_27812,N_27902);
xor U28435 (N_28435,N_27877,N_27668);
xor U28436 (N_28436,N_27784,N_27751);
or U28437 (N_28437,N_27869,N_27156);
and U28438 (N_28438,N_27525,N_27778);
or U28439 (N_28439,N_27075,N_27384);
and U28440 (N_28440,N_27481,N_27713);
and U28441 (N_28441,N_27997,N_27110);
nor U28442 (N_28442,N_27687,N_27746);
and U28443 (N_28443,N_27139,N_27523);
nand U28444 (N_28444,N_27335,N_27989);
xor U28445 (N_28445,N_27821,N_27097);
nand U28446 (N_28446,N_27973,N_27931);
or U28447 (N_28447,N_27622,N_27977);
nand U28448 (N_28448,N_27750,N_27879);
nor U28449 (N_28449,N_27536,N_27888);
and U28450 (N_28450,N_27151,N_27862);
nand U28451 (N_28451,N_27178,N_27333);
nand U28452 (N_28452,N_27175,N_27813);
and U28453 (N_28453,N_27318,N_27016);
and U28454 (N_28454,N_27947,N_27262);
or U28455 (N_28455,N_27406,N_27280);
and U28456 (N_28456,N_27882,N_27929);
and U28457 (N_28457,N_27586,N_27638);
xor U28458 (N_28458,N_27505,N_27797);
and U28459 (N_28459,N_27626,N_27911);
xor U28460 (N_28460,N_27922,N_27014);
or U28461 (N_28461,N_27715,N_27623);
xor U28462 (N_28462,N_27602,N_27364);
xnor U28463 (N_28463,N_27062,N_27654);
nand U28464 (N_28464,N_27555,N_27442);
and U28465 (N_28465,N_27783,N_27289);
and U28466 (N_28466,N_27126,N_27257);
xor U28467 (N_28467,N_27065,N_27113);
and U28468 (N_28468,N_27104,N_27315);
xnor U28469 (N_28469,N_27101,N_27833);
and U28470 (N_28470,N_27627,N_27928);
nor U28471 (N_28471,N_27969,N_27556);
xnor U28472 (N_28472,N_27137,N_27880);
and U28473 (N_28473,N_27837,N_27939);
or U28474 (N_28474,N_27356,N_27908);
nor U28475 (N_28475,N_27001,N_27450);
and U28476 (N_28476,N_27857,N_27283);
or U28477 (N_28477,N_27640,N_27605);
nand U28478 (N_28478,N_27498,N_27714);
and U28479 (N_28479,N_27400,N_27854);
nor U28480 (N_28480,N_27919,N_27818);
nor U28481 (N_28481,N_27256,N_27425);
nand U28482 (N_28482,N_27382,N_27267);
or U28483 (N_28483,N_27248,N_27085);
nand U28484 (N_28484,N_27443,N_27094);
nor U28485 (N_28485,N_27041,N_27606);
nand U28486 (N_28486,N_27189,N_27823);
and U28487 (N_28487,N_27228,N_27272);
nor U28488 (N_28488,N_27899,N_27768);
nand U28489 (N_28489,N_27985,N_27743);
nand U28490 (N_28490,N_27131,N_27757);
or U28491 (N_28491,N_27371,N_27616);
or U28492 (N_28492,N_27107,N_27521);
nor U28493 (N_28493,N_27607,N_27512);
or U28494 (N_28494,N_27013,N_27414);
nand U28495 (N_28495,N_27479,N_27982);
xor U28496 (N_28496,N_27851,N_27582);
nor U28497 (N_28497,N_27019,N_27798);
or U28498 (N_28498,N_27636,N_27230);
and U28499 (N_28499,N_27894,N_27631);
and U28500 (N_28500,N_27499,N_27873);
nand U28501 (N_28501,N_27173,N_27189);
xor U28502 (N_28502,N_27315,N_27390);
and U28503 (N_28503,N_27303,N_27803);
or U28504 (N_28504,N_27924,N_27771);
and U28505 (N_28505,N_27626,N_27343);
nand U28506 (N_28506,N_27953,N_27707);
nand U28507 (N_28507,N_27149,N_27571);
nor U28508 (N_28508,N_27574,N_27507);
nor U28509 (N_28509,N_27300,N_27099);
and U28510 (N_28510,N_27274,N_27158);
and U28511 (N_28511,N_27148,N_27957);
nor U28512 (N_28512,N_27961,N_27953);
xnor U28513 (N_28513,N_27260,N_27242);
xor U28514 (N_28514,N_27002,N_27280);
nand U28515 (N_28515,N_27409,N_27827);
or U28516 (N_28516,N_27727,N_27155);
and U28517 (N_28517,N_27610,N_27409);
or U28518 (N_28518,N_27263,N_27465);
and U28519 (N_28519,N_27654,N_27866);
and U28520 (N_28520,N_27355,N_27914);
nand U28521 (N_28521,N_27535,N_27612);
or U28522 (N_28522,N_27073,N_27745);
nand U28523 (N_28523,N_27368,N_27641);
and U28524 (N_28524,N_27417,N_27508);
nand U28525 (N_28525,N_27075,N_27317);
xnor U28526 (N_28526,N_27879,N_27135);
or U28527 (N_28527,N_27650,N_27258);
or U28528 (N_28528,N_27023,N_27582);
xnor U28529 (N_28529,N_27512,N_27587);
xnor U28530 (N_28530,N_27799,N_27724);
and U28531 (N_28531,N_27835,N_27547);
xor U28532 (N_28532,N_27841,N_27108);
and U28533 (N_28533,N_27126,N_27526);
or U28534 (N_28534,N_27094,N_27973);
or U28535 (N_28535,N_27440,N_27125);
or U28536 (N_28536,N_27107,N_27154);
or U28537 (N_28537,N_27727,N_27426);
nor U28538 (N_28538,N_27256,N_27953);
nand U28539 (N_28539,N_27297,N_27795);
nand U28540 (N_28540,N_27730,N_27195);
or U28541 (N_28541,N_27850,N_27931);
and U28542 (N_28542,N_27004,N_27096);
nor U28543 (N_28543,N_27231,N_27480);
or U28544 (N_28544,N_27554,N_27189);
and U28545 (N_28545,N_27955,N_27973);
or U28546 (N_28546,N_27648,N_27155);
and U28547 (N_28547,N_27573,N_27397);
nor U28548 (N_28548,N_27148,N_27443);
nand U28549 (N_28549,N_27707,N_27353);
nor U28550 (N_28550,N_27118,N_27580);
nor U28551 (N_28551,N_27848,N_27955);
or U28552 (N_28552,N_27977,N_27604);
and U28553 (N_28553,N_27237,N_27381);
and U28554 (N_28554,N_27897,N_27713);
xnor U28555 (N_28555,N_27487,N_27397);
xor U28556 (N_28556,N_27347,N_27446);
and U28557 (N_28557,N_27189,N_27983);
nand U28558 (N_28558,N_27906,N_27967);
or U28559 (N_28559,N_27409,N_27301);
or U28560 (N_28560,N_27372,N_27844);
or U28561 (N_28561,N_27274,N_27285);
nand U28562 (N_28562,N_27043,N_27770);
xnor U28563 (N_28563,N_27524,N_27939);
and U28564 (N_28564,N_27603,N_27134);
and U28565 (N_28565,N_27783,N_27070);
xor U28566 (N_28566,N_27670,N_27012);
nor U28567 (N_28567,N_27375,N_27225);
and U28568 (N_28568,N_27115,N_27852);
nor U28569 (N_28569,N_27658,N_27730);
xnor U28570 (N_28570,N_27080,N_27682);
or U28571 (N_28571,N_27555,N_27190);
and U28572 (N_28572,N_27639,N_27813);
nand U28573 (N_28573,N_27204,N_27513);
or U28574 (N_28574,N_27700,N_27543);
or U28575 (N_28575,N_27795,N_27758);
and U28576 (N_28576,N_27267,N_27355);
or U28577 (N_28577,N_27466,N_27159);
nor U28578 (N_28578,N_27909,N_27654);
nand U28579 (N_28579,N_27112,N_27801);
nor U28580 (N_28580,N_27004,N_27626);
nand U28581 (N_28581,N_27448,N_27822);
nand U28582 (N_28582,N_27250,N_27052);
nand U28583 (N_28583,N_27533,N_27658);
nand U28584 (N_28584,N_27950,N_27333);
and U28585 (N_28585,N_27036,N_27690);
xor U28586 (N_28586,N_27080,N_27895);
or U28587 (N_28587,N_27824,N_27549);
and U28588 (N_28588,N_27175,N_27391);
and U28589 (N_28589,N_27414,N_27293);
nand U28590 (N_28590,N_27313,N_27490);
and U28591 (N_28591,N_27299,N_27786);
nand U28592 (N_28592,N_27887,N_27635);
and U28593 (N_28593,N_27784,N_27916);
nand U28594 (N_28594,N_27758,N_27343);
nand U28595 (N_28595,N_27690,N_27515);
xor U28596 (N_28596,N_27236,N_27475);
and U28597 (N_28597,N_27087,N_27250);
and U28598 (N_28598,N_27912,N_27592);
and U28599 (N_28599,N_27155,N_27372);
and U28600 (N_28600,N_27160,N_27706);
nor U28601 (N_28601,N_27540,N_27338);
nand U28602 (N_28602,N_27141,N_27494);
nand U28603 (N_28603,N_27167,N_27676);
and U28604 (N_28604,N_27076,N_27841);
xnor U28605 (N_28605,N_27131,N_27076);
and U28606 (N_28606,N_27186,N_27481);
xor U28607 (N_28607,N_27257,N_27292);
xor U28608 (N_28608,N_27402,N_27669);
or U28609 (N_28609,N_27759,N_27652);
xnor U28610 (N_28610,N_27976,N_27691);
and U28611 (N_28611,N_27906,N_27747);
nand U28612 (N_28612,N_27183,N_27474);
or U28613 (N_28613,N_27488,N_27920);
and U28614 (N_28614,N_27362,N_27471);
xnor U28615 (N_28615,N_27307,N_27403);
nand U28616 (N_28616,N_27662,N_27891);
or U28617 (N_28617,N_27721,N_27503);
and U28618 (N_28618,N_27044,N_27842);
nand U28619 (N_28619,N_27247,N_27278);
or U28620 (N_28620,N_27408,N_27782);
or U28621 (N_28621,N_27198,N_27100);
xnor U28622 (N_28622,N_27792,N_27711);
and U28623 (N_28623,N_27987,N_27817);
xor U28624 (N_28624,N_27638,N_27511);
nand U28625 (N_28625,N_27056,N_27007);
nand U28626 (N_28626,N_27759,N_27280);
or U28627 (N_28627,N_27812,N_27515);
and U28628 (N_28628,N_27104,N_27339);
or U28629 (N_28629,N_27826,N_27057);
or U28630 (N_28630,N_27821,N_27001);
or U28631 (N_28631,N_27133,N_27237);
nand U28632 (N_28632,N_27718,N_27857);
xnor U28633 (N_28633,N_27894,N_27355);
or U28634 (N_28634,N_27267,N_27142);
nor U28635 (N_28635,N_27644,N_27601);
or U28636 (N_28636,N_27744,N_27149);
and U28637 (N_28637,N_27557,N_27463);
and U28638 (N_28638,N_27693,N_27459);
or U28639 (N_28639,N_27226,N_27190);
nor U28640 (N_28640,N_27744,N_27443);
nor U28641 (N_28641,N_27126,N_27366);
and U28642 (N_28642,N_27221,N_27174);
or U28643 (N_28643,N_27994,N_27725);
nor U28644 (N_28644,N_27183,N_27948);
nor U28645 (N_28645,N_27040,N_27322);
xor U28646 (N_28646,N_27119,N_27978);
nand U28647 (N_28647,N_27230,N_27014);
or U28648 (N_28648,N_27372,N_27700);
xor U28649 (N_28649,N_27452,N_27090);
and U28650 (N_28650,N_27994,N_27756);
xnor U28651 (N_28651,N_27743,N_27739);
nor U28652 (N_28652,N_27866,N_27847);
nand U28653 (N_28653,N_27233,N_27440);
nor U28654 (N_28654,N_27114,N_27288);
nand U28655 (N_28655,N_27758,N_27372);
xor U28656 (N_28656,N_27037,N_27587);
or U28657 (N_28657,N_27739,N_27942);
or U28658 (N_28658,N_27365,N_27668);
nand U28659 (N_28659,N_27752,N_27535);
nand U28660 (N_28660,N_27641,N_27418);
xor U28661 (N_28661,N_27060,N_27011);
xor U28662 (N_28662,N_27858,N_27400);
or U28663 (N_28663,N_27148,N_27401);
xnor U28664 (N_28664,N_27483,N_27775);
xnor U28665 (N_28665,N_27683,N_27662);
nand U28666 (N_28666,N_27093,N_27711);
xor U28667 (N_28667,N_27575,N_27326);
nor U28668 (N_28668,N_27439,N_27142);
nor U28669 (N_28669,N_27990,N_27223);
and U28670 (N_28670,N_27698,N_27726);
nand U28671 (N_28671,N_27146,N_27691);
and U28672 (N_28672,N_27139,N_27901);
nor U28673 (N_28673,N_27126,N_27398);
nor U28674 (N_28674,N_27315,N_27269);
nand U28675 (N_28675,N_27104,N_27882);
xor U28676 (N_28676,N_27265,N_27021);
xor U28677 (N_28677,N_27631,N_27968);
and U28678 (N_28678,N_27694,N_27915);
or U28679 (N_28679,N_27947,N_27888);
nor U28680 (N_28680,N_27589,N_27364);
nor U28681 (N_28681,N_27744,N_27412);
and U28682 (N_28682,N_27741,N_27043);
and U28683 (N_28683,N_27211,N_27659);
nand U28684 (N_28684,N_27053,N_27843);
or U28685 (N_28685,N_27628,N_27017);
nor U28686 (N_28686,N_27634,N_27523);
nand U28687 (N_28687,N_27247,N_27969);
and U28688 (N_28688,N_27551,N_27129);
xor U28689 (N_28689,N_27496,N_27781);
or U28690 (N_28690,N_27188,N_27833);
or U28691 (N_28691,N_27788,N_27641);
nand U28692 (N_28692,N_27314,N_27786);
and U28693 (N_28693,N_27681,N_27000);
nand U28694 (N_28694,N_27953,N_27352);
xnor U28695 (N_28695,N_27035,N_27737);
nand U28696 (N_28696,N_27263,N_27850);
or U28697 (N_28697,N_27380,N_27884);
nor U28698 (N_28698,N_27886,N_27334);
nand U28699 (N_28699,N_27596,N_27103);
xnor U28700 (N_28700,N_27986,N_27924);
nand U28701 (N_28701,N_27364,N_27990);
xor U28702 (N_28702,N_27269,N_27876);
or U28703 (N_28703,N_27173,N_27894);
nand U28704 (N_28704,N_27560,N_27767);
nor U28705 (N_28705,N_27469,N_27346);
nand U28706 (N_28706,N_27667,N_27950);
or U28707 (N_28707,N_27758,N_27428);
nor U28708 (N_28708,N_27282,N_27261);
and U28709 (N_28709,N_27431,N_27881);
nor U28710 (N_28710,N_27364,N_27959);
xnor U28711 (N_28711,N_27662,N_27048);
or U28712 (N_28712,N_27741,N_27708);
and U28713 (N_28713,N_27699,N_27902);
nor U28714 (N_28714,N_27454,N_27141);
nand U28715 (N_28715,N_27792,N_27212);
nor U28716 (N_28716,N_27813,N_27149);
or U28717 (N_28717,N_27423,N_27238);
nor U28718 (N_28718,N_27586,N_27629);
nand U28719 (N_28719,N_27242,N_27726);
xnor U28720 (N_28720,N_27880,N_27837);
and U28721 (N_28721,N_27263,N_27401);
nand U28722 (N_28722,N_27307,N_27786);
xnor U28723 (N_28723,N_27756,N_27391);
and U28724 (N_28724,N_27403,N_27205);
xor U28725 (N_28725,N_27920,N_27027);
xor U28726 (N_28726,N_27716,N_27313);
nor U28727 (N_28727,N_27864,N_27068);
nor U28728 (N_28728,N_27941,N_27270);
nand U28729 (N_28729,N_27179,N_27214);
or U28730 (N_28730,N_27246,N_27871);
or U28731 (N_28731,N_27445,N_27876);
nand U28732 (N_28732,N_27858,N_27448);
and U28733 (N_28733,N_27310,N_27709);
nor U28734 (N_28734,N_27957,N_27767);
nor U28735 (N_28735,N_27335,N_27558);
nor U28736 (N_28736,N_27591,N_27124);
nor U28737 (N_28737,N_27131,N_27305);
xor U28738 (N_28738,N_27201,N_27445);
and U28739 (N_28739,N_27102,N_27132);
nand U28740 (N_28740,N_27981,N_27829);
xnor U28741 (N_28741,N_27543,N_27696);
xnor U28742 (N_28742,N_27758,N_27321);
nor U28743 (N_28743,N_27822,N_27922);
xor U28744 (N_28744,N_27696,N_27128);
nor U28745 (N_28745,N_27628,N_27082);
nand U28746 (N_28746,N_27448,N_27129);
xnor U28747 (N_28747,N_27353,N_27307);
xnor U28748 (N_28748,N_27930,N_27015);
nand U28749 (N_28749,N_27920,N_27306);
nor U28750 (N_28750,N_27204,N_27364);
or U28751 (N_28751,N_27765,N_27535);
xnor U28752 (N_28752,N_27995,N_27896);
or U28753 (N_28753,N_27709,N_27201);
and U28754 (N_28754,N_27167,N_27410);
nor U28755 (N_28755,N_27528,N_27079);
nand U28756 (N_28756,N_27856,N_27282);
nand U28757 (N_28757,N_27983,N_27118);
or U28758 (N_28758,N_27186,N_27033);
nor U28759 (N_28759,N_27649,N_27915);
or U28760 (N_28760,N_27831,N_27425);
xor U28761 (N_28761,N_27555,N_27112);
nand U28762 (N_28762,N_27480,N_27737);
nand U28763 (N_28763,N_27483,N_27508);
xnor U28764 (N_28764,N_27734,N_27959);
nand U28765 (N_28765,N_27984,N_27754);
nor U28766 (N_28766,N_27986,N_27697);
nand U28767 (N_28767,N_27240,N_27276);
or U28768 (N_28768,N_27411,N_27708);
nand U28769 (N_28769,N_27314,N_27615);
or U28770 (N_28770,N_27294,N_27729);
xor U28771 (N_28771,N_27879,N_27783);
xnor U28772 (N_28772,N_27876,N_27455);
and U28773 (N_28773,N_27269,N_27650);
nand U28774 (N_28774,N_27974,N_27232);
nor U28775 (N_28775,N_27575,N_27981);
nor U28776 (N_28776,N_27881,N_27010);
xnor U28777 (N_28777,N_27725,N_27457);
nand U28778 (N_28778,N_27466,N_27574);
nor U28779 (N_28779,N_27497,N_27159);
nor U28780 (N_28780,N_27550,N_27478);
or U28781 (N_28781,N_27455,N_27697);
nand U28782 (N_28782,N_27121,N_27701);
nand U28783 (N_28783,N_27434,N_27053);
and U28784 (N_28784,N_27067,N_27735);
and U28785 (N_28785,N_27958,N_27441);
nand U28786 (N_28786,N_27318,N_27932);
nand U28787 (N_28787,N_27434,N_27293);
nor U28788 (N_28788,N_27492,N_27679);
and U28789 (N_28789,N_27887,N_27195);
nand U28790 (N_28790,N_27926,N_27015);
xor U28791 (N_28791,N_27233,N_27788);
xnor U28792 (N_28792,N_27549,N_27048);
xor U28793 (N_28793,N_27153,N_27336);
nor U28794 (N_28794,N_27655,N_27074);
or U28795 (N_28795,N_27279,N_27643);
xnor U28796 (N_28796,N_27251,N_27500);
and U28797 (N_28797,N_27912,N_27356);
and U28798 (N_28798,N_27402,N_27628);
or U28799 (N_28799,N_27538,N_27096);
xor U28800 (N_28800,N_27825,N_27288);
xnor U28801 (N_28801,N_27160,N_27623);
and U28802 (N_28802,N_27878,N_27128);
xor U28803 (N_28803,N_27228,N_27570);
and U28804 (N_28804,N_27672,N_27048);
nand U28805 (N_28805,N_27394,N_27636);
nand U28806 (N_28806,N_27541,N_27787);
or U28807 (N_28807,N_27375,N_27383);
nand U28808 (N_28808,N_27219,N_27720);
nor U28809 (N_28809,N_27232,N_27786);
nor U28810 (N_28810,N_27148,N_27133);
or U28811 (N_28811,N_27730,N_27015);
nor U28812 (N_28812,N_27097,N_27519);
nand U28813 (N_28813,N_27802,N_27187);
and U28814 (N_28814,N_27345,N_27308);
nand U28815 (N_28815,N_27649,N_27605);
nand U28816 (N_28816,N_27402,N_27477);
nand U28817 (N_28817,N_27403,N_27571);
xnor U28818 (N_28818,N_27884,N_27607);
and U28819 (N_28819,N_27339,N_27984);
xor U28820 (N_28820,N_27695,N_27777);
nor U28821 (N_28821,N_27185,N_27988);
and U28822 (N_28822,N_27329,N_27322);
nand U28823 (N_28823,N_27332,N_27697);
nand U28824 (N_28824,N_27255,N_27960);
and U28825 (N_28825,N_27097,N_27031);
nor U28826 (N_28826,N_27775,N_27233);
xor U28827 (N_28827,N_27744,N_27802);
nand U28828 (N_28828,N_27329,N_27518);
and U28829 (N_28829,N_27543,N_27182);
and U28830 (N_28830,N_27327,N_27655);
or U28831 (N_28831,N_27884,N_27855);
nor U28832 (N_28832,N_27685,N_27285);
or U28833 (N_28833,N_27478,N_27884);
xnor U28834 (N_28834,N_27173,N_27628);
and U28835 (N_28835,N_27912,N_27636);
nor U28836 (N_28836,N_27305,N_27833);
xor U28837 (N_28837,N_27037,N_27640);
xor U28838 (N_28838,N_27457,N_27869);
and U28839 (N_28839,N_27879,N_27308);
nor U28840 (N_28840,N_27877,N_27420);
nand U28841 (N_28841,N_27047,N_27191);
xor U28842 (N_28842,N_27891,N_27091);
or U28843 (N_28843,N_27629,N_27097);
nor U28844 (N_28844,N_27280,N_27675);
xnor U28845 (N_28845,N_27014,N_27767);
and U28846 (N_28846,N_27593,N_27487);
nor U28847 (N_28847,N_27067,N_27848);
and U28848 (N_28848,N_27726,N_27959);
xor U28849 (N_28849,N_27104,N_27224);
nand U28850 (N_28850,N_27316,N_27998);
nand U28851 (N_28851,N_27260,N_27307);
nor U28852 (N_28852,N_27817,N_27463);
nand U28853 (N_28853,N_27197,N_27685);
nand U28854 (N_28854,N_27305,N_27975);
and U28855 (N_28855,N_27694,N_27194);
nor U28856 (N_28856,N_27874,N_27498);
nor U28857 (N_28857,N_27523,N_27175);
or U28858 (N_28858,N_27369,N_27433);
nor U28859 (N_28859,N_27796,N_27957);
or U28860 (N_28860,N_27128,N_27612);
or U28861 (N_28861,N_27663,N_27504);
nand U28862 (N_28862,N_27106,N_27088);
and U28863 (N_28863,N_27719,N_27028);
xor U28864 (N_28864,N_27349,N_27782);
or U28865 (N_28865,N_27864,N_27055);
or U28866 (N_28866,N_27415,N_27265);
nor U28867 (N_28867,N_27123,N_27013);
nand U28868 (N_28868,N_27022,N_27521);
nand U28869 (N_28869,N_27836,N_27564);
or U28870 (N_28870,N_27695,N_27859);
and U28871 (N_28871,N_27876,N_27863);
xnor U28872 (N_28872,N_27511,N_27955);
nor U28873 (N_28873,N_27204,N_27290);
and U28874 (N_28874,N_27732,N_27897);
xor U28875 (N_28875,N_27412,N_27227);
or U28876 (N_28876,N_27888,N_27922);
xnor U28877 (N_28877,N_27105,N_27767);
nor U28878 (N_28878,N_27951,N_27372);
nor U28879 (N_28879,N_27577,N_27900);
nor U28880 (N_28880,N_27066,N_27013);
xnor U28881 (N_28881,N_27528,N_27280);
and U28882 (N_28882,N_27127,N_27713);
and U28883 (N_28883,N_27076,N_27263);
nand U28884 (N_28884,N_27617,N_27037);
nor U28885 (N_28885,N_27495,N_27963);
and U28886 (N_28886,N_27436,N_27510);
and U28887 (N_28887,N_27185,N_27298);
nand U28888 (N_28888,N_27811,N_27927);
or U28889 (N_28889,N_27262,N_27751);
or U28890 (N_28890,N_27067,N_27949);
or U28891 (N_28891,N_27086,N_27224);
xor U28892 (N_28892,N_27429,N_27835);
nor U28893 (N_28893,N_27854,N_27763);
xor U28894 (N_28894,N_27845,N_27772);
nand U28895 (N_28895,N_27166,N_27083);
nor U28896 (N_28896,N_27171,N_27876);
xor U28897 (N_28897,N_27334,N_27244);
nand U28898 (N_28898,N_27208,N_27581);
nand U28899 (N_28899,N_27661,N_27139);
xnor U28900 (N_28900,N_27866,N_27487);
xor U28901 (N_28901,N_27072,N_27142);
nor U28902 (N_28902,N_27888,N_27810);
or U28903 (N_28903,N_27083,N_27399);
or U28904 (N_28904,N_27282,N_27237);
xnor U28905 (N_28905,N_27500,N_27259);
nand U28906 (N_28906,N_27405,N_27516);
nand U28907 (N_28907,N_27634,N_27202);
and U28908 (N_28908,N_27668,N_27319);
or U28909 (N_28909,N_27470,N_27473);
nor U28910 (N_28910,N_27854,N_27469);
and U28911 (N_28911,N_27485,N_27534);
xnor U28912 (N_28912,N_27236,N_27763);
nand U28913 (N_28913,N_27598,N_27060);
and U28914 (N_28914,N_27123,N_27827);
nand U28915 (N_28915,N_27383,N_27039);
or U28916 (N_28916,N_27212,N_27395);
nand U28917 (N_28917,N_27245,N_27927);
nor U28918 (N_28918,N_27701,N_27144);
nor U28919 (N_28919,N_27734,N_27104);
xor U28920 (N_28920,N_27681,N_27738);
and U28921 (N_28921,N_27609,N_27942);
xnor U28922 (N_28922,N_27273,N_27920);
and U28923 (N_28923,N_27509,N_27186);
and U28924 (N_28924,N_27969,N_27405);
nor U28925 (N_28925,N_27232,N_27322);
xnor U28926 (N_28926,N_27873,N_27745);
nand U28927 (N_28927,N_27445,N_27058);
or U28928 (N_28928,N_27420,N_27070);
or U28929 (N_28929,N_27949,N_27352);
and U28930 (N_28930,N_27092,N_27423);
and U28931 (N_28931,N_27332,N_27233);
or U28932 (N_28932,N_27837,N_27537);
nand U28933 (N_28933,N_27670,N_27913);
or U28934 (N_28934,N_27174,N_27253);
xnor U28935 (N_28935,N_27106,N_27798);
nor U28936 (N_28936,N_27838,N_27911);
xor U28937 (N_28937,N_27069,N_27919);
and U28938 (N_28938,N_27282,N_27025);
xnor U28939 (N_28939,N_27957,N_27906);
nand U28940 (N_28940,N_27205,N_27268);
nor U28941 (N_28941,N_27845,N_27197);
nor U28942 (N_28942,N_27345,N_27249);
nand U28943 (N_28943,N_27321,N_27217);
or U28944 (N_28944,N_27905,N_27984);
or U28945 (N_28945,N_27048,N_27850);
nand U28946 (N_28946,N_27847,N_27094);
or U28947 (N_28947,N_27235,N_27988);
and U28948 (N_28948,N_27905,N_27987);
or U28949 (N_28949,N_27619,N_27106);
or U28950 (N_28950,N_27032,N_27064);
nor U28951 (N_28951,N_27215,N_27102);
and U28952 (N_28952,N_27704,N_27171);
and U28953 (N_28953,N_27551,N_27390);
or U28954 (N_28954,N_27260,N_27468);
and U28955 (N_28955,N_27246,N_27338);
nor U28956 (N_28956,N_27964,N_27390);
nor U28957 (N_28957,N_27964,N_27073);
or U28958 (N_28958,N_27755,N_27482);
xnor U28959 (N_28959,N_27416,N_27950);
nand U28960 (N_28960,N_27002,N_27413);
nor U28961 (N_28961,N_27397,N_27825);
xor U28962 (N_28962,N_27337,N_27484);
nor U28963 (N_28963,N_27029,N_27330);
or U28964 (N_28964,N_27672,N_27147);
and U28965 (N_28965,N_27376,N_27413);
nand U28966 (N_28966,N_27183,N_27672);
nor U28967 (N_28967,N_27846,N_27623);
nor U28968 (N_28968,N_27803,N_27578);
nor U28969 (N_28969,N_27440,N_27761);
and U28970 (N_28970,N_27487,N_27602);
nand U28971 (N_28971,N_27460,N_27757);
and U28972 (N_28972,N_27357,N_27344);
nand U28973 (N_28973,N_27529,N_27253);
nand U28974 (N_28974,N_27352,N_27820);
nor U28975 (N_28975,N_27575,N_27410);
xor U28976 (N_28976,N_27965,N_27696);
or U28977 (N_28977,N_27322,N_27796);
and U28978 (N_28978,N_27215,N_27792);
xor U28979 (N_28979,N_27592,N_27675);
xnor U28980 (N_28980,N_27585,N_27735);
nor U28981 (N_28981,N_27701,N_27807);
xnor U28982 (N_28982,N_27486,N_27878);
nor U28983 (N_28983,N_27040,N_27873);
or U28984 (N_28984,N_27192,N_27517);
xor U28985 (N_28985,N_27908,N_27566);
nand U28986 (N_28986,N_27660,N_27680);
nor U28987 (N_28987,N_27262,N_27114);
nand U28988 (N_28988,N_27396,N_27530);
xor U28989 (N_28989,N_27928,N_27620);
and U28990 (N_28990,N_27450,N_27530);
xor U28991 (N_28991,N_27885,N_27603);
nor U28992 (N_28992,N_27042,N_27828);
or U28993 (N_28993,N_27672,N_27515);
nor U28994 (N_28994,N_27937,N_27667);
nor U28995 (N_28995,N_27217,N_27804);
xor U28996 (N_28996,N_27451,N_27416);
nor U28997 (N_28997,N_27356,N_27713);
or U28998 (N_28998,N_27063,N_27427);
or U28999 (N_28999,N_27494,N_27480);
and U29000 (N_29000,N_28940,N_28505);
and U29001 (N_29001,N_28526,N_28694);
xor U29002 (N_29002,N_28370,N_28826);
or U29003 (N_29003,N_28999,N_28088);
nor U29004 (N_29004,N_28126,N_28974);
and U29005 (N_29005,N_28161,N_28047);
nand U29006 (N_29006,N_28313,N_28683);
xnor U29007 (N_29007,N_28704,N_28925);
nor U29008 (N_29008,N_28955,N_28302);
nand U29009 (N_29009,N_28712,N_28506);
or U29010 (N_29010,N_28863,N_28921);
nand U29011 (N_29011,N_28757,N_28667);
nand U29012 (N_29012,N_28249,N_28623);
nor U29013 (N_29013,N_28630,N_28199);
nor U29014 (N_29014,N_28960,N_28225);
xor U29015 (N_29015,N_28379,N_28369);
nor U29016 (N_29016,N_28632,N_28942);
nand U29017 (N_29017,N_28344,N_28166);
and U29018 (N_29018,N_28730,N_28947);
and U29019 (N_29019,N_28777,N_28504);
and U29020 (N_29020,N_28403,N_28056);
and U29021 (N_29021,N_28409,N_28297);
or U29022 (N_29022,N_28152,N_28036);
xnor U29023 (N_29023,N_28258,N_28355);
xnor U29024 (N_29024,N_28223,N_28523);
and U29025 (N_29025,N_28202,N_28842);
or U29026 (N_29026,N_28368,N_28008);
nor U29027 (N_29027,N_28564,N_28348);
nor U29028 (N_29028,N_28354,N_28469);
nor U29029 (N_29029,N_28645,N_28823);
nand U29030 (N_29030,N_28634,N_28480);
and U29031 (N_29031,N_28111,N_28563);
and U29032 (N_29032,N_28383,N_28764);
or U29033 (N_29033,N_28272,N_28359);
nand U29034 (N_29034,N_28477,N_28858);
nor U29035 (N_29035,N_28839,N_28816);
xnor U29036 (N_29036,N_28035,N_28884);
nor U29037 (N_29037,N_28532,N_28930);
nand U29038 (N_29038,N_28615,N_28312);
xor U29039 (N_29039,N_28452,N_28619);
nand U29040 (N_29040,N_28872,N_28525);
xor U29041 (N_29041,N_28647,N_28459);
nand U29042 (N_29042,N_28576,N_28907);
xor U29043 (N_29043,N_28986,N_28649);
or U29044 (N_29044,N_28915,N_28716);
xnor U29045 (N_29045,N_28103,N_28723);
nor U29046 (N_29046,N_28113,N_28291);
xnor U29047 (N_29047,N_28541,N_28473);
and U29048 (N_29048,N_28441,N_28375);
nor U29049 (N_29049,N_28772,N_28701);
xor U29050 (N_29050,N_28766,N_28481);
xor U29051 (N_29051,N_28714,N_28463);
or U29052 (N_29052,N_28635,N_28236);
or U29053 (N_29053,N_28218,N_28700);
nand U29054 (N_29054,N_28901,N_28890);
and U29055 (N_29055,N_28808,N_28625);
or U29056 (N_29056,N_28226,N_28903);
or U29057 (N_29057,N_28274,N_28100);
nor U29058 (N_29058,N_28558,N_28407);
and U29059 (N_29059,N_28350,N_28989);
nor U29060 (N_29060,N_28434,N_28327);
and U29061 (N_29061,N_28596,N_28393);
or U29062 (N_29062,N_28167,N_28460);
nor U29063 (N_29063,N_28096,N_28186);
nor U29064 (N_29064,N_28612,N_28081);
nand U29065 (N_29065,N_28107,N_28484);
or U29066 (N_29066,N_28318,N_28255);
xor U29067 (N_29067,N_28843,N_28963);
nor U29068 (N_29068,N_28191,N_28394);
and U29069 (N_29069,N_28289,N_28796);
nor U29070 (N_29070,N_28495,N_28269);
nor U29071 (N_29071,N_28514,N_28799);
nor U29072 (N_29072,N_28916,N_28372);
and U29073 (N_29073,N_28728,N_28530);
and U29074 (N_29074,N_28817,N_28592);
xor U29075 (N_29075,N_28018,N_28055);
xnor U29076 (N_29076,N_28385,N_28206);
and U29077 (N_29077,N_28471,N_28430);
nand U29078 (N_29078,N_28785,N_28235);
xnor U29079 (N_29079,N_28896,N_28679);
or U29080 (N_29080,N_28024,N_28688);
or U29081 (N_29081,N_28973,N_28172);
or U29082 (N_29082,N_28013,N_28923);
nor U29083 (N_29083,N_28690,N_28412);
or U29084 (N_29084,N_28382,N_28182);
nand U29085 (N_29085,N_28600,N_28445);
and U29086 (N_29086,N_28352,N_28956);
nor U29087 (N_29087,N_28898,N_28954);
xor U29088 (N_29088,N_28391,N_28475);
or U29089 (N_29089,N_28908,N_28565);
nand U29090 (N_29090,N_28680,N_28544);
and U29091 (N_29091,N_28090,N_28945);
or U29092 (N_29092,N_28246,N_28222);
xor U29093 (N_29093,N_28941,N_28158);
and U29094 (N_29094,N_28440,N_28417);
and U29095 (N_29095,N_28579,N_28410);
xor U29096 (N_29096,N_28160,N_28936);
xor U29097 (N_29097,N_28060,N_28735);
nand U29098 (N_29098,N_28467,N_28549);
and U29099 (N_29099,N_28527,N_28092);
xor U29100 (N_29100,N_28201,N_28606);
and U29101 (N_29101,N_28809,N_28432);
nor U29102 (N_29102,N_28566,N_28749);
nor U29103 (N_29103,N_28298,N_28637);
xor U29104 (N_29104,N_28420,N_28847);
xor U29105 (N_29105,N_28075,N_28363);
nor U29106 (N_29106,N_28301,N_28639);
xnor U29107 (N_29107,N_28627,N_28012);
nor U29108 (N_29108,N_28949,N_28244);
and U29109 (N_29109,N_28337,N_28732);
nand U29110 (N_29110,N_28991,N_28065);
and U29111 (N_29111,N_28651,N_28573);
and U29112 (N_29112,N_28374,N_28709);
xnor U29113 (N_29113,N_28795,N_28154);
nand U29114 (N_29114,N_28870,N_28266);
xor U29115 (N_29115,N_28326,N_28052);
nor U29116 (N_29116,N_28132,N_28476);
or U29117 (N_29117,N_28399,N_28602);
or U29118 (N_29118,N_28586,N_28276);
or U29119 (N_29119,N_28436,N_28448);
nand U29120 (N_29120,N_28937,N_28791);
nand U29121 (N_29121,N_28979,N_28768);
xor U29122 (N_29122,N_28125,N_28569);
nor U29123 (N_29123,N_28567,N_28138);
and U29124 (N_29124,N_28806,N_28878);
and U29125 (N_29125,N_28057,N_28622);
nand U29126 (N_29126,N_28224,N_28177);
and U29127 (N_29127,N_28338,N_28015);
or U29128 (N_29128,N_28141,N_28618);
nor U29129 (N_29129,N_28290,N_28102);
nand U29130 (N_29130,N_28275,N_28365);
nand U29131 (N_29131,N_28192,N_28262);
and U29132 (N_29132,N_28773,N_28073);
or U29133 (N_29133,N_28142,N_28265);
xnor U29134 (N_29134,N_28256,N_28413);
nand U29135 (N_29135,N_28204,N_28769);
nor U29136 (N_29136,N_28767,N_28264);
and U29137 (N_29137,N_28756,N_28611);
xnor U29138 (N_29138,N_28707,N_28931);
nand U29139 (N_29139,N_28486,N_28912);
nor U29140 (N_29140,N_28234,N_28282);
xor U29141 (N_29141,N_28252,N_28509);
and U29142 (N_29142,N_28507,N_28361);
nand U29143 (N_29143,N_28129,N_28324);
xnor U29144 (N_29144,N_28388,N_28992);
nand U29145 (N_29145,N_28972,N_28343);
nor U29146 (N_29146,N_28342,N_28014);
nand U29147 (N_29147,N_28299,N_28851);
or U29148 (N_29148,N_28654,N_28577);
or U29149 (N_29149,N_28038,N_28997);
nand U29150 (N_29150,N_28961,N_28743);
and U29151 (N_29151,N_28457,N_28919);
nand U29152 (N_29152,N_28968,N_28351);
or U29153 (N_29153,N_28813,N_28758);
xnor U29154 (N_29154,N_28626,N_28697);
or U29155 (N_29155,N_28239,N_28729);
nor U29156 (N_29156,N_28001,N_28984);
nand U29157 (N_29157,N_28444,N_28561);
nor U29158 (N_29158,N_28660,N_28692);
and U29159 (N_29159,N_28300,N_28832);
xor U29160 (N_29160,N_28411,N_28019);
nor U29161 (N_29161,N_28605,N_28328);
xnor U29162 (N_29162,N_28774,N_28093);
nor U29163 (N_29163,N_28331,N_28016);
nand U29164 (N_29164,N_28496,N_28838);
or U29165 (N_29165,N_28589,N_28491);
nand U29166 (N_29166,N_28939,N_28621);
or U29167 (N_29167,N_28488,N_28115);
nand U29168 (N_29168,N_28454,N_28951);
xnor U29169 (N_29169,N_28010,N_28303);
or U29170 (N_29170,N_28221,N_28455);
xnor U29171 (N_29171,N_28396,N_28283);
or U29172 (N_29172,N_28539,N_28197);
xor U29173 (N_29173,N_28493,N_28489);
nand U29174 (N_29174,N_28286,N_28895);
xnor U29175 (N_29175,N_28557,N_28349);
or U29176 (N_29176,N_28451,N_28325);
nand U29177 (N_29177,N_28068,N_28547);
nand U29178 (N_29178,N_28340,N_28684);
nor U29179 (N_29179,N_28734,N_28831);
and U29180 (N_29180,N_28122,N_28686);
nor U29181 (N_29181,N_28519,N_28428);
nand U29182 (N_29182,N_28028,N_28139);
nor U29183 (N_29183,N_28641,N_28642);
and U29184 (N_29184,N_28702,N_28691);
nor U29185 (N_29185,N_28078,N_28501);
xor U29186 (N_29186,N_28336,N_28150);
xnor U29187 (N_29187,N_28074,N_28879);
and U29188 (N_29188,N_28780,N_28232);
xor U29189 (N_29189,N_28380,N_28636);
xor U29190 (N_29190,N_28442,N_28353);
or U29191 (N_29191,N_28751,N_28810);
nand U29192 (N_29192,N_28738,N_28083);
xor U29193 (N_29193,N_28554,N_28944);
nand U29194 (N_29194,N_28595,N_28775);
nor U29195 (N_29195,N_28560,N_28655);
and U29196 (N_29196,N_28985,N_28401);
and U29197 (N_29197,N_28095,N_28181);
nor U29198 (N_29198,N_28117,N_28064);
nor U29199 (N_29199,N_28120,N_28461);
nand U29200 (N_29200,N_28913,N_28717);
nand U29201 (N_29201,N_28718,N_28082);
nand U29202 (N_29202,N_28423,N_28934);
xnor U29203 (N_29203,N_28840,N_28722);
xor U29204 (N_29204,N_28517,N_28787);
nand U29205 (N_29205,N_28304,N_28362);
xor U29206 (N_29206,N_28248,N_28584);
nor U29207 (N_29207,N_28967,N_28614);
and U29208 (N_29208,N_28849,N_28146);
nand U29209 (N_29209,N_28646,N_28855);
nor U29210 (N_29210,N_28892,N_28296);
xor U29211 (N_29211,N_28850,N_28321);
and U29212 (N_29212,N_28762,N_28971);
nand U29213 (N_29213,N_28883,N_28127);
nand U29214 (N_29214,N_28828,N_28891);
or U29215 (N_29215,N_28969,N_28835);
and U29216 (N_29216,N_28946,N_28000);
and U29217 (N_29217,N_28869,N_28270);
nor U29218 (N_29218,N_28281,N_28169);
and U29219 (N_29219,N_28593,N_28535);
and U29220 (N_29220,N_28315,N_28292);
xnor U29221 (N_29221,N_28433,N_28603);
and U29222 (N_29222,N_28953,N_28957);
nand U29223 (N_29223,N_28040,N_28546);
nor U29224 (N_29224,N_28562,N_28920);
nor U29225 (N_29225,N_28168,N_28695);
nor U29226 (N_29226,N_28906,N_28678);
or U29227 (N_29227,N_28447,N_28833);
nand U29228 (N_29228,N_28776,N_28044);
nor U29229 (N_29229,N_28478,N_28990);
nor U29230 (N_29230,N_28176,N_28824);
nand U29231 (N_29231,N_28508,N_28384);
xnor U29232 (N_29232,N_28594,N_28458);
nand U29233 (N_29233,N_28091,N_28994);
and U29234 (N_29234,N_28449,N_28273);
nor U29235 (N_29235,N_28240,N_28926);
nand U29236 (N_29236,N_28498,N_28609);
and U29237 (N_29237,N_28051,N_28877);
xnor U29238 (N_29238,N_28268,N_28004);
or U29239 (N_29239,N_28727,N_28456);
xor U29240 (N_29240,N_28748,N_28742);
xnor U29241 (N_29241,N_28136,N_28736);
or U29242 (N_29242,N_28002,N_28556);
nand U29243 (N_29243,N_28144,N_28811);
xor U29244 (N_29244,N_28534,N_28807);
and U29245 (N_29245,N_28259,N_28205);
and U29246 (N_29246,N_28978,N_28765);
xnor U29247 (N_29247,N_28149,N_28247);
and U29248 (N_29248,N_28208,N_28426);
nor U29249 (N_29249,N_28101,N_28644);
xor U29250 (N_29250,N_28039,N_28219);
xnor U29251 (N_29251,N_28069,N_28200);
nor U29252 (N_29252,N_28104,N_28882);
and U29253 (N_29253,N_28502,N_28804);
nor U29254 (N_29254,N_28470,N_28613);
and U29255 (N_29255,N_28474,N_28604);
nand U29256 (N_29256,N_28784,N_28744);
or U29257 (N_29257,N_28996,N_28513);
nand U29258 (N_29258,N_28753,N_28750);
nand U29259 (N_29259,N_28251,N_28446);
and U29260 (N_29260,N_28341,N_28285);
nor U29261 (N_29261,N_28468,N_28173);
nand U29262 (N_29262,N_28003,N_28725);
nor U29263 (N_29263,N_28786,N_28076);
or U29264 (N_29264,N_28042,N_28652);
nor U29265 (N_29265,N_28827,N_28376);
and U29266 (N_29266,N_28287,N_28800);
and U29267 (N_29267,N_28425,N_28123);
nor U29268 (N_29268,N_28034,N_28329);
nor U29269 (N_29269,N_28515,N_28114);
or U29270 (N_29270,N_28894,N_28995);
or U29271 (N_29271,N_28211,N_28320);
nor U29272 (N_29272,N_28049,N_28212);
nor U29273 (N_29273,N_28520,N_28797);
nor U29274 (N_29274,N_28875,N_28179);
nand U29275 (N_29275,N_28472,N_28705);
nor U29276 (N_29276,N_28306,N_28213);
or U29277 (N_29277,N_28229,N_28422);
and U29278 (N_29278,N_28771,N_28581);
nor U29279 (N_29279,N_28629,N_28398);
xnor U29280 (N_29280,N_28397,N_28747);
nor U29281 (N_29281,N_28080,N_28007);
or U29282 (N_29282,N_28392,N_28105);
or U29283 (N_29283,N_28097,N_28022);
and U29284 (N_29284,N_28553,N_28572);
or U29285 (N_29285,N_28006,N_28815);
xor U29286 (N_29286,N_28656,N_28531);
xnor U29287 (N_29287,N_28108,N_28148);
nand U29288 (N_29288,N_28360,N_28109);
nand U29289 (N_29289,N_28601,N_28983);
or U29290 (N_29290,N_28050,N_28187);
xnor U29291 (N_29291,N_28373,N_28868);
nor U29292 (N_29292,N_28453,N_28021);
nor U29293 (N_29293,N_28263,N_28437);
xnor U29294 (N_29294,N_28741,N_28171);
xor U29295 (N_29295,N_28190,N_28294);
nor U29296 (N_29296,N_28518,N_28086);
xnor U29297 (N_29297,N_28818,N_28904);
or U29298 (N_29298,N_28402,N_28227);
nand U29299 (N_29299,N_28802,N_28147);
and U29300 (N_29300,N_28308,N_28574);
or U29301 (N_29301,N_28711,N_28072);
nand U29302 (N_29302,N_28077,N_28427);
nor U29303 (N_29303,N_28825,N_28881);
and U29304 (N_29304,N_28617,N_28638);
or U29305 (N_29305,N_28676,N_28793);
and U29306 (N_29306,N_28917,N_28494);
and U29307 (N_29307,N_28922,N_28841);
nand U29308 (N_29308,N_28031,N_28465);
or U29309 (N_29309,N_28788,N_28307);
or U29310 (N_29310,N_28801,N_28233);
xnor U29311 (N_29311,N_28358,N_28070);
or U29312 (N_29312,N_28591,N_28929);
xnor U29313 (N_29313,N_28664,N_28099);
xor U29314 (N_29314,N_28862,N_28054);
xnor U29315 (N_29315,N_28277,N_28438);
nor U29316 (N_29316,N_28366,N_28876);
and U29317 (N_29317,N_28032,N_28880);
nand U29318 (N_29318,N_28046,N_28928);
xor U29319 (N_29319,N_28020,N_28713);
and U29320 (N_29320,N_28681,N_28865);
and U29321 (N_29321,N_28311,N_28322);
nor U29322 (N_29322,N_28689,N_28180);
nor U29323 (N_29323,N_28543,N_28071);
xnor U29324 (N_29324,N_28079,N_28536);
or U29325 (N_29325,N_28976,N_28698);
and U29326 (N_29326,N_28899,N_28053);
nor U29327 (N_29327,N_28378,N_28836);
or U29328 (N_29328,N_28902,N_28216);
and U29329 (N_29329,N_28545,N_28231);
and U29330 (N_29330,N_28552,N_28669);
nor U29331 (N_29331,N_28404,N_28250);
xnor U29332 (N_29332,N_28703,N_28958);
nand U29333 (N_29333,N_28414,N_28682);
and U29334 (N_29334,N_28548,N_28867);
nand U29335 (N_29335,N_28568,N_28314);
xor U29336 (N_29336,N_28253,N_28643);
xor U29337 (N_29337,N_28524,N_28210);
xnor U29338 (N_29338,N_28608,N_28431);
and U29339 (N_29339,N_28790,N_28998);
and U29340 (N_29340,N_28537,N_28106);
or U29341 (N_29341,N_28837,N_28740);
nand U29342 (N_29342,N_28943,N_28779);
nor U29343 (N_29343,N_28668,N_28580);
and U29344 (N_29344,N_28640,N_28209);
or U29345 (N_29345,N_28852,N_28970);
xor U29346 (N_29346,N_28242,N_28677);
and U29347 (N_29347,N_28439,N_28610);
or U29348 (N_29348,N_28633,N_28653);
or U29349 (N_29349,N_28116,N_28885);
and U29350 (N_29350,N_28975,N_28214);
nand U29351 (N_29351,N_28783,N_28759);
nor U29352 (N_29352,N_28217,N_28155);
or U29353 (N_29353,N_28673,N_28571);
or U29354 (N_29354,N_28893,N_28752);
and U29355 (N_29355,N_28721,N_28381);
nor U29356 (N_29356,N_28657,N_28585);
nand U29357 (N_29357,N_28371,N_28932);
and U29358 (N_29358,N_28162,N_28156);
and U29359 (N_29359,N_28829,N_28323);
nand U29360 (N_29360,N_28395,N_28763);
xor U29361 (N_29361,N_28755,N_28966);
xnor U29362 (N_29362,N_28485,N_28821);
or U29363 (N_29363,N_28911,N_28119);
xor U29364 (N_29364,N_28165,N_28066);
xnor U29365 (N_29365,N_28559,N_28196);
or U29366 (N_29366,N_28500,N_28131);
nand U29367 (N_29367,N_28085,N_28859);
or U29368 (N_29368,N_28406,N_28529);
xor U29369 (N_29369,N_28819,N_28230);
nand U29370 (N_29370,N_28087,N_28030);
and U29371 (N_29371,N_28964,N_28220);
nor U29372 (N_29372,N_28174,N_28731);
xnor U29373 (N_29373,N_28708,N_28822);
or U29374 (N_29374,N_28624,N_28587);
xnor U29375 (N_29375,N_28598,N_28853);
xnor U29376 (N_29376,N_28662,N_28720);
and U29377 (N_29377,N_28950,N_28124);
nor U29378 (N_29378,N_28347,N_28663);
xnor U29379 (N_29379,N_28977,N_28261);
nor U29380 (N_29380,N_28650,N_28988);
nand U29381 (N_29381,N_28178,N_28133);
and U29382 (N_29382,N_28089,N_28511);
nand U29383 (N_29383,N_28377,N_28830);
and U29384 (N_29384,N_28450,N_28159);
nor U29385 (N_29385,N_28464,N_28429);
nor U29386 (N_29386,N_28193,N_28948);
and U29387 (N_29387,N_28803,N_28254);
xor U29388 (N_29388,N_28151,N_28888);
or U29389 (N_29389,N_28959,N_28687);
nand U29390 (N_29390,N_28607,N_28267);
nor U29391 (N_29391,N_28198,N_28424);
or U29392 (N_29392,N_28864,N_28027);
nand U29393 (N_29393,N_28243,N_28009);
xor U29394 (N_29394,N_28094,N_28188);
nand U29395 (N_29395,N_28555,N_28789);
nand U29396 (N_29396,N_28356,N_28330);
xor U29397 (N_29397,N_28918,N_28861);
or U29398 (N_29398,N_28130,N_28482);
or U29399 (N_29399,N_28550,N_28062);
nand U29400 (N_29400,N_28737,N_28490);
nand U29401 (N_29401,N_28023,N_28845);
nor U29402 (N_29402,N_28387,N_28048);
xnor U29403 (N_29403,N_28335,N_28134);
and U29404 (N_29404,N_28386,N_28043);
or U29405 (N_29405,N_28037,N_28980);
and U29406 (N_29406,N_28933,N_28710);
or U29407 (N_29407,N_28857,N_28814);
and U29408 (N_29408,N_28164,N_28820);
nor U29409 (N_29409,N_28914,N_28499);
nand U29410 (N_29410,N_28416,N_28583);
xnor U29411 (N_29411,N_28059,N_28616);
and U29412 (N_29412,N_28761,N_28510);
or U29413 (N_29413,N_28540,N_28782);
and U29414 (N_29414,N_28671,N_28860);
xnor U29415 (N_29415,N_28533,N_28245);
nand U29416 (N_29416,N_28389,N_28184);
and U29417 (N_29417,N_28084,N_28658);
and U29418 (N_29418,N_28058,N_28479);
and U29419 (N_29419,N_28271,N_28542);
and U29420 (N_29420,N_28726,N_28487);
xnor U29421 (N_29421,N_28575,N_28163);
and U29422 (N_29422,N_28887,N_28699);
xor U29423 (N_29423,N_28345,N_28145);
and U29424 (N_29424,N_28305,N_28993);
nor U29425 (N_29425,N_28844,N_28551);
xnor U29426 (N_29426,N_28854,N_28719);
xor U29427 (N_29427,N_28153,N_28798);
nor U29428 (N_29428,N_28157,N_28897);
or U29429 (N_29429,N_28848,N_28492);
nand U29430 (N_29430,N_28497,N_28310);
or U29431 (N_29431,N_28874,N_28257);
nand U29432 (N_29432,N_28696,N_28135);
nor U29433 (N_29433,N_28260,N_28026);
nand U29434 (N_29434,N_28812,N_28367);
xor U29435 (N_29435,N_28241,N_28733);
xor U29436 (N_29436,N_28538,N_28628);
nor U29437 (N_29437,N_28962,N_28620);
and U29438 (N_29438,N_28357,N_28659);
nand U29439 (N_29439,N_28293,N_28415);
xnor U29440 (N_29440,N_28185,N_28528);
xnor U29441 (N_29441,N_28207,N_28203);
nor U29442 (N_29442,N_28805,N_28462);
and U29443 (N_29443,N_28183,N_28866);
nor U29444 (N_29444,N_28512,N_28137);
xnor U29445 (N_29445,N_28280,N_28061);
and U29446 (N_29446,N_28284,N_28685);
nor U29447 (N_29447,N_28045,N_28118);
and U29448 (N_29448,N_28905,N_28674);
nor U29449 (N_29449,N_28935,N_28029);
xnor U29450 (N_29450,N_28189,N_28316);
and U29451 (N_29451,N_28794,N_28194);
xor U29452 (N_29452,N_28900,N_28856);
xnor U29453 (N_29453,N_28067,N_28873);
and U29454 (N_29454,N_28746,N_28754);
or U29455 (N_29455,N_28140,N_28981);
nand U29456 (N_29456,N_28228,N_28346);
or U29457 (N_29457,N_28648,N_28390);
nand U29458 (N_29458,N_28670,N_28435);
and U29459 (N_29459,N_28110,N_28570);
nor U29460 (N_29460,N_28339,N_28672);
nor U29461 (N_29461,N_28279,N_28781);
or U29462 (N_29462,N_28760,N_28938);
and U29463 (N_29463,N_28521,N_28483);
or U29464 (N_29464,N_28588,N_28332);
nand U29465 (N_29465,N_28503,N_28982);
or U29466 (N_29466,N_28319,N_28418);
nor U29467 (N_29467,N_28597,N_28364);
or U29468 (N_29468,N_28295,N_28924);
xnor U29469 (N_29469,N_28886,N_28309);
nand U29470 (N_29470,N_28724,N_28693);
xor U29471 (N_29471,N_28578,N_28400);
nor U29472 (N_29472,N_28739,N_28405);
and U29473 (N_29473,N_28128,N_28987);
or U29474 (N_29474,N_28143,N_28846);
nand U29475 (N_29475,N_28952,N_28215);
and U29476 (N_29476,N_28466,N_28631);
and U29477 (N_29477,N_28041,N_28871);
or U29478 (N_29478,N_28582,N_28011);
nor U29479 (N_29479,N_28927,N_28834);
nand U29480 (N_29480,N_28005,N_28675);
xnor U29481 (N_29481,N_28408,N_28317);
nor U29482 (N_29482,N_28661,N_28025);
nor U29483 (N_29483,N_28278,N_28237);
nand U29484 (N_29484,N_28170,N_28666);
xor U29485 (N_29485,N_28590,N_28121);
or U29486 (N_29486,N_28238,N_28965);
nand U29487 (N_29487,N_28288,N_28745);
and U29488 (N_29488,N_28063,N_28792);
nor U29489 (N_29489,N_28195,N_28778);
nand U29490 (N_29490,N_28443,N_28017);
or U29491 (N_29491,N_28770,N_28910);
nor U29492 (N_29492,N_28419,N_28333);
or U29493 (N_29493,N_28098,N_28175);
nand U29494 (N_29494,N_28599,N_28522);
and U29495 (N_29495,N_28909,N_28033);
and U29496 (N_29496,N_28516,N_28421);
xor U29497 (N_29497,N_28706,N_28334);
or U29498 (N_29498,N_28665,N_28715);
or U29499 (N_29499,N_28889,N_28112);
nand U29500 (N_29500,N_28426,N_28468);
nand U29501 (N_29501,N_28609,N_28944);
and U29502 (N_29502,N_28112,N_28273);
xor U29503 (N_29503,N_28250,N_28460);
and U29504 (N_29504,N_28530,N_28987);
or U29505 (N_29505,N_28674,N_28720);
or U29506 (N_29506,N_28640,N_28622);
or U29507 (N_29507,N_28710,N_28632);
nand U29508 (N_29508,N_28498,N_28448);
nor U29509 (N_29509,N_28540,N_28036);
nor U29510 (N_29510,N_28867,N_28551);
and U29511 (N_29511,N_28736,N_28399);
or U29512 (N_29512,N_28281,N_28138);
and U29513 (N_29513,N_28102,N_28616);
nor U29514 (N_29514,N_28048,N_28247);
xor U29515 (N_29515,N_28294,N_28944);
xor U29516 (N_29516,N_28951,N_28576);
nand U29517 (N_29517,N_28949,N_28390);
or U29518 (N_29518,N_28652,N_28663);
nor U29519 (N_29519,N_28991,N_28388);
nor U29520 (N_29520,N_28330,N_28200);
xnor U29521 (N_29521,N_28310,N_28101);
nand U29522 (N_29522,N_28166,N_28671);
and U29523 (N_29523,N_28732,N_28751);
xnor U29524 (N_29524,N_28366,N_28920);
xnor U29525 (N_29525,N_28262,N_28103);
and U29526 (N_29526,N_28334,N_28150);
nand U29527 (N_29527,N_28512,N_28907);
or U29528 (N_29528,N_28747,N_28350);
nand U29529 (N_29529,N_28308,N_28291);
nand U29530 (N_29530,N_28278,N_28045);
xnor U29531 (N_29531,N_28600,N_28037);
xor U29532 (N_29532,N_28628,N_28459);
nor U29533 (N_29533,N_28500,N_28582);
xor U29534 (N_29534,N_28507,N_28157);
and U29535 (N_29535,N_28866,N_28727);
xor U29536 (N_29536,N_28594,N_28981);
nor U29537 (N_29537,N_28446,N_28827);
and U29538 (N_29538,N_28927,N_28844);
nand U29539 (N_29539,N_28007,N_28354);
or U29540 (N_29540,N_28915,N_28689);
nor U29541 (N_29541,N_28462,N_28081);
nor U29542 (N_29542,N_28320,N_28046);
and U29543 (N_29543,N_28765,N_28352);
xnor U29544 (N_29544,N_28058,N_28392);
nor U29545 (N_29545,N_28625,N_28996);
nor U29546 (N_29546,N_28304,N_28673);
nand U29547 (N_29547,N_28219,N_28339);
and U29548 (N_29548,N_28792,N_28746);
xor U29549 (N_29549,N_28756,N_28870);
nand U29550 (N_29550,N_28633,N_28931);
nand U29551 (N_29551,N_28936,N_28791);
xnor U29552 (N_29552,N_28395,N_28004);
nor U29553 (N_29553,N_28988,N_28085);
or U29554 (N_29554,N_28108,N_28316);
xnor U29555 (N_29555,N_28072,N_28455);
or U29556 (N_29556,N_28917,N_28362);
nor U29557 (N_29557,N_28832,N_28793);
nand U29558 (N_29558,N_28865,N_28331);
nand U29559 (N_29559,N_28887,N_28765);
nand U29560 (N_29560,N_28631,N_28946);
or U29561 (N_29561,N_28790,N_28354);
nor U29562 (N_29562,N_28104,N_28173);
or U29563 (N_29563,N_28496,N_28731);
nand U29564 (N_29564,N_28890,N_28566);
nand U29565 (N_29565,N_28293,N_28956);
nor U29566 (N_29566,N_28520,N_28527);
xnor U29567 (N_29567,N_28468,N_28819);
xor U29568 (N_29568,N_28103,N_28356);
and U29569 (N_29569,N_28792,N_28518);
nor U29570 (N_29570,N_28849,N_28342);
and U29571 (N_29571,N_28912,N_28896);
or U29572 (N_29572,N_28299,N_28389);
nor U29573 (N_29573,N_28319,N_28604);
nor U29574 (N_29574,N_28353,N_28875);
nand U29575 (N_29575,N_28666,N_28481);
nand U29576 (N_29576,N_28470,N_28389);
xnor U29577 (N_29577,N_28104,N_28076);
nand U29578 (N_29578,N_28782,N_28229);
and U29579 (N_29579,N_28616,N_28642);
nand U29580 (N_29580,N_28427,N_28767);
or U29581 (N_29581,N_28730,N_28179);
nor U29582 (N_29582,N_28301,N_28084);
and U29583 (N_29583,N_28938,N_28710);
xor U29584 (N_29584,N_28347,N_28395);
nor U29585 (N_29585,N_28073,N_28595);
nor U29586 (N_29586,N_28718,N_28465);
nor U29587 (N_29587,N_28185,N_28797);
nor U29588 (N_29588,N_28434,N_28013);
or U29589 (N_29589,N_28626,N_28157);
xor U29590 (N_29590,N_28004,N_28851);
xnor U29591 (N_29591,N_28573,N_28395);
or U29592 (N_29592,N_28994,N_28975);
and U29593 (N_29593,N_28534,N_28523);
and U29594 (N_29594,N_28488,N_28113);
and U29595 (N_29595,N_28628,N_28423);
xor U29596 (N_29596,N_28481,N_28101);
or U29597 (N_29597,N_28538,N_28477);
xor U29598 (N_29598,N_28533,N_28037);
and U29599 (N_29599,N_28963,N_28261);
nand U29600 (N_29600,N_28053,N_28297);
or U29601 (N_29601,N_28126,N_28195);
or U29602 (N_29602,N_28190,N_28168);
xnor U29603 (N_29603,N_28228,N_28763);
or U29604 (N_29604,N_28515,N_28299);
or U29605 (N_29605,N_28346,N_28642);
or U29606 (N_29606,N_28006,N_28637);
xor U29607 (N_29607,N_28111,N_28480);
nand U29608 (N_29608,N_28086,N_28884);
nand U29609 (N_29609,N_28371,N_28266);
nand U29610 (N_29610,N_28010,N_28403);
nor U29611 (N_29611,N_28554,N_28774);
xor U29612 (N_29612,N_28009,N_28431);
or U29613 (N_29613,N_28354,N_28786);
or U29614 (N_29614,N_28836,N_28193);
and U29615 (N_29615,N_28250,N_28480);
xnor U29616 (N_29616,N_28885,N_28855);
or U29617 (N_29617,N_28732,N_28180);
or U29618 (N_29618,N_28932,N_28506);
nand U29619 (N_29619,N_28061,N_28664);
nor U29620 (N_29620,N_28398,N_28252);
nor U29621 (N_29621,N_28223,N_28643);
or U29622 (N_29622,N_28824,N_28424);
xor U29623 (N_29623,N_28083,N_28268);
and U29624 (N_29624,N_28594,N_28630);
and U29625 (N_29625,N_28636,N_28561);
nor U29626 (N_29626,N_28221,N_28528);
and U29627 (N_29627,N_28537,N_28453);
and U29628 (N_29628,N_28380,N_28694);
or U29629 (N_29629,N_28355,N_28243);
xor U29630 (N_29630,N_28406,N_28473);
nand U29631 (N_29631,N_28051,N_28997);
or U29632 (N_29632,N_28917,N_28395);
nor U29633 (N_29633,N_28769,N_28525);
and U29634 (N_29634,N_28877,N_28358);
xor U29635 (N_29635,N_28945,N_28270);
xor U29636 (N_29636,N_28025,N_28001);
xor U29637 (N_29637,N_28271,N_28588);
and U29638 (N_29638,N_28220,N_28265);
or U29639 (N_29639,N_28335,N_28749);
and U29640 (N_29640,N_28014,N_28099);
or U29641 (N_29641,N_28413,N_28959);
or U29642 (N_29642,N_28992,N_28077);
nor U29643 (N_29643,N_28914,N_28084);
nor U29644 (N_29644,N_28717,N_28412);
nor U29645 (N_29645,N_28284,N_28238);
or U29646 (N_29646,N_28006,N_28908);
xor U29647 (N_29647,N_28118,N_28765);
xnor U29648 (N_29648,N_28251,N_28827);
nor U29649 (N_29649,N_28828,N_28096);
and U29650 (N_29650,N_28051,N_28839);
nor U29651 (N_29651,N_28109,N_28681);
and U29652 (N_29652,N_28392,N_28462);
and U29653 (N_29653,N_28495,N_28231);
and U29654 (N_29654,N_28543,N_28251);
and U29655 (N_29655,N_28531,N_28802);
nor U29656 (N_29656,N_28089,N_28569);
or U29657 (N_29657,N_28860,N_28050);
or U29658 (N_29658,N_28242,N_28070);
or U29659 (N_29659,N_28092,N_28138);
nor U29660 (N_29660,N_28765,N_28078);
xnor U29661 (N_29661,N_28279,N_28480);
or U29662 (N_29662,N_28006,N_28964);
nand U29663 (N_29663,N_28542,N_28566);
nand U29664 (N_29664,N_28434,N_28521);
xor U29665 (N_29665,N_28550,N_28748);
nand U29666 (N_29666,N_28457,N_28704);
nand U29667 (N_29667,N_28206,N_28434);
xnor U29668 (N_29668,N_28194,N_28078);
nor U29669 (N_29669,N_28343,N_28445);
nor U29670 (N_29670,N_28541,N_28368);
and U29671 (N_29671,N_28263,N_28450);
nor U29672 (N_29672,N_28020,N_28475);
or U29673 (N_29673,N_28268,N_28344);
nor U29674 (N_29674,N_28200,N_28897);
xor U29675 (N_29675,N_28097,N_28556);
xnor U29676 (N_29676,N_28161,N_28006);
nand U29677 (N_29677,N_28465,N_28592);
and U29678 (N_29678,N_28203,N_28383);
and U29679 (N_29679,N_28893,N_28565);
or U29680 (N_29680,N_28343,N_28335);
or U29681 (N_29681,N_28825,N_28563);
nand U29682 (N_29682,N_28666,N_28706);
nand U29683 (N_29683,N_28496,N_28723);
xnor U29684 (N_29684,N_28117,N_28113);
or U29685 (N_29685,N_28139,N_28036);
or U29686 (N_29686,N_28070,N_28934);
nor U29687 (N_29687,N_28137,N_28583);
xnor U29688 (N_29688,N_28997,N_28914);
nor U29689 (N_29689,N_28260,N_28978);
nor U29690 (N_29690,N_28273,N_28262);
xor U29691 (N_29691,N_28043,N_28756);
xnor U29692 (N_29692,N_28595,N_28383);
nor U29693 (N_29693,N_28948,N_28711);
nand U29694 (N_29694,N_28475,N_28647);
xnor U29695 (N_29695,N_28457,N_28980);
and U29696 (N_29696,N_28746,N_28476);
and U29697 (N_29697,N_28381,N_28332);
or U29698 (N_29698,N_28574,N_28667);
xnor U29699 (N_29699,N_28155,N_28230);
or U29700 (N_29700,N_28542,N_28088);
and U29701 (N_29701,N_28056,N_28020);
nor U29702 (N_29702,N_28604,N_28459);
xnor U29703 (N_29703,N_28457,N_28229);
or U29704 (N_29704,N_28477,N_28676);
nand U29705 (N_29705,N_28715,N_28656);
and U29706 (N_29706,N_28560,N_28038);
and U29707 (N_29707,N_28249,N_28954);
or U29708 (N_29708,N_28878,N_28062);
nor U29709 (N_29709,N_28849,N_28930);
xnor U29710 (N_29710,N_28266,N_28464);
nand U29711 (N_29711,N_28387,N_28234);
or U29712 (N_29712,N_28398,N_28102);
xnor U29713 (N_29713,N_28307,N_28321);
nand U29714 (N_29714,N_28328,N_28486);
or U29715 (N_29715,N_28411,N_28448);
xor U29716 (N_29716,N_28977,N_28889);
xnor U29717 (N_29717,N_28261,N_28350);
or U29718 (N_29718,N_28590,N_28013);
nand U29719 (N_29719,N_28694,N_28995);
or U29720 (N_29720,N_28777,N_28232);
and U29721 (N_29721,N_28250,N_28953);
xnor U29722 (N_29722,N_28627,N_28880);
and U29723 (N_29723,N_28233,N_28671);
and U29724 (N_29724,N_28712,N_28286);
nor U29725 (N_29725,N_28223,N_28469);
nand U29726 (N_29726,N_28025,N_28607);
and U29727 (N_29727,N_28106,N_28727);
and U29728 (N_29728,N_28790,N_28722);
nand U29729 (N_29729,N_28262,N_28160);
or U29730 (N_29730,N_28126,N_28351);
nand U29731 (N_29731,N_28504,N_28346);
xnor U29732 (N_29732,N_28320,N_28516);
nor U29733 (N_29733,N_28144,N_28733);
or U29734 (N_29734,N_28880,N_28732);
or U29735 (N_29735,N_28241,N_28364);
nor U29736 (N_29736,N_28804,N_28651);
or U29737 (N_29737,N_28785,N_28207);
or U29738 (N_29738,N_28087,N_28170);
nor U29739 (N_29739,N_28974,N_28880);
nor U29740 (N_29740,N_28806,N_28009);
nand U29741 (N_29741,N_28343,N_28545);
nor U29742 (N_29742,N_28365,N_28197);
or U29743 (N_29743,N_28847,N_28759);
xnor U29744 (N_29744,N_28049,N_28228);
or U29745 (N_29745,N_28062,N_28435);
xor U29746 (N_29746,N_28561,N_28304);
and U29747 (N_29747,N_28769,N_28149);
and U29748 (N_29748,N_28787,N_28125);
nor U29749 (N_29749,N_28609,N_28333);
nor U29750 (N_29750,N_28223,N_28687);
or U29751 (N_29751,N_28230,N_28987);
or U29752 (N_29752,N_28240,N_28502);
and U29753 (N_29753,N_28754,N_28092);
nand U29754 (N_29754,N_28291,N_28384);
nor U29755 (N_29755,N_28112,N_28461);
or U29756 (N_29756,N_28049,N_28533);
xnor U29757 (N_29757,N_28367,N_28788);
xor U29758 (N_29758,N_28721,N_28434);
nor U29759 (N_29759,N_28574,N_28168);
nor U29760 (N_29760,N_28485,N_28484);
nand U29761 (N_29761,N_28031,N_28685);
xor U29762 (N_29762,N_28664,N_28562);
xor U29763 (N_29763,N_28690,N_28757);
nand U29764 (N_29764,N_28271,N_28861);
nand U29765 (N_29765,N_28789,N_28364);
and U29766 (N_29766,N_28081,N_28776);
or U29767 (N_29767,N_28889,N_28962);
nand U29768 (N_29768,N_28013,N_28883);
nand U29769 (N_29769,N_28440,N_28783);
or U29770 (N_29770,N_28541,N_28784);
nor U29771 (N_29771,N_28405,N_28176);
or U29772 (N_29772,N_28103,N_28843);
or U29773 (N_29773,N_28631,N_28104);
or U29774 (N_29774,N_28499,N_28162);
nor U29775 (N_29775,N_28726,N_28591);
nand U29776 (N_29776,N_28104,N_28369);
or U29777 (N_29777,N_28130,N_28859);
or U29778 (N_29778,N_28591,N_28377);
nand U29779 (N_29779,N_28758,N_28452);
and U29780 (N_29780,N_28264,N_28036);
nor U29781 (N_29781,N_28013,N_28862);
and U29782 (N_29782,N_28807,N_28224);
nor U29783 (N_29783,N_28337,N_28902);
and U29784 (N_29784,N_28297,N_28509);
or U29785 (N_29785,N_28509,N_28205);
nand U29786 (N_29786,N_28977,N_28767);
nor U29787 (N_29787,N_28347,N_28542);
nor U29788 (N_29788,N_28199,N_28543);
nor U29789 (N_29789,N_28379,N_28391);
nor U29790 (N_29790,N_28850,N_28045);
nand U29791 (N_29791,N_28075,N_28229);
nand U29792 (N_29792,N_28771,N_28579);
or U29793 (N_29793,N_28451,N_28167);
or U29794 (N_29794,N_28936,N_28028);
nand U29795 (N_29795,N_28298,N_28949);
nor U29796 (N_29796,N_28507,N_28175);
xor U29797 (N_29797,N_28931,N_28006);
and U29798 (N_29798,N_28299,N_28517);
nand U29799 (N_29799,N_28596,N_28190);
xor U29800 (N_29800,N_28521,N_28131);
or U29801 (N_29801,N_28624,N_28028);
or U29802 (N_29802,N_28558,N_28440);
nand U29803 (N_29803,N_28276,N_28714);
and U29804 (N_29804,N_28315,N_28959);
or U29805 (N_29805,N_28945,N_28521);
nor U29806 (N_29806,N_28714,N_28153);
or U29807 (N_29807,N_28752,N_28789);
nor U29808 (N_29808,N_28180,N_28301);
nor U29809 (N_29809,N_28582,N_28002);
xor U29810 (N_29810,N_28292,N_28168);
nand U29811 (N_29811,N_28036,N_28069);
and U29812 (N_29812,N_28443,N_28520);
xnor U29813 (N_29813,N_28691,N_28448);
and U29814 (N_29814,N_28311,N_28848);
and U29815 (N_29815,N_28656,N_28320);
nor U29816 (N_29816,N_28478,N_28654);
xnor U29817 (N_29817,N_28858,N_28439);
nor U29818 (N_29818,N_28370,N_28168);
and U29819 (N_29819,N_28360,N_28984);
and U29820 (N_29820,N_28119,N_28221);
nor U29821 (N_29821,N_28541,N_28030);
and U29822 (N_29822,N_28394,N_28367);
xor U29823 (N_29823,N_28923,N_28031);
or U29824 (N_29824,N_28730,N_28897);
xor U29825 (N_29825,N_28316,N_28990);
nand U29826 (N_29826,N_28818,N_28503);
or U29827 (N_29827,N_28892,N_28376);
nor U29828 (N_29828,N_28017,N_28276);
nor U29829 (N_29829,N_28802,N_28927);
nand U29830 (N_29830,N_28142,N_28835);
nor U29831 (N_29831,N_28469,N_28338);
nand U29832 (N_29832,N_28494,N_28598);
nand U29833 (N_29833,N_28855,N_28715);
nand U29834 (N_29834,N_28522,N_28458);
nand U29835 (N_29835,N_28037,N_28075);
nor U29836 (N_29836,N_28921,N_28489);
xnor U29837 (N_29837,N_28773,N_28928);
xnor U29838 (N_29838,N_28974,N_28890);
nand U29839 (N_29839,N_28920,N_28727);
and U29840 (N_29840,N_28970,N_28595);
and U29841 (N_29841,N_28760,N_28852);
or U29842 (N_29842,N_28563,N_28159);
and U29843 (N_29843,N_28558,N_28180);
or U29844 (N_29844,N_28326,N_28581);
xnor U29845 (N_29845,N_28690,N_28356);
or U29846 (N_29846,N_28928,N_28089);
and U29847 (N_29847,N_28770,N_28343);
nor U29848 (N_29848,N_28044,N_28259);
or U29849 (N_29849,N_28788,N_28170);
nand U29850 (N_29850,N_28774,N_28086);
nor U29851 (N_29851,N_28157,N_28582);
nor U29852 (N_29852,N_28444,N_28765);
nand U29853 (N_29853,N_28508,N_28848);
xor U29854 (N_29854,N_28516,N_28307);
or U29855 (N_29855,N_28690,N_28987);
xor U29856 (N_29856,N_28057,N_28115);
or U29857 (N_29857,N_28245,N_28800);
or U29858 (N_29858,N_28465,N_28283);
or U29859 (N_29859,N_28792,N_28648);
nand U29860 (N_29860,N_28972,N_28176);
or U29861 (N_29861,N_28501,N_28670);
and U29862 (N_29862,N_28635,N_28277);
or U29863 (N_29863,N_28708,N_28518);
or U29864 (N_29864,N_28899,N_28304);
xnor U29865 (N_29865,N_28414,N_28268);
nand U29866 (N_29866,N_28045,N_28747);
and U29867 (N_29867,N_28782,N_28094);
or U29868 (N_29868,N_28019,N_28031);
and U29869 (N_29869,N_28239,N_28329);
nor U29870 (N_29870,N_28764,N_28985);
nor U29871 (N_29871,N_28383,N_28186);
nor U29872 (N_29872,N_28337,N_28585);
and U29873 (N_29873,N_28438,N_28608);
xor U29874 (N_29874,N_28194,N_28480);
and U29875 (N_29875,N_28519,N_28084);
nor U29876 (N_29876,N_28129,N_28870);
nand U29877 (N_29877,N_28995,N_28414);
nor U29878 (N_29878,N_28756,N_28088);
nor U29879 (N_29879,N_28468,N_28158);
xor U29880 (N_29880,N_28697,N_28675);
xor U29881 (N_29881,N_28018,N_28585);
or U29882 (N_29882,N_28453,N_28489);
or U29883 (N_29883,N_28120,N_28684);
xor U29884 (N_29884,N_28053,N_28490);
or U29885 (N_29885,N_28040,N_28748);
nor U29886 (N_29886,N_28133,N_28836);
nand U29887 (N_29887,N_28570,N_28020);
xor U29888 (N_29888,N_28791,N_28739);
and U29889 (N_29889,N_28111,N_28893);
nor U29890 (N_29890,N_28819,N_28253);
or U29891 (N_29891,N_28406,N_28202);
and U29892 (N_29892,N_28670,N_28872);
or U29893 (N_29893,N_28315,N_28761);
or U29894 (N_29894,N_28404,N_28282);
or U29895 (N_29895,N_28771,N_28137);
nand U29896 (N_29896,N_28621,N_28366);
nand U29897 (N_29897,N_28211,N_28437);
or U29898 (N_29898,N_28251,N_28788);
nand U29899 (N_29899,N_28298,N_28631);
and U29900 (N_29900,N_28932,N_28587);
and U29901 (N_29901,N_28439,N_28089);
nand U29902 (N_29902,N_28723,N_28227);
nand U29903 (N_29903,N_28309,N_28382);
xor U29904 (N_29904,N_28261,N_28289);
nor U29905 (N_29905,N_28647,N_28227);
nor U29906 (N_29906,N_28459,N_28960);
nor U29907 (N_29907,N_28274,N_28259);
nor U29908 (N_29908,N_28344,N_28399);
nand U29909 (N_29909,N_28589,N_28508);
nor U29910 (N_29910,N_28187,N_28939);
nor U29911 (N_29911,N_28233,N_28843);
and U29912 (N_29912,N_28054,N_28097);
nand U29913 (N_29913,N_28496,N_28370);
nor U29914 (N_29914,N_28967,N_28215);
xnor U29915 (N_29915,N_28742,N_28357);
xnor U29916 (N_29916,N_28224,N_28670);
or U29917 (N_29917,N_28783,N_28960);
and U29918 (N_29918,N_28658,N_28346);
or U29919 (N_29919,N_28310,N_28241);
xor U29920 (N_29920,N_28631,N_28697);
or U29921 (N_29921,N_28660,N_28755);
nand U29922 (N_29922,N_28463,N_28887);
or U29923 (N_29923,N_28394,N_28909);
xor U29924 (N_29924,N_28456,N_28042);
nand U29925 (N_29925,N_28889,N_28886);
or U29926 (N_29926,N_28095,N_28059);
nand U29927 (N_29927,N_28244,N_28805);
or U29928 (N_29928,N_28761,N_28595);
or U29929 (N_29929,N_28482,N_28194);
nor U29930 (N_29930,N_28760,N_28068);
nor U29931 (N_29931,N_28543,N_28312);
nand U29932 (N_29932,N_28208,N_28138);
and U29933 (N_29933,N_28827,N_28174);
and U29934 (N_29934,N_28548,N_28188);
or U29935 (N_29935,N_28766,N_28343);
xor U29936 (N_29936,N_28238,N_28283);
xnor U29937 (N_29937,N_28816,N_28003);
nand U29938 (N_29938,N_28241,N_28153);
and U29939 (N_29939,N_28232,N_28621);
or U29940 (N_29940,N_28434,N_28774);
xor U29941 (N_29941,N_28489,N_28648);
and U29942 (N_29942,N_28337,N_28824);
nor U29943 (N_29943,N_28516,N_28496);
or U29944 (N_29944,N_28674,N_28678);
nand U29945 (N_29945,N_28088,N_28196);
nand U29946 (N_29946,N_28978,N_28966);
nor U29947 (N_29947,N_28267,N_28618);
and U29948 (N_29948,N_28124,N_28646);
and U29949 (N_29949,N_28443,N_28067);
and U29950 (N_29950,N_28935,N_28092);
nand U29951 (N_29951,N_28625,N_28589);
or U29952 (N_29952,N_28519,N_28700);
nand U29953 (N_29953,N_28788,N_28339);
and U29954 (N_29954,N_28649,N_28686);
and U29955 (N_29955,N_28360,N_28428);
nor U29956 (N_29956,N_28368,N_28766);
and U29957 (N_29957,N_28943,N_28833);
nand U29958 (N_29958,N_28668,N_28706);
nand U29959 (N_29959,N_28105,N_28630);
xnor U29960 (N_29960,N_28105,N_28891);
xnor U29961 (N_29961,N_28256,N_28349);
nand U29962 (N_29962,N_28137,N_28687);
nor U29963 (N_29963,N_28062,N_28410);
and U29964 (N_29964,N_28335,N_28079);
and U29965 (N_29965,N_28169,N_28228);
nor U29966 (N_29966,N_28886,N_28397);
xnor U29967 (N_29967,N_28674,N_28705);
nand U29968 (N_29968,N_28783,N_28134);
or U29969 (N_29969,N_28806,N_28023);
or U29970 (N_29970,N_28257,N_28514);
and U29971 (N_29971,N_28375,N_28167);
or U29972 (N_29972,N_28152,N_28119);
xor U29973 (N_29973,N_28858,N_28506);
and U29974 (N_29974,N_28288,N_28951);
xor U29975 (N_29975,N_28254,N_28982);
xnor U29976 (N_29976,N_28088,N_28920);
and U29977 (N_29977,N_28470,N_28257);
xor U29978 (N_29978,N_28868,N_28042);
nand U29979 (N_29979,N_28449,N_28663);
and U29980 (N_29980,N_28127,N_28215);
nor U29981 (N_29981,N_28319,N_28538);
nand U29982 (N_29982,N_28008,N_28619);
nor U29983 (N_29983,N_28310,N_28041);
nor U29984 (N_29984,N_28624,N_28059);
xnor U29985 (N_29985,N_28233,N_28745);
xnor U29986 (N_29986,N_28307,N_28797);
xnor U29987 (N_29987,N_28779,N_28503);
nand U29988 (N_29988,N_28080,N_28263);
and U29989 (N_29989,N_28948,N_28022);
and U29990 (N_29990,N_28830,N_28526);
nand U29991 (N_29991,N_28370,N_28166);
nor U29992 (N_29992,N_28741,N_28983);
nor U29993 (N_29993,N_28336,N_28233);
or U29994 (N_29994,N_28262,N_28320);
xnor U29995 (N_29995,N_28765,N_28379);
or U29996 (N_29996,N_28014,N_28651);
or U29997 (N_29997,N_28428,N_28036);
and U29998 (N_29998,N_28740,N_28394);
nand U29999 (N_29999,N_28591,N_28675);
or UO_0 (O_0,N_29703,N_29146);
or UO_1 (O_1,N_29214,N_29071);
nor UO_2 (O_2,N_29007,N_29283);
or UO_3 (O_3,N_29541,N_29873);
nor UO_4 (O_4,N_29940,N_29474);
or UO_5 (O_5,N_29516,N_29270);
and UO_6 (O_6,N_29257,N_29338);
or UO_7 (O_7,N_29596,N_29408);
xor UO_8 (O_8,N_29409,N_29597);
xnor UO_9 (O_9,N_29442,N_29754);
nand UO_10 (O_10,N_29160,N_29590);
nor UO_11 (O_11,N_29788,N_29238);
xor UO_12 (O_12,N_29499,N_29790);
nand UO_13 (O_13,N_29579,N_29535);
nand UO_14 (O_14,N_29655,N_29271);
nor UO_15 (O_15,N_29981,N_29433);
nand UO_16 (O_16,N_29704,N_29475);
nor UO_17 (O_17,N_29811,N_29679);
nand UO_18 (O_18,N_29642,N_29835);
or UO_19 (O_19,N_29781,N_29102);
nand UO_20 (O_20,N_29201,N_29227);
nand UO_21 (O_21,N_29936,N_29998);
nand UO_22 (O_22,N_29117,N_29090);
xor UO_23 (O_23,N_29309,N_29892);
nand UO_24 (O_24,N_29767,N_29101);
or UO_25 (O_25,N_29565,N_29743);
nor UO_26 (O_26,N_29511,N_29812);
nand UO_27 (O_27,N_29567,N_29387);
nor UO_28 (O_28,N_29691,N_29205);
and UO_29 (O_29,N_29164,N_29791);
nor UO_30 (O_30,N_29467,N_29198);
nor UO_31 (O_31,N_29777,N_29528);
or UO_32 (O_32,N_29938,N_29578);
nand UO_33 (O_33,N_29330,N_29285);
nor UO_34 (O_34,N_29478,N_29111);
xor UO_35 (O_35,N_29540,N_29080);
and UO_36 (O_36,N_29008,N_29904);
or UO_37 (O_37,N_29748,N_29605);
and UO_38 (O_38,N_29750,N_29557);
nor UO_39 (O_39,N_29424,N_29184);
or UO_40 (O_40,N_29952,N_29694);
nor UO_41 (O_41,N_29660,N_29696);
nor UO_42 (O_42,N_29416,N_29473);
nand UO_43 (O_43,N_29663,N_29291);
or UO_44 (O_44,N_29792,N_29664);
nor UO_45 (O_45,N_29690,N_29562);
nor UO_46 (O_46,N_29584,N_29367);
or UO_47 (O_47,N_29732,N_29156);
nand UO_48 (O_48,N_29358,N_29097);
nand UO_49 (O_49,N_29599,N_29228);
and UO_50 (O_50,N_29902,N_29573);
nor UO_51 (O_51,N_29108,N_29692);
xor UO_52 (O_52,N_29971,N_29901);
and UO_53 (O_53,N_29370,N_29091);
and UO_54 (O_54,N_29377,N_29799);
xor UO_55 (O_55,N_29569,N_29103);
xnor UO_56 (O_56,N_29880,N_29680);
nand UO_57 (O_57,N_29328,N_29980);
xnor UO_58 (O_58,N_29064,N_29946);
nor UO_59 (O_59,N_29994,N_29999);
and UO_60 (O_60,N_29484,N_29525);
or UO_61 (O_61,N_29341,N_29052);
and UO_62 (O_62,N_29073,N_29266);
xor UO_63 (O_63,N_29383,N_29045);
xnor UO_64 (O_64,N_29776,N_29864);
and UO_65 (O_65,N_29678,N_29624);
or UO_66 (O_66,N_29333,N_29162);
nor UO_67 (O_67,N_29316,N_29531);
nand UO_68 (O_68,N_29606,N_29312);
xnor UO_69 (O_69,N_29643,N_29012);
or UO_70 (O_70,N_29763,N_29191);
xnor UO_71 (O_71,N_29180,N_29138);
xnor UO_72 (O_72,N_29319,N_29029);
xor UO_73 (O_73,N_29657,N_29490);
nor UO_74 (O_74,N_29404,N_29883);
xor UO_75 (O_75,N_29051,N_29299);
and UO_76 (O_76,N_29083,N_29241);
xor UO_77 (O_77,N_29866,N_29953);
and UO_78 (O_78,N_29297,N_29494);
xnor UO_79 (O_79,N_29558,N_29681);
xor UO_80 (O_80,N_29857,N_29320);
nand UO_81 (O_81,N_29276,N_29649);
and UO_82 (O_82,N_29650,N_29860);
and UO_83 (O_83,N_29592,N_29523);
nor UO_84 (O_84,N_29355,N_29830);
nand UO_85 (O_85,N_29053,N_29104);
and UO_86 (O_86,N_29374,N_29089);
and UO_87 (O_87,N_29034,N_29190);
or UO_88 (O_88,N_29145,N_29520);
nor UO_89 (O_89,N_29448,N_29789);
and UO_90 (O_90,N_29121,N_29171);
xor UO_91 (O_91,N_29668,N_29816);
or UO_92 (O_92,N_29551,N_29095);
or UO_93 (O_93,N_29255,N_29046);
and UO_94 (O_94,N_29165,N_29826);
xnor UO_95 (O_95,N_29002,N_29471);
nand UO_96 (O_96,N_29422,N_29441);
nor UO_97 (O_97,N_29094,N_29311);
and UO_98 (O_98,N_29395,N_29348);
or UO_99 (O_99,N_29527,N_29303);
xnor UO_100 (O_100,N_29878,N_29990);
nor UO_101 (O_101,N_29161,N_29862);
xnor UO_102 (O_102,N_29962,N_29899);
nand UO_103 (O_103,N_29425,N_29059);
xnor UO_104 (O_104,N_29513,N_29518);
and UO_105 (O_105,N_29874,N_29751);
or UO_106 (O_106,N_29100,N_29344);
xor UO_107 (O_107,N_29538,N_29004);
xor UO_108 (O_108,N_29700,N_29987);
xnor UO_109 (O_109,N_29128,N_29598);
nand UO_110 (O_110,N_29495,N_29881);
xor UO_111 (O_111,N_29315,N_29509);
nand UO_112 (O_112,N_29675,N_29993);
or UO_113 (O_113,N_29390,N_29654);
xnor UO_114 (O_114,N_29983,N_29964);
or UO_115 (O_115,N_29453,N_29288);
xor UO_116 (O_116,N_29192,N_29773);
nor UO_117 (O_117,N_29212,N_29877);
or UO_118 (O_118,N_29069,N_29443);
and UO_119 (O_119,N_29419,N_29923);
xnor UO_120 (O_120,N_29208,N_29354);
nand UO_121 (O_121,N_29200,N_29553);
nand UO_122 (O_122,N_29202,N_29250);
xnor UO_123 (O_123,N_29852,N_29410);
nor UO_124 (O_124,N_29740,N_29610);
and UO_125 (O_125,N_29013,N_29614);
xnor UO_126 (O_126,N_29407,N_29019);
nand UO_127 (O_127,N_29403,N_29982);
or UO_128 (O_128,N_29226,N_29016);
and UO_129 (O_129,N_29033,N_29479);
or UO_130 (O_130,N_29697,N_29850);
or UO_131 (O_131,N_29457,N_29392);
and UO_132 (O_132,N_29504,N_29708);
nor UO_133 (O_133,N_29859,N_29028);
and UO_134 (O_134,N_29398,N_29638);
and UO_135 (O_135,N_29988,N_29339);
nor UO_136 (O_136,N_29258,N_29887);
xnor UO_137 (O_137,N_29332,N_29549);
and UO_138 (O_138,N_29782,N_29485);
nand UO_139 (O_139,N_29278,N_29463);
or UO_140 (O_140,N_29336,N_29764);
or UO_141 (O_141,N_29970,N_29742);
nor UO_142 (O_142,N_29583,N_29289);
or UO_143 (O_143,N_29203,N_29452);
and UO_144 (O_144,N_29559,N_29268);
xnor UO_145 (O_145,N_29867,N_29872);
xor UO_146 (O_146,N_29973,N_29353);
nor UO_147 (O_147,N_29948,N_29306);
or UO_148 (O_148,N_29845,N_29838);
xnor UO_149 (O_149,N_29672,N_29607);
xnor UO_150 (O_150,N_29593,N_29086);
or UO_151 (O_151,N_29526,N_29656);
xor UO_152 (O_152,N_29752,N_29294);
or UO_153 (O_153,N_29616,N_29913);
nor UO_154 (O_154,N_29956,N_29965);
and UO_155 (O_155,N_29840,N_29963);
xnor UO_156 (O_156,N_29658,N_29075);
or UO_157 (O_157,N_29861,N_29123);
or UO_158 (O_158,N_29224,N_29262);
nand UO_159 (O_159,N_29920,N_29252);
or UO_160 (O_160,N_29115,N_29134);
and UO_161 (O_161,N_29896,N_29888);
xnor UO_162 (O_162,N_29116,N_29307);
xnor UO_163 (O_163,N_29837,N_29369);
nor UO_164 (O_164,N_29216,N_29785);
or UO_165 (O_165,N_29924,N_29831);
nor UO_166 (O_166,N_29327,N_29093);
nor UO_167 (O_167,N_29155,N_29213);
xor UO_168 (O_168,N_29686,N_29730);
and UO_169 (O_169,N_29456,N_29177);
nor UO_170 (O_170,N_29937,N_29450);
xnor UO_171 (O_171,N_29843,N_29909);
nand UO_172 (O_172,N_29705,N_29635);
nand UO_173 (O_173,N_29817,N_29644);
nor UO_174 (O_174,N_29622,N_29098);
nand UO_175 (O_175,N_29243,N_29169);
and UO_176 (O_176,N_29698,N_29580);
or UO_177 (O_177,N_29186,N_29105);
nand UO_178 (O_178,N_29099,N_29591);
and UO_179 (O_179,N_29359,N_29613);
xnor UO_180 (O_180,N_29349,N_29361);
nand UO_181 (O_181,N_29157,N_29893);
nor UO_182 (O_182,N_29265,N_29652);
nand UO_183 (O_183,N_29173,N_29263);
nor UO_184 (O_184,N_29331,N_29682);
or UO_185 (O_185,N_29068,N_29805);
or UO_186 (O_186,N_29232,N_29346);
nand UO_187 (O_187,N_29056,N_29427);
nor UO_188 (O_188,N_29615,N_29949);
xnor UO_189 (O_189,N_29438,N_29154);
nor UO_190 (O_190,N_29756,N_29833);
or UO_191 (O_191,N_29659,N_29461);
xor UO_192 (O_192,N_29677,N_29889);
nand UO_193 (O_193,N_29293,N_29945);
xnor UO_194 (O_194,N_29365,N_29941);
and UO_195 (O_195,N_29290,N_29914);
nand UO_196 (O_196,N_29564,N_29426);
nand UO_197 (O_197,N_29897,N_29421);
nand UO_198 (O_198,N_29062,N_29806);
nor UO_199 (O_199,N_29211,N_29249);
nor UO_200 (O_200,N_29127,N_29739);
nand UO_201 (O_201,N_29611,N_29366);
nor UO_202 (O_202,N_29026,N_29771);
and UO_203 (O_203,N_29882,N_29502);
xnor UO_204 (O_204,N_29176,N_29522);
xor UO_205 (O_205,N_29295,N_29023);
nor UO_206 (O_206,N_29183,N_29620);
or UO_207 (O_207,N_29738,N_29042);
and UO_208 (O_208,N_29505,N_29546);
nor UO_209 (O_209,N_29119,N_29021);
or UO_210 (O_210,N_29025,N_29038);
and UO_211 (O_211,N_29813,N_29414);
and UO_212 (O_212,N_29930,N_29723);
and UO_213 (O_213,N_29084,N_29239);
nor UO_214 (O_214,N_29735,N_29712);
nor UO_215 (O_215,N_29429,N_29491);
nor UO_216 (O_216,N_29542,N_29997);
and UO_217 (O_217,N_29574,N_29632);
or UO_218 (O_218,N_29444,N_29150);
nand UO_219 (O_219,N_29780,N_29519);
nand UO_220 (O_220,N_29736,N_29006);
and UO_221 (O_221,N_29181,N_29215);
and UO_222 (O_222,N_29666,N_29770);
xor UO_223 (O_223,N_29532,N_29379);
nand UO_224 (O_224,N_29136,N_29876);
or UO_225 (O_225,N_29326,N_29199);
nor UO_226 (O_226,N_29508,N_29633);
and UO_227 (O_227,N_29714,N_29020);
nor UO_228 (O_228,N_29818,N_29178);
xnor UO_229 (O_229,N_29507,N_29462);
nand UO_230 (O_230,N_29281,N_29910);
nand UO_231 (O_231,N_29784,N_29233);
or UO_232 (O_232,N_29547,N_29220);
or UO_233 (O_233,N_29808,N_29489);
nand UO_234 (O_234,N_29032,N_29533);
and UO_235 (O_235,N_29217,N_29786);
and UO_236 (O_236,N_29761,N_29844);
xnor UO_237 (O_237,N_29651,N_29648);
or UO_238 (O_238,N_29741,N_29142);
and UO_239 (O_239,N_29903,N_29572);
xnor UO_240 (O_240,N_29645,N_29063);
nand UO_241 (O_241,N_29125,N_29386);
and UO_242 (O_242,N_29231,N_29885);
or UO_243 (O_243,N_29219,N_29894);
and UO_244 (O_244,N_29673,N_29394);
xnor UO_245 (O_245,N_29148,N_29364);
xnor UO_246 (O_246,N_29802,N_29637);
and UO_247 (O_247,N_29468,N_29017);
nand UO_248 (O_248,N_29236,N_29561);
nand UO_249 (O_249,N_29976,N_29800);
xnor UO_250 (O_250,N_29197,N_29718);
or UO_251 (O_251,N_29676,N_29131);
xnor UO_252 (O_252,N_29671,N_29552);
nor UO_253 (O_253,N_29277,N_29420);
nor UO_254 (O_254,N_29856,N_29688);
or UO_255 (O_255,N_29476,N_29586);
or UO_256 (O_256,N_29259,N_29550);
nand UO_257 (O_257,N_29477,N_29310);
and UO_258 (O_258,N_29720,N_29144);
nor UO_259 (O_259,N_29139,N_29796);
or UO_260 (O_260,N_29768,N_29839);
or UO_261 (O_261,N_29737,N_29702);
nand UO_262 (O_262,N_29109,N_29524);
xor UO_263 (O_263,N_29585,N_29459);
xor UO_264 (O_264,N_29603,N_29396);
nand UO_265 (O_265,N_29061,N_29325);
or UO_266 (O_266,N_29388,N_29906);
xnor UO_267 (O_267,N_29449,N_29218);
and UO_268 (O_268,N_29435,N_29261);
and UO_269 (O_269,N_29634,N_29891);
xnor UO_270 (O_270,N_29929,N_29604);
nor UO_271 (O_271,N_29168,N_29853);
and UO_272 (O_272,N_29003,N_29253);
or UO_273 (O_273,N_29375,N_29048);
nand UO_274 (O_274,N_29382,N_29054);
or UO_275 (O_275,N_29418,N_29464);
nand UO_276 (O_276,N_29158,N_29322);
or UO_277 (O_277,N_29577,N_29699);
and UO_278 (O_278,N_29731,N_29626);
or UO_279 (O_279,N_29821,N_29521);
xor UO_280 (O_280,N_29350,N_29984);
nor UO_281 (O_281,N_29933,N_29460);
nand UO_282 (O_282,N_29907,N_29167);
and UO_283 (O_283,N_29384,N_29163);
and UO_284 (O_284,N_29766,N_29934);
nand UO_285 (O_285,N_29989,N_29807);
or UO_286 (O_286,N_29269,N_29015);
nor UO_287 (O_287,N_29066,N_29267);
or UO_288 (O_288,N_29943,N_29222);
nand UO_289 (O_289,N_29027,N_29472);
xnor UO_290 (O_290,N_29264,N_29589);
or UO_291 (O_291,N_29566,N_29935);
nor UO_292 (O_292,N_29728,N_29405);
and UO_293 (O_293,N_29762,N_29921);
nor UO_294 (O_294,N_29035,N_29724);
and UO_295 (O_295,N_29313,N_29402);
xor UO_296 (O_296,N_29113,N_29321);
or UO_297 (O_297,N_29665,N_29244);
nor UO_298 (O_298,N_29423,N_29129);
and UO_299 (O_299,N_29506,N_29143);
nand UO_300 (O_300,N_29196,N_29337);
nor UO_301 (O_301,N_29568,N_29439);
nand UO_302 (O_302,N_29667,N_29234);
xor UO_303 (O_303,N_29855,N_29814);
xor UO_304 (O_304,N_29555,N_29049);
or UO_305 (O_305,N_29778,N_29760);
or UO_306 (O_306,N_29352,N_29147);
nor UO_307 (O_307,N_29324,N_29030);
nand UO_308 (O_308,N_29246,N_29576);
xor UO_309 (O_309,N_29137,N_29272);
xor UO_310 (O_310,N_29815,N_29371);
nor UO_311 (O_311,N_29001,N_29685);
and UO_312 (O_312,N_29040,N_29480);
nor UO_313 (O_313,N_29329,N_29210);
and UO_314 (O_314,N_29503,N_29908);
nor UO_315 (O_315,N_29759,N_29966);
and UO_316 (O_316,N_29022,N_29978);
and UO_317 (O_317,N_29674,N_29399);
xnor UO_318 (O_318,N_29570,N_29957);
nand UO_319 (O_319,N_29545,N_29820);
nor UO_320 (O_320,N_29755,N_29380);
or UO_321 (O_321,N_29847,N_29958);
nor UO_322 (O_322,N_29483,N_29193);
nand UO_323 (O_323,N_29298,N_29058);
and UO_324 (O_324,N_29969,N_29848);
and UO_325 (O_325,N_29078,N_29070);
and UO_326 (O_326,N_29135,N_29188);
nand UO_327 (O_327,N_29662,N_29846);
and UO_328 (O_328,N_29915,N_29627);
nor UO_329 (O_329,N_29305,N_29230);
or UO_330 (O_330,N_29260,N_29895);
nand UO_331 (O_331,N_29757,N_29719);
and UO_332 (O_332,N_29345,N_29721);
xor UO_333 (O_333,N_29587,N_29254);
or UO_334 (O_334,N_29000,N_29646);
xnor UO_335 (O_335,N_29979,N_29927);
nand UO_336 (O_336,N_29302,N_29729);
nand UO_337 (O_337,N_29653,N_29343);
xor UO_338 (O_338,N_29492,N_29563);
nand UO_339 (O_339,N_29082,N_29974);
nand UO_340 (O_340,N_29235,N_29661);
nor UO_341 (O_341,N_29977,N_29087);
xor UO_342 (O_342,N_29194,N_29795);
and UO_343 (O_343,N_29543,N_29010);
xor UO_344 (O_344,N_29640,N_29372);
nor UO_345 (O_345,N_29709,N_29209);
nor UO_346 (O_346,N_29282,N_29798);
or UO_347 (O_347,N_29400,N_29065);
or UO_348 (O_348,N_29401,N_29865);
or UO_349 (O_349,N_29548,N_29713);
and UO_350 (O_350,N_29207,N_29451);
or UO_351 (O_351,N_29044,N_29018);
nand UO_352 (O_352,N_29446,N_29362);
and UO_353 (O_353,N_29482,N_29465);
nand UO_354 (O_354,N_29669,N_29152);
nor UO_355 (O_355,N_29769,N_29629);
or UO_356 (O_356,N_29793,N_29871);
nand UO_357 (O_357,N_29529,N_29037);
and UO_358 (O_358,N_29618,N_29916);
nor UO_359 (O_359,N_29693,N_29985);
or UO_360 (O_360,N_29500,N_29179);
xnor UO_361 (O_361,N_29092,N_29783);
nand UO_362 (O_362,N_29917,N_29995);
or UO_363 (O_363,N_29647,N_29067);
xor UO_364 (O_364,N_29469,N_29274);
or UO_365 (O_365,N_29991,N_29753);
nor UO_366 (O_366,N_29628,N_29011);
nor UO_367 (O_367,N_29534,N_29836);
xor UO_368 (O_368,N_29050,N_29487);
or UO_369 (O_369,N_29342,N_29076);
nor UO_370 (O_370,N_29470,N_29112);
and UO_371 (O_371,N_29493,N_29955);
xor UO_372 (O_372,N_29107,N_29251);
and UO_373 (O_373,N_29858,N_29120);
xor UO_374 (O_374,N_29706,N_29911);
or UO_375 (O_375,N_29932,N_29581);
xor UO_376 (O_376,N_29195,N_29114);
nor UO_377 (O_377,N_29986,N_29928);
nor UO_378 (O_378,N_29077,N_29481);
and UO_379 (O_379,N_29544,N_29747);
nand UO_380 (O_380,N_29722,N_29707);
nand UO_381 (O_381,N_29630,N_29926);
or UO_382 (O_382,N_29804,N_29683);
xor UO_383 (O_383,N_29560,N_29055);
or UO_384 (O_384,N_29595,N_29151);
nor UO_385 (O_385,N_29832,N_29849);
xnor UO_386 (O_386,N_29950,N_29823);
nand UO_387 (O_387,N_29571,N_29774);
xor UO_388 (O_388,N_29072,N_29140);
and UO_389 (O_389,N_29787,N_29918);
and UO_390 (O_390,N_29824,N_29968);
or UO_391 (O_391,N_29153,N_29539);
nor UO_392 (O_392,N_29744,N_29636);
and UO_393 (O_393,N_29851,N_29185);
nor UO_394 (O_394,N_29256,N_29868);
nand UO_395 (O_395,N_29841,N_29514);
and UO_396 (O_396,N_29381,N_29014);
nor UO_397 (O_397,N_29711,N_29189);
and UO_398 (O_398,N_29939,N_29623);
nand UO_399 (O_399,N_29286,N_29890);
or UO_400 (O_400,N_29466,N_29110);
nor UO_401 (O_401,N_29166,N_29360);
nor UO_402 (O_402,N_29351,N_29081);
nor UO_403 (O_403,N_29869,N_29716);
xnor UO_404 (O_404,N_29822,N_29292);
and UO_405 (O_405,N_29397,N_29515);
nor UO_406 (O_406,N_29436,N_29005);
nor UO_407 (O_407,N_29944,N_29828);
nor UO_408 (O_408,N_29608,N_29710);
or UO_409 (O_409,N_29954,N_29794);
or UO_410 (O_410,N_29919,N_29556);
and UO_411 (O_411,N_29801,N_29440);
xnor UO_412 (O_412,N_29536,N_29886);
xnor UO_413 (O_413,N_29393,N_29308);
or UO_414 (O_414,N_29273,N_29187);
or UO_415 (O_415,N_29417,N_29925);
or UO_416 (O_416,N_29905,N_29854);
nand UO_417 (O_417,N_29582,N_29225);
xnor UO_418 (O_418,N_29746,N_29124);
nor UO_419 (O_419,N_29879,N_29819);
xor UO_420 (O_420,N_29942,N_29863);
nor UO_421 (O_421,N_29842,N_29458);
nand UO_422 (O_422,N_29726,N_29411);
nand UO_423 (O_423,N_29174,N_29088);
and UO_424 (O_424,N_29300,N_29149);
nor UO_425 (O_425,N_29340,N_29412);
and UO_426 (O_426,N_29530,N_29074);
and UO_427 (O_427,N_29619,N_29132);
nor UO_428 (O_428,N_29415,N_29368);
and UO_429 (O_429,N_29900,N_29301);
nand UO_430 (O_430,N_29175,N_29378);
nor UO_431 (O_431,N_29275,N_29237);
xnor UO_432 (O_432,N_29024,N_29617);
and UO_433 (O_433,N_29284,N_29829);
and UO_434 (O_434,N_29413,N_29041);
nor UO_435 (O_435,N_29600,N_29625);
and UO_436 (O_436,N_29715,N_29947);
nor UO_437 (O_437,N_29898,N_29510);
nand UO_438 (O_438,N_29182,N_29159);
and UO_439 (O_439,N_29363,N_29959);
and UO_440 (O_440,N_29870,N_29687);
or UO_441 (O_441,N_29554,N_29631);
xor UO_442 (O_442,N_29172,N_29118);
nor UO_443 (O_443,N_29335,N_29512);
nand UO_444 (O_444,N_29039,N_29447);
xnor UO_445 (O_445,N_29827,N_29498);
nor UO_446 (O_446,N_29280,N_29803);
nand UO_447 (O_447,N_29323,N_29304);
nor UO_448 (O_448,N_29223,N_29996);
nor UO_449 (O_449,N_29057,N_29130);
and UO_450 (O_450,N_29695,N_29612);
nor UO_451 (O_451,N_29609,N_29141);
nor UO_452 (O_452,N_29437,N_29242);
nor UO_453 (O_453,N_29621,N_29961);
xnor UO_454 (O_454,N_29975,N_29497);
and UO_455 (O_455,N_29825,N_29031);
nand UO_456 (O_456,N_29106,N_29967);
nand UO_457 (O_457,N_29455,N_29391);
and UO_458 (O_458,N_29079,N_29318);
nand UO_459 (O_459,N_29248,N_29431);
xnor UO_460 (O_460,N_29749,N_29501);
nor UO_461 (O_461,N_29486,N_29357);
or UO_462 (O_462,N_29245,N_29972);
or UO_463 (O_463,N_29204,N_29060);
nand UO_464 (O_464,N_29389,N_29588);
and UO_465 (O_465,N_29356,N_29279);
nand UO_466 (O_466,N_29085,N_29247);
xnor UO_467 (O_467,N_29575,N_29096);
and UO_468 (O_468,N_29601,N_29745);
and UO_469 (O_469,N_29434,N_29960);
xnor UO_470 (O_470,N_29314,N_29884);
nand UO_471 (O_471,N_29373,N_29594);
or UO_472 (O_472,N_29133,N_29517);
nor UO_473 (O_473,N_29912,N_29775);
nor UO_474 (O_474,N_29334,N_29043);
or UO_475 (O_475,N_29376,N_29922);
or UO_476 (O_476,N_29670,N_29797);
and UO_477 (O_477,N_29809,N_29834);
or UO_478 (O_478,N_29772,N_29428);
nor UO_479 (O_479,N_29206,N_29689);
nand UO_480 (O_480,N_29684,N_29641);
or UO_481 (O_481,N_29122,N_29454);
xnor UO_482 (O_482,N_29229,N_29727);
and UO_483 (O_483,N_29725,N_29036);
nand UO_484 (O_484,N_29221,N_29488);
and UO_485 (O_485,N_29445,N_29779);
or UO_486 (O_486,N_29734,N_29385);
nor UO_487 (O_487,N_29931,N_29287);
xor UO_488 (O_488,N_29406,N_29602);
xor UO_489 (O_489,N_29733,N_29317);
or UO_490 (O_490,N_29537,N_29992);
nor UO_491 (O_491,N_29717,N_29432);
or UO_492 (O_492,N_29347,N_29639);
xnor UO_493 (O_493,N_29875,N_29296);
xnor UO_494 (O_494,N_29701,N_29758);
nand UO_495 (O_495,N_29126,N_29047);
and UO_496 (O_496,N_29240,N_29170);
nand UO_497 (O_497,N_29765,N_29430);
nor UO_498 (O_498,N_29951,N_29009);
xor UO_499 (O_499,N_29496,N_29810);
and UO_500 (O_500,N_29686,N_29114);
nand UO_501 (O_501,N_29503,N_29624);
nand UO_502 (O_502,N_29683,N_29042);
or UO_503 (O_503,N_29507,N_29918);
xnor UO_504 (O_504,N_29309,N_29207);
or UO_505 (O_505,N_29433,N_29792);
xor UO_506 (O_506,N_29508,N_29081);
xor UO_507 (O_507,N_29526,N_29239);
nand UO_508 (O_508,N_29110,N_29817);
nand UO_509 (O_509,N_29345,N_29383);
and UO_510 (O_510,N_29226,N_29498);
or UO_511 (O_511,N_29191,N_29224);
nand UO_512 (O_512,N_29582,N_29733);
and UO_513 (O_513,N_29675,N_29561);
nor UO_514 (O_514,N_29984,N_29132);
nor UO_515 (O_515,N_29843,N_29818);
nand UO_516 (O_516,N_29052,N_29423);
xor UO_517 (O_517,N_29198,N_29229);
or UO_518 (O_518,N_29990,N_29395);
nand UO_519 (O_519,N_29170,N_29735);
and UO_520 (O_520,N_29437,N_29209);
xor UO_521 (O_521,N_29314,N_29443);
nand UO_522 (O_522,N_29881,N_29386);
xnor UO_523 (O_523,N_29983,N_29164);
xnor UO_524 (O_524,N_29114,N_29050);
or UO_525 (O_525,N_29469,N_29923);
nand UO_526 (O_526,N_29476,N_29068);
and UO_527 (O_527,N_29515,N_29021);
or UO_528 (O_528,N_29134,N_29506);
xor UO_529 (O_529,N_29997,N_29571);
nand UO_530 (O_530,N_29737,N_29209);
xor UO_531 (O_531,N_29470,N_29186);
xnor UO_532 (O_532,N_29929,N_29784);
xor UO_533 (O_533,N_29494,N_29980);
and UO_534 (O_534,N_29110,N_29356);
or UO_535 (O_535,N_29193,N_29247);
nand UO_536 (O_536,N_29513,N_29126);
nor UO_537 (O_537,N_29632,N_29300);
or UO_538 (O_538,N_29459,N_29292);
nor UO_539 (O_539,N_29325,N_29171);
or UO_540 (O_540,N_29230,N_29482);
xor UO_541 (O_541,N_29648,N_29978);
xor UO_542 (O_542,N_29235,N_29768);
nor UO_543 (O_543,N_29162,N_29033);
xor UO_544 (O_544,N_29545,N_29957);
xor UO_545 (O_545,N_29861,N_29597);
nor UO_546 (O_546,N_29137,N_29648);
xnor UO_547 (O_547,N_29859,N_29316);
and UO_548 (O_548,N_29100,N_29479);
xor UO_549 (O_549,N_29333,N_29639);
nor UO_550 (O_550,N_29293,N_29428);
nand UO_551 (O_551,N_29908,N_29421);
nor UO_552 (O_552,N_29684,N_29450);
nor UO_553 (O_553,N_29896,N_29368);
nor UO_554 (O_554,N_29971,N_29609);
nor UO_555 (O_555,N_29440,N_29333);
nor UO_556 (O_556,N_29520,N_29725);
and UO_557 (O_557,N_29481,N_29619);
nor UO_558 (O_558,N_29910,N_29703);
and UO_559 (O_559,N_29960,N_29069);
xnor UO_560 (O_560,N_29389,N_29688);
xnor UO_561 (O_561,N_29118,N_29251);
and UO_562 (O_562,N_29748,N_29366);
xor UO_563 (O_563,N_29115,N_29196);
xnor UO_564 (O_564,N_29300,N_29530);
xor UO_565 (O_565,N_29971,N_29198);
or UO_566 (O_566,N_29552,N_29115);
nand UO_567 (O_567,N_29709,N_29256);
or UO_568 (O_568,N_29821,N_29610);
nand UO_569 (O_569,N_29894,N_29917);
or UO_570 (O_570,N_29498,N_29992);
xnor UO_571 (O_571,N_29471,N_29253);
and UO_572 (O_572,N_29767,N_29169);
and UO_573 (O_573,N_29926,N_29405);
nand UO_574 (O_574,N_29223,N_29334);
nand UO_575 (O_575,N_29071,N_29354);
and UO_576 (O_576,N_29214,N_29346);
or UO_577 (O_577,N_29521,N_29946);
nor UO_578 (O_578,N_29606,N_29445);
nor UO_579 (O_579,N_29540,N_29912);
nand UO_580 (O_580,N_29862,N_29659);
xor UO_581 (O_581,N_29570,N_29574);
and UO_582 (O_582,N_29184,N_29929);
xnor UO_583 (O_583,N_29587,N_29655);
nor UO_584 (O_584,N_29628,N_29324);
nand UO_585 (O_585,N_29931,N_29822);
nand UO_586 (O_586,N_29192,N_29751);
xnor UO_587 (O_587,N_29067,N_29128);
nand UO_588 (O_588,N_29577,N_29394);
nand UO_589 (O_589,N_29653,N_29738);
xor UO_590 (O_590,N_29779,N_29295);
and UO_591 (O_591,N_29805,N_29427);
nor UO_592 (O_592,N_29452,N_29353);
nand UO_593 (O_593,N_29866,N_29580);
nor UO_594 (O_594,N_29814,N_29487);
and UO_595 (O_595,N_29113,N_29687);
nand UO_596 (O_596,N_29580,N_29919);
nand UO_597 (O_597,N_29399,N_29789);
nor UO_598 (O_598,N_29531,N_29416);
or UO_599 (O_599,N_29402,N_29881);
and UO_600 (O_600,N_29545,N_29927);
nand UO_601 (O_601,N_29075,N_29458);
or UO_602 (O_602,N_29458,N_29481);
or UO_603 (O_603,N_29511,N_29516);
xnor UO_604 (O_604,N_29976,N_29625);
xor UO_605 (O_605,N_29373,N_29855);
nand UO_606 (O_606,N_29879,N_29786);
nand UO_607 (O_607,N_29633,N_29148);
and UO_608 (O_608,N_29461,N_29935);
nand UO_609 (O_609,N_29688,N_29783);
nand UO_610 (O_610,N_29791,N_29314);
or UO_611 (O_611,N_29698,N_29289);
nor UO_612 (O_612,N_29897,N_29734);
nor UO_613 (O_613,N_29249,N_29787);
nand UO_614 (O_614,N_29515,N_29220);
or UO_615 (O_615,N_29755,N_29508);
and UO_616 (O_616,N_29812,N_29768);
nand UO_617 (O_617,N_29919,N_29461);
xnor UO_618 (O_618,N_29199,N_29184);
nor UO_619 (O_619,N_29770,N_29959);
xor UO_620 (O_620,N_29559,N_29347);
or UO_621 (O_621,N_29269,N_29323);
nand UO_622 (O_622,N_29368,N_29374);
xnor UO_623 (O_623,N_29338,N_29198);
nor UO_624 (O_624,N_29301,N_29263);
xnor UO_625 (O_625,N_29169,N_29590);
or UO_626 (O_626,N_29378,N_29181);
or UO_627 (O_627,N_29568,N_29057);
or UO_628 (O_628,N_29692,N_29225);
or UO_629 (O_629,N_29202,N_29617);
nor UO_630 (O_630,N_29234,N_29928);
and UO_631 (O_631,N_29147,N_29016);
and UO_632 (O_632,N_29261,N_29131);
xor UO_633 (O_633,N_29114,N_29288);
nor UO_634 (O_634,N_29864,N_29259);
or UO_635 (O_635,N_29707,N_29144);
nor UO_636 (O_636,N_29910,N_29995);
and UO_637 (O_637,N_29195,N_29271);
and UO_638 (O_638,N_29995,N_29882);
nor UO_639 (O_639,N_29310,N_29110);
or UO_640 (O_640,N_29861,N_29440);
nor UO_641 (O_641,N_29898,N_29255);
and UO_642 (O_642,N_29101,N_29660);
or UO_643 (O_643,N_29192,N_29233);
nor UO_644 (O_644,N_29434,N_29883);
nor UO_645 (O_645,N_29502,N_29813);
or UO_646 (O_646,N_29594,N_29024);
xor UO_647 (O_647,N_29472,N_29847);
and UO_648 (O_648,N_29819,N_29646);
xnor UO_649 (O_649,N_29750,N_29279);
and UO_650 (O_650,N_29391,N_29395);
or UO_651 (O_651,N_29359,N_29597);
nor UO_652 (O_652,N_29239,N_29090);
and UO_653 (O_653,N_29613,N_29144);
nor UO_654 (O_654,N_29962,N_29403);
xnor UO_655 (O_655,N_29140,N_29133);
and UO_656 (O_656,N_29256,N_29436);
and UO_657 (O_657,N_29052,N_29545);
or UO_658 (O_658,N_29617,N_29604);
or UO_659 (O_659,N_29635,N_29701);
nor UO_660 (O_660,N_29459,N_29166);
nor UO_661 (O_661,N_29260,N_29750);
xor UO_662 (O_662,N_29599,N_29162);
nand UO_663 (O_663,N_29100,N_29621);
or UO_664 (O_664,N_29120,N_29133);
nand UO_665 (O_665,N_29877,N_29487);
nand UO_666 (O_666,N_29092,N_29218);
nand UO_667 (O_667,N_29114,N_29512);
or UO_668 (O_668,N_29237,N_29491);
nand UO_669 (O_669,N_29191,N_29338);
nor UO_670 (O_670,N_29525,N_29740);
or UO_671 (O_671,N_29642,N_29532);
xor UO_672 (O_672,N_29233,N_29967);
nor UO_673 (O_673,N_29521,N_29530);
xor UO_674 (O_674,N_29901,N_29157);
and UO_675 (O_675,N_29230,N_29452);
or UO_676 (O_676,N_29298,N_29322);
or UO_677 (O_677,N_29429,N_29290);
xnor UO_678 (O_678,N_29357,N_29059);
or UO_679 (O_679,N_29826,N_29031);
nand UO_680 (O_680,N_29104,N_29632);
xor UO_681 (O_681,N_29811,N_29275);
nand UO_682 (O_682,N_29827,N_29509);
or UO_683 (O_683,N_29407,N_29390);
and UO_684 (O_684,N_29085,N_29214);
xnor UO_685 (O_685,N_29163,N_29735);
nor UO_686 (O_686,N_29460,N_29267);
nor UO_687 (O_687,N_29320,N_29928);
xnor UO_688 (O_688,N_29891,N_29678);
or UO_689 (O_689,N_29263,N_29149);
and UO_690 (O_690,N_29016,N_29751);
xor UO_691 (O_691,N_29689,N_29189);
or UO_692 (O_692,N_29732,N_29315);
or UO_693 (O_693,N_29847,N_29056);
nand UO_694 (O_694,N_29376,N_29409);
xor UO_695 (O_695,N_29931,N_29697);
nand UO_696 (O_696,N_29022,N_29713);
nand UO_697 (O_697,N_29391,N_29173);
nand UO_698 (O_698,N_29839,N_29135);
nand UO_699 (O_699,N_29509,N_29947);
and UO_700 (O_700,N_29767,N_29431);
nand UO_701 (O_701,N_29800,N_29013);
xnor UO_702 (O_702,N_29316,N_29646);
xnor UO_703 (O_703,N_29457,N_29298);
or UO_704 (O_704,N_29628,N_29704);
or UO_705 (O_705,N_29897,N_29236);
nor UO_706 (O_706,N_29951,N_29055);
nor UO_707 (O_707,N_29332,N_29202);
and UO_708 (O_708,N_29928,N_29101);
nor UO_709 (O_709,N_29516,N_29588);
nand UO_710 (O_710,N_29012,N_29861);
nor UO_711 (O_711,N_29665,N_29085);
or UO_712 (O_712,N_29105,N_29260);
nand UO_713 (O_713,N_29433,N_29284);
and UO_714 (O_714,N_29854,N_29455);
and UO_715 (O_715,N_29006,N_29770);
nand UO_716 (O_716,N_29120,N_29621);
nand UO_717 (O_717,N_29092,N_29860);
and UO_718 (O_718,N_29820,N_29768);
nor UO_719 (O_719,N_29446,N_29342);
xnor UO_720 (O_720,N_29476,N_29414);
and UO_721 (O_721,N_29099,N_29656);
xor UO_722 (O_722,N_29817,N_29841);
or UO_723 (O_723,N_29196,N_29566);
or UO_724 (O_724,N_29296,N_29248);
nor UO_725 (O_725,N_29343,N_29858);
and UO_726 (O_726,N_29269,N_29542);
nor UO_727 (O_727,N_29193,N_29963);
nor UO_728 (O_728,N_29637,N_29885);
nor UO_729 (O_729,N_29728,N_29242);
and UO_730 (O_730,N_29941,N_29800);
xor UO_731 (O_731,N_29161,N_29064);
nand UO_732 (O_732,N_29545,N_29879);
or UO_733 (O_733,N_29267,N_29943);
xor UO_734 (O_734,N_29250,N_29436);
and UO_735 (O_735,N_29645,N_29748);
or UO_736 (O_736,N_29858,N_29634);
nand UO_737 (O_737,N_29409,N_29086);
or UO_738 (O_738,N_29149,N_29555);
and UO_739 (O_739,N_29332,N_29564);
nor UO_740 (O_740,N_29997,N_29726);
or UO_741 (O_741,N_29929,N_29575);
nor UO_742 (O_742,N_29880,N_29885);
nand UO_743 (O_743,N_29928,N_29580);
nor UO_744 (O_744,N_29611,N_29898);
nand UO_745 (O_745,N_29864,N_29984);
and UO_746 (O_746,N_29095,N_29795);
and UO_747 (O_747,N_29526,N_29686);
nor UO_748 (O_748,N_29868,N_29294);
xor UO_749 (O_749,N_29670,N_29139);
and UO_750 (O_750,N_29176,N_29546);
nor UO_751 (O_751,N_29085,N_29830);
or UO_752 (O_752,N_29934,N_29085);
nand UO_753 (O_753,N_29403,N_29984);
and UO_754 (O_754,N_29505,N_29816);
nor UO_755 (O_755,N_29923,N_29871);
and UO_756 (O_756,N_29997,N_29151);
and UO_757 (O_757,N_29567,N_29261);
or UO_758 (O_758,N_29925,N_29151);
or UO_759 (O_759,N_29010,N_29631);
or UO_760 (O_760,N_29683,N_29842);
nor UO_761 (O_761,N_29842,N_29782);
xor UO_762 (O_762,N_29987,N_29432);
nor UO_763 (O_763,N_29700,N_29348);
or UO_764 (O_764,N_29512,N_29784);
xor UO_765 (O_765,N_29204,N_29772);
or UO_766 (O_766,N_29136,N_29195);
nand UO_767 (O_767,N_29699,N_29381);
and UO_768 (O_768,N_29526,N_29934);
nor UO_769 (O_769,N_29418,N_29740);
xor UO_770 (O_770,N_29764,N_29195);
nor UO_771 (O_771,N_29442,N_29122);
and UO_772 (O_772,N_29023,N_29031);
xor UO_773 (O_773,N_29818,N_29783);
nor UO_774 (O_774,N_29938,N_29066);
and UO_775 (O_775,N_29266,N_29899);
nand UO_776 (O_776,N_29531,N_29805);
or UO_777 (O_777,N_29787,N_29838);
nor UO_778 (O_778,N_29859,N_29942);
and UO_779 (O_779,N_29750,N_29445);
or UO_780 (O_780,N_29600,N_29773);
or UO_781 (O_781,N_29858,N_29986);
nand UO_782 (O_782,N_29060,N_29542);
and UO_783 (O_783,N_29028,N_29867);
nand UO_784 (O_784,N_29776,N_29061);
or UO_785 (O_785,N_29665,N_29886);
and UO_786 (O_786,N_29578,N_29671);
and UO_787 (O_787,N_29969,N_29806);
or UO_788 (O_788,N_29841,N_29142);
xor UO_789 (O_789,N_29160,N_29942);
or UO_790 (O_790,N_29986,N_29937);
nor UO_791 (O_791,N_29390,N_29713);
xor UO_792 (O_792,N_29046,N_29761);
or UO_793 (O_793,N_29742,N_29023);
nor UO_794 (O_794,N_29646,N_29185);
or UO_795 (O_795,N_29280,N_29388);
xnor UO_796 (O_796,N_29600,N_29365);
nand UO_797 (O_797,N_29416,N_29513);
or UO_798 (O_798,N_29025,N_29227);
nor UO_799 (O_799,N_29973,N_29643);
and UO_800 (O_800,N_29764,N_29005);
nand UO_801 (O_801,N_29874,N_29535);
xor UO_802 (O_802,N_29501,N_29947);
or UO_803 (O_803,N_29351,N_29426);
nand UO_804 (O_804,N_29431,N_29028);
or UO_805 (O_805,N_29038,N_29858);
nor UO_806 (O_806,N_29365,N_29139);
xnor UO_807 (O_807,N_29622,N_29551);
and UO_808 (O_808,N_29344,N_29797);
nor UO_809 (O_809,N_29721,N_29759);
and UO_810 (O_810,N_29634,N_29797);
and UO_811 (O_811,N_29800,N_29267);
or UO_812 (O_812,N_29081,N_29804);
xnor UO_813 (O_813,N_29122,N_29362);
nand UO_814 (O_814,N_29205,N_29536);
xnor UO_815 (O_815,N_29031,N_29006);
xor UO_816 (O_816,N_29370,N_29129);
or UO_817 (O_817,N_29753,N_29868);
nor UO_818 (O_818,N_29781,N_29311);
and UO_819 (O_819,N_29813,N_29890);
xor UO_820 (O_820,N_29926,N_29790);
nand UO_821 (O_821,N_29478,N_29099);
nand UO_822 (O_822,N_29865,N_29672);
and UO_823 (O_823,N_29845,N_29123);
nand UO_824 (O_824,N_29455,N_29863);
xnor UO_825 (O_825,N_29086,N_29512);
nor UO_826 (O_826,N_29192,N_29199);
xnor UO_827 (O_827,N_29359,N_29026);
and UO_828 (O_828,N_29807,N_29164);
and UO_829 (O_829,N_29777,N_29197);
and UO_830 (O_830,N_29295,N_29438);
and UO_831 (O_831,N_29117,N_29758);
xnor UO_832 (O_832,N_29604,N_29802);
nand UO_833 (O_833,N_29375,N_29867);
xor UO_834 (O_834,N_29758,N_29650);
nor UO_835 (O_835,N_29321,N_29333);
and UO_836 (O_836,N_29222,N_29784);
xor UO_837 (O_837,N_29049,N_29911);
nand UO_838 (O_838,N_29943,N_29440);
xnor UO_839 (O_839,N_29185,N_29495);
xnor UO_840 (O_840,N_29558,N_29098);
nor UO_841 (O_841,N_29345,N_29729);
nor UO_842 (O_842,N_29011,N_29017);
nand UO_843 (O_843,N_29522,N_29764);
xor UO_844 (O_844,N_29963,N_29258);
xnor UO_845 (O_845,N_29435,N_29634);
xnor UO_846 (O_846,N_29426,N_29037);
and UO_847 (O_847,N_29736,N_29046);
nor UO_848 (O_848,N_29403,N_29626);
nor UO_849 (O_849,N_29910,N_29258);
or UO_850 (O_850,N_29965,N_29294);
nor UO_851 (O_851,N_29073,N_29853);
nor UO_852 (O_852,N_29957,N_29579);
and UO_853 (O_853,N_29794,N_29727);
xor UO_854 (O_854,N_29914,N_29046);
and UO_855 (O_855,N_29358,N_29228);
and UO_856 (O_856,N_29578,N_29154);
xor UO_857 (O_857,N_29533,N_29128);
nand UO_858 (O_858,N_29228,N_29018);
nand UO_859 (O_859,N_29557,N_29262);
or UO_860 (O_860,N_29540,N_29670);
xnor UO_861 (O_861,N_29836,N_29073);
nor UO_862 (O_862,N_29168,N_29617);
nand UO_863 (O_863,N_29828,N_29903);
nor UO_864 (O_864,N_29024,N_29839);
or UO_865 (O_865,N_29720,N_29544);
or UO_866 (O_866,N_29821,N_29109);
nand UO_867 (O_867,N_29582,N_29067);
nor UO_868 (O_868,N_29148,N_29488);
or UO_869 (O_869,N_29939,N_29202);
nand UO_870 (O_870,N_29099,N_29452);
nand UO_871 (O_871,N_29823,N_29729);
nor UO_872 (O_872,N_29140,N_29361);
nand UO_873 (O_873,N_29665,N_29256);
and UO_874 (O_874,N_29133,N_29937);
and UO_875 (O_875,N_29083,N_29997);
nand UO_876 (O_876,N_29663,N_29943);
nor UO_877 (O_877,N_29339,N_29885);
and UO_878 (O_878,N_29326,N_29626);
or UO_879 (O_879,N_29868,N_29451);
and UO_880 (O_880,N_29935,N_29987);
xnor UO_881 (O_881,N_29746,N_29312);
nor UO_882 (O_882,N_29423,N_29582);
or UO_883 (O_883,N_29872,N_29276);
or UO_884 (O_884,N_29802,N_29989);
or UO_885 (O_885,N_29028,N_29365);
or UO_886 (O_886,N_29297,N_29730);
or UO_887 (O_887,N_29397,N_29909);
nor UO_888 (O_888,N_29169,N_29685);
nor UO_889 (O_889,N_29342,N_29821);
or UO_890 (O_890,N_29338,N_29900);
nor UO_891 (O_891,N_29130,N_29433);
and UO_892 (O_892,N_29994,N_29458);
xor UO_893 (O_893,N_29231,N_29985);
or UO_894 (O_894,N_29009,N_29906);
xnor UO_895 (O_895,N_29825,N_29073);
xor UO_896 (O_896,N_29747,N_29828);
xor UO_897 (O_897,N_29454,N_29813);
xnor UO_898 (O_898,N_29089,N_29629);
or UO_899 (O_899,N_29080,N_29104);
or UO_900 (O_900,N_29832,N_29691);
or UO_901 (O_901,N_29018,N_29346);
or UO_902 (O_902,N_29469,N_29876);
or UO_903 (O_903,N_29775,N_29737);
xor UO_904 (O_904,N_29948,N_29481);
xor UO_905 (O_905,N_29442,N_29382);
or UO_906 (O_906,N_29165,N_29490);
or UO_907 (O_907,N_29365,N_29730);
xnor UO_908 (O_908,N_29804,N_29437);
nor UO_909 (O_909,N_29567,N_29748);
or UO_910 (O_910,N_29665,N_29113);
and UO_911 (O_911,N_29916,N_29543);
and UO_912 (O_912,N_29830,N_29449);
nor UO_913 (O_913,N_29971,N_29917);
and UO_914 (O_914,N_29176,N_29348);
nor UO_915 (O_915,N_29352,N_29024);
nand UO_916 (O_916,N_29480,N_29414);
and UO_917 (O_917,N_29410,N_29995);
xnor UO_918 (O_918,N_29921,N_29558);
nor UO_919 (O_919,N_29186,N_29568);
xnor UO_920 (O_920,N_29366,N_29874);
or UO_921 (O_921,N_29661,N_29452);
or UO_922 (O_922,N_29444,N_29842);
and UO_923 (O_923,N_29980,N_29235);
or UO_924 (O_924,N_29188,N_29542);
nand UO_925 (O_925,N_29304,N_29496);
nor UO_926 (O_926,N_29533,N_29613);
and UO_927 (O_927,N_29815,N_29391);
nor UO_928 (O_928,N_29126,N_29007);
nand UO_929 (O_929,N_29953,N_29795);
or UO_930 (O_930,N_29344,N_29437);
and UO_931 (O_931,N_29528,N_29221);
xor UO_932 (O_932,N_29496,N_29720);
or UO_933 (O_933,N_29014,N_29253);
or UO_934 (O_934,N_29582,N_29994);
nand UO_935 (O_935,N_29962,N_29849);
nand UO_936 (O_936,N_29743,N_29176);
or UO_937 (O_937,N_29615,N_29686);
nand UO_938 (O_938,N_29585,N_29946);
and UO_939 (O_939,N_29642,N_29557);
nand UO_940 (O_940,N_29958,N_29573);
xnor UO_941 (O_941,N_29592,N_29369);
and UO_942 (O_942,N_29595,N_29941);
nor UO_943 (O_943,N_29622,N_29819);
or UO_944 (O_944,N_29983,N_29134);
or UO_945 (O_945,N_29908,N_29688);
or UO_946 (O_946,N_29808,N_29739);
nor UO_947 (O_947,N_29833,N_29858);
and UO_948 (O_948,N_29817,N_29290);
xor UO_949 (O_949,N_29357,N_29852);
nor UO_950 (O_950,N_29834,N_29820);
xor UO_951 (O_951,N_29530,N_29474);
nand UO_952 (O_952,N_29197,N_29916);
and UO_953 (O_953,N_29110,N_29750);
nand UO_954 (O_954,N_29931,N_29227);
and UO_955 (O_955,N_29097,N_29934);
nand UO_956 (O_956,N_29157,N_29126);
xor UO_957 (O_957,N_29638,N_29804);
nand UO_958 (O_958,N_29645,N_29886);
nor UO_959 (O_959,N_29280,N_29145);
nor UO_960 (O_960,N_29494,N_29637);
nand UO_961 (O_961,N_29466,N_29971);
nor UO_962 (O_962,N_29857,N_29097);
nand UO_963 (O_963,N_29572,N_29551);
xnor UO_964 (O_964,N_29138,N_29761);
xnor UO_965 (O_965,N_29351,N_29438);
and UO_966 (O_966,N_29989,N_29743);
nand UO_967 (O_967,N_29716,N_29536);
and UO_968 (O_968,N_29931,N_29834);
and UO_969 (O_969,N_29907,N_29318);
nand UO_970 (O_970,N_29684,N_29533);
xor UO_971 (O_971,N_29587,N_29382);
or UO_972 (O_972,N_29667,N_29900);
nand UO_973 (O_973,N_29451,N_29376);
nor UO_974 (O_974,N_29082,N_29549);
xnor UO_975 (O_975,N_29319,N_29545);
xnor UO_976 (O_976,N_29928,N_29078);
nand UO_977 (O_977,N_29141,N_29137);
and UO_978 (O_978,N_29152,N_29318);
xnor UO_979 (O_979,N_29515,N_29039);
and UO_980 (O_980,N_29572,N_29888);
xor UO_981 (O_981,N_29114,N_29869);
nand UO_982 (O_982,N_29373,N_29708);
nor UO_983 (O_983,N_29112,N_29831);
or UO_984 (O_984,N_29103,N_29511);
and UO_985 (O_985,N_29160,N_29307);
xor UO_986 (O_986,N_29328,N_29746);
or UO_987 (O_987,N_29541,N_29871);
or UO_988 (O_988,N_29925,N_29244);
and UO_989 (O_989,N_29652,N_29203);
and UO_990 (O_990,N_29352,N_29899);
nor UO_991 (O_991,N_29047,N_29925);
and UO_992 (O_992,N_29209,N_29277);
or UO_993 (O_993,N_29293,N_29113);
nor UO_994 (O_994,N_29635,N_29739);
nand UO_995 (O_995,N_29914,N_29952);
xnor UO_996 (O_996,N_29367,N_29088);
nor UO_997 (O_997,N_29759,N_29486);
nand UO_998 (O_998,N_29157,N_29134);
nor UO_999 (O_999,N_29094,N_29370);
xnor UO_1000 (O_1000,N_29912,N_29555);
xor UO_1001 (O_1001,N_29860,N_29957);
nand UO_1002 (O_1002,N_29415,N_29849);
or UO_1003 (O_1003,N_29129,N_29733);
nand UO_1004 (O_1004,N_29752,N_29663);
nor UO_1005 (O_1005,N_29928,N_29404);
nor UO_1006 (O_1006,N_29512,N_29618);
or UO_1007 (O_1007,N_29904,N_29125);
and UO_1008 (O_1008,N_29338,N_29721);
and UO_1009 (O_1009,N_29567,N_29161);
nor UO_1010 (O_1010,N_29342,N_29937);
nor UO_1011 (O_1011,N_29762,N_29788);
nand UO_1012 (O_1012,N_29226,N_29571);
nor UO_1013 (O_1013,N_29261,N_29616);
nor UO_1014 (O_1014,N_29280,N_29431);
nand UO_1015 (O_1015,N_29078,N_29381);
and UO_1016 (O_1016,N_29276,N_29940);
and UO_1017 (O_1017,N_29666,N_29307);
and UO_1018 (O_1018,N_29912,N_29691);
xor UO_1019 (O_1019,N_29842,N_29106);
nand UO_1020 (O_1020,N_29426,N_29384);
nand UO_1021 (O_1021,N_29089,N_29011);
or UO_1022 (O_1022,N_29296,N_29984);
nor UO_1023 (O_1023,N_29161,N_29528);
xor UO_1024 (O_1024,N_29668,N_29991);
and UO_1025 (O_1025,N_29394,N_29119);
and UO_1026 (O_1026,N_29114,N_29307);
nand UO_1027 (O_1027,N_29571,N_29479);
or UO_1028 (O_1028,N_29039,N_29638);
or UO_1029 (O_1029,N_29224,N_29627);
nor UO_1030 (O_1030,N_29001,N_29715);
or UO_1031 (O_1031,N_29865,N_29066);
nand UO_1032 (O_1032,N_29009,N_29907);
xor UO_1033 (O_1033,N_29040,N_29674);
nand UO_1034 (O_1034,N_29223,N_29782);
xnor UO_1035 (O_1035,N_29009,N_29618);
nor UO_1036 (O_1036,N_29197,N_29772);
or UO_1037 (O_1037,N_29354,N_29342);
or UO_1038 (O_1038,N_29177,N_29992);
nor UO_1039 (O_1039,N_29596,N_29260);
or UO_1040 (O_1040,N_29351,N_29896);
xor UO_1041 (O_1041,N_29691,N_29715);
and UO_1042 (O_1042,N_29723,N_29508);
xnor UO_1043 (O_1043,N_29614,N_29208);
nand UO_1044 (O_1044,N_29061,N_29918);
xor UO_1045 (O_1045,N_29226,N_29500);
nand UO_1046 (O_1046,N_29779,N_29161);
and UO_1047 (O_1047,N_29990,N_29159);
nor UO_1048 (O_1048,N_29877,N_29253);
xor UO_1049 (O_1049,N_29317,N_29544);
or UO_1050 (O_1050,N_29246,N_29841);
and UO_1051 (O_1051,N_29554,N_29993);
and UO_1052 (O_1052,N_29615,N_29191);
nor UO_1053 (O_1053,N_29009,N_29330);
or UO_1054 (O_1054,N_29448,N_29194);
and UO_1055 (O_1055,N_29956,N_29923);
xor UO_1056 (O_1056,N_29694,N_29586);
or UO_1057 (O_1057,N_29610,N_29629);
nor UO_1058 (O_1058,N_29337,N_29717);
nor UO_1059 (O_1059,N_29145,N_29756);
and UO_1060 (O_1060,N_29955,N_29989);
nor UO_1061 (O_1061,N_29480,N_29460);
or UO_1062 (O_1062,N_29371,N_29258);
nand UO_1063 (O_1063,N_29646,N_29309);
nand UO_1064 (O_1064,N_29682,N_29216);
xnor UO_1065 (O_1065,N_29635,N_29567);
nor UO_1066 (O_1066,N_29407,N_29030);
xnor UO_1067 (O_1067,N_29269,N_29768);
and UO_1068 (O_1068,N_29190,N_29735);
or UO_1069 (O_1069,N_29676,N_29234);
xor UO_1070 (O_1070,N_29248,N_29988);
and UO_1071 (O_1071,N_29455,N_29964);
and UO_1072 (O_1072,N_29818,N_29986);
nand UO_1073 (O_1073,N_29657,N_29548);
xor UO_1074 (O_1074,N_29851,N_29190);
xor UO_1075 (O_1075,N_29042,N_29081);
or UO_1076 (O_1076,N_29515,N_29913);
and UO_1077 (O_1077,N_29284,N_29911);
nor UO_1078 (O_1078,N_29447,N_29394);
or UO_1079 (O_1079,N_29921,N_29997);
nor UO_1080 (O_1080,N_29702,N_29343);
or UO_1081 (O_1081,N_29143,N_29690);
xor UO_1082 (O_1082,N_29230,N_29317);
xnor UO_1083 (O_1083,N_29964,N_29167);
and UO_1084 (O_1084,N_29369,N_29674);
nand UO_1085 (O_1085,N_29586,N_29927);
and UO_1086 (O_1086,N_29787,N_29748);
or UO_1087 (O_1087,N_29234,N_29303);
nand UO_1088 (O_1088,N_29284,N_29546);
nand UO_1089 (O_1089,N_29625,N_29016);
and UO_1090 (O_1090,N_29949,N_29257);
and UO_1091 (O_1091,N_29387,N_29563);
or UO_1092 (O_1092,N_29807,N_29336);
and UO_1093 (O_1093,N_29250,N_29046);
or UO_1094 (O_1094,N_29002,N_29733);
xnor UO_1095 (O_1095,N_29677,N_29687);
xnor UO_1096 (O_1096,N_29817,N_29520);
or UO_1097 (O_1097,N_29828,N_29444);
nand UO_1098 (O_1098,N_29652,N_29543);
and UO_1099 (O_1099,N_29176,N_29697);
xor UO_1100 (O_1100,N_29158,N_29842);
nor UO_1101 (O_1101,N_29083,N_29099);
nor UO_1102 (O_1102,N_29679,N_29217);
nor UO_1103 (O_1103,N_29395,N_29406);
or UO_1104 (O_1104,N_29230,N_29490);
nand UO_1105 (O_1105,N_29276,N_29383);
nand UO_1106 (O_1106,N_29873,N_29890);
nand UO_1107 (O_1107,N_29075,N_29939);
xor UO_1108 (O_1108,N_29316,N_29107);
nand UO_1109 (O_1109,N_29235,N_29091);
and UO_1110 (O_1110,N_29418,N_29279);
and UO_1111 (O_1111,N_29795,N_29945);
nor UO_1112 (O_1112,N_29929,N_29699);
xor UO_1113 (O_1113,N_29997,N_29924);
and UO_1114 (O_1114,N_29223,N_29540);
or UO_1115 (O_1115,N_29921,N_29459);
and UO_1116 (O_1116,N_29388,N_29594);
nor UO_1117 (O_1117,N_29208,N_29122);
or UO_1118 (O_1118,N_29712,N_29008);
or UO_1119 (O_1119,N_29641,N_29294);
nand UO_1120 (O_1120,N_29207,N_29327);
xnor UO_1121 (O_1121,N_29342,N_29223);
nor UO_1122 (O_1122,N_29747,N_29736);
or UO_1123 (O_1123,N_29060,N_29304);
nand UO_1124 (O_1124,N_29669,N_29572);
nor UO_1125 (O_1125,N_29463,N_29144);
or UO_1126 (O_1126,N_29433,N_29321);
nor UO_1127 (O_1127,N_29127,N_29752);
xnor UO_1128 (O_1128,N_29014,N_29695);
nand UO_1129 (O_1129,N_29872,N_29012);
and UO_1130 (O_1130,N_29080,N_29513);
nand UO_1131 (O_1131,N_29148,N_29726);
and UO_1132 (O_1132,N_29758,N_29241);
and UO_1133 (O_1133,N_29433,N_29225);
or UO_1134 (O_1134,N_29423,N_29344);
nor UO_1135 (O_1135,N_29068,N_29655);
or UO_1136 (O_1136,N_29687,N_29323);
xor UO_1137 (O_1137,N_29219,N_29576);
nor UO_1138 (O_1138,N_29059,N_29337);
and UO_1139 (O_1139,N_29673,N_29336);
xnor UO_1140 (O_1140,N_29293,N_29500);
nor UO_1141 (O_1141,N_29656,N_29149);
nand UO_1142 (O_1142,N_29112,N_29930);
nor UO_1143 (O_1143,N_29354,N_29421);
and UO_1144 (O_1144,N_29917,N_29291);
and UO_1145 (O_1145,N_29600,N_29628);
xor UO_1146 (O_1146,N_29622,N_29534);
nor UO_1147 (O_1147,N_29572,N_29117);
and UO_1148 (O_1148,N_29569,N_29128);
nor UO_1149 (O_1149,N_29693,N_29710);
or UO_1150 (O_1150,N_29965,N_29345);
and UO_1151 (O_1151,N_29372,N_29907);
nand UO_1152 (O_1152,N_29102,N_29141);
nand UO_1153 (O_1153,N_29801,N_29867);
nand UO_1154 (O_1154,N_29530,N_29914);
or UO_1155 (O_1155,N_29250,N_29330);
xnor UO_1156 (O_1156,N_29492,N_29889);
nor UO_1157 (O_1157,N_29522,N_29691);
nand UO_1158 (O_1158,N_29523,N_29603);
nand UO_1159 (O_1159,N_29806,N_29793);
or UO_1160 (O_1160,N_29689,N_29081);
or UO_1161 (O_1161,N_29824,N_29375);
and UO_1162 (O_1162,N_29515,N_29074);
nor UO_1163 (O_1163,N_29361,N_29713);
and UO_1164 (O_1164,N_29201,N_29801);
xor UO_1165 (O_1165,N_29668,N_29461);
nor UO_1166 (O_1166,N_29758,N_29251);
nor UO_1167 (O_1167,N_29040,N_29861);
nor UO_1168 (O_1168,N_29009,N_29072);
and UO_1169 (O_1169,N_29585,N_29127);
and UO_1170 (O_1170,N_29893,N_29046);
nand UO_1171 (O_1171,N_29486,N_29629);
xnor UO_1172 (O_1172,N_29128,N_29443);
xnor UO_1173 (O_1173,N_29463,N_29568);
nand UO_1174 (O_1174,N_29039,N_29150);
nand UO_1175 (O_1175,N_29112,N_29372);
xor UO_1176 (O_1176,N_29495,N_29976);
xor UO_1177 (O_1177,N_29478,N_29590);
and UO_1178 (O_1178,N_29437,N_29352);
and UO_1179 (O_1179,N_29293,N_29552);
nand UO_1180 (O_1180,N_29959,N_29021);
xor UO_1181 (O_1181,N_29374,N_29304);
xor UO_1182 (O_1182,N_29645,N_29609);
nor UO_1183 (O_1183,N_29455,N_29543);
or UO_1184 (O_1184,N_29101,N_29996);
nor UO_1185 (O_1185,N_29671,N_29789);
or UO_1186 (O_1186,N_29162,N_29338);
nand UO_1187 (O_1187,N_29032,N_29972);
nor UO_1188 (O_1188,N_29777,N_29521);
nand UO_1189 (O_1189,N_29710,N_29546);
or UO_1190 (O_1190,N_29426,N_29409);
and UO_1191 (O_1191,N_29435,N_29761);
or UO_1192 (O_1192,N_29395,N_29731);
nor UO_1193 (O_1193,N_29505,N_29946);
nor UO_1194 (O_1194,N_29028,N_29310);
xnor UO_1195 (O_1195,N_29282,N_29277);
nor UO_1196 (O_1196,N_29982,N_29040);
and UO_1197 (O_1197,N_29462,N_29944);
nand UO_1198 (O_1198,N_29511,N_29091);
and UO_1199 (O_1199,N_29551,N_29751);
nor UO_1200 (O_1200,N_29529,N_29060);
xnor UO_1201 (O_1201,N_29374,N_29765);
nor UO_1202 (O_1202,N_29330,N_29575);
nand UO_1203 (O_1203,N_29816,N_29432);
or UO_1204 (O_1204,N_29280,N_29251);
nand UO_1205 (O_1205,N_29379,N_29750);
nand UO_1206 (O_1206,N_29570,N_29277);
nor UO_1207 (O_1207,N_29901,N_29881);
or UO_1208 (O_1208,N_29704,N_29035);
nor UO_1209 (O_1209,N_29744,N_29902);
or UO_1210 (O_1210,N_29757,N_29926);
nor UO_1211 (O_1211,N_29108,N_29340);
or UO_1212 (O_1212,N_29047,N_29324);
xnor UO_1213 (O_1213,N_29888,N_29641);
nor UO_1214 (O_1214,N_29629,N_29158);
or UO_1215 (O_1215,N_29749,N_29906);
and UO_1216 (O_1216,N_29950,N_29580);
and UO_1217 (O_1217,N_29180,N_29498);
and UO_1218 (O_1218,N_29094,N_29952);
and UO_1219 (O_1219,N_29264,N_29927);
xnor UO_1220 (O_1220,N_29398,N_29182);
xnor UO_1221 (O_1221,N_29446,N_29917);
or UO_1222 (O_1222,N_29835,N_29801);
and UO_1223 (O_1223,N_29677,N_29490);
nor UO_1224 (O_1224,N_29628,N_29374);
nor UO_1225 (O_1225,N_29535,N_29802);
nand UO_1226 (O_1226,N_29271,N_29296);
or UO_1227 (O_1227,N_29988,N_29883);
xor UO_1228 (O_1228,N_29216,N_29189);
nand UO_1229 (O_1229,N_29819,N_29394);
and UO_1230 (O_1230,N_29445,N_29878);
nor UO_1231 (O_1231,N_29498,N_29558);
or UO_1232 (O_1232,N_29155,N_29057);
xnor UO_1233 (O_1233,N_29089,N_29843);
nand UO_1234 (O_1234,N_29350,N_29989);
xor UO_1235 (O_1235,N_29168,N_29455);
nor UO_1236 (O_1236,N_29042,N_29517);
xnor UO_1237 (O_1237,N_29425,N_29640);
or UO_1238 (O_1238,N_29139,N_29098);
or UO_1239 (O_1239,N_29420,N_29899);
nand UO_1240 (O_1240,N_29479,N_29399);
nand UO_1241 (O_1241,N_29700,N_29216);
nand UO_1242 (O_1242,N_29354,N_29165);
nor UO_1243 (O_1243,N_29197,N_29551);
nand UO_1244 (O_1244,N_29300,N_29733);
xnor UO_1245 (O_1245,N_29941,N_29739);
xnor UO_1246 (O_1246,N_29176,N_29568);
nand UO_1247 (O_1247,N_29386,N_29140);
nor UO_1248 (O_1248,N_29388,N_29278);
nor UO_1249 (O_1249,N_29330,N_29290);
xor UO_1250 (O_1250,N_29730,N_29515);
or UO_1251 (O_1251,N_29380,N_29170);
nand UO_1252 (O_1252,N_29072,N_29635);
or UO_1253 (O_1253,N_29331,N_29329);
nand UO_1254 (O_1254,N_29810,N_29752);
nor UO_1255 (O_1255,N_29237,N_29547);
and UO_1256 (O_1256,N_29717,N_29786);
or UO_1257 (O_1257,N_29094,N_29618);
and UO_1258 (O_1258,N_29212,N_29153);
or UO_1259 (O_1259,N_29701,N_29544);
or UO_1260 (O_1260,N_29059,N_29278);
nand UO_1261 (O_1261,N_29878,N_29417);
nand UO_1262 (O_1262,N_29565,N_29274);
nor UO_1263 (O_1263,N_29527,N_29990);
nand UO_1264 (O_1264,N_29302,N_29234);
nor UO_1265 (O_1265,N_29339,N_29573);
xnor UO_1266 (O_1266,N_29892,N_29522);
nand UO_1267 (O_1267,N_29576,N_29176);
nand UO_1268 (O_1268,N_29812,N_29597);
or UO_1269 (O_1269,N_29398,N_29903);
xor UO_1270 (O_1270,N_29325,N_29332);
and UO_1271 (O_1271,N_29433,N_29212);
nor UO_1272 (O_1272,N_29153,N_29340);
nor UO_1273 (O_1273,N_29595,N_29493);
nor UO_1274 (O_1274,N_29842,N_29503);
nor UO_1275 (O_1275,N_29965,N_29138);
xnor UO_1276 (O_1276,N_29110,N_29941);
or UO_1277 (O_1277,N_29747,N_29259);
nand UO_1278 (O_1278,N_29896,N_29177);
or UO_1279 (O_1279,N_29240,N_29660);
nand UO_1280 (O_1280,N_29332,N_29893);
xnor UO_1281 (O_1281,N_29308,N_29342);
xnor UO_1282 (O_1282,N_29654,N_29621);
and UO_1283 (O_1283,N_29333,N_29563);
nand UO_1284 (O_1284,N_29671,N_29665);
nand UO_1285 (O_1285,N_29503,N_29932);
or UO_1286 (O_1286,N_29300,N_29677);
and UO_1287 (O_1287,N_29490,N_29926);
nand UO_1288 (O_1288,N_29674,N_29141);
nand UO_1289 (O_1289,N_29053,N_29922);
or UO_1290 (O_1290,N_29339,N_29157);
xor UO_1291 (O_1291,N_29144,N_29827);
xnor UO_1292 (O_1292,N_29569,N_29553);
nand UO_1293 (O_1293,N_29861,N_29841);
or UO_1294 (O_1294,N_29318,N_29776);
and UO_1295 (O_1295,N_29438,N_29370);
nor UO_1296 (O_1296,N_29523,N_29820);
and UO_1297 (O_1297,N_29008,N_29696);
nor UO_1298 (O_1298,N_29759,N_29700);
nor UO_1299 (O_1299,N_29792,N_29133);
xor UO_1300 (O_1300,N_29713,N_29271);
xnor UO_1301 (O_1301,N_29225,N_29845);
nand UO_1302 (O_1302,N_29502,N_29053);
and UO_1303 (O_1303,N_29260,N_29273);
nor UO_1304 (O_1304,N_29135,N_29393);
and UO_1305 (O_1305,N_29449,N_29658);
nor UO_1306 (O_1306,N_29575,N_29367);
xor UO_1307 (O_1307,N_29073,N_29743);
xor UO_1308 (O_1308,N_29993,N_29930);
nor UO_1309 (O_1309,N_29627,N_29314);
nand UO_1310 (O_1310,N_29231,N_29926);
or UO_1311 (O_1311,N_29601,N_29941);
nand UO_1312 (O_1312,N_29305,N_29308);
nor UO_1313 (O_1313,N_29301,N_29881);
or UO_1314 (O_1314,N_29309,N_29598);
or UO_1315 (O_1315,N_29098,N_29727);
and UO_1316 (O_1316,N_29794,N_29665);
nor UO_1317 (O_1317,N_29503,N_29926);
xnor UO_1318 (O_1318,N_29406,N_29483);
nor UO_1319 (O_1319,N_29850,N_29077);
nor UO_1320 (O_1320,N_29452,N_29421);
nand UO_1321 (O_1321,N_29203,N_29490);
xnor UO_1322 (O_1322,N_29440,N_29178);
xnor UO_1323 (O_1323,N_29692,N_29960);
or UO_1324 (O_1324,N_29134,N_29467);
xor UO_1325 (O_1325,N_29083,N_29703);
xnor UO_1326 (O_1326,N_29694,N_29214);
nor UO_1327 (O_1327,N_29308,N_29835);
nor UO_1328 (O_1328,N_29212,N_29331);
xnor UO_1329 (O_1329,N_29686,N_29810);
nor UO_1330 (O_1330,N_29499,N_29254);
nor UO_1331 (O_1331,N_29690,N_29394);
and UO_1332 (O_1332,N_29886,N_29371);
nor UO_1333 (O_1333,N_29298,N_29104);
or UO_1334 (O_1334,N_29069,N_29422);
or UO_1335 (O_1335,N_29007,N_29836);
xnor UO_1336 (O_1336,N_29033,N_29644);
xnor UO_1337 (O_1337,N_29817,N_29757);
and UO_1338 (O_1338,N_29058,N_29599);
and UO_1339 (O_1339,N_29436,N_29458);
or UO_1340 (O_1340,N_29904,N_29188);
nand UO_1341 (O_1341,N_29894,N_29576);
and UO_1342 (O_1342,N_29079,N_29132);
xor UO_1343 (O_1343,N_29612,N_29372);
or UO_1344 (O_1344,N_29239,N_29902);
or UO_1345 (O_1345,N_29588,N_29552);
or UO_1346 (O_1346,N_29954,N_29840);
or UO_1347 (O_1347,N_29214,N_29060);
nor UO_1348 (O_1348,N_29572,N_29023);
xnor UO_1349 (O_1349,N_29623,N_29650);
and UO_1350 (O_1350,N_29105,N_29351);
xnor UO_1351 (O_1351,N_29050,N_29286);
or UO_1352 (O_1352,N_29394,N_29859);
or UO_1353 (O_1353,N_29862,N_29102);
nor UO_1354 (O_1354,N_29391,N_29709);
xor UO_1355 (O_1355,N_29973,N_29632);
xor UO_1356 (O_1356,N_29032,N_29880);
nand UO_1357 (O_1357,N_29066,N_29712);
and UO_1358 (O_1358,N_29748,N_29263);
nor UO_1359 (O_1359,N_29377,N_29853);
xor UO_1360 (O_1360,N_29743,N_29214);
nor UO_1361 (O_1361,N_29620,N_29735);
nor UO_1362 (O_1362,N_29668,N_29545);
nor UO_1363 (O_1363,N_29083,N_29945);
nor UO_1364 (O_1364,N_29760,N_29420);
nor UO_1365 (O_1365,N_29255,N_29999);
or UO_1366 (O_1366,N_29188,N_29000);
nor UO_1367 (O_1367,N_29402,N_29480);
nor UO_1368 (O_1368,N_29593,N_29476);
or UO_1369 (O_1369,N_29726,N_29874);
nor UO_1370 (O_1370,N_29830,N_29961);
or UO_1371 (O_1371,N_29144,N_29120);
nor UO_1372 (O_1372,N_29392,N_29953);
and UO_1373 (O_1373,N_29773,N_29700);
nand UO_1374 (O_1374,N_29762,N_29893);
nand UO_1375 (O_1375,N_29296,N_29210);
xnor UO_1376 (O_1376,N_29800,N_29580);
nand UO_1377 (O_1377,N_29928,N_29833);
nand UO_1378 (O_1378,N_29354,N_29142);
or UO_1379 (O_1379,N_29963,N_29191);
and UO_1380 (O_1380,N_29189,N_29554);
nor UO_1381 (O_1381,N_29191,N_29272);
nor UO_1382 (O_1382,N_29490,N_29955);
or UO_1383 (O_1383,N_29677,N_29247);
nor UO_1384 (O_1384,N_29129,N_29913);
and UO_1385 (O_1385,N_29677,N_29648);
xor UO_1386 (O_1386,N_29243,N_29155);
xnor UO_1387 (O_1387,N_29431,N_29001);
nor UO_1388 (O_1388,N_29711,N_29822);
xor UO_1389 (O_1389,N_29827,N_29696);
nand UO_1390 (O_1390,N_29657,N_29344);
xor UO_1391 (O_1391,N_29063,N_29290);
nor UO_1392 (O_1392,N_29133,N_29801);
or UO_1393 (O_1393,N_29789,N_29788);
xnor UO_1394 (O_1394,N_29326,N_29989);
nor UO_1395 (O_1395,N_29880,N_29326);
nand UO_1396 (O_1396,N_29089,N_29053);
or UO_1397 (O_1397,N_29333,N_29485);
nor UO_1398 (O_1398,N_29562,N_29108);
xor UO_1399 (O_1399,N_29597,N_29466);
nand UO_1400 (O_1400,N_29517,N_29716);
nor UO_1401 (O_1401,N_29640,N_29809);
xor UO_1402 (O_1402,N_29482,N_29698);
and UO_1403 (O_1403,N_29745,N_29292);
and UO_1404 (O_1404,N_29058,N_29432);
and UO_1405 (O_1405,N_29081,N_29831);
xnor UO_1406 (O_1406,N_29341,N_29926);
nand UO_1407 (O_1407,N_29849,N_29458);
xor UO_1408 (O_1408,N_29780,N_29855);
nor UO_1409 (O_1409,N_29167,N_29968);
nand UO_1410 (O_1410,N_29417,N_29429);
nor UO_1411 (O_1411,N_29660,N_29971);
nand UO_1412 (O_1412,N_29436,N_29530);
or UO_1413 (O_1413,N_29510,N_29527);
xor UO_1414 (O_1414,N_29710,N_29525);
and UO_1415 (O_1415,N_29312,N_29607);
and UO_1416 (O_1416,N_29558,N_29648);
nor UO_1417 (O_1417,N_29805,N_29812);
and UO_1418 (O_1418,N_29912,N_29361);
xnor UO_1419 (O_1419,N_29555,N_29837);
nand UO_1420 (O_1420,N_29352,N_29756);
nand UO_1421 (O_1421,N_29672,N_29080);
xor UO_1422 (O_1422,N_29989,N_29226);
nor UO_1423 (O_1423,N_29423,N_29339);
xnor UO_1424 (O_1424,N_29003,N_29831);
xnor UO_1425 (O_1425,N_29557,N_29633);
and UO_1426 (O_1426,N_29236,N_29021);
xnor UO_1427 (O_1427,N_29086,N_29832);
or UO_1428 (O_1428,N_29561,N_29989);
nand UO_1429 (O_1429,N_29187,N_29515);
and UO_1430 (O_1430,N_29137,N_29011);
nor UO_1431 (O_1431,N_29871,N_29811);
nand UO_1432 (O_1432,N_29749,N_29546);
nor UO_1433 (O_1433,N_29001,N_29292);
nand UO_1434 (O_1434,N_29142,N_29140);
and UO_1435 (O_1435,N_29541,N_29092);
xnor UO_1436 (O_1436,N_29054,N_29611);
xnor UO_1437 (O_1437,N_29259,N_29937);
nand UO_1438 (O_1438,N_29276,N_29611);
nor UO_1439 (O_1439,N_29563,N_29730);
or UO_1440 (O_1440,N_29752,N_29091);
nor UO_1441 (O_1441,N_29430,N_29493);
or UO_1442 (O_1442,N_29435,N_29304);
and UO_1443 (O_1443,N_29115,N_29477);
xnor UO_1444 (O_1444,N_29253,N_29944);
and UO_1445 (O_1445,N_29891,N_29116);
nand UO_1446 (O_1446,N_29732,N_29683);
nor UO_1447 (O_1447,N_29288,N_29181);
xnor UO_1448 (O_1448,N_29553,N_29726);
nor UO_1449 (O_1449,N_29265,N_29676);
nor UO_1450 (O_1450,N_29999,N_29015);
and UO_1451 (O_1451,N_29689,N_29800);
nand UO_1452 (O_1452,N_29641,N_29514);
xor UO_1453 (O_1453,N_29248,N_29593);
and UO_1454 (O_1454,N_29198,N_29108);
or UO_1455 (O_1455,N_29483,N_29368);
xor UO_1456 (O_1456,N_29458,N_29242);
xor UO_1457 (O_1457,N_29735,N_29971);
xor UO_1458 (O_1458,N_29932,N_29799);
nor UO_1459 (O_1459,N_29505,N_29220);
and UO_1460 (O_1460,N_29093,N_29995);
nand UO_1461 (O_1461,N_29152,N_29749);
and UO_1462 (O_1462,N_29897,N_29796);
nand UO_1463 (O_1463,N_29835,N_29404);
nand UO_1464 (O_1464,N_29591,N_29492);
and UO_1465 (O_1465,N_29774,N_29012);
and UO_1466 (O_1466,N_29219,N_29779);
and UO_1467 (O_1467,N_29738,N_29924);
and UO_1468 (O_1468,N_29375,N_29724);
or UO_1469 (O_1469,N_29044,N_29721);
xor UO_1470 (O_1470,N_29887,N_29451);
xor UO_1471 (O_1471,N_29888,N_29129);
and UO_1472 (O_1472,N_29537,N_29828);
and UO_1473 (O_1473,N_29620,N_29318);
nor UO_1474 (O_1474,N_29418,N_29174);
xnor UO_1475 (O_1475,N_29632,N_29415);
nor UO_1476 (O_1476,N_29232,N_29428);
nor UO_1477 (O_1477,N_29805,N_29368);
nand UO_1478 (O_1478,N_29539,N_29693);
xnor UO_1479 (O_1479,N_29272,N_29250);
and UO_1480 (O_1480,N_29831,N_29923);
nor UO_1481 (O_1481,N_29045,N_29561);
xor UO_1482 (O_1482,N_29495,N_29385);
or UO_1483 (O_1483,N_29434,N_29270);
nor UO_1484 (O_1484,N_29410,N_29235);
and UO_1485 (O_1485,N_29210,N_29405);
or UO_1486 (O_1486,N_29246,N_29541);
or UO_1487 (O_1487,N_29304,N_29648);
or UO_1488 (O_1488,N_29228,N_29651);
and UO_1489 (O_1489,N_29124,N_29827);
nand UO_1490 (O_1490,N_29785,N_29602);
or UO_1491 (O_1491,N_29704,N_29647);
or UO_1492 (O_1492,N_29171,N_29139);
xnor UO_1493 (O_1493,N_29050,N_29168);
or UO_1494 (O_1494,N_29677,N_29791);
nor UO_1495 (O_1495,N_29221,N_29320);
nor UO_1496 (O_1496,N_29252,N_29552);
xor UO_1497 (O_1497,N_29221,N_29165);
and UO_1498 (O_1498,N_29451,N_29731);
or UO_1499 (O_1499,N_29312,N_29422);
and UO_1500 (O_1500,N_29038,N_29662);
or UO_1501 (O_1501,N_29547,N_29157);
and UO_1502 (O_1502,N_29329,N_29568);
or UO_1503 (O_1503,N_29586,N_29511);
or UO_1504 (O_1504,N_29913,N_29562);
nor UO_1505 (O_1505,N_29432,N_29497);
nor UO_1506 (O_1506,N_29444,N_29878);
nand UO_1507 (O_1507,N_29113,N_29769);
nor UO_1508 (O_1508,N_29879,N_29461);
nand UO_1509 (O_1509,N_29708,N_29890);
nor UO_1510 (O_1510,N_29959,N_29194);
and UO_1511 (O_1511,N_29194,N_29215);
and UO_1512 (O_1512,N_29656,N_29321);
nor UO_1513 (O_1513,N_29367,N_29422);
or UO_1514 (O_1514,N_29205,N_29697);
and UO_1515 (O_1515,N_29982,N_29560);
and UO_1516 (O_1516,N_29122,N_29615);
nor UO_1517 (O_1517,N_29427,N_29801);
and UO_1518 (O_1518,N_29194,N_29744);
and UO_1519 (O_1519,N_29002,N_29335);
nor UO_1520 (O_1520,N_29830,N_29330);
nor UO_1521 (O_1521,N_29590,N_29879);
xnor UO_1522 (O_1522,N_29740,N_29789);
and UO_1523 (O_1523,N_29596,N_29121);
xor UO_1524 (O_1524,N_29067,N_29433);
or UO_1525 (O_1525,N_29160,N_29524);
xor UO_1526 (O_1526,N_29765,N_29200);
xor UO_1527 (O_1527,N_29782,N_29292);
or UO_1528 (O_1528,N_29199,N_29282);
xor UO_1529 (O_1529,N_29984,N_29947);
or UO_1530 (O_1530,N_29052,N_29724);
nor UO_1531 (O_1531,N_29799,N_29613);
and UO_1532 (O_1532,N_29027,N_29614);
and UO_1533 (O_1533,N_29043,N_29769);
xor UO_1534 (O_1534,N_29351,N_29047);
xnor UO_1535 (O_1535,N_29467,N_29903);
xnor UO_1536 (O_1536,N_29655,N_29557);
and UO_1537 (O_1537,N_29747,N_29148);
or UO_1538 (O_1538,N_29148,N_29483);
xor UO_1539 (O_1539,N_29733,N_29364);
nor UO_1540 (O_1540,N_29355,N_29829);
nand UO_1541 (O_1541,N_29055,N_29243);
xnor UO_1542 (O_1542,N_29077,N_29553);
xor UO_1543 (O_1543,N_29976,N_29122);
xnor UO_1544 (O_1544,N_29220,N_29173);
and UO_1545 (O_1545,N_29283,N_29562);
or UO_1546 (O_1546,N_29192,N_29497);
nor UO_1547 (O_1547,N_29047,N_29959);
nand UO_1548 (O_1548,N_29634,N_29809);
and UO_1549 (O_1549,N_29798,N_29098);
or UO_1550 (O_1550,N_29462,N_29232);
and UO_1551 (O_1551,N_29774,N_29465);
or UO_1552 (O_1552,N_29795,N_29347);
or UO_1553 (O_1553,N_29123,N_29457);
nor UO_1554 (O_1554,N_29206,N_29711);
and UO_1555 (O_1555,N_29392,N_29571);
nor UO_1556 (O_1556,N_29866,N_29245);
nor UO_1557 (O_1557,N_29554,N_29852);
or UO_1558 (O_1558,N_29212,N_29158);
nor UO_1559 (O_1559,N_29516,N_29385);
xnor UO_1560 (O_1560,N_29760,N_29693);
nor UO_1561 (O_1561,N_29990,N_29454);
nand UO_1562 (O_1562,N_29705,N_29967);
and UO_1563 (O_1563,N_29390,N_29450);
nand UO_1564 (O_1564,N_29579,N_29010);
and UO_1565 (O_1565,N_29723,N_29468);
or UO_1566 (O_1566,N_29879,N_29640);
and UO_1567 (O_1567,N_29367,N_29855);
xor UO_1568 (O_1568,N_29143,N_29079);
or UO_1569 (O_1569,N_29744,N_29718);
xnor UO_1570 (O_1570,N_29512,N_29828);
and UO_1571 (O_1571,N_29473,N_29919);
nand UO_1572 (O_1572,N_29379,N_29378);
or UO_1573 (O_1573,N_29133,N_29010);
and UO_1574 (O_1574,N_29591,N_29775);
nand UO_1575 (O_1575,N_29759,N_29285);
nor UO_1576 (O_1576,N_29767,N_29687);
and UO_1577 (O_1577,N_29669,N_29279);
nor UO_1578 (O_1578,N_29621,N_29085);
and UO_1579 (O_1579,N_29280,N_29451);
and UO_1580 (O_1580,N_29564,N_29461);
nor UO_1581 (O_1581,N_29597,N_29936);
xnor UO_1582 (O_1582,N_29764,N_29310);
nor UO_1583 (O_1583,N_29434,N_29949);
nor UO_1584 (O_1584,N_29961,N_29168);
or UO_1585 (O_1585,N_29985,N_29173);
xnor UO_1586 (O_1586,N_29498,N_29439);
xnor UO_1587 (O_1587,N_29999,N_29638);
nor UO_1588 (O_1588,N_29744,N_29394);
or UO_1589 (O_1589,N_29223,N_29564);
nor UO_1590 (O_1590,N_29340,N_29574);
and UO_1591 (O_1591,N_29365,N_29576);
nor UO_1592 (O_1592,N_29733,N_29794);
nand UO_1593 (O_1593,N_29792,N_29289);
nand UO_1594 (O_1594,N_29051,N_29598);
xnor UO_1595 (O_1595,N_29418,N_29760);
nand UO_1596 (O_1596,N_29553,N_29780);
nor UO_1597 (O_1597,N_29960,N_29775);
or UO_1598 (O_1598,N_29256,N_29238);
nor UO_1599 (O_1599,N_29347,N_29912);
nor UO_1600 (O_1600,N_29762,N_29152);
nor UO_1601 (O_1601,N_29541,N_29234);
nor UO_1602 (O_1602,N_29492,N_29340);
or UO_1603 (O_1603,N_29294,N_29122);
and UO_1604 (O_1604,N_29427,N_29398);
nand UO_1605 (O_1605,N_29350,N_29253);
and UO_1606 (O_1606,N_29418,N_29807);
and UO_1607 (O_1607,N_29142,N_29381);
and UO_1608 (O_1608,N_29282,N_29382);
or UO_1609 (O_1609,N_29854,N_29749);
nand UO_1610 (O_1610,N_29125,N_29661);
or UO_1611 (O_1611,N_29724,N_29669);
xnor UO_1612 (O_1612,N_29116,N_29922);
and UO_1613 (O_1613,N_29743,N_29740);
and UO_1614 (O_1614,N_29141,N_29109);
xnor UO_1615 (O_1615,N_29609,N_29520);
nand UO_1616 (O_1616,N_29594,N_29845);
nand UO_1617 (O_1617,N_29504,N_29700);
or UO_1618 (O_1618,N_29474,N_29527);
nand UO_1619 (O_1619,N_29786,N_29228);
and UO_1620 (O_1620,N_29881,N_29632);
or UO_1621 (O_1621,N_29978,N_29409);
xor UO_1622 (O_1622,N_29492,N_29487);
or UO_1623 (O_1623,N_29547,N_29064);
or UO_1624 (O_1624,N_29646,N_29994);
nand UO_1625 (O_1625,N_29291,N_29930);
or UO_1626 (O_1626,N_29693,N_29426);
and UO_1627 (O_1627,N_29710,N_29485);
or UO_1628 (O_1628,N_29348,N_29888);
or UO_1629 (O_1629,N_29541,N_29145);
nand UO_1630 (O_1630,N_29766,N_29395);
or UO_1631 (O_1631,N_29700,N_29785);
or UO_1632 (O_1632,N_29719,N_29078);
nor UO_1633 (O_1633,N_29864,N_29195);
xor UO_1634 (O_1634,N_29333,N_29610);
nand UO_1635 (O_1635,N_29690,N_29839);
xor UO_1636 (O_1636,N_29893,N_29736);
nand UO_1637 (O_1637,N_29584,N_29679);
nand UO_1638 (O_1638,N_29531,N_29885);
xor UO_1639 (O_1639,N_29088,N_29000);
nor UO_1640 (O_1640,N_29636,N_29606);
or UO_1641 (O_1641,N_29408,N_29405);
xnor UO_1642 (O_1642,N_29725,N_29890);
xor UO_1643 (O_1643,N_29463,N_29320);
and UO_1644 (O_1644,N_29355,N_29969);
nand UO_1645 (O_1645,N_29571,N_29477);
nand UO_1646 (O_1646,N_29725,N_29615);
nor UO_1647 (O_1647,N_29506,N_29192);
xor UO_1648 (O_1648,N_29315,N_29128);
nand UO_1649 (O_1649,N_29117,N_29710);
xnor UO_1650 (O_1650,N_29853,N_29957);
nor UO_1651 (O_1651,N_29830,N_29251);
nor UO_1652 (O_1652,N_29935,N_29592);
or UO_1653 (O_1653,N_29828,N_29435);
xnor UO_1654 (O_1654,N_29961,N_29500);
or UO_1655 (O_1655,N_29942,N_29891);
nor UO_1656 (O_1656,N_29756,N_29860);
and UO_1657 (O_1657,N_29333,N_29403);
nor UO_1658 (O_1658,N_29341,N_29367);
nand UO_1659 (O_1659,N_29658,N_29768);
and UO_1660 (O_1660,N_29651,N_29448);
nor UO_1661 (O_1661,N_29992,N_29817);
and UO_1662 (O_1662,N_29537,N_29144);
nand UO_1663 (O_1663,N_29823,N_29036);
nand UO_1664 (O_1664,N_29503,N_29505);
nand UO_1665 (O_1665,N_29683,N_29173);
and UO_1666 (O_1666,N_29104,N_29124);
nand UO_1667 (O_1667,N_29023,N_29359);
and UO_1668 (O_1668,N_29171,N_29634);
nor UO_1669 (O_1669,N_29930,N_29271);
and UO_1670 (O_1670,N_29963,N_29998);
nor UO_1671 (O_1671,N_29977,N_29014);
or UO_1672 (O_1672,N_29628,N_29937);
nand UO_1673 (O_1673,N_29563,N_29522);
xnor UO_1674 (O_1674,N_29380,N_29849);
xnor UO_1675 (O_1675,N_29240,N_29106);
xor UO_1676 (O_1676,N_29774,N_29667);
or UO_1677 (O_1677,N_29295,N_29805);
nor UO_1678 (O_1678,N_29077,N_29841);
and UO_1679 (O_1679,N_29749,N_29595);
nor UO_1680 (O_1680,N_29680,N_29093);
xnor UO_1681 (O_1681,N_29998,N_29787);
or UO_1682 (O_1682,N_29413,N_29570);
or UO_1683 (O_1683,N_29967,N_29568);
and UO_1684 (O_1684,N_29633,N_29415);
xnor UO_1685 (O_1685,N_29308,N_29933);
and UO_1686 (O_1686,N_29555,N_29592);
or UO_1687 (O_1687,N_29094,N_29496);
nand UO_1688 (O_1688,N_29884,N_29928);
and UO_1689 (O_1689,N_29394,N_29728);
or UO_1690 (O_1690,N_29974,N_29607);
and UO_1691 (O_1691,N_29928,N_29310);
and UO_1692 (O_1692,N_29389,N_29469);
and UO_1693 (O_1693,N_29769,N_29567);
or UO_1694 (O_1694,N_29162,N_29575);
nand UO_1695 (O_1695,N_29711,N_29247);
nor UO_1696 (O_1696,N_29748,N_29602);
nor UO_1697 (O_1697,N_29468,N_29101);
xnor UO_1698 (O_1698,N_29229,N_29631);
xnor UO_1699 (O_1699,N_29989,N_29637);
nor UO_1700 (O_1700,N_29123,N_29016);
xnor UO_1701 (O_1701,N_29375,N_29154);
nor UO_1702 (O_1702,N_29553,N_29647);
or UO_1703 (O_1703,N_29948,N_29648);
xor UO_1704 (O_1704,N_29853,N_29466);
or UO_1705 (O_1705,N_29705,N_29523);
nand UO_1706 (O_1706,N_29042,N_29063);
xnor UO_1707 (O_1707,N_29027,N_29075);
or UO_1708 (O_1708,N_29147,N_29665);
and UO_1709 (O_1709,N_29759,N_29515);
nand UO_1710 (O_1710,N_29243,N_29034);
nor UO_1711 (O_1711,N_29635,N_29602);
xnor UO_1712 (O_1712,N_29039,N_29769);
nand UO_1713 (O_1713,N_29764,N_29716);
nand UO_1714 (O_1714,N_29916,N_29573);
xor UO_1715 (O_1715,N_29756,N_29629);
nand UO_1716 (O_1716,N_29004,N_29307);
or UO_1717 (O_1717,N_29069,N_29755);
nand UO_1718 (O_1718,N_29602,N_29885);
nor UO_1719 (O_1719,N_29740,N_29832);
nor UO_1720 (O_1720,N_29722,N_29454);
nor UO_1721 (O_1721,N_29169,N_29390);
and UO_1722 (O_1722,N_29244,N_29011);
or UO_1723 (O_1723,N_29935,N_29784);
and UO_1724 (O_1724,N_29330,N_29086);
nor UO_1725 (O_1725,N_29925,N_29779);
or UO_1726 (O_1726,N_29878,N_29595);
nand UO_1727 (O_1727,N_29086,N_29838);
and UO_1728 (O_1728,N_29159,N_29618);
or UO_1729 (O_1729,N_29550,N_29150);
or UO_1730 (O_1730,N_29885,N_29267);
xnor UO_1731 (O_1731,N_29611,N_29567);
nand UO_1732 (O_1732,N_29553,N_29779);
nand UO_1733 (O_1733,N_29707,N_29054);
nand UO_1734 (O_1734,N_29300,N_29508);
nor UO_1735 (O_1735,N_29131,N_29449);
and UO_1736 (O_1736,N_29370,N_29317);
or UO_1737 (O_1737,N_29558,N_29205);
nor UO_1738 (O_1738,N_29551,N_29100);
or UO_1739 (O_1739,N_29701,N_29333);
nor UO_1740 (O_1740,N_29013,N_29220);
nor UO_1741 (O_1741,N_29496,N_29559);
and UO_1742 (O_1742,N_29350,N_29335);
or UO_1743 (O_1743,N_29313,N_29260);
xnor UO_1744 (O_1744,N_29488,N_29070);
xnor UO_1745 (O_1745,N_29817,N_29628);
and UO_1746 (O_1746,N_29636,N_29223);
nor UO_1747 (O_1747,N_29405,N_29651);
nor UO_1748 (O_1748,N_29378,N_29398);
and UO_1749 (O_1749,N_29536,N_29346);
xor UO_1750 (O_1750,N_29108,N_29866);
and UO_1751 (O_1751,N_29619,N_29855);
xor UO_1752 (O_1752,N_29380,N_29870);
or UO_1753 (O_1753,N_29938,N_29176);
nand UO_1754 (O_1754,N_29566,N_29695);
nor UO_1755 (O_1755,N_29625,N_29896);
xor UO_1756 (O_1756,N_29700,N_29148);
or UO_1757 (O_1757,N_29866,N_29632);
nand UO_1758 (O_1758,N_29317,N_29215);
and UO_1759 (O_1759,N_29771,N_29118);
xnor UO_1760 (O_1760,N_29708,N_29794);
and UO_1761 (O_1761,N_29827,N_29266);
nor UO_1762 (O_1762,N_29781,N_29857);
nand UO_1763 (O_1763,N_29991,N_29435);
xnor UO_1764 (O_1764,N_29762,N_29702);
and UO_1765 (O_1765,N_29179,N_29509);
xor UO_1766 (O_1766,N_29727,N_29434);
nor UO_1767 (O_1767,N_29954,N_29666);
xor UO_1768 (O_1768,N_29172,N_29842);
xor UO_1769 (O_1769,N_29346,N_29464);
and UO_1770 (O_1770,N_29160,N_29734);
or UO_1771 (O_1771,N_29501,N_29028);
nor UO_1772 (O_1772,N_29933,N_29562);
and UO_1773 (O_1773,N_29423,N_29400);
xor UO_1774 (O_1774,N_29152,N_29971);
nand UO_1775 (O_1775,N_29107,N_29976);
and UO_1776 (O_1776,N_29019,N_29953);
and UO_1777 (O_1777,N_29277,N_29159);
and UO_1778 (O_1778,N_29581,N_29253);
xor UO_1779 (O_1779,N_29436,N_29114);
or UO_1780 (O_1780,N_29076,N_29987);
nor UO_1781 (O_1781,N_29912,N_29428);
nand UO_1782 (O_1782,N_29133,N_29056);
nand UO_1783 (O_1783,N_29599,N_29581);
xor UO_1784 (O_1784,N_29046,N_29898);
xnor UO_1785 (O_1785,N_29294,N_29830);
or UO_1786 (O_1786,N_29391,N_29985);
nor UO_1787 (O_1787,N_29090,N_29011);
nand UO_1788 (O_1788,N_29057,N_29408);
or UO_1789 (O_1789,N_29176,N_29562);
nand UO_1790 (O_1790,N_29387,N_29591);
or UO_1791 (O_1791,N_29945,N_29905);
nand UO_1792 (O_1792,N_29443,N_29386);
or UO_1793 (O_1793,N_29350,N_29520);
nor UO_1794 (O_1794,N_29076,N_29083);
nand UO_1795 (O_1795,N_29148,N_29684);
and UO_1796 (O_1796,N_29845,N_29065);
xor UO_1797 (O_1797,N_29936,N_29276);
nor UO_1798 (O_1798,N_29588,N_29919);
xnor UO_1799 (O_1799,N_29799,N_29333);
or UO_1800 (O_1800,N_29760,N_29699);
and UO_1801 (O_1801,N_29901,N_29624);
nand UO_1802 (O_1802,N_29541,N_29882);
or UO_1803 (O_1803,N_29227,N_29716);
nand UO_1804 (O_1804,N_29350,N_29011);
or UO_1805 (O_1805,N_29179,N_29300);
nand UO_1806 (O_1806,N_29265,N_29275);
and UO_1807 (O_1807,N_29627,N_29317);
nand UO_1808 (O_1808,N_29765,N_29439);
xor UO_1809 (O_1809,N_29283,N_29188);
or UO_1810 (O_1810,N_29455,N_29477);
nand UO_1811 (O_1811,N_29653,N_29677);
and UO_1812 (O_1812,N_29570,N_29244);
and UO_1813 (O_1813,N_29814,N_29916);
or UO_1814 (O_1814,N_29332,N_29860);
nand UO_1815 (O_1815,N_29221,N_29831);
or UO_1816 (O_1816,N_29701,N_29902);
nand UO_1817 (O_1817,N_29240,N_29074);
nor UO_1818 (O_1818,N_29048,N_29084);
nand UO_1819 (O_1819,N_29181,N_29950);
or UO_1820 (O_1820,N_29487,N_29376);
nand UO_1821 (O_1821,N_29674,N_29619);
or UO_1822 (O_1822,N_29092,N_29507);
or UO_1823 (O_1823,N_29025,N_29220);
xor UO_1824 (O_1824,N_29637,N_29865);
and UO_1825 (O_1825,N_29253,N_29449);
and UO_1826 (O_1826,N_29518,N_29515);
nor UO_1827 (O_1827,N_29881,N_29675);
xnor UO_1828 (O_1828,N_29745,N_29321);
nand UO_1829 (O_1829,N_29305,N_29513);
nor UO_1830 (O_1830,N_29186,N_29209);
xor UO_1831 (O_1831,N_29421,N_29424);
nand UO_1832 (O_1832,N_29745,N_29285);
nand UO_1833 (O_1833,N_29663,N_29187);
xor UO_1834 (O_1834,N_29141,N_29340);
and UO_1835 (O_1835,N_29025,N_29822);
nor UO_1836 (O_1836,N_29720,N_29500);
nand UO_1837 (O_1837,N_29280,N_29555);
or UO_1838 (O_1838,N_29447,N_29379);
and UO_1839 (O_1839,N_29178,N_29365);
or UO_1840 (O_1840,N_29080,N_29138);
and UO_1841 (O_1841,N_29119,N_29295);
or UO_1842 (O_1842,N_29831,N_29410);
and UO_1843 (O_1843,N_29723,N_29177);
xnor UO_1844 (O_1844,N_29457,N_29629);
nor UO_1845 (O_1845,N_29820,N_29217);
nand UO_1846 (O_1846,N_29819,N_29479);
nand UO_1847 (O_1847,N_29671,N_29458);
nor UO_1848 (O_1848,N_29309,N_29271);
nor UO_1849 (O_1849,N_29092,N_29759);
xor UO_1850 (O_1850,N_29128,N_29267);
xnor UO_1851 (O_1851,N_29372,N_29667);
or UO_1852 (O_1852,N_29674,N_29845);
nor UO_1853 (O_1853,N_29893,N_29884);
and UO_1854 (O_1854,N_29467,N_29883);
and UO_1855 (O_1855,N_29450,N_29600);
nor UO_1856 (O_1856,N_29351,N_29063);
nor UO_1857 (O_1857,N_29857,N_29480);
or UO_1858 (O_1858,N_29333,N_29602);
and UO_1859 (O_1859,N_29296,N_29896);
nor UO_1860 (O_1860,N_29400,N_29802);
or UO_1861 (O_1861,N_29752,N_29200);
xnor UO_1862 (O_1862,N_29830,N_29353);
or UO_1863 (O_1863,N_29659,N_29136);
nor UO_1864 (O_1864,N_29859,N_29767);
nor UO_1865 (O_1865,N_29366,N_29883);
nand UO_1866 (O_1866,N_29094,N_29407);
and UO_1867 (O_1867,N_29500,N_29125);
and UO_1868 (O_1868,N_29771,N_29663);
xnor UO_1869 (O_1869,N_29434,N_29859);
and UO_1870 (O_1870,N_29803,N_29541);
nor UO_1871 (O_1871,N_29653,N_29731);
nand UO_1872 (O_1872,N_29377,N_29460);
nor UO_1873 (O_1873,N_29970,N_29692);
nand UO_1874 (O_1874,N_29044,N_29519);
nand UO_1875 (O_1875,N_29356,N_29096);
or UO_1876 (O_1876,N_29615,N_29117);
xnor UO_1877 (O_1877,N_29882,N_29663);
or UO_1878 (O_1878,N_29987,N_29445);
nor UO_1879 (O_1879,N_29264,N_29328);
and UO_1880 (O_1880,N_29508,N_29413);
or UO_1881 (O_1881,N_29600,N_29311);
xnor UO_1882 (O_1882,N_29267,N_29172);
nor UO_1883 (O_1883,N_29242,N_29686);
xnor UO_1884 (O_1884,N_29216,N_29990);
nand UO_1885 (O_1885,N_29536,N_29116);
nor UO_1886 (O_1886,N_29445,N_29998);
or UO_1887 (O_1887,N_29921,N_29170);
nor UO_1888 (O_1888,N_29645,N_29043);
nor UO_1889 (O_1889,N_29693,N_29835);
xnor UO_1890 (O_1890,N_29115,N_29820);
nand UO_1891 (O_1891,N_29261,N_29214);
nand UO_1892 (O_1892,N_29411,N_29252);
nand UO_1893 (O_1893,N_29506,N_29443);
and UO_1894 (O_1894,N_29690,N_29447);
nor UO_1895 (O_1895,N_29428,N_29141);
or UO_1896 (O_1896,N_29687,N_29492);
and UO_1897 (O_1897,N_29792,N_29769);
nor UO_1898 (O_1898,N_29277,N_29979);
xor UO_1899 (O_1899,N_29198,N_29923);
and UO_1900 (O_1900,N_29427,N_29941);
xnor UO_1901 (O_1901,N_29881,N_29926);
nand UO_1902 (O_1902,N_29025,N_29907);
nor UO_1903 (O_1903,N_29738,N_29548);
or UO_1904 (O_1904,N_29241,N_29543);
xnor UO_1905 (O_1905,N_29097,N_29105);
nor UO_1906 (O_1906,N_29511,N_29989);
xnor UO_1907 (O_1907,N_29891,N_29533);
nor UO_1908 (O_1908,N_29712,N_29417);
and UO_1909 (O_1909,N_29622,N_29193);
and UO_1910 (O_1910,N_29080,N_29251);
nor UO_1911 (O_1911,N_29914,N_29493);
and UO_1912 (O_1912,N_29003,N_29030);
and UO_1913 (O_1913,N_29532,N_29325);
nand UO_1914 (O_1914,N_29555,N_29866);
and UO_1915 (O_1915,N_29592,N_29548);
nor UO_1916 (O_1916,N_29794,N_29338);
and UO_1917 (O_1917,N_29515,N_29764);
xor UO_1918 (O_1918,N_29053,N_29074);
nand UO_1919 (O_1919,N_29575,N_29500);
nand UO_1920 (O_1920,N_29974,N_29509);
nand UO_1921 (O_1921,N_29440,N_29766);
and UO_1922 (O_1922,N_29020,N_29447);
nand UO_1923 (O_1923,N_29946,N_29719);
or UO_1924 (O_1924,N_29308,N_29376);
and UO_1925 (O_1925,N_29728,N_29920);
xnor UO_1926 (O_1926,N_29000,N_29266);
xor UO_1927 (O_1927,N_29542,N_29433);
nor UO_1928 (O_1928,N_29416,N_29200);
or UO_1929 (O_1929,N_29894,N_29521);
xor UO_1930 (O_1930,N_29255,N_29863);
nand UO_1931 (O_1931,N_29602,N_29935);
or UO_1932 (O_1932,N_29882,N_29564);
nor UO_1933 (O_1933,N_29447,N_29201);
or UO_1934 (O_1934,N_29713,N_29047);
or UO_1935 (O_1935,N_29020,N_29487);
xor UO_1936 (O_1936,N_29736,N_29355);
or UO_1937 (O_1937,N_29013,N_29293);
nor UO_1938 (O_1938,N_29875,N_29321);
or UO_1939 (O_1939,N_29532,N_29817);
nor UO_1940 (O_1940,N_29215,N_29570);
and UO_1941 (O_1941,N_29702,N_29903);
nand UO_1942 (O_1942,N_29036,N_29617);
or UO_1943 (O_1943,N_29705,N_29912);
nor UO_1944 (O_1944,N_29777,N_29274);
nand UO_1945 (O_1945,N_29278,N_29371);
nor UO_1946 (O_1946,N_29411,N_29660);
xor UO_1947 (O_1947,N_29067,N_29534);
and UO_1948 (O_1948,N_29411,N_29476);
nand UO_1949 (O_1949,N_29025,N_29217);
and UO_1950 (O_1950,N_29020,N_29065);
nand UO_1951 (O_1951,N_29561,N_29435);
and UO_1952 (O_1952,N_29764,N_29609);
nand UO_1953 (O_1953,N_29987,N_29325);
xor UO_1954 (O_1954,N_29548,N_29214);
and UO_1955 (O_1955,N_29969,N_29795);
xnor UO_1956 (O_1956,N_29635,N_29728);
and UO_1957 (O_1957,N_29803,N_29145);
and UO_1958 (O_1958,N_29001,N_29184);
xor UO_1959 (O_1959,N_29287,N_29775);
or UO_1960 (O_1960,N_29990,N_29274);
xor UO_1961 (O_1961,N_29900,N_29929);
or UO_1962 (O_1962,N_29075,N_29125);
nor UO_1963 (O_1963,N_29512,N_29354);
xnor UO_1964 (O_1964,N_29490,N_29750);
nor UO_1965 (O_1965,N_29971,N_29728);
nor UO_1966 (O_1966,N_29979,N_29145);
and UO_1967 (O_1967,N_29004,N_29200);
and UO_1968 (O_1968,N_29452,N_29025);
or UO_1969 (O_1969,N_29064,N_29388);
or UO_1970 (O_1970,N_29301,N_29579);
xnor UO_1971 (O_1971,N_29588,N_29762);
and UO_1972 (O_1972,N_29083,N_29718);
xnor UO_1973 (O_1973,N_29555,N_29898);
and UO_1974 (O_1974,N_29145,N_29742);
nand UO_1975 (O_1975,N_29805,N_29216);
or UO_1976 (O_1976,N_29099,N_29904);
or UO_1977 (O_1977,N_29323,N_29614);
nand UO_1978 (O_1978,N_29963,N_29182);
and UO_1979 (O_1979,N_29668,N_29639);
nor UO_1980 (O_1980,N_29702,N_29205);
nand UO_1981 (O_1981,N_29300,N_29526);
nor UO_1982 (O_1982,N_29364,N_29483);
or UO_1983 (O_1983,N_29512,N_29736);
and UO_1984 (O_1984,N_29566,N_29286);
or UO_1985 (O_1985,N_29242,N_29221);
or UO_1986 (O_1986,N_29351,N_29518);
nor UO_1987 (O_1987,N_29679,N_29165);
xnor UO_1988 (O_1988,N_29734,N_29707);
and UO_1989 (O_1989,N_29014,N_29595);
and UO_1990 (O_1990,N_29456,N_29505);
xor UO_1991 (O_1991,N_29578,N_29824);
or UO_1992 (O_1992,N_29546,N_29732);
xnor UO_1993 (O_1993,N_29596,N_29793);
and UO_1994 (O_1994,N_29008,N_29070);
nand UO_1995 (O_1995,N_29538,N_29997);
or UO_1996 (O_1996,N_29621,N_29132);
nor UO_1997 (O_1997,N_29456,N_29127);
xor UO_1998 (O_1998,N_29667,N_29225);
xor UO_1999 (O_1999,N_29430,N_29204);
or UO_2000 (O_2000,N_29251,N_29821);
nand UO_2001 (O_2001,N_29028,N_29042);
nor UO_2002 (O_2002,N_29894,N_29728);
xor UO_2003 (O_2003,N_29033,N_29063);
nand UO_2004 (O_2004,N_29989,N_29952);
nand UO_2005 (O_2005,N_29937,N_29274);
nand UO_2006 (O_2006,N_29903,N_29281);
or UO_2007 (O_2007,N_29095,N_29426);
or UO_2008 (O_2008,N_29494,N_29763);
nand UO_2009 (O_2009,N_29057,N_29175);
nor UO_2010 (O_2010,N_29926,N_29290);
xor UO_2011 (O_2011,N_29406,N_29733);
nor UO_2012 (O_2012,N_29613,N_29382);
nor UO_2013 (O_2013,N_29615,N_29843);
and UO_2014 (O_2014,N_29034,N_29124);
nor UO_2015 (O_2015,N_29202,N_29240);
and UO_2016 (O_2016,N_29329,N_29649);
nor UO_2017 (O_2017,N_29486,N_29696);
xnor UO_2018 (O_2018,N_29751,N_29806);
nor UO_2019 (O_2019,N_29066,N_29540);
xor UO_2020 (O_2020,N_29690,N_29844);
or UO_2021 (O_2021,N_29564,N_29402);
and UO_2022 (O_2022,N_29232,N_29946);
nor UO_2023 (O_2023,N_29327,N_29968);
nand UO_2024 (O_2024,N_29707,N_29912);
nor UO_2025 (O_2025,N_29244,N_29938);
and UO_2026 (O_2026,N_29111,N_29388);
and UO_2027 (O_2027,N_29332,N_29312);
nor UO_2028 (O_2028,N_29914,N_29644);
nor UO_2029 (O_2029,N_29323,N_29526);
or UO_2030 (O_2030,N_29856,N_29999);
xor UO_2031 (O_2031,N_29083,N_29141);
nand UO_2032 (O_2032,N_29138,N_29222);
or UO_2033 (O_2033,N_29206,N_29831);
nor UO_2034 (O_2034,N_29750,N_29107);
and UO_2035 (O_2035,N_29669,N_29464);
nand UO_2036 (O_2036,N_29693,N_29468);
nor UO_2037 (O_2037,N_29715,N_29805);
and UO_2038 (O_2038,N_29393,N_29676);
nor UO_2039 (O_2039,N_29996,N_29474);
nand UO_2040 (O_2040,N_29002,N_29892);
xor UO_2041 (O_2041,N_29305,N_29633);
nand UO_2042 (O_2042,N_29516,N_29364);
and UO_2043 (O_2043,N_29784,N_29661);
nor UO_2044 (O_2044,N_29990,N_29936);
nand UO_2045 (O_2045,N_29901,N_29456);
or UO_2046 (O_2046,N_29021,N_29635);
and UO_2047 (O_2047,N_29500,N_29316);
nand UO_2048 (O_2048,N_29113,N_29782);
or UO_2049 (O_2049,N_29138,N_29530);
and UO_2050 (O_2050,N_29304,N_29835);
nand UO_2051 (O_2051,N_29095,N_29741);
or UO_2052 (O_2052,N_29756,N_29813);
or UO_2053 (O_2053,N_29858,N_29760);
and UO_2054 (O_2054,N_29889,N_29282);
or UO_2055 (O_2055,N_29561,N_29899);
nor UO_2056 (O_2056,N_29797,N_29891);
or UO_2057 (O_2057,N_29418,N_29343);
and UO_2058 (O_2058,N_29634,N_29913);
or UO_2059 (O_2059,N_29195,N_29413);
nor UO_2060 (O_2060,N_29193,N_29764);
or UO_2061 (O_2061,N_29234,N_29697);
xnor UO_2062 (O_2062,N_29243,N_29011);
or UO_2063 (O_2063,N_29377,N_29093);
nor UO_2064 (O_2064,N_29533,N_29696);
xnor UO_2065 (O_2065,N_29003,N_29238);
xor UO_2066 (O_2066,N_29739,N_29850);
nor UO_2067 (O_2067,N_29111,N_29114);
or UO_2068 (O_2068,N_29338,N_29923);
or UO_2069 (O_2069,N_29663,N_29634);
nor UO_2070 (O_2070,N_29316,N_29220);
nand UO_2071 (O_2071,N_29819,N_29426);
or UO_2072 (O_2072,N_29121,N_29898);
nor UO_2073 (O_2073,N_29486,N_29196);
and UO_2074 (O_2074,N_29981,N_29677);
and UO_2075 (O_2075,N_29254,N_29299);
or UO_2076 (O_2076,N_29338,N_29102);
or UO_2077 (O_2077,N_29530,N_29135);
nand UO_2078 (O_2078,N_29003,N_29559);
and UO_2079 (O_2079,N_29420,N_29111);
or UO_2080 (O_2080,N_29668,N_29512);
xnor UO_2081 (O_2081,N_29976,N_29410);
nand UO_2082 (O_2082,N_29230,N_29423);
and UO_2083 (O_2083,N_29703,N_29773);
and UO_2084 (O_2084,N_29732,N_29359);
or UO_2085 (O_2085,N_29615,N_29186);
nand UO_2086 (O_2086,N_29391,N_29992);
xnor UO_2087 (O_2087,N_29795,N_29544);
xor UO_2088 (O_2088,N_29593,N_29467);
xor UO_2089 (O_2089,N_29754,N_29281);
nor UO_2090 (O_2090,N_29269,N_29775);
nor UO_2091 (O_2091,N_29387,N_29656);
nand UO_2092 (O_2092,N_29311,N_29281);
xor UO_2093 (O_2093,N_29474,N_29027);
or UO_2094 (O_2094,N_29213,N_29163);
and UO_2095 (O_2095,N_29047,N_29808);
and UO_2096 (O_2096,N_29640,N_29157);
xor UO_2097 (O_2097,N_29371,N_29594);
and UO_2098 (O_2098,N_29882,N_29631);
and UO_2099 (O_2099,N_29944,N_29196);
nand UO_2100 (O_2100,N_29071,N_29293);
or UO_2101 (O_2101,N_29249,N_29938);
nor UO_2102 (O_2102,N_29666,N_29004);
and UO_2103 (O_2103,N_29232,N_29863);
xnor UO_2104 (O_2104,N_29466,N_29137);
and UO_2105 (O_2105,N_29277,N_29289);
xor UO_2106 (O_2106,N_29245,N_29132);
and UO_2107 (O_2107,N_29631,N_29140);
or UO_2108 (O_2108,N_29702,N_29886);
nor UO_2109 (O_2109,N_29914,N_29373);
xnor UO_2110 (O_2110,N_29103,N_29987);
or UO_2111 (O_2111,N_29539,N_29948);
xor UO_2112 (O_2112,N_29921,N_29472);
and UO_2113 (O_2113,N_29828,N_29113);
and UO_2114 (O_2114,N_29835,N_29183);
nor UO_2115 (O_2115,N_29583,N_29227);
xnor UO_2116 (O_2116,N_29039,N_29719);
and UO_2117 (O_2117,N_29443,N_29552);
nand UO_2118 (O_2118,N_29072,N_29538);
xnor UO_2119 (O_2119,N_29489,N_29527);
or UO_2120 (O_2120,N_29832,N_29167);
nand UO_2121 (O_2121,N_29301,N_29611);
nor UO_2122 (O_2122,N_29020,N_29673);
nand UO_2123 (O_2123,N_29617,N_29497);
or UO_2124 (O_2124,N_29629,N_29739);
nand UO_2125 (O_2125,N_29016,N_29497);
nand UO_2126 (O_2126,N_29067,N_29733);
xor UO_2127 (O_2127,N_29856,N_29515);
or UO_2128 (O_2128,N_29734,N_29226);
or UO_2129 (O_2129,N_29978,N_29309);
or UO_2130 (O_2130,N_29346,N_29791);
xor UO_2131 (O_2131,N_29502,N_29223);
or UO_2132 (O_2132,N_29655,N_29867);
xnor UO_2133 (O_2133,N_29237,N_29888);
and UO_2134 (O_2134,N_29081,N_29336);
nand UO_2135 (O_2135,N_29630,N_29076);
nor UO_2136 (O_2136,N_29260,N_29064);
nor UO_2137 (O_2137,N_29722,N_29811);
nand UO_2138 (O_2138,N_29862,N_29342);
and UO_2139 (O_2139,N_29425,N_29491);
and UO_2140 (O_2140,N_29674,N_29481);
nand UO_2141 (O_2141,N_29816,N_29835);
xor UO_2142 (O_2142,N_29853,N_29723);
nand UO_2143 (O_2143,N_29931,N_29940);
xor UO_2144 (O_2144,N_29890,N_29765);
nor UO_2145 (O_2145,N_29464,N_29785);
nor UO_2146 (O_2146,N_29242,N_29649);
nor UO_2147 (O_2147,N_29745,N_29779);
and UO_2148 (O_2148,N_29870,N_29544);
nor UO_2149 (O_2149,N_29072,N_29473);
nand UO_2150 (O_2150,N_29891,N_29267);
and UO_2151 (O_2151,N_29010,N_29641);
nor UO_2152 (O_2152,N_29312,N_29392);
nand UO_2153 (O_2153,N_29906,N_29336);
or UO_2154 (O_2154,N_29296,N_29653);
nand UO_2155 (O_2155,N_29038,N_29827);
xnor UO_2156 (O_2156,N_29918,N_29231);
or UO_2157 (O_2157,N_29509,N_29296);
nor UO_2158 (O_2158,N_29005,N_29511);
or UO_2159 (O_2159,N_29937,N_29159);
xnor UO_2160 (O_2160,N_29668,N_29197);
and UO_2161 (O_2161,N_29083,N_29788);
or UO_2162 (O_2162,N_29848,N_29590);
or UO_2163 (O_2163,N_29386,N_29970);
nand UO_2164 (O_2164,N_29084,N_29794);
or UO_2165 (O_2165,N_29484,N_29519);
nor UO_2166 (O_2166,N_29993,N_29596);
nor UO_2167 (O_2167,N_29690,N_29599);
nand UO_2168 (O_2168,N_29647,N_29341);
xor UO_2169 (O_2169,N_29531,N_29978);
and UO_2170 (O_2170,N_29946,N_29519);
xor UO_2171 (O_2171,N_29543,N_29493);
nor UO_2172 (O_2172,N_29612,N_29287);
or UO_2173 (O_2173,N_29343,N_29376);
xor UO_2174 (O_2174,N_29069,N_29700);
and UO_2175 (O_2175,N_29959,N_29893);
nor UO_2176 (O_2176,N_29279,N_29268);
xor UO_2177 (O_2177,N_29278,N_29991);
or UO_2178 (O_2178,N_29817,N_29780);
nor UO_2179 (O_2179,N_29022,N_29023);
xor UO_2180 (O_2180,N_29590,N_29486);
nor UO_2181 (O_2181,N_29634,N_29764);
or UO_2182 (O_2182,N_29439,N_29030);
and UO_2183 (O_2183,N_29496,N_29277);
nor UO_2184 (O_2184,N_29748,N_29731);
xnor UO_2185 (O_2185,N_29756,N_29859);
xor UO_2186 (O_2186,N_29438,N_29141);
or UO_2187 (O_2187,N_29829,N_29294);
nor UO_2188 (O_2188,N_29867,N_29109);
nor UO_2189 (O_2189,N_29033,N_29091);
nor UO_2190 (O_2190,N_29364,N_29575);
nand UO_2191 (O_2191,N_29523,N_29388);
or UO_2192 (O_2192,N_29696,N_29489);
xnor UO_2193 (O_2193,N_29299,N_29635);
nand UO_2194 (O_2194,N_29680,N_29554);
xor UO_2195 (O_2195,N_29080,N_29875);
nand UO_2196 (O_2196,N_29109,N_29427);
or UO_2197 (O_2197,N_29706,N_29839);
nor UO_2198 (O_2198,N_29673,N_29566);
xnor UO_2199 (O_2199,N_29669,N_29159);
and UO_2200 (O_2200,N_29687,N_29719);
nand UO_2201 (O_2201,N_29531,N_29308);
nand UO_2202 (O_2202,N_29848,N_29609);
xor UO_2203 (O_2203,N_29174,N_29221);
nor UO_2204 (O_2204,N_29340,N_29731);
or UO_2205 (O_2205,N_29439,N_29035);
and UO_2206 (O_2206,N_29500,N_29864);
xor UO_2207 (O_2207,N_29071,N_29281);
xnor UO_2208 (O_2208,N_29617,N_29499);
nor UO_2209 (O_2209,N_29071,N_29349);
nand UO_2210 (O_2210,N_29349,N_29352);
and UO_2211 (O_2211,N_29517,N_29837);
nor UO_2212 (O_2212,N_29751,N_29558);
or UO_2213 (O_2213,N_29445,N_29793);
nand UO_2214 (O_2214,N_29621,N_29462);
nand UO_2215 (O_2215,N_29664,N_29373);
or UO_2216 (O_2216,N_29499,N_29981);
xnor UO_2217 (O_2217,N_29395,N_29637);
nand UO_2218 (O_2218,N_29883,N_29332);
or UO_2219 (O_2219,N_29234,N_29481);
xor UO_2220 (O_2220,N_29278,N_29641);
nand UO_2221 (O_2221,N_29560,N_29451);
nor UO_2222 (O_2222,N_29706,N_29328);
and UO_2223 (O_2223,N_29427,N_29727);
nor UO_2224 (O_2224,N_29711,N_29767);
and UO_2225 (O_2225,N_29845,N_29762);
nor UO_2226 (O_2226,N_29256,N_29108);
and UO_2227 (O_2227,N_29898,N_29803);
or UO_2228 (O_2228,N_29385,N_29606);
nor UO_2229 (O_2229,N_29004,N_29930);
nand UO_2230 (O_2230,N_29412,N_29397);
nor UO_2231 (O_2231,N_29443,N_29720);
and UO_2232 (O_2232,N_29942,N_29090);
or UO_2233 (O_2233,N_29160,N_29228);
and UO_2234 (O_2234,N_29912,N_29526);
xor UO_2235 (O_2235,N_29421,N_29729);
nor UO_2236 (O_2236,N_29121,N_29429);
and UO_2237 (O_2237,N_29301,N_29432);
nor UO_2238 (O_2238,N_29472,N_29612);
or UO_2239 (O_2239,N_29106,N_29295);
nand UO_2240 (O_2240,N_29031,N_29959);
xor UO_2241 (O_2241,N_29619,N_29045);
xor UO_2242 (O_2242,N_29395,N_29963);
nand UO_2243 (O_2243,N_29662,N_29061);
or UO_2244 (O_2244,N_29317,N_29048);
nand UO_2245 (O_2245,N_29446,N_29260);
nand UO_2246 (O_2246,N_29431,N_29095);
nor UO_2247 (O_2247,N_29561,N_29311);
and UO_2248 (O_2248,N_29387,N_29182);
nand UO_2249 (O_2249,N_29172,N_29226);
and UO_2250 (O_2250,N_29785,N_29539);
and UO_2251 (O_2251,N_29166,N_29508);
xnor UO_2252 (O_2252,N_29547,N_29409);
xor UO_2253 (O_2253,N_29314,N_29220);
nor UO_2254 (O_2254,N_29431,N_29308);
or UO_2255 (O_2255,N_29780,N_29402);
nor UO_2256 (O_2256,N_29188,N_29632);
or UO_2257 (O_2257,N_29216,N_29050);
or UO_2258 (O_2258,N_29954,N_29138);
and UO_2259 (O_2259,N_29015,N_29468);
xor UO_2260 (O_2260,N_29432,N_29071);
xnor UO_2261 (O_2261,N_29894,N_29838);
nand UO_2262 (O_2262,N_29354,N_29411);
xnor UO_2263 (O_2263,N_29062,N_29871);
nand UO_2264 (O_2264,N_29362,N_29314);
or UO_2265 (O_2265,N_29744,N_29409);
or UO_2266 (O_2266,N_29062,N_29608);
xnor UO_2267 (O_2267,N_29572,N_29080);
or UO_2268 (O_2268,N_29373,N_29461);
xor UO_2269 (O_2269,N_29597,N_29992);
nor UO_2270 (O_2270,N_29536,N_29149);
and UO_2271 (O_2271,N_29988,N_29513);
or UO_2272 (O_2272,N_29062,N_29475);
nor UO_2273 (O_2273,N_29670,N_29074);
and UO_2274 (O_2274,N_29236,N_29632);
and UO_2275 (O_2275,N_29265,N_29253);
xnor UO_2276 (O_2276,N_29459,N_29979);
xnor UO_2277 (O_2277,N_29601,N_29213);
or UO_2278 (O_2278,N_29405,N_29783);
xor UO_2279 (O_2279,N_29999,N_29643);
xor UO_2280 (O_2280,N_29380,N_29035);
nor UO_2281 (O_2281,N_29544,N_29206);
xnor UO_2282 (O_2282,N_29034,N_29871);
nor UO_2283 (O_2283,N_29984,N_29853);
nor UO_2284 (O_2284,N_29211,N_29285);
and UO_2285 (O_2285,N_29055,N_29498);
xnor UO_2286 (O_2286,N_29037,N_29504);
xor UO_2287 (O_2287,N_29492,N_29167);
nor UO_2288 (O_2288,N_29333,N_29549);
or UO_2289 (O_2289,N_29640,N_29318);
or UO_2290 (O_2290,N_29183,N_29048);
or UO_2291 (O_2291,N_29822,N_29017);
or UO_2292 (O_2292,N_29267,N_29324);
xnor UO_2293 (O_2293,N_29885,N_29883);
or UO_2294 (O_2294,N_29463,N_29157);
or UO_2295 (O_2295,N_29729,N_29133);
xnor UO_2296 (O_2296,N_29760,N_29570);
or UO_2297 (O_2297,N_29087,N_29248);
xnor UO_2298 (O_2298,N_29746,N_29106);
nand UO_2299 (O_2299,N_29325,N_29700);
nor UO_2300 (O_2300,N_29610,N_29110);
or UO_2301 (O_2301,N_29947,N_29549);
and UO_2302 (O_2302,N_29027,N_29104);
xor UO_2303 (O_2303,N_29827,N_29143);
xnor UO_2304 (O_2304,N_29664,N_29629);
xor UO_2305 (O_2305,N_29120,N_29571);
or UO_2306 (O_2306,N_29070,N_29506);
and UO_2307 (O_2307,N_29413,N_29810);
or UO_2308 (O_2308,N_29386,N_29299);
and UO_2309 (O_2309,N_29039,N_29747);
nor UO_2310 (O_2310,N_29130,N_29588);
nand UO_2311 (O_2311,N_29262,N_29095);
xor UO_2312 (O_2312,N_29468,N_29815);
nor UO_2313 (O_2313,N_29373,N_29827);
or UO_2314 (O_2314,N_29808,N_29630);
xor UO_2315 (O_2315,N_29295,N_29193);
or UO_2316 (O_2316,N_29981,N_29064);
or UO_2317 (O_2317,N_29574,N_29141);
xor UO_2318 (O_2318,N_29942,N_29786);
and UO_2319 (O_2319,N_29274,N_29546);
xor UO_2320 (O_2320,N_29696,N_29180);
xor UO_2321 (O_2321,N_29784,N_29902);
and UO_2322 (O_2322,N_29586,N_29796);
nor UO_2323 (O_2323,N_29172,N_29286);
nand UO_2324 (O_2324,N_29702,N_29824);
nand UO_2325 (O_2325,N_29665,N_29913);
xnor UO_2326 (O_2326,N_29212,N_29325);
or UO_2327 (O_2327,N_29281,N_29202);
and UO_2328 (O_2328,N_29889,N_29128);
nor UO_2329 (O_2329,N_29887,N_29238);
nor UO_2330 (O_2330,N_29675,N_29236);
xnor UO_2331 (O_2331,N_29636,N_29894);
xnor UO_2332 (O_2332,N_29935,N_29721);
or UO_2333 (O_2333,N_29455,N_29995);
nor UO_2334 (O_2334,N_29440,N_29484);
xor UO_2335 (O_2335,N_29993,N_29501);
nor UO_2336 (O_2336,N_29575,N_29164);
or UO_2337 (O_2337,N_29918,N_29098);
or UO_2338 (O_2338,N_29925,N_29350);
and UO_2339 (O_2339,N_29224,N_29362);
or UO_2340 (O_2340,N_29656,N_29982);
nand UO_2341 (O_2341,N_29878,N_29735);
nor UO_2342 (O_2342,N_29081,N_29389);
nor UO_2343 (O_2343,N_29355,N_29205);
nand UO_2344 (O_2344,N_29367,N_29401);
nand UO_2345 (O_2345,N_29925,N_29671);
nor UO_2346 (O_2346,N_29835,N_29920);
nor UO_2347 (O_2347,N_29337,N_29662);
and UO_2348 (O_2348,N_29507,N_29913);
xor UO_2349 (O_2349,N_29776,N_29148);
nor UO_2350 (O_2350,N_29816,N_29617);
nor UO_2351 (O_2351,N_29356,N_29289);
and UO_2352 (O_2352,N_29449,N_29432);
or UO_2353 (O_2353,N_29031,N_29127);
xor UO_2354 (O_2354,N_29893,N_29448);
nor UO_2355 (O_2355,N_29657,N_29265);
nor UO_2356 (O_2356,N_29158,N_29154);
xor UO_2357 (O_2357,N_29107,N_29566);
and UO_2358 (O_2358,N_29501,N_29267);
and UO_2359 (O_2359,N_29811,N_29444);
nand UO_2360 (O_2360,N_29019,N_29627);
xor UO_2361 (O_2361,N_29469,N_29784);
nor UO_2362 (O_2362,N_29828,N_29330);
nor UO_2363 (O_2363,N_29089,N_29123);
or UO_2364 (O_2364,N_29951,N_29887);
nand UO_2365 (O_2365,N_29655,N_29316);
nand UO_2366 (O_2366,N_29174,N_29653);
and UO_2367 (O_2367,N_29910,N_29550);
or UO_2368 (O_2368,N_29984,N_29697);
nor UO_2369 (O_2369,N_29697,N_29670);
or UO_2370 (O_2370,N_29038,N_29520);
xnor UO_2371 (O_2371,N_29154,N_29019);
or UO_2372 (O_2372,N_29210,N_29089);
nor UO_2373 (O_2373,N_29770,N_29283);
and UO_2374 (O_2374,N_29670,N_29003);
or UO_2375 (O_2375,N_29545,N_29355);
or UO_2376 (O_2376,N_29798,N_29433);
xnor UO_2377 (O_2377,N_29006,N_29999);
and UO_2378 (O_2378,N_29158,N_29114);
nand UO_2379 (O_2379,N_29827,N_29624);
and UO_2380 (O_2380,N_29994,N_29021);
nand UO_2381 (O_2381,N_29388,N_29547);
nand UO_2382 (O_2382,N_29546,N_29871);
and UO_2383 (O_2383,N_29128,N_29296);
nor UO_2384 (O_2384,N_29284,N_29119);
nor UO_2385 (O_2385,N_29986,N_29705);
xnor UO_2386 (O_2386,N_29827,N_29575);
or UO_2387 (O_2387,N_29344,N_29642);
and UO_2388 (O_2388,N_29166,N_29192);
and UO_2389 (O_2389,N_29994,N_29410);
nor UO_2390 (O_2390,N_29704,N_29518);
nor UO_2391 (O_2391,N_29818,N_29300);
or UO_2392 (O_2392,N_29254,N_29076);
and UO_2393 (O_2393,N_29541,N_29192);
and UO_2394 (O_2394,N_29095,N_29708);
xor UO_2395 (O_2395,N_29640,N_29139);
nor UO_2396 (O_2396,N_29875,N_29410);
and UO_2397 (O_2397,N_29015,N_29722);
and UO_2398 (O_2398,N_29816,N_29093);
or UO_2399 (O_2399,N_29507,N_29255);
nand UO_2400 (O_2400,N_29081,N_29286);
nand UO_2401 (O_2401,N_29551,N_29217);
xnor UO_2402 (O_2402,N_29581,N_29129);
or UO_2403 (O_2403,N_29858,N_29641);
and UO_2404 (O_2404,N_29418,N_29785);
or UO_2405 (O_2405,N_29509,N_29520);
or UO_2406 (O_2406,N_29819,N_29447);
nor UO_2407 (O_2407,N_29611,N_29710);
or UO_2408 (O_2408,N_29663,N_29776);
nor UO_2409 (O_2409,N_29034,N_29953);
or UO_2410 (O_2410,N_29147,N_29881);
nor UO_2411 (O_2411,N_29482,N_29057);
nor UO_2412 (O_2412,N_29617,N_29942);
and UO_2413 (O_2413,N_29001,N_29007);
and UO_2414 (O_2414,N_29918,N_29462);
nand UO_2415 (O_2415,N_29400,N_29314);
or UO_2416 (O_2416,N_29866,N_29736);
and UO_2417 (O_2417,N_29308,N_29634);
nand UO_2418 (O_2418,N_29027,N_29917);
and UO_2419 (O_2419,N_29914,N_29534);
nand UO_2420 (O_2420,N_29628,N_29683);
nor UO_2421 (O_2421,N_29372,N_29796);
nand UO_2422 (O_2422,N_29745,N_29994);
nor UO_2423 (O_2423,N_29178,N_29331);
nand UO_2424 (O_2424,N_29726,N_29056);
or UO_2425 (O_2425,N_29963,N_29720);
xor UO_2426 (O_2426,N_29317,N_29664);
and UO_2427 (O_2427,N_29662,N_29188);
xor UO_2428 (O_2428,N_29769,N_29501);
nor UO_2429 (O_2429,N_29470,N_29866);
or UO_2430 (O_2430,N_29215,N_29476);
xnor UO_2431 (O_2431,N_29955,N_29576);
and UO_2432 (O_2432,N_29282,N_29871);
nand UO_2433 (O_2433,N_29537,N_29793);
xnor UO_2434 (O_2434,N_29506,N_29665);
xnor UO_2435 (O_2435,N_29568,N_29652);
nor UO_2436 (O_2436,N_29852,N_29574);
or UO_2437 (O_2437,N_29331,N_29124);
nand UO_2438 (O_2438,N_29027,N_29658);
and UO_2439 (O_2439,N_29858,N_29862);
or UO_2440 (O_2440,N_29458,N_29131);
nand UO_2441 (O_2441,N_29973,N_29113);
nor UO_2442 (O_2442,N_29906,N_29129);
or UO_2443 (O_2443,N_29408,N_29497);
or UO_2444 (O_2444,N_29891,N_29041);
and UO_2445 (O_2445,N_29655,N_29146);
nand UO_2446 (O_2446,N_29267,N_29587);
nor UO_2447 (O_2447,N_29157,N_29503);
xnor UO_2448 (O_2448,N_29045,N_29551);
or UO_2449 (O_2449,N_29240,N_29731);
nor UO_2450 (O_2450,N_29093,N_29721);
and UO_2451 (O_2451,N_29654,N_29053);
xnor UO_2452 (O_2452,N_29706,N_29681);
nor UO_2453 (O_2453,N_29455,N_29697);
nand UO_2454 (O_2454,N_29829,N_29830);
nand UO_2455 (O_2455,N_29520,N_29940);
nor UO_2456 (O_2456,N_29473,N_29958);
nor UO_2457 (O_2457,N_29153,N_29516);
xnor UO_2458 (O_2458,N_29169,N_29771);
xnor UO_2459 (O_2459,N_29294,N_29568);
nand UO_2460 (O_2460,N_29004,N_29335);
nand UO_2461 (O_2461,N_29938,N_29490);
or UO_2462 (O_2462,N_29434,N_29736);
or UO_2463 (O_2463,N_29076,N_29414);
and UO_2464 (O_2464,N_29736,N_29263);
or UO_2465 (O_2465,N_29438,N_29109);
or UO_2466 (O_2466,N_29989,N_29323);
and UO_2467 (O_2467,N_29286,N_29156);
or UO_2468 (O_2468,N_29742,N_29279);
and UO_2469 (O_2469,N_29754,N_29083);
nand UO_2470 (O_2470,N_29165,N_29633);
or UO_2471 (O_2471,N_29303,N_29360);
or UO_2472 (O_2472,N_29970,N_29427);
xnor UO_2473 (O_2473,N_29493,N_29761);
nand UO_2474 (O_2474,N_29273,N_29620);
xnor UO_2475 (O_2475,N_29638,N_29459);
or UO_2476 (O_2476,N_29034,N_29939);
and UO_2477 (O_2477,N_29901,N_29221);
or UO_2478 (O_2478,N_29914,N_29846);
nor UO_2479 (O_2479,N_29546,N_29409);
nand UO_2480 (O_2480,N_29785,N_29592);
xor UO_2481 (O_2481,N_29659,N_29879);
or UO_2482 (O_2482,N_29090,N_29158);
and UO_2483 (O_2483,N_29162,N_29414);
or UO_2484 (O_2484,N_29168,N_29615);
nand UO_2485 (O_2485,N_29300,N_29838);
xor UO_2486 (O_2486,N_29000,N_29948);
and UO_2487 (O_2487,N_29376,N_29778);
xor UO_2488 (O_2488,N_29753,N_29198);
and UO_2489 (O_2489,N_29020,N_29208);
xor UO_2490 (O_2490,N_29519,N_29148);
and UO_2491 (O_2491,N_29688,N_29860);
or UO_2492 (O_2492,N_29364,N_29786);
xor UO_2493 (O_2493,N_29151,N_29942);
and UO_2494 (O_2494,N_29915,N_29849);
nand UO_2495 (O_2495,N_29061,N_29689);
nor UO_2496 (O_2496,N_29726,N_29866);
nand UO_2497 (O_2497,N_29277,N_29377);
xnor UO_2498 (O_2498,N_29135,N_29615);
and UO_2499 (O_2499,N_29032,N_29489);
and UO_2500 (O_2500,N_29319,N_29226);
and UO_2501 (O_2501,N_29674,N_29285);
and UO_2502 (O_2502,N_29482,N_29156);
and UO_2503 (O_2503,N_29631,N_29379);
or UO_2504 (O_2504,N_29308,N_29154);
and UO_2505 (O_2505,N_29619,N_29856);
or UO_2506 (O_2506,N_29983,N_29186);
nand UO_2507 (O_2507,N_29378,N_29822);
and UO_2508 (O_2508,N_29933,N_29419);
xor UO_2509 (O_2509,N_29719,N_29905);
nand UO_2510 (O_2510,N_29941,N_29660);
or UO_2511 (O_2511,N_29762,N_29631);
or UO_2512 (O_2512,N_29612,N_29490);
nor UO_2513 (O_2513,N_29125,N_29177);
and UO_2514 (O_2514,N_29143,N_29796);
and UO_2515 (O_2515,N_29378,N_29781);
and UO_2516 (O_2516,N_29964,N_29362);
xor UO_2517 (O_2517,N_29767,N_29612);
or UO_2518 (O_2518,N_29414,N_29204);
or UO_2519 (O_2519,N_29271,N_29032);
and UO_2520 (O_2520,N_29370,N_29771);
and UO_2521 (O_2521,N_29698,N_29822);
nand UO_2522 (O_2522,N_29373,N_29271);
nand UO_2523 (O_2523,N_29069,N_29314);
nand UO_2524 (O_2524,N_29984,N_29020);
nand UO_2525 (O_2525,N_29451,N_29069);
and UO_2526 (O_2526,N_29502,N_29705);
xnor UO_2527 (O_2527,N_29533,N_29194);
nand UO_2528 (O_2528,N_29136,N_29470);
and UO_2529 (O_2529,N_29331,N_29937);
nand UO_2530 (O_2530,N_29799,N_29666);
nand UO_2531 (O_2531,N_29902,N_29241);
or UO_2532 (O_2532,N_29836,N_29024);
nor UO_2533 (O_2533,N_29643,N_29831);
xor UO_2534 (O_2534,N_29253,N_29059);
and UO_2535 (O_2535,N_29079,N_29500);
xor UO_2536 (O_2536,N_29197,N_29765);
nor UO_2537 (O_2537,N_29341,N_29576);
and UO_2538 (O_2538,N_29700,N_29092);
and UO_2539 (O_2539,N_29882,N_29628);
xor UO_2540 (O_2540,N_29810,N_29411);
nand UO_2541 (O_2541,N_29255,N_29275);
and UO_2542 (O_2542,N_29385,N_29618);
and UO_2543 (O_2543,N_29670,N_29352);
xnor UO_2544 (O_2544,N_29006,N_29283);
nor UO_2545 (O_2545,N_29833,N_29242);
xnor UO_2546 (O_2546,N_29678,N_29779);
or UO_2547 (O_2547,N_29076,N_29196);
nor UO_2548 (O_2548,N_29287,N_29702);
nand UO_2549 (O_2549,N_29288,N_29283);
nand UO_2550 (O_2550,N_29886,N_29298);
nand UO_2551 (O_2551,N_29052,N_29698);
nand UO_2552 (O_2552,N_29234,N_29983);
nand UO_2553 (O_2553,N_29392,N_29287);
nor UO_2554 (O_2554,N_29901,N_29891);
nand UO_2555 (O_2555,N_29474,N_29893);
xor UO_2556 (O_2556,N_29169,N_29571);
nand UO_2557 (O_2557,N_29330,N_29050);
and UO_2558 (O_2558,N_29679,N_29163);
xor UO_2559 (O_2559,N_29539,N_29227);
and UO_2560 (O_2560,N_29972,N_29864);
nor UO_2561 (O_2561,N_29342,N_29426);
or UO_2562 (O_2562,N_29885,N_29425);
or UO_2563 (O_2563,N_29604,N_29300);
nor UO_2564 (O_2564,N_29020,N_29345);
xnor UO_2565 (O_2565,N_29365,N_29597);
nand UO_2566 (O_2566,N_29192,N_29015);
nand UO_2567 (O_2567,N_29831,N_29550);
xnor UO_2568 (O_2568,N_29623,N_29393);
xor UO_2569 (O_2569,N_29887,N_29907);
or UO_2570 (O_2570,N_29429,N_29109);
xor UO_2571 (O_2571,N_29569,N_29035);
or UO_2572 (O_2572,N_29639,N_29496);
and UO_2573 (O_2573,N_29743,N_29663);
xnor UO_2574 (O_2574,N_29063,N_29529);
xor UO_2575 (O_2575,N_29574,N_29080);
and UO_2576 (O_2576,N_29240,N_29633);
and UO_2577 (O_2577,N_29310,N_29367);
xor UO_2578 (O_2578,N_29917,N_29969);
or UO_2579 (O_2579,N_29873,N_29449);
xnor UO_2580 (O_2580,N_29082,N_29979);
and UO_2581 (O_2581,N_29859,N_29640);
and UO_2582 (O_2582,N_29838,N_29379);
or UO_2583 (O_2583,N_29940,N_29858);
and UO_2584 (O_2584,N_29067,N_29631);
and UO_2585 (O_2585,N_29372,N_29217);
or UO_2586 (O_2586,N_29710,N_29431);
nand UO_2587 (O_2587,N_29047,N_29304);
xnor UO_2588 (O_2588,N_29986,N_29476);
nand UO_2589 (O_2589,N_29159,N_29089);
nor UO_2590 (O_2590,N_29961,N_29726);
or UO_2591 (O_2591,N_29289,N_29503);
xor UO_2592 (O_2592,N_29437,N_29007);
nor UO_2593 (O_2593,N_29250,N_29715);
nor UO_2594 (O_2594,N_29722,N_29782);
xor UO_2595 (O_2595,N_29476,N_29899);
nand UO_2596 (O_2596,N_29178,N_29431);
nand UO_2597 (O_2597,N_29797,N_29112);
nor UO_2598 (O_2598,N_29032,N_29588);
or UO_2599 (O_2599,N_29830,N_29711);
xnor UO_2600 (O_2600,N_29228,N_29708);
xor UO_2601 (O_2601,N_29771,N_29616);
xnor UO_2602 (O_2602,N_29154,N_29732);
and UO_2603 (O_2603,N_29469,N_29668);
nor UO_2604 (O_2604,N_29432,N_29737);
or UO_2605 (O_2605,N_29612,N_29063);
or UO_2606 (O_2606,N_29174,N_29263);
or UO_2607 (O_2607,N_29565,N_29852);
nor UO_2608 (O_2608,N_29947,N_29251);
and UO_2609 (O_2609,N_29850,N_29615);
nand UO_2610 (O_2610,N_29587,N_29855);
and UO_2611 (O_2611,N_29276,N_29770);
and UO_2612 (O_2612,N_29351,N_29258);
and UO_2613 (O_2613,N_29402,N_29168);
or UO_2614 (O_2614,N_29158,N_29899);
or UO_2615 (O_2615,N_29912,N_29941);
and UO_2616 (O_2616,N_29104,N_29727);
and UO_2617 (O_2617,N_29029,N_29380);
and UO_2618 (O_2618,N_29799,N_29682);
nor UO_2619 (O_2619,N_29306,N_29966);
and UO_2620 (O_2620,N_29009,N_29968);
xor UO_2621 (O_2621,N_29256,N_29753);
and UO_2622 (O_2622,N_29231,N_29873);
or UO_2623 (O_2623,N_29354,N_29619);
xor UO_2624 (O_2624,N_29941,N_29813);
or UO_2625 (O_2625,N_29040,N_29222);
nand UO_2626 (O_2626,N_29540,N_29982);
and UO_2627 (O_2627,N_29138,N_29218);
nor UO_2628 (O_2628,N_29723,N_29014);
and UO_2629 (O_2629,N_29553,N_29452);
and UO_2630 (O_2630,N_29881,N_29915);
xnor UO_2631 (O_2631,N_29178,N_29450);
xnor UO_2632 (O_2632,N_29576,N_29060);
or UO_2633 (O_2633,N_29874,N_29892);
nor UO_2634 (O_2634,N_29434,N_29024);
xor UO_2635 (O_2635,N_29235,N_29952);
and UO_2636 (O_2636,N_29355,N_29981);
nand UO_2637 (O_2637,N_29130,N_29414);
xnor UO_2638 (O_2638,N_29344,N_29803);
xnor UO_2639 (O_2639,N_29872,N_29996);
nor UO_2640 (O_2640,N_29895,N_29688);
and UO_2641 (O_2641,N_29800,N_29838);
nor UO_2642 (O_2642,N_29471,N_29462);
nand UO_2643 (O_2643,N_29108,N_29668);
or UO_2644 (O_2644,N_29556,N_29303);
nand UO_2645 (O_2645,N_29930,N_29108);
nor UO_2646 (O_2646,N_29808,N_29201);
and UO_2647 (O_2647,N_29222,N_29929);
nor UO_2648 (O_2648,N_29003,N_29996);
nand UO_2649 (O_2649,N_29174,N_29952);
and UO_2650 (O_2650,N_29706,N_29048);
and UO_2651 (O_2651,N_29314,N_29847);
or UO_2652 (O_2652,N_29022,N_29879);
and UO_2653 (O_2653,N_29073,N_29103);
xor UO_2654 (O_2654,N_29455,N_29114);
or UO_2655 (O_2655,N_29388,N_29840);
nor UO_2656 (O_2656,N_29289,N_29850);
xor UO_2657 (O_2657,N_29945,N_29996);
and UO_2658 (O_2658,N_29785,N_29043);
and UO_2659 (O_2659,N_29415,N_29424);
nand UO_2660 (O_2660,N_29649,N_29500);
nor UO_2661 (O_2661,N_29978,N_29019);
xor UO_2662 (O_2662,N_29338,N_29009);
xnor UO_2663 (O_2663,N_29388,N_29544);
nor UO_2664 (O_2664,N_29591,N_29880);
nor UO_2665 (O_2665,N_29077,N_29942);
nor UO_2666 (O_2666,N_29498,N_29203);
or UO_2667 (O_2667,N_29834,N_29373);
and UO_2668 (O_2668,N_29580,N_29730);
xor UO_2669 (O_2669,N_29865,N_29113);
or UO_2670 (O_2670,N_29796,N_29194);
and UO_2671 (O_2671,N_29568,N_29530);
xor UO_2672 (O_2672,N_29845,N_29206);
and UO_2673 (O_2673,N_29528,N_29358);
xnor UO_2674 (O_2674,N_29992,N_29502);
and UO_2675 (O_2675,N_29079,N_29268);
xor UO_2676 (O_2676,N_29311,N_29229);
xor UO_2677 (O_2677,N_29681,N_29025);
xnor UO_2678 (O_2678,N_29241,N_29428);
nor UO_2679 (O_2679,N_29613,N_29419);
nor UO_2680 (O_2680,N_29843,N_29448);
and UO_2681 (O_2681,N_29642,N_29926);
nor UO_2682 (O_2682,N_29711,N_29765);
and UO_2683 (O_2683,N_29975,N_29154);
nor UO_2684 (O_2684,N_29311,N_29089);
nor UO_2685 (O_2685,N_29150,N_29117);
nor UO_2686 (O_2686,N_29087,N_29194);
or UO_2687 (O_2687,N_29990,N_29333);
and UO_2688 (O_2688,N_29401,N_29226);
nor UO_2689 (O_2689,N_29204,N_29304);
nand UO_2690 (O_2690,N_29690,N_29598);
nand UO_2691 (O_2691,N_29970,N_29436);
xor UO_2692 (O_2692,N_29703,N_29225);
nand UO_2693 (O_2693,N_29413,N_29330);
xnor UO_2694 (O_2694,N_29814,N_29950);
and UO_2695 (O_2695,N_29144,N_29546);
or UO_2696 (O_2696,N_29662,N_29792);
nor UO_2697 (O_2697,N_29553,N_29015);
nor UO_2698 (O_2698,N_29572,N_29319);
nand UO_2699 (O_2699,N_29351,N_29641);
and UO_2700 (O_2700,N_29228,N_29813);
nor UO_2701 (O_2701,N_29682,N_29992);
nor UO_2702 (O_2702,N_29691,N_29020);
xor UO_2703 (O_2703,N_29427,N_29846);
or UO_2704 (O_2704,N_29219,N_29716);
xnor UO_2705 (O_2705,N_29002,N_29418);
nand UO_2706 (O_2706,N_29726,N_29370);
and UO_2707 (O_2707,N_29586,N_29729);
and UO_2708 (O_2708,N_29121,N_29165);
nand UO_2709 (O_2709,N_29815,N_29913);
nor UO_2710 (O_2710,N_29878,N_29350);
and UO_2711 (O_2711,N_29973,N_29861);
and UO_2712 (O_2712,N_29296,N_29614);
nand UO_2713 (O_2713,N_29082,N_29540);
or UO_2714 (O_2714,N_29861,N_29986);
and UO_2715 (O_2715,N_29482,N_29899);
nand UO_2716 (O_2716,N_29884,N_29532);
xor UO_2717 (O_2717,N_29900,N_29981);
or UO_2718 (O_2718,N_29060,N_29172);
and UO_2719 (O_2719,N_29258,N_29237);
nor UO_2720 (O_2720,N_29871,N_29709);
nand UO_2721 (O_2721,N_29287,N_29541);
nor UO_2722 (O_2722,N_29836,N_29327);
nor UO_2723 (O_2723,N_29857,N_29455);
nor UO_2724 (O_2724,N_29329,N_29006);
nor UO_2725 (O_2725,N_29852,N_29552);
or UO_2726 (O_2726,N_29982,N_29944);
xor UO_2727 (O_2727,N_29368,N_29610);
nor UO_2728 (O_2728,N_29608,N_29414);
nor UO_2729 (O_2729,N_29334,N_29616);
and UO_2730 (O_2730,N_29393,N_29803);
nor UO_2731 (O_2731,N_29734,N_29286);
nand UO_2732 (O_2732,N_29746,N_29808);
and UO_2733 (O_2733,N_29679,N_29458);
and UO_2734 (O_2734,N_29391,N_29202);
xor UO_2735 (O_2735,N_29798,N_29378);
or UO_2736 (O_2736,N_29538,N_29024);
nor UO_2737 (O_2737,N_29332,N_29204);
xor UO_2738 (O_2738,N_29921,N_29258);
or UO_2739 (O_2739,N_29174,N_29721);
or UO_2740 (O_2740,N_29782,N_29684);
and UO_2741 (O_2741,N_29585,N_29214);
nand UO_2742 (O_2742,N_29733,N_29934);
nor UO_2743 (O_2743,N_29274,N_29116);
nor UO_2744 (O_2744,N_29057,N_29143);
nand UO_2745 (O_2745,N_29334,N_29722);
or UO_2746 (O_2746,N_29999,N_29946);
nand UO_2747 (O_2747,N_29854,N_29500);
and UO_2748 (O_2748,N_29467,N_29459);
and UO_2749 (O_2749,N_29344,N_29302);
nand UO_2750 (O_2750,N_29743,N_29400);
or UO_2751 (O_2751,N_29704,N_29958);
nand UO_2752 (O_2752,N_29548,N_29291);
nor UO_2753 (O_2753,N_29447,N_29027);
and UO_2754 (O_2754,N_29914,N_29598);
and UO_2755 (O_2755,N_29544,N_29796);
or UO_2756 (O_2756,N_29863,N_29461);
or UO_2757 (O_2757,N_29865,N_29990);
nor UO_2758 (O_2758,N_29877,N_29476);
nand UO_2759 (O_2759,N_29196,N_29610);
and UO_2760 (O_2760,N_29266,N_29973);
xnor UO_2761 (O_2761,N_29702,N_29643);
and UO_2762 (O_2762,N_29215,N_29211);
nand UO_2763 (O_2763,N_29493,N_29433);
or UO_2764 (O_2764,N_29971,N_29974);
nor UO_2765 (O_2765,N_29729,N_29165);
or UO_2766 (O_2766,N_29693,N_29315);
or UO_2767 (O_2767,N_29418,N_29645);
xnor UO_2768 (O_2768,N_29413,N_29169);
and UO_2769 (O_2769,N_29038,N_29818);
nor UO_2770 (O_2770,N_29089,N_29419);
nor UO_2771 (O_2771,N_29484,N_29305);
nand UO_2772 (O_2772,N_29613,N_29748);
and UO_2773 (O_2773,N_29276,N_29766);
nand UO_2774 (O_2774,N_29682,N_29183);
nor UO_2775 (O_2775,N_29611,N_29600);
nor UO_2776 (O_2776,N_29639,N_29336);
xnor UO_2777 (O_2777,N_29761,N_29633);
and UO_2778 (O_2778,N_29750,N_29042);
nand UO_2779 (O_2779,N_29915,N_29937);
xor UO_2780 (O_2780,N_29274,N_29866);
nor UO_2781 (O_2781,N_29604,N_29095);
nor UO_2782 (O_2782,N_29908,N_29654);
or UO_2783 (O_2783,N_29899,N_29403);
and UO_2784 (O_2784,N_29700,N_29351);
nand UO_2785 (O_2785,N_29062,N_29322);
nand UO_2786 (O_2786,N_29484,N_29837);
xnor UO_2787 (O_2787,N_29564,N_29880);
nor UO_2788 (O_2788,N_29087,N_29039);
nand UO_2789 (O_2789,N_29863,N_29343);
xnor UO_2790 (O_2790,N_29427,N_29129);
or UO_2791 (O_2791,N_29659,N_29318);
nor UO_2792 (O_2792,N_29816,N_29024);
and UO_2793 (O_2793,N_29491,N_29567);
or UO_2794 (O_2794,N_29015,N_29653);
nor UO_2795 (O_2795,N_29691,N_29525);
or UO_2796 (O_2796,N_29421,N_29004);
nand UO_2797 (O_2797,N_29826,N_29764);
nor UO_2798 (O_2798,N_29754,N_29551);
xnor UO_2799 (O_2799,N_29037,N_29826);
nand UO_2800 (O_2800,N_29709,N_29789);
and UO_2801 (O_2801,N_29305,N_29091);
nor UO_2802 (O_2802,N_29461,N_29931);
and UO_2803 (O_2803,N_29829,N_29303);
xor UO_2804 (O_2804,N_29549,N_29303);
xnor UO_2805 (O_2805,N_29229,N_29526);
nor UO_2806 (O_2806,N_29749,N_29666);
or UO_2807 (O_2807,N_29561,N_29242);
xor UO_2808 (O_2808,N_29747,N_29870);
xor UO_2809 (O_2809,N_29598,N_29145);
and UO_2810 (O_2810,N_29459,N_29187);
or UO_2811 (O_2811,N_29800,N_29482);
nand UO_2812 (O_2812,N_29670,N_29784);
xnor UO_2813 (O_2813,N_29491,N_29784);
and UO_2814 (O_2814,N_29180,N_29220);
nor UO_2815 (O_2815,N_29808,N_29357);
nor UO_2816 (O_2816,N_29709,N_29842);
or UO_2817 (O_2817,N_29989,N_29732);
nand UO_2818 (O_2818,N_29501,N_29206);
xor UO_2819 (O_2819,N_29490,N_29939);
xnor UO_2820 (O_2820,N_29221,N_29102);
or UO_2821 (O_2821,N_29560,N_29688);
nor UO_2822 (O_2822,N_29750,N_29096);
or UO_2823 (O_2823,N_29943,N_29796);
nor UO_2824 (O_2824,N_29603,N_29181);
nor UO_2825 (O_2825,N_29400,N_29705);
nand UO_2826 (O_2826,N_29831,N_29661);
nand UO_2827 (O_2827,N_29014,N_29113);
or UO_2828 (O_2828,N_29939,N_29380);
and UO_2829 (O_2829,N_29409,N_29176);
nand UO_2830 (O_2830,N_29727,N_29844);
nand UO_2831 (O_2831,N_29120,N_29692);
nor UO_2832 (O_2832,N_29871,N_29402);
nor UO_2833 (O_2833,N_29164,N_29829);
and UO_2834 (O_2834,N_29580,N_29362);
nand UO_2835 (O_2835,N_29998,N_29019);
or UO_2836 (O_2836,N_29490,N_29408);
or UO_2837 (O_2837,N_29693,N_29904);
nor UO_2838 (O_2838,N_29336,N_29119);
xor UO_2839 (O_2839,N_29094,N_29475);
xor UO_2840 (O_2840,N_29302,N_29026);
nor UO_2841 (O_2841,N_29166,N_29308);
or UO_2842 (O_2842,N_29862,N_29185);
nor UO_2843 (O_2843,N_29614,N_29604);
xnor UO_2844 (O_2844,N_29411,N_29892);
nor UO_2845 (O_2845,N_29652,N_29909);
xnor UO_2846 (O_2846,N_29134,N_29731);
xnor UO_2847 (O_2847,N_29580,N_29693);
nand UO_2848 (O_2848,N_29190,N_29874);
nor UO_2849 (O_2849,N_29477,N_29015);
or UO_2850 (O_2850,N_29543,N_29998);
nor UO_2851 (O_2851,N_29029,N_29736);
or UO_2852 (O_2852,N_29440,N_29648);
nor UO_2853 (O_2853,N_29911,N_29216);
or UO_2854 (O_2854,N_29197,N_29096);
or UO_2855 (O_2855,N_29938,N_29523);
and UO_2856 (O_2856,N_29538,N_29659);
and UO_2857 (O_2857,N_29061,N_29004);
xor UO_2858 (O_2858,N_29281,N_29803);
or UO_2859 (O_2859,N_29755,N_29265);
xnor UO_2860 (O_2860,N_29125,N_29419);
xor UO_2861 (O_2861,N_29635,N_29792);
nand UO_2862 (O_2862,N_29450,N_29211);
nor UO_2863 (O_2863,N_29812,N_29480);
or UO_2864 (O_2864,N_29880,N_29202);
nand UO_2865 (O_2865,N_29080,N_29603);
nand UO_2866 (O_2866,N_29531,N_29569);
nor UO_2867 (O_2867,N_29249,N_29620);
nand UO_2868 (O_2868,N_29772,N_29482);
nor UO_2869 (O_2869,N_29243,N_29631);
nor UO_2870 (O_2870,N_29930,N_29199);
and UO_2871 (O_2871,N_29770,N_29399);
or UO_2872 (O_2872,N_29243,N_29370);
or UO_2873 (O_2873,N_29928,N_29453);
and UO_2874 (O_2874,N_29895,N_29690);
xor UO_2875 (O_2875,N_29755,N_29699);
nor UO_2876 (O_2876,N_29889,N_29761);
and UO_2877 (O_2877,N_29041,N_29285);
xor UO_2878 (O_2878,N_29336,N_29697);
nor UO_2879 (O_2879,N_29741,N_29352);
xor UO_2880 (O_2880,N_29188,N_29251);
nor UO_2881 (O_2881,N_29399,N_29543);
nor UO_2882 (O_2882,N_29081,N_29039);
nor UO_2883 (O_2883,N_29000,N_29522);
nor UO_2884 (O_2884,N_29810,N_29128);
and UO_2885 (O_2885,N_29777,N_29006);
xor UO_2886 (O_2886,N_29014,N_29685);
xnor UO_2887 (O_2887,N_29049,N_29934);
nor UO_2888 (O_2888,N_29959,N_29985);
nor UO_2889 (O_2889,N_29708,N_29015);
xnor UO_2890 (O_2890,N_29200,N_29487);
nand UO_2891 (O_2891,N_29284,N_29405);
nand UO_2892 (O_2892,N_29466,N_29169);
nor UO_2893 (O_2893,N_29846,N_29050);
or UO_2894 (O_2894,N_29948,N_29773);
or UO_2895 (O_2895,N_29094,N_29912);
and UO_2896 (O_2896,N_29732,N_29150);
or UO_2897 (O_2897,N_29928,N_29689);
nor UO_2898 (O_2898,N_29006,N_29494);
xnor UO_2899 (O_2899,N_29197,N_29712);
or UO_2900 (O_2900,N_29225,N_29665);
xor UO_2901 (O_2901,N_29780,N_29830);
or UO_2902 (O_2902,N_29300,N_29764);
and UO_2903 (O_2903,N_29307,N_29490);
xor UO_2904 (O_2904,N_29383,N_29222);
nand UO_2905 (O_2905,N_29667,N_29038);
nand UO_2906 (O_2906,N_29312,N_29792);
and UO_2907 (O_2907,N_29631,N_29980);
nand UO_2908 (O_2908,N_29344,N_29026);
xnor UO_2909 (O_2909,N_29869,N_29229);
nor UO_2910 (O_2910,N_29013,N_29773);
nand UO_2911 (O_2911,N_29635,N_29860);
and UO_2912 (O_2912,N_29282,N_29924);
and UO_2913 (O_2913,N_29421,N_29193);
or UO_2914 (O_2914,N_29505,N_29333);
nand UO_2915 (O_2915,N_29276,N_29280);
and UO_2916 (O_2916,N_29012,N_29193);
xnor UO_2917 (O_2917,N_29615,N_29018);
nand UO_2918 (O_2918,N_29069,N_29115);
nand UO_2919 (O_2919,N_29992,N_29915);
or UO_2920 (O_2920,N_29199,N_29824);
or UO_2921 (O_2921,N_29357,N_29716);
xor UO_2922 (O_2922,N_29066,N_29299);
and UO_2923 (O_2923,N_29039,N_29839);
xor UO_2924 (O_2924,N_29272,N_29284);
or UO_2925 (O_2925,N_29882,N_29566);
nand UO_2926 (O_2926,N_29617,N_29446);
nand UO_2927 (O_2927,N_29490,N_29724);
nand UO_2928 (O_2928,N_29172,N_29078);
nor UO_2929 (O_2929,N_29681,N_29088);
nor UO_2930 (O_2930,N_29927,N_29988);
or UO_2931 (O_2931,N_29424,N_29964);
xnor UO_2932 (O_2932,N_29792,N_29995);
nor UO_2933 (O_2933,N_29610,N_29596);
nand UO_2934 (O_2934,N_29479,N_29070);
or UO_2935 (O_2935,N_29098,N_29186);
or UO_2936 (O_2936,N_29141,N_29183);
nand UO_2937 (O_2937,N_29531,N_29964);
nand UO_2938 (O_2938,N_29115,N_29925);
and UO_2939 (O_2939,N_29584,N_29932);
xor UO_2940 (O_2940,N_29907,N_29491);
nor UO_2941 (O_2941,N_29868,N_29974);
or UO_2942 (O_2942,N_29093,N_29459);
or UO_2943 (O_2943,N_29963,N_29121);
and UO_2944 (O_2944,N_29158,N_29507);
or UO_2945 (O_2945,N_29261,N_29318);
or UO_2946 (O_2946,N_29402,N_29031);
nor UO_2947 (O_2947,N_29889,N_29525);
nor UO_2948 (O_2948,N_29896,N_29907);
nand UO_2949 (O_2949,N_29078,N_29565);
or UO_2950 (O_2950,N_29730,N_29018);
and UO_2951 (O_2951,N_29809,N_29088);
or UO_2952 (O_2952,N_29724,N_29219);
and UO_2953 (O_2953,N_29503,N_29728);
xnor UO_2954 (O_2954,N_29749,N_29393);
or UO_2955 (O_2955,N_29182,N_29380);
nand UO_2956 (O_2956,N_29632,N_29908);
nand UO_2957 (O_2957,N_29127,N_29619);
and UO_2958 (O_2958,N_29840,N_29354);
nor UO_2959 (O_2959,N_29626,N_29579);
and UO_2960 (O_2960,N_29526,N_29979);
nand UO_2961 (O_2961,N_29297,N_29239);
or UO_2962 (O_2962,N_29597,N_29062);
and UO_2963 (O_2963,N_29798,N_29624);
nand UO_2964 (O_2964,N_29211,N_29192);
or UO_2965 (O_2965,N_29623,N_29098);
nor UO_2966 (O_2966,N_29771,N_29010);
nor UO_2967 (O_2967,N_29809,N_29089);
nor UO_2968 (O_2968,N_29329,N_29873);
xnor UO_2969 (O_2969,N_29288,N_29721);
xor UO_2970 (O_2970,N_29467,N_29220);
nor UO_2971 (O_2971,N_29844,N_29204);
xor UO_2972 (O_2972,N_29246,N_29748);
nand UO_2973 (O_2973,N_29594,N_29958);
or UO_2974 (O_2974,N_29631,N_29808);
or UO_2975 (O_2975,N_29633,N_29284);
xor UO_2976 (O_2976,N_29201,N_29056);
or UO_2977 (O_2977,N_29905,N_29099);
nand UO_2978 (O_2978,N_29580,N_29948);
xor UO_2979 (O_2979,N_29430,N_29330);
and UO_2980 (O_2980,N_29468,N_29310);
and UO_2981 (O_2981,N_29654,N_29299);
or UO_2982 (O_2982,N_29464,N_29260);
or UO_2983 (O_2983,N_29296,N_29572);
nor UO_2984 (O_2984,N_29509,N_29691);
xor UO_2985 (O_2985,N_29860,N_29760);
nand UO_2986 (O_2986,N_29558,N_29058);
nor UO_2987 (O_2987,N_29995,N_29506);
xor UO_2988 (O_2988,N_29065,N_29538);
or UO_2989 (O_2989,N_29156,N_29395);
or UO_2990 (O_2990,N_29599,N_29562);
and UO_2991 (O_2991,N_29412,N_29248);
xor UO_2992 (O_2992,N_29726,N_29059);
or UO_2993 (O_2993,N_29570,N_29120);
or UO_2994 (O_2994,N_29284,N_29354);
and UO_2995 (O_2995,N_29560,N_29540);
and UO_2996 (O_2996,N_29079,N_29552);
and UO_2997 (O_2997,N_29906,N_29537);
and UO_2998 (O_2998,N_29584,N_29913);
and UO_2999 (O_2999,N_29875,N_29204);
nand UO_3000 (O_3000,N_29514,N_29976);
and UO_3001 (O_3001,N_29239,N_29961);
nor UO_3002 (O_3002,N_29480,N_29555);
nand UO_3003 (O_3003,N_29115,N_29577);
xor UO_3004 (O_3004,N_29958,N_29645);
xnor UO_3005 (O_3005,N_29300,N_29860);
nand UO_3006 (O_3006,N_29981,N_29718);
nand UO_3007 (O_3007,N_29427,N_29900);
and UO_3008 (O_3008,N_29457,N_29603);
or UO_3009 (O_3009,N_29087,N_29945);
xnor UO_3010 (O_3010,N_29741,N_29200);
nor UO_3011 (O_3011,N_29812,N_29624);
nand UO_3012 (O_3012,N_29281,N_29030);
nor UO_3013 (O_3013,N_29319,N_29606);
xnor UO_3014 (O_3014,N_29815,N_29342);
and UO_3015 (O_3015,N_29894,N_29088);
xor UO_3016 (O_3016,N_29623,N_29336);
nand UO_3017 (O_3017,N_29727,N_29499);
xor UO_3018 (O_3018,N_29649,N_29758);
nand UO_3019 (O_3019,N_29047,N_29169);
xor UO_3020 (O_3020,N_29823,N_29040);
xnor UO_3021 (O_3021,N_29148,N_29479);
xor UO_3022 (O_3022,N_29475,N_29674);
nand UO_3023 (O_3023,N_29640,N_29652);
nand UO_3024 (O_3024,N_29025,N_29084);
nand UO_3025 (O_3025,N_29825,N_29332);
nand UO_3026 (O_3026,N_29323,N_29220);
or UO_3027 (O_3027,N_29865,N_29038);
or UO_3028 (O_3028,N_29973,N_29410);
nand UO_3029 (O_3029,N_29043,N_29473);
xor UO_3030 (O_3030,N_29963,N_29776);
xor UO_3031 (O_3031,N_29112,N_29815);
nand UO_3032 (O_3032,N_29052,N_29982);
or UO_3033 (O_3033,N_29148,N_29451);
or UO_3034 (O_3034,N_29117,N_29439);
or UO_3035 (O_3035,N_29951,N_29531);
xnor UO_3036 (O_3036,N_29034,N_29966);
and UO_3037 (O_3037,N_29234,N_29696);
nor UO_3038 (O_3038,N_29219,N_29855);
or UO_3039 (O_3039,N_29175,N_29946);
nand UO_3040 (O_3040,N_29236,N_29635);
nor UO_3041 (O_3041,N_29793,N_29548);
or UO_3042 (O_3042,N_29483,N_29247);
nand UO_3043 (O_3043,N_29237,N_29996);
nand UO_3044 (O_3044,N_29723,N_29159);
nand UO_3045 (O_3045,N_29192,N_29605);
and UO_3046 (O_3046,N_29017,N_29200);
nor UO_3047 (O_3047,N_29606,N_29795);
nand UO_3048 (O_3048,N_29576,N_29967);
and UO_3049 (O_3049,N_29824,N_29518);
xnor UO_3050 (O_3050,N_29010,N_29054);
nor UO_3051 (O_3051,N_29243,N_29809);
xor UO_3052 (O_3052,N_29256,N_29748);
or UO_3053 (O_3053,N_29466,N_29489);
xor UO_3054 (O_3054,N_29052,N_29103);
xor UO_3055 (O_3055,N_29682,N_29808);
or UO_3056 (O_3056,N_29590,N_29144);
nand UO_3057 (O_3057,N_29687,N_29346);
nor UO_3058 (O_3058,N_29772,N_29672);
nand UO_3059 (O_3059,N_29492,N_29878);
nor UO_3060 (O_3060,N_29069,N_29417);
nand UO_3061 (O_3061,N_29432,N_29578);
nand UO_3062 (O_3062,N_29187,N_29099);
nand UO_3063 (O_3063,N_29103,N_29098);
and UO_3064 (O_3064,N_29368,N_29757);
xor UO_3065 (O_3065,N_29706,N_29944);
nor UO_3066 (O_3066,N_29122,N_29062);
xor UO_3067 (O_3067,N_29635,N_29595);
nor UO_3068 (O_3068,N_29130,N_29264);
xor UO_3069 (O_3069,N_29570,N_29176);
nand UO_3070 (O_3070,N_29753,N_29270);
nand UO_3071 (O_3071,N_29051,N_29989);
or UO_3072 (O_3072,N_29568,N_29861);
nor UO_3073 (O_3073,N_29429,N_29166);
nand UO_3074 (O_3074,N_29961,N_29778);
and UO_3075 (O_3075,N_29062,N_29427);
xor UO_3076 (O_3076,N_29411,N_29681);
or UO_3077 (O_3077,N_29539,N_29239);
nand UO_3078 (O_3078,N_29234,N_29743);
and UO_3079 (O_3079,N_29063,N_29129);
nand UO_3080 (O_3080,N_29884,N_29232);
nand UO_3081 (O_3081,N_29362,N_29620);
nor UO_3082 (O_3082,N_29768,N_29697);
or UO_3083 (O_3083,N_29874,N_29117);
xnor UO_3084 (O_3084,N_29073,N_29925);
xnor UO_3085 (O_3085,N_29965,N_29244);
nand UO_3086 (O_3086,N_29854,N_29747);
xor UO_3087 (O_3087,N_29892,N_29018);
or UO_3088 (O_3088,N_29967,N_29668);
nor UO_3089 (O_3089,N_29569,N_29694);
nor UO_3090 (O_3090,N_29653,N_29157);
xor UO_3091 (O_3091,N_29963,N_29712);
nand UO_3092 (O_3092,N_29696,N_29994);
xnor UO_3093 (O_3093,N_29757,N_29900);
nand UO_3094 (O_3094,N_29094,N_29587);
nand UO_3095 (O_3095,N_29382,N_29336);
nor UO_3096 (O_3096,N_29711,N_29586);
nand UO_3097 (O_3097,N_29545,N_29994);
xnor UO_3098 (O_3098,N_29193,N_29574);
or UO_3099 (O_3099,N_29086,N_29517);
xnor UO_3100 (O_3100,N_29550,N_29946);
nand UO_3101 (O_3101,N_29696,N_29552);
xnor UO_3102 (O_3102,N_29715,N_29487);
nor UO_3103 (O_3103,N_29419,N_29537);
and UO_3104 (O_3104,N_29428,N_29407);
xor UO_3105 (O_3105,N_29862,N_29577);
or UO_3106 (O_3106,N_29115,N_29755);
nor UO_3107 (O_3107,N_29459,N_29214);
nand UO_3108 (O_3108,N_29209,N_29202);
and UO_3109 (O_3109,N_29482,N_29018);
or UO_3110 (O_3110,N_29131,N_29976);
nor UO_3111 (O_3111,N_29058,N_29740);
nand UO_3112 (O_3112,N_29982,N_29189);
nand UO_3113 (O_3113,N_29518,N_29613);
nor UO_3114 (O_3114,N_29748,N_29679);
or UO_3115 (O_3115,N_29058,N_29472);
and UO_3116 (O_3116,N_29134,N_29963);
xor UO_3117 (O_3117,N_29458,N_29931);
and UO_3118 (O_3118,N_29223,N_29692);
nand UO_3119 (O_3119,N_29064,N_29156);
or UO_3120 (O_3120,N_29080,N_29608);
xor UO_3121 (O_3121,N_29508,N_29960);
nor UO_3122 (O_3122,N_29750,N_29571);
or UO_3123 (O_3123,N_29794,N_29561);
and UO_3124 (O_3124,N_29375,N_29614);
and UO_3125 (O_3125,N_29899,N_29619);
and UO_3126 (O_3126,N_29013,N_29657);
and UO_3127 (O_3127,N_29200,N_29165);
xor UO_3128 (O_3128,N_29108,N_29604);
xor UO_3129 (O_3129,N_29974,N_29671);
and UO_3130 (O_3130,N_29991,N_29571);
or UO_3131 (O_3131,N_29587,N_29816);
or UO_3132 (O_3132,N_29994,N_29384);
nand UO_3133 (O_3133,N_29189,N_29136);
xor UO_3134 (O_3134,N_29649,N_29422);
xor UO_3135 (O_3135,N_29800,N_29921);
nor UO_3136 (O_3136,N_29405,N_29121);
or UO_3137 (O_3137,N_29632,N_29927);
or UO_3138 (O_3138,N_29510,N_29706);
nand UO_3139 (O_3139,N_29562,N_29032);
xor UO_3140 (O_3140,N_29930,N_29185);
nor UO_3141 (O_3141,N_29831,N_29192);
nor UO_3142 (O_3142,N_29265,N_29840);
and UO_3143 (O_3143,N_29813,N_29209);
nand UO_3144 (O_3144,N_29827,N_29420);
and UO_3145 (O_3145,N_29726,N_29100);
and UO_3146 (O_3146,N_29411,N_29725);
nand UO_3147 (O_3147,N_29234,N_29165);
xor UO_3148 (O_3148,N_29328,N_29077);
nand UO_3149 (O_3149,N_29781,N_29195);
or UO_3150 (O_3150,N_29638,N_29627);
xor UO_3151 (O_3151,N_29075,N_29168);
or UO_3152 (O_3152,N_29422,N_29811);
or UO_3153 (O_3153,N_29684,N_29408);
and UO_3154 (O_3154,N_29824,N_29929);
nor UO_3155 (O_3155,N_29593,N_29486);
nand UO_3156 (O_3156,N_29790,N_29157);
and UO_3157 (O_3157,N_29766,N_29196);
and UO_3158 (O_3158,N_29747,N_29783);
or UO_3159 (O_3159,N_29294,N_29951);
nand UO_3160 (O_3160,N_29001,N_29230);
and UO_3161 (O_3161,N_29837,N_29035);
and UO_3162 (O_3162,N_29022,N_29013);
nand UO_3163 (O_3163,N_29117,N_29121);
and UO_3164 (O_3164,N_29701,N_29028);
nor UO_3165 (O_3165,N_29889,N_29465);
and UO_3166 (O_3166,N_29646,N_29206);
nor UO_3167 (O_3167,N_29239,N_29061);
and UO_3168 (O_3168,N_29831,N_29505);
nor UO_3169 (O_3169,N_29777,N_29199);
nor UO_3170 (O_3170,N_29149,N_29047);
nor UO_3171 (O_3171,N_29666,N_29015);
nand UO_3172 (O_3172,N_29500,N_29893);
nor UO_3173 (O_3173,N_29003,N_29483);
nand UO_3174 (O_3174,N_29446,N_29922);
nand UO_3175 (O_3175,N_29467,N_29312);
and UO_3176 (O_3176,N_29264,N_29145);
or UO_3177 (O_3177,N_29612,N_29973);
nand UO_3178 (O_3178,N_29510,N_29242);
and UO_3179 (O_3179,N_29785,N_29559);
nand UO_3180 (O_3180,N_29467,N_29568);
or UO_3181 (O_3181,N_29347,N_29980);
or UO_3182 (O_3182,N_29636,N_29291);
or UO_3183 (O_3183,N_29908,N_29902);
or UO_3184 (O_3184,N_29276,N_29196);
xor UO_3185 (O_3185,N_29313,N_29442);
xor UO_3186 (O_3186,N_29538,N_29428);
nor UO_3187 (O_3187,N_29361,N_29000);
nor UO_3188 (O_3188,N_29320,N_29502);
nand UO_3189 (O_3189,N_29215,N_29105);
nand UO_3190 (O_3190,N_29325,N_29503);
xnor UO_3191 (O_3191,N_29877,N_29373);
nor UO_3192 (O_3192,N_29135,N_29920);
nand UO_3193 (O_3193,N_29650,N_29077);
nand UO_3194 (O_3194,N_29631,N_29164);
and UO_3195 (O_3195,N_29410,N_29461);
nor UO_3196 (O_3196,N_29414,N_29760);
and UO_3197 (O_3197,N_29795,N_29762);
xor UO_3198 (O_3198,N_29336,N_29888);
or UO_3199 (O_3199,N_29435,N_29346);
or UO_3200 (O_3200,N_29876,N_29668);
or UO_3201 (O_3201,N_29057,N_29261);
xor UO_3202 (O_3202,N_29530,N_29451);
nor UO_3203 (O_3203,N_29372,N_29135);
nor UO_3204 (O_3204,N_29915,N_29095);
xor UO_3205 (O_3205,N_29285,N_29053);
and UO_3206 (O_3206,N_29855,N_29267);
nor UO_3207 (O_3207,N_29237,N_29740);
and UO_3208 (O_3208,N_29036,N_29672);
and UO_3209 (O_3209,N_29859,N_29661);
xnor UO_3210 (O_3210,N_29000,N_29170);
nor UO_3211 (O_3211,N_29862,N_29257);
xnor UO_3212 (O_3212,N_29003,N_29771);
and UO_3213 (O_3213,N_29705,N_29667);
nand UO_3214 (O_3214,N_29896,N_29304);
nor UO_3215 (O_3215,N_29775,N_29492);
nand UO_3216 (O_3216,N_29496,N_29064);
or UO_3217 (O_3217,N_29018,N_29266);
or UO_3218 (O_3218,N_29520,N_29687);
and UO_3219 (O_3219,N_29323,N_29673);
or UO_3220 (O_3220,N_29213,N_29009);
or UO_3221 (O_3221,N_29179,N_29531);
xor UO_3222 (O_3222,N_29688,N_29641);
nand UO_3223 (O_3223,N_29334,N_29441);
xnor UO_3224 (O_3224,N_29249,N_29385);
or UO_3225 (O_3225,N_29338,N_29553);
nor UO_3226 (O_3226,N_29214,N_29119);
nand UO_3227 (O_3227,N_29135,N_29392);
nor UO_3228 (O_3228,N_29908,N_29440);
nand UO_3229 (O_3229,N_29191,N_29399);
nor UO_3230 (O_3230,N_29705,N_29148);
or UO_3231 (O_3231,N_29020,N_29731);
nor UO_3232 (O_3232,N_29233,N_29988);
or UO_3233 (O_3233,N_29143,N_29069);
nand UO_3234 (O_3234,N_29549,N_29852);
nor UO_3235 (O_3235,N_29123,N_29860);
and UO_3236 (O_3236,N_29969,N_29163);
or UO_3237 (O_3237,N_29579,N_29761);
nor UO_3238 (O_3238,N_29431,N_29093);
nor UO_3239 (O_3239,N_29594,N_29187);
and UO_3240 (O_3240,N_29636,N_29004);
xnor UO_3241 (O_3241,N_29447,N_29630);
nor UO_3242 (O_3242,N_29111,N_29898);
or UO_3243 (O_3243,N_29945,N_29093);
xnor UO_3244 (O_3244,N_29055,N_29927);
or UO_3245 (O_3245,N_29816,N_29521);
nor UO_3246 (O_3246,N_29957,N_29858);
xnor UO_3247 (O_3247,N_29648,N_29999);
nor UO_3248 (O_3248,N_29915,N_29614);
nor UO_3249 (O_3249,N_29388,N_29248);
and UO_3250 (O_3250,N_29867,N_29053);
xnor UO_3251 (O_3251,N_29246,N_29987);
nor UO_3252 (O_3252,N_29747,N_29737);
xnor UO_3253 (O_3253,N_29172,N_29066);
or UO_3254 (O_3254,N_29871,N_29192);
xor UO_3255 (O_3255,N_29636,N_29382);
nand UO_3256 (O_3256,N_29558,N_29630);
nand UO_3257 (O_3257,N_29671,N_29693);
xnor UO_3258 (O_3258,N_29894,N_29435);
and UO_3259 (O_3259,N_29440,N_29811);
nand UO_3260 (O_3260,N_29481,N_29237);
nand UO_3261 (O_3261,N_29869,N_29335);
or UO_3262 (O_3262,N_29360,N_29779);
xor UO_3263 (O_3263,N_29335,N_29749);
nand UO_3264 (O_3264,N_29196,N_29671);
or UO_3265 (O_3265,N_29178,N_29640);
and UO_3266 (O_3266,N_29040,N_29516);
or UO_3267 (O_3267,N_29089,N_29465);
and UO_3268 (O_3268,N_29413,N_29960);
xor UO_3269 (O_3269,N_29836,N_29397);
xnor UO_3270 (O_3270,N_29053,N_29447);
or UO_3271 (O_3271,N_29848,N_29460);
and UO_3272 (O_3272,N_29468,N_29664);
or UO_3273 (O_3273,N_29455,N_29120);
nand UO_3274 (O_3274,N_29896,N_29944);
or UO_3275 (O_3275,N_29576,N_29078);
or UO_3276 (O_3276,N_29809,N_29942);
or UO_3277 (O_3277,N_29431,N_29873);
or UO_3278 (O_3278,N_29717,N_29034);
or UO_3279 (O_3279,N_29180,N_29902);
nand UO_3280 (O_3280,N_29165,N_29908);
and UO_3281 (O_3281,N_29094,N_29677);
nor UO_3282 (O_3282,N_29757,N_29407);
nor UO_3283 (O_3283,N_29972,N_29786);
and UO_3284 (O_3284,N_29272,N_29968);
and UO_3285 (O_3285,N_29964,N_29045);
nor UO_3286 (O_3286,N_29223,N_29319);
nor UO_3287 (O_3287,N_29632,N_29484);
nand UO_3288 (O_3288,N_29930,N_29092);
and UO_3289 (O_3289,N_29739,N_29331);
nand UO_3290 (O_3290,N_29491,N_29627);
and UO_3291 (O_3291,N_29585,N_29577);
or UO_3292 (O_3292,N_29747,N_29015);
nand UO_3293 (O_3293,N_29209,N_29868);
and UO_3294 (O_3294,N_29198,N_29712);
nor UO_3295 (O_3295,N_29724,N_29757);
xor UO_3296 (O_3296,N_29781,N_29498);
and UO_3297 (O_3297,N_29941,N_29257);
xnor UO_3298 (O_3298,N_29452,N_29583);
xnor UO_3299 (O_3299,N_29490,N_29600);
nor UO_3300 (O_3300,N_29537,N_29164);
and UO_3301 (O_3301,N_29584,N_29314);
xnor UO_3302 (O_3302,N_29697,N_29784);
nand UO_3303 (O_3303,N_29696,N_29933);
and UO_3304 (O_3304,N_29481,N_29450);
and UO_3305 (O_3305,N_29524,N_29859);
nor UO_3306 (O_3306,N_29908,N_29213);
nor UO_3307 (O_3307,N_29256,N_29244);
xor UO_3308 (O_3308,N_29384,N_29833);
or UO_3309 (O_3309,N_29604,N_29000);
and UO_3310 (O_3310,N_29218,N_29945);
xnor UO_3311 (O_3311,N_29911,N_29928);
or UO_3312 (O_3312,N_29491,N_29231);
or UO_3313 (O_3313,N_29334,N_29864);
or UO_3314 (O_3314,N_29424,N_29627);
nand UO_3315 (O_3315,N_29128,N_29570);
nor UO_3316 (O_3316,N_29365,N_29796);
or UO_3317 (O_3317,N_29208,N_29943);
and UO_3318 (O_3318,N_29199,N_29779);
or UO_3319 (O_3319,N_29075,N_29761);
or UO_3320 (O_3320,N_29534,N_29551);
xor UO_3321 (O_3321,N_29168,N_29137);
or UO_3322 (O_3322,N_29006,N_29966);
and UO_3323 (O_3323,N_29142,N_29527);
nor UO_3324 (O_3324,N_29078,N_29055);
nand UO_3325 (O_3325,N_29030,N_29510);
or UO_3326 (O_3326,N_29607,N_29043);
and UO_3327 (O_3327,N_29315,N_29962);
nor UO_3328 (O_3328,N_29355,N_29220);
nand UO_3329 (O_3329,N_29984,N_29044);
and UO_3330 (O_3330,N_29743,N_29419);
and UO_3331 (O_3331,N_29125,N_29292);
and UO_3332 (O_3332,N_29202,N_29981);
nor UO_3333 (O_3333,N_29088,N_29741);
xnor UO_3334 (O_3334,N_29306,N_29518);
and UO_3335 (O_3335,N_29183,N_29122);
nor UO_3336 (O_3336,N_29090,N_29394);
nor UO_3337 (O_3337,N_29107,N_29318);
or UO_3338 (O_3338,N_29910,N_29956);
and UO_3339 (O_3339,N_29238,N_29703);
nand UO_3340 (O_3340,N_29614,N_29369);
or UO_3341 (O_3341,N_29964,N_29927);
nor UO_3342 (O_3342,N_29569,N_29424);
nand UO_3343 (O_3343,N_29171,N_29563);
nor UO_3344 (O_3344,N_29690,N_29015);
nor UO_3345 (O_3345,N_29845,N_29466);
xor UO_3346 (O_3346,N_29707,N_29990);
nand UO_3347 (O_3347,N_29035,N_29220);
xnor UO_3348 (O_3348,N_29553,N_29425);
nor UO_3349 (O_3349,N_29977,N_29358);
or UO_3350 (O_3350,N_29117,N_29811);
and UO_3351 (O_3351,N_29314,N_29578);
and UO_3352 (O_3352,N_29565,N_29806);
nand UO_3353 (O_3353,N_29382,N_29415);
nor UO_3354 (O_3354,N_29636,N_29251);
or UO_3355 (O_3355,N_29327,N_29432);
xor UO_3356 (O_3356,N_29595,N_29698);
or UO_3357 (O_3357,N_29907,N_29375);
nand UO_3358 (O_3358,N_29371,N_29074);
nor UO_3359 (O_3359,N_29957,N_29159);
or UO_3360 (O_3360,N_29305,N_29018);
nor UO_3361 (O_3361,N_29132,N_29099);
xor UO_3362 (O_3362,N_29174,N_29052);
and UO_3363 (O_3363,N_29262,N_29971);
and UO_3364 (O_3364,N_29121,N_29687);
or UO_3365 (O_3365,N_29328,N_29358);
xor UO_3366 (O_3366,N_29317,N_29420);
nand UO_3367 (O_3367,N_29733,N_29341);
and UO_3368 (O_3368,N_29848,N_29934);
xor UO_3369 (O_3369,N_29631,N_29526);
or UO_3370 (O_3370,N_29152,N_29210);
and UO_3371 (O_3371,N_29373,N_29163);
nand UO_3372 (O_3372,N_29125,N_29167);
nor UO_3373 (O_3373,N_29389,N_29329);
nand UO_3374 (O_3374,N_29814,N_29423);
or UO_3375 (O_3375,N_29358,N_29613);
xor UO_3376 (O_3376,N_29073,N_29954);
and UO_3377 (O_3377,N_29984,N_29164);
or UO_3378 (O_3378,N_29473,N_29942);
nand UO_3379 (O_3379,N_29075,N_29963);
or UO_3380 (O_3380,N_29153,N_29676);
or UO_3381 (O_3381,N_29875,N_29019);
nand UO_3382 (O_3382,N_29909,N_29963);
nor UO_3383 (O_3383,N_29393,N_29477);
or UO_3384 (O_3384,N_29760,N_29393);
and UO_3385 (O_3385,N_29171,N_29274);
nor UO_3386 (O_3386,N_29778,N_29735);
or UO_3387 (O_3387,N_29715,N_29933);
nand UO_3388 (O_3388,N_29459,N_29789);
nor UO_3389 (O_3389,N_29938,N_29182);
nand UO_3390 (O_3390,N_29939,N_29461);
xnor UO_3391 (O_3391,N_29850,N_29514);
xor UO_3392 (O_3392,N_29857,N_29750);
or UO_3393 (O_3393,N_29960,N_29554);
or UO_3394 (O_3394,N_29222,N_29467);
nand UO_3395 (O_3395,N_29800,N_29124);
or UO_3396 (O_3396,N_29860,N_29648);
nand UO_3397 (O_3397,N_29815,N_29155);
nor UO_3398 (O_3398,N_29792,N_29611);
and UO_3399 (O_3399,N_29169,N_29279);
nand UO_3400 (O_3400,N_29949,N_29102);
or UO_3401 (O_3401,N_29728,N_29378);
and UO_3402 (O_3402,N_29532,N_29073);
xor UO_3403 (O_3403,N_29250,N_29198);
nand UO_3404 (O_3404,N_29870,N_29115);
nor UO_3405 (O_3405,N_29832,N_29445);
nand UO_3406 (O_3406,N_29911,N_29423);
nor UO_3407 (O_3407,N_29973,N_29789);
or UO_3408 (O_3408,N_29019,N_29533);
nor UO_3409 (O_3409,N_29839,N_29781);
or UO_3410 (O_3410,N_29085,N_29023);
xor UO_3411 (O_3411,N_29224,N_29865);
nand UO_3412 (O_3412,N_29097,N_29551);
or UO_3413 (O_3413,N_29396,N_29674);
nor UO_3414 (O_3414,N_29883,N_29421);
or UO_3415 (O_3415,N_29583,N_29422);
nor UO_3416 (O_3416,N_29774,N_29106);
and UO_3417 (O_3417,N_29275,N_29968);
xnor UO_3418 (O_3418,N_29564,N_29720);
nor UO_3419 (O_3419,N_29458,N_29087);
and UO_3420 (O_3420,N_29372,N_29888);
or UO_3421 (O_3421,N_29878,N_29318);
xor UO_3422 (O_3422,N_29789,N_29264);
and UO_3423 (O_3423,N_29118,N_29244);
xnor UO_3424 (O_3424,N_29143,N_29247);
nor UO_3425 (O_3425,N_29303,N_29044);
or UO_3426 (O_3426,N_29707,N_29374);
or UO_3427 (O_3427,N_29548,N_29392);
xnor UO_3428 (O_3428,N_29698,N_29703);
nand UO_3429 (O_3429,N_29688,N_29357);
and UO_3430 (O_3430,N_29410,N_29055);
and UO_3431 (O_3431,N_29065,N_29423);
and UO_3432 (O_3432,N_29051,N_29078);
nor UO_3433 (O_3433,N_29601,N_29918);
and UO_3434 (O_3434,N_29239,N_29213);
or UO_3435 (O_3435,N_29465,N_29864);
nor UO_3436 (O_3436,N_29230,N_29694);
nand UO_3437 (O_3437,N_29860,N_29703);
nand UO_3438 (O_3438,N_29089,N_29547);
nor UO_3439 (O_3439,N_29520,N_29134);
xor UO_3440 (O_3440,N_29472,N_29906);
xor UO_3441 (O_3441,N_29742,N_29605);
and UO_3442 (O_3442,N_29004,N_29041);
and UO_3443 (O_3443,N_29386,N_29984);
nand UO_3444 (O_3444,N_29051,N_29474);
xor UO_3445 (O_3445,N_29689,N_29571);
xnor UO_3446 (O_3446,N_29126,N_29244);
and UO_3447 (O_3447,N_29616,N_29325);
or UO_3448 (O_3448,N_29110,N_29180);
or UO_3449 (O_3449,N_29641,N_29691);
xnor UO_3450 (O_3450,N_29385,N_29468);
or UO_3451 (O_3451,N_29935,N_29543);
or UO_3452 (O_3452,N_29021,N_29442);
xor UO_3453 (O_3453,N_29450,N_29673);
nor UO_3454 (O_3454,N_29308,N_29999);
or UO_3455 (O_3455,N_29573,N_29578);
nand UO_3456 (O_3456,N_29670,N_29773);
nor UO_3457 (O_3457,N_29934,N_29623);
or UO_3458 (O_3458,N_29228,N_29492);
xor UO_3459 (O_3459,N_29909,N_29102);
or UO_3460 (O_3460,N_29653,N_29728);
nor UO_3461 (O_3461,N_29375,N_29176);
xor UO_3462 (O_3462,N_29063,N_29269);
and UO_3463 (O_3463,N_29886,N_29783);
xnor UO_3464 (O_3464,N_29084,N_29660);
nor UO_3465 (O_3465,N_29156,N_29377);
and UO_3466 (O_3466,N_29373,N_29532);
and UO_3467 (O_3467,N_29652,N_29727);
or UO_3468 (O_3468,N_29667,N_29670);
or UO_3469 (O_3469,N_29827,N_29189);
nand UO_3470 (O_3470,N_29648,N_29872);
nand UO_3471 (O_3471,N_29275,N_29393);
nor UO_3472 (O_3472,N_29662,N_29809);
or UO_3473 (O_3473,N_29431,N_29988);
or UO_3474 (O_3474,N_29972,N_29454);
nand UO_3475 (O_3475,N_29883,N_29407);
and UO_3476 (O_3476,N_29178,N_29775);
nand UO_3477 (O_3477,N_29286,N_29363);
or UO_3478 (O_3478,N_29074,N_29576);
xnor UO_3479 (O_3479,N_29540,N_29095);
nand UO_3480 (O_3480,N_29339,N_29699);
nor UO_3481 (O_3481,N_29041,N_29981);
nor UO_3482 (O_3482,N_29481,N_29074);
or UO_3483 (O_3483,N_29863,N_29385);
and UO_3484 (O_3484,N_29077,N_29949);
and UO_3485 (O_3485,N_29071,N_29339);
xnor UO_3486 (O_3486,N_29904,N_29081);
and UO_3487 (O_3487,N_29594,N_29308);
nor UO_3488 (O_3488,N_29935,N_29270);
xor UO_3489 (O_3489,N_29919,N_29055);
xor UO_3490 (O_3490,N_29428,N_29503);
nor UO_3491 (O_3491,N_29080,N_29706);
nand UO_3492 (O_3492,N_29129,N_29389);
and UO_3493 (O_3493,N_29665,N_29054);
xnor UO_3494 (O_3494,N_29450,N_29073);
nor UO_3495 (O_3495,N_29500,N_29061);
or UO_3496 (O_3496,N_29831,N_29722);
xor UO_3497 (O_3497,N_29767,N_29557);
xnor UO_3498 (O_3498,N_29750,N_29749);
or UO_3499 (O_3499,N_29217,N_29849);
endmodule