module basic_1000_10000_1500_2_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5004,N_5005,N_5007,N_5009,N_5012,N_5014,N_5015,N_5016,N_5017,N_5021,N_5024,N_5025,N_5027,N_5028,N_5030,N_5031,N_5033,N_5034,N_5036,N_5037,N_5038,N_5039,N_5046,N_5047,N_5049,N_5051,N_5052,N_5054,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5063,N_5064,N_5065,N_5067,N_5068,N_5071,N_5072,N_5073,N_5075,N_5076,N_5078,N_5080,N_5081,N_5082,N_5083,N_5086,N_5088,N_5090,N_5091,N_5092,N_5093,N_5096,N_5097,N_5098,N_5099,N_5107,N_5108,N_5109,N_5111,N_5112,N_5116,N_5117,N_5119,N_5120,N_5121,N_5122,N_5124,N_5125,N_5126,N_5128,N_5130,N_5132,N_5133,N_5134,N_5135,N_5136,N_5138,N_5140,N_5141,N_5142,N_5143,N_5147,N_5151,N_5152,N_5154,N_5155,N_5158,N_5159,N_5160,N_5161,N_5163,N_5165,N_5169,N_5170,N_5171,N_5172,N_5174,N_5175,N_5176,N_5177,N_5178,N_5181,N_5182,N_5183,N_5184,N_5186,N_5187,N_5188,N_5193,N_5194,N_5195,N_5197,N_5198,N_5199,N_5200,N_5201,N_5203,N_5204,N_5205,N_5206,N_5207,N_5209,N_5212,N_5214,N_5216,N_5217,N_5218,N_5220,N_5222,N_5225,N_5229,N_5231,N_5234,N_5235,N_5236,N_5239,N_5240,N_5241,N_5243,N_5244,N_5251,N_5252,N_5253,N_5254,N_5257,N_5259,N_5261,N_5262,N_5263,N_5265,N_5267,N_5270,N_5271,N_5272,N_5273,N_5274,N_5278,N_5279,N_5280,N_5281,N_5282,N_5286,N_5288,N_5289,N_5290,N_5292,N_5295,N_5296,N_5299,N_5300,N_5303,N_5305,N_5306,N_5307,N_5308,N_5310,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5335,N_5337,N_5338,N_5341,N_5342,N_5343,N_5345,N_5346,N_5347,N_5348,N_5349,N_5353,N_5355,N_5358,N_5359,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5368,N_5369,N_5371,N_5373,N_5375,N_5377,N_5379,N_5380,N_5381,N_5384,N_5385,N_5386,N_5387,N_5388,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5402,N_5403,N_5405,N_5406,N_5411,N_5414,N_5416,N_5418,N_5419,N_5422,N_5424,N_5426,N_5427,N_5428,N_5431,N_5433,N_5434,N_5437,N_5438,N_5439,N_5441,N_5442,N_5443,N_5446,N_5447,N_5449,N_5450,N_5451,N_5453,N_5455,N_5456,N_5457,N_5458,N_5463,N_5464,N_5465,N_5466,N_5472,N_5476,N_5477,N_5478,N_5479,N_5480,N_5483,N_5485,N_5487,N_5489,N_5490,N_5492,N_5493,N_5494,N_5495,N_5498,N_5499,N_5500,N_5505,N_5506,N_5508,N_5510,N_5511,N_5512,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5526,N_5527,N_5528,N_5529,N_5532,N_5533,N_5534,N_5535,N_5536,N_5538,N_5539,N_5540,N_5543,N_5544,N_5545,N_5551,N_5552,N_5555,N_5556,N_5557,N_5558,N_5560,N_5561,N_5563,N_5566,N_5567,N_5568,N_5570,N_5571,N_5572,N_5574,N_5575,N_5577,N_5583,N_5584,N_5587,N_5588,N_5590,N_5591,N_5592,N_5594,N_5596,N_5597,N_5601,N_5602,N_5604,N_5606,N_5607,N_5609,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5621,N_5622,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5634,N_5635,N_5636,N_5638,N_5640,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5651,N_5652,N_5655,N_5658,N_5660,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5671,N_5674,N_5677,N_5678,N_5680,N_5681,N_5683,N_5684,N_5685,N_5686,N_5687,N_5689,N_5690,N_5692,N_5694,N_5696,N_5698,N_5699,N_5700,N_5701,N_5704,N_5705,N_5707,N_5709,N_5710,N_5711,N_5714,N_5719,N_5720,N_5721,N_5722,N_5724,N_5727,N_5731,N_5732,N_5734,N_5738,N_5741,N_5743,N_5746,N_5747,N_5748,N_5750,N_5751,N_5752,N_5753,N_5754,N_5756,N_5757,N_5758,N_5761,N_5763,N_5764,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5777,N_5778,N_5780,N_5781,N_5782,N_5783,N_5784,N_5786,N_5788,N_5790,N_5791,N_5792,N_5794,N_5796,N_5797,N_5798,N_5800,N_5803,N_5805,N_5807,N_5808,N_5810,N_5812,N_5813,N_5814,N_5817,N_5818,N_5819,N_5821,N_5823,N_5826,N_5828,N_5836,N_5837,N_5838,N_5839,N_5842,N_5846,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5855,N_5856,N_5857,N_5858,N_5859,N_5861,N_5862,N_5863,N_5865,N_5867,N_5868,N_5869,N_5871,N_5873,N_5874,N_5876,N_5879,N_5880,N_5882,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5891,N_5892,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5909,N_5911,N_5912,N_5913,N_5914,N_5916,N_5917,N_5919,N_5920,N_5921,N_5922,N_5923,N_5927,N_5929,N_5936,N_5937,N_5939,N_5943,N_5944,N_5945,N_5946,N_5947,N_5949,N_5950,N_5951,N_5952,N_5954,N_5956,N_5958,N_5959,N_5960,N_5962,N_5963,N_5964,N_5966,N_5967,N_5968,N_5969,N_5971,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5985,N_5991,N_5992,N_5993,N_5994,N_5996,N_5997,N_6001,N_6002,N_6003,N_6005,N_6006,N_6007,N_6009,N_6011,N_6012,N_6015,N_6016,N_6017,N_6018,N_6021,N_6022,N_6024,N_6025,N_6028,N_6029,N_6033,N_6034,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6049,N_6053,N_6059,N_6061,N_6062,N_6067,N_6068,N_6071,N_6072,N_6073,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6083,N_6084,N_6087,N_6089,N_6090,N_6091,N_6093,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6122,N_6125,N_6126,N_6128,N_6129,N_6132,N_6134,N_6138,N_6139,N_6140,N_6141,N_6145,N_6146,N_6147,N_6148,N_6150,N_6153,N_6154,N_6155,N_6156,N_6159,N_6160,N_6161,N_6162,N_6164,N_6165,N_6166,N_6167,N_6169,N_6170,N_6172,N_6174,N_6176,N_6179,N_6180,N_6181,N_6182,N_6183,N_6185,N_6187,N_6188,N_6189,N_6190,N_6192,N_6193,N_6194,N_6195,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6213,N_6215,N_6216,N_6217,N_6218,N_6220,N_6221,N_6222,N_6223,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6235,N_6236,N_6237,N_6238,N_6241,N_6242,N_6243,N_6245,N_6246,N_6249,N_6259,N_6260,N_6261,N_6262,N_6265,N_6266,N_6268,N_6269,N_6271,N_6272,N_6273,N_6275,N_6278,N_6280,N_6282,N_6286,N_6287,N_6289,N_6290,N_6294,N_6295,N_6296,N_6298,N_6299,N_6302,N_6303,N_6305,N_6306,N_6308,N_6310,N_6311,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6322,N_6323,N_6324,N_6327,N_6330,N_6332,N_6333,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6352,N_6353,N_6355,N_6356,N_6361,N_6362,N_6363,N_6364,N_6366,N_6368,N_6370,N_6371,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6404,N_6407,N_6408,N_6411,N_6413,N_6414,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6438,N_6439,N_6444,N_6445,N_6448,N_6451,N_6454,N_6458,N_6460,N_6461,N_6462,N_6463,N_6465,N_6466,N_6468,N_6470,N_6471,N_6474,N_6476,N_6477,N_6478,N_6479,N_6480,N_6482,N_6484,N_6485,N_6487,N_6488,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6499,N_6501,N_6503,N_6505,N_6508,N_6509,N_6511,N_6513,N_6514,N_6515,N_6516,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6530,N_6534,N_6535,N_6537,N_6543,N_6545,N_6546,N_6547,N_6548,N_6550,N_6552,N_6553,N_6555,N_6556,N_6560,N_6561,N_6562,N_6563,N_6566,N_6567,N_6571,N_6575,N_6576,N_6577,N_6580,N_6584,N_6586,N_6590,N_6591,N_6596,N_6597,N_6600,N_6603,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6614,N_6616,N_6617,N_6619,N_6621,N_6622,N_6623,N_6626,N_6627,N_6629,N_6630,N_6631,N_6632,N_6633,N_6635,N_6636,N_6637,N_6641,N_6643,N_6644,N_6645,N_6646,N_6648,N_6651,N_6653,N_6655,N_6656,N_6658,N_6659,N_6661,N_6664,N_6666,N_6667,N_6668,N_6669,N_6674,N_6675,N_6676,N_6678,N_6679,N_6685,N_6690,N_6691,N_6692,N_6694,N_6695,N_6696,N_6697,N_6699,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6713,N_6715,N_6717,N_6720,N_6721,N_6722,N_6723,N_6726,N_6727,N_6729,N_6730,N_6731,N_6732,N_6735,N_6740,N_6742,N_6744,N_6745,N_6746,N_6747,N_6748,N_6750,N_6753,N_6755,N_6756,N_6757,N_6760,N_6761,N_6766,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6788,N_6792,N_6793,N_6796,N_6797,N_6799,N_6801,N_6802,N_6803,N_6805,N_6806,N_6807,N_6809,N_6810,N_6813,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6823,N_6825,N_6827,N_6833,N_6834,N_6835,N_6838,N_6840,N_6841,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6856,N_6857,N_6859,N_6860,N_6861,N_6862,N_6864,N_6867,N_6868,N_6871,N_6874,N_6875,N_6876,N_6879,N_6881,N_6882,N_6884,N_6886,N_6889,N_6890,N_6891,N_6892,N_6893,N_6895,N_6896,N_6897,N_6898,N_6900,N_6901,N_6904,N_6906,N_6909,N_6910,N_6911,N_6912,N_6915,N_6916,N_6917,N_6918,N_6919,N_6921,N_6924,N_6925,N_6926,N_6928,N_6929,N_6930,N_6932,N_6934,N_6935,N_6936,N_6938,N_6939,N_6940,N_6941,N_6943,N_6944,N_6945,N_6948,N_6950,N_6953,N_6954,N_6955,N_6956,N_6959,N_6960,N_6961,N_6962,N_6964,N_6965,N_6967,N_6968,N_6969,N_6970,N_6971,N_6973,N_6975,N_6976,N_6979,N_6980,N_6982,N_6984,N_6986,N_6987,N_6990,N_6992,N_6993,N_6996,N_6997,N_6998,N_6999,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7011,N_7012,N_7014,N_7016,N_7017,N_7019,N_7020,N_7021,N_7022,N_7024,N_7025,N_7027,N_7028,N_7030,N_7031,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7042,N_7043,N_7044,N_7045,N_7048,N_7049,N_7050,N_7053,N_7055,N_7056,N_7057,N_7063,N_7064,N_7065,N_7067,N_7068,N_7069,N_7070,N_7072,N_7073,N_7074,N_7076,N_7078,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7087,N_7094,N_7095,N_7100,N_7101,N_7103,N_7105,N_7108,N_7112,N_7113,N_7115,N_7117,N_7119,N_7120,N_7121,N_7124,N_7125,N_7126,N_7127,N_7130,N_7132,N_7135,N_7136,N_7138,N_7140,N_7141,N_7144,N_7145,N_7146,N_7148,N_7149,N_7151,N_7152,N_7153,N_7154,N_7155,N_7158,N_7160,N_7161,N_7162,N_7165,N_7167,N_7168,N_7169,N_7170,N_7171,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7183,N_7185,N_7187,N_7188,N_7189,N_7190,N_7191,N_7193,N_7194,N_7195,N_7198,N_7199,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7213,N_7215,N_7217,N_7218,N_7221,N_7222,N_7224,N_7225,N_7226,N_7228,N_7229,N_7232,N_7233,N_7235,N_7236,N_7237,N_7239,N_7241,N_7242,N_7243,N_7244,N_7245,N_7247,N_7250,N_7253,N_7254,N_7255,N_7256,N_7259,N_7261,N_7266,N_7268,N_7271,N_7272,N_7273,N_7274,N_7279,N_7281,N_7282,N_7283,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7293,N_7294,N_7295,N_7296,N_7300,N_7301,N_7303,N_7304,N_7306,N_7307,N_7308,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7318,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7328,N_7331,N_7332,N_7336,N_7338,N_7340,N_7341,N_7342,N_7343,N_7345,N_7347,N_7348,N_7349,N_7351,N_7352,N_7354,N_7356,N_7357,N_7358,N_7360,N_7362,N_7363,N_7367,N_7368,N_7369,N_7370,N_7373,N_7375,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7387,N_7390,N_7391,N_7394,N_7395,N_7396,N_7397,N_7399,N_7402,N_7403,N_7405,N_7407,N_7409,N_7411,N_7416,N_7417,N_7418,N_7419,N_7420,N_7422,N_7423,N_7426,N_7427,N_7428,N_7434,N_7436,N_7437,N_7438,N_7440,N_7442,N_7443,N_7445,N_7447,N_7449,N_7450,N_7451,N_7456,N_7457,N_7459,N_7462,N_7463,N_7464,N_7468,N_7469,N_7470,N_7471,N_7473,N_7474,N_7476,N_7478,N_7479,N_7480,N_7482,N_7483,N_7485,N_7487,N_7488,N_7489,N_7490,N_7492,N_7493,N_7494,N_7496,N_7497,N_7498,N_7501,N_7502,N_7505,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7518,N_7520,N_7522,N_7523,N_7524,N_7526,N_7527,N_7528,N_7531,N_7532,N_7533,N_7534,N_7537,N_7539,N_7540,N_7541,N_7543,N_7545,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7563,N_7566,N_7569,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7583,N_7584,N_7585,N_7587,N_7588,N_7589,N_7591,N_7592,N_7595,N_7600,N_7602,N_7604,N_7605,N_7607,N_7615,N_7616,N_7618,N_7619,N_7620,N_7621,N_7623,N_7624,N_7625,N_7628,N_7629,N_7630,N_7631,N_7632,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7649,N_7650,N_7651,N_7652,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7663,N_7664,N_7666,N_7667,N_7668,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7678,N_7681,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7691,N_7692,N_7694,N_7695,N_7702,N_7703,N_7704,N_7705,N_7706,N_7708,N_7709,N_7711,N_7712,N_7715,N_7716,N_7717,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7736,N_7738,N_7739,N_7740,N_7742,N_7745,N_7746,N_7747,N_7748,N_7749,N_7751,N_7752,N_7754,N_7755,N_7756,N_7758,N_7760,N_7761,N_7762,N_7763,N_7765,N_7766,N_7767,N_7772,N_7775,N_7776,N_7777,N_7779,N_7780,N_7781,N_7783,N_7784,N_7787,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7797,N_7798,N_7799,N_7801,N_7802,N_7803,N_7804,N_7807,N_7808,N_7809,N_7811,N_7812,N_7817,N_7819,N_7820,N_7822,N_7825,N_7826,N_7827,N_7829,N_7830,N_7832,N_7833,N_7835,N_7836,N_7838,N_7839,N_7842,N_7843,N_7845,N_7846,N_7851,N_7854,N_7855,N_7856,N_7859,N_7861,N_7863,N_7867,N_7870,N_7871,N_7872,N_7875,N_7876,N_7880,N_7881,N_7883,N_7884,N_7885,N_7887,N_7890,N_7891,N_7892,N_7895,N_7897,N_7901,N_7902,N_7903,N_7904,N_7906,N_7908,N_7909,N_7911,N_7912,N_7913,N_7914,N_7917,N_7919,N_7920,N_7921,N_7923,N_7925,N_7929,N_7930,N_7931,N_7932,N_7933,N_7936,N_7939,N_7944,N_7945,N_7946,N_7947,N_7948,N_7950,N_7951,N_7953,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7965,N_7966,N_7969,N_7970,N_7971,N_7974,N_7975,N_7978,N_7979,N_7980,N_7982,N_7983,N_7988,N_7989,N_7990,N_7991,N_7994,N_7995,N_7997,N_8001,N_8002,N_8003,N_8005,N_8006,N_8007,N_8008,N_8015,N_8016,N_8017,N_8021,N_8022,N_8023,N_8024,N_8027,N_8029,N_8030,N_8031,N_8034,N_8036,N_8037,N_8038,N_8040,N_8041,N_8042,N_8043,N_8045,N_8047,N_8048,N_8050,N_8051,N_8054,N_8056,N_8057,N_8058,N_8059,N_8060,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8076,N_8077,N_8078,N_8080,N_8082,N_8083,N_8084,N_8088,N_8089,N_8090,N_8092,N_8093,N_8094,N_8095,N_8098,N_8101,N_8105,N_8107,N_8108,N_8109,N_8111,N_8114,N_8116,N_8117,N_8120,N_8121,N_8122,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8134,N_8135,N_8137,N_8138,N_8141,N_8143,N_8144,N_8145,N_8146,N_8147,N_8149,N_8150,N_8153,N_8154,N_8155,N_8157,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8169,N_8170,N_8171,N_8172,N_8173,N_8176,N_8182,N_8183,N_8184,N_8185,N_8187,N_8189,N_8191,N_8192,N_8196,N_8197,N_8198,N_8199,N_8200,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8211,N_8212,N_8213,N_8214,N_8216,N_8217,N_8218,N_8219,N_8221,N_8223,N_8229,N_8231,N_8232,N_8234,N_8235,N_8236,N_8238,N_8240,N_8241,N_8242,N_8244,N_8250,N_8251,N_8254,N_8257,N_8258,N_8260,N_8262,N_8268,N_8270,N_8272,N_8273,N_8275,N_8277,N_8280,N_8281,N_8282,N_8285,N_8287,N_8289,N_8291,N_8293,N_8297,N_8298,N_8299,N_8300,N_8303,N_8305,N_8307,N_8312,N_8314,N_8315,N_8316,N_8318,N_8321,N_8322,N_8327,N_8330,N_8331,N_8332,N_8333,N_8335,N_8336,N_8340,N_8341,N_8342,N_8343,N_8348,N_8350,N_8351,N_8352,N_8353,N_8357,N_8358,N_8360,N_8361,N_8363,N_8365,N_8366,N_8367,N_8369,N_8371,N_8373,N_8375,N_8377,N_8378,N_8379,N_8380,N_8382,N_8386,N_8387,N_8388,N_8389,N_8391,N_8392,N_8397,N_8398,N_8399,N_8400,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8410,N_8411,N_8413,N_8414,N_8417,N_8418,N_8419,N_8420,N_8421,N_8423,N_8426,N_8427,N_8428,N_8429,N_8430,N_8433,N_8434,N_8436,N_8437,N_8438,N_8441,N_8442,N_8443,N_8445,N_8446,N_8449,N_8450,N_8454,N_8455,N_8459,N_8462,N_8463,N_8465,N_8466,N_8468,N_8471,N_8472,N_8473,N_8474,N_8475,N_8478,N_8479,N_8480,N_8481,N_8482,N_8484,N_8485,N_8486,N_8488,N_8489,N_8490,N_8492,N_8494,N_8495,N_8499,N_8502,N_8503,N_8504,N_8506,N_8507,N_8508,N_8511,N_8513,N_8514,N_8515,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8527,N_8528,N_8531,N_8534,N_8537,N_8541,N_8542,N_8544,N_8550,N_8551,N_8552,N_8553,N_8560,N_8562,N_8563,N_8564,N_8565,N_8568,N_8569,N_8570,N_8573,N_8575,N_8577,N_8580,N_8581,N_8583,N_8584,N_8585,N_8586,N_8588,N_8590,N_8591,N_8592,N_8593,N_8595,N_8596,N_8598,N_8600,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8623,N_8624,N_8625,N_8626,N_8628,N_8629,N_8632,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8642,N_8646,N_8647,N_8648,N_8650,N_8651,N_8652,N_8653,N_8655,N_8656,N_8658,N_8659,N_8660,N_8661,N_8662,N_8668,N_8672,N_8675,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8685,N_8687,N_8688,N_8689,N_8691,N_8692,N_8694,N_8696,N_8697,N_8699,N_8700,N_8701,N_8703,N_8705,N_8706,N_8707,N_8711,N_8715,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8726,N_8727,N_8728,N_8731,N_8734,N_8737,N_8738,N_8741,N_8744,N_8745,N_8748,N_8749,N_8751,N_8753,N_8758,N_8759,N_8761,N_8765,N_8766,N_8769,N_8772,N_8773,N_8774,N_8777,N_8778,N_8779,N_8780,N_8782,N_8784,N_8785,N_8787,N_8788,N_8796,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8807,N_8808,N_8809,N_8810,N_8812,N_8815,N_8816,N_8817,N_8819,N_8821,N_8822,N_8823,N_8826,N_8829,N_8831,N_8832,N_8835,N_8838,N_8844,N_8845,N_8846,N_8847,N_8848,N_8850,N_8851,N_8853,N_8857,N_8859,N_8860,N_8861,N_8864,N_8865,N_8866,N_8867,N_8870,N_8871,N_8873,N_8874,N_8877,N_8878,N_8880,N_8881,N_8886,N_8887,N_8888,N_8889,N_8890,N_8892,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8908,N_8911,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8920,N_8921,N_8923,N_8924,N_8926,N_8927,N_8929,N_8930,N_8932,N_8933,N_8934,N_8935,N_8937,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8950,N_8951,N_8952,N_8954,N_8955,N_8958,N_8960,N_8961,N_8964,N_8966,N_8967,N_8968,N_8970,N_8971,N_8972,N_8974,N_8976,N_8977,N_8979,N_8980,N_8981,N_8982,N_8983,N_8986,N_8987,N_8988,N_8993,N_8995,N_8996,N_8997,N_8998,N_9000,N_9001,N_9003,N_9004,N_9005,N_9006,N_9007,N_9013,N_9014,N_9015,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9026,N_9029,N_9030,N_9032,N_9033,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9048,N_9051,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9063,N_9064,N_9065,N_9066,N_9068,N_9070,N_9071,N_9072,N_9076,N_9077,N_9078,N_9080,N_9085,N_9087,N_9091,N_9093,N_9095,N_9096,N_9098,N_9099,N_9100,N_9101,N_9103,N_9105,N_9106,N_9107,N_9108,N_9109,N_9112,N_9113,N_9115,N_9116,N_9118,N_9120,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9134,N_9137,N_9140,N_9142,N_9144,N_9145,N_9146,N_9148,N_9149,N_9150,N_9152,N_9154,N_9155,N_9157,N_9158,N_9159,N_9161,N_9163,N_9165,N_9166,N_9169,N_9175,N_9176,N_9177,N_9182,N_9186,N_9189,N_9190,N_9192,N_9195,N_9196,N_9198,N_9199,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9209,N_9210,N_9213,N_9214,N_9216,N_9217,N_9218,N_9219,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9234,N_9235,N_9237,N_9240,N_9244,N_9245,N_9246,N_9248,N_9254,N_9256,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9266,N_9271,N_9272,N_9273,N_9274,N_9276,N_9277,N_9278,N_9280,N_9283,N_9284,N_9286,N_9290,N_9291,N_9292,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9317,N_9320,N_9322,N_9324,N_9325,N_9327,N_9329,N_9331,N_9332,N_9333,N_9336,N_9337,N_9338,N_9341,N_9342,N_9344,N_9345,N_9346,N_9348,N_9349,N_9350,N_9351,N_9352,N_9356,N_9358,N_9359,N_9360,N_9361,N_9365,N_9366,N_9368,N_9369,N_9370,N_9373,N_9374,N_9375,N_9376,N_9378,N_9379,N_9380,N_9383,N_9386,N_9389,N_9395,N_9396,N_9399,N_9400,N_9402,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9420,N_9424,N_9426,N_9432,N_9433,N_9434,N_9436,N_9438,N_9440,N_9441,N_9442,N_9443,N_9444,N_9446,N_9447,N_9449,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9459,N_9460,N_9461,N_9462,N_9463,N_9467,N_9468,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9481,N_9482,N_9485,N_9487,N_9488,N_9490,N_9491,N_9492,N_9494,N_9497,N_9499,N_9501,N_9506,N_9509,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9519,N_9520,N_9522,N_9525,N_9526,N_9531,N_9533,N_9534,N_9536,N_9538,N_9540,N_9541,N_9542,N_9546,N_9548,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9558,N_9560,N_9562,N_9565,N_9570,N_9572,N_9574,N_9575,N_9576,N_9577,N_9579,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9590,N_9591,N_9593,N_9595,N_9596,N_9600,N_9601,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9610,N_9613,N_9614,N_9615,N_9616,N_9618,N_9619,N_9622,N_9626,N_9627,N_9629,N_9633,N_9634,N_9635,N_9636,N_9637,N_9639,N_9640,N_9641,N_9643,N_9644,N_9647,N_9648,N_9649,N_9651,N_9652,N_9653,N_9657,N_9658,N_9659,N_9663,N_9667,N_9668,N_9669,N_9671,N_9673,N_9675,N_9677,N_9678,N_9682,N_9684,N_9685,N_9686,N_9690,N_9691,N_9692,N_9694,N_9696,N_9698,N_9703,N_9704,N_9705,N_9707,N_9708,N_9709,N_9710,N_9711,N_9713,N_9714,N_9715,N_9717,N_9718,N_9721,N_9722,N_9723,N_9724,N_9725,N_9727,N_9728,N_9730,N_9731,N_9732,N_9738,N_9739,N_9740,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9757,N_9759,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9771,N_9772,N_9773,N_9775,N_9776,N_9777,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9787,N_9788,N_9789,N_9790,N_9791,N_9793,N_9794,N_9795,N_9797,N_9799,N_9801,N_9803,N_9805,N_9807,N_9808,N_9812,N_9813,N_9814,N_9816,N_9818,N_9823,N_9824,N_9825,N_9827,N_9829,N_9830,N_9831,N_9834,N_9836,N_9838,N_9840,N_9843,N_9845,N_9846,N_9847,N_9848,N_9849,N_9853,N_9854,N_9855,N_9857,N_9858,N_9859,N_9860,N_9863,N_9864,N_9866,N_9867,N_9868,N_9869,N_9870,N_9874,N_9877,N_9878,N_9879,N_9880,N_9883,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9893,N_9897,N_9898,N_9899,N_9900,N_9901,N_9904,N_9905,N_9906,N_9907,N_9908,N_9911,N_9912,N_9917,N_9920,N_9921,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9931,N_9932,N_9934,N_9935,N_9940,N_9941,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9956,N_9957,N_9959,N_9960,N_9961,N_9964,N_9969,N_9971,N_9976,N_9977,N_9979,N_9984,N_9990,N_9992,N_9996,N_9997,N_9998;
nor U0 (N_0,In_589,In_981);
or U1 (N_1,In_874,In_71);
or U2 (N_2,In_163,In_19);
or U3 (N_3,In_285,In_298);
xnor U4 (N_4,In_819,In_100);
xor U5 (N_5,In_446,In_711);
or U6 (N_6,In_788,In_289);
nor U7 (N_7,In_770,In_707);
nor U8 (N_8,In_849,In_101);
nand U9 (N_9,In_161,In_207);
nor U10 (N_10,In_274,In_303);
nor U11 (N_11,In_840,In_66);
or U12 (N_12,In_259,In_629);
and U13 (N_13,In_975,In_103);
or U14 (N_14,In_179,In_605);
nor U15 (N_15,In_215,In_954);
nor U16 (N_16,In_909,In_65);
or U17 (N_17,In_539,In_190);
nand U18 (N_18,In_160,In_483);
or U19 (N_19,In_762,In_678);
nor U20 (N_20,In_169,In_24);
nor U21 (N_21,In_21,In_991);
nand U22 (N_22,In_280,In_292);
nor U23 (N_23,In_372,In_794);
and U24 (N_24,In_481,In_33);
nand U25 (N_25,In_513,In_971);
and U26 (N_26,In_703,In_574);
nand U27 (N_27,In_412,In_815);
nand U28 (N_28,In_168,In_772);
or U29 (N_29,In_959,In_296);
or U30 (N_30,In_369,In_524);
or U31 (N_31,In_955,In_440);
or U32 (N_32,In_778,In_804);
nand U33 (N_33,In_246,In_8);
nand U34 (N_34,In_150,In_308);
or U35 (N_35,In_905,In_630);
nand U36 (N_36,In_699,In_45);
nand U37 (N_37,In_88,In_514);
or U38 (N_38,In_698,In_40);
or U39 (N_39,In_758,In_58);
or U40 (N_40,In_950,In_706);
and U41 (N_41,In_293,In_716);
or U42 (N_42,In_127,In_352);
and U43 (N_43,In_198,In_561);
nor U44 (N_44,In_55,In_805);
nand U45 (N_45,In_133,In_847);
and U46 (N_46,In_976,In_32);
nor U47 (N_47,In_339,In_202);
or U48 (N_48,In_204,In_535);
or U49 (N_49,In_683,In_764);
nand U50 (N_50,In_428,In_261);
or U51 (N_51,In_573,In_624);
nand U52 (N_52,In_121,In_744);
and U53 (N_53,In_516,In_7);
nand U54 (N_54,In_690,In_183);
and U55 (N_55,In_149,In_266);
and U56 (N_56,In_526,In_374);
xor U57 (N_57,In_827,In_789);
nor U58 (N_58,In_432,In_970);
or U59 (N_59,In_37,In_326);
or U60 (N_60,In_852,In_858);
xor U61 (N_61,In_410,In_31);
and U62 (N_62,In_503,In_260);
or U63 (N_63,In_816,In_527);
nor U64 (N_64,In_579,In_155);
or U65 (N_65,In_164,In_502);
or U66 (N_66,In_128,In_418);
nor U67 (N_67,In_748,In_22);
or U68 (N_68,In_845,In_750);
or U69 (N_69,In_757,In_802);
or U70 (N_70,In_294,In_433);
and U71 (N_71,In_893,In_554);
xor U72 (N_72,In_17,In_830);
and U73 (N_73,In_69,In_391);
and U74 (N_74,In_906,In_67);
and U75 (N_75,In_814,In_619);
xor U76 (N_76,In_512,In_60);
and U77 (N_77,In_27,In_543);
or U78 (N_78,In_913,In_413);
nor U79 (N_79,In_91,In_158);
or U80 (N_80,In_140,In_415);
nor U81 (N_81,In_910,In_730);
nand U82 (N_82,In_295,In_299);
or U83 (N_83,In_90,In_242);
nor U84 (N_84,In_931,In_405);
and U85 (N_85,In_315,In_26);
nand U86 (N_86,In_217,In_193);
and U87 (N_87,In_468,In_603);
or U88 (N_88,In_461,In_286);
nand U89 (N_89,In_85,In_776);
nor U90 (N_90,In_640,In_426);
nor U91 (N_91,In_115,In_739);
nand U92 (N_92,In_643,In_325);
or U93 (N_93,In_575,In_321);
or U94 (N_94,In_884,In_466);
and U95 (N_95,In_438,In_663);
and U96 (N_96,In_851,In_634);
or U97 (N_97,In_113,In_137);
or U98 (N_98,In_36,In_928);
nand U99 (N_99,In_701,In_244);
nand U100 (N_100,In_964,In_279);
and U101 (N_101,In_824,In_826);
or U102 (N_102,In_742,In_798);
nand U103 (N_103,In_856,In_612);
or U104 (N_104,In_367,In_552);
xor U105 (N_105,In_329,In_907);
nor U106 (N_106,In_112,In_59);
nand U107 (N_107,In_403,In_474);
and U108 (N_108,In_590,In_153);
or U109 (N_109,In_599,In_685);
nor U110 (N_110,In_616,In_173);
or U111 (N_111,In_876,In_187);
nand U112 (N_112,In_771,In_951);
xnor U113 (N_113,In_201,In_675);
nand U114 (N_114,In_883,In_718);
xor U115 (N_115,In_584,In_598);
and U116 (N_116,In_77,In_602);
nor U117 (N_117,In_16,In_175);
nand U118 (N_118,In_505,In_831);
and U119 (N_119,In_189,In_694);
or U120 (N_120,In_312,In_536);
or U121 (N_121,In_559,In_920);
nand U122 (N_122,In_877,In_277);
nor U123 (N_123,In_427,In_281);
and U124 (N_124,In_562,In_449);
and U125 (N_125,In_867,In_806);
nand U126 (N_126,In_317,In_823);
or U127 (N_127,In_681,In_854);
nand U128 (N_128,In_611,In_324);
nand U129 (N_129,In_741,In_200);
nor U130 (N_130,In_371,In_111);
nor U131 (N_131,In_390,In_857);
nand U132 (N_132,In_366,In_491);
or U133 (N_133,In_737,In_496);
nand U134 (N_134,In_541,In_689);
nand U135 (N_135,In_28,In_769);
and U136 (N_136,In_3,In_566);
and U137 (N_137,In_615,In_754);
or U138 (N_138,In_287,In_900);
nand U139 (N_139,In_779,In_985);
or U140 (N_140,In_662,In_75);
and U141 (N_141,In_887,In_196);
or U142 (N_142,In_822,In_987);
or U143 (N_143,In_763,In_650);
nor U144 (N_144,In_73,In_891);
nor U145 (N_145,In_398,In_923);
nor U146 (N_146,In_469,In_719);
or U147 (N_147,In_64,In_185);
and U148 (N_148,In_444,In_633);
nor U149 (N_149,In_362,In_386);
or U150 (N_150,In_607,In_734);
or U151 (N_151,In_151,In_387);
nand U152 (N_152,In_838,In_656);
nand U153 (N_153,In_264,In_123);
nor U154 (N_154,In_921,In_904);
nor U155 (N_155,In_708,In_34);
nor U156 (N_156,In_839,In_233);
or U157 (N_157,In_447,In_560);
and U158 (N_158,In_903,In_87);
and U159 (N_159,In_862,In_177);
or U160 (N_160,In_389,In_759);
or U161 (N_161,In_382,In_842);
nor U162 (N_162,In_182,In_270);
nand U163 (N_163,In_517,In_866);
or U164 (N_164,In_493,In_546);
or U165 (N_165,In_47,In_458);
nand U166 (N_166,In_143,In_157);
nor U167 (N_167,In_43,In_340);
or U168 (N_168,In_729,In_996);
or U169 (N_169,In_79,In_63);
nor U170 (N_170,In_947,In_765);
nand U171 (N_171,In_829,In_29);
or U172 (N_172,In_859,In_380);
and U173 (N_173,In_869,In_235);
xnor U174 (N_174,In_228,In_338);
and U175 (N_175,In_545,In_646);
nor U176 (N_176,In_635,In_453);
or U177 (N_177,In_747,In_256);
nand U178 (N_178,In_897,In_746);
nor U179 (N_179,In_288,In_948);
nor U180 (N_180,In_14,In_888);
and U181 (N_181,In_820,In_625);
and U182 (N_182,In_728,In_471);
or U183 (N_183,In_333,In_577);
or U184 (N_184,In_732,In_178);
xnor U185 (N_185,In_872,In_231);
and U186 (N_186,In_654,In_301);
nand U187 (N_187,In_636,In_12);
and U188 (N_188,In_214,In_434);
or U189 (N_189,In_655,In_247);
and U190 (N_190,In_376,In_997);
and U191 (N_191,In_585,In_506);
or U192 (N_192,In_457,In_501);
nor U193 (N_193,In_523,In_125);
nor U194 (N_194,In_817,In_930);
nand U195 (N_195,In_530,In_620);
and U196 (N_196,In_966,In_166);
nor U197 (N_197,In_323,In_351);
nand U198 (N_198,In_538,In_870);
nand U199 (N_199,In_430,In_74);
and U200 (N_200,In_138,In_886);
and U201 (N_201,In_709,In_319);
or U202 (N_202,In_249,In_318);
nand U203 (N_203,In_146,In_495);
or U204 (N_204,In_11,In_238);
nand U205 (N_205,In_368,In_54);
and U206 (N_206,In_464,In_642);
and U207 (N_207,In_250,In_600);
nand U208 (N_208,In_652,In_409);
or U209 (N_209,In_253,In_373);
nor U210 (N_210,In_223,In_420);
nor U211 (N_211,In_393,In_686);
nand U212 (N_212,In_898,In_417);
and U213 (N_213,In_199,In_358);
or U214 (N_214,In_555,In_665);
or U215 (N_215,In_937,In_962);
and U216 (N_216,In_509,In_723);
nor U217 (N_217,In_375,In_812);
nand U218 (N_218,In_832,In_484);
xor U219 (N_219,In_775,In_343);
and U220 (N_220,In_745,In_786);
and U221 (N_221,In_861,In_52);
nor U222 (N_222,In_365,In_347);
nor U223 (N_223,In_508,In_676);
or U224 (N_224,In_226,In_855);
nand U225 (N_225,In_572,In_693);
nand U226 (N_226,In_846,In_557);
and U227 (N_227,In_197,In_442);
or U228 (N_228,In_422,In_480);
or U229 (N_229,In_126,In_960);
or U230 (N_230,In_229,In_743);
nand U231 (N_231,In_212,In_334);
and U232 (N_232,In_184,In_682);
or U233 (N_233,In_721,In_592);
nor U234 (N_234,In_632,In_850);
and U235 (N_235,In_623,In_740);
nor U236 (N_236,In_567,In_455);
or U237 (N_237,In_83,In_932);
xnor U238 (N_238,In_116,In_377);
nand U239 (N_239,In_205,In_306);
and U240 (N_240,In_738,In_498);
nor U241 (N_241,In_307,In_582);
and U242 (N_242,In_245,In_606);
or U243 (N_243,In_156,In_96);
and U244 (N_244,In_482,In_176);
and U245 (N_245,In_674,In_853);
nand U246 (N_246,In_548,In_811);
xor U247 (N_247,In_20,In_622);
nor U248 (N_248,In_222,In_320);
or U249 (N_249,In_132,In_349);
nor U250 (N_250,In_594,In_983);
or U251 (N_251,In_843,In_401);
nand U252 (N_252,In_194,In_86);
nand U253 (N_253,In_702,In_97);
or U254 (N_254,In_973,In_467);
nor U255 (N_255,In_206,In_595);
nand U256 (N_256,In_188,In_396);
nor U257 (N_257,In_441,In_980);
nor U258 (N_258,In_477,In_300);
nand U259 (N_259,In_218,In_357);
or U260 (N_260,In_672,In_961);
nor U261 (N_261,In_265,In_551);
and U262 (N_262,In_863,In_916);
or U263 (N_263,In_117,In_72);
nand U264 (N_264,In_549,In_518);
and U265 (N_265,In_82,In_10);
nor U266 (N_266,In_547,In_912);
or U267 (N_267,In_221,In_448);
nor U268 (N_268,In_531,In_472);
and U269 (N_269,In_726,In_70);
nand U270 (N_270,In_337,In_475);
or U271 (N_271,In_998,In_171);
nor U272 (N_272,In_208,In_783);
or U273 (N_273,In_381,In_492);
nor U274 (N_274,In_346,In_684);
nand U275 (N_275,In_774,In_297);
nor U276 (N_276,In_302,In_565);
nor U277 (N_277,In_152,In_416);
or U278 (N_278,In_649,In_813);
and U279 (N_279,In_141,In_570);
nor U280 (N_280,In_735,In_715);
or U281 (N_281,In_658,In_924);
nor U282 (N_282,In_345,In_407);
or U283 (N_283,In_553,In_569);
or U284 (N_284,In_435,In_986);
or U285 (N_285,In_515,In_645);
and U286 (N_286,In_56,In_679);
nor U287 (N_287,In_142,In_353);
and U288 (N_288,In_341,In_563);
or U289 (N_289,In_220,In_618);
or U290 (N_290,In_882,In_62);
or U291 (N_291,In_940,In_470);
nand U292 (N_292,In_136,In_258);
nand U293 (N_293,In_773,In_425);
nor U294 (N_294,In_972,In_692);
nor U295 (N_295,In_94,In_49);
nand U296 (N_296,In_348,In_236);
or U297 (N_297,In_239,In_439);
or U298 (N_298,In_473,In_76);
nand U299 (N_299,In_408,In_118);
or U300 (N_300,In_13,In_993);
and U301 (N_301,In_313,In_958);
nor U302 (N_302,In_613,In_792);
and U303 (N_303,In_946,In_587);
or U304 (N_304,In_934,In_465);
nor U305 (N_305,In_801,In_880);
or U306 (N_306,In_450,In_808);
nand U307 (N_307,In_105,In_532);
nand U308 (N_308,In_568,In_511);
nor U309 (N_309,In_915,In_889);
nand U310 (N_310,In_942,In_35);
or U311 (N_311,In_489,In_174);
and U312 (N_312,In_219,In_578);
and U313 (N_313,In_363,In_456);
nor U314 (N_314,In_310,In_952);
nand U315 (N_315,In_271,In_104);
xor U316 (N_316,In_660,In_195);
or U317 (N_317,In_688,In_305);
nor U318 (N_318,In_476,In_637);
nand U319 (N_319,In_782,In_130);
nor U320 (N_320,In_712,In_167);
nand U321 (N_321,In_938,In_571);
or U322 (N_322,In_925,In_664);
and U323 (N_323,In_99,In_478);
nor U324 (N_324,In_626,In_922);
and U325 (N_325,In_180,In_507);
or U326 (N_326,In_644,In_134);
nand U327 (N_327,In_963,In_225);
and U328 (N_328,In_53,In_5);
nor U329 (N_329,In_81,In_454);
or U330 (N_330,In_879,In_429);
nand U331 (N_331,In_935,In_841);
and U332 (N_332,In_360,In_901);
and U333 (N_333,In_825,In_404);
or U334 (N_334,In_673,In_810);
nor U335 (N_335,In_576,In_895);
nor U336 (N_336,In_6,In_550);
or U337 (N_337,In_165,In_525);
nor U338 (N_338,In_821,In_790);
nor U339 (N_339,In_278,In_596);
and U340 (N_340,In_544,In_537);
or U341 (N_341,In_350,In_172);
nor U342 (N_342,In_314,In_283);
nand U343 (N_343,In_593,In_240);
nand U344 (N_344,In_868,In_443);
nand U345 (N_345,In_361,In_399);
nor U346 (N_346,In_601,In_918);
or U347 (N_347,In_908,In_704);
xnor U348 (N_348,In_990,In_392);
nand U349 (N_349,In_186,In_41);
nor U350 (N_350,In_9,In_979);
or U351 (N_351,In_713,In_795);
nand U352 (N_352,In_275,In_272);
or U353 (N_353,In_809,In_497);
or U354 (N_354,In_753,In_38);
or U355 (N_355,In_490,In_385);
and U356 (N_356,In_147,In_761);
or U357 (N_357,In_108,In_423);
nand U358 (N_358,In_731,In_965);
and U359 (N_359,In_462,In_500);
nand U360 (N_360,In_51,In_252);
or U361 (N_361,In_641,In_230);
nand U362 (N_362,In_974,In_680);
or U363 (N_363,In_639,In_628);
and U364 (N_364,In_988,In_720);
or U365 (N_365,In_799,In_335);
nor U366 (N_366,In_463,In_631);
and U367 (N_367,In_638,In_1);
or U368 (N_368,In_4,In_322);
nand U369 (N_369,In_793,In_833);
and U370 (N_370,In_944,In_591);
and U371 (N_371,In_402,In_755);
or U372 (N_372,In_556,In_522);
nor U373 (N_373,In_659,In_837);
or U374 (N_374,In_273,In_336);
xnor U375 (N_375,In_989,In_92);
or U376 (N_376,In_785,In_733);
nand U377 (N_377,In_209,In_995);
or U378 (N_378,In_784,In_949);
nor U379 (N_379,In_44,In_263);
and U380 (N_380,In_95,In_50);
or U381 (N_381,In_604,In_46);
or U382 (N_382,In_98,In_871);
nand U383 (N_383,In_929,In_316);
nor U384 (N_384,In_330,In_445);
nor U385 (N_385,In_529,In_648);
nor U386 (N_386,In_583,In_257);
nor U387 (N_387,In_885,In_621);
nand U388 (N_388,In_896,In_120);
nand U389 (N_389,In_276,In_42);
nor U390 (N_390,In_807,In_327);
and U391 (N_391,In_129,In_145);
and U392 (N_392,In_344,In_653);
nand U393 (N_393,In_677,In_521);
nor U394 (N_394,In_394,In_397);
nand U395 (N_395,In_192,In_982);
nand U396 (N_396,In_647,In_107);
nand U397 (N_397,In_356,In_864);
nor U398 (N_398,In_234,In_452);
xor U399 (N_399,In_332,In_170);
and U400 (N_400,In_388,In_714);
nor U401 (N_401,In_580,In_213);
and U402 (N_402,In_227,In_736);
nor U403 (N_403,In_902,In_78);
nand U404 (N_404,In_967,In_777);
or U405 (N_405,In_370,In_666);
nand U406 (N_406,In_119,In_57);
nor U407 (N_407,In_834,In_917);
nor U408 (N_408,In_384,In_926);
nand U409 (N_409,In_597,In_558);
xor U410 (N_410,In_796,In_224);
or U411 (N_411,In_255,In_749);
nand U412 (N_412,In_860,In_400);
and U413 (N_413,In_110,In_705);
or U414 (N_414,In_135,In_608);
or U415 (N_415,In_700,In_309);
nand U416 (N_416,In_978,In_520);
or U417 (N_417,In_210,In_766);
nor U418 (N_418,In_781,In_767);
and U419 (N_419,In_487,In_939);
nand U420 (N_420,In_941,In_378);
nor U421 (N_421,In_328,In_459);
nor U422 (N_422,In_803,In_379);
and U423 (N_423,In_267,In_994);
and U424 (N_424,In_984,In_486);
and U425 (N_425,In_211,In_80);
or U426 (N_426,In_181,In_534);
and U427 (N_427,In_881,In_93);
xnor U428 (N_428,In_667,In_460);
nand U429 (N_429,In_945,In_451);
nor U430 (N_430,In_724,In_878);
and U431 (N_431,In_436,In_943);
or U432 (N_432,In_268,In_844);
or U433 (N_433,In_581,In_61);
nor U434 (N_434,In_395,In_354);
or U435 (N_435,In_203,In_751);
or U436 (N_436,In_124,In_890);
or U437 (N_437,In_424,In_494);
nand U438 (N_438,In_254,In_953);
or U439 (N_439,In_614,In_725);
nor U440 (N_440,In_162,In_0);
or U441 (N_441,In_610,In_586);
nand U442 (N_442,In_2,In_691);
nand U443 (N_443,In_668,In_437);
and U444 (N_444,In_710,In_669);
nand U445 (N_445,In_144,In_957);
nand U446 (N_446,In_717,In_89);
nand U447 (N_447,In_421,In_919);
or U448 (N_448,In_695,In_102);
nor U449 (N_449,In_800,In_760);
nand U450 (N_450,In_139,In_311);
nand U451 (N_451,In_836,In_383);
xnor U452 (N_452,In_927,In_122);
or U453 (N_453,In_875,In_414);
nor U454 (N_454,In_342,In_892);
xor U455 (N_455,In_232,In_911);
or U456 (N_456,In_670,In_787);
nand U457 (N_457,In_18,In_488);
or U458 (N_458,In_791,In_564);
nor U459 (N_459,In_504,In_894);
or U460 (N_460,In_84,In_304);
nor U461 (N_461,In_331,In_431);
or U462 (N_462,In_848,In_657);
or U463 (N_463,In_533,In_627);
nand U464 (N_464,In_899,In_977);
nand U465 (N_465,In_828,In_499);
nand U466 (N_466,In_109,In_291);
nor U467 (N_467,In_243,In_479);
and U468 (N_468,In_154,In_780);
nor U469 (N_469,In_835,In_756);
or U470 (N_470,In_933,In_114);
nand U471 (N_471,In_510,In_914);
nor U472 (N_472,In_106,In_609);
nand U473 (N_473,In_671,In_248);
nor U474 (N_474,In_419,In_355);
nor U475 (N_475,In_485,In_696);
nor U476 (N_476,In_290,In_617);
and U477 (N_477,In_727,In_25);
nand U478 (N_478,In_999,In_540);
nand U479 (N_479,In_406,In_48);
nand U480 (N_480,In_30,In_411);
or U481 (N_481,In_661,In_797);
or U482 (N_482,In_269,In_873);
and U483 (N_483,In_216,In_191);
nand U484 (N_484,In_68,In_282);
nor U485 (N_485,In_818,In_251);
nand U486 (N_486,In_651,In_159);
nor U487 (N_487,In_284,In_528);
nor U488 (N_488,In_131,In_992);
nand U489 (N_489,In_359,In_519);
nand U490 (N_490,In_936,In_148);
or U491 (N_491,In_768,In_364);
nand U492 (N_492,In_15,In_241);
nor U493 (N_493,In_956,In_237);
or U494 (N_494,In_262,In_865);
nand U495 (N_495,In_697,In_969);
xor U496 (N_496,In_968,In_23);
nor U497 (N_497,In_588,In_39);
nand U498 (N_498,In_752,In_542);
nand U499 (N_499,In_687,In_722);
nand U500 (N_500,In_314,In_865);
and U501 (N_501,In_954,In_535);
nor U502 (N_502,In_527,In_600);
or U503 (N_503,In_453,In_817);
nand U504 (N_504,In_76,In_732);
or U505 (N_505,In_932,In_236);
nand U506 (N_506,In_266,In_765);
xor U507 (N_507,In_243,In_365);
and U508 (N_508,In_406,In_973);
nand U509 (N_509,In_710,In_217);
and U510 (N_510,In_300,In_275);
and U511 (N_511,In_831,In_4);
nor U512 (N_512,In_842,In_574);
xor U513 (N_513,In_527,In_78);
nor U514 (N_514,In_66,In_690);
or U515 (N_515,In_507,In_945);
or U516 (N_516,In_67,In_705);
nor U517 (N_517,In_40,In_204);
or U518 (N_518,In_408,In_813);
or U519 (N_519,In_183,In_112);
nand U520 (N_520,In_658,In_559);
nor U521 (N_521,In_914,In_94);
nand U522 (N_522,In_882,In_442);
nor U523 (N_523,In_237,In_96);
nand U524 (N_524,In_147,In_266);
or U525 (N_525,In_556,In_244);
xnor U526 (N_526,In_965,In_886);
xnor U527 (N_527,In_724,In_209);
nand U528 (N_528,In_448,In_39);
nor U529 (N_529,In_33,In_17);
nand U530 (N_530,In_676,In_68);
or U531 (N_531,In_613,In_662);
or U532 (N_532,In_852,In_687);
or U533 (N_533,In_170,In_151);
or U534 (N_534,In_371,In_975);
nand U535 (N_535,In_971,In_905);
nor U536 (N_536,In_857,In_117);
nor U537 (N_537,In_193,In_804);
or U538 (N_538,In_418,In_89);
nand U539 (N_539,In_867,In_17);
and U540 (N_540,In_157,In_5);
and U541 (N_541,In_271,In_136);
xor U542 (N_542,In_990,In_744);
nand U543 (N_543,In_782,In_191);
or U544 (N_544,In_287,In_39);
and U545 (N_545,In_342,In_139);
nand U546 (N_546,In_303,In_583);
nor U547 (N_547,In_537,In_747);
and U548 (N_548,In_282,In_681);
nor U549 (N_549,In_772,In_821);
nand U550 (N_550,In_781,In_488);
nor U551 (N_551,In_149,In_666);
nand U552 (N_552,In_90,In_256);
and U553 (N_553,In_476,In_725);
nor U554 (N_554,In_133,In_80);
nor U555 (N_555,In_86,In_589);
nor U556 (N_556,In_33,In_919);
or U557 (N_557,In_541,In_950);
or U558 (N_558,In_591,In_464);
and U559 (N_559,In_645,In_503);
or U560 (N_560,In_368,In_707);
and U561 (N_561,In_147,In_557);
nand U562 (N_562,In_996,In_315);
nand U563 (N_563,In_230,In_622);
nor U564 (N_564,In_753,In_136);
nand U565 (N_565,In_991,In_609);
nor U566 (N_566,In_874,In_428);
nand U567 (N_567,In_465,In_585);
and U568 (N_568,In_995,In_109);
nor U569 (N_569,In_121,In_311);
or U570 (N_570,In_363,In_550);
nand U571 (N_571,In_972,In_856);
or U572 (N_572,In_932,In_691);
nor U573 (N_573,In_138,In_487);
nand U574 (N_574,In_881,In_235);
or U575 (N_575,In_782,In_767);
nand U576 (N_576,In_620,In_520);
and U577 (N_577,In_743,In_823);
nand U578 (N_578,In_78,In_714);
or U579 (N_579,In_746,In_728);
or U580 (N_580,In_815,In_385);
nor U581 (N_581,In_258,In_180);
nor U582 (N_582,In_883,In_451);
and U583 (N_583,In_874,In_835);
and U584 (N_584,In_562,In_978);
xor U585 (N_585,In_183,In_387);
or U586 (N_586,In_371,In_296);
nor U587 (N_587,In_497,In_251);
and U588 (N_588,In_605,In_846);
and U589 (N_589,In_17,In_777);
nand U590 (N_590,In_593,In_790);
nor U591 (N_591,In_532,In_347);
nor U592 (N_592,In_735,In_789);
and U593 (N_593,In_773,In_524);
and U594 (N_594,In_91,In_455);
nand U595 (N_595,In_132,In_274);
or U596 (N_596,In_722,In_69);
nand U597 (N_597,In_898,In_90);
nor U598 (N_598,In_430,In_573);
and U599 (N_599,In_64,In_813);
nand U600 (N_600,In_257,In_855);
and U601 (N_601,In_454,In_186);
or U602 (N_602,In_190,In_498);
or U603 (N_603,In_169,In_16);
nand U604 (N_604,In_536,In_643);
and U605 (N_605,In_500,In_233);
and U606 (N_606,In_7,In_874);
nor U607 (N_607,In_15,In_689);
nor U608 (N_608,In_377,In_747);
nor U609 (N_609,In_229,In_860);
nand U610 (N_610,In_749,In_748);
or U611 (N_611,In_329,In_250);
and U612 (N_612,In_544,In_86);
or U613 (N_613,In_69,In_430);
and U614 (N_614,In_927,In_185);
or U615 (N_615,In_374,In_340);
nor U616 (N_616,In_984,In_925);
nor U617 (N_617,In_962,In_627);
xnor U618 (N_618,In_704,In_44);
nand U619 (N_619,In_757,In_52);
or U620 (N_620,In_402,In_671);
nor U621 (N_621,In_17,In_311);
nand U622 (N_622,In_546,In_858);
nor U623 (N_623,In_595,In_98);
nand U624 (N_624,In_551,In_538);
nor U625 (N_625,In_545,In_428);
and U626 (N_626,In_594,In_602);
nor U627 (N_627,In_635,In_792);
nand U628 (N_628,In_513,In_749);
nand U629 (N_629,In_724,In_449);
nand U630 (N_630,In_73,In_324);
nand U631 (N_631,In_783,In_450);
nor U632 (N_632,In_157,In_405);
xor U633 (N_633,In_440,In_270);
and U634 (N_634,In_940,In_529);
and U635 (N_635,In_574,In_113);
nand U636 (N_636,In_975,In_24);
and U637 (N_637,In_715,In_627);
and U638 (N_638,In_903,In_595);
or U639 (N_639,In_391,In_867);
nand U640 (N_640,In_113,In_422);
or U641 (N_641,In_121,In_867);
nand U642 (N_642,In_588,In_937);
or U643 (N_643,In_965,In_602);
or U644 (N_644,In_573,In_105);
nor U645 (N_645,In_631,In_209);
and U646 (N_646,In_215,In_14);
and U647 (N_647,In_554,In_434);
and U648 (N_648,In_121,In_214);
or U649 (N_649,In_89,In_84);
or U650 (N_650,In_793,In_66);
nand U651 (N_651,In_388,In_917);
nor U652 (N_652,In_848,In_742);
nand U653 (N_653,In_785,In_740);
or U654 (N_654,In_58,In_424);
nor U655 (N_655,In_553,In_762);
and U656 (N_656,In_33,In_46);
nand U657 (N_657,In_502,In_273);
nor U658 (N_658,In_367,In_804);
or U659 (N_659,In_501,In_356);
and U660 (N_660,In_826,In_436);
nand U661 (N_661,In_832,In_596);
and U662 (N_662,In_55,In_259);
nor U663 (N_663,In_709,In_143);
or U664 (N_664,In_982,In_650);
or U665 (N_665,In_875,In_179);
or U666 (N_666,In_138,In_780);
and U667 (N_667,In_436,In_399);
nor U668 (N_668,In_434,In_595);
or U669 (N_669,In_490,In_537);
nand U670 (N_670,In_616,In_342);
nand U671 (N_671,In_569,In_917);
nor U672 (N_672,In_665,In_33);
or U673 (N_673,In_579,In_31);
nand U674 (N_674,In_247,In_298);
nand U675 (N_675,In_978,In_568);
nand U676 (N_676,In_837,In_420);
nor U677 (N_677,In_28,In_843);
and U678 (N_678,In_797,In_392);
nand U679 (N_679,In_986,In_551);
nor U680 (N_680,In_430,In_301);
or U681 (N_681,In_928,In_584);
nand U682 (N_682,In_679,In_659);
nor U683 (N_683,In_117,In_261);
nand U684 (N_684,In_865,In_10);
and U685 (N_685,In_219,In_968);
or U686 (N_686,In_953,In_877);
and U687 (N_687,In_922,In_77);
and U688 (N_688,In_9,In_51);
nand U689 (N_689,In_844,In_972);
nor U690 (N_690,In_464,In_781);
nor U691 (N_691,In_175,In_582);
and U692 (N_692,In_758,In_121);
nor U693 (N_693,In_681,In_610);
and U694 (N_694,In_453,In_859);
or U695 (N_695,In_153,In_188);
and U696 (N_696,In_80,In_103);
nand U697 (N_697,In_938,In_642);
nor U698 (N_698,In_25,In_30);
nand U699 (N_699,In_921,In_614);
and U700 (N_700,In_526,In_798);
and U701 (N_701,In_963,In_261);
and U702 (N_702,In_86,In_921);
and U703 (N_703,In_464,In_876);
or U704 (N_704,In_478,In_243);
nor U705 (N_705,In_670,In_442);
nand U706 (N_706,In_338,In_22);
nor U707 (N_707,In_748,In_123);
nand U708 (N_708,In_400,In_837);
nor U709 (N_709,In_42,In_142);
and U710 (N_710,In_239,In_90);
nor U711 (N_711,In_904,In_506);
or U712 (N_712,In_659,In_581);
and U713 (N_713,In_18,In_750);
or U714 (N_714,In_832,In_507);
and U715 (N_715,In_514,In_756);
nor U716 (N_716,In_208,In_877);
nand U717 (N_717,In_470,In_107);
nor U718 (N_718,In_269,In_567);
nand U719 (N_719,In_523,In_852);
and U720 (N_720,In_82,In_956);
nor U721 (N_721,In_379,In_156);
and U722 (N_722,In_541,In_755);
nand U723 (N_723,In_503,In_89);
or U724 (N_724,In_817,In_779);
or U725 (N_725,In_772,In_776);
and U726 (N_726,In_625,In_68);
nand U727 (N_727,In_9,In_475);
or U728 (N_728,In_603,In_747);
or U729 (N_729,In_374,In_527);
or U730 (N_730,In_839,In_127);
nor U731 (N_731,In_530,In_464);
nand U732 (N_732,In_193,In_94);
xor U733 (N_733,In_950,In_610);
or U734 (N_734,In_265,In_174);
or U735 (N_735,In_703,In_177);
and U736 (N_736,In_169,In_698);
nor U737 (N_737,In_735,In_418);
nand U738 (N_738,In_875,In_793);
and U739 (N_739,In_154,In_923);
nor U740 (N_740,In_418,In_64);
nand U741 (N_741,In_659,In_908);
and U742 (N_742,In_456,In_145);
or U743 (N_743,In_230,In_448);
nand U744 (N_744,In_630,In_593);
nor U745 (N_745,In_912,In_216);
or U746 (N_746,In_670,In_559);
nand U747 (N_747,In_385,In_492);
nor U748 (N_748,In_752,In_950);
nor U749 (N_749,In_884,In_720);
or U750 (N_750,In_579,In_891);
nor U751 (N_751,In_179,In_988);
or U752 (N_752,In_875,In_947);
nand U753 (N_753,In_369,In_668);
nand U754 (N_754,In_980,In_737);
xor U755 (N_755,In_24,In_841);
and U756 (N_756,In_901,In_745);
or U757 (N_757,In_434,In_320);
nand U758 (N_758,In_355,In_397);
and U759 (N_759,In_174,In_638);
nand U760 (N_760,In_891,In_438);
and U761 (N_761,In_959,In_982);
and U762 (N_762,In_61,In_262);
or U763 (N_763,In_93,In_277);
and U764 (N_764,In_415,In_938);
or U765 (N_765,In_480,In_897);
or U766 (N_766,In_984,In_358);
nand U767 (N_767,In_815,In_560);
and U768 (N_768,In_557,In_934);
nand U769 (N_769,In_439,In_757);
or U770 (N_770,In_794,In_855);
and U771 (N_771,In_469,In_73);
or U772 (N_772,In_347,In_159);
or U773 (N_773,In_542,In_626);
and U774 (N_774,In_416,In_685);
nor U775 (N_775,In_845,In_518);
nor U776 (N_776,In_844,In_920);
and U777 (N_777,In_50,In_714);
and U778 (N_778,In_658,In_586);
and U779 (N_779,In_991,In_133);
or U780 (N_780,In_303,In_633);
and U781 (N_781,In_181,In_712);
nand U782 (N_782,In_145,In_313);
nor U783 (N_783,In_107,In_231);
nand U784 (N_784,In_922,In_592);
or U785 (N_785,In_397,In_864);
or U786 (N_786,In_444,In_791);
xnor U787 (N_787,In_358,In_243);
and U788 (N_788,In_132,In_565);
xnor U789 (N_789,In_137,In_77);
nand U790 (N_790,In_864,In_718);
nor U791 (N_791,In_717,In_841);
nor U792 (N_792,In_329,In_395);
nand U793 (N_793,In_550,In_919);
nand U794 (N_794,In_126,In_512);
or U795 (N_795,In_770,In_278);
and U796 (N_796,In_717,In_19);
or U797 (N_797,In_896,In_274);
xor U798 (N_798,In_944,In_64);
and U799 (N_799,In_895,In_122);
nand U800 (N_800,In_820,In_8);
or U801 (N_801,In_150,In_729);
or U802 (N_802,In_797,In_701);
and U803 (N_803,In_91,In_696);
nor U804 (N_804,In_507,In_570);
nand U805 (N_805,In_912,In_260);
or U806 (N_806,In_263,In_223);
nor U807 (N_807,In_599,In_324);
and U808 (N_808,In_501,In_379);
or U809 (N_809,In_837,In_938);
nor U810 (N_810,In_545,In_460);
nor U811 (N_811,In_588,In_471);
and U812 (N_812,In_669,In_982);
and U813 (N_813,In_142,In_419);
nor U814 (N_814,In_647,In_368);
nand U815 (N_815,In_422,In_910);
nor U816 (N_816,In_30,In_677);
nand U817 (N_817,In_938,In_489);
or U818 (N_818,In_176,In_724);
and U819 (N_819,In_802,In_162);
nor U820 (N_820,In_791,In_178);
nor U821 (N_821,In_689,In_37);
nand U822 (N_822,In_12,In_39);
or U823 (N_823,In_432,In_651);
nand U824 (N_824,In_562,In_785);
or U825 (N_825,In_824,In_588);
nand U826 (N_826,In_753,In_565);
nor U827 (N_827,In_573,In_958);
nand U828 (N_828,In_737,In_382);
nor U829 (N_829,In_769,In_568);
nor U830 (N_830,In_465,In_240);
nand U831 (N_831,In_165,In_831);
nor U832 (N_832,In_138,In_634);
and U833 (N_833,In_306,In_576);
and U834 (N_834,In_798,In_437);
nor U835 (N_835,In_674,In_866);
nand U836 (N_836,In_61,In_448);
xnor U837 (N_837,In_526,In_917);
nand U838 (N_838,In_806,In_402);
nor U839 (N_839,In_353,In_80);
nor U840 (N_840,In_583,In_3);
nand U841 (N_841,In_905,In_245);
and U842 (N_842,In_140,In_671);
xnor U843 (N_843,In_497,In_486);
or U844 (N_844,In_129,In_896);
nand U845 (N_845,In_646,In_450);
nor U846 (N_846,In_482,In_332);
nand U847 (N_847,In_794,In_355);
xor U848 (N_848,In_841,In_989);
nor U849 (N_849,In_130,In_908);
or U850 (N_850,In_100,In_696);
nor U851 (N_851,In_263,In_8);
nand U852 (N_852,In_964,In_65);
nor U853 (N_853,In_868,In_289);
nand U854 (N_854,In_488,In_581);
nand U855 (N_855,In_793,In_62);
and U856 (N_856,In_720,In_597);
and U857 (N_857,In_575,In_58);
or U858 (N_858,In_430,In_189);
and U859 (N_859,In_180,In_39);
or U860 (N_860,In_478,In_931);
nand U861 (N_861,In_532,In_76);
nand U862 (N_862,In_852,In_812);
nand U863 (N_863,In_855,In_125);
and U864 (N_864,In_903,In_611);
nand U865 (N_865,In_480,In_298);
and U866 (N_866,In_894,In_536);
and U867 (N_867,In_950,In_558);
nor U868 (N_868,In_340,In_740);
nor U869 (N_869,In_607,In_288);
and U870 (N_870,In_411,In_150);
and U871 (N_871,In_410,In_293);
or U872 (N_872,In_707,In_136);
nor U873 (N_873,In_762,In_948);
and U874 (N_874,In_90,In_466);
nor U875 (N_875,In_514,In_33);
nand U876 (N_876,In_525,In_386);
or U877 (N_877,In_345,In_172);
nor U878 (N_878,In_825,In_211);
nand U879 (N_879,In_2,In_561);
nor U880 (N_880,In_292,In_99);
and U881 (N_881,In_576,In_124);
nor U882 (N_882,In_788,In_694);
nor U883 (N_883,In_816,In_965);
nor U884 (N_884,In_209,In_728);
xnor U885 (N_885,In_780,In_237);
nand U886 (N_886,In_819,In_896);
or U887 (N_887,In_485,In_257);
or U888 (N_888,In_429,In_482);
nor U889 (N_889,In_719,In_21);
nand U890 (N_890,In_108,In_181);
and U891 (N_891,In_961,In_0);
nand U892 (N_892,In_814,In_390);
and U893 (N_893,In_707,In_246);
nor U894 (N_894,In_110,In_703);
or U895 (N_895,In_800,In_125);
or U896 (N_896,In_988,In_927);
nand U897 (N_897,In_293,In_23);
and U898 (N_898,In_76,In_110);
nand U899 (N_899,In_406,In_271);
nand U900 (N_900,In_149,In_676);
nor U901 (N_901,In_695,In_298);
or U902 (N_902,In_562,In_74);
and U903 (N_903,In_530,In_109);
nand U904 (N_904,In_659,In_583);
nor U905 (N_905,In_626,In_855);
nor U906 (N_906,In_273,In_783);
nand U907 (N_907,In_252,In_209);
nor U908 (N_908,In_390,In_570);
or U909 (N_909,In_874,In_892);
xnor U910 (N_910,In_698,In_61);
nand U911 (N_911,In_879,In_540);
nor U912 (N_912,In_34,In_711);
nor U913 (N_913,In_610,In_284);
nor U914 (N_914,In_913,In_302);
nand U915 (N_915,In_811,In_498);
and U916 (N_916,In_967,In_136);
or U917 (N_917,In_294,In_632);
nor U918 (N_918,In_152,In_882);
nor U919 (N_919,In_865,In_71);
and U920 (N_920,In_891,In_478);
nor U921 (N_921,In_743,In_284);
and U922 (N_922,In_579,In_787);
xnor U923 (N_923,In_719,In_779);
and U924 (N_924,In_302,In_271);
nor U925 (N_925,In_817,In_202);
nor U926 (N_926,In_680,In_70);
xnor U927 (N_927,In_381,In_711);
nand U928 (N_928,In_191,In_894);
nand U929 (N_929,In_57,In_918);
xnor U930 (N_930,In_831,In_700);
nor U931 (N_931,In_753,In_839);
and U932 (N_932,In_98,In_604);
or U933 (N_933,In_988,In_13);
nand U934 (N_934,In_731,In_284);
nand U935 (N_935,In_663,In_530);
nand U936 (N_936,In_371,In_505);
or U937 (N_937,In_336,In_481);
and U938 (N_938,In_22,In_160);
nor U939 (N_939,In_587,In_59);
or U940 (N_940,In_619,In_928);
nand U941 (N_941,In_987,In_697);
or U942 (N_942,In_859,In_349);
or U943 (N_943,In_740,In_493);
or U944 (N_944,In_797,In_231);
or U945 (N_945,In_694,In_281);
or U946 (N_946,In_374,In_102);
and U947 (N_947,In_410,In_364);
xor U948 (N_948,In_684,In_743);
nand U949 (N_949,In_639,In_278);
or U950 (N_950,In_809,In_610);
and U951 (N_951,In_846,In_513);
and U952 (N_952,In_134,In_212);
and U953 (N_953,In_659,In_320);
nor U954 (N_954,In_158,In_766);
nand U955 (N_955,In_504,In_372);
or U956 (N_956,In_562,In_679);
and U957 (N_957,In_466,In_579);
nand U958 (N_958,In_276,In_126);
or U959 (N_959,In_926,In_661);
nand U960 (N_960,In_852,In_137);
nor U961 (N_961,In_691,In_173);
and U962 (N_962,In_88,In_806);
or U963 (N_963,In_144,In_912);
or U964 (N_964,In_763,In_383);
nand U965 (N_965,In_361,In_52);
nor U966 (N_966,In_551,In_700);
and U967 (N_967,In_614,In_29);
nor U968 (N_968,In_751,In_218);
nand U969 (N_969,In_755,In_395);
and U970 (N_970,In_118,In_759);
or U971 (N_971,In_361,In_46);
and U972 (N_972,In_338,In_565);
or U973 (N_973,In_319,In_622);
nor U974 (N_974,In_527,In_700);
or U975 (N_975,In_457,In_723);
and U976 (N_976,In_534,In_437);
nor U977 (N_977,In_144,In_532);
nand U978 (N_978,In_593,In_838);
nand U979 (N_979,In_421,In_29);
or U980 (N_980,In_748,In_895);
or U981 (N_981,In_702,In_323);
and U982 (N_982,In_771,In_611);
or U983 (N_983,In_160,In_231);
nand U984 (N_984,In_866,In_959);
or U985 (N_985,In_328,In_211);
nand U986 (N_986,In_161,In_112);
nand U987 (N_987,In_512,In_396);
nor U988 (N_988,In_377,In_708);
nor U989 (N_989,In_545,In_160);
nand U990 (N_990,In_188,In_301);
and U991 (N_991,In_430,In_281);
nor U992 (N_992,In_451,In_200);
nand U993 (N_993,In_483,In_362);
xnor U994 (N_994,In_30,In_891);
nor U995 (N_995,In_533,In_521);
or U996 (N_996,In_447,In_32);
nor U997 (N_997,In_367,In_286);
nor U998 (N_998,In_180,In_25);
nor U999 (N_999,In_657,In_314);
nor U1000 (N_1000,In_891,In_321);
or U1001 (N_1001,In_357,In_676);
nor U1002 (N_1002,In_191,In_994);
nand U1003 (N_1003,In_261,In_589);
nor U1004 (N_1004,In_995,In_830);
nand U1005 (N_1005,In_944,In_147);
nand U1006 (N_1006,In_560,In_64);
and U1007 (N_1007,In_36,In_940);
and U1008 (N_1008,In_313,In_386);
nor U1009 (N_1009,In_764,In_570);
or U1010 (N_1010,In_174,In_836);
nand U1011 (N_1011,In_519,In_126);
nand U1012 (N_1012,In_83,In_804);
or U1013 (N_1013,In_206,In_498);
and U1014 (N_1014,In_170,In_493);
nor U1015 (N_1015,In_850,In_289);
nand U1016 (N_1016,In_414,In_406);
or U1017 (N_1017,In_173,In_937);
or U1018 (N_1018,In_112,In_64);
or U1019 (N_1019,In_913,In_415);
nor U1020 (N_1020,In_342,In_659);
or U1021 (N_1021,In_356,In_443);
and U1022 (N_1022,In_709,In_384);
nor U1023 (N_1023,In_240,In_185);
nand U1024 (N_1024,In_311,In_679);
or U1025 (N_1025,In_505,In_799);
and U1026 (N_1026,In_624,In_465);
and U1027 (N_1027,In_856,In_102);
and U1028 (N_1028,In_778,In_945);
nand U1029 (N_1029,In_92,In_469);
nor U1030 (N_1030,In_339,In_146);
xor U1031 (N_1031,In_285,In_129);
or U1032 (N_1032,In_19,In_649);
or U1033 (N_1033,In_3,In_712);
nor U1034 (N_1034,In_312,In_874);
nand U1035 (N_1035,In_736,In_550);
nor U1036 (N_1036,In_610,In_628);
or U1037 (N_1037,In_17,In_518);
nor U1038 (N_1038,In_97,In_770);
or U1039 (N_1039,In_978,In_588);
nand U1040 (N_1040,In_379,In_216);
and U1041 (N_1041,In_438,In_371);
and U1042 (N_1042,In_472,In_875);
nand U1043 (N_1043,In_103,In_629);
xor U1044 (N_1044,In_976,In_367);
xnor U1045 (N_1045,In_377,In_133);
nor U1046 (N_1046,In_313,In_101);
nor U1047 (N_1047,In_9,In_262);
nor U1048 (N_1048,In_291,In_976);
or U1049 (N_1049,In_324,In_126);
or U1050 (N_1050,In_778,In_104);
or U1051 (N_1051,In_419,In_865);
nor U1052 (N_1052,In_122,In_924);
nor U1053 (N_1053,In_755,In_483);
xor U1054 (N_1054,In_120,In_825);
nor U1055 (N_1055,In_747,In_495);
nand U1056 (N_1056,In_952,In_188);
nand U1057 (N_1057,In_393,In_335);
or U1058 (N_1058,In_910,In_773);
or U1059 (N_1059,In_766,In_687);
or U1060 (N_1060,In_826,In_816);
nand U1061 (N_1061,In_118,In_7);
nor U1062 (N_1062,In_238,In_961);
and U1063 (N_1063,In_69,In_258);
nand U1064 (N_1064,In_378,In_325);
xnor U1065 (N_1065,In_811,In_293);
nor U1066 (N_1066,In_87,In_661);
nand U1067 (N_1067,In_866,In_505);
or U1068 (N_1068,In_144,In_677);
or U1069 (N_1069,In_396,In_619);
nor U1070 (N_1070,In_226,In_314);
and U1071 (N_1071,In_307,In_445);
nand U1072 (N_1072,In_98,In_600);
nand U1073 (N_1073,In_215,In_608);
and U1074 (N_1074,In_353,In_932);
or U1075 (N_1075,In_885,In_99);
nor U1076 (N_1076,In_68,In_239);
nor U1077 (N_1077,In_509,In_109);
xnor U1078 (N_1078,In_210,In_880);
nor U1079 (N_1079,In_942,In_404);
and U1080 (N_1080,In_920,In_723);
and U1081 (N_1081,In_646,In_80);
or U1082 (N_1082,In_949,In_462);
and U1083 (N_1083,In_88,In_573);
nand U1084 (N_1084,In_672,In_793);
or U1085 (N_1085,In_707,In_602);
and U1086 (N_1086,In_58,In_962);
nor U1087 (N_1087,In_364,In_882);
nand U1088 (N_1088,In_825,In_819);
and U1089 (N_1089,In_408,In_200);
nand U1090 (N_1090,In_227,In_871);
and U1091 (N_1091,In_480,In_662);
nand U1092 (N_1092,In_195,In_911);
or U1093 (N_1093,In_305,In_854);
or U1094 (N_1094,In_578,In_93);
or U1095 (N_1095,In_77,In_737);
nor U1096 (N_1096,In_955,In_832);
and U1097 (N_1097,In_242,In_310);
nand U1098 (N_1098,In_419,In_228);
and U1099 (N_1099,In_687,In_542);
and U1100 (N_1100,In_473,In_325);
nor U1101 (N_1101,In_955,In_550);
nor U1102 (N_1102,In_143,In_846);
nand U1103 (N_1103,In_348,In_302);
xor U1104 (N_1104,In_983,In_870);
or U1105 (N_1105,In_563,In_168);
nand U1106 (N_1106,In_970,In_543);
and U1107 (N_1107,In_887,In_130);
or U1108 (N_1108,In_791,In_952);
and U1109 (N_1109,In_681,In_279);
and U1110 (N_1110,In_650,In_138);
nor U1111 (N_1111,In_211,In_138);
xnor U1112 (N_1112,In_73,In_268);
nand U1113 (N_1113,In_578,In_210);
or U1114 (N_1114,In_96,In_567);
and U1115 (N_1115,In_336,In_25);
and U1116 (N_1116,In_547,In_385);
nand U1117 (N_1117,In_742,In_855);
or U1118 (N_1118,In_879,In_678);
nor U1119 (N_1119,In_659,In_727);
or U1120 (N_1120,In_884,In_558);
or U1121 (N_1121,In_74,In_285);
nand U1122 (N_1122,In_0,In_166);
nor U1123 (N_1123,In_599,In_560);
or U1124 (N_1124,In_100,In_601);
nand U1125 (N_1125,In_536,In_941);
nor U1126 (N_1126,In_387,In_853);
nand U1127 (N_1127,In_762,In_836);
nor U1128 (N_1128,In_733,In_742);
nor U1129 (N_1129,In_8,In_243);
or U1130 (N_1130,In_94,In_913);
and U1131 (N_1131,In_251,In_15);
nand U1132 (N_1132,In_645,In_399);
or U1133 (N_1133,In_816,In_914);
nor U1134 (N_1134,In_866,In_363);
xor U1135 (N_1135,In_948,In_382);
nor U1136 (N_1136,In_94,In_761);
nor U1137 (N_1137,In_168,In_554);
xnor U1138 (N_1138,In_41,In_597);
and U1139 (N_1139,In_400,In_42);
nand U1140 (N_1140,In_771,In_32);
nor U1141 (N_1141,In_244,In_937);
or U1142 (N_1142,In_842,In_657);
or U1143 (N_1143,In_995,In_854);
and U1144 (N_1144,In_751,In_639);
or U1145 (N_1145,In_723,In_736);
nand U1146 (N_1146,In_423,In_207);
nor U1147 (N_1147,In_5,In_849);
nor U1148 (N_1148,In_53,In_252);
nand U1149 (N_1149,In_328,In_292);
nand U1150 (N_1150,In_210,In_468);
nand U1151 (N_1151,In_861,In_511);
nor U1152 (N_1152,In_244,In_317);
nor U1153 (N_1153,In_782,In_237);
and U1154 (N_1154,In_601,In_878);
xor U1155 (N_1155,In_984,In_205);
nor U1156 (N_1156,In_632,In_133);
nand U1157 (N_1157,In_739,In_658);
xnor U1158 (N_1158,In_673,In_695);
nand U1159 (N_1159,In_657,In_380);
nor U1160 (N_1160,In_392,In_108);
nor U1161 (N_1161,In_580,In_950);
and U1162 (N_1162,In_829,In_647);
nor U1163 (N_1163,In_868,In_627);
or U1164 (N_1164,In_68,In_495);
nor U1165 (N_1165,In_440,In_335);
nor U1166 (N_1166,In_899,In_816);
or U1167 (N_1167,In_251,In_209);
or U1168 (N_1168,In_969,In_496);
and U1169 (N_1169,In_977,In_508);
nor U1170 (N_1170,In_778,In_80);
nor U1171 (N_1171,In_825,In_349);
or U1172 (N_1172,In_459,In_370);
nand U1173 (N_1173,In_557,In_168);
and U1174 (N_1174,In_785,In_69);
nor U1175 (N_1175,In_170,In_892);
nand U1176 (N_1176,In_321,In_477);
and U1177 (N_1177,In_435,In_545);
and U1178 (N_1178,In_966,In_315);
and U1179 (N_1179,In_30,In_15);
and U1180 (N_1180,In_545,In_703);
and U1181 (N_1181,In_92,In_246);
nand U1182 (N_1182,In_81,In_690);
or U1183 (N_1183,In_504,In_473);
and U1184 (N_1184,In_560,In_377);
or U1185 (N_1185,In_223,In_496);
nand U1186 (N_1186,In_741,In_982);
and U1187 (N_1187,In_59,In_868);
nor U1188 (N_1188,In_926,In_51);
xor U1189 (N_1189,In_886,In_870);
nor U1190 (N_1190,In_291,In_204);
nand U1191 (N_1191,In_173,In_392);
or U1192 (N_1192,In_327,In_716);
and U1193 (N_1193,In_412,In_579);
and U1194 (N_1194,In_247,In_359);
or U1195 (N_1195,In_349,In_173);
nor U1196 (N_1196,In_819,In_782);
xor U1197 (N_1197,In_670,In_345);
nor U1198 (N_1198,In_441,In_398);
and U1199 (N_1199,In_778,In_500);
or U1200 (N_1200,In_382,In_750);
or U1201 (N_1201,In_882,In_201);
nand U1202 (N_1202,In_130,In_566);
nand U1203 (N_1203,In_348,In_61);
or U1204 (N_1204,In_753,In_69);
and U1205 (N_1205,In_721,In_364);
nor U1206 (N_1206,In_511,In_124);
or U1207 (N_1207,In_265,In_534);
nand U1208 (N_1208,In_499,In_360);
nand U1209 (N_1209,In_514,In_826);
nand U1210 (N_1210,In_687,In_154);
xor U1211 (N_1211,In_712,In_240);
nand U1212 (N_1212,In_565,In_435);
and U1213 (N_1213,In_39,In_399);
and U1214 (N_1214,In_344,In_829);
and U1215 (N_1215,In_941,In_723);
nand U1216 (N_1216,In_530,In_518);
nor U1217 (N_1217,In_884,In_388);
and U1218 (N_1218,In_582,In_212);
nand U1219 (N_1219,In_877,In_319);
and U1220 (N_1220,In_478,In_530);
nand U1221 (N_1221,In_37,In_47);
xor U1222 (N_1222,In_980,In_277);
and U1223 (N_1223,In_995,In_912);
nor U1224 (N_1224,In_333,In_433);
and U1225 (N_1225,In_77,In_64);
nand U1226 (N_1226,In_531,In_488);
nand U1227 (N_1227,In_802,In_523);
or U1228 (N_1228,In_22,In_513);
and U1229 (N_1229,In_666,In_501);
nor U1230 (N_1230,In_811,In_438);
nand U1231 (N_1231,In_231,In_462);
nand U1232 (N_1232,In_680,In_577);
xor U1233 (N_1233,In_531,In_752);
nand U1234 (N_1234,In_680,In_214);
and U1235 (N_1235,In_327,In_101);
and U1236 (N_1236,In_303,In_433);
or U1237 (N_1237,In_793,In_389);
or U1238 (N_1238,In_859,In_430);
nor U1239 (N_1239,In_689,In_252);
or U1240 (N_1240,In_784,In_559);
nor U1241 (N_1241,In_620,In_692);
or U1242 (N_1242,In_950,In_303);
nor U1243 (N_1243,In_828,In_808);
nand U1244 (N_1244,In_544,In_567);
or U1245 (N_1245,In_305,In_925);
nand U1246 (N_1246,In_479,In_807);
nand U1247 (N_1247,In_175,In_46);
or U1248 (N_1248,In_720,In_29);
and U1249 (N_1249,In_52,In_55);
nor U1250 (N_1250,In_17,In_199);
nand U1251 (N_1251,In_322,In_208);
nor U1252 (N_1252,In_420,In_613);
nor U1253 (N_1253,In_923,In_878);
nor U1254 (N_1254,In_570,In_168);
or U1255 (N_1255,In_108,In_704);
and U1256 (N_1256,In_19,In_182);
nand U1257 (N_1257,In_994,In_315);
or U1258 (N_1258,In_300,In_611);
and U1259 (N_1259,In_390,In_72);
or U1260 (N_1260,In_742,In_648);
or U1261 (N_1261,In_72,In_790);
nor U1262 (N_1262,In_784,In_477);
nor U1263 (N_1263,In_615,In_855);
and U1264 (N_1264,In_97,In_255);
nor U1265 (N_1265,In_960,In_629);
nor U1266 (N_1266,In_568,In_67);
or U1267 (N_1267,In_892,In_396);
nor U1268 (N_1268,In_933,In_158);
or U1269 (N_1269,In_277,In_400);
nor U1270 (N_1270,In_544,In_360);
and U1271 (N_1271,In_351,In_964);
and U1272 (N_1272,In_550,In_591);
and U1273 (N_1273,In_548,In_761);
and U1274 (N_1274,In_382,In_919);
nand U1275 (N_1275,In_473,In_572);
nand U1276 (N_1276,In_643,In_458);
nand U1277 (N_1277,In_821,In_415);
or U1278 (N_1278,In_520,In_602);
or U1279 (N_1279,In_381,In_443);
nand U1280 (N_1280,In_288,In_528);
or U1281 (N_1281,In_840,In_599);
nor U1282 (N_1282,In_160,In_151);
and U1283 (N_1283,In_50,In_145);
or U1284 (N_1284,In_863,In_494);
or U1285 (N_1285,In_712,In_638);
or U1286 (N_1286,In_610,In_827);
and U1287 (N_1287,In_778,In_419);
or U1288 (N_1288,In_289,In_381);
nand U1289 (N_1289,In_330,In_730);
or U1290 (N_1290,In_45,In_597);
nor U1291 (N_1291,In_439,In_91);
or U1292 (N_1292,In_427,In_111);
nand U1293 (N_1293,In_464,In_569);
nand U1294 (N_1294,In_665,In_180);
nor U1295 (N_1295,In_407,In_375);
nor U1296 (N_1296,In_214,In_18);
or U1297 (N_1297,In_268,In_287);
and U1298 (N_1298,In_690,In_538);
nand U1299 (N_1299,In_127,In_70);
xnor U1300 (N_1300,In_530,In_953);
or U1301 (N_1301,In_750,In_575);
or U1302 (N_1302,In_461,In_605);
nor U1303 (N_1303,In_931,In_552);
and U1304 (N_1304,In_984,In_819);
nor U1305 (N_1305,In_530,In_94);
xnor U1306 (N_1306,In_600,In_187);
or U1307 (N_1307,In_829,In_918);
nand U1308 (N_1308,In_974,In_156);
and U1309 (N_1309,In_322,In_351);
and U1310 (N_1310,In_147,In_938);
or U1311 (N_1311,In_393,In_269);
nand U1312 (N_1312,In_194,In_602);
nor U1313 (N_1313,In_28,In_430);
and U1314 (N_1314,In_195,In_626);
or U1315 (N_1315,In_243,In_33);
nor U1316 (N_1316,In_428,In_126);
nor U1317 (N_1317,In_299,In_810);
and U1318 (N_1318,In_89,In_700);
nor U1319 (N_1319,In_816,In_160);
or U1320 (N_1320,In_754,In_972);
and U1321 (N_1321,In_974,In_949);
nand U1322 (N_1322,In_564,In_459);
nand U1323 (N_1323,In_89,In_656);
or U1324 (N_1324,In_369,In_543);
nor U1325 (N_1325,In_667,In_549);
nand U1326 (N_1326,In_789,In_813);
and U1327 (N_1327,In_563,In_973);
nand U1328 (N_1328,In_439,In_196);
xor U1329 (N_1329,In_804,In_194);
or U1330 (N_1330,In_222,In_200);
nor U1331 (N_1331,In_964,In_10);
nand U1332 (N_1332,In_152,In_183);
xnor U1333 (N_1333,In_699,In_350);
nand U1334 (N_1334,In_826,In_403);
nand U1335 (N_1335,In_723,In_243);
or U1336 (N_1336,In_489,In_758);
nor U1337 (N_1337,In_522,In_801);
nor U1338 (N_1338,In_822,In_167);
or U1339 (N_1339,In_352,In_520);
or U1340 (N_1340,In_596,In_845);
and U1341 (N_1341,In_88,In_395);
nor U1342 (N_1342,In_68,In_735);
nor U1343 (N_1343,In_25,In_136);
or U1344 (N_1344,In_717,In_396);
or U1345 (N_1345,In_751,In_983);
and U1346 (N_1346,In_945,In_403);
nor U1347 (N_1347,In_647,In_599);
and U1348 (N_1348,In_549,In_522);
nor U1349 (N_1349,In_975,In_224);
and U1350 (N_1350,In_950,In_491);
or U1351 (N_1351,In_507,In_94);
nor U1352 (N_1352,In_375,In_828);
and U1353 (N_1353,In_571,In_249);
nand U1354 (N_1354,In_45,In_131);
nor U1355 (N_1355,In_920,In_713);
or U1356 (N_1356,In_897,In_721);
nor U1357 (N_1357,In_712,In_693);
and U1358 (N_1358,In_396,In_383);
nor U1359 (N_1359,In_761,In_926);
and U1360 (N_1360,In_969,In_388);
nand U1361 (N_1361,In_477,In_936);
nand U1362 (N_1362,In_81,In_152);
nor U1363 (N_1363,In_689,In_418);
nor U1364 (N_1364,In_667,In_903);
and U1365 (N_1365,In_401,In_999);
and U1366 (N_1366,In_964,In_458);
and U1367 (N_1367,In_591,In_120);
or U1368 (N_1368,In_296,In_949);
or U1369 (N_1369,In_681,In_571);
nand U1370 (N_1370,In_649,In_806);
and U1371 (N_1371,In_740,In_570);
nor U1372 (N_1372,In_173,In_955);
nand U1373 (N_1373,In_431,In_736);
or U1374 (N_1374,In_589,In_472);
nand U1375 (N_1375,In_206,In_688);
and U1376 (N_1376,In_817,In_601);
and U1377 (N_1377,In_715,In_571);
or U1378 (N_1378,In_378,In_380);
nand U1379 (N_1379,In_474,In_642);
nor U1380 (N_1380,In_511,In_958);
or U1381 (N_1381,In_188,In_821);
nor U1382 (N_1382,In_615,In_340);
nand U1383 (N_1383,In_466,In_432);
nor U1384 (N_1384,In_629,In_372);
or U1385 (N_1385,In_176,In_793);
nand U1386 (N_1386,In_399,In_16);
or U1387 (N_1387,In_187,In_502);
and U1388 (N_1388,In_256,In_547);
nand U1389 (N_1389,In_579,In_441);
or U1390 (N_1390,In_77,In_305);
and U1391 (N_1391,In_822,In_515);
nor U1392 (N_1392,In_301,In_258);
and U1393 (N_1393,In_931,In_973);
nand U1394 (N_1394,In_957,In_147);
and U1395 (N_1395,In_805,In_389);
and U1396 (N_1396,In_524,In_395);
nor U1397 (N_1397,In_903,In_784);
nand U1398 (N_1398,In_47,In_540);
and U1399 (N_1399,In_70,In_130);
and U1400 (N_1400,In_739,In_12);
or U1401 (N_1401,In_917,In_934);
nand U1402 (N_1402,In_275,In_202);
or U1403 (N_1403,In_310,In_931);
nand U1404 (N_1404,In_704,In_830);
xor U1405 (N_1405,In_384,In_568);
and U1406 (N_1406,In_728,In_982);
nor U1407 (N_1407,In_938,In_373);
nor U1408 (N_1408,In_655,In_137);
xor U1409 (N_1409,In_43,In_804);
and U1410 (N_1410,In_358,In_227);
nor U1411 (N_1411,In_935,In_2);
xor U1412 (N_1412,In_150,In_810);
xor U1413 (N_1413,In_348,In_287);
nor U1414 (N_1414,In_505,In_374);
nand U1415 (N_1415,In_239,In_894);
nand U1416 (N_1416,In_370,In_968);
and U1417 (N_1417,In_18,In_765);
or U1418 (N_1418,In_748,In_843);
nand U1419 (N_1419,In_214,In_788);
or U1420 (N_1420,In_578,In_214);
nor U1421 (N_1421,In_458,In_411);
or U1422 (N_1422,In_536,In_241);
and U1423 (N_1423,In_538,In_44);
nand U1424 (N_1424,In_274,In_317);
nor U1425 (N_1425,In_917,In_154);
nand U1426 (N_1426,In_498,In_675);
or U1427 (N_1427,In_138,In_917);
nand U1428 (N_1428,In_844,In_478);
and U1429 (N_1429,In_532,In_977);
nor U1430 (N_1430,In_418,In_348);
or U1431 (N_1431,In_384,In_323);
and U1432 (N_1432,In_636,In_617);
nand U1433 (N_1433,In_101,In_424);
and U1434 (N_1434,In_137,In_907);
nand U1435 (N_1435,In_337,In_699);
or U1436 (N_1436,In_28,In_897);
and U1437 (N_1437,In_815,In_136);
and U1438 (N_1438,In_343,In_532);
and U1439 (N_1439,In_541,In_710);
xnor U1440 (N_1440,In_509,In_871);
or U1441 (N_1441,In_714,In_979);
nor U1442 (N_1442,In_752,In_475);
and U1443 (N_1443,In_577,In_61);
nor U1444 (N_1444,In_632,In_80);
nand U1445 (N_1445,In_357,In_483);
or U1446 (N_1446,In_159,In_982);
nand U1447 (N_1447,In_336,In_823);
nor U1448 (N_1448,In_207,In_389);
nand U1449 (N_1449,In_988,In_735);
nand U1450 (N_1450,In_169,In_195);
nand U1451 (N_1451,In_584,In_301);
or U1452 (N_1452,In_971,In_854);
or U1453 (N_1453,In_135,In_79);
and U1454 (N_1454,In_498,In_716);
nand U1455 (N_1455,In_400,In_266);
nand U1456 (N_1456,In_897,In_566);
nor U1457 (N_1457,In_151,In_454);
nand U1458 (N_1458,In_670,In_7);
and U1459 (N_1459,In_787,In_860);
nand U1460 (N_1460,In_606,In_536);
and U1461 (N_1461,In_566,In_721);
or U1462 (N_1462,In_917,In_317);
nor U1463 (N_1463,In_326,In_682);
nor U1464 (N_1464,In_719,In_548);
or U1465 (N_1465,In_676,In_252);
and U1466 (N_1466,In_342,In_467);
and U1467 (N_1467,In_2,In_290);
nor U1468 (N_1468,In_81,In_320);
nor U1469 (N_1469,In_368,In_160);
or U1470 (N_1470,In_443,In_883);
or U1471 (N_1471,In_259,In_986);
nor U1472 (N_1472,In_499,In_425);
nor U1473 (N_1473,In_941,In_889);
nor U1474 (N_1474,In_10,In_930);
and U1475 (N_1475,In_842,In_75);
and U1476 (N_1476,In_402,In_710);
nor U1477 (N_1477,In_788,In_284);
nand U1478 (N_1478,In_638,In_778);
and U1479 (N_1479,In_967,In_30);
or U1480 (N_1480,In_287,In_578);
or U1481 (N_1481,In_216,In_373);
nand U1482 (N_1482,In_285,In_339);
or U1483 (N_1483,In_315,In_730);
or U1484 (N_1484,In_234,In_702);
and U1485 (N_1485,In_891,In_611);
or U1486 (N_1486,In_182,In_171);
or U1487 (N_1487,In_195,In_527);
nand U1488 (N_1488,In_253,In_858);
nor U1489 (N_1489,In_708,In_23);
nand U1490 (N_1490,In_839,In_326);
or U1491 (N_1491,In_810,In_371);
nor U1492 (N_1492,In_917,In_235);
and U1493 (N_1493,In_119,In_582);
and U1494 (N_1494,In_304,In_355);
nor U1495 (N_1495,In_189,In_738);
nand U1496 (N_1496,In_209,In_167);
or U1497 (N_1497,In_333,In_223);
and U1498 (N_1498,In_37,In_140);
nand U1499 (N_1499,In_193,In_976);
nor U1500 (N_1500,In_224,In_771);
nand U1501 (N_1501,In_515,In_280);
and U1502 (N_1502,In_259,In_66);
nand U1503 (N_1503,In_669,In_929);
nor U1504 (N_1504,In_876,In_329);
or U1505 (N_1505,In_580,In_470);
nor U1506 (N_1506,In_88,In_407);
or U1507 (N_1507,In_182,In_908);
nor U1508 (N_1508,In_786,In_415);
or U1509 (N_1509,In_982,In_538);
nand U1510 (N_1510,In_859,In_491);
and U1511 (N_1511,In_229,In_891);
or U1512 (N_1512,In_693,In_939);
nand U1513 (N_1513,In_103,In_995);
nor U1514 (N_1514,In_17,In_775);
nor U1515 (N_1515,In_409,In_255);
or U1516 (N_1516,In_668,In_31);
and U1517 (N_1517,In_414,In_711);
nor U1518 (N_1518,In_527,In_703);
or U1519 (N_1519,In_922,In_946);
nand U1520 (N_1520,In_112,In_875);
nor U1521 (N_1521,In_543,In_702);
and U1522 (N_1522,In_417,In_109);
nand U1523 (N_1523,In_220,In_265);
and U1524 (N_1524,In_783,In_547);
or U1525 (N_1525,In_555,In_695);
and U1526 (N_1526,In_791,In_36);
nand U1527 (N_1527,In_893,In_924);
nor U1528 (N_1528,In_251,In_338);
or U1529 (N_1529,In_751,In_103);
or U1530 (N_1530,In_864,In_125);
or U1531 (N_1531,In_24,In_609);
xor U1532 (N_1532,In_465,In_719);
nor U1533 (N_1533,In_837,In_598);
or U1534 (N_1534,In_136,In_105);
nor U1535 (N_1535,In_881,In_981);
or U1536 (N_1536,In_127,In_540);
nand U1537 (N_1537,In_67,In_708);
nor U1538 (N_1538,In_202,In_437);
nand U1539 (N_1539,In_361,In_104);
and U1540 (N_1540,In_918,In_324);
nand U1541 (N_1541,In_75,In_338);
or U1542 (N_1542,In_304,In_383);
and U1543 (N_1543,In_238,In_71);
or U1544 (N_1544,In_322,In_607);
and U1545 (N_1545,In_193,In_263);
nand U1546 (N_1546,In_210,In_660);
and U1547 (N_1547,In_579,In_999);
or U1548 (N_1548,In_318,In_843);
or U1549 (N_1549,In_60,In_319);
nor U1550 (N_1550,In_964,In_309);
nor U1551 (N_1551,In_318,In_458);
and U1552 (N_1552,In_828,In_504);
nand U1553 (N_1553,In_712,In_475);
nor U1554 (N_1554,In_456,In_553);
nand U1555 (N_1555,In_291,In_942);
nor U1556 (N_1556,In_691,In_73);
and U1557 (N_1557,In_672,In_214);
or U1558 (N_1558,In_358,In_182);
and U1559 (N_1559,In_859,In_896);
or U1560 (N_1560,In_943,In_206);
nor U1561 (N_1561,In_474,In_274);
nor U1562 (N_1562,In_589,In_184);
nand U1563 (N_1563,In_194,In_891);
xor U1564 (N_1564,In_62,In_841);
nor U1565 (N_1565,In_459,In_599);
and U1566 (N_1566,In_322,In_154);
nor U1567 (N_1567,In_135,In_644);
and U1568 (N_1568,In_27,In_268);
nor U1569 (N_1569,In_270,In_877);
and U1570 (N_1570,In_357,In_994);
and U1571 (N_1571,In_721,In_452);
or U1572 (N_1572,In_843,In_820);
nor U1573 (N_1573,In_44,In_157);
or U1574 (N_1574,In_52,In_854);
nor U1575 (N_1575,In_275,In_850);
or U1576 (N_1576,In_664,In_884);
or U1577 (N_1577,In_107,In_778);
nand U1578 (N_1578,In_247,In_992);
nor U1579 (N_1579,In_810,In_696);
nor U1580 (N_1580,In_538,In_257);
and U1581 (N_1581,In_675,In_294);
and U1582 (N_1582,In_286,In_490);
or U1583 (N_1583,In_131,In_882);
nand U1584 (N_1584,In_877,In_344);
and U1585 (N_1585,In_872,In_805);
and U1586 (N_1586,In_944,In_529);
nor U1587 (N_1587,In_588,In_554);
nor U1588 (N_1588,In_498,In_260);
and U1589 (N_1589,In_991,In_500);
or U1590 (N_1590,In_518,In_581);
and U1591 (N_1591,In_875,In_750);
or U1592 (N_1592,In_927,In_47);
nor U1593 (N_1593,In_982,In_425);
or U1594 (N_1594,In_33,In_253);
nor U1595 (N_1595,In_5,In_595);
or U1596 (N_1596,In_722,In_944);
nor U1597 (N_1597,In_450,In_524);
nor U1598 (N_1598,In_797,In_580);
xor U1599 (N_1599,In_904,In_924);
and U1600 (N_1600,In_552,In_38);
or U1601 (N_1601,In_483,In_986);
xnor U1602 (N_1602,In_49,In_972);
nand U1603 (N_1603,In_773,In_911);
and U1604 (N_1604,In_339,In_227);
or U1605 (N_1605,In_524,In_284);
nand U1606 (N_1606,In_745,In_272);
and U1607 (N_1607,In_95,In_341);
or U1608 (N_1608,In_787,In_69);
or U1609 (N_1609,In_820,In_224);
nand U1610 (N_1610,In_576,In_64);
nor U1611 (N_1611,In_76,In_337);
nand U1612 (N_1612,In_157,In_408);
nand U1613 (N_1613,In_822,In_165);
nor U1614 (N_1614,In_129,In_367);
nor U1615 (N_1615,In_435,In_939);
xor U1616 (N_1616,In_45,In_481);
nand U1617 (N_1617,In_521,In_907);
or U1618 (N_1618,In_687,In_704);
nand U1619 (N_1619,In_692,In_241);
nand U1620 (N_1620,In_610,In_463);
nand U1621 (N_1621,In_49,In_604);
and U1622 (N_1622,In_904,In_997);
and U1623 (N_1623,In_417,In_788);
or U1624 (N_1624,In_318,In_874);
nand U1625 (N_1625,In_37,In_477);
nand U1626 (N_1626,In_908,In_512);
nor U1627 (N_1627,In_810,In_576);
or U1628 (N_1628,In_277,In_386);
nor U1629 (N_1629,In_552,In_10);
nor U1630 (N_1630,In_213,In_100);
or U1631 (N_1631,In_340,In_512);
and U1632 (N_1632,In_595,In_150);
nand U1633 (N_1633,In_261,In_78);
nor U1634 (N_1634,In_863,In_59);
nor U1635 (N_1635,In_413,In_404);
and U1636 (N_1636,In_223,In_355);
nand U1637 (N_1637,In_884,In_16);
nor U1638 (N_1638,In_123,In_961);
xnor U1639 (N_1639,In_253,In_269);
and U1640 (N_1640,In_635,In_874);
xor U1641 (N_1641,In_261,In_336);
or U1642 (N_1642,In_248,In_91);
nand U1643 (N_1643,In_802,In_147);
or U1644 (N_1644,In_723,In_365);
nand U1645 (N_1645,In_841,In_683);
or U1646 (N_1646,In_888,In_965);
nand U1647 (N_1647,In_620,In_899);
and U1648 (N_1648,In_678,In_462);
nor U1649 (N_1649,In_848,In_144);
and U1650 (N_1650,In_67,In_580);
nor U1651 (N_1651,In_873,In_186);
xor U1652 (N_1652,In_199,In_381);
or U1653 (N_1653,In_906,In_370);
nor U1654 (N_1654,In_489,In_281);
nand U1655 (N_1655,In_360,In_283);
or U1656 (N_1656,In_471,In_667);
and U1657 (N_1657,In_222,In_780);
and U1658 (N_1658,In_741,In_105);
nor U1659 (N_1659,In_775,In_481);
xor U1660 (N_1660,In_502,In_636);
nor U1661 (N_1661,In_32,In_824);
xnor U1662 (N_1662,In_843,In_929);
nand U1663 (N_1663,In_379,In_942);
nor U1664 (N_1664,In_168,In_20);
and U1665 (N_1665,In_876,In_195);
or U1666 (N_1666,In_103,In_643);
or U1667 (N_1667,In_407,In_531);
nor U1668 (N_1668,In_678,In_670);
nor U1669 (N_1669,In_289,In_319);
or U1670 (N_1670,In_480,In_873);
nor U1671 (N_1671,In_803,In_996);
and U1672 (N_1672,In_445,In_203);
or U1673 (N_1673,In_618,In_593);
nand U1674 (N_1674,In_204,In_270);
and U1675 (N_1675,In_862,In_240);
and U1676 (N_1676,In_564,In_301);
xor U1677 (N_1677,In_594,In_685);
nand U1678 (N_1678,In_23,In_958);
and U1679 (N_1679,In_571,In_382);
and U1680 (N_1680,In_187,In_35);
and U1681 (N_1681,In_913,In_977);
and U1682 (N_1682,In_726,In_260);
nor U1683 (N_1683,In_323,In_986);
or U1684 (N_1684,In_744,In_366);
and U1685 (N_1685,In_958,In_680);
or U1686 (N_1686,In_274,In_797);
nand U1687 (N_1687,In_46,In_187);
and U1688 (N_1688,In_838,In_658);
and U1689 (N_1689,In_342,In_751);
or U1690 (N_1690,In_169,In_93);
nor U1691 (N_1691,In_135,In_174);
nand U1692 (N_1692,In_381,In_303);
nor U1693 (N_1693,In_70,In_252);
nand U1694 (N_1694,In_12,In_112);
or U1695 (N_1695,In_588,In_30);
nor U1696 (N_1696,In_371,In_271);
nand U1697 (N_1697,In_310,In_437);
nand U1698 (N_1698,In_990,In_282);
or U1699 (N_1699,In_952,In_79);
and U1700 (N_1700,In_702,In_315);
and U1701 (N_1701,In_818,In_993);
nor U1702 (N_1702,In_86,In_824);
or U1703 (N_1703,In_489,In_307);
nor U1704 (N_1704,In_28,In_526);
or U1705 (N_1705,In_168,In_269);
nand U1706 (N_1706,In_244,In_800);
or U1707 (N_1707,In_209,In_731);
nor U1708 (N_1708,In_608,In_258);
or U1709 (N_1709,In_298,In_562);
nor U1710 (N_1710,In_764,In_800);
nand U1711 (N_1711,In_41,In_884);
or U1712 (N_1712,In_165,In_349);
nor U1713 (N_1713,In_325,In_15);
xnor U1714 (N_1714,In_54,In_395);
nand U1715 (N_1715,In_34,In_219);
and U1716 (N_1716,In_610,In_812);
or U1717 (N_1717,In_688,In_436);
nor U1718 (N_1718,In_327,In_640);
or U1719 (N_1719,In_26,In_919);
nor U1720 (N_1720,In_809,In_631);
or U1721 (N_1721,In_142,In_938);
nand U1722 (N_1722,In_884,In_382);
xor U1723 (N_1723,In_602,In_91);
or U1724 (N_1724,In_213,In_725);
and U1725 (N_1725,In_52,In_82);
and U1726 (N_1726,In_986,In_268);
and U1727 (N_1727,In_64,In_318);
or U1728 (N_1728,In_162,In_806);
nor U1729 (N_1729,In_54,In_461);
nand U1730 (N_1730,In_602,In_268);
nand U1731 (N_1731,In_579,In_781);
xor U1732 (N_1732,In_888,In_786);
nor U1733 (N_1733,In_683,In_305);
or U1734 (N_1734,In_524,In_289);
and U1735 (N_1735,In_104,In_791);
and U1736 (N_1736,In_99,In_77);
nor U1737 (N_1737,In_408,In_197);
nor U1738 (N_1738,In_612,In_881);
nor U1739 (N_1739,In_235,In_926);
nand U1740 (N_1740,In_308,In_355);
nand U1741 (N_1741,In_792,In_216);
nand U1742 (N_1742,In_653,In_770);
nand U1743 (N_1743,In_335,In_552);
nand U1744 (N_1744,In_910,In_393);
or U1745 (N_1745,In_695,In_13);
or U1746 (N_1746,In_819,In_472);
nor U1747 (N_1747,In_851,In_473);
and U1748 (N_1748,In_254,In_308);
and U1749 (N_1749,In_961,In_785);
nor U1750 (N_1750,In_402,In_465);
or U1751 (N_1751,In_571,In_456);
and U1752 (N_1752,In_82,In_357);
and U1753 (N_1753,In_35,In_156);
or U1754 (N_1754,In_543,In_161);
or U1755 (N_1755,In_967,In_449);
nand U1756 (N_1756,In_891,In_861);
nor U1757 (N_1757,In_921,In_542);
nor U1758 (N_1758,In_876,In_523);
or U1759 (N_1759,In_120,In_720);
or U1760 (N_1760,In_428,In_732);
or U1761 (N_1761,In_582,In_970);
nand U1762 (N_1762,In_552,In_163);
nand U1763 (N_1763,In_911,In_517);
or U1764 (N_1764,In_833,In_660);
or U1765 (N_1765,In_618,In_368);
and U1766 (N_1766,In_709,In_609);
or U1767 (N_1767,In_63,In_509);
and U1768 (N_1768,In_786,In_267);
and U1769 (N_1769,In_500,In_249);
nand U1770 (N_1770,In_385,In_931);
nand U1771 (N_1771,In_793,In_746);
xnor U1772 (N_1772,In_846,In_535);
and U1773 (N_1773,In_2,In_26);
nand U1774 (N_1774,In_12,In_404);
and U1775 (N_1775,In_209,In_249);
or U1776 (N_1776,In_119,In_737);
xnor U1777 (N_1777,In_771,In_253);
or U1778 (N_1778,In_943,In_873);
or U1779 (N_1779,In_425,In_372);
nand U1780 (N_1780,In_250,In_147);
and U1781 (N_1781,In_665,In_449);
nor U1782 (N_1782,In_55,In_229);
and U1783 (N_1783,In_662,In_206);
nor U1784 (N_1784,In_852,In_838);
and U1785 (N_1785,In_175,In_827);
nor U1786 (N_1786,In_960,In_596);
nor U1787 (N_1787,In_604,In_811);
or U1788 (N_1788,In_55,In_634);
or U1789 (N_1789,In_614,In_492);
nand U1790 (N_1790,In_251,In_608);
or U1791 (N_1791,In_367,In_121);
and U1792 (N_1792,In_505,In_346);
and U1793 (N_1793,In_948,In_887);
nand U1794 (N_1794,In_470,In_316);
and U1795 (N_1795,In_530,In_713);
nor U1796 (N_1796,In_214,In_330);
nor U1797 (N_1797,In_292,In_504);
or U1798 (N_1798,In_250,In_222);
nor U1799 (N_1799,In_789,In_926);
nor U1800 (N_1800,In_486,In_140);
or U1801 (N_1801,In_847,In_848);
or U1802 (N_1802,In_761,In_993);
nand U1803 (N_1803,In_740,In_458);
nand U1804 (N_1804,In_336,In_779);
xnor U1805 (N_1805,In_96,In_471);
nor U1806 (N_1806,In_455,In_156);
or U1807 (N_1807,In_148,In_973);
nor U1808 (N_1808,In_895,In_375);
or U1809 (N_1809,In_594,In_61);
or U1810 (N_1810,In_133,In_32);
xor U1811 (N_1811,In_879,In_134);
and U1812 (N_1812,In_249,In_856);
nand U1813 (N_1813,In_898,In_25);
or U1814 (N_1814,In_180,In_190);
nor U1815 (N_1815,In_409,In_103);
nor U1816 (N_1816,In_743,In_692);
and U1817 (N_1817,In_449,In_119);
nor U1818 (N_1818,In_588,In_234);
or U1819 (N_1819,In_882,In_927);
or U1820 (N_1820,In_901,In_309);
nand U1821 (N_1821,In_675,In_595);
nand U1822 (N_1822,In_504,In_60);
nor U1823 (N_1823,In_379,In_784);
nor U1824 (N_1824,In_788,In_305);
nor U1825 (N_1825,In_415,In_652);
and U1826 (N_1826,In_514,In_946);
nand U1827 (N_1827,In_131,In_403);
nand U1828 (N_1828,In_16,In_536);
or U1829 (N_1829,In_224,In_82);
or U1830 (N_1830,In_135,In_992);
nor U1831 (N_1831,In_831,In_472);
nand U1832 (N_1832,In_595,In_418);
and U1833 (N_1833,In_818,In_586);
or U1834 (N_1834,In_814,In_775);
and U1835 (N_1835,In_380,In_944);
or U1836 (N_1836,In_876,In_242);
or U1837 (N_1837,In_540,In_586);
or U1838 (N_1838,In_501,In_277);
nor U1839 (N_1839,In_357,In_921);
and U1840 (N_1840,In_214,In_785);
or U1841 (N_1841,In_338,In_355);
xor U1842 (N_1842,In_194,In_137);
nand U1843 (N_1843,In_91,In_881);
or U1844 (N_1844,In_642,In_568);
nand U1845 (N_1845,In_43,In_328);
nor U1846 (N_1846,In_369,In_829);
nand U1847 (N_1847,In_934,In_137);
nor U1848 (N_1848,In_122,In_196);
and U1849 (N_1849,In_57,In_225);
xor U1850 (N_1850,In_195,In_570);
and U1851 (N_1851,In_432,In_476);
or U1852 (N_1852,In_177,In_2);
nor U1853 (N_1853,In_91,In_250);
nor U1854 (N_1854,In_962,In_931);
or U1855 (N_1855,In_749,In_232);
nand U1856 (N_1856,In_433,In_479);
nand U1857 (N_1857,In_269,In_997);
nand U1858 (N_1858,In_815,In_631);
or U1859 (N_1859,In_152,In_642);
nor U1860 (N_1860,In_732,In_440);
and U1861 (N_1861,In_209,In_203);
nand U1862 (N_1862,In_768,In_126);
and U1863 (N_1863,In_259,In_604);
and U1864 (N_1864,In_3,In_15);
or U1865 (N_1865,In_455,In_316);
or U1866 (N_1866,In_356,In_76);
and U1867 (N_1867,In_316,In_591);
nor U1868 (N_1868,In_596,In_356);
and U1869 (N_1869,In_937,In_880);
or U1870 (N_1870,In_370,In_978);
and U1871 (N_1871,In_994,In_853);
xnor U1872 (N_1872,In_204,In_484);
and U1873 (N_1873,In_823,In_410);
nor U1874 (N_1874,In_870,In_285);
or U1875 (N_1875,In_865,In_200);
nand U1876 (N_1876,In_476,In_564);
and U1877 (N_1877,In_838,In_606);
nand U1878 (N_1878,In_519,In_820);
nand U1879 (N_1879,In_122,In_850);
nor U1880 (N_1880,In_520,In_937);
and U1881 (N_1881,In_453,In_244);
or U1882 (N_1882,In_542,In_955);
nor U1883 (N_1883,In_313,In_319);
or U1884 (N_1884,In_558,In_920);
nand U1885 (N_1885,In_271,In_924);
or U1886 (N_1886,In_122,In_516);
nand U1887 (N_1887,In_65,In_434);
and U1888 (N_1888,In_437,In_518);
or U1889 (N_1889,In_423,In_934);
nor U1890 (N_1890,In_187,In_901);
or U1891 (N_1891,In_341,In_265);
or U1892 (N_1892,In_805,In_636);
nand U1893 (N_1893,In_208,In_247);
nand U1894 (N_1894,In_856,In_419);
nor U1895 (N_1895,In_232,In_867);
and U1896 (N_1896,In_72,In_766);
xor U1897 (N_1897,In_828,In_224);
or U1898 (N_1898,In_35,In_7);
nand U1899 (N_1899,In_775,In_713);
nor U1900 (N_1900,In_965,In_347);
nor U1901 (N_1901,In_493,In_549);
or U1902 (N_1902,In_978,In_192);
nand U1903 (N_1903,In_734,In_212);
or U1904 (N_1904,In_336,In_193);
nor U1905 (N_1905,In_8,In_278);
nand U1906 (N_1906,In_306,In_721);
or U1907 (N_1907,In_375,In_19);
and U1908 (N_1908,In_970,In_438);
nor U1909 (N_1909,In_805,In_622);
nor U1910 (N_1910,In_304,In_399);
nor U1911 (N_1911,In_511,In_554);
and U1912 (N_1912,In_675,In_185);
nor U1913 (N_1913,In_737,In_805);
or U1914 (N_1914,In_66,In_565);
nor U1915 (N_1915,In_96,In_407);
and U1916 (N_1916,In_422,In_467);
nand U1917 (N_1917,In_495,In_599);
nand U1918 (N_1918,In_49,In_372);
or U1919 (N_1919,In_626,In_526);
nand U1920 (N_1920,In_370,In_523);
nor U1921 (N_1921,In_512,In_9);
and U1922 (N_1922,In_891,In_95);
nand U1923 (N_1923,In_609,In_870);
nor U1924 (N_1924,In_981,In_557);
nand U1925 (N_1925,In_163,In_614);
or U1926 (N_1926,In_671,In_121);
and U1927 (N_1927,In_959,In_384);
nand U1928 (N_1928,In_920,In_987);
and U1929 (N_1929,In_582,In_239);
and U1930 (N_1930,In_941,In_319);
or U1931 (N_1931,In_688,In_788);
or U1932 (N_1932,In_581,In_34);
nor U1933 (N_1933,In_40,In_341);
nor U1934 (N_1934,In_98,In_398);
and U1935 (N_1935,In_340,In_965);
or U1936 (N_1936,In_167,In_328);
nor U1937 (N_1937,In_129,In_964);
or U1938 (N_1938,In_223,In_721);
nand U1939 (N_1939,In_607,In_653);
nor U1940 (N_1940,In_607,In_841);
and U1941 (N_1941,In_297,In_433);
and U1942 (N_1942,In_603,In_690);
or U1943 (N_1943,In_583,In_390);
and U1944 (N_1944,In_793,In_95);
nand U1945 (N_1945,In_670,In_289);
and U1946 (N_1946,In_310,In_444);
nor U1947 (N_1947,In_80,In_148);
or U1948 (N_1948,In_461,In_962);
or U1949 (N_1949,In_515,In_306);
nor U1950 (N_1950,In_397,In_179);
and U1951 (N_1951,In_96,In_132);
and U1952 (N_1952,In_986,In_977);
and U1953 (N_1953,In_522,In_989);
and U1954 (N_1954,In_862,In_813);
nand U1955 (N_1955,In_47,In_911);
and U1956 (N_1956,In_826,In_773);
nand U1957 (N_1957,In_514,In_589);
nand U1958 (N_1958,In_418,In_652);
nor U1959 (N_1959,In_181,In_995);
and U1960 (N_1960,In_643,In_92);
and U1961 (N_1961,In_306,In_981);
nor U1962 (N_1962,In_57,In_354);
or U1963 (N_1963,In_735,In_2);
or U1964 (N_1964,In_873,In_590);
and U1965 (N_1965,In_937,In_102);
or U1966 (N_1966,In_81,In_898);
nor U1967 (N_1967,In_968,In_332);
or U1968 (N_1968,In_988,In_929);
nor U1969 (N_1969,In_153,In_832);
nand U1970 (N_1970,In_615,In_378);
and U1971 (N_1971,In_305,In_137);
nor U1972 (N_1972,In_377,In_371);
or U1973 (N_1973,In_847,In_487);
and U1974 (N_1974,In_687,In_696);
and U1975 (N_1975,In_22,In_178);
or U1976 (N_1976,In_188,In_48);
or U1977 (N_1977,In_304,In_662);
nand U1978 (N_1978,In_77,In_430);
nor U1979 (N_1979,In_803,In_417);
and U1980 (N_1980,In_901,In_483);
and U1981 (N_1981,In_661,In_686);
or U1982 (N_1982,In_551,In_468);
nand U1983 (N_1983,In_339,In_368);
xor U1984 (N_1984,In_671,In_652);
nand U1985 (N_1985,In_305,In_159);
and U1986 (N_1986,In_345,In_371);
nor U1987 (N_1987,In_554,In_339);
xnor U1988 (N_1988,In_839,In_437);
or U1989 (N_1989,In_663,In_307);
nand U1990 (N_1990,In_226,In_156);
nor U1991 (N_1991,In_789,In_796);
nand U1992 (N_1992,In_952,In_75);
or U1993 (N_1993,In_640,In_274);
nand U1994 (N_1994,In_246,In_474);
nor U1995 (N_1995,In_839,In_3);
or U1996 (N_1996,In_908,In_681);
or U1997 (N_1997,In_658,In_774);
and U1998 (N_1998,In_924,In_415);
nor U1999 (N_1999,In_958,In_16);
nor U2000 (N_2000,In_264,In_333);
and U2001 (N_2001,In_895,In_33);
or U2002 (N_2002,In_994,In_961);
xor U2003 (N_2003,In_277,In_410);
and U2004 (N_2004,In_167,In_937);
nand U2005 (N_2005,In_141,In_29);
nand U2006 (N_2006,In_50,In_162);
nor U2007 (N_2007,In_337,In_490);
and U2008 (N_2008,In_68,In_595);
and U2009 (N_2009,In_183,In_794);
and U2010 (N_2010,In_66,In_905);
and U2011 (N_2011,In_464,In_489);
and U2012 (N_2012,In_60,In_11);
or U2013 (N_2013,In_178,In_459);
or U2014 (N_2014,In_32,In_163);
nor U2015 (N_2015,In_295,In_879);
and U2016 (N_2016,In_468,In_397);
nand U2017 (N_2017,In_365,In_928);
or U2018 (N_2018,In_683,In_230);
nand U2019 (N_2019,In_989,In_642);
nand U2020 (N_2020,In_754,In_171);
nor U2021 (N_2021,In_842,In_542);
nor U2022 (N_2022,In_486,In_274);
nor U2023 (N_2023,In_278,In_324);
nand U2024 (N_2024,In_666,In_820);
or U2025 (N_2025,In_863,In_80);
nor U2026 (N_2026,In_769,In_979);
or U2027 (N_2027,In_476,In_799);
nand U2028 (N_2028,In_18,In_252);
nand U2029 (N_2029,In_698,In_10);
nor U2030 (N_2030,In_109,In_188);
and U2031 (N_2031,In_127,In_49);
nand U2032 (N_2032,In_206,In_873);
nor U2033 (N_2033,In_736,In_935);
or U2034 (N_2034,In_682,In_670);
nand U2035 (N_2035,In_383,In_661);
nor U2036 (N_2036,In_126,In_695);
nand U2037 (N_2037,In_941,In_821);
or U2038 (N_2038,In_871,In_222);
or U2039 (N_2039,In_452,In_966);
or U2040 (N_2040,In_748,In_394);
nor U2041 (N_2041,In_286,In_408);
nand U2042 (N_2042,In_5,In_399);
nand U2043 (N_2043,In_177,In_925);
nand U2044 (N_2044,In_94,In_84);
nor U2045 (N_2045,In_725,In_460);
nor U2046 (N_2046,In_690,In_704);
or U2047 (N_2047,In_109,In_232);
nand U2048 (N_2048,In_103,In_477);
and U2049 (N_2049,In_859,In_433);
nand U2050 (N_2050,In_870,In_945);
or U2051 (N_2051,In_573,In_874);
nor U2052 (N_2052,In_624,In_818);
nor U2053 (N_2053,In_268,In_508);
nor U2054 (N_2054,In_151,In_746);
nor U2055 (N_2055,In_202,In_768);
or U2056 (N_2056,In_251,In_773);
nor U2057 (N_2057,In_214,In_875);
nand U2058 (N_2058,In_548,In_332);
nor U2059 (N_2059,In_675,In_950);
and U2060 (N_2060,In_728,In_787);
or U2061 (N_2061,In_711,In_223);
nand U2062 (N_2062,In_580,In_520);
or U2063 (N_2063,In_219,In_572);
or U2064 (N_2064,In_481,In_445);
nand U2065 (N_2065,In_301,In_778);
nor U2066 (N_2066,In_857,In_278);
or U2067 (N_2067,In_198,In_996);
nor U2068 (N_2068,In_735,In_63);
nand U2069 (N_2069,In_829,In_705);
or U2070 (N_2070,In_642,In_970);
nand U2071 (N_2071,In_223,In_224);
and U2072 (N_2072,In_380,In_219);
or U2073 (N_2073,In_924,In_283);
nand U2074 (N_2074,In_234,In_317);
or U2075 (N_2075,In_705,In_140);
nand U2076 (N_2076,In_194,In_704);
and U2077 (N_2077,In_95,In_358);
nand U2078 (N_2078,In_855,In_457);
or U2079 (N_2079,In_658,In_779);
or U2080 (N_2080,In_837,In_618);
nand U2081 (N_2081,In_42,In_911);
nor U2082 (N_2082,In_168,In_825);
nor U2083 (N_2083,In_893,In_0);
nor U2084 (N_2084,In_945,In_525);
nand U2085 (N_2085,In_692,In_342);
or U2086 (N_2086,In_135,In_173);
nor U2087 (N_2087,In_748,In_695);
nand U2088 (N_2088,In_991,In_112);
and U2089 (N_2089,In_244,In_88);
nand U2090 (N_2090,In_892,In_64);
and U2091 (N_2091,In_480,In_31);
nor U2092 (N_2092,In_407,In_737);
nor U2093 (N_2093,In_418,In_930);
and U2094 (N_2094,In_980,In_564);
nand U2095 (N_2095,In_57,In_461);
nor U2096 (N_2096,In_612,In_678);
or U2097 (N_2097,In_110,In_323);
and U2098 (N_2098,In_605,In_355);
or U2099 (N_2099,In_152,In_920);
and U2100 (N_2100,In_482,In_185);
and U2101 (N_2101,In_989,In_50);
nor U2102 (N_2102,In_872,In_545);
nand U2103 (N_2103,In_763,In_628);
and U2104 (N_2104,In_92,In_547);
nor U2105 (N_2105,In_874,In_662);
nor U2106 (N_2106,In_233,In_232);
or U2107 (N_2107,In_981,In_865);
or U2108 (N_2108,In_683,In_243);
nor U2109 (N_2109,In_183,In_726);
nor U2110 (N_2110,In_583,In_971);
or U2111 (N_2111,In_16,In_982);
or U2112 (N_2112,In_984,In_820);
or U2113 (N_2113,In_897,In_496);
and U2114 (N_2114,In_775,In_917);
nand U2115 (N_2115,In_261,In_412);
and U2116 (N_2116,In_152,In_720);
nor U2117 (N_2117,In_165,In_736);
and U2118 (N_2118,In_614,In_75);
and U2119 (N_2119,In_630,In_146);
xor U2120 (N_2120,In_15,In_914);
nand U2121 (N_2121,In_499,In_602);
and U2122 (N_2122,In_101,In_394);
nor U2123 (N_2123,In_674,In_425);
nor U2124 (N_2124,In_550,In_141);
or U2125 (N_2125,In_996,In_137);
nor U2126 (N_2126,In_26,In_749);
and U2127 (N_2127,In_298,In_214);
and U2128 (N_2128,In_900,In_350);
nor U2129 (N_2129,In_388,In_165);
xor U2130 (N_2130,In_875,In_547);
and U2131 (N_2131,In_829,In_483);
or U2132 (N_2132,In_330,In_147);
nor U2133 (N_2133,In_300,In_688);
or U2134 (N_2134,In_587,In_241);
or U2135 (N_2135,In_199,In_382);
and U2136 (N_2136,In_250,In_196);
or U2137 (N_2137,In_60,In_948);
and U2138 (N_2138,In_888,In_785);
nor U2139 (N_2139,In_610,In_993);
nor U2140 (N_2140,In_639,In_931);
nand U2141 (N_2141,In_276,In_651);
or U2142 (N_2142,In_617,In_428);
and U2143 (N_2143,In_877,In_737);
or U2144 (N_2144,In_487,In_27);
nand U2145 (N_2145,In_26,In_165);
nor U2146 (N_2146,In_417,In_265);
xor U2147 (N_2147,In_872,In_969);
and U2148 (N_2148,In_687,In_84);
nor U2149 (N_2149,In_794,In_683);
nand U2150 (N_2150,In_827,In_613);
nor U2151 (N_2151,In_223,In_805);
and U2152 (N_2152,In_73,In_949);
nor U2153 (N_2153,In_982,In_987);
and U2154 (N_2154,In_377,In_314);
or U2155 (N_2155,In_544,In_947);
nor U2156 (N_2156,In_135,In_835);
nor U2157 (N_2157,In_295,In_546);
nor U2158 (N_2158,In_266,In_595);
or U2159 (N_2159,In_60,In_117);
nor U2160 (N_2160,In_813,In_622);
nand U2161 (N_2161,In_466,In_766);
nand U2162 (N_2162,In_208,In_300);
nor U2163 (N_2163,In_381,In_541);
xnor U2164 (N_2164,In_230,In_866);
or U2165 (N_2165,In_760,In_787);
or U2166 (N_2166,In_866,In_500);
or U2167 (N_2167,In_527,In_850);
and U2168 (N_2168,In_610,In_786);
and U2169 (N_2169,In_533,In_478);
nor U2170 (N_2170,In_902,In_33);
or U2171 (N_2171,In_633,In_407);
and U2172 (N_2172,In_750,In_331);
nor U2173 (N_2173,In_103,In_891);
nor U2174 (N_2174,In_606,In_384);
nor U2175 (N_2175,In_282,In_678);
and U2176 (N_2176,In_179,In_602);
and U2177 (N_2177,In_75,In_192);
nand U2178 (N_2178,In_881,In_19);
nand U2179 (N_2179,In_615,In_802);
or U2180 (N_2180,In_655,In_793);
and U2181 (N_2181,In_765,In_722);
or U2182 (N_2182,In_96,In_961);
and U2183 (N_2183,In_815,In_163);
or U2184 (N_2184,In_831,In_21);
nor U2185 (N_2185,In_148,In_6);
and U2186 (N_2186,In_467,In_14);
nor U2187 (N_2187,In_745,In_321);
and U2188 (N_2188,In_39,In_183);
or U2189 (N_2189,In_552,In_490);
xor U2190 (N_2190,In_305,In_811);
nor U2191 (N_2191,In_239,In_305);
nand U2192 (N_2192,In_757,In_489);
or U2193 (N_2193,In_178,In_403);
and U2194 (N_2194,In_91,In_779);
nand U2195 (N_2195,In_561,In_507);
nor U2196 (N_2196,In_266,In_510);
or U2197 (N_2197,In_902,In_423);
or U2198 (N_2198,In_332,In_436);
nor U2199 (N_2199,In_760,In_231);
and U2200 (N_2200,In_938,In_668);
nand U2201 (N_2201,In_396,In_802);
or U2202 (N_2202,In_647,In_668);
and U2203 (N_2203,In_876,In_361);
or U2204 (N_2204,In_466,In_96);
or U2205 (N_2205,In_61,In_27);
or U2206 (N_2206,In_833,In_386);
and U2207 (N_2207,In_751,In_228);
nand U2208 (N_2208,In_328,In_568);
and U2209 (N_2209,In_537,In_809);
nor U2210 (N_2210,In_683,In_15);
or U2211 (N_2211,In_787,In_656);
nor U2212 (N_2212,In_918,In_838);
and U2213 (N_2213,In_740,In_93);
or U2214 (N_2214,In_900,In_41);
or U2215 (N_2215,In_819,In_885);
or U2216 (N_2216,In_387,In_397);
and U2217 (N_2217,In_384,In_570);
nand U2218 (N_2218,In_697,In_638);
and U2219 (N_2219,In_61,In_826);
nand U2220 (N_2220,In_45,In_874);
or U2221 (N_2221,In_14,In_339);
nor U2222 (N_2222,In_243,In_830);
xor U2223 (N_2223,In_520,In_813);
nand U2224 (N_2224,In_936,In_569);
nor U2225 (N_2225,In_845,In_626);
nand U2226 (N_2226,In_726,In_750);
nand U2227 (N_2227,In_749,In_216);
nand U2228 (N_2228,In_979,In_256);
and U2229 (N_2229,In_73,In_739);
and U2230 (N_2230,In_476,In_282);
or U2231 (N_2231,In_173,In_4);
nor U2232 (N_2232,In_457,In_421);
nand U2233 (N_2233,In_139,In_504);
nor U2234 (N_2234,In_151,In_828);
nor U2235 (N_2235,In_104,In_918);
nand U2236 (N_2236,In_330,In_96);
or U2237 (N_2237,In_346,In_799);
and U2238 (N_2238,In_913,In_26);
nand U2239 (N_2239,In_68,In_438);
nand U2240 (N_2240,In_279,In_112);
and U2241 (N_2241,In_939,In_925);
nand U2242 (N_2242,In_274,In_675);
or U2243 (N_2243,In_402,In_489);
and U2244 (N_2244,In_9,In_898);
and U2245 (N_2245,In_684,In_134);
and U2246 (N_2246,In_181,In_138);
nand U2247 (N_2247,In_949,In_310);
nand U2248 (N_2248,In_530,In_6);
nor U2249 (N_2249,In_385,In_425);
xor U2250 (N_2250,In_164,In_583);
or U2251 (N_2251,In_798,In_217);
and U2252 (N_2252,In_485,In_572);
and U2253 (N_2253,In_364,In_579);
nand U2254 (N_2254,In_162,In_992);
or U2255 (N_2255,In_714,In_759);
or U2256 (N_2256,In_59,In_902);
or U2257 (N_2257,In_335,In_445);
nor U2258 (N_2258,In_88,In_924);
and U2259 (N_2259,In_826,In_11);
and U2260 (N_2260,In_460,In_365);
xor U2261 (N_2261,In_58,In_789);
and U2262 (N_2262,In_608,In_53);
or U2263 (N_2263,In_695,In_750);
or U2264 (N_2264,In_233,In_414);
or U2265 (N_2265,In_77,In_23);
nor U2266 (N_2266,In_667,In_947);
nor U2267 (N_2267,In_562,In_214);
or U2268 (N_2268,In_736,In_279);
nand U2269 (N_2269,In_459,In_541);
or U2270 (N_2270,In_975,In_968);
and U2271 (N_2271,In_256,In_224);
or U2272 (N_2272,In_376,In_813);
or U2273 (N_2273,In_908,In_832);
nor U2274 (N_2274,In_704,In_710);
or U2275 (N_2275,In_290,In_88);
nor U2276 (N_2276,In_644,In_250);
or U2277 (N_2277,In_256,In_954);
and U2278 (N_2278,In_626,In_766);
nor U2279 (N_2279,In_460,In_302);
nand U2280 (N_2280,In_846,In_50);
and U2281 (N_2281,In_518,In_49);
nand U2282 (N_2282,In_636,In_139);
and U2283 (N_2283,In_768,In_18);
nand U2284 (N_2284,In_515,In_255);
nand U2285 (N_2285,In_661,In_876);
nand U2286 (N_2286,In_791,In_323);
nor U2287 (N_2287,In_34,In_351);
nor U2288 (N_2288,In_339,In_643);
nand U2289 (N_2289,In_192,In_289);
nor U2290 (N_2290,In_259,In_666);
or U2291 (N_2291,In_190,In_675);
and U2292 (N_2292,In_467,In_828);
nand U2293 (N_2293,In_458,In_742);
xnor U2294 (N_2294,In_734,In_398);
and U2295 (N_2295,In_309,In_499);
nor U2296 (N_2296,In_329,In_640);
nand U2297 (N_2297,In_322,In_185);
or U2298 (N_2298,In_375,In_106);
and U2299 (N_2299,In_520,In_671);
or U2300 (N_2300,In_258,In_166);
or U2301 (N_2301,In_753,In_967);
or U2302 (N_2302,In_113,In_237);
and U2303 (N_2303,In_50,In_156);
or U2304 (N_2304,In_447,In_416);
nor U2305 (N_2305,In_978,In_243);
and U2306 (N_2306,In_88,In_309);
and U2307 (N_2307,In_999,In_690);
nor U2308 (N_2308,In_734,In_971);
and U2309 (N_2309,In_806,In_451);
nor U2310 (N_2310,In_431,In_798);
nor U2311 (N_2311,In_729,In_149);
nor U2312 (N_2312,In_130,In_845);
and U2313 (N_2313,In_347,In_144);
or U2314 (N_2314,In_886,In_571);
nor U2315 (N_2315,In_539,In_951);
nor U2316 (N_2316,In_905,In_271);
and U2317 (N_2317,In_316,In_342);
or U2318 (N_2318,In_321,In_722);
and U2319 (N_2319,In_970,In_20);
nor U2320 (N_2320,In_555,In_879);
or U2321 (N_2321,In_485,In_359);
and U2322 (N_2322,In_592,In_260);
nand U2323 (N_2323,In_238,In_274);
or U2324 (N_2324,In_980,In_307);
or U2325 (N_2325,In_451,In_208);
nand U2326 (N_2326,In_490,In_350);
nor U2327 (N_2327,In_139,In_499);
and U2328 (N_2328,In_450,In_797);
or U2329 (N_2329,In_562,In_579);
nand U2330 (N_2330,In_944,In_485);
nand U2331 (N_2331,In_519,In_913);
xnor U2332 (N_2332,In_829,In_670);
nor U2333 (N_2333,In_689,In_810);
nand U2334 (N_2334,In_226,In_350);
nor U2335 (N_2335,In_499,In_583);
and U2336 (N_2336,In_241,In_475);
nor U2337 (N_2337,In_947,In_586);
nand U2338 (N_2338,In_608,In_607);
and U2339 (N_2339,In_747,In_960);
or U2340 (N_2340,In_892,In_902);
or U2341 (N_2341,In_191,In_328);
nand U2342 (N_2342,In_35,In_106);
nor U2343 (N_2343,In_825,In_620);
nand U2344 (N_2344,In_448,In_632);
or U2345 (N_2345,In_205,In_522);
or U2346 (N_2346,In_148,In_780);
or U2347 (N_2347,In_435,In_320);
nor U2348 (N_2348,In_154,In_814);
and U2349 (N_2349,In_607,In_171);
xor U2350 (N_2350,In_34,In_559);
or U2351 (N_2351,In_837,In_397);
or U2352 (N_2352,In_429,In_7);
nor U2353 (N_2353,In_32,In_36);
and U2354 (N_2354,In_595,In_748);
or U2355 (N_2355,In_929,In_838);
and U2356 (N_2356,In_351,In_717);
nand U2357 (N_2357,In_410,In_762);
or U2358 (N_2358,In_503,In_590);
nand U2359 (N_2359,In_206,In_980);
nand U2360 (N_2360,In_820,In_711);
nand U2361 (N_2361,In_51,In_224);
nor U2362 (N_2362,In_60,In_47);
nand U2363 (N_2363,In_211,In_682);
nand U2364 (N_2364,In_85,In_219);
nand U2365 (N_2365,In_563,In_214);
nand U2366 (N_2366,In_194,In_640);
nand U2367 (N_2367,In_24,In_899);
and U2368 (N_2368,In_793,In_842);
nand U2369 (N_2369,In_973,In_645);
and U2370 (N_2370,In_795,In_634);
nand U2371 (N_2371,In_905,In_288);
or U2372 (N_2372,In_952,In_326);
xor U2373 (N_2373,In_317,In_236);
or U2374 (N_2374,In_150,In_175);
xnor U2375 (N_2375,In_195,In_387);
xnor U2376 (N_2376,In_792,In_430);
nor U2377 (N_2377,In_747,In_685);
or U2378 (N_2378,In_353,In_620);
nand U2379 (N_2379,In_716,In_926);
or U2380 (N_2380,In_131,In_864);
nor U2381 (N_2381,In_498,In_709);
nor U2382 (N_2382,In_598,In_925);
or U2383 (N_2383,In_537,In_166);
nor U2384 (N_2384,In_612,In_996);
nand U2385 (N_2385,In_310,In_678);
nor U2386 (N_2386,In_469,In_486);
or U2387 (N_2387,In_693,In_798);
and U2388 (N_2388,In_266,In_130);
nor U2389 (N_2389,In_986,In_773);
nand U2390 (N_2390,In_834,In_370);
and U2391 (N_2391,In_733,In_191);
or U2392 (N_2392,In_50,In_155);
nand U2393 (N_2393,In_41,In_850);
nand U2394 (N_2394,In_324,In_799);
nand U2395 (N_2395,In_657,In_807);
nand U2396 (N_2396,In_683,In_193);
or U2397 (N_2397,In_564,In_880);
nand U2398 (N_2398,In_765,In_603);
and U2399 (N_2399,In_230,In_564);
nand U2400 (N_2400,In_964,In_424);
nand U2401 (N_2401,In_649,In_0);
or U2402 (N_2402,In_185,In_922);
nand U2403 (N_2403,In_807,In_586);
nand U2404 (N_2404,In_456,In_568);
nor U2405 (N_2405,In_31,In_811);
or U2406 (N_2406,In_188,In_943);
or U2407 (N_2407,In_114,In_47);
and U2408 (N_2408,In_175,In_21);
nand U2409 (N_2409,In_754,In_645);
xor U2410 (N_2410,In_401,In_844);
and U2411 (N_2411,In_910,In_600);
nor U2412 (N_2412,In_235,In_743);
or U2413 (N_2413,In_815,In_252);
nor U2414 (N_2414,In_768,In_444);
nand U2415 (N_2415,In_752,In_728);
or U2416 (N_2416,In_509,In_617);
nor U2417 (N_2417,In_114,In_400);
nand U2418 (N_2418,In_804,In_986);
or U2419 (N_2419,In_690,In_463);
nor U2420 (N_2420,In_484,In_470);
or U2421 (N_2421,In_696,In_228);
nor U2422 (N_2422,In_278,In_900);
nor U2423 (N_2423,In_685,In_334);
nor U2424 (N_2424,In_375,In_925);
and U2425 (N_2425,In_685,In_815);
nand U2426 (N_2426,In_582,In_538);
nor U2427 (N_2427,In_480,In_467);
nand U2428 (N_2428,In_42,In_199);
or U2429 (N_2429,In_244,In_945);
or U2430 (N_2430,In_153,In_522);
xor U2431 (N_2431,In_166,In_752);
or U2432 (N_2432,In_361,In_478);
and U2433 (N_2433,In_61,In_167);
or U2434 (N_2434,In_439,In_691);
and U2435 (N_2435,In_29,In_5);
nand U2436 (N_2436,In_372,In_633);
nor U2437 (N_2437,In_102,In_19);
nand U2438 (N_2438,In_775,In_757);
or U2439 (N_2439,In_584,In_925);
nand U2440 (N_2440,In_292,In_116);
or U2441 (N_2441,In_372,In_213);
or U2442 (N_2442,In_232,In_126);
or U2443 (N_2443,In_1,In_346);
nor U2444 (N_2444,In_226,In_313);
nand U2445 (N_2445,In_897,In_886);
nand U2446 (N_2446,In_850,In_167);
nand U2447 (N_2447,In_124,In_150);
and U2448 (N_2448,In_342,In_969);
xor U2449 (N_2449,In_135,In_501);
or U2450 (N_2450,In_56,In_674);
or U2451 (N_2451,In_808,In_199);
nor U2452 (N_2452,In_99,In_456);
nand U2453 (N_2453,In_853,In_222);
nand U2454 (N_2454,In_782,In_689);
or U2455 (N_2455,In_345,In_560);
nor U2456 (N_2456,In_196,In_602);
and U2457 (N_2457,In_573,In_153);
nor U2458 (N_2458,In_672,In_470);
nand U2459 (N_2459,In_369,In_47);
and U2460 (N_2460,In_4,In_736);
nor U2461 (N_2461,In_249,In_33);
nor U2462 (N_2462,In_184,In_239);
or U2463 (N_2463,In_313,In_339);
and U2464 (N_2464,In_96,In_836);
and U2465 (N_2465,In_354,In_448);
or U2466 (N_2466,In_749,In_830);
and U2467 (N_2467,In_230,In_629);
and U2468 (N_2468,In_808,In_501);
nand U2469 (N_2469,In_670,In_895);
nand U2470 (N_2470,In_440,In_944);
nor U2471 (N_2471,In_518,In_792);
nor U2472 (N_2472,In_569,In_637);
or U2473 (N_2473,In_959,In_54);
nand U2474 (N_2474,In_280,In_464);
nor U2475 (N_2475,In_890,In_158);
nand U2476 (N_2476,In_503,In_280);
nor U2477 (N_2477,In_371,In_761);
or U2478 (N_2478,In_975,In_32);
and U2479 (N_2479,In_285,In_999);
or U2480 (N_2480,In_986,In_728);
nand U2481 (N_2481,In_327,In_556);
and U2482 (N_2482,In_788,In_120);
or U2483 (N_2483,In_363,In_26);
nand U2484 (N_2484,In_246,In_744);
or U2485 (N_2485,In_323,In_373);
nor U2486 (N_2486,In_787,In_918);
nand U2487 (N_2487,In_773,In_818);
nand U2488 (N_2488,In_168,In_93);
and U2489 (N_2489,In_957,In_43);
nand U2490 (N_2490,In_425,In_677);
nand U2491 (N_2491,In_948,In_121);
nand U2492 (N_2492,In_67,In_189);
and U2493 (N_2493,In_493,In_5);
nor U2494 (N_2494,In_367,In_967);
and U2495 (N_2495,In_592,In_764);
nand U2496 (N_2496,In_508,In_232);
nor U2497 (N_2497,In_379,In_580);
nand U2498 (N_2498,In_275,In_216);
nand U2499 (N_2499,In_531,In_943);
and U2500 (N_2500,In_260,In_163);
nor U2501 (N_2501,In_794,In_77);
xnor U2502 (N_2502,In_589,In_556);
and U2503 (N_2503,In_822,In_278);
or U2504 (N_2504,In_33,In_238);
nand U2505 (N_2505,In_470,In_560);
nor U2506 (N_2506,In_817,In_691);
or U2507 (N_2507,In_60,In_910);
or U2508 (N_2508,In_447,In_169);
or U2509 (N_2509,In_842,In_575);
and U2510 (N_2510,In_973,In_9);
nand U2511 (N_2511,In_278,In_292);
nand U2512 (N_2512,In_176,In_353);
or U2513 (N_2513,In_558,In_592);
and U2514 (N_2514,In_948,In_711);
nor U2515 (N_2515,In_298,In_595);
nor U2516 (N_2516,In_265,In_535);
nor U2517 (N_2517,In_555,In_299);
or U2518 (N_2518,In_330,In_954);
nor U2519 (N_2519,In_38,In_460);
nand U2520 (N_2520,In_698,In_254);
nor U2521 (N_2521,In_76,In_69);
or U2522 (N_2522,In_879,In_72);
nand U2523 (N_2523,In_549,In_640);
and U2524 (N_2524,In_600,In_342);
or U2525 (N_2525,In_604,In_988);
or U2526 (N_2526,In_590,In_620);
nor U2527 (N_2527,In_388,In_572);
or U2528 (N_2528,In_342,In_232);
nand U2529 (N_2529,In_384,In_426);
xnor U2530 (N_2530,In_741,In_457);
nand U2531 (N_2531,In_946,In_48);
or U2532 (N_2532,In_669,In_289);
or U2533 (N_2533,In_356,In_26);
and U2534 (N_2534,In_191,In_561);
or U2535 (N_2535,In_864,In_64);
and U2536 (N_2536,In_389,In_265);
or U2537 (N_2537,In_70,In_763);
and U2538 (N_2538,In_97,In_585);
and U2539 (N_2539,In_427,In_919);
nor U2540 (N_2540,In_498,In_219);
or U2541 (N_2541,In_562,In_584);
nand U2542 (N_2542,In_379,In_66);
nand U2543 (N_2543,In_554,In_700);
or U2544 (N_2544,In_94,In_590);
or U2545 (N_2545,In_328,In_913);
nand U2546 (N_2546,In_361,In_597);
nor U2547 (N_2547,In_956,In_400);
and U2548 (N_2548,In_306,In_680);
or U2549 (N_2549,In_148,In_185);
and U2550 (N_2550,In_128,In_784);
nor U2551 (N_2551,In_862,In_248);
or U2552 (N_2552,In_987,In_885);
nor U2553 (N_2553,In_531,In_279);
and U2554 (N_2554,In_925,In_529);
xor U2555 (N_2555,In_669,In_833);
nand U2556 (N_2556,In_366,In_228);
nand U2557 (N_2557,In_716,In_278);
or U2558 (N_2558,In_367,In_795);
or U2559 (N_2559,In_59,In_448);
and U2560 (N_2560,In_199,In_541);
nand U2561 (N_2561,In_16,In_591);
nand U2562 (N_2562,In_104,In_303);
nand U2563 (N_2563,In_771,In_479);
nand U2564 (N_2564,In_265,In_195);
nor U2565 (N_2565,In_195,In_936);
or U2566 (N_2566,In_268,In_678);
nor U2567 (N_2567,In_457,In_455);
or U2568 (N_2568,In_977,In_249);
and U2569 (N_2569,In_654,In_432);
or U2570 (N_2570,In_101,In_696);
or U2571 (N_2571,In_530,In_532);
nand U2572 (N_2572,In_829,In_798);
nand U2573 (N_2573,In_513,In_332);
nor U2574 (N_2574,In_458,In_542);
nor U2575 (N_2575,In_611,In_951);
nor U2576 (N_2576,In_510,In_806);
nand U2577 (N_2577,In_816,In_636);
or U2578 (N_2578,In_939,In_208);
xor U2579 (N_2579,In_322,In_244);
and U2580 (N_2580,In_638,In_388);
nor U2581 (N_2581,In_25,In_290);
nor U2582 (N_2582,In_355,In_422);
nor U2583 (N_2583,In_656,In_927);
nand U2584 (N_2584,In_614,In_917);
nor U2585 (N_2585,In_807,In_902);
and U2586 (N_2586,In_291,In_443);
nand U2587 (N_2587,In_557,In_409);
nand U2588 (N_2588,In_851,In_498);
and U2589 (N_2589,In_651,In_222);
and U2590 (N_2590,In_999,In_220);
or U2591 (N_2591,In_482,In_935);
nand U2592 (N_2592,In_539,In_869);
nand U2593 (N_2593,In_686,In_298);
and U2594 (N_2594,In_731,In_278);
or U2595 (N_2595,In_121,In_211);
nor U2596 (N_2596,In_767,In_839);
or U2597 (N_2597,In_217,In_490);
nor U2598 (N_2598,In_539,In_161);
nor U2599 (N_2599,In_879,In_968);
and U2600 (N_2600,In_622,In_182);
and U2601 (N_2601,In_458,In_864);
nor U2602 (N_2602,In_97,In_532);
nand U2603 (N_2603,In_930,In_86);
nor U2604 (N_2604,In_163,In_130);
or U2605 (N_2605,In_900,In_973);
or U2606 (N_2606,In_98,In_298);
or U2607 (N_2607,In_993,In_812);
and U2608 (N_2608,In_497,In_511);
nand U2609 (N_2609,In_255,In_803);
and U2610 (N_2610,In_252,In_45);
nor U2611 (N_2611,In_345,In_617);
nand U2612 (N_2612,In_351,In_836);
and U2613 (N_2613,In_2,In_740);
or U2614 (N_2614,In_461,In_577);
or U2615 (N_2615,In_97,In_487);
and U2616 (N_2616,In_525,In_683);
nor U2617 (N_2617,In_806,In_393);
nor U2618 (N_2618,In_314,In_379);
nor U2619 (N_2619,In_272,In_962);
or U2620 (N_2620,In_279,In_413);
or U2621 (N_2621,In_597,In_302);
or U2622 (N_2622,In_563,In_184);
or U2623 (N_2623,In_155,In_219);
and U2624 (N_2624,In_298,In_250);
nor U2625 (N_2625,In_287,In_151);
nand U2626 (N_2626,In_443,In_28);
nand U2627 (N_2627,In_598,In_281);
and U2628 (N_2628,In_850,In_332);
or U2629 (N_2629,In_162,In_205);
nor U2630 (N_2630,In_42,In_229);
xor U2631 (N_2631,In_846,In_404);
and U2632 (N_2632,In_988,In_424);
nand U2633 (N_2633,In_674,In_263);
nor U2634 (N_2634,In_783,In_908);
and U2635 (N_2635,In_736,In_725);
or U2636 (N_2636,In_921,In_172);
and U2637 (N_2637,In_303,In_200);
nor U2638 (N_2638,In_84,In_74);
and U2639 (N_2639,In_872,In_192);
nor U2640 (N_2640,In_956,In_492);
and U2641 (N_2641,In_861,In_475);
nor U2642 (N_2642,In_597,In_385);
nand U2643 (N_2643,In_319,In_732);
and U2644 (N_2644,In_70,In_768);
or U2645 (N_2645,In_615,In_665);
xnor U2646 (N_2646,In_421,In_665);
and U2647 (N_2647,In_775,In_354);
or U2648 (N_2648,In_825,In_15);
or U2649 (N_2649,In_813,In_888);
or U2650 (N_2650,In_722,In_958);
nand U2651 (N_2651,In_93,In_631);
nand U2652 (N_2652,In_697,In_642);
and U2653 (N_2653,In_739,In_754);
and U2654 (N_2654,In_165,In_418);
and U2655 (N_2655,In_980,In_655);
or U2656 (N_2656,In_445,In_760);
nand U2657 (N_2657,In_775,In_344);
nor U2658 (N_2658,In_439,In_353);
and U2659 (N_2659,In_456,In_862);
or U2660 (N_2660,In_494,In_455);
and U2661 (N_2661,In_944,In_11);
and U2662 (N_2662,In_912,In_502);
nor U2663 (N_2663,In_501,In_623);
nor U2664 (N_2664,In_370,In_407);
nor U2665 (N_2665,In_985,In_521);
nor U2666 (N_2666,In_358,In_416);
or U2667 (N_2667,In_232,In_890);
and U2668 (N_2668,In_985,In_509);
nand U2669 (N_2669,In_433,In_607);
and U2670 (N_2670,In_1,In_981);
nor U2671 (N_2671,In_597,In_645);
nand U2672 (N_2672,In_944,In_582);
or U2673 (N_2673,In_23,In_218);
nand U2674 (N_2674,In_948,In_881);
or U2675 (N_2675,In_604,In_867);
nand U2676 (N_2676,In_39,In_526);
and U2677 (N_2677,In_55,In_700);
nand U2678 (N_2678,In_530,In_11);
nor U2679 (N_2679,In_17,In_700);
and U2680 (N_2680,In_358,In_966);
nand U2681 (N_2681,In_890,In_548);
and U2682 (N_2682,In_809,In_16);
and U2683 (N_2683,In_505,In_606);
nor U2684 (N_2684,In_864,In_835);
nand U2685 (N_2685,In_150,In_774);
or U2686 (N_2686,In_785,In_99);
and U2687 (N_2687,In_916,In_486);
and U2688 (N_2688,In_501,In_969);
nor U2689 (N_2689,In_164,In_661);
nand U2690 (N_2690,In_869,In_538);
and U2691 (N_2691,In_573,In_47);
nand U2692 (N_2692,In_339,In_144);
or U2693 (N_2693,In_203,In_344);
or U2694 (N_2694,In_179,In_290);
nor U2695 (N_2695,In_802,In_246);
or U2696 (N_2696,In_446,In_372);
nor U2697 (N_2697,In_721,In_486);
nand U2698 (N_2698,In_701,In_649);
nand U2699 (N_2699,In_843,In_419);
or U2700 (N_2700,In_877,In_410);
and U2701 (N_2701,In_660,In_393);
or U2702 (N_2702,In_834,In_903);
nor U2703 (N_2703,In_810,In_701);
or U2704 (N_2704,In_618,In_402);
nor U2705 (N_2705,In_131,In_486);
or U2706 (N_2706,In_816,In_743);
or U2707 (N_2707,In_440,In_244);
nand U2708 (N_2708,In_242,In_116);
xnor U2709 (N_2709,In_350,In_725);
and U2710 (N_2710,In_598,In_479);
and U2711 (N_2711,In_477,In_6);
nor U2712 (N_2712,In_344,In_457);
nor U2713 (N_2713,In_763,In_389);
xor U2714 (N_2714,In_892,In_651);
nor U2715 (N_2715,In_488,In_707);
nand U2716 (N_2716,In_744,In_191);
nor U2717 (N_2717,In_249,In_96);
xor U2718 (N_2718,In_313,In_898);
or U2719 (N_2719,In_79,In_647);
nor U2720 (N_2720,In_832,In_220);
nand U2721 (N_2721,In_68,In_616);
nand U2722 (N_2722,In_957,In_286);
nand U2723 (N_2723,In_802,In_708);
or U2724 (N_2724,In_712,In_274);
or U2725 (N_2725,In_765,In_64);
nand U2726 (N_2726,In_101,In_287);
nand U2727 (N_2727,In_998,In_335);
nand U2728 (N_2728,In_422,In_589);
nand U2729 (N_2729,In_438,In_697);
and U2730 (N_2730,In_439,In_614);
and U2731 (N_2731,In_784,In_386);
or U2732 (N_2732,In_432,In_429);
nand U2733 (N_2733,In_426,In_121);
or U2734 (N_2734,In_151,In_470);
and U2735 (N_2735,In_840,In_938);
or U2736 (N_2736,In_757,In_350);
and U2737 (N_2737,In_451,In_824);
or U2738 (N_2738,In_574,In_457);
or U2739 (N_2739,In_125,In_60);
or U2740 (N_2740,In_157,In_247);
nand U2741 (N_2741,In_454,In_472);
and U2742 (N_2742,In_548,In_124);
or U2743 (N_2743,In_770,In_999);
nor U2744 (N_2744,In_238,In_13);
nand U2745 (N_2745,In_223,In_775);
nor U2746 (N_2746,In_983,In_845);
and U2747 (N_2747,In_27,In_534);
and U2748 (N_2748,In_438,In_137);
nor U2749 (N_2749,In_260,In_165);
nand U2750 (N_2750,In_366,In_31);
nand U2751 (N_2751,In_777,In_101);
or U2752 (N_2752,In_245,In_395);
nand U2753 (N_2753,In_476,In_575);
nand U2754 (N_2754,In_896,In_487);
nand U2755 (N_2755,In_869,In_567);
nor U2756 (N_2756,In_757,In_353);
or U2757 (N_2757,In_406,In_166);
and U2758 (N_2758,In_941,In_678);
or U2759 (N_2759,In_94,In_854);
and U2760 (N_2760,In_877,In_246);
nand U2761 (N_2761,In_319,In_267);
nand U2762 (N_2762,In_199,In_588);
or U2763 (N_2763,In_332,In_140);
nand U2764 (N_2764,In_156,In_346);
nor U2765 (N_2765,In_476,In_355);
and U2766 (N_2766,In_68,In_109);
and U2767 (N_2767,In_280,In_560);
and U2768 (N_2768,In_71,In_230);
nand U2769 (N_2769,In_704,In_205);
nor U2770 (N_2770,In_75,In_471);
and U2771 (N_2771,In_145,In_674);
nand U2772 (N_2772,In_648,In_804);
and U2773 (N_2773,In_543,In_168);
nand U2774 (N_2774,In_371,In_488);
or U2775 (N_2775,In_965,In_261);
or U2776 (N_2776,In_905,In_794);
and U2777 (N_2777,In_317,In_602);
and U2778 (N_2778,In_931,In_366);
or U2779 (N_2779,In_240,In_78);
nor U2780 (N_2780,In_283,In_474);
and U2781 (N_2781,In_521,In_71);
and U2782 (N_2782,In_441,In_235);
xnor U2783 (N_2783,In_501,In_862);
nand U2784 (N_2784,In_621,In_537);
or U2785 (N_2785,In_760,In_685);
and U2786 (N_2786,In_372,In_968);
and U2787 (N_2787,In_644,In_450);
nand U2788 (N_2788,In_142,In_832);
nor U2789 (N_2789,In_922,In_984);
nor U2790 (N_2790,In_39,In_576);
nor U2791 (N_2791,In_335,In_999);
or U2792 (N_2792,In_940,In_452);
nor U2793 (N_2793,In_754,In_347);
or U2794 (N_2794,In_648,In_470);
nand U2795 (N_2795,In_798,In_499);
nor U2796 (N_2796,In_947,In_693);
and U2797 (N_2797,In_635,In_39);
or U2798 (N_2798,In_357,In_375);
or U2799 (N_2799,In_184,In_875);
nand U2800 (N_2800,In_386,In_922);
and U2801 (N_2801,In_31,In_825);
or U2802 (N_2802,In_719,In_948);
nand U2803 (N_2803,In_534,In_490);
nand U2804 (N_2804,In_662,In_884);
and U2805 (N_2805,In_634,In_36);
nand U2806 (N_2806,In_61,In_854);
and U2807 (N_2807,In_649,In_955);
and U2808 (N_2808,In_126,In_697);
nor U2809 (N_2809,In_387,In_438);
and U2810 (N_2810,In_319,In_152);
nor U2811 (N_2811,In_358,In_664);
nor U2812 (N_2812,In_89,In_349);
nor U2813 (N_2813,In_907,In_215);
xor U2814 (N_2814,In_233,In_874);
nand U2815 (N_2815,In_305,In_95);
or U2816 (N_2816,In_541,In_385);
xor U2817 (N_2817,In_373,In_274);
nor U2818 (N_2818,In_797,In_743);
and U2819 (N_2819,In_591,In_620);
or U2820 (N_2820,In_86,In_543);
and U2821 (N_2821,In_105,In_19);
or U2822 (N_2822,In_865,In_279);
and U2823 (N_2823,In_857,In_826);
nor U2824 (N_2824,In_372,In_824);
nand U2825 (N_2825,In_93,In_795);
nor U2826 (N_2826,In_499,In_993);
nand U2827 (N_2827,In_587,In_836);
nor U2828 (N_2828,In_932,In_55);
or U2829 (N_2829,In_525,In_160);
or U2830 (N_2830,In_867,In_7);
nor U2831 (N_2831,In_819,In_232);
or U2832 (N_2832,In_472,In_398);
and U2833 (N_2833,In_991,In_705);
nand U2834 (N_2834,In_36,In_363);
nor U2835 (N_2835,In_431,In_336);
nand U2836 (N_2836,In_235,In_741);
nor U2837 (N_2837,In_325,In_712);
or U2838 (N_2838,In_792,In_380);
nand U2839 (N_2839,In_940,In_148);
and U2840 (N_2840,In_407,In_935);
nand U2841 (N_2841,In_472,In_776);
nor U2842 (N_2842,In_548,In_938);
nand U2843 (N_2843,In_988,In_43);
or U2844 (N_2844,In_589,In_82);
nor U2845 (N_2845,In_581,In_765);
nor U2846 (N_2846,In_112,In_832);
nor U2847 (N_2847,In_881,In_674);
or U2848 (N_2848,In_371,In_534);
or U2849 (N_2849,In_511,In_866);
nor U2850 (N_2850,In_831,In_309);
and U2851 (N_2851,In_5,In_791);
nand U2852 (N_2852,In_278,In_509);
nor U2853 (N_2853,In_602,In_457);
or U2854 (N_2854,In_222,In_899);
nor U2855 (N_2855,In_429,In_131);
nor U2856 (N_2856,In_232,In_409);
nand U2857 (N_2857,In_879,In_616);
or U2858 (N_2858,In_497,In_284);
nor U2859 (N_2859,In_324,In_777);
nand U2860 (N_2860,In_425,In_734);
or U2861 (N_2861,In_210,In_612);
nand U2862 (N_2862,In_296,In_159);
nor U2863 (N_2863,In_451,In_768);
or U2864 (N_2864,In_25,In_102);
or U2865 (N_2865,In_296,In_431);
or U2866 (N_2866,In_698,In_290);
and U2867 (N_2867,In_733,In_29);
nand U2868 (N_2868,In_668,In_105);
and U2869 (N_2869,In_62,In_728);
or U2870 (N_2870,In_171,In_453);
or U2871 (N_2871,In_48,In_291);
or U2872 (N_2872,In_423,In_756);
nor U2873 (N_2873,In_668,In_628);
nand U2874 (N_2874,In_216,In_18);
nor U2875 (N_2875,In_564,In_231);
nor U2876 (N_2876,In_64,In_745);
nor U2877 (N_2877,In_285,In_268);
nand U2878 (N_2878,In_176,In_238);
and U2879 (N_2879,In_928,In_390);
nor U2880 (N_2880,In_814,In_782);
or U2881 (N_2881,In_522,In_179);
nand U2882 (N_2882,In_229,In_707);
nor U2883 (N_2883,In_354,In_398);
nor U2884 (N_2884,In_966,In_12);
and U2885 (N_2885,In_452,In_919);
and U2886 (N_2886,In_191,In_811);
or U2887 (N_2887,In_415,In_425);
or U2888 (N_2888,In_553,In_530);
nand U2889 (N_2889,In_426,In_268);
or U2890 (N_2890,In_903,In_189);
nand U2891 (N_2891,In_301,In_226);
and U2892 (N_2892,In_414,In_756);
and U2893 (N_2893,In_769,In_650);
and U2894 (N_2894,In_502,In_689);
nor U2895 (N_2895,In_505,In_126);
nor U2896 (N_2896,In_163,In_308);
nor U2897 (N_2897,In_420,In_476);
nor U2898 (N_2898,In_232,In_548);
nor U2899 (N_2899,In_93,In_562);
or U2900 (N_2900,In_651,In_196);
nor U2901 (N_2901,In_800,In_361);
nand U2902 (N_2902,In_293,In_798);
or U2903 (N_2903,In_881,In_324);
nor U2904 (N_2904,In_108,In_652);
nor U2905 (N_2905,In_98,In_64);
nand U2906 (N_2906,In_108,In_616);
and U2907 (N_2907,In_607,In_831);
or U2908 (N_2908,In_946,In_376);
nor U2909 (N_2909,In_51,In_184);
and U2910 (N_2910,In_881,In_666);
or U2911 (N_2911,In_641,In_336);
or U2912 (N_2912,In_545,In_397);
nor U2913 (N_2913,In_240,In_213);
nand U2914 (N_2914,In_827,In_987);
nand U2915 (N_2915,In_588,In_148);
or U2916 (N_2916,In_977,In_953);
nor U2917 (N_2917,In_429,In_454);
or U2918 (N_2918,In_209,In_333);
and U2919 (N_2919,In_923,In_734);
nor U2920 (N_2920,In_535,In_401);
nand U2921 (N_2921,In_348,In_292);
nor U2922 (N_2922,In_345,In_244);
and U2923 (N_2923,In_303,In_772);
and U2924 (N_2924,In_148,In_489);
or U2925 (N_2925,In_780,In_509);
and U2926 (N_2926,In_189,In_647);
nand U2927 (N_2927,In_806,In_726);
and U2928 (N_2928,In_527,In_594);
and U2929 (N_2929,In_772,In_739);
or U2930 (N_2930,In_397,In_48);
and U2931 (N_2931,In_884,In_237);
nor U2932 (N_2932,In_80,In_894);
or U2933 (N_2933,In_55,In_376);
or U2934 (N_2934,In_754,In_591);
nand U2935 (N_2935,In_811,In_202);
nor U2936 (N_2936,In_847,In_855);
nand U2937 (N_2937,In_573,In_688);
or U2938 (N_2938,In_719,In_106);
and U2939 (N_2939,In_205,In_558);
and U2940 (N_2940,In_456,In_477);
nor U2941 (N_2941,In_492,In_783);
and U2942 (N_2942,In_824,In_928);
and U2943 (N_2943,In_399,In_159);
and U2944 (N_2944,In_901,In_812);
and U2945 (N_2945,In_0,In_297);
or U2946 (N_2946,In_352,In_911);
nor U2947 (N_2947,In_371,In_445);
nor U2948 (N_2948,In_14,In_521);
nand U2949 (N_2949,In_906,In_994);
nor U2950 (N_2950,In_860,In_702);
and U2951 (N_2951,In_262,In_632);
and U2952 (N_2952,In_198,In_69);
nand U2953 (N_2953,In_431,In_513);
or U2954 (N_2954,In_576,In_149);
or U2955 (N_2955,In_426,In_798);
and U2956 (N_2956,In_336,In_856);
or U2957 (N_2957,In_126,In_389);
nand U2958 (N_2958,In_589,In_80);
nor U2959 (N_2959,In_115,In_22);
nand U2960 (N_2960,In_383,In_872);
nor U2961 (N_2961,In_585,In_785);
and U2962 (N_2962,In_162,In_133);
or U2963 (N_2963,In_482,In_238);
and U2964 (N_2964,In_623,In_694);
and U2965 (N_2965,In_868,In_377);
nand U2966 (N_2966,In_164,In_394);
nor U2967 (N_2967,In_917,In_747);
and U2968 (N_2968,In_756,In_507);
and U2969 (N_2969,In_174,In_328);
or U2970 (N_2970,In_66,In_595);
and U2971 (N_2971,In_771,In_493);
nand U2972 (N_2972,In_907,In_386);
and U2973 (N_2973,In_418,In_147);
and U2974 (N_2974,In_0,In_908);
nand U2975 (N_2975,In_405,In_968);
nand U2976 (N_2976,In_746,In_587);
nor U2977 (N_2977,In_315,In_710);
nand U2978 (N_2978,In_486,In_161);
or U2979 (N_2979,In_554,In_654);
and U2980 (N_2980,In_417,In_106);
nor U2981 (N_2981,In_710,In_129);
nand U2982 (N_2982,In_147,In_482);
or U2983 (N_2983,In_727,In_655);
xor U2984 (N_2984,In_423,In_427);
and U2985 (N_2985,In_235,In_724);
or U2986 (N_2986,In_637,In_963);
or U2987 (N_2987,In_427,In_430);
and U2988 (N_2988,In_258,In_605);
nor U2989 (N_2989,In_554,In_236);
and U2990 (N_2990,In_633,In_485);
nor U2991 (N_2991,In_425,In_839);
nand U2992 (N_2992,In_438,In_781);
nor U2993 (N_2993,In_684,In_137);
nor U2994 (N_2994,In_680,In_975);
nor U2995 (N_2995,In_409,In_684);
and U2996 (N_2996,In_355,In_768);
and U2997 (N_2997,In_89,In_857);
nor U2998 (N_2998,In_345,In_47);
and U2999 (N_2999,In_134,In_12);
or U3000 (N_3000,In_565,In_673);
nor U3001 (N_3001,In_435,In_591);
nor U3002 (N_3002,In_233,In_117);
and U3003 (N_3003,In_174,In_697);
nor U3004 (N_3004,In_743,In_659);
nor U3005 (N_3005,In_361,In_914);
xor U3006 (N_3006,In_800,In_713);
nor U3007 (N_3007,In_425,In_291);
nor U3008 (N_3008,In_405,In_59);
nand U3009 (N_3009,In_335,In_110);
and U3010 (N_3010,In_625,In_335);
nand U3011 (N_3011,In_528,In_870);
or U3012 (N_3012,In_643,In_505);
or U3013 (N_3013,In_186,In_111);
and U3014 (N_3014,In_836,In_486);
nor U3015 (N_3015,In_855,In_882);
or U3016 (N_3016,In_863,In_963);
nand U3017 (N_3017,In_647,In_567);
nor U3018 (N_3018,In_99,In_317);
and U3019 (N_3019,In_996,In_584);
and U3020 (N_3020,In_721,In_391);
nand U3021 (N_3021,In_910,In_416);
or U3022 (N_3022,In_55,In_878);
or U3023 (N_3023,In_166,In_662);
nor U3024 (N_3024,In_476,In_357);
and U3025 (N_3025,In_407,In_430);
nand U3026 (N_3026,In_719,In_627);
or U3027 (N_3027,In_614,In_97);
nor U3028 (N_3028,In_374,In_468);
nor U3029 (N_3029,In_936,In_849);
nand U3030 (N_3030,In_963,In_217);
and U3031 (N_3031,In_136,In_871);
and U3032 (N_3032,In_567,In_477);
or U3033 (N_3033,In_536,In_274);
and U3034 (N_3034,In_635,In_826);
and U3035 (N_3035,In_429,In_1);
and U3036 (N_3036,In_883,In_113);
and U3037 (N_3037,In_229,In_454);
or U3038 (N_3038,In_822,In_452);
or U3039 (N_3039,In_215,In_829);
nand U3040 (N_3040,In_922,In_860);
nand U3041 (N_3041,In_586,In_467);
and U3042 (N_3042,In_332,In_8);
nand U3043 (N_3043,In_819,In_273);
nand U3044 (N_3044,In_294,In_892);
and U3045 (N_3045,In_213,In_936);
nor U3046 (N_3046,In_499,In_559);
nand U3047 (N_3047,In_924,In_763);
nand U3048 (N_3048,In_506,In_30);
and U3049 (N_3049,In_474,In_845);
or U3050 (N_3050,In_745,In_565);
nand U3051 (N_3051,In_139,In_909);
or U3052 (N_3052,In_385,In_769);
or U3053 (N_3053,In_384,In_497);
and U3054 (N_3054,In_141,In_38);
nor U3055 (N_3055,In_187,In_407);
and U3056 (N_3056,In_314,In_893);
nor U3057 (N_3057,In_877,In_836);
nor U3058 (N_3058,In_588,In_556);
nand U3059 (N_3059,In_608,In_736);
nor U3060 (N_3060,In_429,In_810);
and U3061 (N_3061,In_591,In_327);
or U3062 (N_3062,In_899,In_209);
and U3063 (N_3063,In_393,In_900);
or U3064 (N_3064,In_369,In_805);
nor U3065 (N_3065,In_881,In_986);
nor U3066 (N_3066,In_702,In_852);
or U3067 (N_3067,In_830,In_155);
nor U3068 (N_3068,In_148,In_591);
nand U3069 (N_3069,In_423,In_895);
nor U3070 (N_3070,In_865,In_79);
nor U3071 (N_3071,In_338,In_297);
or U3072 (N_3072,In_839,In_192);
and U3073 (N_3073,In_374,In_649);
nand U3074 (N_3074,In_843,In_909);
nor U3075 (N_3075,In_792,In_338);
nor U3076 (N_3076,In_84,In_608);
nor U3077 (N_3077,In_214,In_255);
nand U3078 (N_3078,In_937,In_945);
or U3079 (N_3079,In_186,In_419);
nand U3080 (N_3080,In_579,In_354);
xor U3081 (N_3081,In_401,In_42);
and U3082 (N_3082,In_420,In_382);
nor U3083 (N_3083,In_803,In_579);
nand U3084 (N_3084,In_63,In_973);
nor U3085 (N_3085,In_518,In_33);
nor U3086 (N_3086,In_968,In_124);
nand U3087 (N_3087,In_314,In_918);
nor U3088 (N_3088,In_918,In_150);
nand U3089 (N_3089,In_596,In_963);
nor U3090 (N_3090,In_141,In_153);
nand U3091 (N_3091,In_16,In_202);
nand U3092 (N_3092,In_383,In_228);
nand U3093 (N_3093,In_736,In_104);
nor U3094 (N_3094,In_30,In_3);
and U3095 (N_3095,In_879,In_335);
nand U3096 (N_3096,In_447,In_640);
nand U3097 (N_3097,In_415,In_327);
or U3098 (N_3098,In_693,In_222);
xor U3099 (N_3099,In_349,In_17);
nor U3100 (N_3100,In_762,In_541);
and U3101 (N_3101,In_484,In_445);
xnor U3102 (N_3102,In_61,In_793);
and U3103 (N_3103,In_4,In_596);
nand U3104 (N_3104,In_263,In_996);
nor U3105 (N_3105,In_580,In_362);
nor U3106 (N_3106,In_635,In_945);
nor U3107 (N_3107,In_635,In_490);
nor U3108 (N_3108,In_531,In_926);
xor U3109 (N_3109,In_266,In_585);
xor U3110 (N_3110,In_746,In_62);
nor U3111 (N_3111,In_458,In_219);
or U3112 (N_3112,In_596,In_373);
or U3113 (N_3113,In_312,In_177);
nand U3114 (N_3114,In_185,In_812);
nand U3115 (N_3115,In_110,In_801);
nor U3116 (N_3116,In_962,In_422);
or U3117 (N_3117,In_890,In_654);
and U3118 (N_3118,In_889,In_688);
and U3119 (N_3119,In_400,In_692);
nor U3120 (N_3120,In_431,In_0);
nand U3121 (N_3121,In_444,In_471);
or U3122 (N_3122,In_541,In_918);
or U3123 (N_3123,In_872,In_239);
nor U3124 (N_3124,In_520,In_491);
nand U3125 (N_3125,In_220,In_287);
or U3126 (N_3126,In_159,In_944);
nor U3127 (N_3127,In_794,In_689);
nand U3128 (N_3128,In_854,In_147);
or U3129 (N_3129,In_658,In_343);
and U3130 (N_3130,In_890,In_710);
nor U3131 (N_3131,In_679,In_332);
or U3132 (N_3132,In_944,In_10);
nand U3133 (N_3133,In_175,In_768);
and U3134 (N_3134,In_809,In_1);
nor U3135 (N_3135,In_743,In_637);
and U3136 (N_3136,In_135,In_341);
or U3137 (N_3137,In_38,In_899);
xor U3138 (N_3138,In_315,In_374);
and U3139 (N_3139,In_55,In_804);
nor U3140 (N_3140,In_627,In_488);
nand U3141 (N_3141,In_257,In_758);
and U3142 (N_3142,In_656,In_254);
nand U3143 (N_3143,In_941,In_40);
nor U3144 (N_3144,In_987,In_28);
and U3145 (N_3145,In_363,In_806);
nor U3146 (N_3146,In_818,In_519);
nor U3147 (N_3147,In_61,In_367);
nor U3148 (N_3148,In_302,In_938);
or U3149 (N_3149,In_306,In_272);
nor U3150 (N_3150,In_341,In_795);
xor U3151 (N_3151,In_413,In_227);
nor U3152 (N_3152,In_165,In_147);
and U3153 (N_3153,In_39,In_385);
or U3154 (N_3154,In_289,In_929);
xnor U3155 (N_3155,In_824,In_589);
nand U3156 (N_3156,In_663,In_546);
nor U3157 (N_3157,In_601,In_929);
nor U3158 (N_3158,In_298,In_642);
nand U3159 (N_3159,In_819,In_752);
nand U3160 (N_3160,In_189,In_411);
xor U3161 (N_3161,In_852,In_887);
and U3162 (N_3162,In_847,In_366);
and U3163 (N_3163,In_228,In_123);
and U3164 (N_3164,In_295,In_289);
nand U3165 (N_3165,In_867,In_438);
nor U3166 (N_3166,In_974,In_121);
and U3167 (N_3167,In_550,In_189);
nor U3168 (N_3168,In_244,In_124);
and U3169 (N_3169,In_584,In_551);
nand U3170 (N_3170,In_808,In_112);
and U3171 (N_3171,In_415,In_221);
or U3172 (N_3172,In_397,In_311);
and U3173 (N_3173,In_0,In_296);
and U3174 (N_3174,In_498,In_898);
or U3175 (N_3175,In_437,In_372);
nand U3176 (N_3176,In_986,In_96);
or U3177 (N_3177,In_152,In_425);
nand U3178 (N_3178,In_404,In_205);
or U3179 (N_3179,In_743,In_364);
nand U3180 (N_3180,In_332,In_365);
and U3181 (N_3181,In_100,In_623);
or U3182 (N_3182,In_664,In_213);
nand U3183 (N_3183,In_355,In_727);
nor U3184 (N_3184,In_435,In_421);
nor U3185 (N_3185,In_828,In_861);
nand U3186 (N_3186,In_559,In_751);
nand U3187 (N_3187,In_941,In_934);
nor U3188 (N_3188,In_37,In_35);
nand U3189 (N_3189,In_430,In_270);
or U3190 (N_3190,In_935,In_273);
nand U3191 (N_3191,In_86,In_193);
or U3192 (N_3192,In_828,In_907);
or U3193 (N_3193,In_429,In_736);
and U3194 (N_3194,In_41,In_280);
nand U3195 (N_3195,In_814,In_475);
and U3196 (N_3196,In_243,In_266);
and U3197 (N_3197,In_533,In_960);
nand U3198 (N_3198,In_22,In_269);
and U3199 (N_3199,In_460,In_608);
or U3200 (N_3200,In_965,In_204);
and U3201 (N_3201,In_200,In_18);
and U3202 (N_3202,In_637,In_364);
nor U3203 (N_3203,In_209,In_250);
nor U3204 (N_3204,In_851,In_954);
nor U3205 (N_3205,In_86,In_206);
or U3206 (N_3206,In_174,In_531);
nand U3207 (N_3207,In_568,In_987);
xor U3208 (N_3208,In_513,In_383);
and U3209 (N_3209,In_467,In_798);
and U3210 (N_3210,In_856,In_995);
nor U3211 (N_3211,In_674,In_419);
nand U3212 (N_3212,In_264,In_513);
or U3213 (N_3213,In_510,In_166);
nor U3214 (N_3214,In_177,In_856);
or U3215 (N_3215,In_889,In_494);
and U3216 (N_3216,In_742,In_698);
or U3217 (N_3217,In_444,In_414);
or U3218 (N_3218,In_971,In_98);
or U3219 (N_3219,In_331,In_828);
or U3220 (N_3220,In_661,In_276);
or U3221 (N_3221,In_37,In_641);
and U3222 (N_3222,In_916,In_952);
or U3223 (N_3223,In_430,In_806);
and U3224 (N_3224,In_355,In_762);
and U3225 (N_3225,In_251,In_501);
and U3226 (N_3226,In_652,In_614);
or U3227 (N_3227,In_811,In_989);
nor U3228 (N_3228,In_684,In_609);
or U3229 (N_3229,In_273,In_171);
nand U3230 (N_3230,In_348,In_556);
nand U3231 (N_3231,In_380,In_255);
and U3232 (N_3232,In_113,In_423);
nand U3233 (N_3233,In_7,In_383);
or U3234 (N_3234,In_188,In_824);
or U3235 (N_3235,In_576,In_960);
or U3236 (N_3236,In_273,In_766);
or U3237 (N_3237,In_596,In_823);
nand U3238 (N_3238,In_142,In_484);
and U3239 (N_3239,In_808,In_881);
or U3240 (N_3240,In_670,In_586);
nor U3241 (N_3241,In_68,In_147);
nor U3242 (N_3242,In_80,In_576);
nor U3243 (N_3243,In_813,In_118);
and U3244 (N_3244,In_248,In_499);
and U3245 (N_3245,In_275,In_308);
nor U3246 (N_3246,In_383,In_398);
nor U3247 (N_3247,In_94,In_667);
or U3248 (N_3248,In_497,In_798);
and U3249 (N_3249,In_843,In_886);
nand U3250 (N_3250,In_472,In_352);
or U3251 (N_3251,In_938,In_275);
and U3252 (N_3252,In_454,In_108);
or U3253 (N_3253,In_664,In_190);
or U3254 (N_3254,In_166,In_437);
and U3255 (N_3255,In_65,In_632);
xor U3256 (N_3256,In_548,In_665);
and U3257 (N_3257,In_145,In_428);
nor U3258 (N_3258,In_55,In_578);
nor U3259 (N_3259,In_317,In_223);
nand U3260 (N_3260,In_733,In_917);
nand U3261 (N_3261,In_117,In_360);
nand U3262 (N_3262,In_511,In_509);
or U3263 (N_3263,In_39,In_906);
or U3264 (N_3264,In_751,In_62);
and U3265 (N_3265,In_577,In_645);
nand U3266 (N_3266,In_199,In_542);
nor U3267 (N_3267,In_916,In_835);
and U3268 (N_3268,In_116,In_622);
and U3269 (N_3269,In_677,In_55);
nand U3270 (N_3270,In_600,In_302);
nand U3271 (N_3271,In_103,In_590);
nand U3272 (N_3272,In_528,In_592);
and U3273 (N_3273,In_53,In_417);
or U3274 (N_3274,In_593,In_913);
and U3275 (N_3275,In_304,In_700);
xor U3276 (N_3276,In_921,In_513);
nor U3277 (N_3277,In_354,In_125);
and U3278 (N_3278,In_400,In_955);
and U3279 (N_3279,In_378,In_187);
nand U3280 (N_3280,In_485,In_384);
or U3281 (N_3281,In_913,In_635);
and U3282 (N_3282,In_576,In_0);
nor U3283 (N_3283,In_85,In_879);
and U3284 (N_3284,In_749,In_243);
and U3285 (N_3285,In_761,In_461);
nand U3286 (N_3286,In_581,In_424);
nand U3287 (N_3287,In_945,In_408);
or U3288 (N_3288,In_875,In_44);
nor U3289 (N_3289,In_895,In_799);
or U3290 (N_3290,In_807,In_139);
nand U3291 (N_3291,In_870,In_815);
nand U3292 (N_3292,In_44,In_761);
nor U3293 (N_3293,In_446,In_380);
nor U3294 (N_3294,In_447,In_86);
nor U3295 (N_3295,In_158,In_388);
or U3296 (N_3296,In_807,In_845);
and U3297 (N_3297,In_824,In_567);
nand U3298 (N_3298,In_938,In_51);
or U3299 (N_3299,In_661,In_608);
and U3300 (N_3300,In_711,In_869);
nand U3301 (N_3301,In_706,In_95);
and U3302 (N_3302,In_28,In_35);
or U3303 (N_3303,In_485,In_483);
and U3304 (N_3304,In_190,In_749);
and U3305 (N_3305,In_553,In_868);
nand U3306 (N_3306,In_843,In_75);
or U3307 (N_3307,In_766,In_618);
or U3308 (N_3308,In_376,In_241);
xnor U3309 (N_3309,In_14,In_7);
nor U3310 (N_3310,In_845,In_577);
or U3311 (N_3311,In_618,In_353);
and U3312 (N_3312,In_53,In_640);
nor U3313 (N_3313,In_137,In_489);
and U3314 (N_3314,In_120,In_128);
or U3315 (N_3315,In_825,In_631);
or U3316 (N_3316,In_333,In_976);
nor U3317 (N_3317,In_647,In_385);
nand U3318 (N_3318,In_704,In_862);
and U3319 (N_3319,In_116,In_744);
xnor U3320 (N_3320,In_327,In_927);
nor U3321 (N_3321,In_604,In_842);
nand U3322 (N_3322,In_978,In_864);
nor U3323 (N_3323,In_940,In_407);
nand U3324 (N_3324,In_728,In_74);
nor U3325 (N_3325,In_361,In_571);
xnor U3326 (N_3326,In_35,In_46);
nand U3327 (N_3327,In_514,In_422);
and U3328 (N_3328,In_588,In_913);
nor U3329 (N_3329,In_772,In_54);
nand U3330 (N_3330,In_921,In_983);
and U3331 (N_3331,In_555,In_319);
nor U3332 (N_3332,In_947,In_929);
and U3333 (N_3333,In_43,In_95);
and U3334 (N_3334,In_752,In_497);
nand U3335 (N_3335,In_955,In_783);
nor U3336 (N_3336,In_268,In_315);
or U3337 (N_3337,In_18,In_284);
nand U3338 (N_3338,In_933,In_565);
nor U3339 (N_3339,In_479,In_28);
and U3340 (N_3340,In_539,In_401);
and U3341 (N_3341,In_960,In_390);
nand U3342 (N_3342,In_386,In_888);
and U3343 (N_3343,In_40,In_317);
nand U3344 (N_3344,In_494,In_619);
and U3345 (N_3345,In_753,In_818);
and U3346 (N_3346,In_723,In_440);
or U3347 (N_3347,In_622,In_317);
nand U3348 (N_3348,In_261,In_839);
and U3349 (N_3349,In_576,In_628);
nor U3350 (N_3350,In_919,In_212);
nand U3351 (N_3351,In_580,In_966);
nand U3352 (N_3352,In_691,In_509);
or U3353 (N_3353,In_624,In_374);
and U3354 (N_3354,In_731,In_516);
or U3355 (N_3355,In_642,In_143);
or U3356 (N_3356,In_540,In_43);
and U3357 (N_3357,In_350,In_153);
and U3358 (N_3358,In_16,In_128);
nand U3359 (N_3359,In_194,In_627);
and U3360 (N_3360,In_414,In_119);
nor U3361 (N_3361,In_663,In_246);
and U3362 (N_3362,In_396,In_839);
nand U3363 (N_3363,In_980,In_21);
xor U3364 (N_3364,In_678,In_105);
nand U3365 (N_3365,In_630,In_260);
nor U3366 (N_3366,In_614,In_232);
or U3367 (N_3367,In_518,In_623);
and U3368 (N_3368,In_683,In_265);
nand U3369 (N_3369,In_972,In_792);
and U3370 (N_3370,In_794,In_511);
or U3371 (N_3371,In_363,In_958);
nand U3372 (N_3372,In_791,In_144);
or U3373 (N_3373,In_796,In_875);
and U3374 (N_3374,In_953,In_993);
or U3375 (N_3375,In_894,In_57);
nand U3376 (N_3376,In_292,In_288);
nor U3377 (N_3377,In_148,In_372);
nand U3378 (N_3378,In_808,In_580);
nor U3379 (N_3379,In_261,In_690);
nor U3380 (N_3380,In_766,In_236);
or U3381 (N_3381,In_940,In_519);
nor U3382 (N_3382,In_35,In_189);
or U3383 (N_3383,In_898,In_912);
nor U3384 (N_3384,In_320,In_147);
and U3385 (N_3385,In_494,In_184);
or U3386 (N_3386,In_392,In_269);
nor U3387 (N_3387,In_462,In_600);
or U3388 (N_3388,In_168,In_775);
nand U3389 (N_3389,In_246,In_111);
and U3390 (N_3390,In_267,In_985);
or U3391 (N_3391,In_163,In_477);
nor U3392 (N_3392,In_352,In_828);
or U3393 (N_3393,In_640,In_168);
or U3394 (N_3394,In_11,In_418);
or U3395 (N_3395,In_226,In_393);
nand U3396 (N_3396,In_385,In_708);
nand U3397 (N_3397,In_668,In_632);
nand U3398 (N_3398,In_460,In_378);
nor U3399 (N_3399,In_134,In_752);
nand U3400 (N_3400,In_53,In_998);
and U3401 (N_3401,In_396,In_69);
nand U3402 (N_3402,In_866,In_905);
xor U3403 (N_3403,In_576,In_24);
nor U3404 (N_3404,In_631,In_588);
or U3405 (N_3405,In_842,In_582);
nor U3406 (N_3406,In_472,In_720);
or U3407 (N_3407,In_219,In_260);
nor U3408 (N_3408,In_749,In_235);
or U3409 (N_3409,In_795,In_717);
or U3410 (N_3410,In_392,In_558);
nor U3411 (N_3411,In_676,In_224);
and U3412 (N_3412,In_830,In_271);
nand U3413 (N_3413,In_675,In_727);
nand U3414 (N_3414,In_341,In_31);
and U3415 (N_3415,In_441,In_146);
and U3416 (N_3416,In_183,In_606);
and U3417 (N_3417,In_643,In_433);
nor U3418 (N_3418,In_447,In_569);
nor U3419 (N_3419,In_436,In_651);
nand U3420 (N_3420,In_716,In_835);
nand U3421 (N_3421,In_625,In_17);
nand U3422 (N_3422,In_670,In_106);
nor U3423 (N_3423,In_572,In_492);
nand U3424 (N_3424,In_34,In_247);
nand U3425 (N_3425,In_146,In_959);
nand U3426 (N_3426,In_285,In_831);
nand U3427 (N_3427,In_518,In_738);
or U3428 (N_3428,In_265,In_488);
and U3429 (N_3429,In_610,In_0);
or U3430 (N_3430,In_233,In_876);
or U3431 (N_3431,In_999,In_919);
nor U3432 (N_3432,In_536,In_202);
or U3433 (N_3433,In_359,In_577);
nand U3434 (N_3434,In_888,In_842);
and U3435 (N_3435,In_844,In_839);
xnor U3436 (N_3436,In_201,In_933);
nor U3437 (N_3437,In_248,In_323);
or U3438 (N_3438,In_220,In_731);
nor U3439 (N_3439,In_805,In_4);
and U3440 (N_3440,In_946,In_728);
nor U3441 (N_3441,In_295,In_537);
nand U3442 (N_3442,In_952,In_312);
or U3443 (N_3443,In_322,In_958);
and U3444 (N_3444,In_588,In_324);
nor U3445 (N_3445,In_864,In_628);
nand U3446 (N_3446,In_659,In_185);
and U3447 (N_3447,In_458,In_947);
nand U3448 (N_3448,In_738,In_237);
nand U3449 (N_3449,In_44,In_342);
nor U3450 (N_3450,In_716,In_928);
and U3451 (N_3451,In_462,In_965);
and U3452 (N_3452,In_153,In_722);
or U3453 (N_3453,In_500,In_41);
or U3454 (N_3454,In_848,In_59);
or U3455 (N_3455,In_579,In_130);
nand U3456 (N_3456,In_650,In_431);
or U3457 (N_3457,In_76,In_747);
or U3458 (N_3458,In_386,In_793);
and U3459 (N_3459,In_148,In_955);
nor U3460 (N_3460,In_611,In_27);
or U3461 (N_3461,In_229,In_114);
nand U3462 (N_3462,In_778,In_605);
or U3463 (N_3463,In_576,In_618);
nand U3464 (N_3464,In_460,In_649);
and U3465 (N_3465,In_955,In_479);
nor U3466 (N_3466,In_760,In_213);
or U3467 (N_3467,In_221,In_173);
or U3468 (N_3468,In_629,In_395);
or U3469 (N_3469,In_28,In_18);
or U3470 (N_3470,In_59,In_813);
and U3471 (N_3471,In_356,In_649);
or U3472 (N_3472,In_322,In_190);
or U3473 (N_3473,In_618,In_993);
or U3474 (N_3474,In_126,In_750);
or U3475 (N_3475,In_889,In_762);
or U3476 (N_3476,In_783,In_639);
xnor U3477 (N_3477,In_696,In_475);
or U3478 (N_3478,In_956,In_781);
and U3479 (N_3479,In_504,In_964);
nand U3480 (N_3480,In_444,In_823);
and U3481 (N_3481,In_479,In_607);
and U3482 (N_3482,In_683,In_11);
nor U3483 (N_3483,In_566,In_393);
nor U3484 (N_3484,In_534,In_775);
or U3485 (N_3485,In_546,In_399);
xor U3486 (N_3486,In_783,In_149);
nor U3487 (N_3487,In_247,In_527);
nor U3488 (N_3488,In_206,In_493);
nor U3489 (N_3489,In_106,In_71);
or U3490 (N_3490,In_966,In_49);
and U3491 (N_3491,In_621,In_634);
nand U3492 (N_3492,In_819,In_645);
nand U3493 (N_3493,In_193,In_743);
nor U3494 (N_3494,In_627,In_654);
or U3495 (N_3495,In_635,In_749);
nor U3496 (N_3496,In_322,In_894);
nand U3497 (N_3497,In_679,In_153);
nor U3498 (N_3498,In_121,In_777);
nand U3499 (N_3499,In_938,In_407);
nand U3500 (N_3500,In_395,In_355);
xor U3501 (N_3501,In_818,In_470);
and U3502 (N_3502,In_275,In_457);
or U3503 (N_3503,In_389,In_476);
or U3504 (N_3504,In_292,In_101);
nor U3505 (N_3505,In_263,In_434);
and U3506 (N_3506,In_980,In_216);
nand U3507 (N_3507,In_8,In_365);
or U3508 (N_3508,In_369,In_969);
nor U3509 (N_3509,In_462,In_860);
and U3510 (N_3510,In_224,In_890);
or U3511 (N_3511,In_576,In_174);
nor U3512 (N_3512,In_622,In_1);
or U3513 (N_3513,In_121,In_373);
and U3514 (N_3514,In_888,In_144);
nand U3515 (N_3515,In_569,In_960);
nand U3516 (N_3516,In_202,In_108);
or U3517 (N_3517,In_813,In_409);
nand U3518 (N_3518,In_519,In_462);
and U3519 (N_3519,In_286,In_748);
nand U3520 (N_3520,In_881,In_339);
nand U3521 (N_3521,In_777,In_502);
or U3522 (N_3522,In_134,In_82);
nor U3523 (N_3523,In_810,In_509);
or U3524 (N_3524,In_54,In_601);
nor U3525 (N_3525,In_313,In_38);
and U3526 (N_3526,In_83,In_807);
nor U3527 (N_3527,In_503,In_936);
or U3528 (N_3528,In_298,In_778);
or U3529 (N_3529,In_569,In_579);
xor U3530 (N_3530,In_172,In_388);
nand U3531 (N_3531,In_8,In_546);
nor U3532 (N_3532,In_985,In_381);
xnor U3533 (N_3533,In_441,In_662);
nor U3534 (N_3534,In_835,In_112);
or U3535 (N_3535,In_96,In_23);
nand U3536 (N_3536,In_490,In_651);
nand U3537 (N_3537,In_175,In_225);
or U3538 (N_3538,In_546,In_958);
and U3539 (N_3539,In_714,In_915);
or U3540 (N_3540,In_508,In_271);
nand U3541 (N_3541,In_74,In_674);
or U3542 (N_3542,In_75,In_821);
nand U3543 (N_3543,In_174,In_529);
or U3544 (N_3544,In_253,In_508);
xnor U3545 (N_3545,In_581,In_100);
nor U3546 (N_3546,In_266,In_49);
or U3547 (N_3547,In_105,In_986);
and U3548 (N_3548,In_728,In_731);
or U3549 (N_3549,In_853,In_313);
and U3550 (N_3550,In_208,In_588);
and U3551 (N_3551,In_773,In_919);
xor U3552 (N_3552,In_651,In_846);
nand U3553 (N_3553,In_913,In_816);
nand U3554 (N_3554,In_284,In_921);
or U3555 (N_3555,In_859,In_40);
nor U3556 (N_3556,In_897,In_13);
nor U3557 (N_3557,In_578,In_170);
and U3558 (N_3558,In_864,In_164);
nand U3559 (N_3559,In_782,In_885);
and U3560 (N_3560,In_730,In_168);
and U3561 (N_3561,In_8,In_978);
or U3562 (N_3562,In_125,In_302);
nor U3563 (N_3563,In_971,In_463);
nand U3564 (N_3564,In_491,In_277);
or U3565 (N_3565,In_831,In_402);
and U3566 (N_3566,In_639,In_591);
nand U3567 (N_3567,In_593,In_21);
nor U3568 (N_3568,In_997,In_884);
nor U3569 (N_3569,In_2,In_866);
nor U3570 (N_3570,In_725,In_388);
and U3571 (N_3571,In_126,In_570);
nor U3572 (N_3572,In_928,In_342);
nor U3573 (N_3573,In_496,In_918);
nand U3574 (N_3574,In_716,In_187);
nand U3575 (N_3575,In_565,In_621);
or U3576 (N_3576,In_907,In_101);
nand U3577 (N_3577,In_521,In_545);
and U3578 (N_3578,In_340,In_569);
nand U3579 (N_3579,In_902,In_719);
and U3580 (N_3580,In_223,In_396);
and U3581 (N_3581,In_302,In_921);
and U3582 (N_3582,In_299,In_807);
nor U3583 (N_3583,In_188,In_24);
or U3584 (N_3584,In_313,In_491);
and U3585 (N_3585,In_302,In_772);
or U3586 (N_3586,In_929,In_682);
and U3587 (N_3587,In_707,In_587);
and U3588 (N_3588,In_764,In_190);
nand U3589 (N_3589,In_504,In_870);
and U3590 (N_3590,In_509,In_402);
nor U3591 (N_3591,In_216,In_239);
or U3592 (N_3592,In_527,In_22);
and U3593 (N_3593,In_235,In_134);
and U3594 (N_3594,In_649,In_567);
nor U3595 (N_3595,In_986,In_100);
nand U3596 (N_3596,In_181,In_590);
nand U3597 (N_3597,In_869,In_293);
nor U3598 (N_3598,In_369,In_157);
or U3599 (N_3599,In_153,In_431);
or U3600 (N_3600,In_223,In_4);
nand U3601 (N_3601,In_101,In_266);
or U3602 (N_3602,In_672,In_498);
nor U3603 (N_3603,In_870,In_720);
and U3604 (N_3604,In_800,In_159);
and U3605 (N_3605,In_312,In_9);
xnor U3606 (N_3606,In_537,In_751);
nand U3607 (N_3607,In_327,In_332);
nand U3608 (N_3608,In_658,In_261);
nor U3609 (N_3609,In_477,In_311);
nor U3610 (N_3610,In_386,In_283);
and U3611 (N_3611,In_576,In_145);
xor U3612 (N_3612,In_294,In_981);
xor U3613 (N_3613,In_472,In_220);
or U3614 (N_3614,In_911,In_994);
nor U3615 (N_3615,In_278,In_437);
nand U3616 (N_3616,In_63,In_13);
nor U3617 (N_3617,In_408,In_454);
or U3618 (N_3618,In_331,In_182);
nand U3619 (N_3619,In_314,In_718);
or U3620 (N_3620,In_714,In_313);
nand U3621 (N_3621,In_534,In_516);
or U3622 (N_3622,In_780,In_336);
and U3623 (N_3623,In_789,In_414);
or U3624 (N_3624,In_142,In_897);
and U3625 (N_3625,In_168,In_684);
or U3626 (N_3626,In_284,In_661);
nor U3627 (N_3627,In_49,In_421);
and U3628 (N_3628,In_469,In_311);
and U3629 (N_3629,In_764,In_487);
or U3630 (N_3630,In_156,In_964);
nand U3631 (N_3631,In_319,In_612);
nand U3632 (N_3632,In_167,In_999);
nor U3633 (N_3633,In_419,In_433);
or U3634 (N_3634,In_349,In_674);
or U3635 (N_3635,In_709,In_304);
nor U3636 (N_3636,In_152,In_354);
and U3637 (N_3637,In_262,In_766);
or U3638 (N_3638,In_697,In_425);
and U3639 (N_3639,In_681,In_481);
nor U3640 (N_3640,In_703,In_241);
or U3641 (N_3641,In_949,In_7);
nand U3642 (N_3642,In_547,In_430);
nand U3643 (N_3643,In_13,In_865);
or U3644 (N_3644,In_499,In_361);
nand U3645 (N_3645,In_355,In_588);
and U3646 (N_3646,In_412,In_145);
and U3647 (N_3647,In_65,In_627);
nand U3648 (N_3648,In_302,In_168);
nor U3649 (N_3649,In_301,In_765);
and U3650 (N_3650,In_809,In_467);
nand U3651 (N_3651,In_156,In_190);
or U3652 (N_3652,In_517,In_340);
nand U3653 (N_3653,In_461,In_195);
nor U3654 (N_3654,In_254,In_300);
nor U3655 (N_3655,In_709,In_54);
and U3656 (N_3656,In_300,In_821);
nand U3657 (N_3657,In_202,In_493);
and U3658 (N_3658,In_65,In_57);
and U3659 (N_3659,In_884,In_691);
nor U3660 (N_3660,In_542,In_454);
or U3661 (N_3661,In_857,In_697);
nand U3662 (N_3662,In_863,In_453);
nor U3663 (N_3663,In_946,In_747);
and U3664 (N_3664,In_63,In_338);
nor U3665 (N_3665,In_595,In_563);
or U3666 (N_3666,In_950,In_701);
and U3667 (N_3667,In_603,In_337);
and U3668 (N_3668,In_593,In_59);
and U3669 (N_3669,In_215,In_950);
nand U3670 (N_3670,In_224,In_185);
nor U3671 (N_3671,In_528,In_500);
and U3672 (N_3672,In_127,In_155);
nand U3673 (N_3673,In_679,In_897);
and U3674 (N_3674,In_252,In_32);
or U3675 (N_3675,In_324,In_867);
nand U3676 (N_3676,In_975,In_744);
or U3677 (N_3677,In_893,In_754);
nor U3678 (N_3678,In_118,In_283);
nor U3679 (N_3679,In_523,In_246);
nand U3680 (N_3680,In_696,In_770);
or U3681 (N_3681,In_611,In_872);
or U3682 (N_3682,In_386,In_987);
nand U3683 (N_3683,In_883,In_911);
and U3684 (N_3684,In_827,In_541);
or U3685 (N_3685,In_684,In_765);
or U3686 (N_3686,In_518,In_5);
or U3687 (N_3687,In_182,In_610);
nor U3688 (N_3688,In_791,In_225);
nor U3689 (N_3689,In_502,In_501);
nor U3690 (N_3690,In_842,In_344);
nor U3691 (N_3691,In_569,In_514);
or U3692 (N_3692,In_214,In_343);
xnor U3693 (N_3693,In_492,In_347);
and U3694 (N_3694,In_549,In_551);
nand U3695 (N_3695,In_260,In_133);
or U3696 (N_3696,In_500,In_593);
or U3697 (N_3697,In_76,In_167);
nor U3698 (N_3698,In_707,In_970);
or U3699 (N_3699,In_791,In_854);
nand U3700 (N_3700,In_895,In_453);
xor U3701 (N_3701,In_354,In_959);
nand U3702 (N_3702,In_630,In_919);
and U3703 (N_3703,In_118,In_612);
and U3704 (N_3704,In_29,In_600);
or U3705 (N_3705,In_76,In_964);
nor U3706 (N_3706,In_393,In_702);
or U3707 (N_3707,In_954,In_381);
or U3708 (N_3708,In_227,In_7);
and U3709 (N_3709,In_686,In_960);
or U3710 (N_3710,In_534,In_109);
nor U3711 (N_3711,In_431,In_855);
or U3712 (N_3712,In_853,In_975);
and U3713 (N_3713,In_922,In_873);
and U3714 (N_3714,In_177,In_212);
and U3715 (N_3715,In_225,In_758);
nor U3716 (N_3716,In_917,In_494);
and U3717 (N_3717,In_491,In_379);
and U3718 (N_3718,In_743,In_59);
nor U3719 (N_3719,In_426,In_445);
nor U3720 (N_3720,In_873,In_418);
nor U3721 (N_3721,In_335,In_709);
and U3722 (N_3722,In_425,In_979);
and U3723 (N_3723,In_857,In_888);
and U3724 (N_3724,In_739,In_309);
or U3725 (N_3725,In_892,In_58);
nand U3726 (N_3726,In_577,In_165);
or U3727 (N_3727,In_580,In_337);
and U3728 (N_3728,In_433,In_170);
or U3729 (N_3729,In_5,In_842);
nor U3730 (N_3730,In_429,In_276);
or U3731 (N_3731,In_124,In_4);
or U3732 (N_3732,In_209,In_287);
nand U3733 (N_3733,In_191,In_162);
nand U3734 (N_3734,In_984,In_757);
nor U3735 (N_3735,In_800,In_945);
and U3736 (N_3736,In_661,In_957);
and U3737 (N_3737,In_881,In_604);
nand U3738 (N_3738,In_771,In_779);
and U3739 (N_3739,In_394,In_231);
and U3740 (N_3740,In_181,In_225);
or U3741 (N_3741,In_61,In_947);
or U3742 (N_3742,In_595,In_781);
nor U3743 (N_3743,In_259,In_915);
nand U3744 (N_3744,In_359,In_459);
nor U3745 (N_3745,In_771,In_25);
or U3746 (N_3746,In_6,In_136);
or U3747 (N_3747,In_853,In_265);
nand U3748 (N_3748,In_568,In_85);
nand U3749 (N_3749,In_3,In_711);
or U3750 (N_3750,In_108,In_651);
and U3751 (N_3751,In_707,In_647);
or U3752 (N_3752,In_384,In_902);
nor U3753 (N_3753,In_558,In_771);
xnor U3754 (N_3754,In_49,In_532);
or U3755 (N_3755,In_787,In_138);
and U3756 (N_3756,In_827,In_284);
and U3757 (N_3757,In_818,In_427);
xor U3758 (N_3758,In_699,In_508);
nand U3759 (N_3759,In_986,In_639);
or U3760 (N_3760,In_842,In_195);
nand U3761 (N_3761,In_694,In_490);
nor U3762 (N_3762,In_346,In_14);
or U3763 (N_3763,In_226,In_995);
nand U3764 (N_3764,In_459,In_933);
or U3765 (N_3765,In_477,In_670);
or U3766 (N_3766,In_769,In_511);
nand U3767 (N_3767,In_900,In_902);
xor U3768 (N_3768,In_850,In_70);
nor U3769 (N_3769,In_352,In_280);
nor U3770 (N_3770,In_77,In_578);
and U3771 (N_3771,In_187,In_376);
nand U3772 (N_3772,In_590,In_242);
nand U3773 (N_3773,In_121,In_229);
nand U3774 (N_3774,In_724,In_103);
or U3775 (N_3775,In_728,In_475);
nor U3776 (N_3776,In_682,In_646);
or U3777 (N_3777,In_457,In_912);
and U3778 (N_3778,In_651,In_917);
nor U3779 (N_3779,In_86,In_330);
or U3780 (N_3780,In_870,In_855);
xor U3781 (N_3781,In_245,In_566);
xnor U3782 (N_3782,In_112,In_185);
nor U3783 (N_3783,In_747,In_204);
or U3784 (N_3784,In_958,In_462);
nor U3785 (N_3785,In_654,In_36);
nor U3786 (N_3786,In_326,In_873);
and U3787 (N_3787,In_534,In_211);
or U3788 (N_3788,In_349,In_69);
nand U3789 (N_3789,In_618,In_493);
or U3790 (N_3790,In_578,In_19);
xnor U3791 (N_3791,In_904,In_348);
and U3792 (N_3792,In_536,In_362);
nor U3793 (N_3793,In_966,In_472);
and U3794 (N_3794,In_744,In_219);
or U3795 (N_3795,In_333,In_512);
or U3796 (N_3796,In_585,In_436);
and U3797 (N_3797,In_787,In_551);
nor U3798 (N_3798,In_707,In_458);
nand U3799 (N_3799,In_990,In_339);
nor U3800 (N_3800,In_519,In_682);
and U3801 (N_3801,In_217,In_47);
or U3802 (N_3802,In_782,In_682);
or U3803 (N_3803,In_968,In_971);
nor U3804 (N_3804,In_311,In_714);
nor U3805 (N_3805,In_167,In_409);
or U3806 (N_3806,In_343,In_188);
or U3807 (N_3807,In_813,In_90);
and U3808 (N_3808,In_562,In_912);
nor U3809 (N_3809,In_661,In_435);
nand U3810 (N_3810,In_706,In_698);
nor U3811 (N_3811,In_23,In_612);
nor U3812 (N_3812,In_114,In_921);
xnor U3813 (N_3813,In_73,In_865);
nor U3814 (N_3814,In_133,In_693);
xnor U3815 (N_3815,In_507,In_159);
and U3816 (N_3816,In_584,In_697);
nor U3817 (N_3817,In_426,In_390);
nand U3818 (N_3818,In_238,In_790);
nand U3819 (N_3819,In_656,In_141);
nor U3820 (N_3820,In_991,In_557);
and U3821 (N_3821,In_773,In_139);
nand U3822 (N_3822,In_31,In_193);
or U3823 (N_3823,In_618,In_140);
or U3824 (N_3824,In_145,In_566);
nand U3825 (N_3825,In_93,In_184);
nand U3826 (N_3826,In_724,In_648);
or U3827 (N_3827,In_963,In_845);
and U3828 (N_3828,In_87,In_254);
or U3829 (N_3829,In_421,In_532);
or U3830 (N_3830,In_75,In_538);
or U3831 (N_3831,In_374,In_67);
nand U3832 (N_3832,In_321,In_457);
and U3833 (N_3833,In_684,In_855);
nor U3834 (N_3834,In_654,In_11);
nand U3835 (N_3835,In_545,In_863);
nand U3836 (N_3836,In_579,In_536);
or U3837 (N_3837,In_912,In_245);
and U3838 (N_3838,In_224,In_378);
nand U3839 (N_3839,In_256,In_259);
nor U3840 (N_3840,In_726,In_778);
nand U3841 (N_3841,In_538,In_97);
xor U3842 (N_3842,In_214,In_998);
nand U3843 (N_3843,In_226,In_721);
and U3844 (N_3844,In_21,In_940);
nand U3845 (N_3845,In_142,In_900);
or U3846 (N_3846,In_647,In_297);
or U3847 (N_3847,In_5,In_462);
nand U3848 (N_3848,In_252,In_567);
or U3849 (N_3849,In_236,In_428);
nor U3850 (N_3850,In_531,In_641);
nor U3851 (N_3851,In_293,In_699);
and U3852 (N_3852,In_623,In_74);
or U3853 (N_3853,In_15,In_945);
nor U3854 (N_3854,In_84,In_896);
or U3855 (N_3855,In_189,In_783);
or U3856 (N_3856,In_348,In_231);
or U3857 (N_3857,In_981,In_399);
nor U3858 (N_3858,In_373,In_325);
and U3859 (N_3859,In_311,In_855);
nor U3860 (N_3860,In_748,In_983);
or U3861 (N_3861,In_361,In_166);
and U3862 (N_3862,In_442,In_118);
nor U3863 (N_3863,In_478,In_786);
or U3864 (N_3864,In_707,In_99);
nor U3865 (N_3865,In_173,In_898);
nand U3866 (N_3866,In_800,In_217);
or U3867 (N_3867,In_591,In_439);
nor U3868 (N_3868,In_773,In_412);
or U3869 (N_3869,In_390,In_368);
or U3870 (N_3870,In_75,In_349);
nand U3871 (N_3871,In_921,In_122);
or U3872 (N_3872,In_284,In_129);
nand U3873 (N_3873,In_764,In_119);
xnor U3874 (N_3874,In_969,In_360);
and U3875 (N_3875,In_726,In_708);
or U3876 (N_3876,In_354,In_246);
nor U3877 (N_3877,In_196,In_466);
nand U3878 (N_3878,In_945,In_915);
nor U3879 (N_3879,In_855,In_426);
and U3880 (N_3880,In_746,In_923);
and U3881 (N_3881,In_685,In_120);
nor U3882 (N_3882,In_837,In_77);
and U3883 (N_3883,In_881,In_399);
nor U3884 (N_3884,In_47,In_958);
nand U3885 (N_3885,In_688,In_583);
nand U3886 (N_3886,In_522,In_671);
nand U3887 (N_3887,In_323,In_137);
and U3888 (N_3888,In_755,In_71);
nand U3889 (N_3889,In_771,In_780);
and U3890 (N_3890,In_539,In_803);
or U3891 (N_3891,In_840,In_256);
nand U3892 (N_3892,In_593,In_539);
nand U3893 (N_3893,In_854,In_855);
and U3894 (N_3894,In_753,In_814);
nor U3895 (N_3895,In_268,In_391);
or U3896 (N_3896,In_66,In_646);
nor U3897 (N_3897,In_277,In_872);
and U3898 (N_3898,In_772,In_899);
and U3899 (N_3899,In_484,In_815);
nor U3900 (N_3900,In_873,In_33);
nor U3901 (N_3901,In_852,In_499);
or U3902 (N_3902,In_467,In_653);
nor U3903 (N_3903,In_802,In_839);
xor U3904 (N_3904,In_939,In_167);
nor U3905 (N_3905,In_535,In_252);
xor U3906 (N_3906,In_144,In_275);
nor U3907 (N_3907,In_282,In_969);
and U3908 (N_3908,In_818,In_924);
nand U3909 (N_3909,In_950,In_929);
or U3910 (N_3910,In_655,In_125);
nand U3911 (N_3911,In_583,In_928);
nand U3912 (N_3912,In_979,In_447);
or U3913 (N_3913,In_606,In_474);
or U3914 (N_3914,In_963,In_518);
nor U3915 (N_3915,In_81,In_43);
or U3916 (N_3916,In_565,In_828);
and U3917 (N_3917,In_372,In_829);
nand U3918 (N_3918,In_612,In_909);
and U3919 (N_3919,In_194,In_595);
or U3920 (N_3920,In_976,In_812);
and U3921 (N_3921,In_537,In_924);
nor U3922 (N_3922,In_24,In_644);
and U3923 (N_3923,In_330,In_857);
nor U3924 (N_3924,In_886,In_54);
nand U3925 (N_3925,In_95,In_680);
nor U3926 (N_3926,In_282,In_772);
or U3927 (N_3927,In_239,In_916);
nand U3928 (N_3928,In_574,In_482);
nor U3929 (N_3929,In_379,In_536);
nand U3930 (N_3930,In_872,In_845);
and U3931 (N_3931,In_798,In_652);
nor U3932 (N_3932,In_629,In_517);
or U3933 (N_3933,In_663,In_65);
and U3934 (N_3934,In_402,In_938);
and U3935 (N_3935,In_913,In_34);
and U3936 (N_3936,In_72,In_200);
nand U3937 (N_3937,In_347,In_916);
and U3938 (N_3938,In_231,In_740);
nor U3939 (N_3939,In_109,In_685);
or U3940 (N_3940,In_54,In_768);
or U3941 (N_3941,In_750,In_472);
or U3942 (N_3942,In_400,In_864);
nor U3943 (N_3943,In_737,In_25);
nor U3944 (N_3944,In_596,In_387);
and U3945 (N_3945,In_610,In_444);
nor U3946 (N_3946,In_82,In_922);
or U3947 (N_3947,In_899,In_757);
or U3948 (N_3948,In_834,In_729);
and U3949 (N_3949,In_110,In_708);
nor U3950 (N_3950,In_65,In_782);
or U3951 (N_3951,In_516,In_92);
nand U3952 (N_3952,In_73,In_358);
xnor U3953 (N_3953,In_545,In_399);
nand U3954 (N_3954,In_212,In_653);
nor U3955 (N_3955,In_413,In_777);
or U3956 (N_3956,In_866,In_974);
nand U3957 (N_3957,In_720,In_935);
and U3958 (N_3958,In_404,In_807);
and U3959 (N_3959,In_16,In_888);
or U3960 (N_3960,In_391,In_907);
and U3961 (N_3961,In_584,In_812);
and U3962 (N_3962,In_777,In_490);
xor U3963 (N_3963,In_584,In_848);
and U3964 (N_3964,In_205,In_189);
or U3965 (N_3965,In_951,In_147);
and U3966 (N_3966,In_575,In_425);
or U3967 (N_3967,In_169,In_554);
xnor U3968 (N_3968,In_543,In_235);
nor U3969 (N_3969,In_627,In_108);
or U3970 (N_3970,In_74,In_775);
nor U3971 (N_3971,In_893,In_426);
or U3972 (N_3972,In_233,In_512);
or U3973 (N_3973,In_82,In_375);
nand U3974 (N_3974,In_955,In_52);
nand U3975 (N_3975,In_584,In_732);
and U3976 (N_3976,In_68,In_161);
or U3977 (N_3977,In_189,In_243);
nor U3978 (N_3978,In_423,In_28);
and U3979 (N_3979,In_91,In_61);
and U3980 (N_3980,In_374,In_992);
and U3981 (N_3981,In_571,In_234);
and U3982 (N_3982,In_173,In_137);
xor U3983 (N_3983,In_244,In_966);
or U3984 (N_3984,In_376,In_634);
nand U3985 (N_3985,In_366,In_374);
or U3986 (N_3986,In_563,In_676);
and U3987 (N_3987,In_26,In_741);
or U3988 (N_3988,In_295,In_635);
or U3989 (N_3989,In_691,In_225);
nor U3990 (N_3990,In_795,In_246);
xnor U3991 (N_3991,In_358,In_145);
nor U3992 (N_3992,In_531,In_14);
nor U3993 (N_3993,In_584,In_901);
nand U3994 (N_3994,In_177,In_73);
or U3995 (N_3995,In_832,In_381);
or U3996 (N_3996,In_162,In_384);
and U3997 (N_3997,In_835,In_70);
nor U3998 (N_3998,In_178,In_883);
nor U3999 (N_3999,In_687,In_473);
nand U4000 (N_4000,In_388,In_126);
nand U4001 (N_4001,In_133,In_849);
or U4002 (N_4002,In_445,In_890);
nor U4003 (N_4003,In_787,In_841);
nor U4004 (N_4004,In_897,In_592);
or U4005 (N_4005,In_174,In_673);
nor U4006 (N_4006,In_598,In_497);
or U4007 (N_4007,In_33,In_263);
nand U4008 (N_4008,In_669,In_920);
or U4009 (N_4009,In_817,In_802);
nor U4010 (N_4010,In_473,In_62);
or U4011 (N_4011,In_276,In_475);
or U4012 (N_4012,In_766,In_19);
nand U4013 (N_4013,In_475,In_368);
nand U4014 (N_4014,In_620,In_22);
nor U4015 (N_4015,In_649,In_795);
nor U4016 (N_4016,In_658,In_690);
or U4017 (N_4017,In_52,In_578);
or U4018 (N_4018,In_133,In_30);
nand U4019 (N_4019,In_672,In_369);
and U4020 (N_4020,In_601,In_493);
or U4021 (N_4021,In_235,In_436);
nor U4022 (N_4022,In_949,In_486);
nor U4023 (N_4023,In_841,In_529);
nor U4024 (N_4024,In_856,In_491);
nand U4025 (N_4025,In_64,In_472);
nor U4026 (N_4026,In_467,In_491);
nand U4027 (N_4027,In_460,In_91);
nand U4028 (N_4028,In_158,In_176);
nor U4029 (N_4029,In_295,In_762);
nand U4030 (N_4030,In_472,In_498);
nand U4031 (N_4031,In_221,In_708);
or U4032 (N_4032,In_916,In_582);
and U4033 (N_4033,In_300,In_151);
nand U4034 (N_4034,In_325,In_802);
nor U4035 (N_4035,In_569,In_217);
or U4036 (N_4036,In_178,In_361);
nor U4037 (N_4037,In_273,In_651);
nor U4038 (N_4038,In_452,In_84);
or U4039 (N_4039,In_837,In_521);
nand U4040 (N_4040,In_189,In_855);
nand U4041 (N_4041,In_470,In_432);
and U4042 (N_4042,In_422,In_922);
and U4043 (N_4043,In_673,In_572);
and U4044 (N_4044,In_660,In_493);
and U4045 (N_4045,In_841,In_933);
and U4046 (N_4046,In_879,In_306);
and U4047 (N_4047,In_592,In_412);
or U4048 (N_4048,In_214,In_153);
nand U4049 (N_4049,In_547,In_389);
or U4050 (N_4050,In_631,In_308);
nand U4051 (N_4051,In_167,In_519);
or U4052 (N_4052,In_213,In_881);
or U4053 (N_4053,In_417,In_117);
or U4054 (N_4054,In_793,In_267);
or U4055 (N_4055,In_10,In_288);
nor U4056 (N_4056,In_613,In_376);
nand U4057 (N_4057,In_995,In_387);
xor U4058 (N_4058,In_775,In_448);
nor U4059 (N_4059,In_816,In_953);
or U4060 (N_4060,In_818,In_401);
nor U4061 (N_4061,In_569,In_98);
nand U4062 (N_4062,In_969,In_885);
nor U4063 (N_4063,In_484,In_424);
nand U4064 (N_4064,In_780,In_946);
and U4065 (N_4065,In_492,In_756);
nor U4066 (N_4066,In_624,In_913);
or U4067 (N_4067,In_408,In_219);
and U4068 (N_4068,In_960,In_397);
or U4069 (N_4069,In_865,In_549);
or U4070 (N_4070,In_409,In_591);
and U4071 (N_4071,In_894,In_696);
nand U4072 (N_4072,In_184,In_723);
or U4073 (N_4073,In_467,In_495);
and U4074 (N_4074,In_576,In_44);
nor U4075 (N_4075,In_132,In_682);
or U4076 (N_4076,In_208,In_503);
nor U4077 (N_4077,In_289,In_47);
and U4078 (N_4078,In_201,In_217);
nand U4079 (N_4079,In_946,In_147);
nand U4080 (N_4080,In_300,In_970);
nor U4081 (N_4081,In_179,In_233);
nand U4082 (N_4082,In_376,In_517);
nand U4083 (N_4083,In_190,In_940);
or U4084 (N_4084,In_931,In_116);
or U4085 (N_4085,In_725,In_817);
nand U4086 (N_4086,In_317,In_539);
nor U4087 (N_4087,In_434,In_613);
nor U4088 (N_4088,In_408,In_670);
and U4089 (N_4089,In_641,In_412);
nand U4090 (N_4090,In_873,In_68);
or U4091 (N_4091,In_177,In_917);
and U4092 (N_4092,In_883,In_360);
and U4093 (N_4093,In_886,In_155);
or U4094 (N_4094,In_552,In_302);
nor U4095 (N_4095,In_22,In_808);
nand U4096 (N_4096,In_501,In_647);
nor U4097 (N_4097,In_447,In_996);
xnor U4098 (N_4098,In_323,In_32);
and U4099 (N_4099,In_371,In_693);
nand U4100 (N_4100,In_361,In_276);
nor U4101 (N_4101,In_47,In_149);
or U4102 (N_4102,In_653,In_576);
nor U4103 (N_4103,In_873,In_488);
nor U4104 (N_4104,In_204,In_339);
nand U4105 (N_4105,In_29,In_453);
nand U4106 (N_4106,In_773,In_559);
nand U4107 (N_4107,In_477,In_884);
nand U4108 (N_4108,In_373,In_798);
and U4109 (N_4109,In_814,In_275);
and U4110 (N_4110,In_452,In_417);
nand U4111 (N_4111,In_961,In_689);
and U4112 (N_4112,In_110,In_14);
nand U4113 (N_4113,In_484,In_825);
or U4114 (N_4114,In_361,In_512);
nand U4115 (N_4115,In_589,In_997);
and U4116 (N_4116,In_138,In_333);
nand U4117 (N_4117,In_429,In_964);
nor U4118 (N_4118,In_169,In_555);
nand U4119 (N_4119,In_140,In_253);
xor U4120 (N_4120,In_498,In_745);
and U4121 (N_4121,In_424,In_86);
nor U4122 (N_4122,In_110,In_146);
or U4123 (N_4123,In_263,In_641);
nand U4124 (N_4124,In_557,In_626);
or U4125 (N_4125,In_681,In_491);
or U4126 (N_4126,In_397,In_919);
and U4127 (N_4127,In_798,In_247);
or U4128 (N_4128,In_112,In_629);
and U4129 (N_4129,In_340,In_283);
nor U4130 (N_4130,In_976,In_912);
nand U4131 (N_4131,In_212,In_451);
and U4132 (N_4132,In_156,In_570);
nand U4133 (N_4133,In_679,In_683);
nand U4134 (N_4134,In_707,In_282);
nand U4135 (N_4135,In_966,In_844);
nor U4136 (N_4136,In_939,In_823);
or U4137 (N_4137,In_33,In_70);
and U4138 (N_4138,In_91,In_876);
or U4139 (N_4139,In_670,In_691);
and U4140 (N_4140,In_794,In_586);
or U4141 (N_4141,In_818,In_629);
xnor U4142 (N_4142,In_179,In_644);
or U4143 (N_4143,In_489,In_23);
nor U4144 (N_4144,In_775,In_183);
nor U4145 (N_4145,In_566,In_865);
nor U4146 (N_4146,In_87,In_77);
or U4147 (N_4147,In_525,In_929);
or U4148 (N_4148,In_757,In_243);
nor U4149 (N_4149,In_861,In_27);
and U4150 (N_4150,In_961,In_196);
and U4151 (N_4151,In_227,In_344);
nand U4152 (N_4152,In_543,In_836);
nor U4153 (N_4153,In_1,In_779);
nand U4154 (N_4154,In_239,In_297);
nor U4155 (N_4155,In_850,In_895);
or U4156 (N_4156,In_813,In_387);
nand U4157 (N_4157,In_7,In_554);
nor U4158 (N_4158,In_110,In_399);
nor U4159 (N_4159,In_5,In_843);
xnor U4160 (N_4160,In_517,In_918);
nand U4161 (N_4161,In_918,In_788);
or U4162 (N_4162,In_406,In_462);
nand U4163 (N_4163,In_392,In_670);
and U4164 (N_4164,In_674,In_620);
nor U4165 (N_4165,In_81,In_47);
xor U4166 (N_4166,In_893,In_761);
or U4167 (N_4167,In_128,In_552);
nand U4168 (N_4168,In_179,In_485);
or U4169 (N_4169,In_216,In_401);
nand U4170 (N_4170,In_983,In_493);
nand U4171 (N_4171,In_638,In_237);
nand U4172 (N_4172,In_179,In_193);
nor U4173 (N_4173,In_32,In_525);
nor U4174 (N_4174,In_934,In_329);
nand U4175 (N_4175,In_100,In_930);
nor U4176 (N_4176,In_155,In_950);
and U4177 (N_4177,In_802,In_20);
or U4178 (N_4178,In_784,In_323);
nor U4179 (N_4179,In_27,In_758);
nor U4180 (N_4180,In_262,In_737);
and U4181 (N_4181,In_423,In_329);
or U4182 (N_4182,In_559,In_493);
and U4183 (N_4183,In_645,In_425);
and U4184 (N_4184,In_620,In_6);
or U4185 (N_4185,In_958,In_985);
or U4186 (N_4186,In_183,In_65);
and U4187 (N_4187,In_93,In_698);
or U4188 (N_4188,In_564,In_379);
and U4189 (N_4189,In_67,In_6);
and U4190 (N_4190,In_910,In_528);
or U4191 (N_4191,In_655,In_296);
or U4192 (N_4192,In_131,In_777);
or U4193 (N_4193,In_840,In_685);
nor U4194 (N_4194,In_273,In_823);
or U4195 (N_4195,In_115,In_191);
or U4196 (N_4196,In_683,In_604);
and U4197 (N_4197,In_339,In_734);
and U4198 (N_4198,In_907,In_530);
nand U4199 (N_4199,In_497,In_2);
and U4200 (N_4200,In_92,In_833);
nor U4201 (N_4201,In_236,In_372);
nand U4202 (N_4202,In_281,In_416);
nor U4203 (N_4203,In_186,In_343);
or U4204 (N_4204,In_879,In_336);
and U4205 (N_4205,In_335,In_912);
or U4206 (N_4206,In_850,In_872);
nand U4207 (N_4207,In_904,In_268);
or U4208 (N_4208,In_724,In_997);
nor U4209 (N_4209,In_771,In_884);
nand U4210 (N_4210,In_690,In_789);
nand U4211 (N_4211,In_793,In_683);
and U4212 (N_4212,In_73,In_87);
or U4213 (N_4213,In_380,In_228);
or U4214 (N_4214,In_404,In_112);
nor U4215 (N_4215,In_356,In_831);
and U4216 (N_4216,In_680,In_900);
nand U4217 (N_4217,In_228,In_272);
and U4218 (N_4218,In_661,In_614);
nand U4219 (N_4219,In_451,In_180);
and U4220 (N_4220,In_541,In_17);
nand U4221 (N_4221,In_955,In_435);
nand U4222 (N_4222,In_806,In_520);
or U4223 (N_4223,In_883,In_490);
or U4224 (N_4224,In_268,In_531);
or U4225 (N_4225,In_972,In_80);
nand U4226 (N_4226,In_842,In_824);
and U4227 (N_4227,In_926,In_591);
and U4228 (N_4228,In_507,In_336);
or U4229 (N_4229,In_177,In_781);
or U4230 (N_4230,In_576,In_335);
nor U4231 (N_4231,In_332,In_83);
nand U4232 (N_4232,In_491,In_710);
nand U4233 (N_4233,In_841,In_551);
or U4234 (N_4234,In_738,In_836);
and U4235 (N_4235,In_6,In_23);
or U4236 (N_4236,In_408,In_472);
nand U4237 (N_4237,In_892,In_563);
or U4238 (N_4238,In_504,In_425);
nand U4239 (N_4239,In_256,In_352);
and U4240 (N_4240,In_548,In_168);
nand U4241 (N_4241,In_142,In_586);
and U4242 (N_4242,In_258,In_615);
or U4243 (N_4243,In_987,In_71);
nand U4244 (N_4244,In_487,In_128);
nand U4245 (N_4245,In_701,In_440);
and U4246 (N_4246,In_951,In_635);
nand U4247 (N_4247,In_431,In_999);
or U4248 (N_4248,In_482,In_881);
or U4249 (N_4249,In_507,In_591);
and U4250 (N_4250,In_485,In_686);
nand U4251 (N_4251,In_549,In_307);
nor U4252 (N_4252,In_842,In_684);
and U4253 (N_4253,In_869,In_643);
nor U4254 (N_4254,In_477,In_472);
or U4255 (N_4255,In_923,In_423);
nor U4256 (N_4256,In_854,In_198);
xnor U4257 (N_4257,In_902,In_464);
and U4258 (N_4258,In_900,In_127);
and U4259 (N_4259,In_598,In_878);
nand U4260 (N_4260,In_636,In_626);
and U4261 (N_4261,In_786,In_275);
and U4262 (N_4262,In_480,In_967);
nand U4263 (N_4263,In_555,In_83);
nand U4264 (N_4264,In_996,In_498);
and U4265 (N_4265,In_368,In_745);
nand U4266 (N_4266,In_489,In_267);
nor U4267 (N_4267,In_102,In_193);
nand U4268 (N_4268,In_368,In_377);
and U4269 (N_4269,In_633,In_895);
nand U4270 (N_4270,In_33,In_235);
nor U4271 (N_4271,In_105,In_174);
or U4272 (N_4272,In_681,In_304);
or U4273 (N_4273,In_492,In_274);
nand U4274 (N_4274,In_108,In_103);
nor U4275 (N_4275,In_486,In_453);
and U4276 (N_4276,In_261,In_313);
and U4277 (N_4277,In_819,In_682);
nor U4278 (N_4278,In_882,In_962);
and U4279 (N_4279,In_366,In_363);
and U4280 (N_4280,In_267,In_735);
nor U4281 (N_4281,In_301,In_955);
or U4282 (N_4282,In_393,In_478);
or U4283 (N_4283,In_285,In_594);
or U4284 (N_4284,In_840,In_740);
nor U4285 (N_4285,In_234,In_966);
and U4286 (N_4286,In_131,In_389);
xor U4287 (N_4287,In_405,In_520);
or U4288 (N_4288,In_460,In_214);
nand U4289 (N_4289,In_257,In_487);
and U4290 (N_4290,In_997,In_992);
nand U4291 (N_4291,In_749,In_800);
nand U4292 (N_4292,In_374,In_835);
or U4293 (N_4293,In_212,In_536);
or U4294 (N_4294,In_922,In_905);
or U4295 (N_4295,In_108,In_269);
or U4296 (N_4296,In_617,In_603);
nand U4297 (N_4297,In_250,In_698);
and U4298 (N_4298,In_892,In_588);
nand U4299 (N_4299,In_552,In_884);
and U4300 (N_4300,In_528,In_448);
nand U4301 (N_4301,In_304,In_365);
or U4302 (N_4302,In_661,In_553);
or U4303 (N_4303,In_209,In_215);
or U4304 (N_4304,In_284,In_667);
nor U4305 (N_4305,In_426,In_825);
nor U4306 (N_4306,In_867,In_583);
nor U4307 (N_4307,In_878,In_943);
nor U4308 (N_4308,In_276,In_465);
or U4309 (N_4309,In_69,In_820);
nand U4310 (N_4310,In_862,In_629);
xnor U4311 (N_4311,In_489,In_684);
and U4312 (N_4312,In_815,In_463);
nor U4313 (N_4313,In_463,In_364);
nor U4314 (N_4314,In_148,In_873);
and U4315 (N_4315,In_13,In_461);
or U4316 (N_4316,In_839,In_76);
and U4317 (N_4317,In_952,In_632);
nand U4318 (N_4318,In_682,In_858);
and U4319 (N_4319,In_897,In_613);
and U4320 (N_4320,In_709,In_911);
nand U4321 (N_4321,In_469,In_1);
and U4322 (N_4322,In_586,In_98);
and U4323 (N_4323,In_998,In_522);
and U4324 (N_4324,In_873,In_502);
nand U4325 (N_4325,In_336,In_501);
nand U4326 (N_4326,In_985,In_748);
nor U4327 (N_4327,In_725,In_333);
and U4328 (N_4328,In_588,In_506);
nor U4329 (N_4329,In_370,In_907);
xnor U4330 (N_4330,In_353,In_54);
or U4331 (N_4331,In_747,In_266);
nor U4332 (N_4332,In_562,In_721);
nor U4333 (N_4333,In_264,In_189);
nand U4334 (N_4334,In_826,In_219);
nand U4335 (N_4335,In_971,In_871);
or U4336 (N_4336,In_945,In_335);
nor U4337 (N_4337,In_535,In_383);
or U4338 (N_4338,In_177,In_916);
and U4339 (N_4339,In_420,In_416);
nor U4340 (N_4340,In_614,In_961);
or U4341 (N_4341,In_670,In_723);
nor U4342 (N_4342,In_653,In_625);
nand U4343 (N_4343,In_461,In_626);
or U4344 (N_4344,In_342,In_623);
nand U4345 (N_4345,In_927,In_394);
nor U4346 (N_4346,In_384,In_906);
or U4347 (N_4347,In_245,In_168);
or U4348 (N_4348,In_999,In_61);
and U4349 (N_4349,In_240,In_186);
and U4350 (N_4350,In_315,In_944);
or U4351 (N_4351,In_387,In_774);
or U4352 (N_4352,In_195,In_978);
nand U4353 (N_4353,In_159,In_202);
and U4354 (N_4354,In_372,In_922);
nor U4355 (N_4355,In_363,In_814);
or U4356 (N_4356,In_2,In_234);
nand U4357 (N_4357,In_675,In_30);
nor U4358 (N_4358,In_103,In_425);
or U4359 (N_4359,In_170,In_421);
or U4360 (N_4360,In_183,In_222);
nor U4361 (N_4361,In_379,In_676);
nor U4362 (N_4362,In_632,In_863);
and U4363 (N_4363,In_57,In_704);
or U4364 (N_4364,In_548,In_883);
nor U4365 (N_4365,In_171,In_541);
nor U4366 (N_4366,In_596,In_46);
or U4367 (N_4367,In_163,In_17);
nand U4368 (N_4368,In_228,In_974);
nand U4369 (N_4369,In_193,In_85);
nand U4370 (N_4370,In_749,In_923);
xnor U4371 (N_4371,In_472,In_801);
and U4372 (N_4372,In_122,In_53);
and U4373 (N_4373,In_499,In_84);
or U4374 (N_4374,In_952,In_793);
and U4375 (N_4375,In_368,In_221);
nand U4376 (N_4376,In_589,In_16);
or U4377 (N_4377,In_737,In_605);
and U4378 (N_4378,In_328,In_2);
or U4379 (N_4379,In_900,In_888);
or U4380 (N_4380,In_51,In_968);
nand U4381 (N_4381,In_601,In_553);
or U4382 (N_4382,In_165,In_246);
and U4383 (N_4383,In_527,In_966);
nor U4384 (N_4384,In_277,In_242);
nor U4385 (N_4385,In_21,In_713);
and U4386 (N_4386,In_65,In_135);
or U4387 (N_4387,In_45,In_493);
nand U4388 (N_4388,In_199,In_690);
nor U4389 (N_4389,In_213,In_183);
nor U4390 (N_4390,In_855,In_455);
nor U4391 (N_4391,In_549,In_548);
nand U4392 (N_4392,In_722,In_6);
or U4393 (N_4393,In_141,In_102);
and U4394 (N_4394,In_216,In_146);
or U4395 (N_4395,In_506,In_581);
nor U4396 (N_4396,In_993,In_27);
nand U4397 (N_4397,In_38,In_222);
nand U4398 (N_4398,In_68,In_153);
or U4399 (N_4399,In_322,In_581);
nor U4400 (N_4400,In_347,In_290);
or U4401 (N_4401,In_259,In_840);
nor U4402 (N_4402,In_837,In_934);
or U4403 (N_4403,In_160,In_358);
and U4404 (N_4404,In_694,In_625);
and U4405 (N_4405,In_85,In_124);
nand U4406 (N_4406,In_920,In_215);
or U4407 (N_4407,In_782,In_156);
nand U4408 (N_4408,In_569,In_562);
or U4409 (N_4409,In_364,In_276);
and U4410 (N_4410,In_184,In_174);
and U4411 (N_4411,In_654,In_682);
nor U4412 (N_4412,In_763,In_59);
nor U4413 (N_4413,In_965,In_982);
nor U4414 (N_4414,In_639,In_990);
nand U4415 (N_4415,In_401,In_52);
nand U4416 (N_4416,In_764,In_491);
nand U4417 (N_4417,In_252,In_154);
or U4418 (N_4418,In_341,In_740);
or U4419 (N_4419,In_561,In_252);
nand U4420 (N_4420,In_188,In_579);
nand U4421 (N_4421,In_833,In_908);
nor U4422 (N_4422,In_748,In_352);
or U4423 (N_4423,In_639,In_469);
and U4424 (N_4424,In_623,In_552);
or U4425 (N_4425,In_286,In_290);
or U4426 (N_4426,In_326,In_786);
nand U4427 (N_4427,In_296,In_460);
and U4428 (N_4428,In_606,In_480);
nor U4429 (N_4429,In_87,In_364);
xor U4430 (N_4430,In_305,In_779);
or U4431 (N_4431,In_841,In_645);
or U4432 (N_4432,In_798,In_322);
nor U4433 (N_4433,In_516,In_368);
or U4434 (N_4434,In_76,In_413);
nor U4435 (N_4435,In_714,In_125);
nand U4436 (N_4436,In_722,In_463);
or U4437 (N_4437,In_892,In_286);
or U4438 (N_4438,In_409,In_86);
nand U4439 (N_4439,In_638,In_901);
nand U4440 (N_4440,In_651,In_715);
and U4441 (N_4441,In_128,In_927);
or U4442 (N_4442,In_882,In_369);
nand U4443 (N_4443,In_735,In_231);
nand U4444 (N_4444,In_680,In_764);
xnor U4445 (N_4445,In_307,In_808);
nor U4446 (N_4446,In_336,In_594);
and U4447 (N_4447,In_97,In_686);
nand U4448 (N_4448,In_22,In_471);
nand U4449 (N_4449,In_958,In_362);
and U4450 (N_4450,In_74,In_896);
and U4451 (N_4451,In_140,In_489);
and U4452 (N_4452,In_873,In_117);
and U4453 (N_4453,In_916,In_902);
or U4454 (N_4454,In_717,In_441);
nand U4455 (N_4455,In_695,In_842);
or U4456 (N_4456,In_816,In_568);
nor U4457 (N_4457,In_627,In_602);
nand U4458 (N_4458,In_339,In_77);
or U4459 (N_4459,In_267,In_594);
or U4460 (N_4460,In_695,In_460);
nand U4461 (N_4461,In_44,In_289);
or U4462 (N_4462,In_59,In_596);
nor U4463 (N_4463,In_843,In_255);
or U4464 (N_4464,In_115,In_217);
and U4465 (N_4465,In_212,In_826);
nand U4466 (N_4466,In_471,In_89);
or U4467 (N_4467,In_135,In_125);
nand U4468 (N_4468,In_705,In_229);
or U4469 (N_4469,In_319,In_707);
and U4470 (N_4470,In_143,In_886);
nand U4471 (N_4471,In_647,In_718);
and U4472 (N_4472,In_399,In_787);
or U4473 (N_4473,In_419,In_176);
nor U4474 (N_4474,In_733,In_930);
nor U4475 (N_4475,In_587,In_618);
nand U4476 (N_4476,In_137,In_220);
xnor U4477 (N_4477,In_518,In_190);
nor U4478 (N_4478,In_414,In_252);
nand U4479 (N_4479,In_548,In_398);
and U4480 (N_4480,In_325,In_829);
nor U4481 (N_4481,In_212,In_835);
and U4482 (N_4482,In_428,In_799);
nand U4483 (N_4483,In_314,In_346);
or U4484 (N_4484,In_882,In_868);
nor U4485 (N_4485,In_757,In_213);
or U4486 (N_4486,In_801,In_637);
and U4487 (N_4487,In_496,In_92);
and U4488 (N_4488,In_408,In_834);
and U4489 (N_4489,In_844,In_113);
and U4490 (N_4490,In_94,In_810);
and U4491 (N_4491,In_215,In_882);
or U4492 (N_4492,In_715,In_842);
nand U4493 (N_4493,In_633,In_676);
nor U4494 (N_4494,In_754,In_69);
nor U4495 (N_4495,In_625,In_317);
nand U4496 (N_4496,In_912,In_419);
and U4497 (N_4497,In_134,In_65);
and U4498 (N_4498,In_119,In_572);
nor U4499 (N_4499,In_818,In_22);
nand U4500 (N_4500,In_367,In_671);
and U4501 (N_4501,In_907,In_970);
and U4502 (N_4502,In_196,In_943);
and U4503 (N_4503,In_316,In_132);
nand U4504 (N_4504,In_0,In_236);
nand U4505 (N_4505,In_364,In_365);
nor U4506 (N_4506,In_903,In_170);
nor U4507 (N_4507,In_531,In_684);
or U4508 (N_4508,In_838,In_734);
or U4509 (N_4509,In_909,In_103);
and U4510 (N_4510,In_304,In_544);
or U4511 (N_4511,In_24,In_143);
nand U4512 (N_4512,In_597,In_470);
nor U4513 (N_4513,In_852,In_520);
xor U4514 (N_4514,In_851,In_940);
or U4515 (N_4515,In_919,In_170);
and U4516 (N_4516,In_905,In_521);
nand U4517 (N_4517,In_153,In_581);
and U4518 (N_4518,In_913,In_469);
xor U4519 (N_4519,In_717,In_418);
or U4520 (N_4520,In_240,In_296);
and U4521 (N_4521,In_702,In_299);
or U4522 (N_4522,In_795,In_37);
or U4523 (N_4523,In_176,In_259);
nor U4524 (N_4524,In_143,In_950);
nand U4525 (N_4525,In_852,In_22);
and U4526 (N_4526,In_577,In_41);
nor U4527 (N_4527,In_15,In_195);
or U4528 (N_4528,In_682,In_562);
or U4529 (N_4529,In_789,In_423);
or U4530 (N_4530,In_115,In_800);
nand U4531 (N_4531,In_679,In_356);
xor U4532 (N_4532,In_555,In_188);
or U4533 (N_4533,In_752,In_168);
or U4534 (N_4534,In_347,In_68);
nand U4535 (N_4535,In_74,In_172);
xor U4536 (N_4536,In_467,In_965);
nor U4537 (N_4537,In_147,In_289);
nor U4538 (N_4538,In_40,In_910);
nand U4539 (N_4539,In_17,In_251);
and U4540 (N_4540,In_940,In_831);
nor U4541 (N_4541,In_543,In_570);
nand U4542 (N_4542,In_745,In_262);
and U4543 (N_4543,In_444,In_697);
and U4544 (N_4544,In_425,In_870);
or U4545 (N_4545,In_581,In_150);
or U4546 (N_4546,In_338,In_981);
xor U4547 (N_4547,In_436,In_785);
nor U4548 (N_4548,In_474,In_754);
nor U4549 (N_4549,In_416,In_244);
xnor U4550 (N_4550,In_664,In_48);
nand U4551 (N_4551,In_738,In_173);
or U4552 (N_4552,In_498,In_50);
or U4553 (N_4553,In_668,In_322);
or U4554 (N_4554,In_178,In_430);
nor U4555 (N_4555,In_562,In_224);
or U4556 (N_4556,In_562,In_545);
nor U4557 (N_4557,In_99,In_644);
nor U4558 (N_4558,In_994,In_654);
and U4559 (N_4559,In_599,In_226);
nor U4560 (N_4560,In_511,In_448);
or U4561 (N_4561,In_567,In_319);
and U4562 (N_4562,In_258,In_274);
xnor U4563 (N_4563,In_163,In_252);
and U4564 (N_4564,In_0,In_478);
and U4565 (N_4565,In_868,In_845);
and U4566 (N_4566,In_737,In_173);
and U4567 (N_4567,In_74,In_587);
nand U4568 (N_4568,In_384,In_257);
nor U4569 (N_4569,In_907,In_2);
or U4570 (N_4570,In_731,In_709);
nand U4571 (N_4571,In_245,In_149);
nor U4572 (N_4572,In_332,In_268);
and U4573 (N_4573,In_33,In_228);
nand U4574 (N_4574,In_828,In_893);
or U4575 (N_4575,In_709,In_131);
nand U4576 (N_4576,In_922,In_276);
nand U4577 (N_4577,In_56,In_195);
nand U4578 (N_4578,In_149,In_788);
and U4579 (N_4579,In_269,In_976);
nor U4580 (N_4580,In_116,In_52);
nand U4581 (N_4581,In_256,In_988);
nand U4582 (N_4582,In_701,In_127);
nand U4583 (N_4583,In_300,In_831);
or U4584 (N_4584,In_491,In_685);
or U4585 (N_4585,In_893,In_707);
and U4586 (N_4586,In_995,In_94);
xor U4587 (N_4587,In_449,In_441);
or U4588 (N_4588,In_289,In_264);
and U4589 (N_4589,In_988,In_270);
and U4590 (N_4590,In_289,In_546);
nand U4591 (N_4591,In_172,In_23);
and U4592 (N_4592,In_649,In_530);
nand U4593 (N_4593,In_323,In_183);
and U4594 (N_4594,In_897,In_53);
or U4595 (N_4595,In_148,In_834);
or U4596 (N_4596,In_677,In_18);
nor U4597 (N_4597,In_605,In_398);
nor U4598 (N_4598,In_727,In_332);
nand U4599 (N_4599,In_186,In_225);
and U4600 (N_4600,In_362,In_29);
nand U4601 (N_4601,In_921,In_125);
nor U4602 (N_4602,In_45,In_624);
or U4603 (N_4603,In_402,In_573);
and U4604 (N_4604,In_984,In_552);
nand U4605 (N_4605,In_754,In_512);
nor U4606 (N_4606,In_554,In_646);
xor U4607 (N_4607,In_688,In_994);
or U4608 (N_4608,In_135,In_494);
or U4609 (N_4609,In_76,In_192);
and U4610 (N_4610,In_617,In_573);
nor U4611 (N_4611,In_222,In_291);
nand U4612 (N_4612,In_233,In_660);
and U4613 (N_4613,In_290,In_501);
nand U4614 (N_4614,In_285,In_955);
nand U4615 (N_4615,In_69,In_740);
or U4616 (N_4616,In_399,In_284);
or U4617 (N_4617,In_620,In_84);
nand U4618 (N_4618,In_370,In_333);
nand U4619 (N_4619,In_247,In_552);
nor U4620 (N_4620,In_108,In_122);
nor U4621 (N_4621,In_782,In_184);
or U4622 (N_4622,In_333,In_740);
and U4623 (N_4623,In_249,In_718);
nor U4624 (N_4624,In_237,In_641);
or U4625 (N_4625,In_758,In_389);
nand U4626 (N_4626,In_662,In_526);
and U4627 (N_4627,In_427,In_896);
nand U4628 (N_4628,In_755,In_413);
nor U4629 (N_4629,In_565,In_780);
and U4630 (N_4630,In_658,In_880);
or U4631 (N_4631,In_969,In_937);
nor U4632 (N_4632,In_298,In_211);
and U4633 (N_4633,In_53,In_257);
and U4634 (N_4634,In_712,In_324);
nor U4635 (N_4635,In_398,In_865);
nand U4636 (N_4636,In_374,In_720);
nand U4637 (N_4637,In_997,In_485);
or U4638 (N_4638,In_107,In_777);
nor U4639 (N_4639,In_750,In_637);
xor U4640 (N_4640,In_188,In_295);
or U4641 (N_4641,In_403,In_812);
or U4642 (N_4642,In_944,In_508);
and U4643 (N_4643,In_272,In_544);
and U4644 (N_4644,In_845,In_885);
nor U4645 (N_4645,In_365,In_489);
nand U4646 (N_4646,In_758,In_655);
or U4647 (N_4647,In_129,In_958);
or U4648 (N_4648,In_354,In_298);
and U4649 (N_4649,In_993,In_475);
or U4650 (N_4650,In_74,In_162);
nand U4651 (N_4651,In_441,In_437);
and U4652 (N_4652,In_956,In_923);
nand U4653 (N_4653,In_144,In_168);
or U4654 (N_4654,In_955,In_455);
nor U4655 (N_4655,In_481,In_68);
nand U4656 (N_4656,In_381,In_444);
or U4657 (N_4657,In_407,In_937);
nor U4658 (N_4658,In_797,In_272);
or U4659 (N_4659,In_8,In_718);
or U4660 (N_4660,In_868,In_680);
nand U4661 (N_4661,In_113,In_940);
and U4662 (N_4662,In_397,In_405);
and U4663 (N_4663,In_290,In_856);
xnor U4664 (N_4664,In_229,In_718);
nor U4665 (N_4665,In_949,In_979);
and U4666 (N_4666,In_100,In_506);
and U4667 (N_4667,In_565,In_733);
and U4668 (N_4668,In_453,In_741);
and U4669 (N_4669,In_542,In_432);
and U4670 (N_4670,In_862,In_985);
and U4671 (N_4671,In_415,In_632);
or U4672 (N_4672,In_667,In_55);
nor U4673 (N_4673,In_59,In_980);
nand U4674 (N_4674,In_827,In_54);
xor U4675 (N_4675,In_649,In_711);
or U4676 (N_4676,In_460,In_111);
or U4677 (N_4677,In_824,In_618);
nor U4678 (N_4678,In_511,In_380);
nand U4679 (N_4679,In_539,In_30);
nor U4680 (N_4680,In_604,In_12);
nand U4681 (N_4681,In_456,In_290);
nand U4682 (N_4682,In_923,In_340);
and U4683 (N_4683,In_160,In_935);
nor U4684 (N_4684,In_865,In_380);
nor U4685 (N_4685,In_157,In_708);
and U4686 (N_4686,In_125,In_14);
or U4687 (N_4687,In_247,In_216);
nor U4688 (N_4688,In_699,In_950);
and U4689 (N_4689,In_141,In_471);
nor U4690 (N_4690,In_154,In_326);
nor U4691 (N_4691,In_501,In_713);
nand U4692 (N_4692,In_867,In_758);
nor U4693 (N_4693,In_820,In_819);
nor U4694 (N_4694,In_643,In_27);
nor U4695 (N_4695,In_348,In_530);
nor U4696 (N_4696,In_915,In_3);
nor U4697 (N_4697,In_96,In_121);
nand U4698 (N_4698,In_675,In_692);
nand U4699 (N_4699,In_600,In_533);
xnor U4700 (N_4700,In_825,In_357);
nand U4701 (N_4701,In_391,In_696);
and U4702 (N_4702,In_814,In_908);
or U4703 (N_4703,In_290,In_932);
nor U4704 (N_4704,In_841,In_587);
nand U4705 (N_4705,In_853,In_319);
nand U4706 (N_4706,In_543,In_117);
xnor U4707 (N_4707,In_942,In_72);
and U4708 (N_4708,In_665,In_314);
nand U4709 (N_4709,In_363,In_278);
xnor U4710 (N_4710,In_44,In_156);
and U4711 (N_4711,In_39,In_573);
or U4712 (N_4712,In_781,In_348);
nand U4713 (N_4713,In_493,In_432);
nand U4714 (N_4714,In_272,In_427);
xor U4715 (N_4715,In_15,In_404);
or U4716 (N_4716,In_321,In_374);
nand U4717 (N_4717,In_665,In_308);
nand U4718 (N_4718,In_724,In_236);
or U4719 (N_4719,In_258,In_577);
or U4720 (N_4720,In_472,In_795);
and U4721 (N_4721,In_565,In_919);
nor U4722 (N_4722,In_234,In_213);
or U4723 (N_4723,In_756,In_160);
nor U4724 (N_4724,In_303,In_820);
xor U4725 (N_4725,In_169,In_187);
and U4726 (N_4726,In_849,In_217);
and U4727 (N_4727,In_765,In_832);
or U4728 (N_4728,In_43,In_353);
nor U4729 (N_4729,In_29,In_370);
nand U4730 (N_4730,In_36,In_258);
nand U4731 (N_4731,In_918,In_735);
nor U4732 (N_4732,In_770,In_929);
or U4733 (N_4733,In_77,In_774);
or U4734 (N_4734,In_54,In_142);
xor U4735 (N_4735,In_463,In_232);
or U4736 (N_4736,In_211,In_917);
nand U4737 (N_4737,In_846,In_562);
or U4738 (N_4738,In_597,In_663);
nor U4739 (N_4739,In_8,In_440);
nand U4740 (N_4740,In_743,In_863);
nor U4741 (N_4741,In_810,In_61);
and U4742 (N_4742,In_366,In_350);
or U4743 (N_4743,In_409,In_830);
nand U4744 (N_4744,In_403,In_941);
or U4745 (N_4745,In_931,In_474);
and U4746 (N_4746,In_404,In_855);
xor U4747 (N_4747,In_794,In_288);
and U4748 (N_4748,In_229,In_148);
nor U4749 (N_4749,In_429,In_678);
or U4750 (N_4750,In_95,In_178);
nand U4751 (N_4751,In_689,In_998);
nand U4752 (N_4752,In_288,In_625);
or U4753 (N_4753,In_329,In_886);
or U4754 (N_4754,In_992,In_213);
nor U4755 (N_4755,In_154,In_49);
nor U4756 (N_4756,In_122,In_747);
and U4757 (N_4757,In_338,In_141);
nand U4758 (N_4758,In_757,In_628);
nand U4759 (N_4759,In_126,In_658);
and U4760 (N_4760,In_800,In_958);
and U4761 (N_4761,In_752,In_782);
or U4762 (N_4762,In_888,In_179);
nand U4763 (N_4763,In_917,In_679);
nor U4764 (N_4764,In_154,In_417);
xnor U4765 (N_4765,In_756,In_616);
nor U4766 (N_4766,In_960,In_242);
or U4767 (N_4767,In_593,In_947);
nand U4768 (N_4768,In_58,In_872);
nand U4769 (N_4769,In_968,In_564);
nand U4770 (N_4770,In_517,In_12);
and U4771 (N_4771,In_625,In_650);
nor U4772 (N_4772,In_883,In_536);
nor U4773 (N_4773,In_408,In_750);
and U4774 (N_4774,In_552,In_619);
and U4775 (N_4775,In_875,In_109);
and U4776 (N_4776,In_281,In_178);
or U4777 (N_4777,In_712,In_137);
nand U4778 (N_4778,In_457,In_403);
nand U4779 (N_4779,In_285,In_600);
and U4780 (N_4780,In_923,In_907);
nor U4781 (N_4781,In_633,In_252);
nor U4782 (N_4782,In_186,In_978);
nor U4783 (N_4783,In_744,In_999);
and U4784 (N_4784,In_17,In_262);
and U4785 (N_4785,In_742,In_841);
and U4786 (N_4786,In_698,In_937);
or U4787 (N_4787,In_312,In_71);
and U4788 (N_4788,In_234,In_463);
nand U4789 (N_4789,In_750,In_956);
nor U4790 (N_4790,In_803,In_934);
nor U4791 (N_4791,In_131,In_769);
and U4792 (N_4792,In_582,In_198);
and U4793 (N_4793,In_512,In_618);
nand U4794 (N_4794,In_917,In_189);
xor U4795 (N_4795,In_842,In_457);
nand U4796 (N_4796,In_894,In_795);
or U4797 (N_4797,In_578,In_58);
and U4798 (N_4798,In_922,In_428);
nand U4799 (N_4799,In_652,In_533);
or U4800 (N_4800,In_274,In_889);
or U4801 (N_4801,In_739,In_751);
or U4802 (N_4802,In_203,In_612);
nor U4803 (N_4803,In_793,In_894);
and U4804 (N_4804,In_343,In_610);
or U4805 (N_4805,In_47,In_164);
or U4806 (N_4806,In_898,In_63);
nor U4807 (N_4807,In_110,In_338);
nor U4808 (N_4808,In_540,In_251);
nor U4809 (N_4809,In_471,In_99);
or U4810 (N_4810,In_780,In_574);
or U4811 (N_4811,In_273,In_354);
nand U4812 (N_4812,In_885,In_288);
and U4813 (N_4813,In_694,In_629);
and U4814 (N_4814,In_222,In_835);
nand U4815 (N_4815,In_369,In_8);
nor U4816 (N_4816,In_338,In_347);
xnor U4817 (N_4817,In_740,In_177);
or U4818 (N_4818,In_225,In_527);
and U4819 (N_4819,In_931,In_598);
or U4820 (N_4820,In_984,In_66);
nor U4821 (N_4821,In_547,In_778);
nand U4822 (N_4822,In_843,In_452);
and U4823 (N_4823,In_288,In_681);
or U4824 (N_4824,In_355,In_952);
or U4825 (N_4825,In_499,In_287);
and U4826 (N_4826,In_980,In_61);
or U4827 (N_4827,In_866,In_878);
and U4828 (N_4828,In_210,In_454);
nor U4829 (N_4829,In_600,In_613);
or U4830 (N_4830,In_84,In_198);
nor U4831 (N_4831,In_218,In_354);
nor U4832 (N_4832,In_931,In_36);
nand U4833 (N_4833,In_528,In_708);
nor U4834 (N_4834,In_754,In_163);
and U4835 (N_4835,In_374,In_748);
or U4836 (N_4836,In_633,In_617);
and U4837 (N_4837,In_941,In_496);
and U4838 (N_4838,In_375,In_712);
or U4839 (N_4839,In_816,In_569);
nor U4840 (N_4840,In_84,In_996);
and U4841 (N_4841,In_19,In_459);
nand U4842 (N_4842,In_345,In_193);
nor U4843 (N_4843,In_256,In_7);
and U4844 (N_4844,In_635,In_329);
and U4845 (N_4845,In_120,In_583);
and U4846 (N_4846,In_284,In_203);
nor U4847 (N_4847,In_968,In_530);
nor U4848 (N_4848,In_333,In_92);
nand U4849 (N_4849,In_649,In_80);
and U4850 (N_4850,In_456,In_34);
nor U4851 (N_4851,In_998,In_517);
nand U4852 (N_4852,In_736,In_524);
and U4853 (N_4853,In_815,In_586);
and U4854 (N_4854,In_56,In_985);
nand U4855 (N_4855,In_485,In_353);
nand U4856 (N_4856,In_978,In_205);
nand U4857 (N_4857,In_500,In_954);
nor U4858 (N_4858,In_417,In_141);
nand U4859 (N_4859,In_966,In_762);
or U4860 (N_4860,In_404,In_969);
or U4861 (N_4861,In_714,In_466);
nor U4862 (N_4862,In_762,In_132);
nor U4863 (N_4863,In_849,In_989);
nand U4864 (N_4864,In_310,In_865);
or U4865 (N_4865,In_560,In_501);
nor U4866 (N_4866,In_400,In_888);
and U4867 (N_4867,In_332,In_756);
nor U4868 (N_4868,In_444,In_101);
and U4869 (N_4869,In_254,In_54);
and U4870 (N_4870,In_219,In_26);
or U4871 (N_4871,In_599,In_776);
and U4872 (N_4872,In_153,In_99);
nor U4873 (N_4873,In_330,In_235);
and U4874 (N_4874,In_104,In_829);
nor U4875 (N_4875,In_896,In_485);
or U4876 (N_4876,In_527,In_967);
and U4877 (N_4877,In_664,In_26);
nor U4878 (N_4878,In_25,In_872);
and U4879 (N_4879,In_865,In_92);
or U4880 (N_4880,In_363,In_507);
and U4881 (N_4881,In_564,In_216);
nand U4882 (N_4882,In_569,In_525);
or U4883 (N_4883,In_440,In_100);
and U4884 (N_4884,In_434,In_813);
or U4885 (N_4885,In_919,In_676);
nor U4886 (N_4886,In_276,In_263);
or U4887 (N_4887,In_848,In_747);
and U4888 (N_4888,In_575,In_804);
or U4889 (N_4889,In_479,In_523);
nand U4890 (N_4890,In_977,In_670);
nor U4891 (N_4891,In_490,In_790);
nand U4892 (N_4892,In_174,In_526);
nor U4893 (N_4893,In_410,In_476);
nor U4894 (N_4894,In_988,In_344);
nand U4895 (N_4895,In_332,In_633);
nand U4896 (N_4896,In_257,In_794);
and U4897 (N_4897,In_856,In_937);
nor U4898 (N_4898,In_953,In_698);
nand U4899 (N_4899,In_863,In_974);
or U4900 (N_4900,In_755,In_544);
nor U4901 (N_4901,In_556,In_609);
xor U4902 (N_4902,In_742,In_105);
nand U4903 (N_4903,In_977,In_189);
or U4904 (N_4904,In_576,In_248);
nand U4905 (N_4905,In_395,In_162);
and U4906 (N_4906,In_547,In_985);
nor U4907 (N_4907,In_411,In_515);
nor U4908 (N_4908,In_320,In_224);
nand U4909 (N_4909,In_293,In_283);
or U4910 (N_4910,In_200,In_270);
nor U4911 (N_4911,In_833,In_79);
and U4912 (N_4912,In_287,In_748);
or U4913 (N_4913,In_719,In_264);
or U4914 (N_4914,In_732,In_951);
nand U4915 (N_4915,In_20,In_362);
nand U4916 (N_4916,In_678,In_513);
nor U4917 (N_4917,In_604,In_829);
nor U4918 (N_4918,In_26,In_199);
or U4919 (N_4919,In_647,In_433);
xor U4920 (N_4920,In_759,In_278);
or U4921 (N_4921,In_783,In_308);
nor U4922 (N_4922,In_49,In_846);
nor U4923 (N_4923,In_607,In_9);
and U4924 (N_4924,In_462,In_407);
xnor U4925 (N_4925,In_225,In_873);
nand U4926 (N_4926,In_55,In_716);
and U4927 (N_4927,In_908,In_789);
nand U4928 (N_4928,In_648,In_679);
and U4929 (N_4929,In_928,In_447);
or U4930 (N_4930,In_703,In_673);
nand U4931 (N_4931,In_533,In_590);
or U4932 (N_4932,In_804,In_715);
nor U4933 (N_4933,In_650,In_69);
or U4934 (N_4934,In_678,In_14);
and U4935 (N_4935,In_698,In_115);
nand U4936 (N_4936,In_59,In_873);
and U4937 (N_4937,In_645,In_222);
nor U4938 (N_4938,In_338,In_119);
nand U4939 (N_4939,In_502,In_370);
and U4940 (N_4940,In_612,In_180);
nor U4941 (N_4941,In_392,In_628);
nor U4942 (N_4942,In_340,In_201);
or U4943 (N_4943,In_114,In_646);
and U4944 (N_4944,In_309,In_392);
nor U4945 (N_4945,In_299,In_723);
nor U4946 (N_4946,In_669,In_881);
and U4947 (N_4947,In_749,In_734);
nor U4948 (N_4948,In_55,In_861);
or U4949 (N_4949,In_623,In_669);
or U4950 (N_4950,In_612,In_940);
or U4951 (N_4951,In_64,In_728);
or U4952 (N_4952,In_7,In_210);
nand U4953 (N_4953,In_24,In_723);
xor U4954 (N_4954,In_199,In_698);
nor U4955 (N_4955,In_136,In_807);
nand U4956 (N_4956,In_782,In_703);
nor U4957 (N_4957,In_221,In_200);
nor U4958 (N_4958,In_281,In_125);
nor U4959 (N_4959,In_161,In_293);
nand U4960 (N_4960,In_335,In_758);
and U4961 (N_4961,In_818,In_130);
or U4962 (N_4962,In_824,In_354);
nor U4963 (N_4963,In_472,In_735);
or U4964 (N_4964,In_955,In_699);
nand U4965 (N_4965,In_571,In_975);
or U4966 (N_4966,In_781,In_336);
xnor U4967 (N_4967,In_943,In_662);
nor U4968 (N_4968,In_916,In_79);
nand U4969 (N_4969,In_930,In_225);
nand U4970 (N_4970,In_869,In_18);
and U4971 (N_4971,In_300,In_209);
nor U4972 (N_4972,In_366,In_195);
nand U4973 (N_4973,In_832,In_503);
or U4974 (N_4974,In_140,In_983);
nor U4975 (N_4975,In_244,In_268);
nand U4976 (N_4976,In_847,In_797);
nand U4977 (N_4977,In_334,In_322);
or U4978 (N_4978,In_132,In_418);
or U4979 (N_4979,In_428,In_750);
and U4980 (N_4980,In_643,In_154);
or U4981 (N_4981,In_244,In_209);
nor U4982 (N_4982,In_835,In_308);
nand U4983 (N_4983,In_588,In_709);
xor U4984 (N_4984,In_174,In_844);
nand U4985 (N_4985,In_755,In_534);
nand U4986 (N_4986,In_138,In_714);
or U4987 (N_4987,In_30,In_944);
and U4988 (N_4988,In_624,In_761);
and U4989 (N_4989,In_339,In_49);
or U4990 (N_4990,In_574,In_60);
nand U4991 (N_4991,In_177,In_77);
nor U4992 (N_4992,In_194,In_304);
and U4993 (N_4993,In_838,In_640);
nand U4994 (N_4994,In_520,In_995);
or U4995 (N_4995,In_514,In_495);
nand U4996 (N_4996,In_910,In_336);
nand U4997 (N_4997,In_201,In_42);
or U4998 (N_4998,In_93,In_705);
and U4999 (N_4999,In_788,In_476);
nand U5000 (N_5000,N_3868,N_4909);
nand U5001 (N_5001,N_2165,N_2916);
and U5002 (N_5002,N_243,N_3082);
nor U5003 (N_5003,N_2374,N_2655);
or U5004 (N_5004,N_1749,N_1784);
and U5005 (N_5005,N_105,N_294);
and U5006 (N_5006,N_4361,N_1551);
nor U5007 (N_5007,N_4512,N_3555);
nand U5008 (N_5008,N_454,N_4059);
or U5009 (N_5009,N_3591,N_1108);
nor U5010 (N_5010,N_3375,N_3959);
nand U5011 (N_5011,N_2336,N_1729);
or U5012 (N_5012,N_1812,N_4408);
nor U5013 (N_5013,N_3283,N_3987);
nand U5014 (N_5014,N_415,N_277);
nor U5015 (N_5015,N_4127,N_3753);
and U5016 (N_5016,N_309,N_2547);
nor U5017 (N_5017,N_3739,N_3636);
nor U5018 (N_5018,N_3382,N_3589);
and U5019 (N_5019,N_3991,N_1403);
nor U5020 (N_5020,N_4885,N_1752);
xnor U5021 (N_5021,N_318,N_112);
and U5022 (N_5022,N_4939,N_972);
and U5023 (N_5023,N_4578,N_4207);
or U5024 (N_5024,N_1430,N_409);
xnor U5025 (N_5025,N_3440,N_3666);
and U5026 (N_5026,N_1191,N_2856);
nor U5027 (N_5027,N_2543,N_3139);
nor U5028 (N_5028,N_4052,N_4312);
nand U5029 (N_5029,N_1653,N_3757);
nor U5030 (N_5030,N_1634,N_2662);
and U5031 (N_5031,N_2199,N_1346);
nor U5032 (N_5032,N_4302,N_537);
nand U5033 (N_5033,N_2465,N_3136);
nand U5034 (N_5034,N_2051,N_4595);
nand U5035 (N_5035,N_130,N_1562);
and U5036 (N_5036,N_2839,N_2701);
or U5037 (N_5037,N_4426,N_2891);
and U5038 (N_5038,N_1724,N_297);
nor U5039 (N_5039,N_4145,N_43);
and U5040 (N_5040,N_2949,N_4739);
or U5041 (N_5041,N_1094,N_3367);
nand U5042 (N_5042,N_4093,N_3779);
nor U5043 (N_5043,N_2933,N_374);
and U5044 (N_5044,N_4161,N_1319);
xnor U5045 (N_5045,N_4109,N_4536);
or U5046 (N_5046,N_3904,N_3063);
nor U5047 (N_5047,N_1861,N_4611);
and U5048 (N_5048,N_2578,N_4508);
and U5049 (N_5049,N_1185,N_786);
and U5050 (N_5050,N_2231,N_4676);
and U5051 (N_5051,N_1605,N_1090);
and U5052 (N_5052,N_1523,N_3008);
or U5053 (N_5053,N_3651,N_2031);
nand U5054 (N_5054,N_1371,N_522);
nand U5055 (N_5055,N_4637,N_2544);
nand U5056 (N_5056,N_4754,N_102);
nand U5057 (N_5057,N_2260,N_2598);
and U5058 (N_5058,N_4405,N_4363);
nand U5059 (N_5059,N_4397,N_1950);
nor U5060 (N_5060,N_390,N_548);
nand U5061 (N_5061,N_1601,N_2132);
and U5062 (N_5062,N_3869,N_1199);
nor U5063 (N_5063,N_4131,N_4884);
nor U5064 (N_5064,N_2119,N_1258);
and U5065 (N_5065,N_4496,N_2833);
or U5066 (N_5066,N_3160,N_3342);
and U5067 (N_5067,N_191,N_4530);
or U5068 (N_5068,N_72,N_540);
and U5069 (N_5069,N_1461,N_97);
nor U5070 (N_5070,N_312,N_4745);
nand U5071 (N_5071,N_2163,N_3125);
and U5072 (N_5072,N_2185,N_2315);
and U5073 (N_5073,N_950,N_4857);
and U5074 (N_5074,N_2085,N_1168);
or U5075 (N_5075,N_2718,N_3054);
nand U5076 (N_5076,N_917,N_4417);
and U5077 (N_5077,N_3781,N_84);
nor U5078 (N_5078,N_1277,N_1619);
or U5079 (N_5079,N_559,N_4951);
or U5080 (N_5080,N_891,N_2780);
nor U5081 (N_5081,N_3413,N_3265);
or U5082 (N_5082,N_209,N_2563);
and U5083 (N_5083,N_2939,N_2018);
and U5084 (N_5084,N_1487,N_2675);
nand U5085 (N_5085,N_3627,N_2134);
nor U5086 (N_5086,N_4101,N_2133);
nand U5087 (N_5087,N_800,N_4490);
or U5088 (N_5088,N_4241,N_539);
or U5089 (N_5089,N_500,N_2641);
and U5090 (N_5090,N_1607,N_2552);
or U5091 (N_5091,N_4500,N_2836);
nand U5092 (N_5092,N_1955,N_1522);
and U5093 (N_5093,N_2243,N_3643);
nand U5094 (N_5094,N_2028,N_1069);
nor U5095 (N_5095,N_2511,N_480);
nand U5096 (N_5096,N_2184,N_1170);
xnor U5097 (N_5097,N_2900,N_2265);
or U5098 (N_5098,N_207,N_2424);
nor U5099 (N_5099,N_1034,N_3941);
or U5100 (N_5100,N_2913,N_427);
nor U5101 (N_5101,N_2129,N_4625);
and U5102 (N_5102,N_2645,N_247);
and U5103 (N_5103,N_613,N_2301);
nand U5104 (N_5104,N_2379,N_4516);
nand U5105 (N_5105,N_941,N_1010);
nor U5106 (N_5106,N_4874,N_2510);
nor U5107 (N_5107,N_4802,N_4376);
nor U5108 (N_5108,N_4971,N_2468);
and U5109 (N_5109,N_2521,N_1545);
nand U5110 (N_5110,N_3046,N_3242);
and U5111 (N_5111,N_1716,N_298);
or U5112 (N_5112,N_3354,N_25);
nor U5113 (N_5113,N_2647,N_4088);
nand U5114 (N_5114,N_3765,N_4114);
or U5115 (N_5115,N_3864,N_2015);
and U5116 (N_5116,N_1374,N_1356);
nand U5117 (N_5117,N_3123,N_245);
nand U5118 (N_5118,N_4137,N_4091);
nor U5119 (N_5119,N_3386,N_1706);
nor U5120 (N_5120,N_2053,N_3185);
nor U5121 (N_5121,N_980,N_4049);
nor U5122 (N_5122,N_395,N_2588);
nor U5123 (N_5123,N_2887,N_3993);
nand U5124 (N_5124,N_4463,N_1883);
nand U5125 (N_5125,N_3142,N_3190);
nor U5126 (N_5126,N_3023,N_4314);
nand U5127 (N_5127,N_372,N_2760);
and U5128 (N_5128,N_4236,N_3405);
or U5129 (N_5129,N_4650,N_4069);
nand U5130 (N_5130,N_1934,N_4348);
or U5131 (N_5131,N_3919,N_3790);
nand U5132 (N_5132,N_1966,N_2125);
nor U5133 (N_5133,N_568,N_1288);
nand U5134 (N_5134,N_3061,N_734);
nand U5135 (N_5135,N_1492,N_4605);
nor U5136 (N_5136,N_3542,N_3866);
or U5137 (N_5137,N_2773,N_4094);
nor U5138 (N_5138,N_3490,N_2771);
nor U5139 (N_5139,N_2843,N_4660);
nor U5140 (N_5140,N_216,N_3925);
nand U5141 (N_5141,N_724,N_3645);
or U5142 (N_5142,N_1206,N_2342);
or U5143 (N_5143,N_255,N_1328);
and U5144 (N_5144,N_4471,N_3122);
or U5145 (N_5145,N_2932,N_1313);
and U5146 (N_5146,N_706,N_3568);
nor U5147 (N_5147,N_4203,N_771);
or U5148 (N_5148,N_4324,N_4535);
or U5149 (N_5149,N_3252,N_4195);
nand U5150 (N_5150,N_2976,N_1312);
nand U5151 (N_5151,N_1783,N_1173);
and U5152 (N_5152,N_3224,N_3742);
nand U5153 (N_5153,N_2435,N_4225);
and U5154 (N_5154,N_1622,N_1662);
nand U5155 (N_5155,N_4529,N_1334);
nand U5156 (N_5156,N_2012,N_4820);
nand U5157 (N_5157,N_2448,N_711);
or U5158 (N_5158,N_1681,N_171);
or U5159 (N_5159,N_1774,N_4062);
or U5160 (N_5160,N_3554,N_1731);
and U5161 (N_5161,N_2264,N_3289);
or U5162 (N_5162,N_1887,N_4954);
nand U5163 (N_5163,N_3510,N_3079);
nand U5164 (N_5164,N_4035,N_3258);
nand U5165 (N_5165,N_1058,N_3797);
or U5166 (N_5166,N_3321,N_3646);
and U5167 (N_5167,N_1370,N_2661);
nor U5168 (N_5168,N_4394,N_3557);
and U5169 (N_5169,N_2558,N_1448);
nor U5170 (N_5170,N_3710,N_3691);
and U5171 (N_5171,N_1047,N_3196);
or U5172 (N_5172,N_574,N_2206);
nand U5173 (N_5173,N_4333,N_2036);
nor U5174 (N_5174,N_2633,N_3768);
nand U5175 (N_5175,N_3719,N_546);
nor U5176 (N_5176,N_3389,N_2364);
or U5177 (N_5177,N_4944,N_710);
nor U5178 (N_5178,N_2101,N_2312);
nor U5179 (N_5179,N_1560,N_1903);
nand U5180 (N_5180,N_2546,N_4429);
nand U5181 (N_5181,N_976,N_2501);
and U5182 (N_5182,N_2621,N_1439);
or U5183 (N_5183,N_2237,N_3736);
or U5184 (N_5184,N_2077,N_39);
nor U5185 (N_5185,N_2288,N_2951);
nand U5186 (N_5186,N_4711,N_819);
nor U5187 (N_5187,N_2726,N_554);
nor U5188 (N_5188,N_4838,N_4890);
or U5189 (N_5189,N_2162,N_2369);
nor U5190 (N_5190,N_68,N_4663);
nor U5191 (N_5191,N_4355,N_2750);
xnor U5192 (N_5192,N_3102,N_3671);
or U5193 (N_5193,N_3482,N_2466);
and U5194 (N_5194,N_1152,N_175);
nor U5195 (N_5195,N_2948,N_361);
and U5196 (N_5196,N_3276,N_571);
and U5197 (N_5197,N_2355,N_4881);
and U5198 (N_5198,N_618,N_1411);
or U5199 (N_5199,N_2504,N_1621);
nand U5200 (N_5200,N_2135,N_4449);
and U5201 (N_5201,N_3932,N_2110);
nand U5202 (N_5202,N_4823,N_4958);
nand U5203 (N_5203,N_3502,N_1916);
xor U5204 (N_5204,N_110,N_2961);
or U5205 (N_5205,N_3347,N_12);
and U5206 (N_5206,N_3293,N_4855);
nand U5207 (N_5207,N_2581,N_2236);
or U5208 (N_5208,N_11,N_73);
or U5209 (N_5209,N_1514,N_2892);
nor U5210 (N_5210,N_1423,N_2888);
and U5211 (N_5211,N_3170,N_639);
and U5212 (N_5212,N_4260,N_2094);
xnor U5213 (N_5213,N_3526,N_4713);
and U5214 (N_5214,N_4840,N_4180);
xnor U5215 (N_5215,N_1329,N_3240);
or U5216 (N_5216,N_3501,N_864);
nor U5217 (N_5217,N_1825,N_4528);
or U5218 (N_5218,N_1184,N_179);
and U5219 (N_5219,N_2562,N_4515);
nor U5220 (N_5220,N_2982,N_1945);
or U5221 (N_5221,N_760,N_4072);
nor U5222 (N_5222,N_4896,N_4372);
or U5223 (N_5223,N_2895,N_1115);
and U5224 (N_5224,N_3100,N_2140);
or U5225 (N_5225,N_2953,N_1464);
or U5226 (N_5226,N_3949,N_4119);
nor U5227 (N_5227,N_4387,N_2014);
nand U5228 (N_5228,N_1787,N_3496);
or U5229 (N_5229,N_2361,N_3667);
nor U5230 (N_5230,N_2883,N_4278);
and U5231 (N_5231,N_3107,N_24);
or U5232 (N_5232,N_2318,N_4416);
nor U5233 (N_5233,N_491,N_4570);
and U5234 (N_5234,N_473,N_3493);
and U5235 (N_5235,N_1111,N_2160);
and U5236 (N_5236,N_2564,N_4189);
nand U5237 (N_5237,N_1958,N_4111);
nor U5238 (N_5238,N_2327,N_2984);
nor U5239 (N_5239,N_3295,N_3514);
nor U5240 (N_5240,N_1056,N_350);
nand U5241 (N_5241,N_1134,N_4919);
nor U5242 (N_5242,N_4340,N_4075);
nor U5243 (N_5243,N_853,N_2256);
nand U5244 (N_5244,N_3882,N_2849);
nor U5245 (N_5245,N_2934,N_2003);
nand U5246 (N_5246,N_2207,N_3137);
nor U5247 (N_5247,N_748,N_1208);
or U5248 (N_5248,N_4994,N_236);
nand U5249 (N_5249,N_1211,N_1466);
nand U5250 (N_5250,N_2181,N_2560);
nand U5251 (N_5251,N_1956,N_4977);
nor U5252 (N_5252,N_3734,N_2349);
nand U5253 (N_5253,N_825,N_4157);
or U5254 (N_5254,N_1766,N_2317);
nand U5255 (N_5255,N_2149,N_60);
or U5256 (N_5256,N_3519,N_4803);
and U5257 (N_5257,N_757,N_2057);
nor U5258 (N_5258,N_871,N_4753);
and U5259 (N_5259,N_3393,N_966);
nand U5260 (N_5260,N_1529,N_4374);
xnor U5261 (N_5261,N_489,N_2357);
or U5262 (N_5262,N_1198,N_1557);
nor U5263 (N_5263,N_3085,N_1420);
and U5264 (N_5264,N_4606,N_4327);
nor U5265 (N_5265,N_693,N_1459);
or U5266 (N_5266,N_1264,N_3730);
or U5267 (N_5267,N_2286,N_1882);
and U5268 (N_5268,N_1011,N_3194);
nor U5269 (N_5269,N_1652,N_2746);
and U5270 (N_5270,N_4021,N_3371);
nor U5271 (N_5271,N_866,N_3004);
or U5272 (N_5272,N_1092,N_4593);
or U5273 (N_5273,N_1556,N_1892);
nand U5274 (N_5274,N_1162,N_2532);
and U5275 (N_5275,N_2820,N_2765);
and U5276 (N_5276,N_3447,N_2409);
nor U5277 (N_5277,N_1996,N_4704);
nand U5278 (N_5278,N_2296,N_364);
and U5279 (N_5279,N_387,N_3305);
or U5280 (N_5280,N_1990,N_1895);
or U5281 (N_5281,N_1323,N_1614);
nor U5282 (N_5282,N_708,N_3217);
nor U5283 (N_5283,N_1359,N_1878);
and U5284 (N_5284,N_765,N_217);
or U5285 (N_5285,N_342,N_2295);
nand U5286 (N_5286,N_3893,N_3564);
or U5287 (N_5287,N_584,N_2824);
nand U5288 (N_5288,N_2047,N_3307);
nor U5289 (N_5289,N_3433,N_1665);
xnor U5290 (N_5290,N_4023,N_2489);
nor U5291 (N_5291,N_2004,N_1383);
and U5292 (N_5292,N_1482,N_2289);
or U5293 (N_5293,N_98,N_4828);
nand U5294 (N_5294,N_4583,N_2550);
nand U5295 (N_5295,N_2007,N_4297);
nor U5296 (N_5296,N_2962,N_2522);
and U5297 (N_5297,N_3927,N_4859);
nand U5298 (N_5298,N_3895,N_3678);
nand U5299 (N_5299,N_3598,N_2396);
nand U5300 (N_5300,N_1151,N_3425);
and U5301 (N_5301,N_3124,N_4889);
or U5302 (N_5302,N_4081,N_4796);
nand U5303 (N_5303,N_335,N_3620);
and U5304 (N_5304,N_4003,N_3674);
nor U5305 (N_5305,N_1564,N_3962);
and U5306 (N_5306,N_1532,N_1525);
nand U5307 (N_5307,N_647,N_4947);
or U5308 (N_5308,N_1847,N_1046);
nand U5309 (N_5309,N_4614,N_4725);
nor U5310 (N_5310,N_4158,N_2920);
nor U5311 (N_5311,N_923,N_2131);
nand U5312 (N_5312,N_3346,N_2845);
nand U5313 (N_5313,N_2965,N_4549);
and U5314 (N_5314,N_661,N_2091);
xor U5315 (N_5315,N_10,N_3251);
or U5316 (N_5316,N_3648,N_1119);
or U5317 (N_5317,N_2612,N_1072);
or U5318 (N_5318,N_4102,N_2107);
nor U5319 (N_5319,N_1477,N_1538);
and U5320 (N_5320,N_3944,N_4474);
nand U5321 (N_5321,N_4247,N_9);
or U5322 (N_5322,N_2749,N_723);
and U5323 (N_5323,N_3318,N_482);
nor U5324 (N_5324,N_4099,N_435);
nand U5325 (N_5325,N_2535,N_1876);
nor U5326 (N_5326,N_4569,N_1458);
nand U5327 (N_5327,N_1123,N_1381);
and U5328 (N_5328,N_4092,N_674);
nor U5329 (N_5329,N_3961,N_2247);
or U5330 (N_5330,N_3458,N_1097);
nand U5331 (N_5331,N_1991,N_2690);
and U5332 (N_5332,N_4651,N_4707);
or U5333 (N_5333,N_1326,N_3036);
nand U5334 (N_5334,N_3049,N_2627);
nand U5335 (N_5335,N_3844,N_1480);
and U5336 (N_5336,N_636,N_963);
and U5337 (N_5337,N_3958,N_2067);
or U5338 (N_5338,N_4862,N_2724);
nor U5339 (N_5339,N_4329,N_1303);
nor U5340 (N_5340,N_1138,N_4983);
nand U5341 (N_5341,N_987,N_2373);
or U5342 (N_5342,N_580,N_2438);
xor U5343 (N_5343,N_3284,N_964);
and U5344 (N_5344,N_1169,N_1979);
nand U5345 (N_5345,N_2899,N_4544);
and U5346 (N_5346,N_1165,N_1321);
or U5347 (N_5347,N_3848,N_2141);
or U5348 (N_5348,N_3909,N_1164);
nand U5349 (N_5349,N_3398,N_1540);
nand U5350 (N_5350,N_295,N_3560);
or U5351 (N_5351,N_549,N_1535);
or U5352 (N_5352,N_2879,N_1009);
and U5353 (N_5353,N_1949,N_1566);
nand U5354 (N_5354,N_3,N_663);
and U5355 (N_5355,N_3520,N_2828);
or U5356 (N_5356,N_1068,N_2798);
nand U5357 (N_5357,N_839,N_4342);
or U5358 (N_5358,N_4357,N_4585);
or U5359 (N_5359,N_363,N_339);
or U5360 (N_5360,N_6,N_4431);
nand U5361 (N_5361,N_3806,N_4171);
or U5362 (N_5362,N_2486,N_2197);
or U5363 (N_5363,N_481,N_893);
and U5364 (N_5364,N_1554,N_1145);
xor U5365 (N_5365,N_4044,N_2853);
and U5366 (N_5366,N_1579,N_4852);
nand U5367 (N_5367,N_2224,N_31);
and U5368 (N_5368,N_125,N_2164);
nor U5369 (N_5369,N_205,N_3450);
nand U5370 (N_5370,N_4304,N_1526);
nand U5371 (N_5371,N_4851,N_1516);
and U5372 (N_5372,N_2994,N_4048);
nor U5373 (N_5373,N_1132,N_263);
nand U5374 (N_5374,N_2383,N_3906);
nor U5375 (N_5375,N_4441,N_2559);
and U5376 (N_5376,N_3917,N_3632);
xor U5377 (N_5377,N_677,N_2493);
nor U5378 (N_5378,N_1933,N_3888);
and U5379 (N_5379,N_459,N_3403);
nor U5380 (N_5380,N_1040,N_1479);
and U5381 (N_5381,N_1929,N_99);
or U5382 (N_5382,N_114,N_2539);
or U5383 (N_5383,N_3696,N_3161);
nand U5384 (N_5384,N_2587,N_4275);
nand U5385 (N_5385,N_2166,N_4927);
nand U5386 (N_5386,N_4755,N_1486);
xnor U5387 (N_5387,N_3208,N_1623);
xnor U5388 (N_5388,N_536,N_3565);
nor U5389 (N_5389,N_447,N_3416);
xor U5390 (N_5390,N_4883,N_3740);
nor U5391 (N_5391,N_3411,N_256);
nor U5392 (N_5392,N_1278,N_3058);
or U5393 (N_5393,N_3296,N_529);
nor U5394 (N_5394,N_1874,N_3395);
and U5395 (N_5395,N_4226,N_2688);
and U5396 (N_5396,N_3798,N_2738);
and U5397 (N_5397,N_398,N_4425);
nor U5398 (N_5398,N_1820,N_944);
nor U5399 (N_5399,N_2278,N_1266);
or U5400 (N_5400,N_913,N_4795);
nor U5401 (N_5401,N_4074,N_1864);
and U5402 (N_5402,N_4214,N_1937);
and U5403 (N_5403,N_356,N_2039);
and U5404 (N_5404,N_3595,N_2755);
or U5405 (N_5405,N_3780,N_2421);
xor U5406 (N_5406,N_2371,N_3172);
or U5407 (N_5407,N_414,N_1224);
nand U5408 (N_5408,N_4732,N_3698);
nand U5409 (N_5409,N_521,N_4100);
or U5410 (N_5410,N_842,N_1967);
nand U5411 (N_5411,N_3525,N_3400);
or U5412 (N_5412,N_2060,N_2758);
and U5413 (N_5413,N_895,N_4871);
and U5414 (N_5414,N_3504,N_1689);
nand U5415 (N_5415,N_1147,N_3613);
nor U5416 (N_5416,N_2080,N_3697);
nand U5417 (N_5417,N_1037,N_1962);
or U5418 (N_5418,N_3660,N_2178);
or U5419 (N_5419,N_2009,N_2191);
and U5420 (N_5420,N_3563,N_1829);
or U5421 (N_5421,N_4369,N_3392);
nor U5422 (N_5422,N_3585,N_3873);
or U5423 (N_5423,N_1028,N_4928);
or U5424 (N_5424,N_945,N_1672);
xnor U5425 (N_5425,N_1019,N_4334);
nor U5426 (N_5426,N_3074,N_1914);
or U5427 (N_5427,N_911,N_2830);
and U5428 (N_5428,N_4198,N_1921);
nand U5429 (N_5429,N_4974,N_937);
and U5430 (N_5430,N_4934,N_2360);
nand U5431 (N_5431,N_1307,N_2046);
or U5432 (N_5432,N_1983,N_1909);
nand U5433 (N_5433,N_4296,N_3047);
nor U5434 (N_5434,N_3033,N_4669);
or U5435 (N_5435,N_4779,N_1304);
nor U5436 (N_5436,N_3328,N_4308);
nor U5437 (N_5437,N_66,N_4009);
and U5438 (N_5438,N_3750,N_1243);
and U5439 (N_5439,N_4981,N_4481);
and U5440 (N_5440,N_4607,N_2029);
nand U5441 (N_5441,N_1204,N_3638);
nor U5442 (N_5442,N_1840,N_715);
nand U5443 (N_5443,N_3191,N_1039);
or U5444 (N_5444,N_4462,N_2065);
and U5445 (N_5445,N_1748,N_4192);
nor U5446 (N_5446,N_4580,N_901);
or U5447 (N_5447,N_2235,N_4891);
and U5448 (N_5448,N_4001,N_867);
nor U5449 (N_5449,N_2034,N_38);
and U5450 (N_5450,N_2699,N_41);
or U5451 (N_5451,N_3010,N_666);
nor U5452 (N_5452,N_566,N_802);
or U5453 (N_5453,N_3593,N_2650);
nand U5454 (N_5454,N_2707,N_2764);
and U5455 (N_5455,N_4724,N_2453);
nand U5456 (N_5456,N_2854,N_3515);
nand U5457 (N_5457,N_2052,N_957);
and U5458 (N_5458,N_570,N_4103);
nand U5459 (N_5459,N_3417,N_2592);
or U5460 (N_5460,N_2326,N_1600);
or U5461 (N_5461,N_308,N_657);
and U5462 (N_5462,N_4729,N_3836);
nor U5463 (N_5463,N_2671,N_4992);
nor U5464 (N_5464,N_3616,N_3007);
nor U5465 (N_5465,N_1995,N_4897);
and U5466 (N_5466,N_3694,N_1142);
and U5467 (N_5467,N_1137,N_3197);
or U5468 (N_5468,N_1693,N_3577);
and U5469 (N_5469,N_402,N_996);
nor U5470 (N_5470,N_1942,N_3971);
or U5471 (N_5471,N_2637,N_4518);
nand U5472 (N_5472,N_2159,N_4117);
nand U5473 (N_5473,N_4338,N_1045);
and U5474 (N_5474,N_2041,N_3380);
nor U5475 (N_5475,N_4448,N_3227);
nor U5476 (N_5476,N_2574,N_926);
and U5477 (N_5477,N_1632,N_2450);
nor U5478 (N_5478,N_3484,N_644);
or U5479 (N_5479,N_405,N_1181);
and U5480 (N_5480,N_2784,N_334);
and U5481 (N_5481,N_3244,N_3266);
and U5482 (N_5482,N_1505,N_4228);
nor U5483 (N_5483,N_1331,N_1320);
and U5484 (N_5484,N_1799,N_74);
nand U5485 (N_5485,N_4980,N_54);
nand U5486 (N_5486,N_1435,N_2555);
and U5487 (N_5487,N_1106,N_4356);
nand U5488 (N_5488,N_2461,N_1391);
nor U5489 (N_5489,N_4948,N_2803);
xor U5490 (N_5490,N_965,N_3947);
and U5491 (N_5491,N_1823,N_955);
nor U5492 (N_5492,N_3628,N_1252);
nand U5493 (N_5493,N_3220,N_624);
nor U5494 (N_5494,N_4805,N_1865);
nand U5495 (N_5495,N_2792,N_3826);
and U5496 (N_5496,N_1989,N_887);
and U5497 (N_5497,N_158,N_820);
nor U5498 (N_5498,N_2037,N_3357);
nor U5499 (N_5499,N_991,N_3090);
nor U5500 (N_5500,N_86,N_1118);
and U5501 (N_5501,N_46,N_2499);
nor U5502 (N_5502,N_147,N_3473);
nor U5503 (N_5503,N_1210,N_694);
or U5504 (N_5504,N_1163,N_4152);
or U5505 (N_5505,N_2640,N_4952);
or U5506 (N_5506,N_2056,N_1628);
and U5507 (N_5507,N_1860,N_3777);
and U5508 (N_5508,N_1735,N_3083);
nand U5509 (N_5509,N_2048,N_4067);
or U5510 (N_5510,N_4972,N_4723);
and U5511 (N_5511,N_2019,N_2702);
nand U5512 (N_5512,N_4830,N_550);
or U5513 (N_5513,N_3145,N_240);
nand U5514 (N_5514,N_3350,N_921);
or U5515 (N_5515,N_2395,N_1598);
and U5516 (N_5516,N_592,N_2152);
or U5517 (N_5517,N_3141,N_2418);
nand U5518 (N_5518,N_3624,N_4888);
nand U5519 (N_5519,N_909,N_1259);
and U5520 (N_5520,N_749,N_1182);
nor U5521 (N_5521,N_2911,N_2956);
and U5522 (N_5522,N_3056,N_4744);
or U5523 (N_5523,N_4507,N_2514);
nor U5524 (N_5524,N_1660,N_2343);
nand U5525 (N_5525,N_2710,N_4126);
or U5526 (N_5526,N_2692,N_4298);
nor U5527 (N_5527,N_3749,N_1465);
nand U5528 (N_5528,N_2391,N_3278);
nand U5529 (N_5529,N_1875,N_4984);
nor U5530 (N_5530,N_3737,N_3219);
and U5531 (N_5531,N_3255,N_1678);
nand U5532 (N_5532,N_2429,N_3158);
xor U5533 (N_5533,N_883,N_3333);
and U5534 (N_5534,N_4717,N_1593);
nand U5535 (N_5535,N_4016,N_620);
or U5536 (N_5536,N_2208,N_4273);
or U5537 (N_5537,N_4941,N_1732);
nor U5538 (N_5538,N_2331,N_3875);
and U5539 (N_5539,N_4353,N_1498);
or U5540 (N_5540,N_2902,N_1073);
or U5541 (N_5541,N_2144,N_2174);
and U5542 (N_5542,N_4701,N_615);
and U5543 (N_5543,N_2593,N_4819);
nor U5544 (N_5544,N_1835,N_3279);
or U5545 (N_5545,N_1041,N_2275);
nor U5546 (N_5546,N_4261,N_4277);
nand U5547 (N_5547,N_4143,N_3982);
nand U5548 (N_5548,N_671,N_107);
or U5549 (N_5549,N_3202,N_983);
nand U5550 (N_5550,N_1572,N_101);
and U5551 (N_5551,N_3329,N_675);
or U5552 (N_5552,N_3796,N_1074);
nand U5553 (N_5553,N_1488,N_2938);
and U5554 (N_5554,N_1188,N_3457);
nor U5555 (N_5555,N_2713,N_3081);
nor U5556 (N_5556,N_3960,N_3561);
xor U5557 (N_5557,N_1581,N_461);
nand U5558 (N_5558,N_3299,N_1692);
or U5559 (N_5559,N_4281,N_332);
nand U5560 (N_5560,N_1755,N_2335);
nor U5561 (N_5561,N_3931,N_3973);
and U5562 (N_5562,N_2303,N_2772);
and U5563 (N_5563,N_1379,N_1975);
and U5564 (N_5564,N_3566,N_3397);
and U5565 (N_5565,N_2473,N_219);
or U5566 (N_5566,N_3022,N_4837);
or U5567 (N_5567,N_1077,N_4780);
nand U5568 (N_5568,N_4064,N_4877);
nor U5569 (N_5569,N_4720,N_4122);
or U5570 (N_5570,N_215,N_3127);
nor U5571 (N_5571,N_3231,N_1963);
and U5572 (N_5572,N_1207,N_2958);
and U5573 (N_5573,N_4182,N_3871);
nand U5574 (N_5574,N_1997,N_3975);
or U5575 (N_5575,N_184,N_1740);
or U5576 (N_5576,N_1930,N_2021);
and U5577 (N_5577,N_2198,N_301);
or U5578 (N_5578,N_2372,N_2926);
nand U5579 (N_5579,N_3420,N_607);
or U5580 (N_5580,N_4488,N_2927);
xor U5581 (N_5581,N_3485,N_1954);
and U5582 (N_5582,N_1808,N_2192);
nand U5583 (N_5583,N_1590,N_1908);
or U5584 (N_5584,N_4211,N_2666);
xnor U5585 (N_5585,N_131,N_1322);
nand U5586 (N_5586,N_2363,N_42);
nand U5587 (N_5587,N_141,N_4268);
or U5588 (N_5588,N_2096,N_3783);
nor U5589 (N_5589,N_587,N_3617);
nor U5590 (N_5590,N_4063,N_795);
xnor U5591 (N_5591,N_3272,N_3096);
or U5592 (N_5592,N_4604,N_920);
and U5593 (N_5593,N_640,N_244);
or U5594 (N_5594,N_4413,N_3453);
nand U5595 (N_5595,N_166,N_3001);
nand U5596 (N_5596,N_3339,N_1769);
nand U5597 (N_5597,N_148,N_4567);
nand U5598 (N_5598,N_4087,N_3434);
and U5599 (N_5599,N_668,N_3746);
and U5600 (N_5600,N_4041,N_3997);
and U5601 (N_5601,N_4525,N_1744);
nand U5602 (N_5602,N_4550,N_1005);
nand U5603 (N_5603,N_4443,N_4594);
nand U5604 (N_5604,N_1770,N_4221);
nand U5605 (N_5605,N_3039,N_1446);
nand U5606 (N_5606,N_496,N_123);
and U5607 (N_5607,N_3690,N_476);
and U5608 (N_5608,N_3250,N_3112);
nand U5609 (N_5609,N_3302,N_2413);
or U5610 (N_5610,N_2253,N_1896);
nor U5611 (N_5611,N_377,N_3338);
or U5612 (N_5612,N_4310,N_1254);
nand U5613 (N_5613,N_1711,N_3020);
and U5614 (N_5614,N_3778,N_2074);
nand U5615 (N_5615,N_1049,N_4708);
and U5616 (N_5616,N_3106,N_1282);
nor U5617 (N_5617,N_1483,N_2635);
xor U5618 (N_5618,N_2660,N_2022);
nor U5619 (N_5619,N_40,N_4188);
nor U5620 (N_5620,N_57,N_1180);
or U5621 (N_5621,N_266,N_1597);
or U5622 (N_5622,N_1580,N_2925);
nand U5623 (N_5623,N_4364,N_324);
and U5624 (N_5624,N_792,N_3150);
nor U5625 (N_5625,N_1508,N_1733);
or U5626 (N_5626,N_3574,N_3770);
or U5627 (N_5627,N_1442,N_2850);
and U5628 (N_5628,N_1154,N_1054);
and U5629 (N_5629,N_3174,N_721);
and U5630 (N_5630,N_52,N_279);
nor U5631 (N_5631,N_3017,N_2914);
nand U5632 (N_5632,N_1059,N_385);
nand U5633 (N_5633,N_3476,N_2687);
nand U5634 (N_5634,N_4599,N_1410);
and U5635 (N_5635,N_4849,N_635);
nor U5636 (N_5636,N_1325,N_1830);
or U5637 (N_5637,N_1986,N_351);
or U5638 (N_5638,N_1104,N_1506);
nand U5639 (N_5639,N_2273,N_811);
nand U5640 (N_5640,N_280,N_2027);
nor U5641 (N_5641,N_2201,N_1246);
nor U5642 (N_5642,N_572,N_1972);
nand U5643 (N_5643,N_1635,N_3111);
or U5644 (N_5644,N_2344,N_4690);
or U5645 (N_5645,N_1555,N_1399);
nand U5646 (N_5646,N_3516,N_1826);
nor U5647 (N_5647,N_268,N_327);
nand U5648 (N_5648,N_1128,N_237);
nor U5649 (N_5649,N_4046,N_3865);
and U5650 (N_5650,N_3084,N_3748);
or U5651 (N_5651,N_272,N_1797);
nand U5652 (N_5652,N_2594,N_4437);
nand U5653 (N_5653,N_4485,N_392);
and U5654 (N_5654,N_3175,N_4183);
and U5655 (N_5655,N_3630,N_4799);
and U5656 (N_5656,N_208,N_4499);
or U5657 (N_5657,N_691,N_1035);
or U5658 (N_5658,N_1202,N_4204);
nand U5659 (N_5659,N_206,N_1150);
nor U5660 (N_5660,N_4531,N_3825);
nor U5661 (N_5661,N_3480,N_3966);
nand U5662 (N_5662,N_2423,N_667);
nand U5663 (N_5663,N_2426,N_3976);
and U5664 (N_5664,N_1952,N_1504);
nand U5665 (N_5665,N_14,N_1226);
nand U5666 (N_5666,N_3978,N_1531);
and U5667 (N_5667,N_4710,N_1273);
nand U5668 (N_5668,N_653,N_3654);
or U5669 (N_5669,N_704,N_4243);
or U5670 (N_5670,N_4902,N_2251);
xor U5671 (N_5671,N_4370,N_2488);
or U5672 (N_5672,N_413,N_736);
and U5673 (N_5673,N_1904,N_3314);
and U5674 (N_5674,N_1274,N_173);
nor U5675 (N_5675,N_695,N_2276);
xor U5676 (N_5676,N_4039,N_3863);
or U5677 (N_5677,N_3967,N_3353);
and U5678 (N_5678,N_4794,N_2400);
nand U5679 (N_5679,N_2703,N_1174);
nor U5680 (N_5680,N_1265,N_4756);
and U5681 (N_5681,N_1494,N_371);
and U5682 (N_5682,N_4254,N_4621);
and U5683 (N_5683,N_1287,N_4240);
and U5684 (N_5684,N_2822,N_4377);
nor U5685 (N_5685,N_3012,N_2410);
and U5686 (N_5686,N_3897,N_170);
nor U5687 (N_5687,N_444,N_69);
or U5688 (N_5688,N_4661,N_3062);
and U5689 (N_5689,N_3211,N_3360);
or U5690 (N_5690,N_235,N_2795);
and U5691 (N_5691,N_1890,N_854);
nand U5692 (N_5692,N_3803,N_1585);
nand U5693 (N_5693,N_2775,N_4045);
or U5694 (N_5694,N_3665,N_4808);
nor U5695 (N_5695,N_538,N_3233);
or U5696 (N_5696,N_89,N_4523);
and U5697 (N_5697,N_238,N_1712);
nand U5698 (N_5698,N_203,N_4289);
nor U5699 (N_5699,N_4999,N_4673);
and U5700 (N_5700,N_747,N_956);
and U5701 (N_5701,N_4659,N_845);
nor U5702 (N_5702,N_4534,N_679);
nand U5703 (N_5703,N_2240,N_352);
nor U5704 (N_5704,N_3262,N_2536);
or U5705 (N_5705,N_4132,N_1788);
nor U5706 (N_5706,N_2686,N_1703);
nor U5707 (N_5707,N_4826,N_3459);
nand U5708 (N_5708,N_149,N_3985);
and U5709 (N_5709,N_3388,N_4258);
nand U5710 (N_5710,N_4656,N_138);
and U5711 (N_5711,N_3604,N_1833);
and U5712 (N_5712,N_3312,N_456);
or U5713 (N_5713,N_4938,N_2805);
and U5714 (N_5714,N_2061,N_1055);
and U5715 (N_5715,N_3157,N_1527);
and U5716 (N_5716,N_3438,N_2339);
and U5717 (N_5717,N_3035,N_2407);
and U5718 (N_5718,N_2392,N_3006);
nand U5719 (N_5719,N_595,N_1400);
or U5720 (N_5720,N_2763,N_1081);
nand U5721 (N_5721,N_1004,N_3760);
nor U5722 (N_5722,N_2487,N_688);
nor U5723 (N_5723,N_2300,N_3881);
nor U5724 (N_5724,N_381,N_3198);
or U5725 (N_5725,N_4098,N_2347);
and U5726 (N_5726,N_4784,N_3639);
and U5727 (N_5727,N_2590,N_2787);
and U5728 (N_5728,N_63,N_597);
nand U5729 (N_5729,N_851,N_1038);
nand U5730 (N_5730,N_464,N_2219);
or U5731 (N_5731,N_1853,N_807);
nor U5732 (N_5732,N_830,N_1831);
and U5733 (N_5733,N_2569,N_2623);
nand U5734 (N_5734,N_3315,N_3503);
and U5735 (N_5735,N_1064,N_3068);
and U5736 (N_5736,N_3094,N_189);
nand U5737 (N_5737,N_90,N_614);
nor U5738 (N_5738,N_3933,N_3215);
nor U5739 (N_5739,N_4545,N_4224);
nor U5740 (N_5740,N_1587,N_1676);
nor U5741 (N_5741,N_3965,N_877);
nand U5742 (N_5742,N_1708,N_3274);
nand U5743 (N_5743,N_3065,N_642);
nor U5744 (N_5744,N_2991,N_1239);
and U5745 (N_5745,N_4561,N_577);
nand U5746 (N_5746,N_2748,N_2025);
and U5747 (N_5747,N_2523,N_3366);
nand U5748 (N_5748,N_2102,N_3536);
nor U5749 (N_5749,N_471,N_3486);
and U5750 (N_5750,N_4412,N_4781);
nor U5751 (N_5751,N_4588,N_1375);
nor U5752 (N_5752,N_3681,N_3070);
nor U5753 (N_5753,N_2282,N_1146);
nand U5754 (N_5754,N_3572,N_2676);
nor U5755 (N_5755,N_4995,N_34);
and U5756 (N_5756,N_1421,N_168);
nand U5757 (N_5757,N_870,N_1719);
nand U5758 (N_5758,N_2579,N_1721);
and U5759 (N_5759,N_1219,N_2669);
or U5760 (N_5760,N_349,N_545);
nor U5761 (N_5761,N_1382,N_1528);
nand U5762 (N_5762,N_4287,N_773);
or U5763 (N_5763,N_2090,N_995);
nand U5764 (N_5764,N_4337,N_547);
or U5765 (N_5765,N_2337,N_3118);
nand U5766 (N_5766,N_873,N_3601);
or U5767 (N_5767,N_4011,N_264);
nand U5768 (N_5768,N_1603,N_875);
or U5769 (N_5769,N_2492,N_4616);
nor U5770 (N_5770,N_1656,N_1427);
or U5771 (N_5771,N_1900,N_1884);
nor U5772 (N_5772,N_4300,N_3498);
nand U5773 (N_5773,N_430,N_4924);
nor U5774 (N_5774,N_4649,N_4190);
or U5775 (N_5775,N_4362,N_3575);
nor U5776 (N_5776,N_4982,N_2472);
nor U5777 (N_5777,N_4033,N_4538);
or U5778 (N_5778,N_2330,N_3747);
or U5779 (N_5779,N_4451,N_199);
and U5780 (N_5780,N_317,N_2187);
and U5781 (N_5781,N_3528,N_4060);
nand U5782 (N_5782,N_1023,N_2729);
nor U5783 (N_5783,N_4773,N_2695);
or U5784 (N_5784,N_2503,N_1497);
or U5785 (N_5785,N_3003,N_445);
nand U5786 (N_5786,N_3317,N_4219);
and U5787 (N_5787,N_1839,N_1372);
nand U5788 (N_5788,N_2245,N_2173);
nor U5789 (N_5789,N_4577,N_669);
and U5790 (N_5790,N_2947,N_474);
and U5791 (N_5791,N_766,N_2813);
or U5792 (N_5792,N_4309,N_4502);
xnor U5793 (N_5793,N_156,N_210);
or U5794 (N_5794,N_4581,N_288);
and U5795 (N_5795,N_3943,N_290);
and U5796 (N_5796,N_1918,N_1649);
nor U5797 (N_5797,N_1608,N_3492);
nor U5798 (N_5798,N_81,N_3069);
nand U5799 (N_5799,N_4231,N_3248);
or U5800 (N_5800,N_3384,N_4572);
and U5801 (N_5801,N_1779,N_3241);
nor U5802 (N_5802,N_4787,N_709);
or U5803 (N_5803,N_599,N_3531);
nand U5804 (N_5804,N_1398,N_2229);
or U5805 (N_5805,N_3479,N_2736);
nor U5806 (N_5806,N_935,N_159);
and U5807 (N_5807,N_2271,N_4949);
nor U5808 (N_5808,N_4554,N_4602);
or U5809 (N_5809,N_4395,N_345);
and U5810 (N_5810,N_4438,N_1153);
nor U5811 (N_5811,N_1611,N_2769);
and U5812 (N_5812,N_3883,N_2155);
xnor U5813 (N_5813,N_3337,N_2322);
xor U5814 (N_5814,N_4666,N_3922);
nand U5815 (N_5815,N_2115,N_604);
or U5816 (N_5816,N_1261,N_2768);
nand U5817 (N_5817,N_172,N_1222);
and U5818 (N_5818,N_2387,N_333);
xor U5819 (N_5819,N_790,N_129);
and U5820 (N_5820,N_1302,N_3300);
nor U5821 (N_5821,N_3183,N_4466);
nor U5822 (N_5822,N_3002,N_4645);
or U5823 (N_5823,N_1520,N_436);
nand U5824 (N_5824,N_4085,N_3850);
nand U5825 (N_5825,N_1898,N_4603);
nand U5826 (N_5826,N_4946,N_3451);
nor U5827 (N_5827,N_713,N_1369);
nand U5828 (N_5828,N_1057,N_4696);
or U5829 (N_5829,N_3109,N_1730);
nand U5830 (N_5830,N_4343,N_3963);
or U5831 (N_5831,N_1913,N_262);
or U5832 (N_5832,N_1363,N_1714);
or U5833 (N_5833,N_4800,N_2665);
nand U5834 (N_5834,N_2211,N_1985);
or U5835 (N_5835,N_2643,N_3097);
nand U5836 (N_5836,N_3735,N_4774);
nor U5837 (N_5837,N_1679,N_742);
and U5838 (N_5838,N_4248,N_4699);
or U5839 (N_5839,N_2279,N_3693);
and U5840 (N_5840,N_598,N_2068);
or U5841 (N_5841,N_3467,N_1395);
nand U5842 (N_5842,N_2143,N_992);
and U5843 (N_5843,N_2517,N_3821);
and U5844 (N_5844,N_2055,N_1793);
nor U5845 (N_5845,N_3652,N_2464);
or U5846 (N_5846,N_664,N_1396);
and U5847 (N_5847,N_1547,N_3675);
nand U5848 (N_5848,N_304,N_888);
or U5849 (N_5849,N_316,N_3684);
nor U5850 (N_5850,N_3679,N_2230);
or U5851 (N_5851,N_4597,N_1083);
nor U5852 (N_5852,N_4688,N_336);
and U5853 (N_5853,N_1866,N_1377);
and U5854 (N_5854,N_4793,N_4082);
and U5855 (N_5855,N_30,N_879);
or U5856 (N_5856,N_4873,N_439);
and U5857 (N_5857,N_1969,N_2302);
xnor U5858 (N_5858,N_2367,N_1221);
and U5859 (N_5859,N_4172,N_2901);
or U5860 (N_5860,N_971,N_1782);
or U5861 (N_5861,N_221,N_1105);
nor U5862 (N_5862,N_4389,N_4921);
nand U5863 (N_5863,N_1414,N_2194);
or U5864 (N_5864,N_2242,N_2557);
nand U5865 (N_5865,N_2533,N_3064);
or U5866 (N_5866,N_2691,N_4054);
and U5867 (N_5867,N_3764,N_396);
or U5868 (N_5868,N_1192,N_1926);
or U5869 (N_5869,N_4815,N_4153);
or U5870 (N_5870,N_4406,N_3114);
and U5871 (N_5871,N_2716,N_3316);
nor U5872 (N_5872,N_4547,N_3055);
nor U5873 (N_5873,N_4269,N_761);
nor U5874 (N_5874,N_649,N_4501);
nor U5875 (N_5875,N_2483,N_1112);
nor U5876 (N_5876,N_1868,N_3910);
xnor U5877 (N_5877,N_108,N_2870);
and U5878 (N_5878,N_4790,N_2528);
nor U5879 (N_5879,N_1633,N_2341);
or U5880 (N_5880,N_1588,N_1822);
nand U5881 (N_5881,N_4487,N_4685);
and U5882 (N_5882,N_2113,N_1683);
and U5883 (N_5883,N_2834,N_2823);
and U5884 (N_5884,N_4227,N_466);
nor U5885 (N_5885,N_1776,N_4668);
nor U5886 (N_5886,N_406,N_3713);
nand U5887 (N_5887,N_789,N_1938);
nand U5888 (N_5888,N_4315,N_1976);
and U5889 (N_5889,N_424,N_533);
nand U5890 (N_5890,N_4742,N_2705);
or U5891 (N_5891,N_3587,N_3622);
nand U5892 (N_5892,N_3325,N_137);
and U5893 (N_5893,N_1021,N_251);
nand U5894 (N_5894,N_2613,N_1801);
and U5895 (N_5895,N_340,N_643);
nand U5896 (N_5896,N_2818,N_3009);
or U5897 (N_5897,N_541,N_629);
nor U5898 (N_5898,N_3352,N_4255);
nand U5899 (N_5899,N_344,N_1339);
nor U5900 (N_5900,N_4166,N_2513);
or U5901 (N_5901,N_2066,N_1810);
nand U5902 (N_5902,N_4199,N_3285);
and U5903 (N_5903,N_858,N_4747);
and U5904 (N_5904,N_4760,N_4806);
xor U5905 (N_5905,N_4731,N_3364);
and U5906 (N_5906,N_3209,N_2087);
nor U5907 (N_5907,N_2906,N_1715);
nand U5908 (N_5908,N_3551,N_3268);
and U5909 (N_5909,N_3867,N_951);
nand U5910 (N_5910,N_3301,N_281);
or U5911 (N_5911,N_1176,N_357);
xor U5912 (N_5912,N_1629,N_814);
and U5913 (N_5913,N_319,N_3399);
and U5914 (N_5914,N_3188,N_4886);
nor U5915 (N_5915,N_154,N_3271);
and U5916 (N_5916,N_2017,N_4391);
nor U5917 (N_5917,N_1789,N_1984);
nand U5918 (N_5918,N_4038,N_1238);
nor U5919 (N_5919,N_2694,N_3345);
nand U5920 (N_5920,N_4913,N_968);
or U5921 (N_5921,N_115,N_1798);
or U5922 (N_5922,N_490,N_4869);
nand U5923 (N_5923,N_4336,N_528);
or U5924 (N_5924,N_3619,N_1964);
and U5925 (N_5925,N_135,N_1216);
nor U5926 (N_5926,N_781,N_535);
and U5927 (N_5927,N_2706,N_3828);
or U5928 (N_5928,N_1576,N_3802);
and U5929 (N_5929,N_903,N_3990);
or U5930 (N_5930,N_428,N_198);
or U5931 (N_5931,N_626,N_826);
nand U5932 (N_5932,N_3722,N_1114);
nor U5933 (N_5933,N_1845,N_726);
and U5934 (N_5934,N_3858,N_919);
nor U5935 (N_5935,N_889,N_1308);
nand U5936 (N_5936,N_1753,N_1807);
or U5937 (N_5937,N_2596,N_3218);
nand U5938 (N_5938,N_3060,N_2819);
and U5939 (N_5939,N_1741,N_3464);
and U5940 (N_5940,N_3015,N_4019);
nand U5941 (N_5941,N_4191,N_1365);
nor U5942 (N_5942,N_1102,N_407);
or U5943 (N_5943,N_3098,N_2393);
nand U5944 (N_5944,N_897,N_2722);
or U5945 (N_5945,N_2801,N_1768);
and U5946 (N_5946,N_2737,N_591);
nand U5947 (N_5947,N_772,N_2670);
nand U5948 (N_5948,N_1214,N_4727);
or U5949 (N_5949,N_259,N_2506);
nor U5950 (N_5950,N_2624,N_812);
nor U5951 (N_5951,N_4392,N_4601);
or U5952 (N_5952,N_358,N_4825);
nor U5953 (N_5953,N_3543,N_2239);
and U5954 (N_5954,N_4266,N_3815);
or U5955 (N_5955,N_2960,N_596);
nor U5956 (N_5956,N_4115,N_1166);
nor U5957 (N_5957,N_144,N_3119);
nor U5958 (N_5958,N_3596,N_2735);
or U5959 (N_5959,N_2088,N_586);
nand U5960 (N_5960,N_2512,N_3711);
xor U5961 (N_5961,N_511,N_4674);
and U5962 (N_5962,N_4382,N_2332);
or U5963 (N_5963,N_2791,N_4018);
or U5964 (N_5964,N_619,N_4396);
nand U5965 (N_5965,N_3275,N_2989);
and U5966 (N_5966,N_2542,N_1444);
nand U5967 (N_5967,N_3680,N_1397);
and U5968 (N_5968,N_1276,N_822);
or U5969 (N_5969,N_2281,N_3348);
nand U5970 (N_5970,N_1225,N_2280);
or U5971 (N_5971,N_809,N_4887);
and U5972 (N_5972,N_4196,N_2782);
nor U5973 (N_5973,N_3042,N_1422);
or U5974 (N_5974,N_3972,N_3071);
and U5975 (N_5975,N_1120,N_2180);
or U5976 (N_5976,N_4520,N_4903);
nor U5977 (N_5977,N_4155,N_3647);
or U5978 (N_5978,N_648,N_2725);
or U5979 (N_5979,N_2157,N_2292);
nor U5980 (N_5980,N_303,N_4521);
and U5981 (N_5981,N_4788,N_4931);
and U5982 (N_5982,N_2639,N_3571);
or U5983 (N_5983,N_2937,N_2615);
and U5984 (N_5984,N_3028,N_1869);
xnor U5985 (N_5985,N_4700,N_701);
or U5986 (N_5986,N_4108,N_1149);
nor U5987 (N_5987,N_373,N_4624);
or U5988 (N_5988,N_3984,N_2859);
nand U5989 (N_5989,N_1231,N_1177);
or U5990 (N_5990,N_1570,N_3762);
nor U5991 (N_5991,N_4208,N_3940);
nand U5992 (N_5992,N_4953,N_4445);
nand U5993 (N_5993,N_3212,N_4209);
nor U5994 (N_5994,N_1393,N_4469);
or U5995 (N_5995,N_3410,N_3246);
and U5996 (N_5996,N_341,N_1947);
or U5997 (N_5997,N_3581,N_4942);
nor U5998 (N_5998,N_1893,N_4482);
nor U5999 (N_5999,N_3456,N_3914);
and U6000 (N_6000,N_65,N_4272);
and U6001 (N_6001,N_1837,N_3419);
and U6002 (N_6002,N_2584,N_526);
or U6003 (N_6003,N_633,N_4945);
xor U6004 (N_6004,N_3609,N_2213);
nand U6005 (N_6005,N_3126,N_4031);
and U6006 (N_6006,N_3956,N_4450);
or U6007 (N_6007,N_3822,N_2457);
nand U6008 (N_6008,N_1999,N_791);
nand U6009 (N_6009,N_1795,N_4223);
or U6010 (N_6010,N_51,N_4912);
or U6011 (N_6011,N_1720,N_2757);
or U6012 (N_6012,N_3290,N_174);
and U6013 (N_6013,N_2952,N_768);
xnor U6014 (N_6014,N_2527,N_214);
xor U6015 (N_6015,N_18,N_3835);
or U6016 (N_6016,N_1453,N_4767);
nand U6017 (N_6017,N_994,N_4139);
nor U6018 (N_6018,N_3653,N_1489);
nand U6019 (N_6019,N_1450,N_4029);
and U6020 (N_6020,N_4194,N_4703);
nand U6021 (N_6021,N_1385,N_2505);
nand U6022 (N_6022,N_3939,N_3774);
and U6023 (N_6023,N_3475,N_3685);
or U6024 (N_6024,N_1852,N_3166);
and U6025 (N_6025,N_2583,N_705);
nand U6026 (N_6026,N_1849,N_4555);
and U6027 (N_6027,N_4311,N_507);
or U6028 (N_6028,N_739,N_193);
or U6029 (N_6029,N_4002,N_4106);
or U6030 (N_6030,N_904,N_2700);
nor U6031 (N_6031,N_1386,N_3655);
nand U6032 (N_6032,N_3788,N_4670);
nor U6033 (N_6033,N_4510,N_3772);
xor U6034 (N_6034,N_418,N_467);
and U6035 (N_6035,N_1502,N_2405);
nor U6036 (N_6036,N_2311,N_225);
nand U6037 (N_6037,N_4969,N_797);
nand U6038 (N_6038,N_3247,N_1885);
or U6039 (N_6039,N_3313,N_3207);
xor U6040 (N_6040,N_553,N_1327);
nand U6041 (N_6041,N_2681,N_2963);
and U6042 (N_6042,N_2319,N_224);
nor U6043 (N_6043,N_106,N_1283);
nand U6044 (N_6044,N_20,N_1534);
and U6045 (N_6045,N_2297,N_735);
nor U6046 (N_6046,N_2139,N_4527);
nor U6047 (N_6047,N_1763,N_717);
nor U6048 (N_6048,N_504,N_4824);
nor U6049 (N_6049,N_2999,N_2611);
or U6050 (N_6050,N_1171,N_2644);
nand U6051 (N_6051,N_906,N_2399);
or U6052 (N_6052,N_4358,N_2109);
nor U6053 (N_6053,N_3310,N_2500);
nor U6054 (N_6054,N_2882,N_612);
and U6055 (N_6055,N_1474,N_169);
nand U6056 (N_6056,N_1800,N_119);
nor U6057 (N_6057,N_2382,N_1121);
and U6058 (N_6058,N_375,N_2188);
nand U6059 (N_6059,N_2054,N_1616);
and U6060 (N_6060,N_1255,N_465);
nand U6061 (N_6061,N_4447,N_3041);
and U6062 (N_6062,N_2714,N_878);
or U6063 (N_6063,N_4613,N_850);
and U6064 (N_6064,N_3854,N_874);
nor U6065 (N_6065,N_3529,N_3974);
nor U6066 (N_6066,N_2978,N_4096);
nand U6067 (N_6067,N_2362,N_246);
and U6068 (N_6068,N_4301,N_1695);
and U6069 (N_6069,N_2985,N_1617);
and U6070 (N_6070,N_4420,N_1336);
nand U6071 (N_6071,N_2804,N_2436);
and U6072 (N_6072,N_2740,N_1583);
and U6073 (N_6073,N_1227,N_835);
and U6074 (N_6074,N_2111,N_934);
or U6075 (N_6075,N_4622,N_4907);
and U6076 (N_6076,N_1901,N_3178);
and U6077 (N_6077,N_4737,N_4875);
nor U6078 (N_6078,N_2170,N_233);
nor U6079 (N_6079,N_2225,N_4979);
and U6080 (N_6080,N_3235,N_3657);
nand U6081 (N_6081,N_4142,N_2881);
nor U6082 (N_6082,N_1079,N_2711);
nor U6083 (N_6083,N_1677,N_4652);
and U6084 (N_6084,N_627,N_686);
and U6085 (N_6085,N_1536,N_3856);
and U6086 (N_6086,N_3996,N_4505);
nor U6087 (N_6087,N_4872,N_7);
nor U6088 (N_6088,N_2105,N_3600);
nand U6089 (N_6089,N_1992,N_3323);
or U6090 (N_6090,N_3361,N_1910);
and U6091 (N_6091,N_818,N_1780);
or U6092 (N_6092,N_33,N_186);
and U6093 (N_6093,N_1844,N_2747);
and U6094 (N_6094,N_0,N_3663);
or U6095 (N_6095,N_2414,N_2324);
or U6096 (N_6096,N_3728,N_4286);
nor U6097 (N_6097,N_2630,N_3884);
and U6098 (N_6098,N_2366,N_4987);
or U6099 (N_6099,N_4608,N_4618);
nand U6100 (N_6100,N_562,N_2944);
and U6101 (N_6101,N_2137,N_645);
xor U6102 (N_6102,N_1542,N_2979);
or U6103 (N_6103,N_36,N_458);
nor U6104 (N_6104,N_2044,N_3130);
nand U6105 (N_6105,N_1449,N_775);
nand U6106 (N_6106,N_1699,N_330);
nand U6107 (N_6107,N_1205,N_841);
nand U6108 (N_6108,N_799,N_3950);
nand U6109 (N_6109,N_1922,N_499);
and U6110 (N_6110,N_3998,N_703);
or U6111 (N_6111,N_2226,N_4678);
and U6112 (N_6112,N_3186,N_4325);
nor U6113 (N_6113,N_3378,N_3462);
or U6114 (N_6114,N_4472,N_3298);
nor U6115 (N_6115,N_1065,N_1594);
nand U6116 (N_6116,N_2375,N_1098);
and U6117 (N_6117,N_4213,N_3903);
nor U6118 (N_6118,N_4162,N_3368);
or U6119 (N_6119,N_3452,N_423);
and U6120 (N_6120,N_383,N_3408);
or U6121 (N_6121,N_3754,N_2790);
nor U6122 (N_6122,N_2651,N_2816);
and U6123 (N_6123,N_984,N_949);
nand U6124 (N_6124,N_1848,N_2035);
and U6125 (N_6125,N_885,N_3330);
and U6126 (N_6126,N_4279,N_1939);
nand U6127 (N_6127,N_2917,N_492);
and U6128 (N_6128,N_4193,N_856);
and U6129 (N_6129,N_3631,N_3103);
nor U6130 (N_6130,N_4922,N_2942);
and U6131 (N_6131,N_658,N_3847);
or U6132 (N_6132,N_1032,N_4961);
nand U6133 (N_6133,N_755,N_3817);
nor U6134 (N_6134,N_2855,N_3104);
nand U6135 (N_6135,N_2274,N_833);
nand U6136 (N_6136,N_1710,N_961);
xor U6137 (N_6137,N_4777,N_4514);
or U6138 (N_6138,N_3813,N_3537);
nand U6139 (N_6139,N_3162,N_3341);
nand U6140 (N_6140,N_2667,N_1031);
nand U6141 (N_6141,N_2032,N_719);
nor U6142 (N_6142,N_2601,N_2443);
or U6143 (N_6143,N_3874,N_265);
and U6144 (N_6144,N_416,N_4929);
nor U6145 (N_6145,N_2063,N_307);
or U6146 (N_6146,N_1140,N_1682);
or U6147 (N_6147,N_714,N_4138);
and U6148 (N_6148,N_3072,N_53);
and U6149 (N_6149,N_1879,N_4844);
or U6150 (N_6150,N_4253,N_4776);
nand U6151 (N_6151,N_4489,N_3148);
nor U6152 (N_6152,N_3177,N_4684);
or U6153 (N_6153,N_4483,N_3390);
and U6154 (N_6154,N_2777,N_2449);
or U6155 (N_6155,N_3930,N_4133);
nor U6156 (N_6156,N_3763,N_2114);
nand U6157 (N_6157,N_3532,N_4323);
nor U6158 (N_6158,N_2572,N_1894);
nand U6159 (N_6159,N_1433,N_4910);
or U6160 (N_6160,N_4865,N_2998);
or U6161 (N_6161,N_2719,N_252);
and U6162 (N_6162,N_4498,N_3011);
nor U6163 (N_6163,N_1510,N_4722);
nand U6164 (N_6164,N_242,N_3402);
and U6165 (N_6165,N_3099,N_3253);
nand U6166 (N_6166,N_3530,N_4347);
nor U6167 (N_6167,N_2995,N_886);
or U6168 (N_6168,N_509,N_2477);
nor U6169 (N_6169,N_2390,N_120);
nand U6170 (N_6170,N_1796,N_1380);
nand U6171 (N_6171,N_798,N_4233);
nor U6172 (N_6172,N_1244,N_2977);
nor U6173 (N_6173,N_2831,N_3934);
nor U6174 (N_6174,N_270,N_4560);
and U6175 (N_6175,N_672,N_603);
nand U6176 (N_6176,N_1686,N_4313);
nor U6177 (N_6177,N_2595,N_201);
nand U6178 (N_6178,N_3448,N_1175);
nor U6179 (N_6179,N_4433,N_3469);
and U6180 (N_6180,N_1827,N_4691);
or U6181 (N_6181,N_3173,N_4383);
and U6182 (N_6182,N_2381,N_2868);
or U6183 (N_6183,N_1242,N_2142);
nand U6184 (N_6184,N_3969,N_2089);
or U6185 (N_6185,N_4032,N_3146);
nand U6186 (N_6186,N_1036,N_3494);
and U6187 (N_6187,N_1408,N_4968);
nor U6188 (N_6188,N_2228,N_4112);
or U6189 (N_6189,N_1299,N_1944);
nor U6190 (N_6190,N_1657,N_3995);
or U6191 (N_6191,N_4976,N_3626);
or U6192 (N_6192,N_1158,N_296);
nor U6193 (N_6193,N_1517,N_1361);
or U6194 (N_6194,N_1348,N_134);
nand U6195 (N_6195,N_328,N_1443);
and U6196 (N_6196,N_3044,N_1432);
or U6197 (N_6197,N_2398,N_600);
nand U6198 (N_6198,N_368,N_2767);
and U6199 (N_6199,N_1338,N_4197);
or U6200 (N_6200,N_4596,N_420);
nor U6201 (N_6201,N_139,N_3206);
or U6202 (N_6202,N_4167,N_22);
nand U6203 (N_6203,N_4216,N_4326);
or U6204 (N_6204,N_4812,N_3793);
nand U6205 (N_6205,N_3723,N_2128);
or U6206 (N_6206,N_2401,N_4442);
xnor U6207 (N_6207,N_3829,N_3128);
xnor U6208 (N_6208,N_1854,N_3831);
and U6209 (N_6209,N_3132,N_4642);
or U6210 (N_6210,N_3692,N_2918);
nor U6211 (N_6211,N_4850,N_967);
nor U6212 (N_6212,N_4403,N_3131);
nor U6213 (N_6213,N_365,N_3841);
nor U6214 (N_6214,N_3970,N_4073);
nor U6215 (N_6215,N_220,N_787);
or U6216 (N_6216,N_197,N_4863);
xor U6217 (N_6217,N_4339,N_2840);
nand U6218 (N_6218,N_2646,N_75);
or U6219 (N_6219,N_3115,N_1673);
or U6220 (N_6220,N_3535,N_412);
nand U6221 (N_6221,N_1388,N_1067);
and U6222 (N_6222,N_2496,N_2249);
nor U6223 (N_6223,N_3182,N_4562);
or U6224 (N_6224,N_2001,N_2910);
or U6225 (N_6225,N_4935,N_394);
and U6226 (N_6226,N_2672,N_740);
nand U6227 (N_6227,N_1337,N_2310);
nor U6228 (N_6228,N_2441,N_2968);
nand U6229 (N_6229,N_3488,N_1193);
or U6230 (N_6230,N_1493,N_1957);
and U6231 (N_6231,N_3929,N_1643);
and U6232 (N_6232,N_4239,N_1027);
nand U6233 (N_6233,N_3474,N_4130);
or U6234 (N_6234,N_3517,N_1314);
nand U6235 (N_6235,N_1544,N_1606);
and U6236 (N_6236,N_4168,N_2313);
nor U6237 (N_6237,N_3699,N_654);
or U6238 (N_6238,N_117,N_2183);
or U6239 (N_6239,N_3135,N_3633);
nor U6240 (N_6240,N_753,N_2415);
nand U6241 (N_6241,N_3846,N_673);
nand U6242 (N_6242,N_974,N_3369);
nand U6243 (N_6243,N_4444,N_4565);
nor U6244 (N_6244,N_485,N_3842);
and U6245 (N_6245,N_3487,N_2002);
and U6246 (N_6246,N_4962,N_4821);
and U6247 (N_6247,N_525,N_2799);
nand U6248 (N_6248,N_1668,N_49);
nand U6249 (N_6249,N_4232,N_2403);
nand U6250 (N_6250,N_2618,N_1862);
nand U6251 (N_6251,N_326,N_273);
nor U6252 (N_6252,N_4959,N_4176);
and U6253 (N_6253,N_37,N_4940);
nand U6254 (N_6254,N_1271,N_3851);
or U6255 (N_6255,N_646,N_2277);
or U6256 (N_6256,N_4177,N_239);
and U6257 (N_6257,N_759,N_518);
nor U6258 (N_6258,N_4090,N_440);
xnor U6259 (N_6259,N_2717,N_2720);
and U6260 (N_6260,N_3441,N_4480);
and U6261 (N_6261,N_2940,N_2957);
nand U6262 (N_6262,N_4926,N_1235);
nand U6263 (N_6263,N_3228,N_2865);
or U6264 (N_6264,N_2475,N_2524);
or U6265 (N_6265,N_3905,N_2605);
and U6266 (N_6266,N_202,N_178);
nand U6267 (N_6267,N_2568,N_1324);
and U6268 (N_6268,N_4318,N_2733);
nor U6269 (N_6269,N_3615,N_3708);
or U6270 (N_6270,N_3852,N_3559);
xnor U6271 (N_6271,N_4385,N_588);
and U6272 (N_6272,N_3470,N_593);
nand U6273 (N_6273,N_3549,N_1013);
nor U6274 (N_6274,N_4990,N_3886);
or U6275 (N_6275,N_785,N_3759);
nand U6276 (N_6276,N_2254,N_3151);
or U6277 (N_6277,N_660,N_3377);
or U6278 (N_6278,N_3057,N_2083);
nor U6279 (N_6279,N_2079,N_515);
nand U6280 (N_6280,N_1691,N_2304);
or U6281 (N_6281,N_659,N_289);
nand U6282 (N_6282,N_257,N_725);
or U6283 (N_6283,N_3365,N_2986);
or U6284 (N_6284,N_551,N_978);
nor U6285 (N_6285,N_3379,N_3541);
and U6286 (N_6286,N_4446,N_4160);
xor U6287 (N_6287,N_1646,N_4156);
nand U6288 (N_6288,N_1620,N_2215);
nor U6289 (N_6289,N_3823,N_4532);
nor U6290 (N_6290,N_4070,N_4084);
and U6291 (N_6291,N_3362,N_2261);
nor U6292 (N_6292,N_3129,N_1233);
and U6293 (N_6293,N_152,N_2551);
nor U6294 (N_6294,N_729,N_4836);
and U6295 (N_6295,N_2167,N_836);
nand U6296 (N_6296,N_3733,N_2428);
nand U6297 (N_6297,N_4218,N_738);
and U6298 (N_6298,N_2338,N_4234);
nor U6299 (N_6299,N_55,N_8);
nor U6300 (N_6300,N_2043,N_180);
and U6301 (N_6301,N_3935,N_3355);
nand U6302 (N_6302,N_4116,N_1818);
nand U6303 (N_6303,N_4354,N_3885);
and U6304 (N_6304,N_1846,N_241);
or U6305 (N_6305,N_4662,N_813);
or U6306 (N_6306,N_848,N_2168);
or U6307 (N_6307,N_2257,N_4766);
or U6308 (N_6308,N_1931,N_4411);
nand U6309 (N_6309,N_1524,N_2011);
xor U6310 (N_6310,N_2467,N_1469);
or U6311 (N_6311,N_3837,N_2990);
or U6312 (N_6312,N_3695,N_126);
and U6313 (N_6313,N_2050,N_1792);
nor U6314 (N_6314,N_4399,N_222);
nand U6315 (N_6315,N_1463,N_4856);
nand U6316 (N_6316,N_3743,N_561);
or U6317 (N_6317,N_1549,N_1200);
nand U6318 (N_6318,N_2980,N_3421);
nor U6319 (N_6319,N_2334,N_3924);
nand U6320 (N_6320,N_4689,N_1131);
or U6321 (N_6321,N_4892,N_1599);
or U6322 (N_6322,N_4390,N_4095);
nand U6323 (N_6323,N_3025,N_1917);
nand U6324 (N_6324,N_3644,N_4709);
nand U6325 (N_6325,N_4807,N_1773);
and U6326 (N_6326,N_3439,N_4542);
nand U6327 (N_6327,N_1201,N_2433);
xnor U6328 (N_6328,N_3239,N_1015);
nand U6329 (N_6329,N_1511,N_2394);
nand U6330 (N_6330,N_2024,N_3767);
nor U6331 (N_6331,N_4895,N_3701);
nor U6332 (N_6332,N_182,N_185);
and U6333 (N_6333,N_741,N_2871);
or U6334 (N_6334,N_3524,N_1636);
nor U6335 (N_6335,N_3051,N_1925);
and U6336 (N_6336,N_3335,N_2796);
nand U6337 (N_6337,N_1537,N_3795);
or U6338 (N_6338,N_1053,N_3230);
and U6339 (N_6339,N_3163,N_3048);
and U6340 (N_6340,N_2246,N_4568);
nor U6341 (N_6341,N_4764,N_1160);
nand U6342 (N_6342,N_1785,N_4320);
and U6343 (N_6343,N_2586,N_3845);
nand U6344 (N_6344,N_3324,N_4571);
nand U6345 (N_6345,N_2283,N_2100);
nor U6346 (N_6346,N_354,N_3269);
nand U6347 (N_6347,N_4769,N_306);
nand U6348 (N_6348,N_3992,N_2446);
nand U6349 (N_6349,N_989,N_652);
or U6350 (N_6350,N_3153,N_683);
or U6351 (N_6351,N_3444,N_3234);
nand U6352 (N_6352,N_1392,N_767);
or U6353 (N_6353,N_3562,N_2321);
nor U6354 (N_6354,N_3249,N_543);
and U6355 (N_6355,N_908,N_3576);
or U6356 (N_6356,N_3034,N_322);
nor U6357 (N_6357,N_1007,N_384);
and U6358 (N_6358,N_1994,N_656);
or U6359 (N_6359,N_3320,N_821);
and U6360 (N_6360,N_1764,N_3030);
and U6361 (N_6361,N_4455,N_882);
or U6362 (N_6362,N_3442,N_922);
and U6363 (N_6363,N_4066,N_2272);
and U6364 (N_6364,N_1790,N_95);
and U6365 (N_6365,N_2075,N_2603);
or U6366 (N_6366,N_4695,N_325);
and U6367 (N_6367,N_1436,N_4763);
nand U6368 (N_6368,N_1737,N_4284);
or U6369 (N_6369,N_2190,N_2599);
or U6370 (N_6370,N_2210,N_2238);
and U6371 (N_6371,N_865,N_2108);
nand U6372 (N_6372,N_3687,N_3891);
and U6373 (N_6373,N_1778,N_1746);
nand U6374 (N_6374,N_3507,N_924);
or U6375 (N_6375,N_505,N_764);
or U6376 (N_6376,N_2507,N_3556);
or U6377 (N_6377,N_4770,N_1262);
nor U6378 (N_6378,N_930,N_3838);
nor U6379 (N_6379,N_2919,N_3704);
and U6380 (N_6380,N_712,N_3859);
and U6381 (N_6381,N_2205,N_2179);
xor U6382 (N_6382,N_3618,N_4321);
and U6383 (N_6383,N_1415,N_278);
and U6384 (N_6384,N_3095,N_1624);
nand U6385 (N_6385,N_4519,N_4245);
xor U6386 (N_6386,N_35,N_876);
or U6387 (N_6387,N_4575,N_3834);
or U6388 (N_6388,N_3640,N_1189);
and U6389 (N_6389,N_300,N_2653);
or U6390 (N_6390,N_579,N_3508);
nor U6391 (N_6391,N_1305,N_801);
and U6392 (N_6392,N_4816,N_3926);
and U6393 (N_6393,N_1573,N_1495);
nand U6394 (N_6394,N_3073,N_4409);
or U6395 (N_6395,N_4665,N_2566);
nor U6396 (N_6396,N_3853,N_1296);
or U6397 (N_6397,N_2861,N_1974);
and U6398 (N_6398,N_3189,N_3727);
or U6399 (N_6399,N_3205,N_187);
and U6400 (N_6400,N_1941,N_4468);
or U6401 (N_6401,N_431,N_4113);
nor U6402 (N_6402,N_1701,N_2452);
or U6403 (N_6403,N_4128,N_4582);
nor U6404 (N_6404,N_1232,N_2679);
or U6405 (N_6405,N_1330,N_2378);
or U6406 (N_6406,N_3782,N_4692);
nand U6407 (N_6407,N_4619,N_3088);
xor U6408 (N_6408,N_3067,N_3870);
and U6409 (N_6409,N_422,N_1117);
or U6410 (N_6410,N_88,N_2797);
and U6411 (N_6411,N_1726,N_1157);
nand U6412 (N_6412,N_3446,N_223);
and U6413 (N_6413,N_927,N_2785);
nor U6414 (N_6414,N_2649,N_2175);
or U6415 (N_6415,N_2307,N_1183);
xor U6416 (N_6416,N_1697,N_1762);
or U6417 (N_6417,N_2147,N_3553);
xnor U6418 (N_6418,N_4051,N_512);
nor U6419 (N_6419,N_4345,N_3602);
or U6420 (N_6420,N_2975,N_1101);
nor U6421 (N_6421,N_3256,N_3688);
nor U6422 (N_6422,N_4178,N_4853);
or U6423 (N_6423,N_2907,N_183);
nor U6424 (N_6424,N_353,N_4484);
nor U6425 (N_6425,N_1086,N_136);
nor U6426 (N_6426,N_360,N_3597);
or U6427 (N_6427,N_2928,N_3791);
and U6428 (N_6428,N_1666,N_4748);
nand U6429 (N_6429,N_1384,N_2020);
nand U6430 (N_6430,N_4151,N_2538);
and U6431 (N_6431,N_2872,N_1828);
nand U6432 (N_6432,N_2884,N_4079);
nor U6433 (N_6433,N_3430,N_1452);
and U6434 (N_6434,N_1515,N_4436);
nand U6435 (N_6435,N_3396,N_1217);
or U6436 (N_6436,N_3093,N_442);
nor U6437 (N_6437,N_1569,N_2320);
nor U6438 (N_6438,N_1017,N_2571);
and U6439 (N_6439,N_575,N_3489);
nand U6440 (N_6440,N_1179,N_441);
nand U6441 (N_6441,N_1987,N_3732);
or U6442 (N_6442,N_2430,N_2742);
nor U6443 (N_6443,N_3839,N_3579);
or U6444 (N_6444,N_716,N_4846);
nor U6445 (N_6445,N_4242,N_3264);
and U6446 (N_6446,N_952,N_4464);
nand U6447 (N_6447,N_4726,N_3455);
and U6448 (N_6448,N_2589,N_3149);
and U6449 (N_6449,N_3478,N_124);
or U6450 (N_6450,N_985,N_2223);
and U6451 (N_6451,N_4641,N_3918);
or U6452 (N_6452,N_85,N_3670);
nand U6453 (N_6453,N_3794,N_1553);
nor U6454 (N_6454,N_362,N_959);
nor U6455 (N_6455,N_892,N_1546);
or U6456 (N_6456,N_3799,N_4076);
nor U6457 (N_6457,N_1943,N_2625);
nor U6458 (N_6458,N_3860,N_4000);
and U6459 (N_6459,N_1704,N_1602);
and U6460 (N_6460,N_1447,N_2715);
and U6461 (N_6461,N_2809,N_3426);
nand U6462 (N_6462,N_1237,N_3518);
nand U6463 (N_6463,N_4350,N_2969);
or U6464 (N_6464,N_1791,N_3986);
nand U6465 (N_6465,N_3606,N_1042);
nor U6466 (N_6466,N_4014,N_4163);
or U6467 (N_6467,N_3513,N_1419);
nor U6468 (N_6468,N_2013,N_3843);
nand U6469 (N_6469,N_2898,N_1125);
or U6470 (N_6470,N_2866,N_3578);
nor U6471 (N_6471,N_902,N_655);
or U6472 (N_6472,N_915,N_676);
or U6473 (N_6473,N_3424,N_754);
nor U6474 (N_6474,N_2459,N_2732);
nor U6475 (N_6475,N_3024,N_3857);
and U6476 (N_6476,N_988,N_3861);
nor U6477 (N_6477,N_4964,N_1284);
or U6478 (N_6478,N_1109,N_2753);
and U6479 (N_6479,N_1297,N_153);
nor U6480 (N_6480,N_3394,N_3911);
or U6481 (N_6481,N_3226,N_4366);
nor U6482 (N_6482,N_446,N_1223);
or U6483 (N_6483,N_195,N_3872);
xnor U6484 (N_6484,N_576,N_3236);
or U6485 (N_6485,N_434,N_1409);
and U6486 (N_6486,N_3223,N_3907);
and U6487 (N_6487,N_834,N_4305);
nor U6488 (N_6488,N_1977,N_3358);
and U6489 (N_6489,N_2698,N_218);
nor U6490 (N_6490,N_3731,N_804);
and U6491 (N_6491,N_165,N_4854);
and U6492 (N_6492,N_4657,N_1136);
nand U6493 (N_6493,N_3143,N_4801);
nor U6494 (N_6494,N_2541,N_756);
or U6495 (N_6495,N_3066,N_1728);
or U6496 (N_6496,N_2759,N_1811);
or U6497 (N_6497,N_3259,N_4626);
and U6498 (N_6498,N_3641,N_1781);
and U6499 (N_6499,N_1260,N_4901);
nand U6500 (N_6500,N_2811,N_780);
nor U6501 (N_6501,N_3294,N_4592);
nand U6502 (N_6502,N_1513,N_2770);
or U6503 (N_6503,N_563,N_4706);
xnor U6504 (N_6504,N_2431,N_4632);
or U6505 (N_6505,N_3539,N_2329);
nor U6506 (N_6506,N_2293,N_4368);
and U6507 (N_6507,N_3816,N_3898);
or U6508 (N_6508,N_17,N_4647);
nor U6509 (N_6509,N_1218,N_4071);
xnor U6510 (N_6510,N_2890,N_3968);
nand U6511 (N_6511,N_1638,N_4998);
and U6512 (N_6512,N_4860,N_3669);
nand U6513 (N_6513,N_4457,N_3147);
nor U6514 (N_6514,N_2176,N_4012);
or U6515 (N_6515,N_3005,N_2837);
and U6516 (N_6516,N_3714,N_2609);
or U6517 (N_6517,N_743,N_1717);
nor U6518 (N_6518,N_4834,N_2262);
nor U6519 (N_6519,N_3415,N_2673);
and U6520 (N_6520,N_4937,N_3807);
nor U6521 (N_6521,N_1203,N_1091);
and U6522 (N_6522,N_2867,N_3558);
nand U6523 (N_6523,N_2730,N_2808);
nor U6524 (N_6524,N_2754,N_3332);
and U6525 (N_6525,N_3720,N_3800);
and U6526 (N_6526,N_4118,N_4917);
and U6527 (N_6527,N_1215,N_692);
nor U6528 (N_6528,N_497,N_2305);
and U6529 (N_6529,N_4352,N_56);
and U6530 (N_6530,N_2565,N_432);
or U6531 (N_6531,N_641,N_1096);
nand U6532 (N_6532,N_1267,N_3954);
xor U6533 (N_6533,N_631,N_560);
nor U6534 (N_6534,N_3288,N_1309);
nand U6535 (N_6535,N_4140,N_111);
or U6536 (N_6536,N_3181,N_3988);
nand U6537 (N_6537,N_1863,N_2810);
nand U6538 (N_6538,N_2545,N_1457);
nor U6539 (N_6539,N_4879,N_3952);
nor U6540 (N_6540,N_3894,N_1389);
nor U6541 (N_6541,N_2234,N_3908);
nor U6542 (N_6542,N_234,N_4633);
or U6543 (N_6543,N_1085,N_2456);
nor U6544 (N_6544,N_3979,N_4978);
or U6545 (N_6545,N_343,N_514);
and U6546 (N_6546,N_1625,N_1018);
nand U6547 (N_6547,N_3027,N_194);
or U6548 (N_6548,N_2447,N_61);
nor U6549 (N_6549,N_3477,N_1642);
nand U6550 (N_6550,N_3014,N_2781);
nand U6551 (N_6551,N_386,N_4861);
and U6552 (N_6552,N_2520,N_4319);
nand U6553 (N_6553,N_4612,N_3832);
nand U6554 (N_6554,N_4811,N_4378);
or U6555 (N_6555,N_2774,N_2151);
xor U6556 (N_6556,N_484,N_3546);
or U6557 (N_6557,N_3401,N_1767);
or U6558 (N_6558,N_510,N_2600);
and U6559 (N_6559,N_2556,N_680);
nand U6560 (N_6560,N_3552,N_3786);
nand U6561 (N_6561,N_2082,N_3210);
nand U6562 (N_6562,N_1490,N_1687);
nand U6563 (N_6563,N_1417,N_552);
and U6564 (N_6564,N_1604,N_975);
nor U6565 (N_6565,N_83,N_3621);
nand U6566 (N_6566,N_64,N_3771);
nand U6567 (N_6567,N_3304,N_4384);
nor U6568 (N_6568,N_4920,N_2935);
and U6569 (N_6569,N_4598,N_3580);
nor U6570 (N_6570,N_4027,N_140);
and U6571 (N_6571,N_4026,N_4360);
or U6572 (N_6572,N_3237,N_4170);
or U6573 (N_6573,N_3029,N_4454);
and U6574 (N_6574,N_4491,N_3637);
nor U6575 (N_6575,N_4504,N_3445);
xnor U6576 (N_6576,N_2794,N_2385);
xnor U6577 (N_6577,N_4259,N_4299);
and U6578 (N_6578,N_3363,N_2974);
nor U6579 (N_6579,N_4077,N_1071);
and U6580 (N_6580,N_1357,N_2117);
nand U6581 (N_6581,N_4459,N_2380);
nor U6582 (N_6582,N_3156,N_1552);
or U6583 (N_6583,N_71,N_2993);
nand U6584 (N_6584,N_2812,N_3043);
nor U6585 (N_6585,N_868,N_4973);
nand U6586 (N_6586,N_2186,N_844);
nor U6587 (N_6587,N_1786,N_19);
xor U6588 (N_6588,N_2864,N_151);
or U6589 (N_6589,N_2495,N_4835);
or U6590 (N_6590,N_1133,N_2683);
and U6591 (N_6591,N_2458,N_954);
or U6592 (N_6592,N_4201,N_1052);
xor U6593 (N_6593,N_4293,N_914);
nor U6594 (N_6594,N_1029,N_662);
nand U6595 (N_6595,N_925,N_1360);
or U6596 (N_6596,N_3013,N_2093);
nand U6597 (N_6597,N_82,N_2815);
nand U6598 (N_6598,N_2516,N_1195);
nor U6599 (N_6599,N_3428,N_2553);
nand U6600 (N_6600,N_145,N_998);
or U6601 (N_6601,N_1659,N_3673);
and U6602 (N_6602,N_2912,N_1167);
and U6603 (N_6603,N_687,N_1742);
nor U6604 (N_6604,N_3340,N_503);
or U6605 (N_6605,N_2708,N_2626);
nand U6606 (N_6606,N_44,N_258);
nand U6607 (N_6607,N_3548,N_4997);
nand U6608 (N_6608,N_2104,N_4557);
nand U6609 (N_6609,N_634,N_4697);
nand U6610 (N_6610,N_2576,N_2745);
nand U6611 (N_6611,N_2474,N_1476);
xnor U6612 (N_6612,N_1843,N_1026);
or U6613 (N_6613,N_2789,N_3761);
nand U6614 (N_6614,N_1772,N_3709);
and U6615 (N_6615,N_2878,N_1407);
and U6616 (N_6616,N_4543,N_1249);
nand U6617 (N_6617,N_4493,N_4235);
and U6618 (N_6618,N_2370,N_2704);
and U6619 (N_6619,N_27,N_4036);
or U6620 (N_6620,N_4276,N_1298);
and U6621 (N_6621,N_2608,N_1654);
nor U6622 (N_6622,N_1001,N_4831);
or U6623 (N_6623,N_699,N_4434);
and U6624 (N_6624,N_2145,N_3105);
and U6625 (N_6625,N_4015,N_2406);
nor U6626 (N_6626,N_3460,N_2807);
and U6627 (N_6627,N_3724,N_3356);
nand U6628 (N_6628,N_1961,N_157);
nor U6629 (N_6629,N_2267,N_1187);
nand U6630 (N_6630,N_817,N_2909);
and U6631 (N_6631,N_2788,N_2200);
nand U6632 (N_6632,N_118,N_1481);
nor U6633 (N_6633,N_828,N_4564);
or U6634 (N_6634,N_2709,N_3260);
xor U6635 (N_6635,N_827,N_1571);
nor U6636 (N_6636,N_3214,N_1819);
or U6637 (N_6637,N_2434,N_3164);
or U6638 (N_6638,N_912,N_869);
or U6639 (N_6639,N_3497,N_1473);
nand U6640 (N_6640,N_3443,N_3391);
nor U6641 (N_6641,N_3121,N_4256);
and U6642 (N_6642,N_1306,N_2955);
nor U6643 (N_6643,N_3019,N_4460);
or U6644 (N_6644,N_4024,N_78);
nor U6645 (N_6645,N_4477,N_557);
nor U6646 (N_6646,N_758,N_4868);
nor U6647 (N_6647,N_608,N_3892);
and U6648 (N_6648,N_4960,N_2863);
or U6649 (N_6649,N_4061,N_513);
or U6650 (N_6650,N_2069,N_3432);
and U6651 (N_6651,N_4832,N_2182);
or U6652 (N_6652,N_2290,N_1247);
or U6653 (N_6653,N_400,N_4375);
nor U6654 (N_6654,N_2642,N_1851);
nand U6655 (N_6655,N_1559,N_1451);
or U6656 (N_6656,N_4428,N_3168);
nand U6657 (N_6657,N_1993,N_388);
or U6658 (N_6658,N_2971,N_531);
nand U6659 (N_6659,N_1641,N_2092);
xor U6660 (N_6660,N_4736,N_2006);
nor U6661 (N_6661,N_1354,N_1739);
nor U6662 (N_6662,N_1578,N_29);
nor U6663 (N_6663,N_860,N_1873);
nand U6664 (N_6664,N_2076,N_4238);
and U6665 (N_6665,N_4750,N_2827);
nor U6666 (N_6666,N_3037,N_2604);
nand U6667 (N_6667,N_274,N_977);
or U6668 (N_6668,N_4316,N_1595);
or U6669 (N_6669,N_4295,N_1367);
nand U6670 (N_6670,N_2470,N_2896);
nor U6671 (N_6671,N_769,N_2567);
or U6672 (N_6672,N_4058,N_3179);
and U6673 (N_6673,N_4634,N_3169);
and U6674 (N_6674,N_2353,N_3994);
or U6675 (N_6675,N_3117,N_3527);
nand U6676 (N_6676,N_87,N_3495);
or U6677 (N_6677,N_2241,N_204);
or U6678 (N_6678,N_502,N_4989);
nor U6679 (N_6679,N_1353,N_1197);
nand U6680 (N_6680,N_231,N_1727);
nor U6681 (N_6681,N_2216,N_4285);
and U6682 (N_6682,N_894,N_443);
or U6683 (N_6683,N_3649,N_2663);
and U6684 (N_6684,N_1771,N_4476);
and U6685 (N_6685,N_1775,N_1816);
nor U6686 (N_6686,N_1368,N_331);
nor U6687 (N_6687,N_4735,N_3059);
nor U6688 (N_6688,N_832,N_4380);
nand U6689 (N_6689,N_2970,N_3878);
nand U6690 (N_6690,N_291,N_378);
or U6691 (N_6691,N_2721,N_2268);
nand U6692 (N_6692,N_4008,N_2515);
and U6693 (N_6693,N_4640,N_3718);
and U6694 (N_6694,N_2478,N_3776);
xor U6695 (N_6695,N_1478,N_4566);
nor U6696 (N_6696,N_2744,N_93);
nor U6697 (N_6697,N_2905,N_3712);
nand U6698 (N_6698,N_3946,N_763);
or U6699 (N_6699,N_4967,N_3785);
and U6700 (N_6700,N_837,N_2741);
nor U6701 (N_6701,N_690,N_1658);
nand U6702 (N_6702,N_1888,N_2005);
nand U6703 (N_6703,N_916,N_4057);
nand U6704 (N_6704,N_4165,N_3089);
nor U6705 (N_6705,N_2161,N_1936);
nand U6706 (N_6706,N_3721,N_3303);
nand U6707 (N_6707,N_700,N_4159);
nor U6708 (N_6708,N_1405,N_4623);
nand U6709 (N_6709,N_2404,N_4993);
or U6710 (N_6710,N_4671,N_1317);
and U6711 (N_6711,N_2097,N_4878);
or U6712 (N_6712,N_401,N_4373);
nor U6713 (N_6713,N_4332,N_1836);
nand U6714 (N_6714,N_1940,N_229);
nand U6715 (N_6715,N_3547,N_4629);
and U6716 (N_6716,N_2658,N_1236);
nor U6717 (N_6717,N_1020,N_4147);
and U6718 (N_6718,N_4870,N_4761);
or U6719 (N_6719,N_4381,N_3216);
nand U6720 (N_6720,N_4419,N_4533);
nor U6721 (N_6721,N_3811,N_1803);
nor U6722 (N_6722,N_2614,N_3707);
nor U6723 (N_6723,N_3277,N_815);
or U6724 (N_6724,N_1475,N_3273);
nor U6725 (N_6725,N_1592,N_1577);
or U6726 (N_6726,N_1355,N_594);
or U6727 (N_6727,N_3658,N_2233);
and U6728 (N_6728,N_3031,N_3725);
and U6729 (N_6729,N_4809,N_4089);
nand U6730 (N_6730,N_4620,N_3980);
and U6731 (N_6731,N_4440,N_3436);
nor U6732 (N_6732,N_249,N_2130);
nor U6733 (N_6733,N_4421,N_2258);
or U6734 (N_6734,N_3756,N_1230);
or U6735 (N_6735,N_2172,N_314);
and U6736 (N_6736,N_1684,N_493);
or U6737 (N_6737,N_4906,N_408);
nand U6738 (N_6738,N_2723,N_321);
nand U6739 (N_6739,N_3830,N_872);
nand U6740 (N_6740,N_2800,N_143);
nor U6741 (N_6741,N_2072,N_4386);
and U6742 (N_6742,N_196,N_1159);
and U6743 (N_6743,N_1765,N_4291);
or U6744 (N_6744,N_4388,N_483);
or U6745 (N_6745,N_1509,N_4341);
and U6746 (N_6746,N_4752,N_1738);
or U6747 (N_6747,N_299,N_3625);
or U6748 (N_6748,N_1912,N_4822);
and U6749 (N_6749,N_2778,N_2743);
or U6750 (N_6750,N_849,N_452);
or U6751 (N_6751,N_2540,N_1025);
or U6752 (N_6752,N_2358,N_1734);
nand U6753 (N_6753,N_2124,N_3521);
nor U6754 (N_6754,N_4751,N_808);
and U6755 (N_6755,N_3937,N_1971);
or U6756 (N_6756,N_3213,N_2232);
and U6757 (N_6757,N_4653,N_2664);
nor U6758 (N_6758,N_4110,N_1148);
nand U6759 (N_6759,N_4741,N_1084);
and U6760 (N_6760,N_1060,N_310);
or U6761 (N_6761,N_4470,N_1856);
nand U6762 (N_6762,N_948,N_2580);
nand U6763 (N_6763,N_4494,N_433);
and U6764 (N_6764,N_4322,N_4771);
nor U6765 (N_6765,N_3505,N_1143);
nand U6766 (N_6766,N_3689,N_3152);
and U6767 (N_6767,N_1613,N_1899);
nand U6768 (N_6768,N_495,N_3656);
nor U6769 (N_6769,N_162,N_684);
nand U6770 (N_6770,N_2078,N_1358);
nand U6771 (N_6771,N_23,N_3418);
nor U6772 (N_6772,N_936,N_3523);
or U6773 (N_6773,N_411,N_3306);
nand U6774 (N_6774,N_1832,N_2106);
nand U6775 (N_6775,N_4789,N_3533);
and U6776 (N_6776,N_3199,N_4975);
nor U6777 (N_6777,N_1582,N_803);
nor U6778 (N_6778,N_4028,N_973);
xor U6779 (N_6779,N_3936,N_3381);
and U6780 (N_6780,N_4772,N_4552);
nor U6781 (N_6781,N_4679,N_1499);
and U6782 (N_6782,N_4475,N_3387);
nand U6783 (N_6783,N_2734,N_993);
nor U6784 (N_6784,N_176,N_1813);
and U6785 (N_6785,N_3282,N_1126);
nor U6786 (N_6786,N_1186,N_4563);
xnor U6787 (N_6787,N_4237,N_2786);
nand U6788 (N_6788,N_4453,N_4765);
and U6789 (N_6789,N_287,N_1723);
nand U6790 (N_6790,N_4055,N_2417);
or U6791 (N_6791,N_2678,N_3755);
nand U6792 (N_6792,N_4415,N_4174);
nor U6793 (N_6793,N_1982,N_146);
and U6794 (N_6794,N_2266,N_4120);
and U6795 (N_6795,N_4217,N_1316);
and U6796 (N_6796,N_4733,N_4306);
and U6797 (N_6797,N_4526,N_2561);
and U6798 (N_6798,N_1824,N_2316);
and U6799 (N_6799,N_4734,N_3086);
nand U6800 (N_6800,N_4759,N_2981);
or U6801 (N_6801,N_4330,N_1935);
and U6802 (N_6802,N_3512,N_2494);
nor U6803 (N_6803,N_478,N_4043);
nor U6804 (N_6804,N_602,N_4932);
or U6805 (N_6805,N_4497,N_616);
nor U6806 (N_6806,N_4914,N_3928);
and U6807 (N_6807,N_744,N_698);
or U6808 (N_6808,N_2095,N_286);
nor U6809 (N_6809,N_4134,N_4262);
nor U6810 (N_6810,N_4864,N_1694);
and U6811 (N_6811,N_1434,N_2682);
and U6812 (N_6812,N_1301,N_4365);
nand U6813 (N_6813,N_1418,N_1674);
nor U6814 (N_6814,N_3819,N_267);
nor U6815 (N_6815,N_2752,N_3021);
and U6816 (N_6816,N_2386,N_3588);
nand U6817 (N_6817,N_1051,N_3573);
nor U6818 (N_6818,N_4141,N_1541);
nor U6819 (N_6819,N_2631,N_4393);
and U6820 (N_6820,N_4893,N_1124);
or U6821 (N_6821,N_2607,N_1518);
nor U6822 (N_6822,N_1713,N_3471);
nor U6823 (N_6823,N_4556,N_1413);
nand U6824 (N_6824,N_3818,N_816);
and U6825 (N_6825,N_399,N_2255);
and U6826 (N_6826,N_569,N_2674);
nor U6827 (N_6827,N_1698,N_4424);
or U6828 (N_6828,N_2000,N_981);
and U6829 (N_6829,N_520,N_4107);
or U6830 (N_6830,N_2950,N_4175);
nand U6831 (N_6831,N_1591,N_2306);
nand U6832 (N_6832,N_426,N_67);
nand U6833 (N_6833,N_3804,N_1998);
nor U6834 (N_6834,N_2038,N_1902);
nand U6835 (N_6835,N_4537,N_3407);
nor U6836 (N_6836,N_762,N_3245);
nor U6837 (N_6837,N_421,N_1343);
nand U6838 (N_6838,N_2519,N_1530);
nand U6839 (N_6839,N_1615,N_4900);
nor U6840 (N_6840,N_2222,N_4876);
nand U6841 (N_6841,N_565,N_2885);
or U6842 (N_6842,N_3890,N_2585);
and U6843 (N_6843,N_1016,N_3608);
or U6844 (N_6844,N_315,N_80);
and U6845 (N_6845,N_751,N_4792);
or U6846 (N_6846,N_3745,N_4681);
nor U6847 (N_6847,N_1315,N_486);
and U6848 (N_6848,N_898,N_2454);
nand U6849 (N_6849,N_2936,N_1194);
nor U6850 (N_6850,N_722,N_3091);
nand U6851 (N_6851,N_2846,N_907);
or U6852 (N_6852,N_4042,N_2476);
nor U6853 (N_6853,N_4738,N_2299);
nand U6854 (N_6854,N_2156,N_4743);
and U6855 (N_6855,N_4714,N_3586);
or U6856 (N_6856,N_3824,N_4829);
nand U6857 (N_6857,N_3481,N_1725);
or U6858 (N_6858,N_1190,N_2654);
and U6859 (N_6859,N_4782,N_2636);
nor U6860 (N_6860,N_1920,N_3232);
nand U6861 (N_6861,N_2806,N_534);
and U6862 (N_6862,N_4559,N_4551);
and U6863 (N_6863,N_625,N_4600);
nor U6864 (N_6864,N_3717,N_4511);
nand U6865 (N_6865,N_3326,N_2783);
and U6866 (N_6866,N_3913,N_3877);
nand U6867 (N_6867,N_2591,N_2959);
or U6868 (N_6868,N_776,N_348);
nor U6869 (N_6869,N_253,N_2460);
nor U6870 (N_6870,N_3018,N_2620);
xnor U6871 (N_6871,N_1821,N_2323);
nor U6872 (N_6872,N_4930,N_3343);
nor U6873 (N_6873,N_3078,N_2127);
nand U6874 (N_6874,N_1144,N_928);
nand U6875 (N_6875,N_523,N_1809);
or U6876 (N_6876,N_1366,N_737);
nor U6877 (N_6877,N_4346,N_2582);
or U6878 (N_6878,N_355,N_2416);
and U6879 (N_6879,N_2420,N_4654);
or U6880 (N_6880,N_682,N_1161);
and U6881 (N_6881,N_167,N_4418);
nand U6882 (N_6882,N_2480,N_4693);
nor U6883 (N_6883,N_696,N_4848);
or U6884 (N_6884,N_1062,N_2874);
xnor U6885 (N_6885,N_3373,N_3611);
or U6886 (N_6886,N_1558,N_2526);
and U6887 (N_6887,N_397,N_1454);
and U6888 (N_6888,N_1428,N_1696);
and U6889 (N_6889,N_3184,N_1503);
and U6890 (N_6890,N_778,N_2622);
or U6891 (N_6891,N_1745,N_250);
nor U6892 (N_6892,N_4249,N_3092);
xnor U6893 (N_6893,N_460,N_4290);
and U6894 (N_6894,N_970,N_4655);
nand U6895 (N_6895,N_2922,N_3359);
nand U6896 (N_6896,N_2203,N_2153);
or U6897 (N_6897,N_3203,N_3077);
or U6898 (N_6898,N_1736,N_284);
nor U6899 (N_6899,N_1980,N_3263);
xnor U6900 (N_6900,N_4205,N_3404);
nand U6901 (N_6901,N_1340,N_3752);
or U6902 (N_6902,N_589,N_2189);
nand U6903 (N_6903,N_1946,N_2437);
and U6904 (N_6904,N_2439,N_450);
xor U6905 (N_6905,N_4712,N_718);
nand U6906 (N_6906,N_4524,N_1932);
xnor U6907 (N_6907,N_3592,N_4558);
nor U6908 (N_6908,N_4677,N_4252);
and U6909 (N_6909,N_3594,N_2365);
nor U6910 (N_6910,N_1290,N_4615);
and U6911 (N_6911,N_2869,N_4244);
or U6912 (N_6912,N_2793,N_369);
nand U6913 (N_6913,N_4988,N_3683);
and U6914 (N_6914,N_1248,N_366);
or U6915 (N_6915,N_462,N_4078);
nand U6916 (N_6916,N_2204,N_155);
and U6917 (N_6917,N_665,N_3912);
or U6918 (N_6918,N_1245,N_3540);
or U6919 (N_6919,N_1445,N_1280);
nor U6920 (N_6920,N_4686,N_1647);
and U6921 (N_6921,N_181,N_3409);
or U6922 (N_6922,N_4680,N_2120);
and U6923 (N_6923,N_3899,N_4148);
nand U6924 (N_6924,N_1438,N_4587);
or U6925 (N_6925,N_4757,N_585);
nand U6926 (N_6926,N_900,N_2419);
nand U6927 (N_6927,N_2689,N_4270);
or U6928 (N_6928,N_4985,N_3437);
nand U6929 (N_6929,N_707,N_2146);
nor U6930 (N_6930,N_4229,N_1880);
nor U6931 (N_6931,N_2325,N_3261);
and U6932 (N_6932,N_2118,N_1838);
nand U6933 (N_6933,N_1257,N_4344);
nand U6934 (N_6934,N_1066,N_4022);
nor U6935 (N_6935,N_213,N_1959);
xnor U6936 (N_6936,N_1376,N_2954);
nor U6937 (N_6937,N_4473,N_943);
and U6938 (N_6938,N_1951,N_4294);
or U6939 (N_6939,N_2531,N_2554);
and U6940 (N_6940,N_2356,N_4908);
nor U6941 (N_6941,N_1756,N_2);
nor U6942 (N_6942,N_3138,N_292);
nor U6943 (N_6943,N_3225,N_4215);
or U6944 (N_6944,N_3336,N_1012);
nor U6945 (N_6945,N_4548,N_3951);
and U6946 (N_6946,N_449,N_3677);
and U6947 (N_6947,N_4427,N_2537);
nor U6948 (N_6948,N_4966,N_4904);
nand U6949 (N_6949,N_2862,N_4590);
or U6950 (N_6950,N_62,N_2502);
or U6951 (N_6951,N_488,N_720);
nand U6952 (N_6952,N_3406,N_1268);
and U6953 (N_6953,N_15,N_4068);
or U6954 (N_6954,N_2471,N_1335);
nor U6955 (N_6955,N_2218,N_1156);
or U6956 (N_6956,N_3465,N_4956);
nor U6957 (N_6957,N_2455,N_2873);
or U6958 (N_6958,N_2941,N_4056);
and U6959 (N_6959,N_4465,N_4025);
or U6960 (N_6960,N_2903,N_3281);
nor U6961 (N_6961,N_4053,N_4718);
nor U6962 (N_6962,N_4251,N_1000);
nand U6963 (N_6963,N_1341,N_3374);
nor U6964 (N_6964,N_3792,N_745);
nor U6965 (N_6965,N_4925,N_1333);
nand U6966 (N_6966,N_161,N_3567);
or U6967 (N_6967,N_4367,N_2485);
and U6968 (N_6968,N_783,N_793);
and U6969 (N_6969,N_3915,N_4083);
or U6970 (N_6970,N_3383,N_3880);
or U6971 (N_6971,N_857,N_3267);
or U6972 (N_6972,N_2751,N_1618);
nor U6973 (N_6973,N_2597,N_824);
nor U6974 (N_6974,N_1841,N_4923);
or U6975 (N_6975,N_1050,N_4173);
nor U6976 (N_6976,N_3766,N_4257);
or U6977 (N_6977,N_3953,N_1639);
nand U6978 (N_6978,N_477,N_359);
nand U6979 (N_6979,N_3599,N_1404);
nor U6980 (N_6980,N_590,N_2817);
nand U6981 (N_6981,N_1220,N_4422);
and U6982 (N_6982,N_1178,N_2841);
nor U6983 (N_6983,N_2064,N_1342);
and U6984 (N_6984,N_3176,N_1754);
and U6985 (N_6985,N_2158,N_2070);
and U6986 (N_6986,N_1139,N_4898);
nor U6987 (N_6987,N_4963,N_1670);
or U6988 (N_6988,N_4955,N_1645);
nor U6989 (N_6989,N_4034,N_3706);
nand U6990 (N_6990,N_3200,N_26);
or U6991 (N_6991,N_4635,N_1281);
nand U6992 (N_6992,N_4818,N_1561);
nor U6993 (N_6993,N_1318,N_4847);
nand U6994 (N_6994,N_3159,N_404);
nor U6995 (N_6995,N_1644,N_4827);
or U6996 (N_6996,N_1924,N_4400);
and U6997 (N_6997,N_113,N_4030);
nor U6998 (N_6998,N_4687,N_4716);
or U6999 (N_6999,N_4682,N_2148);
nand U7000 (N_7000,N_1519,N_4905);
and U7001 (N_7001,N_2761,N_4123);
and U7002 (N_7002,N_3726,N_4007);
and U7003 (N_7003,N_1275,N_3840);
nand U7004 (N_7004,N_2422,N_2196);
and U7005 (N_7005,N_2402,N_4740);
nor U7006 (N_7006,N_3422,N_3945);
and U7007 (N_7007,N_4797,N_4331);
or U7008 (N_7008,N_2762,N_4439);
nand U7009 (N_7009,N_3820,N_3154);
or U7010 (N_7010,N_3385,N_788);
nor U7011 (N_7011,N_1080,N_403);
and U7012 (N_7012,N_2202,N_3334);
and U7013 (N_7013,N_4065,N_2739);
nor U7014 (N_7014,N_982,N_4149);
and U7015 (N_7015,N_1911,N_13);
xor U7016 (N_7016,N_3957,N_1685);
nor U7017 (N_7017,N_4267,N_3120);
and U7018 (N_7018,N_3702,N_1626);
or U7019 (N_7019,N_3291,N_2575);
and U7020 (N_7020,N_4758,N_881);
nand U7021 (N_7021,N_4721,N_4020);
or U7022 (N_7022,N_3989,N_1352);
and U7023 (N_7023,N_3414,N_4591);
xnor U7024 (N_7024,N_583,N_605);
nand U7025 (N_7025,N_1630,N_2010);
or U7026 (N_7026,N_3050,N_190);
or U7027 (N_7027,N_4430,N_794);
and U7028 (N_7028,N_4553,N_2440);
or U7029 (N_7029,N_2350,N_3331);
nor U7030 (N_7030,N_918,N_730);
and U7031 (N_7031,N_3435,N_1209);
and U7032 (N_7032,N_4817,N_1293);
or U7033 (N_7033,N_2508,N_3116);
and U7034 (N_7034,N_2728,N_3376);
and U7035 (N_7035,N_581,N_3204);
nor U7036 (N_7036,N_2518,N_260);
nor U7037 (N_7037,N_4222,N_556);
or U7038 (N_7038,N_1867,N_28);
or U7039 (N_7039,N_121,N_4576);
nand U7040 (N_7040,N_3662,N_3238);
and U7041 (N_7041,N_79,N_226);
xor U7042 (N_7042,N_4610,N_3466);
and U7043 (N_7043,N_3787,N_2677);
and U7044 (N_7044,N_376,N_3534);
nor U7045 (N_7045,N_45,N_1024);
nand U7046 (N_7046,N_1664,N_271);
xor U7047 (N_7047,N_4206,N_1596);
nor U7048 (N_7048,N_311,N_4292);
or U7049 (N_7049,N_3427,N_2996);
nand U7050 (N_7050,N_2033,N_2214);
nand U7051 (N_7051,N_4263,N_2121);
or U7052 (N_7052,N_2309,N_1928);
or U7053 (N_7053,N_2988,N_1044);
nand U7054 (N_7054,N_3292,N_1548);
or U7055 (N_7055,N_3789,N_4730);
and U7056 (N_7056,N_4746,N_1263);
nand U7057 (N_7057,N_230,N_2221);
or U7058 (N_7058,N_1008,N_2377);
nor U7059 (N_7059,N_2348,N_1311);
and U7060 (N_7060,N_380,N_1345);
or U7061 (N_7061,N_4136,N_391);
nand U7062 (N_7062,N_389,N_4911);
and U7063 (N_7063,N_1802,N_2930);
nand U7064 (N_7064,N_211,N_4648);
or U7065 (N_7065,N_4646,N_2826);
nor U7066 (N_7066,N_810,N_3254);
and U7067 (N_7067,N_1953,N_2023);
nor U7068 (N_7068,N_212,N_2388);
nand U7069 (N_7069,N_1675,N_347);
and U7070 (N_7070,N_77,N_4702);
nor U7071 (N_7071,N_4414,N_2875);
and U7072 (N_7072,N_4842,N_4636);
or U7073 (N_7073,N_3964,N_2333);
nor U7074 (N_7074,N_2389,N_3472);
or U7075 (N_7075,N_890,N_2923);
and U7076 (N_7076,N_4467,N_4936);
nand U7077 (N_7077,N_501,N_2298);
nand U7078 (N_7078,N_1805,N_1680);
or U7079 (N_7079,N_859,N_425);
nor U7080 (N_7080,N_2112,N_2964);
or U7081 (N_7081,N_132,N_4503);
nand U7082 (N_7082,N_1650,N_2617);
or U7083 (N_7083,N_2479,N_455);
nand U7084 (N_7084,N_3682,N_4762);
and U7085 (N_7085,N_829,N_468);
nand U7086 (N_7086,N_3192,N_254);
nand U7087 (N_7087,N_3133,N_4202);
or U7088 (N_7088,N_4486,N_2482);
or U7089 (N_7089,N_1373,N_4664);
or U7090 (N_7090,N_21,N_2756);
and U7091 (N_7091,N_2026,N_379);
xnor U7092 (N_7092,N_1722,N_437);
nor U7093 (N_7093,N_3257,N_3849);
or U7094 (N_7094,N_2638,N_1897);
nor U7095 (N_7095,N_1402,N_3522);
nor U7096 (N_7096,N_3902,N_774);
nor U7097 (N_7097,N_3583,N_2071);
nand U7098 (N_7098,N_3000,N_1467);
nand U7099 (N_7099,N_3463,N_4991);
nand U7100 (N_7100,N_3483,N_4200);
nand U7101 (N_7101,N_1130,N_2269);
or U7102 (N_7102,N_3280,N_838);
nand U7103 (N_7103,N_880,N_4589);
nand U7104 (N_7104,N_3570,N_4398);
xnor U7105 (N_7105,N_2904,N_2945);
nor U7106 (N_7106,N_94,N_2997);
and U7107 (N_7107,N_2632,N_530);
or U7108 (N_7108,N_2525,N_4728);
and U7109 (N_7109,N_3634,N_248);
nand U7110 (N_7110,N_4586,N_1250);
nor U7111 (N_7111,N_3308,N_855);
nor U7112 (N_7112,N_2619,N_578);
or U7113 (N_7113,N_4246,N_282);
or U7114 (N_7114,N_457,N_2629);
nand U7115 (N_7115,N_4037,N_1512);
or U7116 (N_7116,N_4810,N_2832);
xor U7117 (N_7117,N_448,N_100);
xor U7118 (N_7118,N_2877,N_393);
and U7119 (N_7119,N_3977,N_3623);
or U7120 (N_7120,N_4124,N_2838);
nor U7121 (N_7121,N_2150,N_1760);
and U7122 (N_7122,N_601,N_1470);
or U7123 (N_7123,N_4880,N_2059);
and U7124 (N_7124,N_678,N_2171);
nor U7125 (N_7125,N_2648,N_1351);
or U7126 (N_7126,N_2244,N_4186);
xor U7127 (N_7127,N_1870,N_122);
nand U7128 (N_7128,N_4785,N_2081);
or U7129 (N_7129,N_3603,N_2442);
or U7130 (N_7130,N_969,N_4423);
nor U7131 (N_7131,N_884,N_1589);
nor U7132 (N_7132,N_2193,N_1429);
and U7133 (N_7133,N_1471,N_3511);
or U7134 (N_7134,N_3431,N_1871);
and U7135 (N_7135,N_932,N_2427);
nand U7136 (N_7136,N_517,N_1567);
and U7137 (N_7137,N_2314,N_1240);
and U7138 (N_7138,N_429,N_1110);
and U7139 (N_7139,N_796,N_962);
nand U7140 (N_7140,N_1349,N_59);
nand U7141 (N_7141,N_2084,N_2530);
and U7142 (N_7142,N_2445,N_1229);
and U7143 (N_7143,N_609,N_116);
nand U7144 (N_7144,N_3981,N_2652);
nor U7145 (N_7145,N_1923,N_160);
or U7146 (N_7146,N_2814,N_1960);
nor U7147 (N_7147,N_1228,N_805);
nor U7148 (N_7148,N_2684,N_76);
nand U7149 (N_7149,N_3983,N_4574);
nor U7150 (N_7150,N_1565,N_1116);
nor U7151 (N_7151,N_2444,N_2352);
and U7152 (N_7152,N_4814,N_3582);
nor U7153 (N_7153,N_3738,N_1294);
nor U7154 (N_7154,N_275,N_899);
and U7155 (N_7155,N_4804,N_2628);
or U7156 (N_7156,N_4265,N_4841);
nand U7157 (N_7157,N_3664,N_2987);
or U7158 (N_7158,N_1988,N_1279);
and U7159 (N_7159,N_4916,N_1141);
xor U7160 (N_7160,N_1817,N_558);
nor U7161 (N_7161,N_1750,N_2346);
nand U7162 (N_7162,N_861,N_4129);
nand U7163 (N_7163,N_2529,N_438);
nand U7164 (N_7164,N_689,N_4957);
nand U7165 (N_7165,N_4672,N_70);
nand U7166 (N_7166,N_746,N_1286);
and U7167 (N_7167,N_3999,N_2123);
and U7168 (N_7168,N_3814,N_4719);
or U7169 (N_7169,N_2469,N_1344);
and U7170 (N_7170,N_276,N_3809);
and U7171 (N_7171,N_2169,N_1272);
or U7172 (N_7172,N_3053,N_3900);
and U7173 (N_7173,N_1087,N_5);
or U7174 (N_7174,N_1804,N_469);
nand U7175 (N_7175,N_3229,N_4351);
and U7176 (N_7176,N_3920,N_1747);
and U7177 (N_7177,N_320,N_843);
and U7178 (N_7178,N_1196,N_1401);
and U7179 (N_7179,N_4698,N_3605);
or U7180 (N_7180,N_3167,N_2802);
nor U7181 (N_7181,N_1234,N_4866);
and U7182 (N_7182,N_1758,N_3741);
and U7183 (N_7183,N_2462,N_2463);
nor U7184 (N_7184,N_840,N_939);
nand U7185 (N_7185,N_3887,N_3110);
or U7186 (N_7186,N_4584,N_4918);
nor U7187 (N_7187,N_2411,N_4833);
or U7188 (N_7188,N_4005,N_2412);
and U7189 (N_7189,N_4317,N_3193);
nand U7190 (N_7190,N_3423,N_1362);
or U7191 (N_7191,N_2847,N_1886);
nand U7192 (N_7192,N_1814,N_2354);
and U7193 (N_7193,N_4950,N_3686);
and U7194 (N_7194,N_3506,N_4506);
nand U7195 (N_7195,N_2880,N_4638);
or U7196 (N_7196,N_1907,N_4456);
or U7197 (N_7197,N_4705,N_4461);
nand U7198 (N_7198,N_2549,N_1394);
and U7199 (N_7199,N_3155,N_1);
nand U7200 (N_7200,N_2857,N_4996);
or U7201 (N_7201,N_1690,N_1172);
xor U7202 (N_7202,N_2259,N_806);
and U7203 (N_7203,N_1364,N_4288);
nor U7204 (N_7204,N_940,N_905);
nand U7205 (N_7205,N_2659,N_527);
or U7206 (N_7206,N_2451,N_2384);
or U7207 (N_7207,N_733,N_1842);
and U7208 (N_7208,N_2727,N_784);
nor U7209 (N_7209,N_1574,N_4683);
nor U7210 (N_7210,N_2291,N_1834);
nor U7211 (N_7211,N_2570,N_4813);
and U7212 (N_7212,N_4643,N_1455);
and U7213 (N_7213,N_2876,N_91);
or U7214 (N_7214,N_852,N_2573);
nor U7215 (N_7215,N_269,N_4965);
or U7216 (N_7216,N_3509,N_4715);
xor U7217 (N_7217,N_2425,N_3769);
or U7218 (N_7218,N_3454,N_2285);
nand U7219 (N_7219,N_2177,N_313);
or U7220 (N_7220,N_1919,N_2656);
and U7221 (N_7221,N_3923,N_1970);
and U7222 (N_7222,N_2073,N_4933);
or U7223 (N_7223,N_4839,N_1350);
or U7224 (N_7224,N_942,N_3703);
nand U7225 (N_7225,N_752,N_524);
or U7226 (N_7226,N_4628,N_3584);
nor U7227 (N_7227,N_1099,N_4435);
nor U7228 (N_7228,N_2766,N_4786);
and U7229 (N_7229,N_1107,N_4791);
nand U7230 (N_7230,N_3612,N_3808);
nor U7231 (N_7231,N_58,N_997);
and U7232 (N_7232,N_1858,N_382);
or U7233 (N_7233,N_164,N_4540);
and U7234 (N_7234,N_1563,N_3700);
and U7235 (N_7235,N_1291,N_4250);
and U7236 (N_7236,N_4307,N_2284);
and U7237 (N_7237,N_1610,N_555);
nor U7238 (N_7238,N_4882,N_508);
nand U7239 (N_7239,N_128,N_1543);
or U7240 (N_7240,N_4894,N_4479);
nor U7241 (N_7241,N_2921,N_4010);
nand U7242 (N_7242,N_628,N_2376);
and U7243 (N_7243,N_4513,N_4146);
nand U7244 (N_7244,N_4154,N_3080);
and U7245 (N_7245,N_3758,N_2693);
nand U7246 (N_7246,N_470,N_3344);
or U7247 (N_7247,N_1533,N_910);
nor U7248 (N_7248,N_1815,N_1387);
and U7249 (N_7249,N_1500,N_3171);
and U7250 (N_7250,N_4410,N_1881);
nand U7251 (N_7251,N_2287,N_103);
nand U7252 (N_7252,N_2049,N_261);
and U7253 (N_7253,N_487,N_3569);
nand U7254 (N_7254,N_979,N_4579);
or U7255 (N_7255,N_346,N_4181);
nand U7256 (N_7256,N_1063,N_4121);
and U7257 (N_7257,N_16,N_929);
or U7258 (N_7258,N_1003,N_142);
or U7259 (N_7259,N_1440,N_3716);
nor U7260 (N_7260,N_1213,N_1424);
nor U7261 (N_7261,N_4858,N_4407);
nand U7262 (N_7262,N_4050,N_2263);
or U7263 (N_7263,N_986,N_4040);
or U7264 (N_7264,N_611,N_567);
nor U7265 (N_7265,N_4328,N_1043);
or U7266 (N_7266,N_3590,N_109);
nand U7267 (N_7267,N_637,N_4135);
or U7268 (N_7268,N_1761,N_4778);
nand U7269 (N_7269,N_4546,N_1968);
nand U7270 (N_7270,N_4125,N_3916);
or U7271 (N_7271,N_1501,N_1456);
nor U7272 (N_7272,N_1757,N_4768);
nand U7273 (N_7273,N_3165,N_188);
nand U7274 (N_7274,N_1640,N_1651);
and U7275 (N_7275,N_4179,N_1700);
or U7276 (N_7276,N_1014,N_1981);
nand U7277 (N_7277,N_1251,N_1378);
nand U7278 (N_7278,N_2696,N_847);
xnor U7279 (N_7279,N_472,N_3327);
and U7280 (N_7280,N_4658,N_4517);
nand U7281 (N_7281,N_1667,N_2345);
nand U7282 (N_7282,N_2122,N_3180);
and U7283 (N_7283,N_3026,N_1462);
and U7284 (N_7284,N_621,N_2842);
or U7285 (N_7285,N_47,N_3449);
nor U7286 (N_7286,N_1468,N_4371);
nand U7287 (N_7287,N_1022,N_2220);
and U7288 (N_7288,N_3016,N_1093);
nand U7289 (N_7289,N_1550,N_4644);
and U7290 (N_7290,N_2138,N_3805);
xor U7291 (N_7291,N_3311,N_4212);
nand U7292 (N_7292,N_2929,N_1496);
or U7293 (N_7293,N_3705,N_3610);
nor U7294 (N_7294,N_2908,N_1948);
nor U7295 (N_7295,N_1390,N_293);
nor U7296 (N_7296,N_4970,N_2983);
nor U7297 (N_7297,N_2992,N_732);
nand U7298 (N_7298,N_3243,N_2062);
and U7299 (N_7299,N_4004,N_3751);
or U7300 (N_7300,N_4006,N_542);
nand U7301 (N_7301,N_104,N_862);
nor U7302 (N_7302,N_4303,N_3672);
nand U7303 (N_7303,N_3052,N_4749);
or U7304 (N_7304,N_4845,N_779);
nor U7305 (N_7305,N_4899,N_3075);
and U7306 (N_7306,N_4667,N_305);
nand U7307 (N_7307,N_2825,N_1048);
nand U7308 (N_7308,N_232,N_953);
nand U7309 (N_7309,N_1292,N_2889);
and U7310 (N_7310,N_4164,N_770);
or U7311 (N_7311,N_573,N_1584);
and U7312 (N_7312,N_933,N_3661);
nand U7313 (N_7313,N_727,N_2116);
or U7314 (N_7314,N_283,N_2016);
nor U7315 (N_7315,N_4630,N_3309);
nor U7316 (N_7316,N_227,N_1061);
and U7317 (N_7317,N_1705,N_1412);
nand U7318 (N_7318,N_2657,N_3286);
or U7319 (N_7319,N_2490,N_2829);
nand U7320 (N_7320,N_506,N_2136);
and U7321 (N_7321,N_3635,N_127);
and U7322 (N_7322,N_3221,N_150);
and U7323 (N_7323,N_494,N_4509);
or U7324 (N_7324,N_831,N_2966);
and U7325 (N_7325,N_731,N_2195);
nor U7326 (N_7326,N_2852,N_947);
nor U7327 (N_7327,N_1965,N_697);
or U7328 (N_7328,N_3896,N_1850);
nand U7329 (N_7329,N_2931,N_632);
or U7330 (N_7330,N_1095,N_1431);
or U7331 (N_7331,N_419,N_2509);
or U7332 (N_7332,N_863,N_1441);
and U7333 (N_7333,N_417,N_3801);
nor U7334 (N_7334,N_3270,N_1586);
and U7335 (N_7335,N_1485,N_3144);
nand U7336 (N_7336,N_2481,N_4675);
and U7337 (N_7337,N_544,N_1669);
nor U7338 (N_7338,N_3629,N_3550);
nand U7339 (N_7339,N_3729,N_1671);
nand U7340 (N_7340,N_2973,N_1100);
or U7341 (N_7341,N_1759,N_728);
or U7342 (N_7342,N_323,N_3538);
nor U7343 (N_7343,N_2851,N_1425);
nand U7344 (N_7344,N_4017,N_2098);
nor U7345 (N_7345,N_1609,N_4495);
and U7346 (N_7346,N_4097,N_1663);
or U7347 (N_7347,N_2616,N_3938);
nor U7348 (N_7348,N_2408,N_133);
or U7349 (N_7349,N_1285,N_4271);
and U7350 (N_7350,N_1877,N_3461);
and U7351 (N_7351,N_3676,N_1270);
and U7352 (N_7352,N_1507,N_990);
nand U7353 (N_7353,N_2368,N_2042);
and U7354 (N_7354,N_92,N_3784);
and U7355 (N_7355,N_1076,N_1078);
and U7356 (N_7356,N_3319,N_3351);
nand U7357 (N_7357,N_2602,N_2103);
or U7358 (N_7358,N_1127,N_3901);
and U7359 (N_7359,N_4843,N_1089);
nand U7360 (N_7360,N_302,N_2946);
nand U7361 (N_7361,N_4086,N_2548);
nand U7362 (N_7362,N_1113,N_2045);
nor U7363 (N_7363,N_1702,N_2252);
nand U7364 (N_7364,N_685,N_4867);
nand U7365 (N_7365,N_4184,N_370);
or U7366 (N_7366,N_2844,N_2154);
nand U7367 (N_7367,N_582,N_1648);
or U7368 (N_7368,N_3812,N_1289);
nor U7369 (N_7369,N_610,N_1631);
and U7370 (N_7370,N_1718,N_4783);
or U7371 (N_7371,N_3659,N_4185);
nor U7372 (N_7372,N_3827,N_2209);
nand U7373 (N_7373,N_4104,N_2577);
nand U7374 (N_7374,N_650,N_2099);
or U7375 (N_7375,N_4798,N_1033);
and U7376 (N_7376,N_1484,N_2491);
and U7377 (N_7377,N_2270,N_3222);
nand U7378 (N_7378,N_1002,N_958);
nand U7379 (N_7379,N_4220,N_1777);
nor U7380 (N_7380,N_4541,N_3833);
and U7381 (N_7381,N_3545,N_2294);
or U7382 (N_7382,N_4187,N_2779);
nand U7383 (N_7383,N_1751,N_463);
nand U7384 (N_7384,N_4573,N_4150);
nand U7385 (N_7385,N_1269,N_2397);
and U7386 (N_7386,N_1155,N_4458);
and U7387 (N_7387,N_2250,N_4210);
or U7388 (N_7388,N_564,N_1491);
nor U7389 (N_7389,N_4402,N_3499);
and U7390 (N_7390,N_2924,N_475);
or U7391 (N_7391,N_3134,N_1406);
or U7392 (N_7392,N_1426,N_2227);
xor U7393 (N_7393,N_2484,N_3955);
nor U7394 (N_7394,N_4274,N_3201);
and U7395 (N_7395,N_2894,N_1806);
nand U7396 (N_7396,N_451,N_163);
nand U7397 (N_7397,N_3607,N_4144);
and U7398 (N_7398,N_3108,N_4013);
and U7399 (N_7399,N_4280,N_2835);
or U7400 (N_7400,N_1122,N_2634);
nand U7401 (N_7401,N_4401,N_4404);
and U7402 (N_7402,N_2712,N_1927);
or U7403 (N_7403,N_338,N_1906);
nand U7404 (N_7404,N_3349,N_410);
nor U7405 (N_7405,N_2858,N_2606);
nand U7406 (N_7406,N_3810,N_1889);
nor U7407 (N_7407,N_3744,N_1905);
nand U7408 (N_7408,N_1241,N_3038);
nor U7409 (N_7409,N_1857,N_2351);
nand U7410 (N_7410,N_1612,N_3855);
nand U7411 (N_7411,N_2860,N_617);
nand U7412 (N_7412,N_938,N_2058);
nor U7413 (N_7413,N_50,N_4379);
nor U7414 (N_7414,N_2893,N_3322);
nand U7415 (N_7415,N_2498,N_2731);
and U7416 (N_7416,N_4617,N_4639);
nor U7417 (N_7417,N_4986,N_1030);
and U7418 (N_7418,N_1688,N_823);
nand U7419 (N_7419,N_3045,N_4);
and U7420 (N_7420,N_638,N_2328);
and U7421 (N_7421,N_2008,N_4694);
nand U7422 (N_7422,N_1915,N_1575);
nand U7423 (N_7423,N_1082,N_1637);
nand U7424 (N_7424,N_4335,N_1437);
nand U7425 (N_7425,N_1661,N_1088);
nand U7426 (N_7426,N_1891,N_516);
nor U7427 (N_7427,N_2086,N_1075);
nor U7428 (N_7428,N_1006,N_2340);
nor U7429 (N_7429,N_651,N_4943);
or U7430 (N_7430,N_3468,N_1460);
nand U7431 (N_7431,N_2680,N_2915);
nand U7432 (N_7432,N_750,N_1212);
and U7433 (N_7433,N_3297,N_4349);
and U7434 (N_7434,N_4359,N_1709);
nand U7435 (N_7435,N_931,N_3195);
nor U7436 (N_7436,N_1300,N_4105);
nand U7437 (N_7437,N_192,N_630);
nand U7438 (N_7438,N_702,N_3773);
nand U7439 (N_7439,N_2821,N_4627);
nand U7440 (N_7440,N_3032,N_681);
or U7441 (N_7441,N_2212,N_3140);
nor U7442 (N_7442,N_782,N_3429);
or U7443 (N_7443,N_1129,N_4080);
nand U7444 (N_7444,N_1568,N_3642);
and U7445 (N_7445,N_2943,N_4539);
nand U7446 (N_7446,N_4915,N_3862);
or U7447 (N_7447,N_2610,N_96);
and U7448 (N_7448,N_3614,N_532);
and U7449 (N_7449,N_3187,N_1347);
or U7450 (N_7450,N_3889,N_1855);
nor U7451 (N_7451,N_4432,N_3948);
nor U7452 (N_7452,N_1135,N_846);
or U7453 (N_7453,N_2126,N_228);
or U7454 (N_7454,N_1332,N_1253);
nand U7455 (N_7455,N_2685,N_670);
nand U7456 (N_7456,N_4522,N_4478);
nand U7457 (N_7457,N_4047,N_285);
or U7458 (N_7458,N_2497,N_3076);
or U7459 (N_7459,N_2776,N_3876);
nand U7460 (N_7460,N_3101,N_367);
nor U7461 (N_7461,N_200,N_1872);
and U7462 (N_7462,N_2217,N_3879);
nor U7463 (N_7463,N_4775,N_177);
or U7464 (N_7464,N_337,N_2432);
nand U7465 (N_7465,N_1521,N_1295);
nor U7466 (N_7466,N_4492,N_1707);
nor U7467 (N_7467,N_2972,N_3087);
nor U7468 (N_7468,N_1256,N_3668);
and U7469 (N_7469,N_4283,N_3412);
or U7470 (N_7470,N_3921,N_1310);
or U7471 (N_7471,N_960,N_999);
and U7472 (N_7472,N_3942,N_777);
or U7473 (N_7473,N_622,N_2308);
or U7474 (N_7474,N_2668,N_1859);
and U7475 (N_7475,N_3715,N_1472);
or U7476 (N_7476,N_1539,N_2897);
nand U7477 (N_7477,N_3287,N_1743);
or U7478 (N_7478,N_1416,N_3040);
nor U7479 (N_7479,N_4230,N_3113);
and U7480 (N_7480,N_3775,N_623);
or U7481 (N_7481,N_498,N_453);
nor U7482 (N_7482,N_3500,N_1978);
or U7483 (N_7483,N_1070,N_48);
and U7484 (N_7484,N_3544,N_3491);
nor U7485 (N_7485,N_329,N_2248);
nor U7486 (N_7486,N_2030,N_4609);
nand U7487 (N_7487,N_2697,N_2967);
and U7488 (N_7488,N_1103,N_946);
or U7489 (N_7489,N_1973,N_1655);
nor U7490 (N_7490,N_606,N_479);
nand U7491 (N_7491,N_519,N_2359);
or U7492 (N_7492,N_2534,N_4169);
nor U7493 (N_7493,N_4264,N_4452);
nand U7494 (N_7494,N_1794,N_1627);
and U7495 (N_7495,N_896,N_2040);
or U7496 (N_7496,N_3370,N_4282);
nor U7497 (N_7497,N_2886,N_2848);
nand U7498 (N_7498,N_4631,N_32);
or U7499 (N_7499,N_3372,N_3650);
nor U7500 (N_7500,N_4550,N_1430);
or U7501 (N_7501,N_2597,N_1494);
or U7502 (N_7502,N_4733,N_3401);
and U7503 (N_7503,N_2969,N_1083);
nand U7504 (N_7504,N_4876,N_2540);
or U7505 (N_7505,N_2597,N_3578);
or U7506 (N_7506,N_1741,N_2584);
nand U7507 (N_7507,N_2657,N_1975);
nor U7508 (N_7508,N_4793,N_627);
and U7509 (N_7509,N_1975,N_211);
nor U7510 (N_7510,N_4895,N_2912);
or U7511 (N_7511,N_2300,N_2102);
nor U7512 (N_7512,N_4549,N_1020);
nor U7513 (N_7513,N_1067,N_1899);
nor U7514 (N_7514,N_4103,N_2419);
and U7515 (N_7515,N_1171,N_3908);
or U7516 (N_7516,N_756,N_3803);
or U7517 (N_7517,N_3512,N_685);
and U7518 (N_7518,N_2923,N_709);
nand U7519 (N_7519,N_1668,N_1504);
nor U7520 (N_7520,N_4892,N_1850);
nor U7521 (N_7521,N_2811,N_2069);
nor U7522 (N_7522,N_1355,N_3010);
nor U7523 (N_7523,N_3456,N_157);
or U7524 (N_7524,N_2242,N_2146);
nand U7525 (N_7525,N_4431,N_1369);
nor U7526 (N_7526,N_3845,N_2773);
and U7527 (N_7527,N_743,N_1097);
xnor U7528 (N_7528,N_267,N_4463);
and U7529 (N_7529,N_4069,N_1116);
or U7530 (N_7530,N_554,N_2494);
nor U7531 (N_7531,N_3907,N_4318);
nor U7532 (N_7532,N_229,N_4050);
or U7533 (N_7533,N_3623,N_1305);
or U7534 (N_7534,N_3565,N_3796);
nand U7535 (N_7535,N_4662,N_3287);
nand U7536 (N_7536,N_4071,N_2017);
and U7537 (N_7537,N_2120,N_485);
and U7538 (N_7538,N_2156,N_3698);
nor U7539 (N_7539,N_3700,N_2248);
and U7540 (N_7540,N_3519,N_3926);
or U7541 (N_7541,N_3815,N_1591);
nor U7542 (N_7542,N_2372,N_168);
and U7543 (N_7543,N_4703,N_2505);
nand U7544 (N_7544,N_1651,N_1628);
or U7545 (N_7545,N_2415,N_2480);
nor U7546 (N_7546,N_4784,N_4833);
and U7547 (N_7547,N_863,N_2680);
or U7548 (N_7548,N_4467,N_2809);
nor U7549 (N_7549,N_2048,N_3251);
and U7550 (N_7550,N_4540,N_4101);
nor U7551 (N_7551,N_4261,N_3971);
and U7552 (N_7552,N_460,N_4849);
and U7553 (N_7553,N_3926,N_2586);
or U7554 (N_7554,N_253,N_3917);
or U7555 (N_7555,N_2889,N_3129);
nor U7556 (N_7556,N_4751,N_1558);
and U7557 (N_7557,N_2488,N_4547);
or U7558 (N_7558,N_4012,N_838);
xor U7559 (N_7559,N_3243,N_1466);
or U7560 (N_7560,N_1359,N_2643);
or U7561 (N_7561,N_2338,N_1938);
or U7562 (N_7562,N_3943,N_3307);
nand U7563 (N_7563,N_2520,N_1820);
nor U7564 (N_7564,N_1781,N_3688);
nand U7565 (N_7565,N_3059,N_4690);
nand U7566 (N_7566,N_126,N_2360);
and U7567 (N_7567,N_4781,N_2452);
nor U7568 (N_7568,N_1578,N_2301);
and U7569 (N_7569,N_4535,N_180);
xnor U7570 (N_7570,N_1168,N_2123);
nor U7571 (N_7571,N_3210,N_3803);
and U7572 (N_7572,N_1023,N_3546);
nand U7573 (N_7573,N_4709,N_3505);
and U7574 (N_7574,N_1213,N_514);
nand U7575 (N_7575,N_1563,N_959);
and U7576 (N_7576,N_1890,N_4230);
nor U7577 (N_7577,N_1152,N_427);
nor U7578 (N_7578,N_93,N_3760);
nand U7579 (N_7579,N_4807,N_4264);
nor U7580 (N_7580,N_4588,N_1289);
or U7581 (N_7581,N_4837,N_4566);
or U7582 (N_7582,N_2191,N_1527);
nand U7583 (N_7583,N_93,N_2228);
nor U7584 (N_7584,N_3767,N_1052);
nor U7585 (N_7585,N_699,N_4332);
nand U7586 (N_7586,N_3099,N_1057);
nand U7587 (N_7587,N_1207,N_497);
nor U7588 (N_7588,N_4758,N_1721);
and U7589 (N_7589,N_4302,N_3845);
and U7590 (N_7590,N_3265,N_1467);
nand U7591 (N_7591,N_552,N_2986);
and U7592 (N_7592,N_3863,N_234);
nor U7593 (N_7593,N_1574,N_2696);
nor U7594 (N_7594,N_3777,N_3556);
nor U7595 (N_7595,N_1325,N_1426);
and U7596 (N_7596,N_739,N_3610);
or U7597 (N_7597,N_3505,N_897);
and U7598 (N_7598,N_4766,N_1356);
nor U7599 (N_7599,N_3209,N_1748);
nand U7600 (N_7600,N_2554,N_3201);
and U7601 (N_7601,N_2552,N_4047);
nor U7602 (N_7602,N_3288,N_932);
nor U7603 (N_7603,N_3955,N_4242);
nor U7604 (N_7604,N_3971,N_4352);
nor U7605 (N_7605,N_4437,N_3729);
and U7606 (N_7606,N_714,N_3993);
or U7607 (N_7607,N_2903,N_3322);
and U7608 (N_7608,N_2382,N_1971);
xnor U7609 (N_7609,N_2069,N_1266);
nor U7610 (N_7610,N_2170,N_3005);
nand U7611 (N_7611,N_4791,N_1270);
and U7612 (N_7612,N_2074,N_2946);
and U7613 (N_7613,N_3347,N_4490);
or U7614 (N_7614,N_3688,N_4916);
nor U7615 (N_7615,N_1287,N_4002);
nand U7616 (N_7616,N_443,N_3531);
nor U7617 (N_7617,N_439,N_4788);
nor U7618 (N_7618,N_2741,N_3551);
and U7619 (N_7619,N_2079,N_1608);
nor U7620 (N_7620,N_3814,N_2717);
or U7621 (N_7621,N_2432,N_958);
and U7622 (N_7622,N_1777,N_2444);
and U7623 (N_7623,N_3098,N_3980);
nand U7624 (N_7624,N_570,N_3942);
and U7625 (N_7625,N_368,N_3460);
nand U7626 (N_7626,N_2004,N_1618);
nand U7627 (N_7627,N_632,N_4621);
nor U7628 (N_7628,N_4639,N_1);
and U7629 (N_7629,N_1061,N_546);
and U7630 (N_7630,N_157,N_2602);
or U7631 (N_7631,N_3142,N_3134);
nor U7632 (N_7632,N_3902,N_256);
or U7633 (N_7633,N_2892,N_4647);
and U7634 (N_7634,N_3532,N_3990);
and U7635 (N_7635,N_3010,N_4030);
nor U7636 (N_7636,N_4893,N_192);
nor U7637 (N_7637,N_4647,N_3152);
nand U7638 (N_7638,N_3427,N_1147);
nand U7639 (N_7639,N_2206,N_987);
or U7640 (N_7640,N_1019,N_2166);
nand U7641 (N_7641,N_1883,N_3339);
nand U7642 (N_7642,N_13,N_962);
or U7643 (N_7643,N_1605,N_909);
nor U7644 (N_7644,N_3560,N_2481);
nor U7645 (N_7645,N_485,N_3328);
or U7646 (N_7646,N_2078,N_3950);
or U7647 (N_7647,N_2556,N_880);
or U7648 (N_7648,N_110,N_959);
nor U7649 (N_7649,N_4124,N_2719);
xor U7650 (N_7650,N_1731,N_1772);
nor U7651 (N_7651,N_1913,N_3947);
nor U7652 (N_7652,N_1756,N_1878);
or U7653 (N_7653,N_4007,N_633);
nor U7654 (N_7654,N_2123,N_1293);
nand U7655 (N_7655,N_2557,N_267);
and U7656 (N_7656,N_2719,N_1014);
or U7657 (N_7657,N_1278,N_3603);
and U7658 (N_7658,N_1684,N_3338);
or U7659 (N_7659,N_3849,N_1371);
nand U7660 (N_7660,N_80,N_2447);
nand U7661 (N_7661,N_2053,N_457);
nor U7662 (N_7662,N_1195,N_2486);
and U7663 (N_7663,N_4338,N_320);
and U7664 (N_7664,N_3665,N_4177);
nand U7665 (N_7665,N_2262,N_2463);
or U7666 (N_7666,N_2758,N_4374);
nand U7667 (N_7667,N_4839,N_2746);
nor U7668 (N_7668,N_2684,N_2742);
nor U7669 (N_7669,N_2583,N_1119);
and U7670 (N_7670,N_4114,N_1423);
or U7671 (N_7671,N_4849,N_3347);
nor U7672 (N_7672,N_306,N_1774);
or U7673 (N_7673,N_2848,N_4223);
nand U7674 (N_7674,N_4725,N_269);
or U7675 (N_7675,N_611,N_2704);
nand U7676 (N_7676,N_2875,N_1075);
or U7677 (N_7677,N_3394,N_294);
nor U7678 (N_7678,N_1408,N_2286);
and U7679 (N_7679,N_699,N_3262);
or U7680 (N_7680,N_1379,N_3331);
nand U7681 (N_7681,N_3757,N_1754);
nor U7682 (N_7682,N_1873,N_2513);
and U7683 (N_7683,N_3310,N_2553);
nand U7684 (N_7684,N_3888,N_2398);
xnor U7685 (N_7685,N_3925,N_3594);
nand U7686 (N_7686,N_3996,N_3543);
or U7687 (N_7687,N_4776,N_3534);
nor U7688 (N_7688,N_643,N_4551);
nand U7689 (N_7689,N_1843,N_3506);
and U7690 (N_7690,N_269,N_3210);
nor U7691 (N_7691,N_3540,N_2311);
and U7692 (N_7692,N_3698,N_2949);
or U7693 (N_7693,N_1729,N_4694);
or U7694 (N_7694,N_3615,N_2042);
or U7695 (N_7695,N_1371,N_3279);
or U7696 (N_7696,N_2402,N_79);
and U7697 (N_7697,N_4035,N_2536);
xnor U7698 (N_7698,N_4074,N_17);
nor U7699 (N_7699,N_1453,N_2774);
and U7700 (N_7700,N_4793,N_3817);
nand U7701 (N_7701,N_1946,N_1597);
nor U7702 (N_7702,N_1539,N_1585);
or U7703 (N_7703,N_513,N_2170);
xor U7704 (N_7704,N_3320,N_2404);
or U7705 (N_7705,N_3182,N_178);
or U7706 (N_7706,N_3875,N_2903);
nor U7707 (N_7707,N_111,N_1500);
nand U7708 (N_7708,N_4962,N_2663);
and U7709 (N_7709,N_3816,N_3850);
nand U7710 (N_7710,N_2356,N_1185);
nor U7711 (N_7711,N_3970,N_2518);
and U7712 (N_7712,N_3926,N_1941);
nand U7713 (N_7713,N_2968,N_3476);
nand U7714 (N_7714,N_1931,N_553);
or U7715 (N_7715,N_1783,N_2427);
or U7716 (N_7716,N_1836,N_2716);
or U7717 (N_7717,N_2456,N_4183);
nor U7718 (N_7718,N_3584,N_348);
or U7719 (N_7719,N_2672,N_3866);
and U7720 (N_7720,N_4802,N_3649);
nor U7721 (N_7721,N_4161,N_4625);
and U7722 (N_7722,N_1656,N_1555);
nand U7723 (N_7723,N_1499,N_2242);
xnor U7724 (N_7724,N_247,N_1229);
nor U7725 (N_7725,N_1588,N_4350);
nand U7726 (N_7726,N_4678,N_4672);
and U7727 (N_7727,N_1096,N_1935);
nor U7728 (N_7728,N_102,N_4388);
and U7729 (N_7729,N_828,N_1964);
and U7730 (N_7730,N_1010,N_1992);
nand U7731 (N_7731,N_1758,N_3801);
and U7732 (N_7732,N_2009,N_1009);
and U7733 (N_7733,N_239,N_4082);
nand U7734 (N_7734,N_1070,N_2320);
nand U7735 (N_7735,N_75,N_1032);
or U7736 (N_7736,N_1591,N_2942);
nor U7737 (N_7737,N_2508,N_357);
xor U7738 (N_7738,N_4434,N_683);
xor U7739 (N_7739,N_4453,N_3333);
or U7740 (N_7740,N_4328,N_975);
or U7741 (N_7741,N_4208,N_3902);
nor U7742 (N_7742,N_1969,N_1643);
nor U7743 (N_7743,N_3488,N_1634);
and U7744 (N_7744,N_2209,N_4610);
or U7745 (N_7745,N_4537,N_3445);
nand U7746 (N_7746,N_3374,N_2592);
nand U7747 (N_7747,N_3893,N_4828);
nor U7748 (N_7748,N_1278,N_2635);
or U7749 (N_7749,N_3158,N_1536);
or U7750 (N_7750,N_802,N_4643);
xor U7751 (N_7751,N_193,N_1594);
nor U7752 (N_7752,N_783,N_1460);
or U7753 (N_7753,N_1888,N_555);
or U7754 (N_7754,N_2356,N_4156);
xor U7755 (N_7755,N_2205,N_2584);
or U7756 (N_7756,N_514,N_4646);
or U7757 (N_7757,N_843,N_2379);
nor U7758 (N_7758,N_2265,N_471);
and U7759 (N_7759,N_3887,N_4813);
xor U7760 (N_7760,N_178,N_4908);
and U7761 (N_7761,N_3111,N_3507);
or U7762 (N_7762,N_3389,N_1182);
nor U7763 (N_7763,N_2523,N_4848);
and U7764 (N_7764,N_2386,N_3750);
or U7765 (N_7765,N_3600,N_3238);
nand U7766 (N_7766,N_1698,N_799);
nand U7767 (N_7767,N_1414,N_1822);
nor U7768 (N_7768,N_1441,N_2262);
and U7769 (N_7769,N_3374,N_2219);
and U7770 (N_7770,N_879,N_644);
and U7771 (N_7771,N_3457,N_3893);
and U7772 (N_7772,N_333,N_4467);
nand U7773 (N_7773,N_4652,N_4636);
or U7774 (N_7774,N_4645,N_760);
nand U7775 (N_7775,N_2820,N_2865);
nor U7776 (N_7776,N_1380,N_4595);
nand U7777 (N_7777,N_714,N_3184);
nand U7778 (N_7778,N_3934,N_1387);
xor U7779 (N_7779,N_2252,N_2820);
and U7780 (N_7780,N_4782,N_3071);
nor U7781 (N_7781,N_37,N_1423);
nor U7782 (N_7782,N_4897,N_2669);
and U7783 (N_7783,N_2581,N_3934);
nor U7784 (N_7784,N_3710,N_2618);
and U7785 (N_7785,N_4899,N_2001);
nand U7786 (N_7786,N_677,N_2576);
nor U7787 (N_7787,N_458,N_3699);
xnor U7788 (N_7788,N_1870,N_326);
nor U7789 (N_7789,N_1034,N_1018);
nand U7790 (N_7790,N_404,N_3400);
or U7791 (N_7791,N_1652,N_1287);
nand U7792 (N_7792,N_4946,N_2314);
or U7793 (N_7793,N_2282,N_3248);
or U7794 (N_7794,N_1995,N_3345);
or U7795 (N_7795,N_1467,N_1058);
or U7796 (N_7796,N_4756,N_4645);
and U7797 (N_7797,N_3650,N_2037);
nor U7798 (N_7798,N_3397,N_284);
nor U7799 (N_7799,N_73,N_4750);
nand U7800 (N_7800,N_4067,N_560);
and U7801 (N_7801,N_264,N_527);
and U7802 (N_7802,N_416,N_1521);
nor U7803 (N_7803,N_75,N_4104);
and U7804 (N_7804,N_3931,N_2372);
or U7805 (N_7805,N_3408,N_4769);
nor U7806 (N_7806,N_2507,N_440);
xnor U7807 (N_7807,N_2392,N_2296);
or U7808 (N_7808,N_480,N_229);
and U7809 (N_7809,N_3154,N_1523);
nand U7810 (N_7810,N_3479,N_3842);
and U7811 (N_7811,N_4114,N_4547);
and U7812 (N_7812,N_851,N_3731);
nor U7813 (N_7813,N_4564,N_4051);
nand U7814 (N_7814,N_2307,N_4761);
and U7815 (N_7815,N_2391,N_2327);
xnor U7816 (N_7816,N_373,N_2163);
and U7817 (N_7817,N_41,N_3229);
nand U7818 (N_7818,N_1289,N_3512);
nor U7819 (N_7819,N_962,N_2548);
nand U7820 (N_7820,N_2490,N_1973);
nand U7821 (N_7821,N_392,N_2527);
or U7822 (N_7822,N_907,N_4814);
nand U7823 (N_7823,N_2991,N_3744);
nor U7824 (N_7824,N_3907,N_2042);
and U7825 (N_7825,N_864,N_3275);
nand U7826 (N_7826,N_4551,N_3673);
nand U7827 (N_7827,N_807,N_3537);
nor U7828 (N_7828,N_2131,N_1659);
or U7829 (N_7829,N_955,N_926);
nand U7830 (N_7830,N_1729,N_2392);
nor U7831 (N_7831,N_164,N_4651);
or U7832 (N_7832,N_26,N_3584);
and U7833 (N_7833,N_4171,N_3567);
nand U7834 (N_7834,N_4821,N_1958);
or U7835 (N_7835,N_3254,N_1706);
or U7836 (N_7836,N_1173,N_4616);
or U7837 (N_7837,N_3560,N_4711);
nand U7838 (N_7838,N_762,N_2357);
nor U7839 (N_7839,N_3504,N_932);
nand U7840 (N_7840,N_133,N_1018);
and U7841 (N_7841,N_3986,N_642);
and U7842 (N_7842,N_1392,N_1074);
nor U7843 (N_7843,N_4777,N_3364);
nand U7844 (N_7844,N_1032,N_1795);
or U7845 (N_7845,N_3447,N_2086);
nand U7846 (N_7846,N_3653,N_2409);
or U7847 (N_7847,N_3088,N_4999);
and U7848 (N_7848,N_3415,N_4565);
or U7849 (N_7849,N_1021,N_1579);
and U7850 (N_7850,N_1005,N_353);
and U7851 (N_7851,N_3335,N_1148);
nand U7852 (N_7852,N_4382,N_490);
and U7853 (N_7853,N_660,N_4755);
or U7854 (N_7854,N_4683,N_1644);
nand U7855 (N_7855,N_4147,N_4777);
or U7856 (N_7856,N_3442,N_633);
nor U7857 (N_7857,N_2163,N_3540);
nor U7858 (N_7858,N_3605,N_4792);
or U7859 (N_7859,N_1067,N_514);
nand U7860 (N_7860,N_2976,N_2844);
or U7861 (N_7861,N_1257,N_3331);
or U7862 (N_7862,N_3331,N_1804);
nand U7863 (N_7863,N_1806,N_777);
or U7864 (N_7864,N_2002,N_3463);
nand U7865 (N_7865,N_3995,N_916);
or U7866 (N_7866,N_4597,N_915);
and U7867 (N_7867,N_431,N_253);
nand U7868 (N_7868,N_4602,N_3293);
and U7869 (N_7869,N_2170,N_1862);
xnor U7870 (N_7870,N_1515,N_3081);
nand U7871 (N_7871,N_3385,N_2530);
nor U7872 (N_7872,N_1514,N_4638);
nor U7873 (N_7873,N_1423,N_613);
nor U7874 (N_7874,N_41,N_4789);
or U7875 (N_7875,N_3779,N_4772);
and U7876 (N_7876,N_701,N_1066);
nor U7877 (N_7877,N_2424,N_3174);
or U7878 (N_7878,N_2603,N_3195);
nor U7879 (N_7879,N_1579,N_1995);
nor U7880 (N_7880,N_342,N_4744);
and U7881 (N_7881,N_2971,N_1968);
nand U7882 (N_7882,N_383,N_1883);
nor U7883 (N_7883,N_1918,N_3172);
and U7884 (N_7884,N_3450,N_3195);
nand U7885 (N_7885,N_1730,N_1440);
nor U7886 (N_7886,N_2736,N_3222);
and U7887 (N_7887,N_2775,N_2137);
or U7888 (N_7888,N_2362,N_3847);
nand U7889 (N_7889,N_707,N_485);
nand U7890 (N_7890,N_3965,N_2762);
nor U7891 (N_7891,N_3048,N_3153);
and U7892 (N_7892,N_2202,N_166);
or U7893 (N_7893,N_3638,N_766);
nand U7894 (N_7894,N_600,N_4955);
and U7895 (N_7895,N_2520,N_451);
nand U7896 (N_7896,N_2019,N_4056);
and U7897 (N_7897,N_2711,N_4025);
and U7898 (N_7898,N_3319,N_4373);
and U7899 (N_7899,N_2095,N_3812);
nor U7900 (N_7900,N_2389,N_663);
or U7901 (N_7901,N_1790,N_2881);
nor U7902 (N_7902,N_60,N_1147);
nand U7903 (N_7903,N_1828,N_1843);
and U7904 (N_7904,N_4431,N_3913);
or U7905 (N_7905,N_619,N_335);
or U7906 (N_7906,N_4337,N_1395);
or U7907 (N_7907,N_2976,N_1847);
nor U7908 (N_7908,N_2500,N_332);
or U7909 (N_7909,N_2400,N_1921);
nand U7910 (N_7910,N_1444,N_120);
and U7911 (N_7911,N_4751,N_3130);
nor U7912 (N_7912,N_4012,N_2073);
and U7913 (N_7913,N_4076,N_532);
nor U7914 (N_7914,N_4941,N_2245);
nor U7915 (N_7915,N_2188,N_3342);
nor U7916 (N_7916,N_3207,N_346);
and U7917 (N_7917,N_600,N_4378);
or U7918 (N_7918,N_4858,N_2919);
or U7919 (N_7919,N_4502,N_4151);
nor U7920 (N_7920,N_4994,N_4565);
and U7921 (N_7921,N_3626,N_2267);
or U7922 (N_7922,N_1042,N_1396);
nand U7923 (N_7923,N_2302,N_80);
or U7924 (N_7924,N_462,N_2524);
nand U7925 (N_7925,N_2619,N_4513);
or U7926 (N_7926,N_1866,N_290);
or U7927 (N_7927,N_1637,N_1422);
or U7928 (N_7928,N_4964,N_222);
nand U7929 (N_7929,N_1617,N_835);
xnor U7930 (N_7930,N_1745,N_1002);
or U7931 (N_7931,N_2671,N_1440);
and U7932 (N_7932,N_3301,N_2958);
or U7933 (N_7933,N_631,N_1729);
nor U7934 (N_7934,N_1266,N_2020);
nand U7935 (N_7935,N_3670,N_2424);
nand U7936 (N_7936,N_4341,N_1928);
nor U7937 (N_7937,N_3255,N_944);
nand U7938 (N_7938,N_3479,N_829);
and U7939 (N_7939,N_4807,N_950);
nor U7940 (N_7940,N_2977,N_4249);
and U7941 (N_7941,N_1686,N_2207);
and U7942 (N_7942,N_1436,N_3642);
or U7943 (N_7943,N_2271,N_2107);
or U7944 (N_7944,N_2730,N_717);
or U7945 (N_7945,N_17,N_372);
nand U7946 (N_7946,N_3929,N_1609);
nor U7947 (N_7947,N_4217,N_1776);
nor U7948 (N_7948,N_2862,N_241);
nand U7949 (N_7949,N_2314,N_4772);
and U7950 (N_7950,N_1268,N_2742);
and U7951 (N_7951,N_2686,N_153);
and U7952 (N_7952,N_404,N_3629);
xnor U7953 (N_7953,N_4438,N_4120);
nand U7954 (N_7954,N_2419,N_4904);
nor U7955 (N_7955,N_3088,N_755);
or U7956 (N_7956,N_393,N_286);
nand U7957 (N_7957,N_1601,N_3205);
nor U7958 (N_7958,N_4143,N_3813);
nor U7959 (N_7959,N_3090,N_2170);
nor U7960 (N_7960,N_2996,N_4290);
and U7961 (N_7961,N_2261,N_2376);
and U7962 (N_7962,N_3234,N_924);
and U7963 (N_7963,N_1300,N_2003);
nand U7964 (N_7964,N_1547,N_756);
or U7965 (N_7965,N_1021,N_1610);
or U7966 (N_7966,N_565,N_2548);
nand U7967 (N_7967,N_3573,N_1158);
nor U7968 (N_7968,N_1002,N_4443);
or U7969 (N_7969,N_1572,N_1437);
nand U7970 (N_7970,N_3519,N_289);
or U7971 (N_7971,N_4256,N_3014);
and U7972 (N_7972,N_4159,N_1411);
and U7973 (N_7973,N_1001,N_2167);
nor U7974 (N_7974,N_216,N_533);
or U7975 (N_7975,N_3279,N_1641);
or U7976 (N_7976,N_423,N_4938);
or U7977 (N_7977,N_3095,N_2273);
nor U7978 (N_7978,N_2943,N_445);
and U7979 (N_7979,N_1405,N_1329);
nor U7980 (N_7980,N_1086,N_1605);
nand U7981 (N_7981,N_4309,N_2107);
nand U7982 (N_7982,N_97,N_2754);
nand U7983 (N_7983,N_3626,N_312);
or U7984 (N_7984,N_3003,N_2636);
nor U7985 (N_7985,N_2650,N_4615);
nor U7986 (N_7986,N_1741,N_268);
and U7987 (N_7987,N_1396,N_1466);
nand U7988 (N_7988,N_1755,N_873);
nor U7989 (N_7989,N_1051,N_2738);
and U7990 (N_7990,N_1956,N_2716);
and U7991 (N_7991,N_2757,N_1293);
nor U7992 (N_7992,N_4005,N_4670);
and U7993 (N_7993,N_1761,N_3186);
or U7994 (N_7994,N_1950,N_2404);
and U7995 (N_7995,N_1052,N_1205);
or U7996 (N_7996,N_4474,N_2437);
nand U7997 (N_7997,N_4873,N_623);
or U7998 (N_7998,N_723,N_768);
and U7999 (N_7999,N_1795,N_4375);
or U8000 (N_8000,N_4248,N_577);
and U8001 (N_8001,N_3808,N_787);
nor U8002 (N_8002,N_762,N_4836);
or U8003 (N_8003,N_1063,N_3);
nand U8004 (N_8004,N_2980,N_1137);
nand U8005 (N_8005,N_3492,N_4418);
nand U8006 (N_8006,N_2584,N_1540);
and U8007 (N_8007,N_1796,N_1504);
nor U8008 (N_8008,N_444,N_4485);
nand U8009 (N_8009,N_2238,N_1385);
or U8010 (N_8010,N_2646,N_3075);
nor U8011 (N_8011,N_2145,N_4648);
nor U8012 (N_8012,N_4491,N_2052);
nor U8013 (N_8013,N_4340,N_742);
or U8014 (N_8014,N_3546,N_4253);
or U8015 (N_8015,N_3522,N_1989);
nand U8016 (N_8016,N_1844,N_3536);
or U8017 (N_8017,N_512,N_4228);
nand U8018 (N_8018,N_1703,N_767);
nand U8019 (N_8019,N_1414,N_915);
nand U8020 (N_8020,N_1360,N_1705);
or U8021 (N_8021,N_1246,N_786);
nand U8022 (N_8022,N_348,N_3118);
and U8023 (N_8023,N_4924,N_745);
and U8024 (N_8024,N_3450,N_643);
and U8025 (N_8025,N_3819,N_4500);
nand U8026 (N_8026,N_220,N_651);
nand U8027 (N_8027,N_1791,N_3177);
and U8028 (N_8028,N_4733,N_2694);
nand U8029 (N_8029,N_554,N_548);
and U8030 (N_8030,N_1998,N_1854);
and U8031 (N_8031,N_2498,N_2725);
or U8032 (N_8032,N_3826,N_3099);
nand U8033 (N_8033,N_3166,N_3134);
and U8034 (N_8034,N_446,N_3439);
nor U8035 (N_8035,N_659,N_4005);
nor U8036 (N_8036,N_4490,N_3740);
and U8037 (N_8037,N_2798,N_290);
or U8038 (N_8038,N_3894,N_4987);
and U8039 (N_8039,N_2765,N_894);
nor U8040 (N_8040,N_6,N_3360);
or U8041 (N_8041,N_2129,N_1050);
and U8042 (N_8042,N_2322,N_4718);
and U8043 (N_8043,N_2403,N_145);
nor U8044 (N_8044,N_3887,N_4689);
or U8045 (N_8045,N_4552,N_1198);
or U8046 (N_8046,N_2552,N_1075);
or U8047 (N_8047,N_4354,N_1668);
and U8048 (N_8048,N_2763,N_1363);
nand U8049 (N_8049,N_4608,N_4062);
and U8050 (N_8050,N_115,N_125);
and U8051 (N_8051,N_4024,N_2520);
nor U8052 (N_8052,N_2757,N_2559);
or U8053 (N_8053,N_335,N_3957);
or U8054 (N_8054,N_4083,N_280);
and U8055 (N_8055,N_2067,N_507);
nor U8056 (N_8056,N_959,N_4399);
nand U8057 (N_8057,N_529,N_765);
nor U8058 (N_8058,N_1051,N_2934);
and U8059 (N_8059,N_1605,N_2500);
or U8060 (N_8060,N_4030,N_3729);
and U8061 (N_8061,N_4367,N_1930);
or U8062 (N_8062,N_4667,N_457);
nor U8063 (N_8063,N_3496,N_3300);
nor U8064 (N_8064,N_862,N_3526);
nor U8065 (N_8065,N_3258,N_2539);
nor U8066 (N_8066,N_3471,N_559);
xnor U8067 (N_8067,N_4563,N_3648);
nor U8068 (N_8068,N_2870,N_2038);
or U8069 (N_8069,N_4170,N_4629);
and U8070 (N_8070,N_2803,N_1897);
or U8071 (N_8071,N_956,N_2743);
and U8072 (N_8072,N_756,N_2008);
and U8073 (N_8073,N_4022,N_3959);
or U8074 (N_8074,N_3595,N_4022);
nor U8075 (N_8075,N_403,N_2520);
and U8076 (N_8076,N_2944,N_3339);
and U8077 (N_8077,N_3700,N_1885);
and U8078 (N_8078,N_1990,N_4839);
nand U8079 (N_8079,N_382,N_76);
and U8080 (N_8080,N_4777,N_645);
or U8081 (N_8081,N_3586,N_1730);
or U8082 (N_8082,N_1392,N_1485);
nand U8083 (N_8083,N_1984,N_1155);
or U8084 (N_8084,N_381,N_1468);
or U8085 (N_8085,N_1015,N_1510);
nand U8086 (N_8086,N_1456,N_3460);
nand U8087 (N_8087,N_327,N_183);
xnor U8088 (N_8088,N_3340,N_1998);
and U8089 (N_8089,N_4626,N_30);
or U8090 (N_8090,N_922,N_4675);
nand U8091 (N_8091,N_2133,N_1997);
or U8092 (N_8092,N_3931,N_6);
xnor U8093 (N_8093,N_1763,N_4737);
nand U8094 (N_8094,N_3561,N_3192);
nor U8095 (N_8095,N_1949,N_2820);
nand U8096 (N_8096,N_2330,N_3605);
and U8097 (N_8097,N_4408,N_2472);
and U8098 (N_8098,N_1999,N_2398);
or U8099 (N_8099,N_128,N_914);
or U8100 (N_8100,N_2635,N_131);
nand U8101 (N_8101,N_9,N_4104);
and U8102 (N_8102,N_2493,N_4428);
or U8103 (N_8103,N_3304,N_3025);
or U8104 (N_8104,N_3824,N_4139);
nand U8105 (N_8105,N_125,N_247);
nand U8106 (N_8106,N_2559,N_4702);
nand U8107 (N_8107,N_1157,N_1605);
nand U8108 (N_8108,N_2316,N_2254);
nand U8109 (N_8109,N_2206,N_3060);
and U8110 (N_8110,N_4268,N_3505);
nor U8111 (N_8111,N_2475,N_3036);
and U8112 (N_8112,N_236,N_3669);
nor U8113 (N_8113,N_3750,N_3236);
or U8114 (N_8114,N_1394,N_4697);
nor U8115 (N_8115,N_1181,N_2558);
nor U8116 (N_8116,N_4961,N_1415);
nor U8117 (N_8117,N_271,N_711);
nand U8118 (N_8118,N_135,N_618);
nor U8119 (N_8119,N_1926,N_3307);
and U8120 (N_8120,N_2936,N_4438);
or U8121 (N_8121,N_3968,N_3352);
nand U8122 (N_8122,N_4542,N_1231);
nand U8123 (N_8123,N_4377,N_3741);
xnor U8124 (N_8124,N_808,N_1313);
nand U8125 (N_8125,N_842,N_4466);
and U8126 (N_8126,N_3731,N_4542);
and U8127 (N_8127,N_4946,N_2963);
nand U8128 (N_8128,N_1773,N_4868);
or U8129 (N_8129,N_3961,N_619);
and U8130 (N_8130,N_949,N_3762);
nor U8131 (N_8131,N_2799,N_1786);
or U8132 (N_8132,N_2914,N_4749);
or U8133 (N_8133,N_4857,N_4036);
nand U8134 (N_8134,N_3530,N_4027);
or U8135 (N_8135,N_3619,N_3797);
and U8136 (N_8136,N_3279,N_922);
and U8137 (N_8137,N_1649,N_1195);
or U8138 (N_8138,N_835,N_2718);
nor U8139 (N_8139,N_2766,N_1859);
and U8140 (N_8140,N_773,N_3718);
and U8141 (N_8141,N_2878,N_610);
nor U8142 (N_8142,N_4176,N_4769);
and U8143 (N_8143,N_4401,N_180);
nand U8144 (N_8144,N_2119,N_4133);
nand U8145 (N_8145,N_1247,N_1381);
nand U8146 (N_8146,N_100,N_2904);
or U8147 (N_8147,N_2305,N_4255);
xnor U8148 (N_8148,N_261,N_2449);
nand U8149 (N_8149,N_2592,N_4373);
nor U8150 (N_8150,N_1559,N_2019);
and U8151 (N_8151,N_4161,N_462);
or U8152 (N_8152,N_2698,N_3010);
nand U8153 (N_8153,N_1741,N_833);
or U8154 (N_8154,N_2191,N_4505);
or U8155 (N_8155,N_2050,N_2538);
nor U8156 (N_8156,N_2740,N_4320);
nor U8157 (N_8157,N_311,N_4678);
or U8158 (N_8158,N_327,N_1993);
or U8159 (N_8159,N_2788,N_1106);
nor U8160 (N_8160,N_425,N_1332);
nor U8161 (N_8161,N_2039,N_3189);
nor U8162 (N_8162,N_330,N_4625);
and U8163 (N_8163,N_2919,N_3229);
nor U8164 (N_8164,N_75,N_3101);
or U8165 (N_8165,N_2822,N_4075);
nand U8166 (N_8166,N_1934,N_691);
or U8167 (N_8167,N_3295,N_3598);
and U8168 (N_8168,N_1165,N_4957);
and U8169 (N_8169,N_1297,N_1940);
or U8170 (N_8170,N_2673,N_662);
nor U8171 (N_8171,N_3981,N_2146);
nor U8172 (N_8172,N_1355,N_1690);
nor U8173 (N_8173,N_1763,N_2831);
or U8174 (N_8174,N_3291,N_4734);
and U8175 (N_8175,N_34,N_2713);
or U8176 (N_8176,N_4038,N_886);
xor U8177 (N_8177,N_3672,N_4094);
nand U8178 (N_8178,N_892,N_2754);
nor U8179 (N_8179,N_3915,N_1496);
nand U8180 (N_8180,N_2607,N_1743);
and U8181 (N_8181,N_4054,N_2592);
nor U8182 (N_8182,N_4037,N_288);
nor U8183 (N_8183,N_4546,N_4413);
nor U8184 (N_8184,N_3827,N_3852);
and U8185 (N_8185,N_322,N_2435);
xor U8186 (N_8186,N_4397,N_2643);
or U8187 (N_8187,N_862,N_1827);
nand U8188 (N_8188,N_3823,N_4098);
nand U8189 (N_8189,N_911,N_1156);
and U8190 (N_8190,N_1573,N_3527);
or U8191 (N_8191,N_1364,N_1418);
and U8192 (N_8192,N_2141,N_3299);
and U8193 (N_8193,N_1373,N_3385);
and U8194 (N_8194,N_256,N_4754);
nor U8195 (N_8195,N_4071,N_3507);
and U8196 (N_8196,N_4375,N_770);
nor U8197 (N_8197,N_1405,N_2973);
and U8198 (N_8198,N_686,N_1304);
or U8199 (N_8199,N_4093,N_3396);
and U8200 (N_8200,N_1517,N_136);
nor U8201 (N_8201,N_1884,N_4619);
nor U8202 (N_8202,N_4680,N_104);
or U8203 (N_8203,N_4505,N_2192);
nand U8204 (N_8204,N_2486,N_2646);
or U8205 (N_8205,N_1375,N_3209);
nor U8206 (N_8206,N_3602,N_4323);
nand U8207 (N_8207,N_3904,N_1478);
nand U8208 (N_8208,N_3573,N_4179);
nand U8209 (N_8209,N_3341,N_3024);
and U8210 (N_8210,N_1552,N_363);
and U8211 (N_8211,N_3634,N_80);
or U8212 (N_8212,N_2993,N_74);
and U8213 (N_8213,N_3781,N_1447);
nand U8214 (N_8214,N_4556,N_1584);
nand U8215 (N_8215,N_3846,N_2662);
nand U8216 (N_8216,N_3951,N_3851);
or U8217 (N_8217,N_2828,N_3561);
and U8218 (N_8218,N_1559,N_4525);
nand U8219 (N_8219,N_3598,N_1021);
nand U8220 (N_8220,N_867,N_3398);
or U8221 (N_8221,N_3840,N_1177);
nand U8222 (N_8222,N_3345,N_3899);
nor U8223 (N_8223,N_123,N_3778);
and U8224 (N_8224,N_4938,N_3483);
and U8225 (N_8225,N_4862,N_4517);
nand U8226 (N_8226,N_965,N_2853);
nand U8227 (N_8227,N_3092,N_4563);
or U8228 (N_8228,N_528,N_3405);
or U8229 (N_8229,N_4801,N_3397);
or U8230 (N_8230,N_4571,N_4586);
or U8231 (N_8231,N_381,N_1794);
and U8232 (N_8232,N_907,N_4415);
or U8233 (N_8233,N_3751,N_1476);
and U8234 (N_8234,N_1320,N_1605);
nand U8235 (N_8235,N_3357,N_2074);
or U8236 (N_8236,N_2597,N_3211);
and U8237 (N_8237,N_4099,N_3488);
or U8238 (N_8238,N_4219,N_2218);
nand U8239 (N_8239,N_3266,N_2957);
nor U8240 (N_8240,N_4507,N_2050);
or U8241 (N_8241,N_4077,N_713);
and U8242 (N_8242,N_2950,N_955);
nand U8243 (N_8243,N_622,N_2572);
nor U8244 (N_8244,N_3772,N_576);
and U8245 (N_8245,N_966,N_3989);
nor U8246 (N_8246,N_1997,N_924);
and U8247 (N_8247,N_256,N_39);
nand U8248 (N_8248,N_3101,N_4101);
or U8249 (N_8249,N_4980,N_4060);
nor U8250 (N_8250,N_1772,N_4630);
and U8251 (N_8251,N_4479,N_4388);
nor U8252 (N_8252,N_1944,N_1373);
and U8253 (N_8253,N_574,N_3357);
or U8254 (N_8254,N_4674,N_4109);
and U8255 (N_8255,N_1919,N_581);
or U8256 (N_8256,N_386,N_80);
and U8257 (N_8257,N_2800,N_1532);
nand U8258 (N_8258,N_4051,N_250);
nand U8259 (N_8259,N_2729,N_860);
nand U8260 (N_8260,N_1453,N_2945);
or U8261 (N_8261,N_4110,N_2254);
nand U8262 (N_8262,N_3200,N_515);
nor U8263 (N_8263,N_3928,N_4852);
nand U8264 (N_8264,N_2031,N_819);
and U8265 (N_8265,N_476,N_912);
or U8266 (N_8266,N_1812,N_2098);
nor U8267 (N_8267,N_1452,N_2077);
nor U8268 (N_8268,N_1277,N_1005);
nand U8269 (N_8269,N_1255,N_1276);
nand U8270 (N_8270,N_1100,N_1927);
or U8271 (N_8271,N_4172,N_2222);
nand U8272 (N_8272,N_4778,N_1646);
nor U8273 (N_8273,N_2544,N_918);
and U8274 (N_8274,N_1074,N_4844);
or U8275 (N_8275,N_185,N_1695);
nand U8276 (N_8276,N_4686,N_624);
nor U8277 (N_8277,N_1673,N_3680);
nor U8278 (N_8278,N_2058,N_2701);
and U8279 (N_8279,N_4652,N_3842);
and U8280 (N_8280,N_4732,N_996);
and U8281 (N_8281,N_3443,N_4746);
or U8282 (N_8282,N_3035,N_448);
nand U8283 (N_8283,N_4038,N_4681);
nor U8284 (N_8284,N_2208,N_2956);
nor U8285 (N_8285,N_1985,N_1525);
or U8286 (N_8286,N_2289,N_3700);
nand U8287 (N_8287,N_3074,N_658);
or U8288 (N_8288,N_351,N_2467);
and U8289 (N_8289,N_2535,N_4056);
nor U8290 (N_8290,N_4998,N_2056);
nand U8291 (N_8291,N_3565,N_557);
and U8292 (N_8292,N_1068,N_1117);
nor U8293 (N_8293,N_4888,N_3797);
or U8294 (N_8294,N_4362,N_833);
nand U8295 (N_8295,N_1768,N_529);
or U8296 (N_8296,N_1809,N_2551);
nand U8297 (N_8297,N_4065,N_4336);
and U8298 (N_8298,N_1621,N_1545);
nand U8299 (N_8299,N_4019,N_1091);
nor U8300 (N_8300,N_4054,N_3653);
nor U8301 (N_8301,N_2419,N_1505);
nand U8302 (N_8302,N_208,N_3895);
or U8303 (N_8303,N_2925,N_3643);
nor U8304 (N_8304,N_1579,N_2403);
nand U8305 (N_8305,N_3239,N_3349);
or U8306 (N_8306,N_4532,N_3424);
nand U8307 (N_8307,N_1669,N_1173);
nor U8308 (N_8308,N_3282,N_4916);
xnor U8309 (N_8309,N_687,N_1312);
or U8310 (N_8310,N_4546,N_303);
nand U8311 (N_8311,N_21,N_1375);
nand U8312 (N_8312,N_4319,N_19);
or U8313 (N_8313,N_4697,N_2919);
nor U8314 (N_8314,N_4941,N_4921);
and U8315 (N_8315,N_1579,N_3037);
and U8316 (N_8316,N_3339,N_215);
or U8317 (N_8317,N_2000,N_4907);
nand U8318 (N_8318,N_2138,N_1721);
nor U8319 (N_8319,N_2558,N_454);
nor U8320 (N_8320,N_2096,N_1352);
or U8321 (N_8321,N_4237,N_2604);
xnor U8322 (N_8322,N_3662,N_4760);
nor U8323 (N_8323,N_4978,N_431);
nand U8324 (N_8324,N_445,N_4674);
xor U8325 (N_8325,N_3991,N_4221);
or U8326 (N_8326,N_2953,N_2682);
nand U8327 (N_8327,N_4088,N_2676);
and U8328 (N_8328,N_1249,N_2799);
nand U8329 (N_8329,N_378,N_3561);
xnor U8330 (N_8330,N_295,N_3847);
or U8331 (N_8331,N_4929,N_4893);
nor U8332 (N_8332,N_1582,N_504);
nand U8333 (N_8333,N_3581,N_237);
and U8334 (N_8334,N_1660,N_1581);
xnor U8335 (N_8335,N_2285,N_8);
and U8336 (N_8336,N_876,N_813);
or U8337 (N_8337,N_3985,N_4766);
or U8338 (N_8338,N_2691,N_643);
or U8339 (N_8339,N_131,N_4339);
and U8340 (N_8340,N_3603,N_4610);
or U8341 (N_8341,N_3456,N_129);
nor U8342 (N_8342,N_1333,N_2893);
and U8343 (N_8343,N_313,N_3205);
or U8344 (N_8344,N_1107,N_3347);
nor U8345 (N_8345,N_1574,N_2574);
or U8346 (N_8346,N_4552,N_1107);
and U8347 (N_8347,N_3678,N_4884);
or U8348 (N_8348,N_1824,N_547);
and U8349 (N_8349,N_1326,N_3350);
or U8350 (N_8350,N_855,N_4072);
nor U8351 (N_8351,N_1275,N_2823);
nand U8352 (N_8352,N_1529,N_3096);
xnor U8353 (N_8353,N_3871,N_884);
nand U8354 (N_8354,N_614,N_1408);
nor U8355 (N_8355,N_2554,N_2315);
xor U8356 (N_8356,N_1667,N_1988);
and U8357 (N_8357,N_3542,N_3619);
nor U8358 (N_8358,N_1428,N_2694);
or U8359 (N_8359,N_636,N_369);
nor U8360 (N_8360,N_2646,N_136);
or U8361 (N_8361,N_2367,N_4193);
nand U8362 (N_8362,N_4253,N_4729);
and U8363 (N_8363,N_3096,N_4314);
nand U8364 (N_8364,N_4354,N_4951);
nand U8365 (N_8365,N_2393,N_1370);
nand U8366 (N_8366,N_4360,N_2350);
or U8367 (N_8367,N_3596,N_3861);
and U8368 (N_8368,N_4078,N_466);
or U8369 (N_8369,N_3338,N_3583);
or U8370 (N_8370,N_1952,N_750);
or U8371 (N_8371,N_3775,N_357);
nor U8372 (N_8372,N_2023,N_134);
or U8373 (N_8373,N_1350,N_619);
nor U8374 (N_8374,N_1590,N_4305);
nor U8375 (N_8375,N_1836,N_4141);
nor U8376 (N_8376,N_2159,N_4979);
and U8377 (N_8377,N_1291,N_1740);
or U8378 (N_8378,N_2169,N_3396);
nor U8379 (N_8379,N_3161,N_3500);
and U8380 (N_8380,N_86,N_708);
or U8381 (N_8381,N_4873,N_1190);
nand U8382 (N_8382,N_3803,N_1814);
and U8383 (N_8383,N_3011,N_1463);
or U8384 (N_8384,N_4245,N_449);
nor U8385 (N_8385,N_4588,N_4251);
or U8386 (N_8386,N_3279,N_4136);
nand U8387 (N_8387,N_1218,N_4751);
and U8388 (N_8388,N_2859,N_2409);
or U8389 (N_8389,N_1981,N_4368);
nor U8390 (N_8390,N_3403,N_2468);
or U8391 (N_8391,N_1019,N_2816);
nand U8392 (N_8392,N_515,N_863);
or U8393 (N_8393,N_1908,N_1569);
and U8394 (N_8394,N_2723,N_4525);
and U8395 (N_8395,N_1037,N_3404);
or U8396 (N_8396,N_1733,N_3637);
nand U8397 (N_8397,N_2219,N_2070);
or U8398 (N_8398,N_3319,N_2825);
or U8399 (N_8399,N_4499,N_2879);
nor U8400 (N_8400,N_3360,N_4402);
nand U8401 (N_8401,N_3785,N_3649);
nand U8402 (N_8402,N_4223,N_3774);
and U8403 (N_8403,N_2774,N_2907);
and U8404 (N_8404,N_3126,N_1890);
nand U8405 (N_8405,N_811,N_1657);
nor U8406 (N_8406,N_3414,N_224);
or U8407 (N_8407,N_597,N_1225);
and U8408 (N_8408,N_728,N_1345);
nor U8409 (N_8409,N_1145,N_817);
and U8410 (N_8410,N_925,N_2859);
and U8411 (N_8411,N_1551,N_242);
nor U8412 (N_8412,N_2935,N_2481);
and U8413 (N_8413,N_3264,N_45);
nand U8414 (N_8414,N_564,N_2762);
nand U8415 (N_8415,N_1724,N_1133);
nor U8416 (N_8416,N_2185,N_246);
nand U8417 (N_8417,N_2916,N_4193);
nand U8418 (N_8418,N_1848,N_3242);
nor U8419 (N_8419,N_2845,N_1340);
or U8420 (N_8420,N_1578,N_1279);
and U8421 (N_8421,N_4876,N_4630);
or U8422 (N_8422,N_2553,N_277);
and U8423 (N_8423,N_31,N_3645);
and U8424 (N_8424,N_3082,N_3045);
nand U8425 (N_8425,N_2030,N_1199);
and U8426 (N_8426,N_2377,N_4721);
nor U8427 (N_8427,N_550,N_1337);
nor U8428 (N_8428,N_2864,N_2067);
nor U8429 (N_8429,N_728,N_2081);
nand U8430 (N_8430,N_578,N_2995);
or U8431 (N_8431,N_842,N_2203);
nand U8432 (N_8432,N_4082,N_2348);
and U8433 (N_8433,N_11,N_1029);
nand U8434 (N_8434,N_4957,N_1788);
nor U8435 (N_8435,N_3432,N_1747);
and U8436 (N_8436,N_1101,N_2229);
nor U8437 (N_8437,N_3499,N_153);
nand U8438 (N_8438,N_2509,N_148);
and U8439 (N_8439,N_1044,N_4086);
nand U8440 (N_8440,N_456,N_2223);
and U8441 (N_8441,N_4654,N_550);
or U8442 (N_8442,N_1309,N_3492);
nand U8443 (N_8443,N_559,N_1912);
nor U8444 (N_8444,N_4089,N_4288);
nand U8445 (N_8445,N_3162,N_3543);
nor U8446 (N_8446,N_2012,N_3700);
and U8447 (N_8447,N_678,N_1015);
nor U8448 (N_8448,N_160,N_553);
or U8449 (N_8449,N_3350,N_221);
nor U8450 (N_8450,N_3884,N_4356);
or U8451 (N_8451,N_2242,N_3083);
or U8452 (N_8452,N_928,N_4518);
nor U8453 (N_8453,N_3670,N_191);
and U8454 (N_8454,N_4998,N_3506);
and U8455 (N_8455,N_3327,N_4338);
and U8456 (N_8456,N_841,N_4725);
nor U8457 (N_8457,N_3782,N_2137);
or U8458 (N_8458,N_1433,N_3861);
or U8459 (N_8459,N_4153,N_2445);
and U8460 (N_8460,N_1371,N_2198);
and U8461 (N_8461,N_1798,N_750);
and U8462 (N_8462,N_3211,N_3835);
or U8463 (N_8463,N_1615,N_3725);
nand U8464 (N_8464,N_238,N_4734);
and U8465 (N_8465,N_4030,N_4016);
nor U8466 (N_8466,N_108,N_964);
nor U8467 (N_8467,N_2297,N_435);
nor U8468 (N_8468,N_2461,N_1537);
and U8469 (N_8469,N_601,N_2603);
or U8470 (N_8470,N_2123,N_1217);
nor U8471 (N_8471,N_1986,N_4168);
nand U8472 (N_8472,N_3218,N_3092);
and U8473 (N_8473,N_1655,N_3186);
nand U8474 (N_8474,N_1565,N_2241);
nor U8475 (N_8475,N_1309,N_2297);
or U8476 (N_8476,N_4448,N_2766);
or U8477 (N_8477,N_3718,N_4648);
nand U8478 (N_8478,N_2017,N_2738);
nand U8479 (N_8479,N_4598,N_1101);
nor U8480 (N_8480,N_975,N_2887);
xor U8481 (N_8481,N_287,N_610);
and U8482 (N_8482,N_3886,N_595);
or U8483 (N_8483,N_2024,N_2134);
nand U8484 (N_8484,N_3134,N_4798);
and U8485 (N_8485,N_2067,N_1575);
nand U8486 (N_8486,N_393,N_2937);
nor U8487 (N_8487,N_2119,N_1283);
nor U8488 (N_8488,N_1175,N_4903);
nor U8489 (N_8489,N_3417,N_3100);
and U8490 (N_8490,N_3796,N_1924);
and U8491 (N_8491,N_1915,N_1737);
or U8492 (N_8492,N_1610,N_3708);
and U8493 (N_8493,N_103,N_206);
nor U8494 (N_8494,N_3510,N_4888);
and U8495 (N_8495,N_1906,N_632);
nand U8496 (N_8496,N_3771,N_1855);
and U8497 (N_8497,N_1958,N_1069);
and U8498 (N_8498,N_2203,N_3237);
nor U8499 (N_8499,N_1016,N_2142);
nand U8500 (N_8500,N_1192,N_2580);
nand U8501 (N_8501,N_510,N_1905);
or U8502 (N_8502,N_2321,N_4651);
or U8503 (N_8503,N_726,N_2803);
nand U8504 (N_8504,N_2871,N_2607);
nand U8505 (N_8505,N_719,N_1533);
or U8506 (N_8506,N_4440,N_1157);
nor U8507 (N_8507,N_3203,N_1615);
or U8508 (N_8508,N_3976,N_98);
and U8509 (N_8509,N_1366,N_794);
and U8510 (N_8510,N_812,N_942);
nand U8511 (N_8511,N_1004,N_3935);
and U8512 (N_8512,N_2745,N_1790);
xnor U8513 (N_8513,N_2388,N_464);
and U8514 (N_8514,N_1275,N_4810);
or U8515 (N_8515,N_2856,N_2212);
or U8516 (N_8516,N_2533,N_986);
nor U8517 (N_8517,N_797,N_1931);
and U8518 (N_8518,N_2753,N_1787);
or U8519 (N_8519,N_3041,N_772);
and U8520 (N_8520,N_4328,N_3476);
nand U8521 (N_8521,N_4338,N_2130);
and U8522 (N_8522,N_1599,N_2526);
xor U8523 (N_8523,N_570,N_3213);
xor U8524 (N_8524,N_669,N_1728);
and U8525 (N_8525,N_3401,N_4789);
or U8526 (N_8526,N_140,N_3191);
or U8527 (N_8527,N_1706,N_1197);
and U8528 (N_8528,N_875,N_785);
nor U8529 (N_8529,N_2241,N_1543);
nand U8530 (N_8530,N_1822,N_2819);
or U8531 (N_8531,N_120,N_2872);
or U8532 (N_8532,N_400,N_4345);
nor U8533 (N_8533,N_2169,N_2288);
nor U8534 (N_8534,N_2845,N_1033);
and U8535 (N_8535,N_3363,N_826);
nand U8536 (N_8536,N_4254,N_3336);
or U8537 (N_8537,N_4318,N_3466);
nand U8538 (N_8538,N_3176,N_4762);
and U8539 (N_8539,N_2716,N_4963);
nand U8540 (N_8540,N_4527,N_2047);
or U8541 (N_8541,N_1156,N_765);
nand U8542 (N_8542,N_4119,N_4938);
and U8543 (N_8543,N_4686,N_4502);
or U8544 (N_8544,N_3726,N_554);
nor U8545 (N_8545,N_4543,N_3083);
nor U8546 (N_8546,N_1061,N_2225);
or U8547 (N_8547,N_64,N_3860);
and U8548 (N_8548,N_2748,N_1929);
and U8549 (N_8549,N_3221,N_2906);
xnor U8550 (N_8550,N_1607,N_1230);
nor U8551 (N_8551,N_4466,N_3503);
nand U8552 (N_8552,N_1316,N_319);
or U8553 (N_8553,N_1939,N_326);
nor U8554 (N_8554,N_2152,N_4139);
and U8555 (N_8555,N_1181,N_3847);
or U8556 (N_8556,N_1900,N_4456);
nor U8557 (N_8557,N_1172,N_503);
and U8558 (N_8558,N_1018,N_1105);
nand U8559 (N_8559,N_1179,N_1222);
and U8560 (N_8560,N_2557,N_1373);
and U8561 (N_8561,N_4585,N_3558);
nand U8562 (N_8562,N_913,N_437);
xnor U8563 (N_8563,N_4771,N_3484);
nor U8564 (N_8564,N_110,N_1090);
nor U8565 (N_8565,N_2866,N_3412);
nor U8566 (N_8566,N_1676,N_637);
or U8567 (N_8567,N_4733,N_1044);
nand U8568 (N_8568,N_604,N_4731);
nand U8569 (N_8569,N_4024,N_1341);
nor U8570 (N_8570,N_4592,N_2059);
or U8571 (N_8571,N_2218,N_1165);
and U8572 (N_8572,N_1674,N_3489);
nor U8573 (N_8573,N_3532,N_4197);
nor U8574 (N_8574,N_2709,N_4652);
or U8575 (N_8575,N_4933,N_2027);
and U8576 (N_8576,N_4740,N_1678);
nor U8577 (N_8577,N_1606,N_1434);
and U8578 (N_8578,N_695,N_1916);
or U8579 (N_8579,N_1161,N_4506);
and U8580 (N_8580,N_1450,N_2203);
or U8581 (N_8581,N_1018,N_803);
and U8582 (N_8582,N_4393,N_1748);
and U8583 (N_8583,N_4273,N_2946);
and U8584 (N_8584,N_4456,N_4627);
nand U8585 (N_8585,N_2386,N_1779);
nor U8586 (N_8586,N_572,N_1066);
or U8587 (N_8587,N_3734,N_978);
xor U8588 (N_8588,N_3061,N_3356);
and U8589 (N_8589,N_2374,N_1669);
nor U8590 (N_8590,N_3578,N_4344);
and U8591 (N_8591,N_1281,N_537);
nor U8592 (N_8592,N_2121,N_573);
and U8593 (N_8593,N_3182,N_709);
and U8594 (N_8594,N_948,N_2415);
nand U8595 (N_8595,N_3753,N_500);
nand U8596 (N_8596,N_1830,N_2503);
and U8597 (N_8597,N_2298,N_1849);
nand U8598 (N_8598,N_584,N_669);
nor U8599 (N_8599,N_3411,N_3892);
nor U8600 (N_8600,N_2461,N_3770);
and U8601 (N_8601,N_1283,N_1452);
nor U8602 (N_8602,N_4868,N_4871);
nand U8603 (N_8603,N_4012,N_463);
and U8604 (N_8604,N_1093,N_4674);
or U8605 (N_8605,N_1570,N_4767);
or U8606 (N_8606,N_154,N_2042);
and U8607 (N_8607,N_1072,N_219);
nand U8608 (N_8608,N_906,N_3901);
and U8609 (N_8609,N_2060,N_4434);
or U8610 (N_8610,N_2840,N_245);
nor U8611 (N_8611,N_2136,N_588);
or U8612 (N_8612,N_757,N_1404);
or U8613 (N_8613,N_4117,N_2049);
nor U8614 (N_8614,N_1755,N_3371);
nand U8615 (N_8615,N_4492,N_938);
xor U8616 (N_8616,N_1280,N_3693);
nand U8617 (N_8617,N_1964,N_355);
nor U8618 (N_8618,N_1960,N_2834);
nor U8619 (N_8619,N_4859,N_855);
nor U8620 (N_8620,N_4111,N_4652);
nand U8621 (N_8621,N_3810,N_1954);
or U8622 (N_8622,N_1271,N_4602);
nor U8623 (N_8623,N_4729,N_3540);
or U8624 (N_8624,N_4872,N_1288);
and U8625 (N_8625,N_2263,N_102);
nand U8626 (N_8626,N_1958,N_4133);
and U8627 (N_8627,N_4565,N_634);
nor U8628 (N_8628,N_1575,N_4212);
or U8629 (N_8629,N_1356,N_1927);
nor U8630 (N_8630,N_2058,N_2268);
and U8631 (N_8631,N_3259,N_663);
nand U8632 (N_8632,N_1897,N_2784);
or U8633 (N_8633,N_3034,N_2410);
or U8634 (N_8634,N_127,N_4291);
nand U8635 (N_8635,N_669,N_1730);
or U8636 (N_8636,N_1564,N_740);
and U8637 (N_8637,N_1535,N_3817);
and U8638 (N_8638,N_4005,N_2698);
nand U8639 (N_8639,N_4024,N_799);
nor U8640 (N_8640,N_4318,N_196);
nor U8641 (N_8641,N_3673,N_4545);
nor U8642 (N_8642,N_3287,N_59);
and U8643 (N_8643,N_872,N_2998);
nor U8644 (N_8644,N_953,N_3900);
and U8645 (N_8645,N_1412,N_1954);
nand U8646 (N_8646,N_492,N_3890);
nor U8647 (N_8647,N_1314,N_8);
and U8648 (N_8648,N_1496,N_1905);
nand U8649 (N_8649,N_791,N_234);
nor U8650 (N_8650,N_259,N_3300);
or U8651 (N_8651,N_4650,N_1934);
nand U8652 (N_8652,N_2408,N_3992);
nor U8653 (N_8653,N_546,N_2181);
nor U8654 (N_8654,N_100,N_4599);
or U8655 (N_8655,N_2827,N_738);
or U8656 (N_8656,N_2366,N_2866);
or U8657 (N_8657,N_1242,N_4452);
and U8658 (N_8658,N_2562,N_56);
nand U8659 (N_8659,N_3172,N_382);
or U8660 (N_8660,N_3484,N_4293);
and U8661 (N_8661,N_1374,N_2611);
nand U8662 (N_8662,N_4062,N_4206);
nor U8663 (N_8663,N_1388,N_2657);
or U8664 (N_8664,N_2485,N_1651);
or U8665 (N_8665,N_4745,N_1363);
or U8666 (N_8666,N_901,N_2157);
or U8667 (N_8667,N_4834,N_3032);
nor U8668 (N_8668,N_2029,N_4631);
nand U8669 (N_8669,N_3982,N_2128);
nand U8670 (N_8670,N_2403,N_3169);
nand U8671 (N_8671,N_1538,N_3260);
nand U8672 (N_8672,N_4160,N_4481);
nor U8673 (N_8673,N_1616,N_3467);
nor U8674 (N_8674,N_3766,N_2933);
or U8675 (N_8675,N_3213,N_3624);
and U8676 (N_8676,N_2311,N_737);
and U8677 (N_8677,N_238,N_137);
nand U8678 (N_8678,N_2673,N_1969);
or U8679 (N_8679,N_4930,N_3470);
or U8680 (N_8680,N_1190,N_4552);
or U8681 (N_8681,N_4367,N_1816);
and U8682 (N_8682,N_354,N_1235);
or U8683 (N_8683,N_984,N_4466);
nand U8684 (N_8684,N_3813,N_4907);
nand U8685 (N_8685,N_1458,N_4150);
nor U8686 (N_8686,N_3825,N_2965);
nor U8687 (N_8687,N_3961,N_4367);
nand U8688 (N_8688,N_4043,N_4432);
and U8689 (N_8689,N_1999,N_1816);
nor U8690 (N_8690,N_674,N_4383);
and U8691 (N_8691,N_261,N_4831);
nand U8692 (N_8692,N_4951,N_1908);
and U8693 (N_8693,N_98,N_2967);
or U8694 (N_8694,N_3776,N_4545);
or U8695 (N_8695,N_4992,N_3716);
nor U8696 (N_8696,N_4619,N_4294);
and U8697 (N_8697,N_862,N_249);
and U8698 (N_8698,N_3694,N_2823);
nand U8699 (N_8699,N_3644,N_4346);
nand U8700 (N_8700,N_61,N_407);
or U8701 (N_8701,N_694,N_3900);
nand U8702 (N_8702,N_1529,N_3930);
nand U8703 (N_8703,N_3776,N_290);
and U8704 (N_8704,N_1207,N_142);
nor U8705 (N_8705,N_2289,N_4796);
nor U8706 (N_8706,N_721,N_2241);
and U8707 (N_8707,N_4781,N_1238);
and U8708 (N_8708,N_3136,N_2270);
or U8709 (N_8709,N_3458,N_1003);
and U8710 (N_8710,N_3424,N_4160);
nor U8711 (N_8711,N_1492,N_262);
and U8712 (N_8712,N_2807,N_1639);
or U8713 (N_8713,N_775,N_353);
nor U8714 (N_8714,N_3577,N_3286);
nand U8715 (N_8715,N_4412,N_2205);
xor U8716 (N_8716,N_1353,N_2935);
nor U8717 (N_8717,N_739,N_1159);
and U8718 (N_8718,N_79,N_4362);
or U8719 (N_8719,N_4672,N_3306);
nor U8720 (N_8720,N_4777,N_3929);
nand U8721 (N_8721,N_239,N_434);
nor U8722 (N_8722,N_4147,N_1139);
xnor U8723 (N_8723,N_2806,N_3776);
or U8724 (N_8724,N_1448,N_3826);
nor U8725 (N_8725,N_3828,N_3390);
xor U8726 (N_8726,N_1309,N_3941);
or U8727 (N_8727,N_382,N_4026);
or U8728 (N_8728,N_1271,N_882);
or U8729 (N_8729,N_3015,N_3959);
nand U8730 (N_8730,N_3886,N_62);
or U8731 (N_8731,N_3403,N_958);
or U8732 (N_8732,N_421,N_4683);
nor U8733 (N_8733,N_775,N_2725);
or U8734 (N_8734,N_1566,N_1797);
and U8735 (N_8735,N_4725,N_43);
or U8736 (N_8736,N_4863,N_1322);
nand U8737 (N_8737,N_43,N_3271);
and U8738 (N_8738,N_882,N_1771);
or U8739 (N_8739,N_3601,N_2954);
nand U8740 (N_8740,N_1924,N_2182);
and U8741 (N_8741,N_4882,N_81);
and U8742 (N_8742,N_866,N_3615);
or U8743 (N_8743,N_92,N_504);
nand U8744 (N_8744,N_1977,N_3607);
and U8745 (N_8745,N_139,N_1332);
or U8746 (N_8746,N_1309,N_4718);
nor U8747 (N_8747,N_2941,N_811);
nor U8748 (N_8748,N_4688,N_1564);
and U8749 (N_8749,N_1089,N_1745);
nand U8750 (N_8750,N_1859,N_1024);
and U8751 (N_8751,N_1279,N_4025);
or U8752 (N_8752,N_4761,N_3562);
nand U8753 (N_8753,N_297,N_4209);
nor U8754 (N_8754,N_779,N_3513);
or U8755 (N_8755,N_949,N_4303);
nor U8756 (N_8756,N_2267,N_2439);
or U8757 (N_8757,N_2309,N_4701);
and U8758 (N_8758,N_4677,N_873);
and U8759 (N_8759,N_2299,N_3712);
nand U8760 (N_8760,N_1753,N_1651);
nand U8761 (N_8761,N_3834,N_2045);
or U8762 (N_8762,N_3213,N_1730);
nand U8763 (N_8763,N_3786,N_976);
xnor U8764 (N_8764,N_3110,N_1136);
nand U8765 (N_8765,N_670,N_2473);
and U8766 (N_8766,N_957,N_4573);
nand U8767 (N_8767,N_3050,N_2304);
nor U8768 (N_8768,N_4085,N_2672);
or U8769 (N_8769,N_3496,N_1083);
nor U8770 (N_8770,N_2138,N_1380);
nor U8771 (N_8771,N_3569,N_3208);
and U8772 (N_8772,N_156,N_4762);
nand U8773 (N_8773,N_2937,N_1005);
nor U8774 (N_8774,N_1892,N_1336);
nor U8775 (N_8775,N_4160,N_1769);
or U8776 (N_8776,N_1537,N_1300);
nor U8777 (N_8777,N_4048,N_3924);
and U8778 (N_8778,N_3613,N_3102);
nor U8779 (N_8779,N_4180,N_1513);
and U8780 (N_8780,N_1515,N_1268);
and U8781 (N_8781,N_4850,N_731);
xnor U8782 (N_8782,N_830,N_2217);
nand U8783 (N_8783,N_1776,N_4415);
nor U8784 (N_8784,N_229,N_2711);
or U8785 (N_8785,N_1416,N_1250);
nand U8786 (N_8786,N_4890,N_4812);
or U8787 (N_8787,N_3564,N_822);
or U8788 (N_8788,N_2581,N_2380);
nor U8789 (N_8789,N_2692,N_3196);
or U8790 (N_8790,N_3710,N_4302);
or U8791 (N_8791,N_3459,N_3664);
xor U8792 (N_8792,N_1049,N_1069);
nand U8793 (N_8793,N_3836,N_423);
nand U8794 (N_8794,N_1314,N_2051);
or U8795 (N_8795,N_1624,N_3928);
or U8796 (N_8796,N_4879,N_1406);
and U8797 (N_8797,N_4230,N_3537);
nand U8798 (N_8798,N_3929,N_1551);
and U8799 (N_8799,N_1407,N_1012);
and U8800 (N_8800,N_2324,N_4536);
nand U8801 (N_8801,N_1601,N_4486);
nor U8802 (N_8802,N_2976,N_4717);
nand U8803 (N_8803,N_4714,N_2126);
or U8804 (N_8804,N_3490,N_4401);
nor U8805 (N_8805,N_3921,N_3969);
nor U8806 (N_8806,N_3021,N_3651);
nand U8807 (N_8807,N_2128,N_3613);
and U8808 (N_8808,N_151,N_1644);
and U8809 (N_8809,N_2768,N_3798);
and U8810 (N_8810,N_1721,N_2388);
and U8811 (N_8811,N_4997,N_1442);
nand U8812 (N_8812,N_3499,N_3181);
or U8813 (N_8813,N_2751,N_2747);
or U8814 (N_8814,N_3837,N_3300);
nor U8815 (N_8815,N_1238,N_3439);
and U8816 (N_8816,N_2805,N_4119);
or U8817 (N_8817,N_4536,N_3457);
nand U8818 (N_8818,N_1607,N_4269);
or U8819 (N_8819,N_4246,N_1591);
nor U8820 (N_8820,N_984,N_238);
and U8821 (N_8821,N_4388,N_4334);
and U8822 (N_8822,N_2004,N_1924);
and U8823 (N_8823,N_2001,N_1392);
nor U8824 (N_8824,N_816,N_4779);
xnor U8825 (N_8825,N_4126,N_3509);
nand U8826 (N_8826,N_3546,N_2000);
nor U8827 (N_8827,N_3935,N_2359);
and U8828 (N_8828,N_2219,N_4646);
and U8829 (N_8829,N_3006,N_3460);
nor U8830 (N_8830,N_3760,N_249);
and U8831 (N_8831,N_4861,N_247);
or U8832 (N_8832,N_1686,N_252);
xnor U8833 (N_8833,N_1255,N_1395);
nand U8834 (N_8834,N_1190,N_2808);
nand U8835 (N_8835,N_2129,N_1794);
nor U8836 (N_8836,N_2312,N_4362);
nand U8837 (N_8837,N_3736,N_727);
nor U8838 (N_8838,N_2146,N_2372);
nand U8839 (N_8839,N_1143,N_2875);
nor U8840 (N_8840,N_849,N_4952);
nand U8841 (N_8841,N_4630,N_3488);
or U8842 (N_8842,N_794,N_870);
nand U8843 (N_8843,N_2679,N_2294);
or U8844 (N_8844,N_857,N_4992);
and U8845 (N_8845,N_1875,N_3413);
or U8846 (N_8846,N_2724,N_3314);
nand U8847 (N_8847,N_3635,N_2668);
nor U8848 (N_8848,N_4797,N_2876);
nand U8849 (N_8849,N_570,N_1367);
and U8850 (N_8850,N_3984,N_2474);
and U8851 (N_8851,N_1714,N_4211);
and U8852 (N_8852,N_3049,N_4611);
nor U8853 (N_8853,N_660,N_725);
and U8854 (N_8854,N_843,N_2611);
nor U8855 (N_8855,N_3428,N_4912);
and U8856 (N_8856,N_3137,N_2027);
and U8857 (N_8857,N_969,N_3954);
nor U8858 (N_8858,N_4346,N_255);
nor U8859 (N_8859,N_2185,N_2280);
nor U8860 (N_8860,N_4538,N_4382);
and U8861 (N_8861,N_1025,N_2914);
or U8862 (N_8862,N_1532,N_2751);
and U8863 (N_8863,N_2566,N_291);
nand U8864 (N_8864,N_2761,N_2105);
and U8865 (N_8865,N_4643,N_4654);
and U8866 (N_8866,N_3336,N_4387);
nor U8867 (N_8867,N_2283,N_3273);
nor U8868 (N_8868,N_2454,N_450);
and U8869 (N_8869,N_2374,N_1282);
or U8870 (N_8870,N_4770,N_3064);
and U8871 (N_8871,N_1993,N_100);
or U8872 (N_8872,N_2122,N_908);
xnor U8873 (N_8873,N_4159,N_2758);
or U8874 (N_8874,N_793,N_849);
nor U8875 (N_8875,N_189,N_4986);
nor U8876 (N_8876,N_2068,N_721);
nor U8877 (N_8877,N_3940,N_524);
and U8878 (N_8878,N_3997,N_2643);
nor U8879 (N_8879,N_3339,N_4209);
and U8880 (N_8880,N_1825,N_473);
and U8881 (N_8881,N_280,N_703);
and U8882 (N_8882,N_3813,N_2156);
nand U8883 (N_8883,N_676,N_3493);
or U8884 (N_8884,N_3926,N_4733);
or U8885 (N_8885,N_1008,N_3101);
nand U8886 (N_8886,N_3063,N_4488);
nand U8887 (N_8887,N_4298,N_4730);
or U8888 (N_8888,N_2206,N_4032);
nand U8889 (N_8889,N_1646,N_362);
or U8890 (N_8890,N_216,N_975);
and U8891 (N_8891,N_2215,N_261);
or U8892 (N_8892,N_3026,N_2408);
nor U8893 (N_8893,N_63,N_1647);
or U8894 (N_8894,N_2397,N_110);
nand U8895 (N_8895,N_2562,N_964);
nor U8896 (N_8896,N_2091,N_2684);
nand U8897 (N_8897,N_4370,N_3221);
and U8898 (N_8898,N_4807,N_1343);
or U8899 (N_8899,N_4262,N_3362);
nand U8900 (N_8900,N_419,N_2037);
or U8901 (N_8901,N_3717,N_1363);
nand U8902 (N_8902,N_576,N_3092);
or U8903 (N_8903,N_3464,N_2509);
or U8904 (N_8904,N_3896,N_1722);
or U8905 (N_8905,N_1298,N_3072);
nand U8906 (N_8906,N_4937,N_1996);
nor U8907 (N_8907,N_3949,N_2719);
or U8908 (N_8908,N_3534,N_629);
nand U8909 (N_8909,N_4086,N_4931);
nor U8910 (N_8910,N_3233,N_4956);
nand U8911 (N_8911,N_827,N_2947);
nand U8912 (N_8912,N_472,N_460);
nor U8913 (N_8913,N_2178,N_3655);
nor U8914 (N_8914,N_4485,N_3844);
or U8915 (N_8915,N_2609,N_1742);
nor U8916 (N_8916,N_3168,N_4032);
nand U8917 (N_8917,N_4723,N_4833);
nand U8918 (N_8918,N_759,N_541);
nor U8919 (N_8919,N_708,N_4317);
and U8920 (N_8920,N_1380,N_673);
nand U8921 (N_8921,N_4591,N_3765);
nor U8922 (N_8922,N_156,N_3309);
and U8923 (N_8923,N_4346,N_1517);
and U8924 (N_8924,N_4472,N_4702);
nand U8925 (N_8925,N_3919,N_4604);
xor U8926 (N_8926,N_3401,N_3239);
or U8927 (N_8927,N_4515,N_4366);
or U8928 (N_8928,N_2363,N_279);
and U8929 (N_8929,N_4467,N_3449);
and U8930 (N_8930,N_597,N_549);
nor U8931 (N_8931,N_4968,N_3823);
nor U8932 (N_8932,N_4738,N_768);
and U8933 (N_8933,N_3018,N_3615);
and U8934 (N_8934,N_2175,N_2524);
xor U8935 (N_8935,N_1932,N_756);
nand U8936 (N_8936,N_2617,N_1697);
and U8937 (N_8937,N_1346,N_838);
nor U8938 (N_8938,N_4244,N_1477);
nor U8939 (N_8939,N_839,N_2946);
or U8940 (N_8940,N_671,N_994);
nand U8941 (N_8941,N_2226,N_4021);
nand U8942 (N_8942,N_3002,N_1985);
nor U8943 (N_8943,N_4154,N_608);
and U8944 (N_8944,N_3156,N_4270);
or U8945 (N_8945,N_3503,N_4742);
or U8946 (N_8946,N_979,N_3035);
and U8947 (N_8947,N_4113,N_3835);
nor U8948 (N_8948,N_4819,N_2498);
nand U8949 (N_8949,N_4650,N_3646);
xor U8950 (N_8950,N_2872,N_1562);
nor U8951 (N_8951,N_3567,N_670);
nand U8952 (N_8952,N_1570,N_3264);
nand U8953 (N_8953,N_402,N_940);
and U8954 (N_8954,N_1738,N_139);
nor U8955 (N_8955,N_3529,N_2946);
or U8956 (N_8956,N_2965,N_1368);
nor U8957 (N_8957,N_3964,N_503);
and U8958 (N_8958,N_4633,N_3186);
or U8959 (N_8959,N_4307,N_748);
and U8960 (N_8960,N_1898,N_1765);
nor U8961 (N_8961,N_2013,N_1118);
nand U8962 (N_8962,N_2155,N_1879);
or U8963 (N_8963,N_1804,N_3497);
or U8964 (N_8964,N_3903,N_1255);
or U8965 (N_8965,N_2070,N_591);
or U8966 (N_8966,N_583,N_2836);
or U8967 (N_8967,N_869,N_2245);
nand U8968 (N_8968,N_1169,N_3138);
nand U8969 (N_8969,N_1965,N_2729);
or U8970 (N_8970,N_3853,N_801);
and U8971 (N_8971,N_1513,N_1173);
xor U8972 (N_8972,N_807,N_99);
and U8973 (N_8973,N_1473,N_2992);
nand U8974 (N_8974,N_4025,N_2223);
nor U8975 (N_8975,N_1829,N_1673);
nand U8976 (N_8976,N_816,N_2645);
or U8977 (N_8977,N_2445,N_4771);
nor U8978 (N_8978,N_4601,N_4720);
nor U8979 (N_8979,N_1247,N_1534);
xor U8980 (N_8980,N_4463,N_2169);
or U8981 (N_8981,N_2799,N_2595);
and U8982 (N_8982,N_4880,N_1373);
nand U8983 (N_8983,N_440,N_2994);
nand U8984 (N_8984,N_206,N_1525);
nor U8985 (N_8985,N_528,N_2991);
nor U8986 (N_8986,N_1960,N_2900);
or U8987 (N_8987,N_2803,N_3174);
nand U8988 (N_8988,N_4198,N_2232);
or U8989 (N_8989,N_1754,N_4448);
nor U8990 (N_8990,N_2086,N_2566);
nor U8991 (N_8991,N_3377,N_3803);
nor U8992 (N_8992,N_3270,N_1075);
nand U8993 (N_8993,N_1253,N_2588);
and U8994 (N_8994,N_3672,N_2871);
nor U8995 (N_8995,N_973,N_4888);
and U8996 (N_8996,N_98,N_4313);
nand U8997 (N_8997,N_75,N_2203);
and U8998 (N_8998,N_3667,N_4967);
or U8999 (N_8999,N_1663,N_4725);
nor U9000 (N_9000,N_3584,N_801);
nand U9001 (N_9001,N_2031,N_4552);
nand U9002 (N_9002,N_3246,N_1687);
and U9003 (N_9003,N_3683,N_2890);
or U9004 (N_9004,N_2848,N_1552);
and U9005 (N_9005,N_3357,N_3486);
and U9006 (N_9006,N_2719,N_4759);
nor U9007 (N_9007,N_512,N_210);
and U9008 (N_9008,N_1262,N_1491);
and U9009 (N_9009,N_3294,N_3811);
nand U9010 (N_9010,N_203,N_2672);
nand U9011 (N_9011,N_3779,N_3715);
and U9012 (N_9012,N_44,N_4065);
and U9013 (N_9013,N_3275,N_1196);
nand U9014 (N_9014,N_3649,N_4969);
nand U9015 (N_9015,N_3901,N_4306);
nor U9016 (N_9016,N_158,N_367);
nor U9017 (N_9017,N_820,N_307);
and U9018 (N_9018,N_4561,N_3731);
xnor U9019 (N_9019,N_4048,N_4288);
and U9020 (N_9020,N_2605,N_1409);
and U9021 (N_9021,N_3842,N_2259);
xnor U9022 (N_9022,N_2904,N_1534);
nor U9023 (N_9023,N_853,N_4228);
and U9024 (N_9024,N_3606,N_2823);
and U9025 (N_9025,N_2975,N_4910);
or U9026 (N_9026,N_4514,N_2852);
nand U9027 (N_9027,N_4749,N_1154);
nand U9028 (N_9028,N_3846,N_1119);
nand U9029 (N_9029,N_2572,N_365);
nand U9030 (N_9030,N_1069,N_2035);
nor U9031 (N_9031,N_1629,N_1954);
or U9032 (N_9032,N_987,N_1379);
and U9033 (N_9033,N_4196,N_4802);
or U9034 (N_9034,N_475,N_3758);
nand U9035 (N_9035,N_3089,N_3611);
nor U9036 (N_9036,N_976,N_3791);
nor U9037 (N_9037,N_1545,N_725);
nor U9038 (N_9038,N_1319,N_4152);
nor U9039 (N_9039,N_4453,N_4445);
nand U9040 (N_9040,N_149,N_1766);
and U9041 (N_9041,N_136,N_3791);
and U9042 (N_9042,N_589,N_2896);
nor U9043 (N_9043,N_3856,N_2137);
nor U9044 (N_9044,N_2768,N_4776);
nor U9045 (N_9045,N_3778,N_3156);
and U9046 (N_9046,N_4651,N_217);
nand U9047 (N_9047,N_3688,N_105);
nor U9048 (N_9048,N_2422,N_3139);
and U9049 (N_9049,N_4462,N_1075);
nand U9050 (N_9050,N_4507,N_4368);
nand U9051 (N_9051,N_394,N_2465);
nand U9052 (N_9052,N_2169,N_826);
and U9053 (N_9053,N_1722,N_4574);
or U9054 (N_9054,N_4762,N_2306);
or U9055 (N_9055,N_4226,N_1141);
or U9056 (N_9056,N_1598,N_2572);
nor U9057 (N_9057,N_763,N_4127);
nand U9058 (N_9058,N_808,N_395);
and U9059 (N_9059,N_4102,N_2146);
nand U9060 (N_9060,N_4523,N_29);
and U9061 (N_9061,N_133,N_1381);
nor U9062 (N_9062,N_974,N_546);
or U9063 (N_9063,N_1006,N_1428);
and U9064 (N_9064,N_222,N_4543);
or U9065 (N_9065,N_2705,N_3460);
nand U9066 (N_9066,N_4895,N_2090);
nand U9067 (N_9067,N_1129,N_1383);
or U9068 (N_9068,N_2381,N_4274);
nand U9069 (N_9069,N_3856,N_2342);
or U9070 (N_9070,N_3916,N_198);
or U9071 (N_9071,N_4138,N_130);
and U9072 (N_9072,N_1500,N_3999);
and U9073 (N_9073,N_2521,N_91);
and U9074 (N_9074,N_853,N_2299);
and U9075 (N_9075,N_1681,N_387);
nand U9076 (N_9076,N_4702,N_4809);
nand U9077 (N_9077,N_1562,N_4899);
or U9078 (N_9078,N_2323,N_2457);
and U9079 (N_9079,N_4576,N_549);
or U9080 (N_9080,N_2888,N_3274);
or U9081 (N_9081,N_4071,N_2624);
nor U9082 (N_9082,N_2578,N_3030);
or U9083 (N_9083,N_1977,N_1483);
and U9084 (N_9084,N_2980,N_1967);
nand U9085 (N_9085,N_1804,N_339);
and U9086 (N_9086,N_4254,N_3543);
nor U9087 (N_9087,N_363,N_572);
nand U9088 (N_9088,N_1381,N_2201);
nor U9089 (N_9089,N_889,N_2987);
nand U9090 (N_9090,N_1181,N_2273);
or U9091 (N_9091,N_3201,N_1570);
or U9092 (N_9092,N_3421,N_2717);
nor U9093 (N_9093,N_204,N_869);
and U9094 (N_9094,N_2242,N_2891);
or U9095 (N_9095,N_4629,N_3303);
and U9096 (N_9096,N_624,N_3684);
and U9097 (N_9097,N_3976,N_4248);
xnor U9098 (N_9098,N_2284,N_2074);
and U9099 (N_9099,N_3015,N_1344);
and U9100 (N_9100,N_4731,N_4389);
and U9101 (N_9101,N_3171,N_3744);
and U9102 (N_9102,N_883,N_3387);
nand U9103 (N_9103,N_3635,N_4184);
nor U9104 (N_9104,N_1047,N_2973);
or U9105 (N_9105,N_490,N_3989);
xor U9106 (N_9106,N_4263,N_3870);
nor U9107 (N_9107,N_2332,N_4596);
nor U9108 (N_9108,N_4507,N_2330);
or U9109 (N_9109,N_4832,N_767);
or U9110 (N_9110,N_2450,N_2672);
nand U9111 (N_9111,N_2200,N_4969);
or U9112 (N_9112,N_4344,N_4191);
or U9113 (N_9113,N_4050,N_3899);
and U9114 (N_9114,N_1100,N_3913);
or U9115 (N_9115,N_4941,N_2273);
nor U9116 (N_9116,N_2233,N_1811);
xor U9117 (N_9117,N_1428,N_373);
or U9118 (N_9118,N_171,N_803);
or U9119 (N_9119,N_1880,N_2753);
xnor U9120 (N_9120,N_2568,N_312);
nand U9121 (N_9121,N_1285,N_839);
nor U9122 (N_9122,N_378,N_2582);
nand U9123 (N_9123,N_1554,N_3521);
xor U9124 (N_9124,N_1518,N_2512);
or U9125 (N_9125,N_257,N_2246);
nand U9126 (N_9126,N_1044,N_491);
and U9127 (N_9127,N_4207,N_836);
nand U9128 (N_9128,N_3438,N_3718);
nor U9129 (N_9129,N_2951,N_2014);
nor U9130 (N_9130,N_3563,N_2174);
nor U9131 (N_9131,N_1387,N_3975);
or U9132 (N_9132,N_3019,N_3264);
and U9133 (N_9133,N_1226,N_2788);
and U9134 (N_9134,N_1284,N_3527);
or U9135 (N_9135,N_3145,N_3201);
or U9136 (N_9136,N_2357,N_590);
nand U9137 (N_9137,N_2483,N_506);
or U9138 (N_9138,N_4092,N_3400);
nand U9139 (N_9139,N_4875,N_1352);
nor U9140 (N_9140,N_4948,N_4625);
nand U9141 (N_9141,N_3166,N_4128);
nor U9142 (N_9142,N_1631,N_3968);
and U9143 (N_9143,N_3194,N_3467);
or U9144 (N_9144,N_509,N_4606);
and U9145 (N_9145,N_1944,N_843);
nand U9146 (N_9146,N_5,N_245);
or U9147 (N_9147,N_4877,N_261);
nand U9148 (N_9148,N_1474,N_2385);
nor U9149 (N_9149,N_3814,N_1757);
or U9150 (N_9150,N_3456,N_4664);
nor U9151 (N_9151,N_4387,N_4201);
nor U9152 (N_9152,N_4249,N_1307);
or U9153 (N_9153,N_949,N_1962);
or U9154 (N_9154,N_2788,N_4126);
nor U9155 (N_9155,N_2789,N_2955);
nor U9156 (N_9156,N_2427,N_513);
or U9157 (N_9157,N_3916,N_1310);
nor U9158 (N_9158,N_796,N_1348);
nand U9159 (N_9159,N_763,N_4436);
and U9160 (N_9160,N_2483,N_4554);
nor U9161 (N_9161,N_1289,N_296);
or U9162 (N_9162,N_1247,N_4165);
nor U9163 (N_9163,N_649,N_4385);
and U9164 (N_9164,N_3815,N_243);
and U9165 (N_9165,N_481,N_2112);
nor U9166 (N_9166,N_307,N_180);
and U9167 (N_9167,N_3648,N_2900);
nand U9168 (N_9168,N_4075,N_4264);
and U9169 (N_9169,N_3468,N_4398);
and U9170 (N_9170,N_1123,N_861);
nor U9171 (N_9171,N_3431,N_1608);
and U9172 (N_9172,N_3096,N_4449);
and U9173 (N_9173,N_583,N_3594);
nor U9174 (N_9174,N_969,N_345);
and U9175 (N_9175,N_949,N_2187);
nor U9176 (N_9176,N_3845,N_4767);
or U9177 (N_9177,N_4204,N_932);
nor U9178 (N_9178,N_4731,N_3494);
nor U9179 (N_9179,N_3531,N_887);
nor U9180 (N_9180,N_3815,N_2641);
nor U9181 (N_9181,N_276,N_1702);
nand U9182 (N_9182,N_814,N_4020);
and U9183 (N_9183,N_1291,N_2957);
nand U9184 (N_9184,N_2505,N_1427);
nand U9185 (N_9185,N_4197,N_4868);
nor U9186 (N_9186,N_3351,N_3752);
and U9187 (N_9187,N_4946,N_3328);
nand U9188 (N_9188,N_2857,N_2871);
or U9189 (N_9189,N_495,N_3250);
nand U9190 (N_9190,N_2889,N_1999);
or U9191 (N_9191,N_137,N_4021);
nand U9192 (N_9192,N_2249,N_4837);
nor U9193 (N_9193,N_539,N_2311);
nor U9194 (N_9194,N_310,N_4531);
nor U9195 (N_9195,N_4398,N_3150);
or U9196 (N_9196,N_317,N_4330);
and U9197 (N_9197,N_4977,N_1230);
or U9198 (N_9198,N_2143,N_2723);
nor U9199 (N_9199,N_4812,N_2227);
or U9200 (N_9200,N_1166,N_3812);
nor U9201 (N_9201,N_64,N_4758);
xnor U9202 (N_9202,N_753,N_4373);
nand U9203 (N_9203,N_4164,N_3912);
nor U9204 (N_9204,N_4850,N_1528);
or U9205 (N_9205,N_4180,N_664);
and U9206 (N_9206,N_688,N_1089);
nand U9207 (N_9207,N_1468,N_857);
xor U9208 (N_9208,N_3845,N_1753);
nand U9209 (N_9209,N_4978,N_289);
and U9210 (N_9210,N_3872,N_2155);
and U9211 (N_9211,N_4715,N_366);
nand U9212 (N_9212,N_2267,N_1041);
nand U9213 (N_9213,N_582,N_4402);
and U9214 (N_9214,N_2246,N_688);
and U9215 (N_9215,N_390,N_2437);
nand U9216 (N_9216,N_303,N_2043);
nor U9217 (N_9217,N_1620,N_2578);
nand U9218 (N_9218,N_3304,N_2416);
nor U9219 (N_9219,N_3103,N_2990);
nor U9220 (N_9220,N_4890,N_1228);
and U9221 (N_9221,N_4975,N_3170);
and U9222 (N_9222,N_226,N_3901);
nand U9223 (N_9223,N_2308,N_2420);
or U9224 (N_9224,N_4898,N_2502);
nand U9225 (N_9225,N_3008,N_4311);
or U9226 (N_9226,N_936,N_4553);
and U9227 (N_9227,N_356,N_4882);
and U9228 (N_9228,N_2275,N_4385);
and U9229 (N_9229,N_2036,N_4298);
nor U9230 (N_9230,N_4706,N_4513);
nor U9231 (N_9231,N_3807,N_574);
nor U9232 (N_9232,N_4345,N_147);
nand U9233 (N_9233,N_3335,N_3468);
and U9234 (N_9234,N_275,N_1990);
nand U9235 (N_9235,N_2571,N_4898);
nor U9236 (N_9236,N_319,N_2133);
nor U9237 (N_9237,N_4784,N_4749);
and U9238 (N_9238,N_3545,N_2047);
or U9239 (N_9239,N_4397,N_4876);
nor U9240 (N_9240,N_1552,N_1135);
or U9241 (N_9241,N_1160,N_2352);
nand U9242 (N_9242,N_1328,N_4025);
nor U9243 (N_9243,N_1819,N_3244);
or U9244 (N_9244,N_3841,N_1337);
or U9245 (N_9245,N_3616,N_3601);
and U9246 (N_9246,N_4623,N_4978);
or U9247 (N_9247,N_2784,N_61);
nor U9248 (N_9248,N_3585,N_2612);
or U9249 (N_9249,N_555,N_3589);
nand U9250 (N_9250,N_4947,N_631);
nor U9251 (N_9251,N_3713,N_1472);
nor U9252 (N_9252,N_872,N_2180);
nand U9253 (N_9253,N_2090,N_463);
nor U9254 (N_9254,N_1606,N_1603);
nand U9255 (N_9255,N_4337,N_4787);
xnor U9256 (N_9256,N_23,N_2213);
or U9257 (N_9257,N_2187,N_653);
xnor U9258 (N_9258,N_4030,N_3327);
and U9259 (N_9259,N_2638,N_2703);
nor U9260 (N_9260,N_2970,N_4310);
nor U9261 (N_9261,N_3724,N_4968);
nor U9262 (N_9262,N_518,N_773);
nor U9263 (N_9263,N_220,N_4374);
nor U9264 (N_9264,N_4581,N_1682);
xnor U9265 (N_9265,N_2285,N_3508);
or U9266 (N_9266,N_838,N_4783);
or U9267 (N_9267,N_4731,N_3755);
nor U9268 (N_9268,N_3650,N_2271);
and U9269 (N_9269,N_2754,N_4078);
or U9270 (N_9270,N_142,N_2079);
xor U9271 (N_9271,N_1685,N_1517);
or U9272 (N_9272,N_4895,N_566);
or U9273 (N_9273,N_3311,N_4135);
or U9274 (N_9274,N_2651,N_3095);
nand U9275 (N_9275,N_3067,N_3894);
or U9276 (N_9276,N_1993,N_1947);
nand U9277 (N_9277,N_950,N_1874);
or U9278 (N_9278,N_674,N_603);
nor U9279 (N_9279,N_1823,N_1610);
nor U9280 (N_9280,N_4220,N_3021);
and U9281 (N_9281,N_2641,N_2501);
nand U9282 (N_9282,N_4667,N_1826);
or U9283 (N_9283,N_105,N_2060);
nor U9284 (N_9284,N_366,N_4134);
nor U9285 (N_9285,N_2116,N_2337);
nand U9286 (N_9286,N_3120,N_4011);
nor U9287 (N_9287,N_1145,N_4545);
xnor U9288 (N_9288,N_242,N_4439);
nand U9289 (N_9289,N_494,N_2366);
nand U9290 (N_9290,N_3857,N_3006);
nand U9291 (N_9291,N_2316,N_4288);
nor U9292 (N_9292,N_1464,N_1357);
nand U9293 (N_9293,N_537,N_2700);
nand U9294 (N_9294,N_1667,N_880);
or U9295 (N_9295,N_4707,N_2470);
or U9296 (N_9296,N_2399,N_1991);
or U9297 (N_9297,N_1636,N_3198);
or U9298 (N_9298,N_2832,N_4544);
nor U9299 (N_9299,N_1709,N_136);
nor U9300 (N_9300,N_2382,N_3591);
or U9301 (N_9301,N_4863,N_932);
xnor U9302 (N_9302,N_4330,N_1315);
nor U9303 (N_9303,N_1604,N_3147);
nand U9304 (N_9304,N_2134,N_4622);
and U9305 (N_9305,N_1041,N_1543);
and U9306 (N_9306,N_3703,N_2481);
and U9307 (N_9307,N_3418,N_3648);
nand U9308 (N_9308,N_1208,N_3219);
and U9309 (N_9309,N_1944,N_3465);
and U9310 (N_9310,N_3083,N_1700);
or U9311 (N_9311,N_4657,N_1401);
nor U9312 (N_9312,N_402,N_3738);
or U9313 (N_9313,N_853,N_4423);
nand U9314 (N_9314,N_3352,N_3486);
or U9315 (N_9315,N_3192,N_1434);
and U9316 (N_9316,N_2639,N_2846);
nor U9317 (N_9317,N_3447,N_2751);
and U9318 (N_9318,N_2573,N_2837);
nor U9319 (N_9319,N_2938,N_3901);
or U9320 (N_9320,N_1260,N_798);
and U9321 (N_9321,N_1903,N_285);
or U9322 (N_9322,N_2064,N_1789);
and U9323 (N_9323,N_2867,N_3185);
nand U9324 (N_9324,N_102,N_2436);
nand U9325 (N_9325,N_4271,N_4624);
or U9326 (N_9326,N_3798,N_3132);
and U9327 (N_9327,N_1282,N_1501);
nand U9328 (N_9328,N_124,N_3375);
nand U9329 (N_9329,N_1182,N_3034);
or U9330 (N_9330,N_3846,N_1775);
nor U9331 (N_9331,N_3626,N_1219);
and U9332 (N_9332,N_193,N_3330);
nor U9333 (N_9333,N_1255,N_558);
nand U9334 (N_9334,N_2294,N_4957);
and U9335 (N_9335,N_3679,N_1747);
nand U9336 (N_9336,N_879,N_106);
nor U9337 (N_9337,N_3707,N_4903);
and U9338 (N_9338,N_4309,N_446);
nor U9339 (N_9339,N_3119,N_1117);
nand U9340 (N_9340,N_2540,N_3343);
and U9341 (N_9341,N_3170,N_106);
or U9342 (N_9342,N_286,N_4567);
or U9343 (N_9343,N_4549,N_1097);
and U9344 (N_9344,N_974,N_126);
nand U9345 (N_9345,N_4769,N_2045);
xnor U9346 (N_9346,N_4379,N_3627);
or U9347 (N_9347,N_1981,N_1257);
or U9348 (N_9348,N_753,N_4937);
nand U9349 (N_9349,N_1859,N_4129);
nor U9350 (N_9350,N_2516,N_3580);
and U9351 (N_9351,N_3050,N_1788);
and U9352 (N_9352,N_2209,N_880);
nand U9353 (N_9353,N_4412,N_3165);
or U9354 (N_9354,N_1010,N_2598);
and U9355 (N_9355,N_2469,N_1542);
or U9356 (N_9356,N_697,N_771);
or U9357 (N_9357,N_4893,N_4054);
nand U9358 (N_9358,N_2596,N_3243);
nor U9359 (N_9359,N_4946,N_3532);
or U9360 (N_9360,N_1790,N_3364);
xor U9361 (N_9361,N_1700,N_3090);
or U9362 (N_9362,N_2044,N_193);
and U9363 (N_9363,N_3554,N_3327);
or U9364 (N_9364,N_3867,N_2300);
and U9365 (N_9365,N_2229,N_707);
nand U9366 (N_9366,N_4422,N_2533);
or U9367 (N_9367,N_2893,N_4882);
or U9368 (N_9368,N_2092,N_3960);
xor U9369 (N_9369,N_2283,N_4326);
nand U9370 (N_9370,N_4604,N_3237);
or U9371 (N_9371,N_2579,N_1218);
nand U9372 (N_9372,N_3492,N_1609);
and U9373 (N_9373,N_3800,N_3771);
nand U9374 (N_9374,N_1461,N_2606);
nand U9375 (N_9375,N_2050,N_2979);
or U9376 (N_9376,N_3437,N_4839);
nor U9377 (N_9377,N_4610,N_3888);
or U9378 (N_9378,N_1763,N_3438);
and U9379 (N_9379,N_4656,N_3776);
nand U9380 (N_9380,N_4480,N_4599);
or U9381 (N_9381,N_1210,N_4576);
nand U9382 (N_9382,N_812,N_1039);
and U9383 (N_9383,N_4833,N_599);
nand U9384 (N_9384,N_817,N_547);
or U9385 (N_9385,N_4181,N_3515);
nand U9386 (N_9386,N_1550,N_730);
and U9387 (N_9387,N_3864,N_1432);
or U9388 (N_9388,N_4871,N_4435);
or U9389 (N_9389,N_4033,N_4280);
nor U9390 (N_9390,N_3996,N_1833);
nand U9391 (N_9391,N_4825,N_805);
or U9392 (N_9392,N_870,N_2586);
and U9393 (N_9393,N_1968,N_3841);
nand U9394 (N_9394,N_3853,N_4632);
nand U9395 (N_9395,N_320,N_2971);
or U9396 (N_9396,N_1666,N_1704);
nand U9397 (N_9397,N_840,N_2373);
or U9398 (N_9398,N_1211,N_2355);
nor U9399 (N_9399,N_612,N_1001);
and U9400 (N_9400,N_4066,N_3934);
xnor U9401 (N_9401,N_740,N_1781);
nand U9402 (N_9402,N_2452,N_1176);
nor U9403 (N_9403,N_4774,N_2731);
or U9404 (N_9404,N_3374,N_3567);
xor U9405 (N_9405,N_4001,N_1516);
and U9406 (N_9406,N_702,N_3161);
or U9407 (N_9407,N_1840,N_649);
or U9408 (N_9408,N_4510,N_2124);
nor U9409 (N_9409,N_2441,N_2722);
and U9410 (N_9410,N_921,N_559);
or U9411 (N_9411,N_4212,N_717);
nand U9412 (N_9412,N_1787,N_4233);
nor U9413 (N_9413,N_553,N_2030);
or U9414 (N_9414,N_4250,N_3816);
or U9415 (N_9415,N_4954,N_4744);
and U9416 (N_9416,N_3379,N_344);
nand U9417 (N_9417,N_68,N_689);
nor U9418 (N_9418,N_2253,N_4206);
nor U9419 (N_9419,N_3300,N_926);
nand U9420 (N_9420,N_1367,N_4145);
nor U9421 (N_9421,N_4265,N_2748);
nand U9422 (N_9422,N_2731,N_606);
or U9423 (N_9423,N_3567,N_82);
nand U9424 (N_9424,N_4584,N_1650);
nor U9425 (N_9425,N_4385,N_512);
and U9426 (N_9426,N_3713,N_1358);
and U9427 (N_9427,N_586,N_2082);
and U9428 (N_9428,N_144,N_3772);
and U9429 (N_9429,N_2995,N_2894);
nand U9430 (N_9430,N_1508,N_917);
or U9431 (N_9431,N_3784,N_3475);
and U9432 (N_9432,N_1125,N_1084);
and U9433 (N_9433,N_2419,N_3355);
and U9434 (N_9434,N_3343,N_2442);
nor U9435 (N_9435,N_952,N_2116);
nor U9436 (N_9436,N_3907,N_4427);
nand U9437 (N_9437,N_1332,N_462);
nand U9438 (N_9438,N_2267,N_4914);
and U9439 (N_9439,N_1912,N_2418);
and U9440 (N_9440,N_3302,N_1977);
nand U9441 (N_9441,N_1975,N_514);
nor U9442 (N_9442,N_1192,N_4110);
nor U9443 (N_9443,N_1466,N_3069);
or U9444 (N_9444,N_4051,N_1577);
nand U9445 (N_9445,N_2802,N_3899);
and U9446 (N_9446,N_2726,N_2521);
nor U9447 (N_9447,N_2406,N_3373);
nand U9448 (N_9448,N_939,N_114);
or U9449 (N_9449,N_1327,N_3897);
nor U9450 (N_9450,N_1429,N_628);
and U9451 (N_9451,N_471,N_1404);
or U9452 (N_9452,N_579,N_4436);
or U9453 (N_9453,N_681,N_3408);
or U9454 (N_9454,N_3159,N_392);
and U9455 (N_9455,N_1892,N_447);
and U9456 (N_9456,N_2883,N_1752);
nor U9457 (N_9457,N_1114,N_2700);
xor U9458 (N_9458,N_4666,N_4171);
nand U9459 (N_9459,N_2471,N_1490);
or U9460 (N_9460,N_3102,N_655);
nand U9461 (N_9461,N_894,N_1938);
nand U9462 (N_9462,N_1648,N_3574);
nor U9463 (N_9463,N_955,N_2861);
nor U9464 (N_9464,N_4766,N_2401);
nand U9465 (N_9465,N_2915,N_2498);
or U9466 (N_9466,N_2431,N_174);
nand U9467 (N_9467,N_155,N_4442);
nand U9468 (N_9468,N_4487,N_4199);
nand U9469 (N_9469,N_401,N_3210);
and U9470 (N_9470,N_2657,N_1182);
nor U9471 (N_9471,N_2468,N_279);
or U9472 (N_9472,N_4491,N_1691);
and U9473 (N_9473,N_2129,N_2784);
and U9474 (N_9474,N_4369,N_982);
and U9475 (N_9475,N_641,N_2243);
nor U9476 (N_9476,N_1786,N_4978);
or U9477 (N_9477,N_3285,N_606);
nand U9478 (N_9478,N_1800,N_1265);
or U9479 (N_9479,N_3736,N_3525);
or U9480 (N_9480,N_3823,N_4374);
or U9481 (N_9481,N_4871,N_669);
and U9482 (N_9482,N_3921,N_3033);
xor U9483 (N_9483,N_4419,N_965);
and U9484 (N_9484,N_3088,N_1342);
or U9485 (N_9485,N_4782,N_1185);
nor U9486 (N_9486,N_685,N_1703);
nor U9487 (N_9487,N_3346,N_676);
nand U9488 (N_9488,N_1776,N_1780);
and U9489 (N_9489,N_209,N_833);
nand U9490 (N_9490,N_702,N_3830);
nand U9491 (N_9491,N_3623,N_4463);
and U9492 (N_9492,N_396,N_4542);
and U9493 (N_9493,N_4813,N_1052);
nor U9494 (N_9494,N_3066,N_4771);
or U9495 (N_9495,N_1846,N_1568);
nor U9496 (N_9496,N_888,N_3656);
nor U9497 (N_9497,N_858,N_3120);
or U9498 (N_9498,N_386,N_411);
nand U9499 (N_9499,N_2936,N_4534);
nand U9500 (N_9500,N_1090,N_3054);
and U9501 (N_9501,N_814,N_341);
xnor U9502 (N_9502,N_245,N_1540);
nand U9503 (N_9503,N_282,N_1292);
nand U9504 (N_9504,N_2850,N_1233);
nor U9505 (N_9505,N_744,N_1860);
or U9506 (N_9506,N_4671,N_1838);
nand U9507 (N_9507,N_210,N_3960);
and U9508 (N_9508,N_710,N_4505);
and U9509 (N_9509,N_3114,N_3896);
and U9510 (N_9510,N_2514,N_1457);
or U9511 (N_9511,N_23,N_3772);
nand U9512 (N_9512,N_3845,N_2397);
nor U9513 (N_9513,N_3399,N_3884);
and U9514 (N_9514,N_2233,N_2640);
and U9515 (N_9515,N_1180,N_736);
nand U9516 (N_9516,N_2051,N_4243);
or U9517 (N_9517,N_2518,N_1612);
nand U9518 (N_9518,N_1374,N_555);
nand U9519 (N_9519,N_1377,N_3753);
nor U9520 (N_9520,N_2971,N_4789);
and U9521 (N_9521,N_2867,N_472);
nand U9522 (N_9522,N_4858,N_371);
or U9523 (N_9523,N_2692,N_4052);
nand U9524 (N_9524,N_721,N_527);
or U9525 (N_9525,N_1347,N_2802);
or U9526 (N_9526,N_1183,N_4493);
nor U9527 (N_9527,N_3726,N_3143);
xor U9528 (N_9528,N_4571,N_4809);
or U9529 (N_9529,N_2669,N_3562);
nor U9530 (N_9530,N_4706,N_357);
or U9531 (N_9531,N_2393,N_2342);
nor U9532 (N_9532,N_967,N_593);
nor U9533 (N_9533,N_614,N_1491);
and U9534 (N_9534,N_4608,N_2765);
nor U9535 (N_9535,N_1391,N_3637);
nor U9536 (N_9536,N_116,N_2089);
xor U9537 (N_9537,N_4026,N_1819);
or U9538 (N_9538,N_2679,N_694);
nand U9539 (N_9539,N_4806,N_1543);
and U9540 (N_9540,N_1214,N_1081);
xor U9541 (N_9541,N_1957,N_4546);
and U9542 (N_9542,N_1630,N_2647);
nand U9543 (N_9543,N_1323,N_3859);
nor U9544 (N_9544,N_3846,N_4120);
or U9545 (N_9545,N_3148,N_1036);
or U9546 (N_9546,N_1531,N_545);
and U9547 (N_9547,N_421,N_1589);
or U9548 (N_9548,N_4946,N_1406);
nor U9549 (N_9549,N_2821,N_3836);
and U9550 (N_9550,N_698,N_4211);
and U9551 (N_9551,N_2887,N_1700);
nor U9552 (N_9552,N_4678,N_1529);
and U9553 (N_9553,N_1427,N_949);
nor U9554 (N_9554,N_3741,N_1820);
nor U9555 (N_9555,N_3258,N_3013);
nand U9556 (N_9556,N_2981,N_2432);
and U9557 (N_9557,N_2351,N_3422);
or U9558 (N_9558,N_157,N_4474);
nor U9559 (N_9559,N_2823,N_4516);
nand U9560 (N_9560,N_552,N_2182);
nand U9561 (N_9561,N_3233,N_4463);
nand U9562 (N_9562,N_3882,N_1250);
nor U9563 (N_9563,N_430,N_2502);
or U9564 (N_9564,N_2373,N_1926);
nor U9565 (N_9565,N_2126,N_227);
nor U9566 (N_9566,N_2271,N_1481);
nor U9567 (N_9567,N_249,N_2634);
or U9568 (N_9568,N_4397,N_4784);
and U9569 (N_9569,N_4154,N_3811);
nor U9570 (N_9570,N_104,N_2717);
nor U9571 (N_9571,N_2965,N_2382);
or U9572 (N_9572,N_1017,N_2891);
nand U9573 (N_9573,N_2835,N_3427);
nor U9574 (N_9574,N_911,N_992);
and U9575 (N_9575,N_2050,N_4295);
and U9576 (N_9576,N_2999,N_1996);
or U9577 (N_9577,N_4115,N_4661);
and U9578 (N_9578,N_311,N_2461);
and U9579 (N_9579,N_1497,N_190);
and U9580 (N_9580,N_2457,N_4678);
and U9581 (N_9581,N_2754,N_2568);
nand U9582 (N_9582,N_1337,N_1975);
nand U9583 (N_9583,N_2482,N_415);
xor U9584 (N_9584,N_1017,N_2059);
or U9585 (N_9585,N_1564,N_2751);
nand U9586 (N_9586,N_2132,N_4715);
or U9587 (N_9587,N_3140,N_4191);
or U9588 (N_9588,N_1096,N_2785);
and U9589 (N_9589,N_4610,N_1511);
nor U9590 (N_9590,N_581,N_2332);
xor U9591 (N_9591,N_1526,N_3347);
nor U9592 (N_9592,N_4824,N_586);
or U9593 (N_9593,N_813,N_2289);
xor U9594 (N_9594,N_1137,N_2141);
or U9595 (N_9595,N_404,N_4025);
and U9596 (N_9596,N_4542,N_3711);
nor U9597 (N_9597,N_1061,N_519);
or U9598 (N_9598,N_3319,N_32);
nor U9599 (N_9599,N_4629,N_4907);
nor U9600 (N_9600,N_1006,N_2590);
nand U9601 (N_9601,N_3340,N_1001);
or U9602 (N_9602,N_1118,N_1583);
or U9603 (N_9603,N_916,N_205);
or U9604 (N_9604,N_835,N_4253);
nand U9605 (N_9605,N_2339,N_934);
or U9606 (N_9606,N_3032,N_4930);
and U9607 (N_9607,N_4719,N_4120);
or U9608 (N_9608,N_2839,N_3323);
and U9609 (N_9609,N_2414,N_4650);
and U9610 (N_9610,N_3037,N_3629);
nand U9611 (N_9611,N_1851,N_3926);
nand U9612 (N_9612,N_4877,N_313);
nor U9613 (N_9613,N_1809,N_1659);
nand U9614 (N_9614,N_3423,N_3728);
and U9615 (N_9615,N_4392,N_2012);
or U9616 (N_9616,N_4327,N_950);
nor U9617 (N_9617,N_4914,N_2382);
and U9618 (N_9618,N_3409,N_160);
or U9619 (N_9619,N_3063,N_4232);
and U9620 (N_9620,N_3703,N_2148);
and U9621 (N_9621,N_2980,N_3147);
nor U9622 (N_9622,N_2001,N_3382);
nor U9623 (N_9623,N_2117,N_4823);
and U9624 (N_9624,N_49,N_1725);
and U9625 (N_9625,N_2420,N_986);
nor U9626 (N_9626,N_4978,N_701);
nor U9627 (N_9627,N_2150,N_3385);
nand U9628 (N_9628,N_2157,N_2741);
nor U9629 (N_9629,N_1898,N_301);
and U9630 (N_9630,N_4265,N_3278);
nand U9631 (N_9631,N_2440,N_331);
and U9632 (N_9632,N_1031,N_4396);
nand U9633 (N_9633,N_3234,N_722);
xor U9634 (N_9634,N_1957,N_4645);
or U9635 (N_9635,N_1470,N_3498);
and U9636 (N_9636,N_3992,N_3680);
xnor U9637 (N_9637,N_3721,N_2480);
nor U9638 (N_9638,N_2215,N_224);
nand U9639 (N_9639,N_2421,N_2970);
or U9640 (N_9640,N_2485,N_2938);
nand U9641 (N_9641,N_4367,N_4491);
nor U9642 (N_9642,N_148,N_4398);
nor U9643 (N_9643,N_724,N_3214);
nand U9644 (N_9644,N_4393,N_4056);
or U9645 (N_9645,N_156,N_3583);
and U9646 (N_9646,N_1258,N_1526);
and U9647 (N_9647,N_270,N_3195);
or U9648 (N_9648,N_1798,N_64);
nor U9649 (N_9649,N_4146,N_1607);
nand U9650 (N_9650,N_1323,N_2558);
or U9651 (N_9651,N_2503,N_1180);
nor U9652 (N_9652,N_2367,N_3752);
nor U9653 (N_9653,N_4060,N_2817);
nor U9654 (N_9654,N_3601,N_682);
or U9655 (N_9655,N_2174,N_3026);
and U9656 (N_9656,N_2204,N_647);
nand U9657 (N_9657,N_4980,N_3710);
or U9658 (N_9658,N_1247,N_1827);
nor U9659 (N_9659,N_2254,N_3894);
nor U9660 (N_9660,N_2074,N_1054);
or U9661 (N_9661,N_2882,N_4572);
and U9662 (N_9662,N_2820,N_2333);
nor U9663 (N_9663,N_1528,N_4534);
or U9664 (N_9664,N_4173,N_4436);
and U9665 (N_9665,N_1968,N_4664);
nor U9666 (N_9666,N_3035,N_4611);
nand U9667 (N_9667,N_4800,N_20);
and U9668 (N_9668,N_2156,N_3569);
nand U9669 (N_9669,N_2195,N_4685);
or U9670 (N_9670,N_4306,N_1913);
xnor U9671 (N_9671,N_518,N_3596);
and U9672 (N_9672,N_792,N_2207);
nand U9673 (N_9673,N_2954,N_2755);
nor U9674 (N_9674,N_3572,N_2668);
nand U9675 (N_9675,N_4873,N_625);
or U9676 (N_9676,N_3716,N_11);
nand U9677 (N_9677,N_389,N_2731);
nand U9678 (N_9678,N_4410,N_2210);
nor U9679 (N_9679,N_3758,N_484);
and U9680 (N_9680,N_4952,N_1880);
or U9681 (N_9681,N_4267,N_2882);
and U9682 (N_9682,N_2876,N_2454);
or U9683 (N_9683,N_2491,N_3548);
and U9684 (N_9684,N_2042,N_2107);
or U9685 (N_9685,N_2389,N_4084);
nand U9686 (N_9686,N_4322,N_4942);
nand U9687 (N_9687,N_2883,N_2579);
nor U9688 (N_9688,N_3718,N_4234);
nor U9689 (N_9689,N_2838,N_3116);
or U9690 (N_9690,N_3925,N_2102);
nand U9691 (N_9691,N_3874,N_4110);
nor U9692 (N_9692,N_4107,N_790);
nor U9693 (N_9693,N_4798,N_3390);
nor U9694 (N_9694,N_1624,N_1224);
and U9695 (N_9695,N_1055,N_839);
nand U9696 (N_9696,N_1363,N_1581);
nor U9697 (N_9697,N_1724,N_4511);
and U9698 (N_9698,N_1073,N_1169);
nand U9699 (N_9699,N_2775,N_4892);
or U9700 (N_9700,N_158,N_3059);
or U9701 (N_9701,N_2861,N_4483);
nor U9702 (N_9702,N_868,N_2177);
and U9703 (N_9703,N_1511,N_4214);
or U9704 (N_9704,N_4410,N_4264);
xnor U9705 (N_9705,N_3961,N_3527);
or U9706 (N_9706,N_394,N_2261);
nor U9707 (N_9707,N_3350,N_2554);
nor U9708 (N_9708,N_785,N_2070);
nor U9709 (N_9709,N_3499,N_2151);
or U9710 (N_9710,N_2969,N_4320);
nand U9711 (N_9711,N_2658,N_829);
nor U9712 (N_9712,N_765,N_23);
nor U9713 (N_9713,N_980,N_4671);
nand U9714 (N_9714,N_2954,N_3324);
or U9715 (N_9715,N_2103,N_1020);
nor U9716 (N_9716,N_3471,N_4896);
and U9717 (N_9717,N_3382,N_1197);
nor U9718 (N_9718,N_3822,N_4621);
nand U9719 (N_9719,N_1012,N_80);
nand U9720 (N_9720,N_495,N_3803);
and U9721 (N_9721,N_237,N_3129);
nor U9722 (N_9722,N_2640,N_2159);
nand U9723 (N_9723,N_2365,N_2032);
and U9724 (N_9724,N_3821,N_3365);
or U9725 (N_9725,N_4074,N_3476);
nand U9726 (N_9726,N_4802,N_4156);
nor U9727 (N_9727,N_4219,N_2006);
or U9728 (N_9728,N_4891,N_261);
or U9729 (N_9729,N_1944,N_2949);
or U9730 (N_9730,N_3164,N_4371);
nand U9731 (N_9731,N_1673,N_1367);
nand U9732 (N_9732,N_2662,N_2485);
nand U9733 (N_9733,N_3741,N_1305);
xor U9734 (N_9734,N_1137,N_3211);
nand U9735 (N_9735,N_4895,N_1367);
or U9736 (N_9736,N_4014,N_3918);
nor U9737 (N_9737,N_3457,N_729);
nor U9738 (N_9738,N_2338,N_2758);
nand U9739 (N_9739,N_3348,N_381);
or U9740 (N_9740,N_3830,N_4965);
or U9741 (N_9741,N_3821,N_2349);
nand U9742 (N_9742,N_822,N_1110);
nor U9743 (N_9743,N_3610,N_978);
and U9744 (N_9744,N_725,N_4155);
or U9745 (N_9745,N_1227,N_4965);
nor U9746 (N_9746,N_3603,N_4918);
nand U9747 (N_9747,N_3123,N_2853);
nand U9748 (N_9748,N_1284,N_1941);
nor U9749 (N_9749,N_2976,N_2324);
or U9750 (N_9750,N_3771,N_1211);
or U9751 (N_9751,N_4036,N_1409);
nor U9752 (N_9752,N_2723,N_383);
and U9753 (N_9753,N_4188,N_3685);
and U9754 (N_9754,N_3121,N_2893);
and U9755 (N_9755,N_2324,N_4663);
and U9756 (N_9756,N_1717,N_2326);
nand U9757 (N_9757,N_221,N_819);
or U9758 (N_9758,N_2161,N_3216);
nand U9759 (N_9759,N_1339,N_3757);
or U9760 (N_9760,N_2281,N_817);
xor U9761 (N_9761,N_1950,N_3821);
nor U9762 (N_9762,N_786,N_2191);
nand U9763 (N_9763,N_2920,N_1615);
or U9764 (N_9764,N_3378,N_102);
nor U9765 (N_9765,N_4780,N_1335);
nand U9766 (N_9766,N_999,N_377);
and U9767 (N_9767,N_3518,N_2749);
and U9768 (N_9768,N_1944,N_2480);
nor U9769 (N_9769,N_1389,N_516);
and U9770 (N_9770,N_2602,N_3494);
nor U9771 (N_9771,N_111,N_1156);
nand U9772 (N_9772,N_3315,N_4173);
nor U9773 (N_9773,N_3375,N_4054);
or U9774 (N_9774,N_929,N_3635);
xor U9775 (N_9775,N_2340,N_3099);
nand U9776 (N_9776,N_2455,N_3130);
nand U9777 (N_9777,N_1784,N_4672);
xnor U9778 (N_9778,N_4558,N_1544);
or U9779 (N_9779,N_1361,N_4283);
nor U9780 (N_9780,N_2737,N_4523);
nor U9781 (N_9781,N_3475,N_2974);
xnor U9782 (N_9782,N_1131,N_3905);
nor U9783 (N_9783,N_960,N_4950);
nand U9784 (N_9784,N_2151,N_4227);
and U9785 (N_9785,N_1642,N_647);
nand U9786 (N_9786,N_3098,N_2121);
nand U9787 (N_9787,N_4949,N_2005);
nand U9788 (N_9788,N_605,N_956);
and U9789 (N_9789,N_2958,N_565);
or U9790 (N_9790,N_3091,N_715);
nor U9791 (N_9791,N_3181,N_1854);
and U9792 (N_9792,N_2788,N_4312);
nor U9793 (N_9793,N_3900,N_3805);
or U9794 (N_9794,N_200,N_2174);
nand U9795 (N_9795,N_4777,N_2797);
nor U9796 (N_9796,N_954,N_1518);
and U9797 (N_9797,N_1113,N_1200);
and U9798 (N_9798,N_1279,N_3270);
or U9799 (N_9799,N_1170,N_1739);
nor U9800 (N_9800,N_2638,N_1157);
nor U9801 (N_9801,N_1540,N_4107);
or U9802 (N_9802,N_2370,N_2143);
nor U9803 (N_9803,N_4447,N_1304);
nand U9804 (N_9804,N_1248,N_505);
nand U9805 (N_9805,N_2309,N_4774);
nor U9806 (N_9806,N_698,N_3536);
and U9807 (N_9807,N_3378,N_1378);
and U9808 (N_9808,N_2045,N_3282);
or U9809 (N_9809,N_2610,N_831);
and U9810 (N_9810,N_294,N_2746);
nor U9811 (N_9811,N_563,N_4364);
nand U9812 (N_9812,N_2647,N_2056);
and U9813 (N_9813,N_1453,N_4416);
nor U9814 (N_9814,N_178,N_3238);
or U9815 (N_9815,N_2733,N_1645);
nand U9816 (N_9816,N_1658,N_678);
nor U9817 (N_9817,N_83,N_145);
or U9818 (N_9818,N_2043,N_4548);
and U9819 (N_9819,N_1953,N_998);
nor U9820 (N_9820,N_924,N_2716);
xor U9821 (N_9821,N_486,N_1095);
and U9822 (N_9822,N_1549,N_4188);
and U9823 (N_9823,N_772,N_2587);
and U9824 (N_9824,N_2089,N_3472);
nand U9825 (N_9825,N_3492,N_4062);
nor U9826 (N_9826,N_3117,N_4204);
nor U9827 (N_9827,N_4921,N_4574);
or U9828 (N_9828,N_1426,N_1502);
or U9829 (N_9829,N_2336,N_1437);
and U9830 (N_9830,N_3263,N_3159);
or U9831 (N_9831,N_2207,N_3702);
or U9832 (N_9832,N_819,N_2509);
nor U9833 (N_9833,N_1306,N_1844);
nor U9834 (N_9834,N_4064,N_3699);
nand U9835 (N_9835,N_2855,N_3963);
nor U9836 (N_9836,N_2952,N_1148);
nand U9837 (N_9837,N_1383,N_4658);
and U9838 (N_9838,N_2826,N_4994);
nand U9839 (N_9839,N_2865,N_1159);
and U9840 (N_9840,N_1473,N_3535);
nor U9841 (N_9841,N_505,N_2475);
nand U9842 (N_9842,N_2513,N_1104);
or U9843 (N_9843,N_2442,N_2899);
or U9844 (N_9844,N_1026,N_1705);
and U9845 (N_9845,N_2692,N_824);
nand U9846 (N_9846,N_4839,N_2459);
and U9847 (N_9847,N_2438,N_3742);
and U9848 (N_9848,N_2710,N_4422);
nor U9849 (N_9849,N_1731,N_820);
nand U9850 (N_9850,N_1089,N_176);
and U9851 (N_9851,N_4581,N_115);
nor U9852 (N_9852,N_967,N_1015);
or U9853 (N_9853,N_1652,N_1653);
nor U9854 (N_9854,N_2774,N_14);
and U9855 (N_9855,N_2032,N_2406);
nor U9856 (N_9856,N_537,N_893);
nand U9857 (N_9857,N_3804,N_3808);
and U9858 (N_9858,N_56,N_1899);
or U9859 (N_9859,N_574,N_2644);
nor U9860 (N_9860,N_4105,N_4914);
nor U9861 (N_9861,N_1439,N_258);
or U9862 (N_9862,N_917,N_2559);
and U9863 (N_9863,N_3097,N_3276);
and U9864 (N_9864,N_4290,N_1901);
or U9865 (N_9865,N_4702,N_4644);
and U9866 (N_9866,N_1412,N_992);
and U9867 (N_9867,N_4226,N_1253);
nand U9868 (N_9868,N_255,N_242);
or U9869 (N_9869,N_3467,N_4283);
and U9870 (N_9870,N_2533,N_4345);
nand U9871 (N_9871,N_2685,N_4784);
or U9872 (N_9872,N_3528,N_4958);
nor U9873 (N_9873,N_2029,N_4129);
nand U9874 (N_9874,N_3350,N_191);
nor U9875 (N_9875,N_2243,N_2618);
nor U9876 (N_9876,N_2599,N_4219);
and U9877 (N_9877,N_4555,N_2102);
nand U9878 (N_9878,N_3890,N_3231);
nor U9879 (N_9879,N_3037,N_4920);
nor U9880 (N_9880,N_554,N_4522);
and U9881 (N_9881,N_1102,N_3333);
xnor U9882 (N_9882,N_993,N_369);
nand U9883 (N_9883,N_4711,N_29);
xnor U9884 (N_9884,N_254,N_4700);
and U9885 (N_9885,N_1439,N_696);
nand U9886 (N_9886,N_4181,N_3722);
nand U9887 (N_9887,N_4497,N_1830);
nor U9888 (N_9888,N_2602,N_2692);
or U9889 (N_9889,N_2300,N_30);
or U9890 (N_9890,N_2829,N_268);
nand U9891 (N_9891,N_1923,N_1099);
nand U9892 (N_9892,N_637,N_4170);
nand U9893 (N_9893,N_755,N_1208);
or U9894 (N_9894,N_4674,N_2847);
and U9895 (N_9895,N_1539,N_4684);
nand U9896 (N_9896,N_4213,N_2588);
and U9897 (N_9897,N_339,N_2820);
and U9898 (N_9898,N_3494,N_413);
or U9899 (N_9899,N_3700,N_1208);
nand U9900 (N_9900,N_746,N_4958);
nand U9901 (N_9901,N_1754,N_3971);
nand U9902 (N_9902,N_4821,N_2500);
and U9903 (N_9903,N_1660,N_2071);
or U9904 (N_9904,N_15,N_1316);
or U9905 (N_9905,N_1658,N_4472);
and U9906 (N_9906,N_1060,N_1666);
nor U9907 (N_9907,N_429,N_3426);
nor U9908 (N_9908,N_90,N_4613);
nand U9909 (N_9909,N_1477,N_2799);
nor U9910 (N_9910,N_1563,N_1814);
nand U9911 (N_9911,N_3636,N_2382);
or U9912 (N_9912,N_3649,N_887);
and U9913 (N_9913,N_2340,N_2871);
nand U9914 (N_9914,N_4378,N_4803);
nor U9915 (N_9915,N_126,N_4012);
or U9916 (N_9916,N_4639,N_3345);
or U9917 (N_9917,N_2440,N_371);
nand U9918 (N_9918,N_468,N_2584);
xor U9919 (N_9919,N_3597,N_2808);
and U9920 (N_9920,N_2785,N_2864);
and U9921 (N_9921,N_1134,N_486);
nor U9922 (N_9922,N_267,N_957);
or U9923 (N_9923,N_2670,N_3952);
nor U9924 (N_9924,N_3546,N_2808);
or U9925 (N_9925,N_1930,N_2925);
nor U9926 (N_9926,N_2426,N_2009);
nor U9927 (N_9927,N_4600,N_1692);
nor U9928 (N_9928,N_911,N_1188);
xor U9929 (N_9929,N_2843,N_4871);
nand U9930 (N_9930,N_823,N_1967);
and U9931 (N_9931,N_195,N_2243);
nand U9932 (N_9932,N_4326,N_1799);
nor U9933 (N_9933,N_669,N_984);
and U9934 (N_9934,N_3036,N_17);
xor U9935 (N_9935,N_2868,N_2321);
nand U9936 (N_9936,N_1494,N_1634);
and U9937 (N_9937,N_425,N_65);
nand U9938 (N_9938,N_1225,N_4078);
nor U9939 (N_9939,N_4409,N_3320);
nor U9940 (N_9940,N_4573,N_2592);
or U9941 (N_9941,N_3964,N_4972);
nand U9942 (N_9942,N_4475,N_2786);
nand U9943 (N_9943,N_3866,N_1784);
nand U9944 (N_9944,N_698,N_3690);
or U9945 (N_9945,N_4706,N_4225);
and U9946 (N_9946,N_2092,N_4086);
nand U9947 (N_9947,N_3354,N_3031);
nand U9948 (N_9948,N_4680,N_2702);
or U9949 (N_9949,N_2257,N_3802);
and U9950 (N_9950,N_4801,N_246);
or U9951 (N_9951,N_964,N_1713);
nor U9952 (N_9952,N_4758,N_4347);
or U9953 (N_9953,N_1696,N_2006);
xnor U9954 (N_9954,N_1382,N_3084);
and U9955 (N_9955,N_4588,N_497);
nand U9956 (N_9956,N_4393,N_4398);
and U9957 (N_9957,N_4453,N_4972);
and U9958 (N_9958,N_4461,N_1500);
nand U9959 (N_9959,N_2842,N_1943);
nor U9960 (N_9960,N_4606,N_1079);
nor U9961 (N_9961,N_4405,N_46);
and U9962 (N_9962,N_3339,N_1419);
or U9963 (N_9963,N_1307,N_139);
nand U9964 (N_9964,N_2962,N_1381);
and U9965 (N_9965,N_4842,N_3357);
or U9966 (N_9966,N_3645,N_1241);
or U9967 (N_9967,N_3953,N_349);
nor U9968 (N_9968,N_1174,N_4143);
and U9969 (N_9969,N_2606,N_4357);
or U9970 (N_9970,N_2658,N_4332);
and U9971 (N_9971,N_2334,N_4047);
nor U9972 (N_9972,N_3576,N_4733);
and U9973 (N_9973,N_1264,N_2828);
and U9974 (N_9974,N_462,N_4969);
nand U9975 (N_9975,N_608,N_1847);
nor U9976 (N_9976,N_3574,N_3647);
nor U9977 (N_9977,N_2775,N_3077);
or U9978 (N_9978,N_4361,N_705);
or U9979 (N_9979,N_2174,N_1183);
nand U9980 (N_9980,N_726,N_3173);
nor U9981 (N_9981,N_3138,N_1379);
and U9982 (N_9982,N_4160,N_4013);
and U9983 (N_9983,N_3467,N_1958);
nand U9984 (N_9984,N_3842,N_2110);
nand U9985 (N_9985,N_1127,N_3837);
and U9986 (N_9986,N_4820,N_2004);
nor U9987 (N_9987,N_637,N_3078);
nor U9988 (N_9988,N_426,N_1272);
nand U9989 (N_9989,N_4216,N_1673);
or U9990 (N_9990,N_4969,N_665);
nor U9991 (N_9991,N_508,N_1784);
nor U9992 (N_9992,N_2979,N_413);
xor U9993 (N_9993,N_1503,N_1036);
or U9994 (N_9994,N_4892,N_2650);
xor U9995 (N_9995,N_3107,N_546);
and U9996 (N_9996,N_3740,N_3989);
or U9997 (N_9997,N_4386,N_3694);
nor U9998 (N_9998,N_4077,N_2647);
or U9999 (N_9999,N_3309,N_4631);
nand UO_0 (O_0,N_6203,N_5288);
or UO_1 (O_1,N_5781,N_9322);
or UO_2 (O_2,N_8217,N_5909);
nor UO_3 (O_3,N_7646,N_8683);
and UO_4 (O_4,N_8888,N_7767);
nand UO_5 (O_5,N_5403,N_9145);
nor UO_6 (O_6,N_6170,N_8639);
or UO_7 (O_7,N_5450,N_7281);
and UO_8 (O_8,N_8400,N_7955);
and UO_9 (O_9,N_6162,N_9408);
and UO_10 (O_10,N_8689,N_8160);
and UO_11 (O_11,N_9730,N_7042);
or UO_12 (O_12,N_6655,N_5993);
nand UO_13 (O_13,N_7600,N_6732);
or UO_14 (O_14,N_9900,N_8473);
or UO_15 (O_15,N_8070,N_8514);
nand UO_16 (O_16,N_7043,N_8945);
nand UO_17 (O_17,N_9460,N_7209);
or UO_18 (O_18,N_5320,N_8375);
nor UO_19 (O_19,N_6641,N_8944);
and UO_20 (O_20,N_6236,N_6485);
nand UO_21 (O_21,N_6527,N_5911);
and UO_22 (O_22,N_6388,N_9686);
and UO_23 (O_23,N_8486,N_6231);
nand UO_24 (O_24,N_7436,N_6816);
or UO_25 (O_25,N_9877,N_9869);
and UO_26 (O_26,N_6623,N_5373);
nand UO_27 (O_27,N_7664,N_7055);
or UO_28 (O_28,N_8450,N_9649);
and UO_29 (O_29,N_6884,N_9246);
and UO_30 (O_30,N_6668,N_9057);
or UO_31 (O_31,N_5446,N_6241);
nor UO_32 (O_32,N_9290,N_6034);
nand UO_33 (O_33,N_6577,N_8489);
and UO_34 (O_34,N_7838,N_7178);
nand UO_35 (O_35,N_8541,N_8590);
or UO_36 (O_36,N_7880,N_5766);
nand UO_37 (O_37,N_5897,N_6556);
nand UO_38 (O_38,N_7250,N_9051);
or UO_39 (O_39,N_7951,N_5437);
nor UO_40 (O_40,N_6061,N_5945);
nor UO_41 (O_41,N_7064,N_6591);
nor UO_42 (O_42,N_9979,N_5064);
or UO_43 (O_43,N_8250,N_9608);
nor UO_44 (O_44,N_8445,N_8105);
or UO_45 (O_45,N_7180,N_9415);
or UO_46 (O_46,N_5289,N_9710);
or UO_47 (O_47,N_7310,N_7947);
and UO_48 (O_48,N_8209,N_8826);
or UO_49 (O_49,N_8335,N_7817);
nand UO_50 (O_50,N_9647,N_5455);
nor UO_51 (O_51,N_5096,N_7982);
nor UO_52 (O_52,N_8617,N_5746);
nand UO_53 (O_53,N_5310,N_6195);
nand UO_54 (O_54,N_8745,N_7854);
nor UO_55 (O_55,N_5379,N_9928);
nand UO_56 (O_56,N_8896,N_5974);
nor UO_57 (O_57,N_7607,N_6228);
nor UO_58 (O_58,N_7416,N_8420);
nand UO_59 (O_59,N_7348,N_6482);
xor UO_60 (O_60,N_6330,N_7273);
nor UO_61 (O_61,N_7901,N_7068);
or UO_62 (O_62,N_6188,N_5734);
and UO_63 (O_63,N_7459,N_5458);
xor UO_64 (O_64,N_5034,N_6376);
xnor UO_65 (O_65,N_8410,N_8679);
nand UO_66 (O_66,N_8027,N_6108);
nand UO_67 (O_67,N_8857,N_9855);
and UO_68 (O_68,N_6303,N_8607);
and UO_69 (O_69,N_9708,N_9175);
nor UO_70 (O_70,N_6797,N_9889);
nand UO_71 (O_71,N_8128,N_9072);
and UO_72 (O_72,N_8759,N_5869);
or UO_73 (O_73,N_7551,N_5996);
or UO_74 (O_74,N_8164,N_8819);
nand UO_75 (O_75,N_9225,N_5214);
or UO_76 (O_76,N_7711,N_6347);
and UO_77 (O_77,N_7338,N_9455);
nand UO_78 (O_78,N_9032,N_8207);
and UO_79 (O_79,N_5792,N_5668);
nor UO_80 (O_80,N_7127,N_7748);
xor UO_81 (O_81,N_7566,N_8659);
nor UO_82 (O_82,N_8176,N_8146);
or UO_83 (O_83,N_5097,N_5386);
and UO_84 (O_84,N_6194,N_7833);
and UO_85 (O_85,N_8744,N_7602);
or UO_86 (O_86,N_7017,N_6397);
or UO_87 (O_87,N_6851,N_5979);
or UO_88 (O_88,N_9784,N_8701);
or UO_89 (O_89,N_5518,N_5009);
or UO_90 (O_90,N_5307,N_8982);
nand UO_91 (O_91,N_7543,N_5239);
nor UO_92 (O_92,N_5418,N_6944);
nand UO_93 (O_93,N_5402,N_5902);
and UO_94 (O_94,N_5126,N_9538);
nor UO_95 (O_95,N_7078,N_7830);
or UO_96 (O_96,N_5975,N_5068);
and UO_97 (O_97,N_7812,N_8838);
nand UO_98 (O_98,N_8974,N_6364);
and UO_99 (O_99,N_8116,N_7331);
nand UO_100 (O_100,N_8769,N_6608);
or UO_101 (O_101,N_8787,N_8980);
and UO_102 (O_102,N_5567,N_5719);
nand UO_103 (O_103,N_5253,N_5414);
or UO_104 (O_104,N_5390,N_6494);
and UO_105 (O_105,N_5584,N_7016);
nand UO_106 (O_106,N_5234,N_8515);
nand UO_107 (O_107,N_6825,N_8600);
nor UO_108 (O_108,N_9048,N_9157);
nor UO_109 (O_109,N_7930,N_9717);
and UO_110 (O_110,N_7141,N_8568);
nand UO_111 (O_111,N_5116,N_5790);
nand UO_112 (O_112,N_6841,N_5577);
and UO_113 (O_113,N_6717,N_6921);
or UO_114 (O_114,N_9926,N_7666);
and UO_115 (O_115,N_6726,N_7974);
xor UO_116 (O_116,N_8379,N_6656);
and UO_117 (O_117,N_8343,N_9908);
nand UO_118 (O_118,N_5449,N_6399);
nor UO_119 (O_119,N_7261,N_6786);
or UO_120 (O_120,N_8082,N_9777);
and UO_121 (O_121,N_9948,N_6950);
nand UO_122 (O_122,N_8198,N_9026);
and UO_123 (O_123,N_9227,N_6073);
xnor UO_124 (O_124,N_6242,N_7576);
nor UO_125 (O_125,N_8772,N_6526);
nand UO_126 (O_126,N_9761,N_8923);
or UO_127 (O_127,N_9907,N_7347);
or UO_128 (O_128,N_7557,N_6269);
and UO_129 (O_129,N_5687,N_5195);
nor UO_130 (O_130,N_6349,N_6327);
and UO_131 (O_131,N_7352,N_6848);
and UO_132 (O_132,N_8699,N_9007);
nor UO_133 (O_133,N_9836,N_9350);
and UO_134 (O_134,N_7906,N_9807);
nor UO_135 (O_135,N_6290,N_7033);
nor UO_136 (O_136,N_6071,N_9078);
and UO_137 (O_137,N_9917,N_7218);
nor UO_138 (O_138,N_9108,N_6757);
nand UO_139 (O_139,N_9395,N_5335);
nor UO_140 (O_140,N_7045,N_6479);
and UO_141 (O_141,N_5342,N_9399);
nor UO_142 (O_142,N_5500,N_6172);
and UO_143 (O_143,N_5968,N_9512);
or UO_144 (O_144,N_7909,N_7279);
nand UO_145 (O_145,N_6723,N_9791);
nand UO_146 (O_146,N_9077,N_5000);
or UO_147 (O_147,N_7921,N_5616);
nand UO_148 (O_148,N_5571,N_8064);
or UO_149 (O_149,N_8144,N_9678);
nor UO_150 (O_150,N_6956,N_5081);
nand UO_151 (O_151,N_8504,N_7554);
nor UO_152 (O_152,N_7675,N_9128);
nor UO_153 (O_153,N_9558,N_5121);
or UO_154 (O_154,N_9581,N_5609);
and UO_155 (O_155,N_7692,N_9853);
nor UO_156 (O_156,N_5704,N_7380);
or UO_157 (O_157,N_8038,N_5711);
nand UO_158 (O_158,N_6049,N_8002);
nor UO_159 (O_159,N_8993,N_6139);
and UO_160 (O_160,N_5212,N_6986);
nand UO_161 (O_161,N_9946,N_7632);
and UO_162 (O_162,N_9284,N_5557);
or UO_163 (O_163,N_6100,N_9531);
and UO_164 (O_164,N_9789,N_8480);
or UO_165 (O_165,N_9337,N_5194);
nor UO_166 (O_166,N_7189,N_9704);
or UO_167 (O_167,N_8275,N_7842);
and UO_168 (O_168,N_7004,N_9420);
and UO_169 (O_169,N_5163,N_6524);
nor UO_170 (O_170,N_6968,N_5898);
or UO_171 (O_171,N_8163,N_9648);
nand UO_172 (O_172,N_7420,N_9438);
nor UO_173 (O_173,N_9905,N_9863);
nand UO_174 (O_174,N_7469,N_9472);
nor UO_175 (O_175,N_7239,N_9003);
or UO_176 (O_176,N_6215,N_8681);
nor UO_177 (O_177,N_7193,N_8692);
nor UO_178 (O_178,N_7356,N_7034);
nor UO_179 (O_179,N_5858,N_5261);
nand UO_180 (O_180,N_7482,N_5337);
and UO_181 (O_181,N_9440,N_9443);
or UO_182 (O_182,N_6324,N_5836);
nand UO_183 (O_183,N_7563,N_6690);
nor UO_184 (O_184,N_6083,N_7673);
or UO_185 (O_185,N_9457,N_8523);
or UO_186 (O_186,N_7210,N_5456);
nor UO_187 (O_187,N_6141,N_6999);
or UO_188 (O_188,N_7136,N_5039);
or UO_189 (O_189,N_7027,N_9870);
or UO_190 (O_190,N_6400,N_9474);
nor UO_191 (O_191,N_9463,N_9788);
nor UO_192 (O_192,N_6159,N_7399);
and UO_193 (O_193,N_5521,N_5680);
nor UO_194 (O_194,N_8167,N_6138);
nor UO_195 (O_195,N_9864,N_7358);
nor UO_196 (O_196,N_6193,N_5689);
nor UO_197 (O_197,N_6911,N_7256);
nand UO_198 (O_198,N_6261,N_6371);
or UO_199 (O_199,N_9112,N_9379);
nor UO_200 (O_200,N_7095,N_8093);
nor UO_201 (O_201,N_6965,N_8933);
or UO_202 (O_202,N_5193,N_8970);
or UO_203 (O_203,N_9485,N_6198);
or UO_204 (O_204,N_7548,N_8632);
or UO_205 (O_205,N_6199,N_8562);
nor UO_206 (O_206,N_9582,N_7792);
and UO_207 (O_207,N_5368,N_7944);
or UO_208 (O_208,N_7533,N_7571);
or UO_209 (O_209,N_8610,N_7162);
nor UO_210 (O_210,N_6209,N_5108);
and UO_211 (O_211,N_8653,N_6619);
nor UO_212 (O_212,N_7631,N_6461);
nor UO_213 (O_213,N_7391,N_8241);
nor UO_214 (O_214,N_8351,N_9879);
and UO_215 (O_215,N_9847,N_7173);
nand UO_216 (O_216,N_7492,N_7130);
nor UO_217 (O_217,N_5767,N_6845);
nand UO_218 (O_218,N_8867,N_7468);
nor UO_219 (O_219,N_8475,N_5093);
or UO_220 (O_220,N_9653,N_6940);
nor UO_221 (O_221,N_9957,N_7057);
and UO_222 (O_222,N_7528,N_9177);
nand UO_223 (O_223,N_6029,N_8413);
or UO_224 (O_224,N_5159,N_6562);
or UO_225 (O_225,N_5138,N_8517);
or UO_226 (O_226,N_6616,N_5472);
nor UO_227 (O_227,N_5002,N_9812);
nand UO_228 (O_228,N_6916,N_7378);
and UO_229 (O_229,N_6362,N_8537);
or UO_230 (O_230,N_8300,N_5545);
nor UO_231 (O_231,N_5873,N_7463);
nor UO_232 (O_232,N_8254,N_6091);
nor UO_233 (O_233,N_9272,N_6729);
or UO_234 (O_234,N_8870,N_7496);
nand UO_235 (O_235,N_5326,N_5572);
nor UO_236 (O_236,N_5808,N_7709);
nor UO_237 (O_237,N_5049,N_8208);
nor UO_238 (O_238,N_9303,N_7037);
and UO_239 (O_239,N_8066,N_5896);
or UO_240 (O_240,N_6705,N_7464);
and UO_241 (O_241,N_8899,N_6930);
nor UO_242 (O_242,N_9308,N_6266);
nor UO_243 (O_243,N_6926,N_7970);
xor UO_244 (O_244,N_7236,N_8553);
nand UO_245 (O_245,N_6165,N_6271);
nand UO_246 (O_246,N_9413,N_8832);
or UO_247 (O_247,N_6111,N_5479);
nor UO_248 (O_248,N_6742,N_7712);
or UO_249 (O_249,N_6948,N_7789);
or UO_250 (O_250,N_9375,N_9106);
and UO_251 (O_251,N_5916,N_8365);
or UO_252 (O_252,N_6394,N_9358);
nand UO_253 (O_253,N_7323,N_6633);
or UO_254 (O_254,N_8126,N_5627);
nor UO_255 (O_255,N_6815,N_6676);
or UO_256 (O_256,N_7957,N_7235);
xor UO_257 (O_257,N_5243,N_6217);
or UO_258 (O_258,N_5170,N_5197);
and UO_259 (O_259,N_5341,N_7036);
nor UO_260 (O_260,N_6929,N_6761);
and UO_261 (O_261,N_9451,N_7876);
or UO_262 (O_262,N_9274,N_9596);
nor UO_263 (O_263,N_6810,N_5165);
nand UO_264 (O_264,N_5556,N_7419);
and UO_265 (O_265,N_9300,N_8127);
xor UO_266 (O_266,N_5330,N_5976);
nor UO_267 (O_267,N_9071,N_9436);
or UO_268 (O_268,N_6128,N_6201);
xor UO_269 (O_269,N_8336,N_5722);
xor UO_270 (O_270,N_6772,N_8042);
nor UO_271 (O_271,N_5721,N_8513);
and UO_272 (O_272,N_5819,N_5526);
or UO_273 (O_273,N_9035,N_8078);
xor UO_274 (O_274,N_8465,N_5645);
or UO_275 (O_275,N_9533,N_7121);
nor UO_276 (O_276,N_5353,N_8799);
or UO_277 (O_277,N_6332,N_6160);
nor UO_278 (O_278,N_7025,N_7715);
or UO_279 (O_279,N_9130,N_5140);
nor UO_280 (O_280,N_9831,N_8573);
nand UO_281 (O_281,N_5800,N_5345);
nand UO_282 (O_282,N_7101,N_9080);
nor UO_283 (O_283,N_5533,N_5849);
nand UO_284 (O_284,N_5220,N_8056);
and UO_285 (O_285,N_7780,N_9196);
nor UO_286 (O_286,N_7474,N_9739);
nor UO_287 (O_287,N_9743,N_6245);
or UO_288 (O_288,N_8150,N_5016);
nor UO_289 (O_289,N_6080,N_7979);
nand UO_290 (O_290,N_8592,N_8873);
and UO_291 (O_291,N_7756,N_9329);
and UO_292 (O_292,N_7259,N_6420);
or UO_293 (O_293,N_9467,N_6272);
or UO_294 (O_294,N_5618,N_9240);
and UO_295 (O_295,N_7245,N_7920);
nand UO_296 (O_296,N_9846,N_5566);
or UO_297 (O_297,N_7514,N_6695);
or UO_298 (O_298,N_6918,N_7367);
and UO_299 (O_299,N_5133,N_7731);
nor UO_300 (O_300,N_6316,N_7917);
nand UO_301 (O_301,N_9091,N_9473);
nor UO_302 (O_302,N_7820,N_8652);
and UO_303 (O_303,N_9235,N_6666);
or UO_304 (O_304,N_6146,N_7144);
and UO_305 (O_305,N_6740,N_8147);
nand UO_306 (O_306,N_8720,N_5463);
and UO_307 (O_307,N_6246,N_5839);
nand UO_308 (O_308,N_5200,N_9553);
nor UO_309 (O_309,N_6919,N_6835);
nor UO_310 (O_310,N_6584,N_6805);
or UO_311 (O_311,N_9560,N_8060);
or UO_312 (O_312,N_8471,N_7351);
xnor UO_313 (O_313,N_7953,N_6727);
xnor UO_314 (O_314,N_6306,N_7595);
nand UO_315 (O_315,N_9471,N_5775);
nor UO_316 (O_316,N_5638,N_6973);
nand UO_317 (O_317,N_7440,N_6998);
nor UO_318 (O_318,N_9511,N_9214);
or UO_319 (O_319,N_9790,N_6097);
or UO_320 (O_320,N_5124,N_7502);
or UO_321 (O_321,N_8650,N_8015);
nand UO_322 (O_322,N_8782,N_6003);
or UO_323 (O_323,N_6774,N_7931);
and UO_324 (O_324,N_6229,N_9155);
nor UO_325 (O_325,N_7108,N_6429);
and UO_326 (O_326,N_7490,N_6876);
and UO_327 (O_327,N_8900,N_9816);
nor UO_328 (O_328,N_6744,N_6635);
and UO_329 (O_329,N_9386,N_5186);
and UO_330 (O_330,N_9731,N_7206);
nand UO_331 (O_331,N_8874,N_9990);
nand UO_332 (O_332,N_5529,N_8442);
and UO_333 (O_333,N_5678,N_8131);
nand UO_334 (O_334,N_9468,N_7730);
xnor UO_335 (O_335,N_6067,N_8468);
and UO_336 (O_336,N_7443,N_7132);
and UO_337 (O_337,N_9412,N_9779);
and UO_338 (O_338,N_7908,N_8753);
nand UO_339 (O_339,N_6997,N_7237);
and UO_340 (O_340,N_5465,N_8499);
nand UO_341 (O_341,N_8404,N_8114);
nor UO_342 (O_342,N_7183,N_9709);
nand UO_343 (O_343,N_6273,N_7978);
or UO_344 (O_344,N_8459,N_6563);
and UO_345 (O_345,N_8758,N_5946);
nand UO_346 (O_346,N_7522,N_7035);
or UO_347 (O_347,N_8662,N_9762);
nand UO_348 (O_348,N_7645,N_8429);
nor UO_349 (O_349,N_7003,N_7758);
or UO_350 (O_350,N_6730,N_7825);
and UO_351 (O_351,N_9897,N_6471);
nand UO_352 (O_352,N_9366,N_5853);
nor UO_353 (O_353,N_9400,N_5271);
nor UO_354 (O_354,N_8360,N_7403);
and UO_355 (O_355,N_7871,N_6678);
nand UO_356 (O_356,N_9492,N_6068);
or UO_357 (O_357,N_8438,N_7450);
and UO_358 (O_358,N_9969,N_9099);
nand UO_359 (O_359,N_6122,N_8273);
and UO_360 (O_360,N_6731,N_5783);
nor UO_361 (O_361,N_9824,N_5510);
and UO_362 (O_362,N_9691,N_7861);
or UO_363 (O_363,N_5073,N_5051);
nand UO_364 (O_364,N_6045,N_7983);
nor UO_365 (O_365,N_5664,N_8495);
nand UO_366 (O_366,N_9960,N_9442);
nor UO_367 (O_367,N_7312,N_6181);
and UO_368 (O_368,N_5021,N_7605);
nand UO_369 (O_369,N_9149,N_7125);
and UO_370 (O_370,N_7487,N_7676);
and UO_371 (O_371,N_5648,N_6788);
nand UO_372 (O_372,N_6499,N_6515);
and UO_373 (O_373,N_7845,N_7958);
or UO_374 (O_374,N_7989,N_9619);
nand UO_375 (O_375,N_7642,N_9482);
or UO_376 (O_376,N_7881,N_9297);
xnor UO_377 (O_377,N_6454,N_9189);
and UO_378 (O_378,N_8717,N_8387);
nand UO_379 (O_379,N_8016,N_9935);
nand UO_380 (O_380,N_5130,N_5570);
nor UO_381 (O_381,N_6208,N_5628);
nand UO_382 (O_382,N_9277,N_5520);
and UO_383 (O_383,N_5606,N_6348);
or UO_384 (O_384,N_7296,N_9475);
or UO_385 (O_385,N_6522,N_8149);
nor UO_386 (O_386,N_9574,N_5823);
nor UO_387 (O_387,N_6513,N_5983);
nor UO_388 (O_388,N_8816,N_9359);
or UO_389 (O_389,N_8373,N_6383);
nor UO_390 (O_390,N_7226,N_7702);
and UO_391 (O_391,N_8109,N_6590);
nand UO_392 (O_392,N_8141,N_7946);
nand UO_393 (O_393,N_8986,N_5615);
and UO_394 (O_394,N_6476,N_7021);
and UO_395 (O_395,N_9724,N_8466);
or UO_396 (O_396,N_5391,N_8436);
or UO_397 (O_397,N_8219,N_7574);
and UO_398 (O_398,N_5442,N_8997);
and UO_399 (O_399,N_8877,N_8107);
nand UO_400 (O_400,N_9076,N_9659);
or UO_401 (O_401,N_5183,N_9577);
nor UO_402 (O_402,N_9244,N_7063);
nor UO_403 (O_403,N_7369,N_5876);
and UO_404 (O_404,N_7685,N_5489);
or UO_405 (O_405,N_7105,N_5791);
or UO_406 (O_406,N_9997,N_5630);
nand UO_407 (O_407,N_6355,N_5364);
or UO_408 (O_408,N_5065,N_6496);
xnor UO_409 (O_409,N_6132,N_6636);
xor UO_410 (O_410,N_8330,N_6707);
and UO_411 (O_411,N_9923,N_9707);
or UO_412 (O_412,N_9949,N_7243);
nor UO_413 (O_413,N_8668,N_6975);
and UO_414 (O_414,N_8182,N_6148);
xor UO_415 (O_415,N_7379,N_9182);
or UO_416 (O_416,N_7560,N_8845);
nor UO_417 (O_417,N_9745,N_5705);
nand UO_418 (O_418,N_9414,N_7044);
nand UO_419 (O_419,N_5813,N_7579);
nand UO_420 (O_420,N_7328,N_6697);
nand UO_421 (O_421,N_9346,N_7846);
nor UO_422 (O_422,N_8189,N_8521);
nand UO_423 (O_423,N_9744,N_5552);
nor UO_424 (O_424,N_9749,N_6235);
nand UO_425 (O_425,N_5700,N_6820);
or UO_426 (O_426,N_6781,N_7733);
and UO_427 (O_427,N_5929,N_6747);
nor UO_428 (O_428,N_7678,N_8784);
nand UO_429 (O_429,N_8591,N_6501);
and UO_430 (O_430,N_9685,N_9858);
or UO_431 (O_431,N_9341,N_6418);
nand UO_432 (O_432,N_8801,N_7618);
or UO_433 (O_433,N_9845,N_6465);
nor UO_434 (O_434,N_5279,N_9740);
nand UO_435 (O_435,N_7747,N_9198);
and UO_436 (O_436,N_8034,N_5433);
nor UO_437 (O_437,N_8071,N_9248);
or UO_438 (O_438,N_9320,N_9103);
nor UO_439 (O_439,N_6120,N_6451);
nand UO_440 (O_440,N_6407,N_5480);
nand UO_441 (O_441,N_5597,N_7360);
or UO_442 (O_442,N_7550,N_8519);
nand UO_443 (O_443,N_7752,N_7945);
nor UO_444 (O_444,N_7168,N_8694);
nand UO_445 (O_445,N_5865,N_6180);
and UO_446 (O_446,N_7995,N_9302);
and UO_447 (O_447,N_6265,N_6745);
nor UO_448 (O_448,N_7956,N_7948);
nor UO_449 (O_449,N_9934,N_7085);
or UO_450 (O_450,N_6259,N_6028);
and UO_451 (O_451,N_5313,N_5099);
nand UO_452 (O_452,N_8138,N_8080);
and UO_453 (O_453,N_6904,N_9956);
and UO_454 (O_454,N_5206,N_9105);
nor UO_455 (O_455,N_8314,N_6769);
nor UO_456 (O_456,N_6571,N_9715);
or UO_457 (O_457,N_9669,N_9087);
or UO_458 (O_458,N_9593,N_8583);
nor UO_459 (O_459,N_6140,N_5184);
nand UO_460 (O_460,N_6969,N_7148);
and UO_461 (O_461,N_5188,N_9795);
or UO_462 (O_462,N_5092,N_7211);
or UO_463 (O_463,N_9148,N_9444);
or UO_464 (O_464,N_8604,N_7656);
nand UO_465 (O_465,N_5257,N_6038);
nor UO_466 (O_466,N_8322,N_9449);
nor UO_467 (O_467,N_5814,N_8073);
nor UO_468 (O_468,N_8635,N_9682);
nor UO_469 (O_469,N_9663,N_8191);
and UO_470 (O_470,N_6115,N_8231);
nor UO_471 (O_471,N_9462,N_9487);
or UO_472 (O_472,N_5613,N_8124);
and UO_473 (O_473,N_8216,N_8625);
nand UO_474 (O_474,N_7708,N_9368);
nand UO_475 (O_475,N_8864,N_6521);
nor UO_476 (O_476,N_5852,N_6237);
nor UO_477 (O_477,N_5204,N_9750);
or UO_478 (O_478,N_7616,N_7175);
and UO_479 (O_479,N_6314,N_9254);
or UO_480 (O_480,N_9446,N_5506);
or UO_481 (O_481,N_7382,N_5967);
nand UO_482 (O_482,N_6990,N_7084);
or UO_483 (O_483,N_5714,N_5887);
or UO_484 (O_484,N_8408,N_7204);
and UO_485 (O_485,N_6982,N_9551);
or UO_486 (O_486,N_5524,N_7851);
nor UO_487 (O_487,N_5380,N_5063);
and UO_488 (O_488,N_5231,N_9312);
nor UO_489 (O_489,N_6044,N_5387);
nand UO_490 (O_490,N_7553,N_7797);
nand UO_491 (O_491,N_8492,N_6661);
or UO_492 (O_492,N_6491,N_7155);
or UO_493 (O_493,N_6753,N_6119);
nor UO_494 (O_494,N_6720,N_5709);
xor UO_495 (O_495,N_6076,N_8051);
or UO_496 (O_496,N_8001,N_7634);
nor UO_497 (O_497,N_7526,N_8534);
nand UO_498 (O_498,N_8120,N_9063);
and UO_499 (O_499,N_6490,N_9959);
or UO_500 (O_500,N_5587,N_6967);
xnor UO_501 (O_501,N_7244,N_9014);
and UO_502 (O_502,N_9548,N_6809);
or UO_503 (O_503,N_9565,N_5394);
or UO_504 (O_504,N_8172,N_8889);
and UO_505 (O_505,N_7638,N_5273);
nand UO_506 (O_506,N_6868,N_7286);
or UO_507 (O_507,N_8094,N_9006);
and UO_508 (O_508,N_9658,N_6126);
or UO_509 (O_509,N_8117,N_9711);
nand UO_510 (O_510,N_8660,N_9555);
nand UO_511 (O_511,N_8232,N_7311);
nand UO_512 (O_512,N_8268,N_6230);
and UO_513 (O_513,N_9245,N_5375);
nand UO_514 (O_514,N_5848,N_5604);
or UO_515 (O_515,N_5457,N_8057);
or UO_516 (O_516,N_6861,N_5686);
or UO_517 (O_517,N_9886,N_6200);
nand UO_518 (O_518,N_9953,N_5971);
and UO_519 (O_519,N_5142,N_9256);
nand UO_520 (O_520,N_7483,N_9763);
or UO_521 (O_521,N_9797,N_8277);
and UO_522 (O_522,N_8724,N_6308);
and UO_523 (O_523,N_8987,N_9218);
or UO_524 (O_524,N_6637,N_8954);
nor UO_525 (O_525,N_7836,N_6511);
nor UO_526 (O_526,N_9232,N_8242);
nand UO_527 (O_527,N_9404,N_9022);
or UO_528 (O_528,N_9056,N_5817);
and UO_529 (O_529,N_5913,N_9231);
and UO_530 (O_530,N_5758,N_5303);
nand UO_531 (O_531,N_5786,N_5944);
or UO_532 (O_532,N_5939,N_9748);
nor UO_533 (O_533,N_6853,N_7395);
and UO_534 (O_534,N_9447,N_5544);
nand UO_535 (O_535,N_8765,N_6553);
and UO_536 (O_536,N_9456,N_8316);
nor UO_537 (O_537,N_7670,N_5015);
or UO_538 (O_538,N_8472,N_5622);
or UO_539 (O_539,N_5267,N_9158);
nor UO_540 (O_540,N_5665,N_8407);
and UO_541 (O_541,N_9773,N_6431);
nand UO_542 (O_542,N_6566,N_6286);
xnor UO_543 (O_543,N_6924,N_7723);
nand UO_544 (O_544,N_7540,N_7561);
nor UO_545 (O_545,N_6381,N_6488);
and UO_546 (O_546,N_5901,N_7724);
and UO_547 (O_547,N_9840,N_6174);
nand UO_548 (O_548,N_5774,N_9998);
and UO_549 (O_549,N_5155,N_5135);
or UO_550 (O_550,N_6555,N_8204);
and UO_551 (O_551,N_9396,N_7485);
nand UO_552 (O_552,N_9874,N_5960);
and UO_553 (O_553,N_6917,N_8088);
or UO_554 (O_554,N_5879,N_9945);
nand UO_555 (O_555,N_5919,N_6477);
nor UO_556 (O_556,N_8661,N_8342);
and UO_557 (O_557,N_6900,N_5280);
or UO_558 (O_558,N_9964,N_6104);
or UO_559 (O_559,N_5080,N_5274);
nand UO_560 (O_560,N_7349,N_8454);
nor UO_561 (O_561,N_9163,N_6424);
and UO_562 (O_562,N_7635,N_9159);
nand UO_563 (O_563,N_8930,N_6596);
and UO_564 (O_564,N_9885,N_5588);
and UO_565 (O_565,N_7912,N_7863);
and UO_566 (O_566,N_5272,N_5385);
nand UO_567 (O_567,N_5508,N_9929);
or UO_568 (O_568,N_7215,N_6882);
xnor UO_569 (O_569,N_9765,N_7153);
nor UO_570 (O_570,N_9764,N_9857);
or UO_571 (O_571,N_5038,N_6939);
xnor UO_572 (O_572,N_8272,N_6847);
nor UO_573 (O_573,N_6679,N_5803);
nand UO_574 (O_574,N_7179,N_5954);
nand UO_575 (O_575,N_6617,N_6015);
nor UO_576 (O_576,N_7304,N_5756);
nand UO_577 (O_577,N_7501,N_8352);
nor UO_578 (O_578,N_9123,N_9291);
xnor UO_579 (O_579,N_5181,N_8405);
nor UO_580 (O_580,N_8880,N_7271);
nor UO_581 (O_581,N_6821,N_5534);
xnor UO_582 (O_582,N_7445,N_5757);
nor UO_583 (O_583,N_9622,N_5061);
nand UO_584 (O_584,N_8958,N_5443);
and UO_585 (O_585,N_7494,N_9859);
nor UO_586 (O_586,N_7729,N_7048);
nor UO_587 (O_587,N_7965,N_9154);
nor UO_588 (O_588,N_5674,N_8705);
or UO_589 (O_589,N_8024,N_8377);
nand UO_590 (O_590,N_6945,N_8964);
and UO_591 (O_591,N_7784,N_7301);
and UO_592 (O_592,N_8433,N_6667);
and UO_593 (O_593,N_9696,N_8614);
nor UO_594 (O_594,N_5871,N_9520);
nor UO_595 (O_595,N_8951,N_9017);
or UO_596 (O_596,N_7067,N_6423);
or UO_597 (O_597,N_6856,N_8298);
or UO_598 (O_598,N_7749,N_7217);
nand UO_599 (O_599,N_9015,N_5478);
or UO_600 (O_600,N_8428,N_7056);
nor UO_601 (O_601,N_8041,N_9369);
and UO_602 (O_602,N_7808,N_7146);
and UO_603 (O_603,N_9751,N_7426);
nand UO_604 (O_604,N_8892,N_6041);
or UO_605 (O_605,N_5788,N_9651);
or UO_606 (O_606,N_6993,N_6627);
and UO_607 (O_607,N_8780,N_6721);
and UO_608 (O_608,N_9237,N_6102);
nor UO_609 (O_609,N_5028,N_5057);
nor UO_610 (O_610,N_5517,N_6694);
and UO_611 (O_611,N_6626,N_6651);
nor UO_612 (O_612,N_9641,N_7588);
or UO_613 (O_613,N_7247,N_6941);
nor UO_614 (O_614,N_9140,N_5005);
nor UO_615 (O_615,N_7188,N_8045);
and UO_616 (O_616,N_9336,N_7019);
and UO_617 (O_617,N_8738,N_7476);
or UO_618 (O_618,N_5240,N_8503);
nor UO_619 (O_619,N_7322,N_7887);
nand UO_620 (O_620,N_7891,N_9260);
nor UO_621 (O_621,N_6862,N_9263);
or UO_622 (O_622,N_7073,N_7694);
nand UO_623 (O_623,N_8577,N_8929);
and UO_624 (O_624,N_5959,N_8229);
or UO_625 (O_625,N_5493,N_7294);
nor UO_626 (O_626,N_6338,N_5058);
nand UO_627 (O_627,N_8647,N_9209);
nand UO_628 (O_628,N_9514,N_8443);
and UO_629 (O_629,N_7288,N_6166);
nor UO_630 (O_630,N_7826,N_6813);
nand UO_631 (O_631,N_8511,N_7539);
nor UO_632 (O_632,N_7980,N_5086);
nor UO_633 (O_633,N_7819,N_6183);
and UO_634 (O_634,N_8021,N_5014);
nor UO_635 (O_635,N_8608,N_7577);
or UO_636 (O_636,N_5199,N_6886);
or UO_637 (O_637,N_9776,N_6438);
or UO_638 (O_638,N_6891,N_5175);
xnor UO_639 (O_639,N_8734,N_5107);
xnor UO_640 (O_640,N_9122,N_9782);
and UO_641 (O_641,N_5505,N_6530);
nand UO_642 (O_642,N_5671,N_8218);
xnor UO_643 (O_643,N_9579,N_9309);
nor UO_644 (O_644,N_6322,N_9019);
nor UO_645 (O_645,N_7620,N_8017);
nor UO_646 (O_646,N_7203,N_6630);
xor UO_647 (O_647,N_5683,N_6474);
nor UO_648 (O_648,N_8258,N_5560);
or UO_649 (O_649,N_5727,N_7387);
or UO_650 (O_650,N_9829,N_7990);
nand UO_651 (O_651,N_5331,N_6892);
nand UO_652 (O_652,N_7318,N_7154);
and UO_653 (O_653,N_5225,N_5419);
nand UO_654 (O_654,N_7306,N_5698);
nor UO_655 (O_655,N_6311,N_6296);
nor UO_656 (O_656,N_6295,N_8183);
nor UO_657 (O_657,N_8637,N_7354);
nor UO_658 (O_658,N_6145,N_8915);
or UO_659 (O_659,N_5647,N_8392);
nand UO_660 (O_660,N_9787,N_9799);
or UO_661 (O_661,N_8778,N_8058);
nand UO_662 (O_662,N_6607,N_7559);
and UO_663 (O_663,N_6699,N_5060);
nand UO_664 (O_664,N_7722,N_9066);
nand UO_665 (O_665,N_7194,N_9517);
nand UO_666 (O_666,N_8803,N_9096);
or UO_667 (O_667,N_5325,N_5136);
or UO_668 (O_668,N_7072,N_5447);
nor UO_669 (O_669,N_8043,N_5985);
or UO_670 (O_670,N_9616,N_6912);
nand UO_671 (O_671,N_7523,N_8369);
nand UO_672 (O_672,N_7229,N_7584);
and UO_673 (O_673,N_6543,N_6936);
or UO_674 (O_674,N_8111,N_5540);
or UO_675 (O_675,N_6691,N_7794);
and UO_676 (O_676,N_9506,N_9931);
nand UO_677 (O_677,N_5601,N_5884);
and UO_678 (O_678,N_9550,N_6938);
nor UO_679 (O_679,N_6022,N_9698);
nand UO_680 (O_680,N_6110,N_9823);
or UO_681 (O_681,N_8815,N_8005);
or UO_682 (O_682,N_5752,N_5981);
nand UO_683 (O_683,N_7160,N_6561);
and UO_684 (O_684,N_7087,N_8388);
xnor UO_685 (O_685,N_6262,N_7167);
nand UO_686 (O_686,N_6021,N_6079);
or UO_687 (O_687,N_8655,N_6928);
or UO_688 (O_688,N_5398,N_6603);
or UO_689 (O_689,N_6390,N_9921);
and UO_690 (O_690,N_9434,N_7511);
or UO_691 (O_691,N_9405,N_6404);
and UO_692 (O_692,N_7647,N_5558);
or UO_693 (O_693,N_9705,N_6840);
or UO_694 (O_694,N_9640,N_5964);
nand UO_695 (O_695,N_9217,N_7411);
and UO_696 (O_696,N_6516,N_9838);
or UO_697 (O_697,N_5381,N_5362);
and UO_698 (O_698,N_5612,N_5361);
nor UO_699 (O_699,N_8157,N_5109);
nand UO_700 (O_700,N_5027,N_7799);
xor UO_701 (O_701,N_8831,N_9314);
nand UO_702 (O_702,N_7783,N_5991);
or UO_703 (O_703,N_9849,N_6722);
or UO_704 (O_704,N_9370,N_6879);
nor UO_705 (O_705,N_8800,N_7313);
nand UO_706 (O_706,N_5607,N_8135);
nand UO_707 (O_707,N_5187,N_9629);
nand UO_708 (O_708,N_8426,N_8616);
nor UO_709 (O_709,N_7703,N_6935);
or UO_710 (O_710,N_8287,N_9694);
nand UO_711 (O_711,N_7643,N_5658);
nor UO_712 (O_712,N_7428,N_7151);
nor UO_713 (O_713,N_6605,N_5317);
or UO_714 (O_714,N_7254,N_9324);
or UO_715 (O_715,N_9344,N_6953);
nor UO_716 (O_716,N_8580,N_5355);
and UO_717 (O_717,N_9848,N_6396);
nor UO_718 (O_718,N_6996,N_9813);
and UO_719 (O_719,N_8484,N_6852);
and UO_720 (O_720,N_7094,N_8728);
and UO_721 (O_721,N_5519,N_5663);
nand UO_722 (O_722,N_7407,N_8887);
nand UO_723 (O_723,N_5128,N_7531);
and UO_724 (O_724,N_7213,N_7885);
nand UO_725 (O_725,N_8563,N_5451);
or UO_726 (O_726,N_8170,N_8072);
nor UO_727 (O_727,N_5851,N_6643);
or UO_728 (O_728,N_9453,N_5295);
xor UO_729 (O_729,N_8262,N_7549);
nand UO_730 (O_730,N_7005,N_5434);
or UO_731 (O_731,N_8624,N_6340);
nor UO_732 (O_732,N_8946,N_7790);
nor UO_733 (O_733,N_5300,N_8318);
or UO_734 (O_734,N_8213,N_5012);
or UO_735 (O_735,N_5082,N_5754);
or UO_736 (O_736,N_9374,N_8581);
or UO_737 (O_737,N_6382,N_7904);
xor UO_738 (O_738,N_9101,N_7161);
and UO_739 (O_739,N_6955,N_8927);
or UO_740 (O_740,N_6081,N_9890);
and UO_741 (O_741,N_6213,N_6421);
nand UO_742 (O_742,N_9228,N_9803);
or UO_743 (O_743,N_6895,N_8851);
xor UO_744 (O_744,N_6756,N_8542);
and UO_745 (O_745,N_9229,N_7742);
nor UO_746 (O_746,N_6007,N_6735);
and UO_747 (O_747,N_9315,N_6934);
or UO_748 (O_748,N_5278,N_5369);
and UO_749 (O_749,N_9166,N_5071);
nor UO_750 (O_750,N_7660,N_9714);
and UO_751 (O_751,N_8446,N_6838);
nor UO_752 (O_752,N_6380,N_8886);
or UO_753 (O_753,N_5347,N_5710);
nor UO_754 (O_754,N_9634,N_5891);
or UO_755 (O_755,N_8943,N_7890);
nor UO_756 (O_756,N_7427,N_8003);
or UO_757 (O_757,N_9601,N_5888);
or UO_758 (O_758,N_8584,N_5666);
nor UO_759 (O_759,N_9607,N_5906);
nor UO_760 (O_760,N_8155,N_5667);
and UO_761 (O_761,N_5495,N_5681);
or UO_762 (O_762,N_6207,N_5025);
and UO_763 (O_763,N_6011,N_5088);
or UO_764 (O_764,N_5907,N_9361);
nor UO_765 (O_765,N_6817,N_6796);
nor UO_766 (O_766,N_5314,N_8389);
nor UO_767 (O_767,N_7208,N_6238);
nor UO_768 (O_768,N_8331,N_5147);
or UO_769 (O_769,N_8165,N_7855);
nor UO_770 (O_770,N_6393,N_9356);
nor UO_771 (O_771,N_9195,N_8050);
nand UO_772 (O_772,N_8427,N_9692);
nand UO_773 (O_773,N_5922,N_5958);
or UO_774 (O_774,N_8846,N_8812);
nor UO_775 (O_775,N_6748,N_6806);
nor UO_776 (O_776,N_5937,N_9061);
nor UO_777 (O_777,N_9278,N_7777);
and UO_778 (O_778,N_9673,N_9221);
nand UO_779 (O_779,N_7969,N_6470);
and UO_780 (O_780,N_8656,N_6411);
and UO_781 (O_781,N_6669,N_6356);
nor UO_782 (O_782,N_8481,N_9109);
and UO_783 (O_783,N_9407,N_9516);
and UO_784 (O_784,N_7705,N_9834);
nor UO_785 (O_785,N_8463,N_7541);
nand UO_786 (O_786,N_5856,N_7591);
xor UO_787 (O_787,N_6182,N_9118);
nor UO_788 (O_788,N_7686,N_5837);
nand UO_789 (O_789,N_5943,N_8696);
xor UO_790 (O_790,N_9040,N_8719);
or UO_791 (O_791,N_5861,N_7470);
nor UO_792 (O_792,N_8934,N_8727);
and UO_793 (O_793,N_5047,N_9878);
nor UO_794 (O_794,N_6155,N_7988);
and UO_795 (O_795,N_7497,N_9952);
or UO_796 (O_796,N_5644,N_8865);
nand UO_797 (O_797,N_6087,N_8726);
nand UO_798 (O_798,N_6033,N_6232);
or UO_799 (O_799,N_9378,N_8629);
and UO_800 (O_800,N_7791,N_5768);
xnor UO_801 (O_801,N_9854,N_7966);
and UO_802 (O_802,N_9013,N_8941);
or UO_803 (O_803,N_8077,N_8419);
nand UO_804 (O_804,N_7028,N_7012);
and UO_805 (O_805,N_7053,N_7835);
nand UO_806 (O_806,N_8981,N_8161);
or UO_807 (O_807,N_9961,N_8866);
xnor UO_808 (O_808,N_7357,N_5761);
nand UO_809 (O_809,N_5209,N_5543);
nand UO_810 (O_810,N_5859,N_9152);
or UO_811 (O_811,N_5914,N_9224);
and UO_812 (O_812,N_6370,N_9307);
or UO_813 (O_813,N_5030,N_9146);
nor UO_814 (O_814,N_5782,N_8490);
and UO_815 (O_815,N_8901,N_8628);
or UO_816 (O_816,N_9552,N_7651);
nor UO_817 (O_817,N_5477,N_5747);
or UO_818 (O_818,N_6205,N_8289);
and UO_819 (O_819,N_7119,N_7065);
or UO_820 (O_820,N_7573,N_8474);
and UO_821 (O_821,N_6318,N_9499);
and UO_822 (O_822,N_7232,N_5083);
and UO_823 (O_823,N_5265,N_9652);
nor UO_824 (O_824,N_9635,N_8205);
xnor UO_825 (O_825,N_8908,N_8805);
or UO_826 (O_826,N_6992,N_5111);
nand UO_827 (O_827,N_8367,N_7321);
and UO_828 (O_828,N_6780,N_5707);
and UO_829 (O_829,N_9522,N_9310);
nand UO_830 (O_830,N_9036,N_7030);
or UO_831 (O_831,N_8047,N_9924);
and UO_832 (O_832,N_8916,N_9606);
nor UO_833 (O_833,N_5969,N_8861);
nand UO_834 (O_834,N_9887,N_6480);
nor UO_835 (O_835,N_7658,N_7480);
or UO_836 (O_836,N_5850,N_7228);
nor UO_837 (O_837,N_7895,N_5951);
nand UO_838 (O_838,N_6336,N_6702);
or UO_839 (O_839,N_5161,N_5892);
or UO_840 (O_840,N_6025,N_7009);
and UO_841 (O_841,N_5296,N_8950);
nor UO_842 (O_842,N_7811,N_7615);
or UO_843 (O_843,N_5818,N_9129);
nand UO_844 (O_844,N_7405,N_9675);
and UO_845 (O_845,N_7140,N_8917);
nand UO_846 (O_846,N_9333,N_8550);
nor UO_847 (O_847,N_9738,N_6427);
or UO_848 (O_848,N_7190,N_5428);
nor UO_849 (O_849,N_7798,N_7925);
and UO_850 (O_850,N_6305,N_7672);
and UO_851 (O_851,N_8307,N_5046);
nand UO_852 (O_852,N_8926,N_6287);
or UO_853 (O_853,N_9276,N_9298);
nor UO_854 (O_854,N_9637,N_7650);
and UO_855 (O_855,N_7644,N_6906);
nand UO_856 (O_856,N_8251,N_8430);
nor UO_857 (O_857,N_5828,N_5784);
nor UO_858 (O_858,N_8940,N_8030);
nor UO_859 (O_859,N_9927,N_8952);
and UO_860 (O_860,N_8282,N_5207);
nor UO_861 (O_861,N_7892,N_7932);
or UO_862 (O_862,N_5292,N_9296);
xor UO_863 (O_863,N_8130,N_5235);
and UO_864 (O_864,N_5031,N_9327);
nor UO_865 (O_865,N_8688,N_8595);
nor UO_866 (O_866,N_7396,N_6164);
or UO_867 (O_867,N_9722,N_9668);
nand UO_868 (O_868,N_5217,N_5229);
or UO_869 (O_869,N_8054,N_9348);
nand UO_870 (O_870,N_6150,N_9332);
or UO_871 (O_871,N_6017,N_6323);
nand UO_872 (O_872,N_8154,N_9060);
or UO_873 (O_873,N_6713,N_6408);
and UO_874 (O_874,N_8211,N_8706);
nor UO_875 (O_875,N_9501,N_8244);
and UO_876 (O_876,N_7315,N_7451);
xnor UO_877 (O_877,N_7149,N_6109);
or UO_878 (O_878,N_9725,N_9971);
or UO_879 (O_879,N_8853,N_5863);
or UO_880 (O_880,N_7775,N_5384);
nor UO_881 (O_881,N_5807,N_5575);
nor UO_882 (O_882,N_6386,N_9100);
or UO_883 (O_883,N_5794,N_5821);
nand UO_884 (O_884,N_5154,N_8293);
or UO_885 (O_885,N_8327,N_7959);
and UO_886 (O_886,N_6560,N_5322);
and UO_887 (O_887,N_7241,N_7505);
or UO_888 (O_888,N_6890,N_9818);
and UO_889 (O_889,N_7314,N_6333);
nand UO_890 (O_890,N_8911,N_8966);
nand UO_891 (O_891,N_9223,N_7751);
and UO_892 (O_892,N_6508,N_5635);
nand UO_893 (O_893,N_6378,N_6298);
nand UO_894 (O_894,N_7534,N_9867);
and UO_895 (O_895,N_9338,N_5692);
nor UO_896 (O_896,N_5282,N_8822);
nand UO_897 (O_897,N_5917,N_8937);
nand UO_898 (O_898,N_8626,N_6460);
nand UO_899 (O_899,N_9373,N_8206);
nand UO_900 (O_900,N_8125,N_6190);
nand UO_901 (O_901,N_6468,N_8967);
nand UO_902 (O_902,N_7558,N_9416);
or UO_903 (O_903,N_8185,N_5900);
or UO_904 (O_904,N_9684,N_7556);
and UO_905 (O_905,N_8948,N_5751);
or UO_906 (O_906,N_6760,N_6310);
and UO_907 (O_907,N_9262,N_7781);
nor UO_908 (O_908,N_7913,N_9292);
or UO_909 (O_909,N_9286,N_5812);
nand UO_910 (O_910,N_9452,N_7493);
or UO_911 (O_911,N_9880,N_9868);
or UO_912 (O_912,N_8455,N_6134);
and UO_913 (O_913,N_8804,N_6576);
nor UO_914 (O_914,N_8680,N_6827);
and UO_915 (O_915,N_9911,N_5171);
nor UO_916 (O_916,N_9126,N_7732);
nand UO_917 (O_917,N_5371,N_8048);
and UO_918 (O_918,N_7719,N_7578);
nor UO_919 (O_919,N_9759,N_5882);
nor UO_920 (O_920,N_6089,N_8606);
nor UO_921 (O_921,N_8305,N_5690);
nor UO_922 (O_922,N_5962,N_7630);
nand UO_923 (O_923,N_7165,N_6445);
xor UO_924 (O_924,N_8303,N_8895);
and UO_925 (O_925,N_7513,N_8240);
nand UO_926 (O_926,N_7960,N_6755);
and UO_927 (O_927,N_8707,N_8399);
nand UO_928 (O_928,N_5536,N_9470);
nand UO_929 (O_929,N_7113,N_9192);
and UO_930 (O_930,N_9219,N_6871);
or UO_931 (O_931,N_5017,N_9767);
nor UO_932 (O_932,N_7449,N_8788);
nor UO_933 (O_933,N_9115,N_6600);
nand UO_934 (O_934,N_8998,N_8972);
nand UO_935 (O_935,N_5646,N_8646);
or UO_936 (O_936,N_8508,N_5741);
nand UO_937 (O_937,N_5699,N_8847);
nand UO_938 (O_938,N_6366,N_6114);
nand UO_939 (O_939,N_7765,N_9342);
nor UO_940 (O_940,N_8588,N_5632);
nand UO_941 (O_941,N_7242,N_9124);
and UO_942 (O_942,N_6964,N_9299);
nor UO_943 (O_943,N_7628,N_7803);
nor UO_944 (O_944,N_8552,N_5172);
or UO_945 (O_945,N_8423,N_8348);
or UO_946 (O_946,N_6345,N_8202);
or UO_947 (O_947,N_8076,N_6645);
or UO_948 (O_948,N_9093,N_6278);
or UO_949 (O_949,N_6093,N_7875);
and UO_950 (O_950,N_9912,N_9004);
or UO_951 (O_951,N_6715,N_7082);
nor UO_952 (O_952,N_7512,N_6552);
or UO_953 (O_953,N_8823,N_6398);
nor UO_954 (O_954,N_7721,N_7637);
and UO_955 (O_955,N_8996,N_7170);
or UO_956 (O_956,N_9860,N_7471);
or UO_957 (O_957,N_9199,N_8068);
or UO_958 (O_958,N_8008,N_7975);
and UO_959 (O_959,N_8418,N_5523);
or UO_960 (O_960,N_6389,N_9590);
or UO_961 (O_961,N_7103,N_8281);
nand UO_962 (O_962,N_6646,N_9098);
nand UO_963 (O_963,N_7024,N_8321);
and UO_964 (O_964,N_8947,N_5750);
nand UO_965 (O_965,N_9481,N_9757);
nor UO_966 (O_966,N_6425,N_9213);
or UO_967 (O_967,N_8417,N_5805);
xnor UO_968 (O_968,N_7569,N_6976);
nand UO_969 (O_969,N_9613,N_8779);
nand UO_970 (O_970,N_6901,N_8386);
nor UO_971 (O_971,N_5516,N_5696);
or UO_972 (O_972,N_6478,N_7872);
and UO_973 (O_973,N_5308,N_6961);
or UO_974 (O_974,N_9932,N_7289);
or UO_975 (O_975,N_9409,N_8037);
nor UO_976 (O_976,N_9996,N_6658);
nand UO_977 (O_977,N_6249,N_9360);
nor UO_978 (O_978,N_5677,N_6280);
nor UO_979 (O_979,N_9144,N_6216);
xnor UO_980 (O_980,N_5720,N_6703);
nor UO_981 (O_981,N_7489,N_9169);
nand UO_982 (O_982,N_5498,N_5490);
and UO_983 (O_983,N_9626,N_6197);
nand UO_984 (O_984,N_8678,N_9186);
and UO_985 (O_985,N_9954,N_9125);
nand UO_986 (O_986,N_6043,N_8398);
and UO_987 (O_987,N_8022,N_7135);
and UO_988 (O_988,N_6548,N_7623);
or UO_989 (O_989,N_6117,N_7199);
and UO_990 (O_990,N_7457,N_6484);
and UO_991 (O_991,N_7994,N_9519);
or UO_992 (O_992,N_6849,N_9554);
nor UO_993 (O_993,N_8777,N_6211);
or UO_994 (O_994,N_7381,N_8520);
or UO_995 (O_995,N_8603,N_6509);
nor UO_996 (O_996,N_7695,N_5312);
and UO_997 (O_997,N_9562,N_5119);
nand UO_998 (O_998,N_6860,N_8363);
nand UO_999 (O_999,N_6302,N_9600);
nand UO_1000 (O_1000,N_9030,N_8722);
nor UO_1001 (O_1001,N_6987,N_5602);
xnor UO_1002 (O_1002,N_6925,N_7687);
xor UO_1003 (O_1003,N_9941,N_9402);
or UO_1004 (O_1004,N_6153,N_6614);
nand UO_1005 (O_1005,N_6223,N_9633);
and UO_1006 (O_1006,N_5134,N_8462);
xnor UO_1007 (O_1007,N_9542,N_7434);
or UO_1008 (O_1008,N_8437,N_9137);
nor UO_1009 (O_1009,N_8084,N_5056);
nor UO_1010 (O_1010,N_8074,N_5346);
nor UO_1011 (O_1011,N_7282,N_7745);
nor UO_1012 (O_1012,N_5405,N_7340);
and UO_1013 (O_1013,N_5771,N_8748);
nor UO_1014 (O_1014,N_9001,N_8711);
and UO_1015 (O_1015,N_5594,N_6444);
xor UO_1016 (O_1016,N_9380,N_8441);
and UO_1017 (O_1017,N_8414,N_7772);
nand UO_1018 (O_1018,N_7266,N_7527);
and UO_1019 (O_1019,N_6147,N_5024);
and UO_1020 (O_1020,N_8506,N_8942);
and UO_1021 (O_1021,N_5141,N_7681);
or UO_1022 (O_1022,N_7006,N_7691);
nor UO_1023 (O_1023,N_6341,N_9643);
nor UO_1024 (O_1024,N_6675,N_8634);
nand UO_1025 (O_1025,N_8525,N_8808);
or UO_1026 (O_1026,N_6154,N_9644);
or UO_1027 (O_1027,N_9107,N_8570);
nor UO_1028 (O_1028,N_9906,N_5796);
nor UO_1029 (O_1029,N_9021,N_9627);
and UO_1030 (O_1030,N_6893,N_7342);
nand UO_1031 (O_1031,N_8859,N_7345);
or UO_1032 (O_1032,N_8878,N_8697);
nand UO_1033 (O_1033,N_7736,N_6523);
nand UO_1034 (O_1034,N_9747,N_6984);
xnor UO_1035 (O_1035,N_7343,N_7375);
or UO_1036 (O_1036,N_5259,N_5778);
nand UO_1037 (O_1037,N_9176,N_6062);
nor UO_1038 (O_1038,N_6040,N_8069);
or UO_1039 (O_1039,N_8083,N_7801);
nor UO_1040 (O_1040,N_7462,N_8918);
nor UO_1041 (O_1041,N_5555,N_8312);
nand UO_1042 (O_1042,N_6881,N_6361);
nand UO_1043 (O_1043,N_6260,N_7287);
or UO_1044 (O_1044,N_9583,N_8731);
nand UO_1045 (O_1045,N_9204,N_9636);
and UO_1046 (O_1046,N_5905,N_6980);
or UO_1047 (O_1047,N_9728,N_7185);
or UO_1048 (O_1048,N_8817,N_5236);
and UO_1049 (O_1049,N_6962,N_5617);
nor UO_1050 (O_1050,N_7746,N_8961);
or UO_1051 (O_1051,N_5359,N_9984);
nand UO_1052 (O_1052,N_9018,N_5348);
and UO_1053 (O_1053,N_8065,N_8196);
nor UO_1054 (O_1054,N_5176,N_7488);
nor UO_1055 (O_1055,N_7914,N_8522);
nor UO_1056 (O_1056,N_6664,N_8371);
or UO_1057 (O_1057,N_5655,N_5117);
and UO_1058 (O_1058,N_8658,N_8988);
or UO_1059 (O_1059,N_7341,N_5492);
nand UO_1060 (O_1060,N_9588,N_8089);
nor UO_1061 (O_1061,N_7629,N_7592);
and UO_1062 (O_1062,N_7368,N_8524);
or UO_1063 (O_1063,N_7754,N_6850);
nand UO_1064 (O_1064,N_5338,N_8184);
or UO_1065 (O_1065,N_6979,N_7663);
or UO_1066 (O_1066,N_6692,N_8785);
xnor UO_1067 (O_1067,N_9587,N_6187);
or UO_1068 (O_1068,N_9029,N_7117);
and UO_1069 (O_1069,N_7717,N_5982);
nand UO_1070 (O_1070,N_5453,N_5764);
and UO_1071 (O_1071,N_5007,N_6567);
nor UO_1072 (O_1072,N_9234,N_8774);
nand UO_1073 (O_1073,N_9490,N_7779);
and UO_1074 (O_1074,N_8507,N_7923);
nor UO_1075 (O_1075,N_8749,N_9814);
nor UO_1076 (O_1076,N_6458,N_5483);
nand UO_1077 (O_1077,N_8260,N_9113);
nand UO_1078 (O_1078,N_8031,N_9459);
nand UO_1079 (O_1079,N_7320,N_9024);
or UO_1080 (O_1080,N_7478,N_7547);
or UO_1081 (O_1081,N_8935,N_8995);
and UO_1082 (O_1082,N_8611,N_8333);
nor UO_1083 (O_1083,N_5318,N_6221);
nand UO_1084 (O_1084,N_5777,N_7402);
nor UO_1085 (O_1085,N_9657,N_6546);
nor UO_1086 (O_1086,N_6294,N_6339);
or UO_1087 (O_1087,N_6783,N_8528);
nand UO_1088 (O_1088,N_5950,N_6116);
or UO_1089 (O_1089,N_8971,N_5151);
nor UO_1090 (O_1090,N_5770,N_9055);
nor UO_1091 (O_1091,N_8029,N_5198);
nor UO_1092 (O_1092,N_7417,N_6413);
or UO_1093 (O_1093,N_5904,N_7725);
nand UO_1094 (O_1094,N_8353,N_5592);
and UO_1095 (O_1095,N_8871,N_7308);
and UO_1096 (O_1096,N_6525,N_9345);
or UO_1097 (O_1097,N_9727,N_6078);
nor UO_1098 (O_1098,N_7671,N_9534);
nand UO_1099 (O_1099,N_7274,N_7080);
or UO_1100 (O_1100,N_5169,N_6701);
and UO_1101 (O_1101,N_9461,N_8751);
nor UO_1102 (O_1102,N_6156,N_5037);
and UO_1103 (O_1103,N_5685,N_7202);
and UO_1104 (O_1104,N_7524,N_5358);
and UO_1105 (O_1105,N_5158,N_7363);
and UO_1106 (O_1106,N_7639,N_6368);
nand UO_1107 (O_1107,N_5305,N_7409);
nor UO_1108 (O_1108,N_7787,N_8810);
nor UO_1109 (O_1109,N_7120,N_5753);
nand UO_1110 (O_1110,N_6387,N_9752);
or UO_1111 (O_1111,N_9526,N_5669);
nor UO_1112 (O_1112,N_5143,N_8166);
or UO_1113 (O_1113,N_9190,N_7115);
and UO_1114 (O_1114,N_8143,N_8040);
or UO_1115 (O_1115,N_5855,N_6042);
nand UO_1116 (O_1116,N_7856,N_8411);
nand UO_1117 (O_1117,N_9120,N_5464);
nor UO_1118 (O_1118,N_7126,N_6009);
nand UO_1119 (O_1119,N_9280,N_9825);
and UO_1120 (O_1120,N_7377,N_5980);
nor UO_1121 (O_1121,N_9925,N_6874);
and UO_1122 (O_1122,N_6167,N_7755);
nor UO_1123 (O_1123,N_8366,N_5252);
and UO_1124 (O_1124,N_5574,N_5583);
nand UO_1125 (O_1125,N_5535,N_7014);
nand UO_1126 (O_1126,N_9781,N_9780);
nand UO_1127 (O_1127,N_9667,N_5738);
or UO_1128 (O_1128,N_7933,N_9317);
and UO_1129 (O_1129,N_5590,N_9432);
nor UO_1130 (O_1130,N_8638,N_6910);
nor UO_1131 (O_1131,N_9576,N_5377);
xnor UO_1132 (O_1132,N_5614,N_6352);
and UO_1133 (O_1133,N_8687,N_9843);
or UO_1134 (O_1134,N_5551,N_6864);
nor UO_1135 (O_1135,N_5122,N_7619);
nor UO_1136 (O_1136,N_5903,N_8358);
nand UO_1137 (O_1137,N_7532,N_6746);
nand UO_1138 (O_1138,N_6463,N_7657);
or UO_1139 (O_1139,N_6002,N_9305);
or UO_1140 (O_1140,N_7373,N_5072);
nor UO_1141 (O_1141,N_6971,N_7867);
or UO_1142 (O_1142,N_9639,N_5511);
nor UO_1143 (O_1143,N_7720,N_6379);
or UO_1144 (O_1144,N_5838,N_8977);
nor UO_1145 (O_1145,N_8270,N_9020);
nor UO_1146 (O_1146,N_9992,N_5874);
nand UO_1147 (O_1147,N_8968,N_9207);
or UO_1148 (O_1148,N_6775,N_5563);
or UO_1149 (O_1149,N_7897,N_6218);
or UO_1150 (O_1150,N_9424,N_5424);
nand UO_1151 (O_1151,N_5328,N_6644);
and UO_1152 (O_1152,N_7316,N_6492);
nand UO_1153 (O_1153,N_5596,N_8121);
nand UO_1154 (O_1154,N_6909,N_6823);
nand UO_1155 (O_1155,N_7081,N_7181);
nor UO_1156 (O_1156,N_9732,N_8494);
nand UO_1157 (O_1157,N_8023,N_5078);
nor UO_1158 (O_1158,N_9515,N_9586);
nand UO_1159 (O_1159,N_6621,N_8586);
nand UO_1160 (O_1160,N_5629,N_6896);
nand UO_1161 (O_1161,N_8200,N_6077);
or UO_1162 (O_1162,N_5810,N_9023);
nor UO_1163 (O_1163,N_5636,N_7205);
nor UO_1164 (O_1164,N_8341,N_6487);
or UO_1165 (O_1165,N_6954,N_8223);
or UO_1166 (O_1166,N_5216,N_6320);
and UO_1167 (O_1167,N_7843,N_7011);
or UO_1168 (O_1168,N_6106,N_8596);
nand UO_1169 (O_1169,N_6960,N_5880);
and UO_1170 (O_1170,N_6505,N_8598);
nand UO_1171 (O_1171,N_7007,N_9426);
and UO_1172 (O_1172,N_7649,N_7390);
nor UO_1173 (O_1173,N_7397,N_7295);
nor UO_1174 (O_1174,N_5152,N_9546);
xnor UO_1175 (O_1175,N_5365,N_5748);
nand UO_1176 (O_1176,N_9304,N_9703);
and UO_1177 (O_1177,N_8979,N_6653);
nand UO_1178 (O_1178,N_5254,N_7222);
nand UO_1179 (O_1179,N_7394,N_7233);
xor UO_1180 (O_1180,N_6006,N_5512);
xor UO_1181 (O_1181,N_6622,N_7285);
or UO_1182 (O_1182,N_5416,N_7124);
or UO_1183 (O_1183,N_7760,N_6210);
or UO_1184 (O_1184,N_8802,N_7859);
nand UO_1185 (O_1185,N_9610,N_9365);
and UO_1186 (O_1186,N_6401,N_9940);
nand UO_1187 (O_1187,N_7456,N_7636);
or UO_1188 (O_1188,N_5857,N_6674);
nor UO_1189 (O_1189,N_7255,N_5936);
and UO_1190 (O_1190,N_5684,N_9603);
or UO_1191 (O_1191,N_5438,N_7659);
and UO_1192 (O_1192,N_8715,N_8378);
or UO_1193 (O_1193,N_7587,N_6610);
nor UO_1194 (O_1194,N_5363,N_5724);
or UO_1195 (O_1195,N_6534,N_7793);
nand UO_1196 (O_1196,N_8544,N_9210);
nor UO_1197 (O_1197,N_7802,N_7763);
or UO_1198 (O_1198,N_7473,N_8835);
or UO_1199 (O_1199,N_5397,N_9389);
and UO_1200 (O_1200,N_5997,N_9721);
and UO_1201 (O_1201,N_7138,N_6803);
nor UO_1202 (O_1202,N_6706,N_8391);
nand UO_1203 (O_1203,N_9540,N_5591);
and UO_1204 (O_1204,N_8382,N_6001);
or UO_1205 (O_1205,N_7008,N_8153);
and UO_1206 (O_1206,N_5132,N_7152);
nor UO_1207 (O_1207,N_5899,N_5316);
and UO_1208 (O_1208,N_5059,N_6773);
and UO_1209 (O_1209,N_6113,N_5923);
nor UO_1210 (O_1210,N_5319,N_7069);
or UO_1211 (O_1211,N_6750,N_6631);
xnor UO_1212 (O_1212,N_9920,N_5290);
nor UO_1213 (O_1213,N_6898,N_6222);
or UO_1214 (O_1214,N_6432,N_6659);
nand UO_1215 (O_1215,N_9070,N_5885);
nand UO_1216 (O_1216,N_6395,N_5076);
nand UO_1217 (O_1217,N_6268,N_6075);
and UO_1218 (O_1218,N_5640,N_9898);
and UO_1219 (O_1219,N_9258,N_8291);
and UO_1220 (O_1220,N_5862,N_8285);
nand UO_1221 (O_1221,N_9351,N_8615);
and UO_1222 (O_1222,N_9033,N_6189);
nor UO_1223 (O_1223,N_6289,N_8821);
and UO_1224 (O_1224,N_8162,N_7726);
nand UO_1225 (O_1225,N_8723,N_6099);
and UO_1226 (O_1226,N_9830,N_5732);
nor UO_1227 (O_1227,N_7225,N_6005);
nand UO_1228 (O_1228,N_6575,N_6834);
and UO_1229 (O_1229,N_7253,N_5977);
nand UO_1230 (O_1230,N_7145,N_6243);
and UO_1231 (O_1231,N_6161,N_6105);
nand UO_1232 (O_1232,N_5947,N_8406);
nor UO_1233 (O_1233,N_6176,N_9604);
or UO_1234 (O_1234,N_9222,N_6493);
and UO_1235 (O_1235,N_5952,N_6275);
nand UO_1236 (O_1236,N_9783,N_8761);
and UO_1237 (O_1237,N_5323,N_6233);
nand UO_1238 (O_1238,N_8332,N_6875);
nor UO_1239 (O_1239,N_8623,N_6514);
or UO_1240 (O_1240,N_8092,N_7332);
nor UO_1241 (O_1241,N_6859,N_8214);
and UO_1242 (O_1242,N_8565,N_9383);
and UO_1243 (O_1243,N_8932,N_9671);
and UO_1244 (O_1244,N_7621,N_8090);
nand UO_1245 (O_1245,N_8983,N_8187);
nand UO_1246 (O_1246,N_5515,N_9899);
nand UO_1247 (O_1247,N_9785,N_5286);
nand UO_1248 (O_1248,N_5660,N_9947);
or UO_1249 (O_1249,N_9411,N_7545);
nor UO_1250 (O_1250,N_5743,N_8315);
xor UO_1251 (O_1251,N_9127,N_6915);
or UO_1252 (O_1252,N_9349,N_9266);
nand UO_1253 (O_1253,N_6192,N_7903);
nand UO_1254 (O_1254,N_6782,N_7418);
and UO_1255 (O_1255,N_5251,N_6422);
or UO_1256 (O_1256,N_5001,N_5174);
or UO_1257 (O_1257,N_7076,N_7776);
nor UO_1258 (O_1258,N_6550,N_6537);
nor UO_1259 (O_1259,N_6535,N_7822);
nor UO_1260 (O_1260,N_5125,N_7884);
nand UO_1261 (O_1261,N_8960,N_9131);
and UO_1262 (O_1262,N_8575,N_7174);
or UO_1263 (O_1263,N_6704,N_8403);
nand UO_1264 (O_1264,N_7293,N_8569);
nand UO_1265 (O_1265,N_8829,N_5763);
nor UO_1266 (O_1266,N_9541,N_7950);
and UO_1267 (O_1267,N_9441,N_8238);
nor UO_1268 (O_1268,N_8914,N_8006);
or UO_1269 (O_1269,N_7324,N_5244);
and UO_1270 (O_1270,N_5036,N_9766);
nand UO_1271 (O_1271,N_6337,N_6084);
or UO_1272 (O_1272,N_8955,N_9901);
nor UO_1273 (O_1273,N_8890,N_9039);
nand UO_1274 (O_1274,N_9134,N_9808);
and UO_1275 (O_1275,N_6685,N_6299);
nor UO_1276 (O_1276,N_9058,N_5388);
and UO_1277 (O_1277,N_5772,N_7624);
nor UO_1278 (O_1278,N_7604,N_6428);
and UO_1279 (O_1279,N_5643,N_9888);
nor UO_1280 (O_1280,N_5532,N_7652);
and UO_1281 (O_1281,N_8485,N_6696);
nand UO_1282 (O_1282,N_6016,N_9352);
or UO_1283 (O_1283,N_5112,N_8585);
nor UO_1284 (O_1284,N_7207,N_8203);
nand UO_1285 (O_1285,N_5949,N_7221);
nand UO_1286 (O_1286,N_7552,N_5701);
and UO_1287 (O_1287,N_8059,N_7655);
nor UO_1288 (O_1288,N_5522,N_8672);
or UO_1289 (O_1289,N_5241,N_5439);
nor UO_1290 (O_1290,N_7585,N_6785);
nand UO_1291 (O_1291,N_8920,N_6118);
nor UO_1292 (O_1292,N_8976,N_8036);
and UO_1293 (O_1293,N_7224,N_7074);
xor UO_1294 (O_1294,N_7479,N_7575);
or UO_1295 (O_1295,N_7370,N_9064);
or UO_1296 (O_1296,N_8531,N_9866);
and UO_1297 (O_1297,N_5426,N_6047);
and UO_1298 (O_1298,N_7667,N_5004);
or UO_1299 (O_1299,N_9095,N_7070);
nand UO_1300 (O_1300,N_6606,N_6889);
nor UO_1301 (O_1301,N_7939,N_5422);
nand UO_1302 (O_1302,N_5324,N_5886);
nand UO_1303 (O_1303,N_6353,N_9801);
and UO_1304 (O_1304,N_6430,N_8721);
nand UO_1305 (O_1305,N_6282,N_5178);
and UO_1306 (O_1306,N_5966,N_8134);
nor UO_1307 (O_1307,N_6802,N_6024);
nand UO_1308 (O_1308,N_7498,N_7325);
or UO_1309 (O_1309,N_8809,N_8685);
nand UO_1310 (O_1310,N_9264,N_8212);
nor UO_1311 (O_1311,N_6462,N_7929);
or UO_1312 (O_1312,N_5561,N_5427);
and UO_1313 (O_1313,N_5920,N_7589);
nand UO_1314 (O_1314,N_7809,N_6597);
or UO_1315 (O_1315,N_5343,N_9525);
nor UO_1316 (O_1316,N_5329,N_7883);
and UO_1317 (O_1317,N_5912,N_5992);
nand UO_1318 (O_1318,N_8636,N_5098);
nand UO_1319 (O_1319,N_5406,N_7038);
and UO_1320 (O_1320,N_6072,N_8807);
nor UO_1321 (O_1321,N_9202,N_5466);
and UO_1322 (O_1322,N_7827,N_7300);
nor UO_1323 (O_1323,N_5921,N_7362);
nand UO_1324 (O_1324,N_8844,N_7520);
and UO_1325 (O_1325,N_8350,N_8898);
nand UO_1326 (O_1326,N_5978,N_7829);
and UO_1327 (O_1327,N_8518,N_5182);
nand UO_1328 (O_1328,N_9615,N_9313);
or UO_1329 (O_1329,N_9203,N_9000);
and UO_1330 (O_1330,N_6801,N_7022);
and UO_1331 (O_1331,N_9904,N_7583);
and UO_1332 (O_1332,N_5649,N_7112);
nor UO_1333 (O_1333,N_6629,N_8527);
and UO_1334 (O_1334,N_9491,N_7919);
nor UO_1335 (O_1335,N_9085,N_7437);
and UO_1336 (O_1336,N_9509,N_8860);
and UO_1337 (O_1337,N_5395,N_7169);
and UO_1338 (O_1338,N_7268,N_6466);
nor UO_1339 (O_1339,N_6609,N_6503);
or UO_1340 (O_1340,N_6090,N_7191);
and UO_1341 (O_1341,N_5075,N_7509);
nand UO_1342 (O_1342,N_6206,N_8640);
nor UO_1343 (O_1343,N_8850,N_8108);
or UO_1344 (O_1344,N_5177,N_7839);
nand UO_1345 (O_1345,N_6844,N_8234);
xor UO_1346 (O_1346,N_7158,N_6792);
xnor UO_1347 (O_1347,N_8642,N_8095);
or UO_1348 (O_1348,N_7020,N_5393);
nor UO_1349 (O_1349,N_9570,N_9150);
and UO_1350 (O_1350,N_6169,N_9259);
nor UO_1351 (O_1351,N_5396,N_5160);
xnor UO_1352 (O_1352,N_5769,N_8257);
nand UO_1353 (O_1353,N_6833,N_9488);
or UO_1354 (O_1354,N_6098,N_7187);
or UO_1355 (O_1355,N_7307,N_6943);
and UO_1356 (O_1356,N_5052,N_5798);
nor UO_1357 (O_1357,N_8449,N_6547);
nor UO_1358 (O_1358,N_7911,N_8221);
and UO_1359 (O_1359,N_7668,N_9205);
or UO_1360 (O_1360,N_6819,N_6818);
nor UO_1361 (O_1361,N_9893,N_8691);
xor UO_1362 (O_1362,N_8651,N_9283);
or UO_1363 (O_1363,N_7654,N_8129);
nor UO_1364 (O_1364,N_5694,N_8741);
nand UO_1365 (O_1365,N_5205,N_8421);
nor UO_1366 (O_1366,N_9793,N_9161);
nor UO_1367 (O_1367,N_7674,N_8280);
nor UO_1368 (O_1368,N_6350,N_7031);
nand UO_1369 (O_1369,N_8173,N_8340);
and UO_1370 (O_1370,N_6385,N_5528);
nand UO_1371 (O_1371,N_7438,N_6227);
nand UO_1372 (O_1372,N_6784,N_8737);
nor UO_1373 (O_1373,N_5652,N_8605);
nand UO_1374 (O_1374,N_5963,N_7991);
and UO_1375 (O_1375,N_9605,N_5327);
or UO_1376 (O_1376,N_6179,N_9059);
or UO_1377 (O_1377,N_5527,N_5306);
and UO_1378 (O_1378,N_9494,N_6932);
nor UO_1379 (O_1379,N_5927,N_8397);
and UO_1380 (O_1380,N_9065,N_8593);
nand UO_1381 (O_1381,N_6107,N_8171);
and UO_1382 (O_1382,N_5538,N_5867);
nor UO_1383 (O_1383,N_5826,N_6101);
nor UO_1384 (O_1384,N_7176,N_5392);
nor UO_1385 (O_1385,N_6586,N_8921);
and UO_1386 (O_1386,N_8479,N_7422);
xnor UO_1387 (O_1387,N_8137,N_8067);
or UO_1388 (O_1388,N_6448,N_6315);
nor UO_1389 (O_1389,N_5797,N_5222);
nor UO_1390 (O_1390,N_9068,N_8101);
nand UO_1391 (O_1391,N_6419,N_7936);
or UO_1392 (O_1392,N_9584,N_6346);
nor UO_1393 (O_1393,N_7625,N_9116);
nand UO_1394 (O_1394,N_5731,N_7290);
nand UO_1395 (O_1395,N_5366,N_8007);
nor UO_1396 (O_1396,N_6632,N_9261);
nor UO_1397 (O_1397,N_5091,N_6793);
and UO_1398 (O_1398,N_7704,N_5262);
and UO_1399 (O_1399,N_7572,N_9775);
nor UO_1400 (O_1400,N_5332,N_7171);
nor UO_1401 (O_1401,N_8235,N_7997);
or UO_1402 (O_1402,N_9976,N_5201);
or UO_1403 (O_1403,N_6202,N_7515);
and UO_1404 (O_1404,N_8299,N_8297);
or UO_1405 (O_1405,N_7832,N_6018);
or UO_1406 (O_1406,N_5270,N_7716);
nand UO_1407 (O_1407,N_9536,N_9038);
nor UO_1408 (O_1408,N_5090,N_8897);
nor UO_1409 (O_1409,N_9206,N_5846);
nor UO_1410 (O_1410,N_6970,N_6059);
nand UO_1411 (O_1411,N_8488,N_5485);
nor UO_1412 (O_1412,N_5411,N_8609);
nand UO_1413 (O_1413,N_6414,N_9977);
nand UO_1414 (O_1414,N_8924,N_5568);
nand UO_1415 (O_1415,N_7518,N_8145);
or UO_1416 (O_1416,N_9226,N_9618);
and UO_1417 (O_1417,N_5780,N_9497);
nor UO_1418 (O_1418,N_9575,N_9772);
and UO_1419 (O_1419,N_8502,N_9037);
and UO_1420 (O_1420,N_7442,N_7050);
nand UO_1421 (O_1421,N_7083,N_9595);
and UO_1422 (O_1422,N_8613,N_5625);
nor UO_1423 (O_1423,N_7272,N_8482);
nor UO_1424 (O_1424,N_7761,N_9718);
nor UO_1425 (O_1425,N_9794,N_5218);
nor UO_1426 (O_1426,N_9406,N_7177);
or UO_1427 (O_1427,N_7740,N_6012);
and UO_1428 (O_1428,N_9614,N_9585);
and UO_1429 (O_1429,N_8648,N_5895);
nand UO_1430 (O_1430,N_9771,N_8098);
nand UO_1431 (O_1431,N_8551,N_6220);
and UO_1432 (O_1432,N_7734,N_5621);
or UO_1433 (O_1433,N_8682,N_9951);
and UO_1434 (O_1434,N_7684,N_5399);
and UO_1435 (O_1435,N_5476,N_8564);
or UO_1436 (O_1436,N_7100,N_8773);
nand UO_1437 (O_1437,N_5634,N_7049);
and UO_1438 (O_1438,N_6770,N_5263);
and UO_1439 (O_1439,N_6545,N_7336);
nor UO_1440 (O_1440,N_7195,N_6495);
nor UO_1441 (O_1441,N_5626,N_7423);
nand UO_1442 (O_1442,N_7291,N_9713);
nand UO_1443 (O_1443,N_5441,N_9325);
nor UO_1444 (O_1444,N_9677,N_8703);
and UO_1445 (O_1445,N_9230,N_9950);
and UO_1446 (O_1446,N_9513,N_7870);
nand UO_1447 (O_1447,N_6580,N_6319);
or UO_1448 (O_1448,N_5773,N_7706);
and UO_1449 (O_1449,N_7766,N_8718);
nor UO_1450 (O_1450,N_5868,N_6363);
nand UO_1451 (O_1451,N_9805,N_6417);
nor UO_1452 (O_1452,N_7971,N_9433);
and UO_1453 (O_1453,N_9376,N_6799);
nor UO_1454 (O_1454,N_6317,N_8361);
or UO_1455 (O_1455,N_5281,N_5315);
or UO_1456 (O_1456,N_5842,N_9271);
and UO_1457 (O_1457,N_6867,N_7738);
or UO_1458 (O_1458,N_5431,N_9142);
nor UO_1459 (O_1459,N_7807,N_8199);
nor UO_1460 (O_1460,N_6846,N_7804);
or UO_1461 (O_1461,N_7739,N_8357);
nor UO_1462 (O_1462,N_9005,N_9827);
nor UO_1463 (O_1463,N_9311,N_9883);
or UO_1464 (O_1464,N_7283,N_6897);
nor UO_1465 (O_1465,N_5120,N_7762);
and UO_1466 (O_1466,N_7198,N_8881);
and UO_1467 (O_1467,N_5487,N_5956);
nand UO_1468 (O_1468,N_6039,N_8700);
or UO_1469 (O_1469,N_6611,N_6129);
or UO_1470 (O_1470,N_5889,N_8796);
xor UO_1471 (O_1471,N_8766,N_8197);
nand UO_1472 (O_1472,N_9331,N_5631);
nand UO_1473 (O_1473,N_9165,N_8122);
nor UO_1474 (O_1474,N_7902,N_8236);
nor UO_1475 (O_1475,N_8192,N_5067);
nand UO_1476 (O_1476,N_8434,N_7683);
or UO_1477 (O_1477,N_5054,N_8848);
and UO_1478 (O_1478,N_7303,N_8602);
nor UO_1479 (O_1479,N_6053,N_6439);
and UO_1480 (O_1480,N_6046,N_8380);
nor UO_1481 (O_1481,N_9690,N_9216);
nor UO_1482 (O_1482,N_8560,N_7688);
nor UO_1483 (O_1483,N_8478,N_5349);
nand UO_1484 (O_1484,N_9572,N_7447);
nand UO_1485 (O_1485,N_5994,N_9591);
nand UO_1486 (O_1486,N_6959,N_5651);
or UO_1487 (O_1487,N_9746,N_6843);
xnor UO_1488 (O_1488,N_6766,N_7510);
or UO_1489 (O_1489,N_6857,N_8169);
nand UO_1490 (O_1490,N_6185,N_9723);
or UO_1491 (O_1491,N_8618,N_9301);
or UO_1492 (O_1492,N_5499,N_9273);
nand UO_1493 (O_1493,N_6771,N_5203);
xor UO_1494 (O_1494,N_5494,N_7537);
and UO_1495 (O_1495,N_8913,N_6807);
nor UO_1496 (O_1496,N_5539,N_9454);
nor UO_1497 (O_1497,N_6125,N_6377);
and UO_1498 (O_1498,N_5033,N_5299);
nand UO_1499 (O_1499,N_8675,N_6648);
endmodule