module basic_750_5000_1000_25_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_266,In_615);
nor U1 (N_1,In_169,In_619);
nand U2 (N_2,In_692,In_141);
or U3 (N_3,In_666,In_437);
and U4 (N_4,In_200,In_560);
nor U5 (N_5,In_360,In_729);
nor U6 (N_6,In_458,In_353);
or U7 (N_7,In_580,In_261);
and U8 (N_8,In_478,In_318);
and U9 (N_9,In_155,In_139);
or U10 (N_10,In_383,In_613);
and U11 (N_11,In_628,In_441);
or U12 (N_12,In_146,In_40);
xnor U13 (N_13,In_133,In_173);
xnor U14 (N_14,In_26,In_711);
and U15 (N_15,In_625,In_23);
and U16 (N_16,In_269,In_45);
xor U17 (N_17,In_514,In_305);
and U18 (N_18,In_22,In_278);
and U19 (N_19,In_587,In_591);
and U20 (N_20,In_4,In_290);
nor U21 (N_21,In_41,In_681);
or U22 (N_22,In_714,In_398);
nor U23 (N_23,In_12,In_355);
nand U24 (N_24,In_338,In_109);
nand U25 (N_25,In_612,In_724);
nor U26 (N_26,In_2,In_137);
or U27 (N_27,In_391,In_396);
nor U28 (N_28,In_542,In_361);
nand U29 (N_29,In_245,In_6);
nor U30 (N_30,In_250,In_302);
nand U31 (N_31,In_224,In_185);
nand U32 (N_32,In_199,In_241);
and U33 (N_33,In_470,In_674);
nand U34 (N_34,In_140,In_521);
or U35 (N_35,In_256,In_747);
nor U36 (N_36,In_10,In_722);
or U37 (N_37,In_659,In_616);
or U38 (N_38,In_610,In_225);
nand U39 (N_39,In_392,In_21);
or U40 (N_40,In_648,In_663);
or U41 (N_41,In_452,In_161);
nor U42 (N_42,In_322,In_236);
nand U43 (N_43,In_601,In_198);
nor U44 (N_44,In_201,In_60);
and U45 (N_45,In_152,In_216);
xnor U46 (N_46,In_286,In_43);
xor U47 (N_47,In_545,In_637);
nand U48 (N_48,In_49,In_550);
nand U49 (N_49,In_158,In_489);
or U50 (N_50,In_260,In_394);
nand U51 (N_51,In_519,In_429);
nor U52 (N_52,In_484,In_691);
nor U53 (N_53,In_264,In_268);
nor U54 (N_54,In_682,In_237);
xnor U55 (N_55,In_157,In_459);
nand U56 (N_56,In_189,In_535);
and U57 (N_57,In_678,In_719);
nor U58 (N_58,In_455,In_186);
nor U59 (N_59,In_377,In_288);
nand U60 (N_60,In_639,In_276);
xnor U61 (N_61,In_39,In_407);
xor U62 (N_62,In_346,In_16);
or U63 (N_63,In_246,In_243);
nor U64 (N_64,In_138,In_488);
nor U65 (N_65,In_147,In_235);
and U66 (N_66,In_124,In_79);
nand U67 (N_67,In_569,In_480);
nor U68 (N_68,In_351,In_425);
nor U69 (N_69,In_727,In_638);
nand U70 (N_70,In_510,In_700);
nor U71 (N_71,In_176,In_544);
nand U72 (N_72,In_702,In_378);
or U73 (N_73,In_512,In_645);
or U74 (N_74,In_136,In_617);
nor U75 (N_75,In_403,In_369);
and U76 (N_76,In_98,In_597);
xnor U77 (N_77,In_18,In_270);
or U78 (N_78,In_144,In_151);
or U79 (N_79,In_603,In_502);
or U80 (N_80,In_609,In_233);
xor U81 (N_81,In_15,In_431);
xor U82 (N_82,In_527,In_29);
or U83 (N_83,In_611,In_704);
or U84 (N_84,In_149,In_238);
or U85 (N_85,In_731,In_668);
or U86 (N_86,In_585,In_63);
or U87 (N_87,In_640,In_449);
xor U88 (N_88,In_337,In_568);
nand U89 (N_89,In_249,In_232);
xor U90 (N_90,In_127,In_24);
nor U91 (N_91,In_490,In_194);
nor U92 (N_92,In_107,In_366);
xnor U93 (N_93,In_183,In_165);
or U94 (N_94,In_234,In_385);
and U95 (N_95,In_633,In_5);
nand U96 (N_96,In_556,In_229);
nand U97 (N_97,In_306,In_148);
nor U98 (N_98,In_523,In_104);
and U99 (N_99,In_81,In_82);
and U100 (N_100,In_536,In_742);
and U101 (N_101,In_606,In_273);
nor U102 (N_102,In_287,In_664);
xor U103 (N_103,In_558,In_421);
nor U104 (N_104,In_390,In_142);
or U105 (N_105,In_740,In_240);
nor U106 (N_106,In_406,In_472);
xnor U107 (N_107,In_461,In_543);
nor U108 (N_108,In_53,In_333);
nor U109 (N_109,In_426,In_358);
and U110 (N_110,In_415,In_516);
and U111 (N_111,In_631,In_145);
nor U112 (N_112,In_710,In_414);
nor U113 (N_113,In_258,In_319);
and U114 (N_114,In_654,In_172);
and U115 (N_115,In_177,In_596);
or U116 (N_116,In_715,In_65);
and U117 (N_117,In_326,In_373);
and U118 (N_118,In_283,In_301);
nand U119 (N_119,In_693,In_584);
and U120 (N_120,In_365,In_683);
nand U121 (N_121,In_744,In_47);
and U122 (N_122,In_528,In_393);
and U123 (N_123,In_670,In_552);
or U124 (N_124,In_422,In_450);
nor U125 (N_125,In_713,In_299);
nand U126 (N_126,In_749,In_275);
or U127 (N_127,In_336,In_563);
and U128 (N_128,In_745,In_447);
nor U129 (N_129,In_531,In_518);
and U130 (N_130,In_561,In_120);
nand U131 (N_131,In_471,In_718);
nand U132 (N_132,In_341,In_402);
nand U133 (N_133,In_62,In_94);
or U134 (N_134,In_347,In_254);
or U135 (N_135,In_297,In_119);
nand U136 (N_136,In_323,In_72);
or U137 (N_137,In_190,In_181);
nand U138 (N_138,In_537,In_741);
or U139 (N_139,In_85,In_187);
nand U140 (N_140,In_36,In_624);
and U141 (N_141,In_382,In_32);
or U142 (N_142,In_20,In_413);
nand U143 (N_143,In_367,In_313);
nand U144 (N_144,In_70,In_52);
nor U145 (N_145,In_272,In_122);
nor U146 (N_146,In_226,In_412);
and U147 (N_147,In_457,In_105);
or U148 (N_148,In_474,In_706);
or U149 (N_149,In_325,In_445);
nand U150 (N_150,In_384,In_463);
and U151 (N_151,In_281,In_202);
nor U152 (N_152,In_661,In_466);
nor U153 (N_153,In_493,In_332);
nand U154 (N_154,In_168,In_33);
nor U155 (N_155,In_419,In_737);
nand U156 (N_156,In_634,In_228);
nand U157 (N_157,In_476,In_3);
nor U158 (N_158,In_126,In_635);
nor U159 (N_159,In_357,In_331);
or U160 (N_160,In_191,In_453);
or U161 (N_161,In_643,In_443);
nor U162 (N_162,In_223,In_477);
nand U163 (N_163,In_428,In_75);
and U164 (N_164,In_685,In_559);
or U165 (N_165,In_698,In_629);
nor U166 (N_166,In_581,In_651);
xnor U167 (N_167,In_91,In_28);
nor U168 (N_168,In_34,In_354);
nor U169 (N_169,In_248,In_78);
nor U170 (N_170,In_77,In_195);
and U171 (N_171,In_300,In_511);
nand U172 (N_172,In_469,In_686);
nand U173 (N_173,In_71,In_178);
nor U174 (N_174,In_370,In_374);
nand U175 (N_175,In_99,In_9);
nand U176 (N_176,In_646,In_388);
xnor U177 (N_177,In_503,In_513);
or U178 (N_178,In_219,In_196);
or U179 (N_179,In_676,In_58);
and U180 (N_180,In_604,In_123);
or U181 (N_181,In_7,In_436);
nand U182 (N_182,In_732,In_557);
and U183 (N_183,In_193,In_541);
nand U184 (N_184,In_409,In_626);
or U185 (N_185,In_296,In_592);
nor U186 (N_186,In_117,In_66);
xor U187 (N_187,In_709,In_498);
and U188 (N_188,In_594,In_106);
nor U189 (N_189,In_595,In_314);
nor U190 (N_190,In_285,In_92);
xnor U191 (N_191,In_19,In_289);
nand U192 (N_192,In_174,In_166);
xnor U193 (N_193,In_221,In_100);
nand U194 (N_194,In_340,In_408);
nor U195 (N_195,In_239,In_184);
nand U196 (N_196,In_534,In_0);
xor U197 (N_197,In_156,In_725);
or U198 (N_198,In_231,In_339);
and U199 (N_199,In_74,In_1);
or U200 (N_200,In_227,In_620);
and U201 (N_201,In_214,In_131);
nor U202 (N_202,In_647,N_127);
nand U203 (N_203,N_168,In_451);
and U204 (N_204,In_208,In_68);
or U205 (N_205,N_144,In_547);
nand U206 (N_206,N_170,In_102);
nand U207 (N_207,In_282,In_562);
and U208 (N_208,In_649,In_121);
nor U209 (N_209,N_107,In_101);
nand U210 (N_210,In_416,In_736);
nand U211 (N_211,In_204,N_77);
or U212 (N_212,In_197,N_37);
and U213 (N_213,N_63,In_263);
or U214 (N_214,N_150,In_672);
or U215 (N_215,In_87,In_621);
nand U216 (N_216,N_198,N_35);
nor U217 (N_217,In_315,N_49);
xor U218 (N_218,In_575,N_101);
nor U219 (N_219,In_247,In_485);
or U220 (N_220,N_45,N_94);
nor U221 (N_221,In_362,In_673);
or U222 (N_222,N_38,In_192);
and U223 (N_223,N_100,In_252);
or U224 (N_224,In_748,In_170);
or U225 (N_225,In_669,In_423);
nand U226 (N_226,In_627,In_548);
and U227 (N_227,In_303,N_120);
xor U228 (N_228,N_90,N_56);
and U229 (N_229,N_183,N_27);
or U230 (N_230,In_712,In_150);
xnor U231 (N_231,In_690,In_11);
nand U232 (N_232,In_522,N_187);
nor U233 (N_233,In_397,N_123);
nor U234 (N_234,In_310,In_658);
nand U235 (N_235,In_586,In_293);
and U236 (N_236,In_515,In_345);
or U237 (N_237,In_335,In_159);
and U238 (N_238,In_707,N_137);
or U239 (N_239,In_456,N_160);
nor U240 (N_240,In_97,N_171);
xnor U241 (N_241,In_342,In_524);
nand U242 (N_242,In_589,In_371);
nor U243 (N_243,In_465,In_687);
nor U244 (N_244,In_162,N_33);
nand U245 (N_245,N_40,In_464);
or U246 (N_246,In_506,N_46);
xor U247 (N_247,In_577,In_520);
xnor U248 (N_248,N_10,N_4);
nor U249 (N_249,In_188,In_317);
xor U250 (N_250,In_481,N_71);
nand U251 (N_251,In_130,In_701);
nand U252 (N_252,In_372,N_164);
nor U253 (N_253,In_641,In_111);
xnor U254 (N_254,N_85,In_538);
and U255 (N_255,N_116,In_128);
nand U256 (N_256,In_205,In_381);
and U257 (N_257,In_573,In_572);
xnor U258 (N_258,In_86,In_433);
nor U259 (N_259,N_53,In_467);
and U260 (N_260,In_438,In_344);
nand U261 (N_261,In_51,In_73);
or U262 (N_262,N_65,N_88);
nor U263 (N_263,N_131,In_675);
nor U264 (N_264,In_37,N_51);
and U265 (N_265,In_376,In_588);
and U266 (N_266,N_50,N_43);
nand U267 (N_267,In_486,N_162);
nor U268 (N_268,In_180,In_48);
nand U269 (N_269,In_14,In_89);
nor U270 (N_270,In_375,In_112);
nand U271 (N_271,N_7,N_108);
and U272 (N_272,In_636,In_17);
nor U273 (N_273,N_32,N_130);
nand U274 (N_274,N_145,N_109);
and U275 (N_275,N_189,In_316);
nand U276 (N_276,N_80,In_386);
and U277 (N_277,In_38,N_99);
and U278 (N_278,In_509,In_671);
xnor U279 (N_279,In_656,In_230);
or U280 (N_280,N_6,In_571);
nand U281 (N_281,N_58,In_46);
nor U282 (N_282,In_652,N_193);
nand U283 (N_283,In_504,N_61);
nand U284 (N_284,In_598,N_12);
xor U285 (N_285,N_185,In_363);
or U286 (N_286,In_460,N_176);
or U287 (N_287,In_80,N_184);
nor U288 (N_288,N_103,In_76);
nand U289 (N_289,In_582,In_153);
nor U290 (N_290,In_726,N_140);
nor U291 (N_291,N_70,In_309);
nor U292 (N_292,N_196,N_158);
nand U293 (N_293,In_350,In_321);
or U294 (N_294,In_44,In_88);
nor U295 (N_295,N_175,In_209);
and U296 (N_296,In_526,N_17);
nand U297 (N_297,In_220,N_15);
or U298 (N_298,In_242,In_507);
and U299 (N_299,In_689,In_262);
xor U300 (N_300,In_175,N_96);
or U301 (N_301,In_280,In_623);
xor U302 (N_302,N_169,In_90);
or U303 (N_303,In_8,In_271);
and U304 (N_304,In_539,In_277);
nand U305 (N_305,In_607,N_178);
or U306 (N_306,In_655,In_405);
or U307 (N_307,In_696,In_650);
nand U308 (N_308,In_55,In_448);
xor U309 (N_309,In_442,N_20);
and U310 (N_310,In_61,In_677);
nor U311 (N_311,N_98,In_118);
nor U312 (N_312,N_48,N_156);
and U313 (N_313,In_135,N_54);
or U314 (N_314,In_600,In_328);
or U315 (N_315,N_92,In_108);
and U316 (N_316,In_129,In_67);
and U317 (N_317,N_36,N_139);
and U318 (N_318,N_129,In_475);
nor U319 (N_319,In_103,In_329);
nor U320 (N_320,In_349,In_434);
nor U321 (N_321,In_251,N_11);
nor U322 (N_322,In_739,In_379);
nor U323 (N_323,N_114,In_213);
or U324 (N_324,In_716,In_717);
and U325 (N_325,In_13,N_2);
nand U326 (N_326,In_125,In_253);
and U327 (N_327,In_487,N_93);
or U328 (N_328,In_501,N_55);
or U329 (N_329,N_74,In_171);
nor U330 (N_330,In_279,In_222);
nor U331 (N_331,N_16,N_133);
or U332 (N_332,In_267,In_56);
xor U333 (N_333,In_27,In_114);
and U334 (N_334,N_186,N_181);
nor U335 (N_335,In_25,In_163);
nand U336 (N_336,In_680,In_667);
nand U337 (N_337,N_141,In_435);
nor U338 (N_338,In_294,In_565);
nand U339 (N_339,In_244,In_399);
xnor U340 (N_340,In_420,In_593);
and U341 (N_341,N_122,In_430);
nor U342 (N_342,N_1,N_89);
nor U343 (N_343,N_146,In_496);
or U344 (N_344,N_13,N_167);
and U345 (N_345,N_153,N_149);
xor U346 (N_346,In_320,N_112);
nor U347 (N_347,N_102,In_298);
nand U348 (N_348,In_179,In_327);
or U349 (N_349,In_738,N_179);
and U350 (N_350,In_630,In_644);
nor U351 (N_351,In_662,In_614);
nand U352 (N_352,In_695,N_174);
and U353 (N_353,N_194,In_479);
and U354 (N_354,In_312,In_602);
nand U355 (N_355,N_125,In_497);
and U356 (N_356,N_23,N_44);
or U357 (N_357,In_215,In_330);
nor U358 (N_358,In_93,In_400);
or U359 (N_359,N_81,In_533);
nand U360 (N_360,In_579,In_84);
or U361 (N_361,In_440,In_307);
nand U362 (N_362,N_57,N_104);
or U363 (N_363,N_21,N_154);
or U364 (N_364,In_110,N_161);
or U365 (N_365,In_30,N_195);
or U366 (N_366,In_64,In_508);
nor U367 (N_367,N_39,In_31);
and U368 (N_368,In_554,N_182);
nand U369 (N_369,In_427,N_73);
or U370 (N_370,In_368,N_110);
nand U371 (N_371,In_622,N_132);
nor U372 (N_372,In_35,In_705);
and U373 (N_373,N_47,In_274);
nor U374 (N_374,In_608,In_308);
nor U375 (N_375,In_182,In_499);
nand U376 (N_376,In_599,N_165);
and U377 (N_377,N_177,N_59);
and U378 (N_378,In_632,In_549);
nand U379 (N_379,In_653,In_500);
nand U380 (N_380,N_124,In_570);
xor U381 (N_381,N_79,N_113);
xnor U382 (N_382,N_69,In_54);
and U383 (N_383,In_83,In_660);
and U384 (N_384,N_91,In_255);
nor U385 (N_385,N_0,In_57);
or U386 (N_386,In_743,N_148);
and U387 (N_387,In_207,N_64);
xnor U388 (N_388,N_87,N_83);
and U389 (N_389,N_42,In_95);
nor U390 (N_390,In_404,N_126);
and U391 (N_391,In_311,In_567);
xor U392 (N_392,In_42,N_119);
and U393 (N_393,In_432,N_111);
or U394 (N_394,In_540,N_115);
and U395 (N_395,N_190,N_24);
nand U396 (N_396,In_699,In_352);
nor U397 (N_397,In_694,In_387);
and U398 (N_398,In_578,N_199);
or U399 (N_399,N_41,In_164);
or U400 (N_400,N_223,N_246);
nand U401 (N_401,N_337,N_373);
and U402 (N_402,N_272,In_295);
xnor U403 (N_403,N_235,N_52);
or U404 (N_404,In_334,In_218);
or U405 (N_405,N_339,In_417);
or U406 (N_406,N_368,N_215);
nand U407 (N_407,N_34,N_117);
nor U408 (N_408,In_439,N_324);
and U409 (N_409,N_371,In_59);
nor U410 (N_410,N_212,N_218);
or U411 (N_411,N_298,N_352);
and U412 (N_412,N_281,N_67);
nor U413 (N_413,N_227,N_313);
nand U414 (N_414,N_391,In_495);
and U415 (N_415,N_277,In_576);
and U416 (N_416,N_206,N_247);
nor U417 (N_417,N_306,N_345);
nor U418 (N_418,In_730,N_192);
nand U419 (N_419,In_734,In_134);
nor U420 (N_420,N_76,N_5);
nand U421 (N_421,In_483,In_721);
or U422 (N_422,N_335,In_454);
or U423 (N_423,N_321,In_217);
nor U424 (N_424,In_566,N_322);
or U425 (N_425,N_211,N_163);
nand U426 (N_426,N_279,In_116);
or U427 (N_427,In_733,N_332);
nor U428 (N_428,N_263,N_383);
or U429 (N_429,In_50,N_260);
nand U430 (N_430,N_268,In_343);
or U431 (N_431,N_251,N_294);
nor U432 (N_432,N_173,N_22);
or U433 (N_433,In_530,N_286);
xnor U434 (N_434,N_265,N_261);
and U435 (N_435,N_387,N_293);
nor U436 (N_436,N_304,In_553);
nor U437 (N_437,N_14,N_318);
xnor U438 (N_438,In_348,N_393);
or U439 (N_439,N_280,N_209);
nor U440 (N_440,N_62,N_244);
nor U441 (N_441,N_312,N_26);
nor U442 (N_442,N_346,In_720);
and U443 (N_443,N_202,In_679);
or U444 (N_444,In_132,N_365);
nand U445 (N_445,N_292,N_9);
or U446 (N_446,N_309,N_317);
xor U447 (N_447,In_665,In_688);
xnor U448 (N_448,N_299,N_361);
and U449 (N_449,N_331,N_232);
nor U450 (N_450,N_325,N_97);
nor U451 (N_451,N_273,N_390);
xnor U452 (N_452,N_297,N_264);
nand U453 (N_453,In_517,N_296);
nand U454 (N_454,N_301,N_236);
and U455 (N_455,N_283,N_311);
nand U456 (N_456,N_230,N_367);
or U457 (N_457,N_363,N_398);
or U458 (N_458,N_348,In_115);
nor U459 (N_459,In_257,N_172);
nor U460 (N_460,N_316,N_267);
and U461 (N_461,In_462,N_289);
nor U462 (N_462,In_424,N_319);
nor U463 (N_463,N_381,In_657);
and U464 (N_464,N_303,N_31);
or U465 (N_465,N_191,In_491);
nand U466 (N_466,In_359,In_605);
nand U467 (N_467,N_106,In_684);
nand U468 (N_468,N_166,N_315);
or U469 (N_469,N_291,N_254);
or U470 (N_470,N_344,N_343);
nor U471 (N_471,N_210,N_341);
or U472 (N_472,In_590,N_152);
or U473 (N_473,N_266,In_505);
and U474 (N_474,N_307,N_147);
and U475 (N_475,N_395,N_330);
and U476 (N_476,In_735,N_397);
or U477 (N_477,N_159,N_334);
or U478 (N_478,N_328,N_382);
xnor U479 (N_479,N_396,N_19);
nor U480 (N_480,N_60,In_259);
nor U481 (N_481,In_492,N_220);
or U482 (N_482,N_394,N_225);
nor U483 (N_483,In_468,N_228);
nor U484 (N_484,In_574,N_369);
and U485 (N_485,N_357,N_278);
or U486 (N_486,N_242,N_270);
and U487 (N_487,N_78,N_327);
and U488 (N_488,N_349,N_3);
nand U489 (N_489,N_82,In_206);
or U490 (N_490,N_233,N_284);
nand U491 (N_491,N_329,In_697);
nand U492 (N_492,N_213,N_384);
or U493 (N_493,In_703,N_326);
nand U494 (N_494,N_290,N_214);
nand U495 (N_495,N_259,N_30);
nor U496 (N_496,N_95,N_392);
nand U497 (N_497,N_68,N_208);
nand U498 (N_498,N_305,N_276);
or U499 (N_499,In_212,N_205);
or U500 (N_500,N_310,N_342);
or U501 (N_501,In_265,In_746);
and U502 (N_502,N_155,N_243);
xnor U503 (N_503,In_203,N_300);
nor U504 (N_504,N_372,N_29);
and U505 (N_505,N_86,In_532);
nor U506 (N_506,N_360,N_386);
or U507 (N_507,N_200,N_229);
or U508 (N_508,In_154,N_375);
nand U509 (N_509,N_320,In_292);
nor U510 (N_510,In_389,N_203);
and U511 (N_511,In_555,N_380);
nor U512 (N_512,In_618,N_252);
or U513 (N_513,N_201,N_347);
xnor U514 (N_514,N_121,N_258);
nand U515 (N_515,N_8,N_142);
nand U516 (N_516,N_399,In_143);
nor U517 (N_517,N_388,In_446);
xor U518 (N_518,N_302,N_239);
xnor U519 (N_519,N_180,N_188);
nor U520 (N_520,N_354,N_245);
xor U521 (N_521,N_389,N_353);
nor U522 (N_522,In_113,In_210);
nor U523 (N_523,In_525,In_728);
or U524 (N_524,N_308,N_217);
nor U525 (N_525,N_350,In_380);
or U526 (N_526,In_167,In_708);
or U527 (N_527,N_75,N_359);
xnor U528 (N_528,In_494,N_237);
nand U529 (N_529,In_291,N_285);
nand U530 (N_530,N_385,N_287);
or U531 (N_531,In_564,N_157);
or U532 (N_532,N_271,N_25);
nand U533 (N_533,N_231,N_338);
nor U534 (N_534,N_376,N_379);
nor U535 (N_535,N_336,N_355);
nor U536 (N_536,N_378,N_84);
nand U537 (N_537,N_134,N_28);
xor U538 (N_538,N_118,N_224);
nand U539 (N_539,In_546,N_66);
and U540 (N_540,In_723,N_207);
or U541 (N_541,N_314,N_257);
xnor U542 (N_542,N_351,N_216);
nor U543 (N_543,N_204,N_374);
or U544 (N_544,N_333,N_282);
or U545 (N_545,In_364,N_221);
nor U546 (N_546,N_249,In_529);
or U547 (N_547,N_275,N_295);
nand U548 (N_548,N_143,N_105);
or U549 (N_549,In_411,N_356);
and U550 (N_550,In_160,N_135);
or U551 (N_551,N_138,N_197);
nor U552 (N_552,N_255,In_96);
and U553 (N_553,N_238,N_364);
xnor U554 (N_554,N_128,N_226);
or U555 (N_555,N_136,N_323);
or U556 (N_556,In_401,N_370);
nand U557 (N_557,In_473,N_240);
nor U558 (N_558,N_269,In_444);
or U559 (N_559,In_304,N_256);
nor U560 (N_560,N_250,N_222);
nand U561 (N_561,N_151,N_219);
and U562 (N_562,N_358,In_395);
nor U563 (N_563,N_366,N_274);
nand U564 (N_564,In_356,N_377);
and U565 (N_565,In_642,N_340);
and U566 (N_566,In_284,N_362);
xnor U567 (N_567,N_253,N_288);
nor U568 (N_568,In_69,In_583);
xor U569 (N_569,N_248,N_72);
and U570 (N_570,N_234,In_482);
nor U571 (N_571,In_410,N_241);
nand U572 (N_572,In_551,In_324);
or U573 (N_573,In_211,In_418);
nor U574 (N_574,N_262,N_18);
xnor U575 (N_575,N_230,In_292);
nor U576 (N_576,In_566,In_113);
xnor U577 (N_577,N_350,In_304);
and U578 (N_578,N_320,In_50);
nor U579 (N_579,N_29,N_371);
and U580 (N_580,N_166,N_142);
nor U581 (N_581,N_355,N_163);
and U582 (N_582,N_290,N_348);
xnor U583 (N_583,N_285,N_95);
nor U584 (N_584,In_684,In_132);
or U585 (N_585,N_398,In_473);
xor U586 (N_586,N_371,N_138);
xor U587 (N_587,N_271,N_377);
or U588 (N_588,In_495,N_385);
nor U589 (N_589,N_393,In_529);
nor U590 (N_590,In_292,N_347);
and U591 (N_591,In_96,N_351);
or U592 (N_592,N_152,In_720);
or U593 (N_593,N_308,N_134);
nand U594 (N_594,N_242,N_361);
nor U595 (N_595,N_14,In_553);
and U596 (N_596,N_266,N_296);
nand U597 (N_597,N_118,N_157);
or U598 (N_598,In_708,N_320);
nand U599 (N_599,In_132,N_256);
and U600 (N_600,N_463,N_557);
and U601 (N_601,N_477,N_435);
and U602 (N_602,N_407,N_531);
nor U603 (N_603,N_479,N_537);
nand U604 (N_604,N_588,N_598);
and U605 (N_605,N_418,N_578);
xor U606 (N_606,N_595,N_561);
and U607 (N_607,N_528,N_425);
or U608 (N_608,N_474,N_587);
or U609 (N_609,N_486,N_582);
and U610 (N_610,N_424,N_417);
or U611 (N_611,N_568,N_596);
and U612 (N_612,N_524,N_507);
or U613 (N_613,N_404,N_453);
nand U614 (N_614,N_481,N_408);
and U615 (N_615,N_471,N_452);
nand U616 (N_616,N_567,N_580);
or U617 (N_617,N_569,N_488);
or U618 (N_618,N_508,N_516);
and U619 (N_619,N_592,N_440);
and U620 (N_620,N_546,N_415);
xnor U621 (N_621,N_583,N_489);
nor U622 (N_622,N_503,N_437);
nor U623 (N_623,N_514,N_534);
or U624 (N_624,N_439,N_403);
or U625 (N_625,N_430,N_436);
nor U626 (N_626,N_540,N_594);
nand U627 (N_627,N_444,N_527);
nor U628 (N_628,N_491,N_443);
nand U629 (N_629,N_522,N_562);
or U630 (N_630,N_559,N_454);
and U631 (N_631,N_570,N_506);
nor U632 (N_632,N_574,N_542);
nor U633 (N_633,N_523,N_513);
or U634 (N_634,N_420,N_564);
or U635 (N_635,N_466,N_462);
nand U636 (N_636,N_448,N_402);
or U637 (N_637,N_460,N_585);
or U638 (N_638,N_400,N_593);
or U639 (N_639,N_543,N_427);
or U640 (N_640,N_549,N_539);
xor U641 (N_641,N_442,N_476);
nand U642 (N_642,N_597,N_554);
nand U643 (N_643,N_566,N_500);
or U644 (N_644,N_449,N_480);
nor U645 (N_645,N_412,N_532);
or U646 (N_646,N_461,N_494);
and U647 (N_647,N_552,N_538);
nand U648 (N_648,N_450,N_590);
and U649 (N_649,N_533,N_521);
and U650 (N_650,N_497,N_501);
and U651 (N_651,N_411,N_465);
or U652 (N_652,N_413,N_515);
nand U653 (N_653,N_493,N_558);
and U654 (N_654,N_550,N_426);
or U655 (N_655,N_423,N_529);
xnor U656 (N_656,N_599,N_421);
nor U657 (N_657,N_473,N_545);
and U658 (N_658,N_496,N_555);
or U659 (N_659,N_576,N_405);
nand U660 (N_660,N_441,N_518);
and U661 (N_661,N_575,N_556);
xnor U662 (N_662,N_504,N_560);
or U663 (N_663,N_483,N_485);
nand U664 (N_664,N_551,N_487);
xnor U665 (N_665,N_455,N_526);
nand U666 (N_666,N_525,N_548);
or U667 (N_667,N_456,N_475);
nor U668 (N_668,N_535,N_446);
nand U669 (N_669,N_472,N_478);
or U670 (N_670,N_457,N_505);
and U671 (N_671,N_429,N_519);
or U672 (N_672,N_541,N_410);
nor U673 (N_673,N_490,N_495);
xor U674 (N_674,N_484,N_572);
or U675 (N_675,N_433,N_553);
nor U676 (N_676,N_447,N_431);
or U677 (N_677,N_584,N_591);
nor U678 (N_678,N_502,N_536);
nand U679 (N_679,N_547,N_419);
and U680 (N_680,N_510,N_469);
nand U681 (N_681,N_432,N_482);
and U682 (N_682,N_434,N_544);
nand U683 (N_683,N_509,N_401);
or U684 (N_684,N_468,N_577);
and U685 (N_685,N_589,N_571);
nand U686 (N_686,N_406,N_464);
or U687 (N_687,N_422,N_445);
nand U688 (N_688,N_459,N_565);
nor U689 (N_689,N_470,N_416);
xor U690 (N_690,N_492,N_586);
and U691 (N_691,N_563,N_414);
and U692 (N_692,N_530,N_467);
nor U693 (N_693,N_499,N_579);
nand U694 (N_694,N_517,N_428);
nand U695 (N_695,N_511,N_498);
nand U696 (N_696,N_458,N_573);
nor U697 (N_697,N_581,N_438);
and U698 (N_698,N_520,N_451);
nor U699 (N_699,N_512,N_409);
nor U700 (N_700,N_532,N_585);
and U701 (N_701,N_491,N_427);
and U702 (N_702,N_413,N_463);
and U703 (N_703,N_535,N_439);
and U704 (N_704,N_588,N_465);
and U705 (N_705,N_533,N_542);
nor U706 (N_706,N_412,N_589);
nand U707 (N_707,N_413,N_416);
and U708 (N_708,N_588,N_450);
nand U709 (N_709,N_541,N_580);
or U710 (N_710,N_510,N_427);
and U711 (N_711,N_446,N_447);
xor U712 (N_712,N_593,N_517);
or U713 (N_713,N_566,N_552);
nor U714 (N_714,N_596,N_425);
nor U715 (N_715,N_568,N_465);
nand U716 (N_716,N_578,N_597);
nand U717 (N_717,N_437,N_581);
and U718 (N_718,N_446,N_596);
nor U719 (N_719,N_543,N_585);
and U720 (N_720,N_582,N_444);
or U721 (N_721,N_540,N_586);
nor U722 (N_722,N_551,N_552);
nor U723 (N_723,N_451,N_501);
nor U724 (N_724,N_400,N_459);
xnor U725 (N_725,N_536,N_426);
and U726 (N_726,N_540,N_451);
nor U727 (N_727,N_553,N_419);
and U728 (N_728,N_475,N_402);
or U729 (N_729,N_507,N_437);
and U730 (N_730,N_473,N_406);
or U731 (N_731,N_495,N_476);
nand U732 (N_732,N_403,N_584);
or U733 (N_733,N_546,N_471);
nor U734 (N_734,N_563,N_524);
nor U735 (N_735,N_523,N_550);
nand U736 (N_736,N_415,N_565);
and U737 (N_737,N_494,N_508);
and U738 (N_738,N_405,N_432);
and U739 (N_739,N_489,N_419);
nand U740 (N_740,N_441,N_403);
nand U741 (N_741,N_512,N_472);
or U742 (N_742,N_546,N_596);
nor U743 (N_743,N_559,N_537);
nand U744 (N_744,N_436,N_567);
nor U745 (N_745,N_483,N_435);
or U746 (N_746,N_559,N_530);
nor U747 (N_747,N_578,N_505);
nand U748 (N_748,N_537,N_451);
or U749 (N_749,N_544,N_454);
or U750 (N_750,N_450,N_562);
or U751 (N_751,N_423,N_447);
or U752 (N_752,N_537,N_507);
and U753 (N_753,N_479,N_520);
or U754 (N_754,N_423,N_474);
and U755 (N_755,N_489,N_523);
nor U756 (N_756,N_434,N_526);
nor U757 (N_757,N_420,N_458);
nor U758 (N_758,N_561,N_405);
xor U759 (N_759,N_567,N_560);
or U760 (N_760,N_415,N_419);
nand U761 (N_761,N_434,N_473);
or U762 (N_762,N_528,N_466);
nor U763 (N_763,N_510,N_497);
or U764 (N_764,N_515,N_551);
and U765 (N_765,N_557,N_427);
nand U766 (N_766,N_429,N_556);
nand U767 (N_767,N_420,N_566);
nor U768 (N_768,N_442,N_512);
nand U769 (N_769,N_402,N_512);
xor U770 (N_770,N_527,N_515);
xnor U771 (N_771,N_492,N_428);
nand U772 (N_772,N_477,N_595);
nand U773 (N_773,N_432,N_546);
and U774 (N_774,N_575,N_574);
nor U775 (N_775,N_472,N_528);
or U776 (N_776,N_573,N_596);
or U777 (N_777,N_506,N_586);
xor U778 (N_778,N_565,N_458);
and U779 (N_779,N_435,N_561);
and U780 (N_780,N_532,N_484);
nand U781 (N_781,N_434,N_480);
and U782 (N_782,N_444,N_544);
and U783 (N_783,N_496,N_543);
and U784 (N_784,N_541,N_469);
nor U785 (N_785,N_455,N_542);
nand U786 (N_786,N_444,N_455);
or U787 (N_787,N_473,N_554);
xor U788 (N_788,N_412,N_473);
nor U789 (N_789,N_481,N_507);
and U790 (N_790,N_466,N_542);
xor U791 (N_791,N_463,N_424);
nand U792 (N_792,N_562,N_581);
nor U793 (N_793,N_575,N_573);
nor U794 (N_794,N_470,N_570);
nor U795 (N_795,N_597,N_577);
or U796 (N_796,N_592,N_451);
or U797 (N_797,N_559,N_545);
nand U798 (N_798,N_479,N_462);
nand U799 (N_799,N_538,N_442);
nor U800 (N_800,N_717,N_611);
and U801 (N_801,N_613,N_691);
nor U802 (N_802,N_772,N_692);
or U803 (N_803,N_625,N_603);
nor U804 (N_804,N_715,N_762);
or U805 (N_805,N_724,N_657);
and U806 (N_806,N_765,N_616);
and U807 (N_807,N_670,N_734);
or U808 (N_808,N_700,N_770);
and U809 (N_809,N_761,N_759);
and U810 (N_810,N_784,N_658);
nand U811 (N_811,N_758,N_632);
or U812 (N_812,N_656,N_720);
nor U813 (N_813,N_614,N_681);
or U814 (N_814,N_620,N_755);
nand U815 (N_815,N_747,N_600);
or U816 (N_816,N_757,N_605);
and U817 (N_817,N_650,N_756);
and U818 (N_818,N_666,N_689);
or U819 (N_819,N_746,N_749);
xor U820 (N_820,N_708,N_766);
nor U821 (N_821,N_795,N_723);
nor U822 (N_822,N_667,N_793);
nand U823 (N_823,N_675,N_649);
nand U824 (N_824,N_682,N_783);
nor U825 (N_825,N_663,N_610);
xnor U826 (N_826,N_705,N_693);
nor U827 (N_827,N_760,N_641);
and U828 (N_828,N_647,N_773);
nor U829 (N_829,N_754,N_782);
and U830 (N_830,N_768,N_619);
nor U831 (N_831,N_753,N_771);
or U832 (N_832,N_609,N_653);
nor U833 (N_833,N_799,N_668);
and U834 (N_834,N_786,N_671);
or U835 (N_835,N_690,N_785);
nor U836 (N_836,N_792,N_726);
xor U837 (N_837,N_624,N_750);
and U838 (N_838,N_763,N_788);
or U839 (N_839,N_683,N_798);
or U840 (N_840,N_731,N_645);
or U841 (N_841,N_679,N_779);
and U842 (N_842,N_669,N_639);
nor U843 (N_843,N_677,N_767);
nor U844 (N_844,N_697,N_727);
nand U845 (N_845,N_626,N_643);
or U846 (N_846,N_703,N_661);
and U847 (N_847,N_642,N_737);
or U848 (N_848,N_710,N_686);
or U849 (N_849,N_797,N_751);
xnor U850 (N_850,N_638,N_790);
nand U851 (N_851,N_777,N_622);
nand U852 (N_852,N_796,N_730);
or U853 (N_853,N_601,N_718);
and U854 (N_854,N_712,N_711);
nand U855 (N_855,N_698,N_752);
xnor U856 (N_856,N_662,N_652);
nor U857 (N_857,N_633,N_764);
or U858 (N_858,N_728,N_604);
and U859 (N_859,N_744,N_635);
and U860 (N_860,N_655,N_615);
or U861 (N_861,N_636,N_660);
nand U862 (N_862,N_627,N_780);
nand U863 (N_863,N_787,N_602);
nand U864 (N_864,N_719,N_740);
or U865 (N_865,N_738,N_617);
and U866 (N_866,N_733,N_707);
or U867 (N_867,N_608,N_729);
or U868 (N_868,N_789,N_640);
nand U869 (N_869,N_741,N_646);
or U870 (N_870,N_776,N_629);
nand U871 (N_871,N_774,N_680);
nand U872 (N_872,N_775,N_612);
nor U873 (N_873,N_695,N_623);
and U874 (N_874,N_634,N_659);
nand U875 (N_875,N_654,N_676);
xor U876 (N_876,N_778,N_706);
and U877 (N_877,N_621,N_688);
nand U878 (N_878,N_713,N_685);
and U879 (N_879,N_637,N_769);
and U880 (N_880,N_699,N_648);
and U881 (N_881,N_748,N_716);
or U882 (N_882,N_702,N_791);
or U883 (N_883,N_665,N_725);
xnor U884 (N_884,N_696,N_644);
or U885 (N_885,N_739,N_736);
nand U886 (N_886,N_684,N_673);
and U887 (N_887,N_735,N_732);
nor U888 (N_888,N_672,N_722);
nor U889 (N_889,N_651,N_701);
and U890 (N_890,N_743,N_674);
nand U891 (N_891,N_721,N_687);
nand U892 (N_892,N_618,N_714);
nor U893 (N_893,N_709,N_607);
or U894 (N_894,N_630,N_704);
and U895 (N_895,N_694,N_781);
nand U896 (N_896,N_742,N_628);
or U897 (N_897,N_745,N_606);
nor U898 (N_898,N_664,N_678);
and U899 (N_899,N_631,N_794);
nand U900 (N_900,N_600,N_736);
xnor U901 (N_901,N_745,N_748);
nor U902 (N_902,N_760,N_739);
or U903 (N_903,N_659,N_755);
or U904 (N_904,N_696,N_658);
nor U905 (N_905,N_693,N_759);
and U906 (N_906,N_722,N_776);
nand U907 (N_907,N_798,N_672);
and U908 (N_908,N_650,N_620);
nand U909 (N_909,N_737,N_730);
and U910 (N_910,N_666,N_618);
nand U911 (N_911,N_774,N_626);
or U912 (N_912,N_689,N_761);
or U913 (N_913,N_796,N_656);
or U914 (N_914,N_742,N_699);
xor U915 (N_915,N_614,N_764);
or U916 (N_916,N_642,N_784);
nand U917 (N_917,N_673,N_730);
and U918 (N_918,N_772,N_671);
nor U919 (N_919,N_684,N_721);
or U920 (N_920,N_726,N_671);
xnor U921 (N_921,N_668,N_760);
nand U922 (N_922,N_681,N_639);
nand U923 (N_923,N_630,N_628);
and U924 (N_924,N_746,N_682);
or U925 (N_925,N_672,N_734);
or U926 (N_926,N_665,N_620);
and U927 (N_927,N_646,N_739);
or U928 (N_928,N_685,N_789);
and U929 (N_929,N_756,N_729);
nor U930 (N_930,N_638,N_644);
or U931 (N_931,N_764,N_615);
nor U932 (N_932,N_709,N_670);
nor U933 (N_933,N_621,N_765);
and U934 (N_934,N_751,N_772);
nor U935 (N_935,N_652,N_602);
or U936 (N_936,N_616,N_680);
nor U937 (N_937,N_672,N_688);
and U938 (N_938,N_754,N_762);
and U939 (N_939,N_726,N_665);
nand U940 (N_940,N_637,N_647);
and U941 (N_941,N_749,N_660);
or U942 (N_942,N_643,N_617);
nor U943 (N_943,N_623,N_735);
and U944 (N_944,N_726,N_629);
nand U945 (N_945,N_674,N_664);
nor U946 (N_946,N_733,N_706);
or U947 (N_947,N_606,N_669);
and U948 (N_948,N_653,N_758);
xnor U949 (N_949,N_683,N_786);
nand U950 (N_950,N_742,N_609);
or U951 (N_951,N_708,N_736);
nand U952 (N_952,N_714,N_767);
and U953 (N_953,N_623,N_635);
or U954 (N_954,N_747,N_680);
and U955 (N_955,N_781,N_713);
nand U956 (N_956,N_753,N_793);
nor U957 (N_957,N_627,N_795);
and U958 (N_958,N_680,N_778);
nand U959 (N_959,N_731,N_796);
nand U960 (N_960,N_781,N_799);
and U961 (N_961,N_664,N_731);
xor U962 (N_962,N_725,N_688);
nor U963 (N_963,N_736,N_683);
and U964 (N_964,N_733,N_734);
or U965 (N_965,N_660,N_796);
and U966 (N_966,N_633,N_680);
and U967 (N_967,N_691,N_660);
or U968 (N_968,N_696,N_637);
nor U969 (N_969,N_619,N_761);
and U970 (N_970,N_614,N_783);
nor U971 (N_971,N_683,N_627);
nand U972 (N_972,N_667,N_649);
and U973 (N_973,N_765,N_792);
nor U974 (N_974,N_705,N_787);
nand U975 (N_975,N_641,N_742);
and U976 (N_976,N_786,N_653);
and U977 (N_977,N_774,N_741);
or U978 (N_978,N_717,N_624);
nor U979 (N_979,N_650,N_680);
and U980 (N_980,N_608,N_702);
nor U981 (N_981,N_666,N_605);
and U982 (N_982,N_706,N_789);
xnor U983 (N_983,N_670,N_676);
nand U984 (N_984,N_729,N_660);
nor U985 (N_985,N_649,N_669);
or U986 (N_986,N_645,N_744);
and U987 (N_987,N_629,N_739);
or U988 (N_988,N_730,N_718);
xor U989 (N_989,N_763,N_600);
and U990 (N_990,N_770,N_749);
and U991 (N_991,N_658,N_721);
nor U992 (N_992,N_674,N_629);
or U993 (N_993,N_665,N_789);
xnor U994 (N_994,N_799,N_684);
nor U995 (N_995,N_656,N_704);
or U996 (N_996,N_631,N_696);
or U997 (N_997,N_784,N_789);
nor U998 (N_998,N_600,N_706);
nand U999 (N_999,N_751,N_674);
nor U1000 (N_1000,N_891,N_880);
and U1001 (N_1001,N_860,N_994);
or U1002 (N_1002,N_984,N_900);
nor U1003 (N_1003,N_955,N_960);
xor U1004 (N_1004,N_863,N_950);
xor U1005 (N_1005,N_818,N_911);
or U1006 (N_1006,N_872,N_892);
or U1007 (N_1007,N_839,N_884);
nand U1008 (N_1008,N_901,N_967);
and U1009 (N_1009,N_992,N_837);
nand U1010 (N_1010,N_938,N_931);
nor U1011 (N_1011,N_914,N_954);
or U1012 (N_1012,N_831,N_993);
nor U1013 (N_1013,N_951,N_867);
or U1014 (N_1014,N_824,N_963);
nand U1015 (N_1015,N_836,N_856);
and U1016 (N_1016,N_919,N_943);
nor U1017 (N_1017,N_851,N_999);
nand U1018 (N_1018,N_998,N_897);
or U1019 (N_1019,N_945,N_826);
nand U1020 (N_1020,N_811,N_959);
or U1021 (N_1021,N_868,N_940);
and U1022 (N_1022,N_822,N_847);
and U1023 (N_1023,N_854,N_991);
and U1024 (N_1024,N_917,N_965);
nand U1025 (N_1025,N_935,N_913);
nor U1026 (N_1026,N_934,N_846);
nor U1027 (N_1027,N_923,N_823);
and U1028 (N_1028,N_812,N_870);
nor U1029 (N_1029,N_980,N_956);
nand U1030 (N_1030,N_842,N_909);
and U1031 (N_1031,N_835,N_930);
or U1032 (N_1032,N_850,N_804);
and U1033 (N_1033,N_838,N_957);
or U1034 (N_1034,N_876,N_948);
and U1035 (N_1035,N_875,N_982);
and U1036 (N_1036,N_849,N_886);
xnor U1037 (N_1037,N_926,N_979);
nor U1038 (N_1038,N_987,N_974);
or U1039 (N_1039,N_918,N_820);
or U1040 (N_1040,N_933,N_903);
nand U1041 (N_1041,N_962,N_958);
nand U1042 (N_1042,N_883,N_888);
nand U1043 (N_1043,N_882,N_961);
nand U1044 (N_1044,N_809,N_869);
or U1045 (N_1045,N_852,N_893);
nand U1046 (N_1046,N_819,N_977);
nand U1047 (N_1047,N_828,N_830);
or U1048 (N_1048,N_827,N_801);
nand U1049 (N_1049,N_898,N_953);
nor U1050 (N_1050,N_966,N_881);
xnor U1051 (N_1051,N_952,N_825);
nand U1052 (N_1052,N_928,N_990);
or U1053 (N_1053,N_920,N_871);
nand U1054 (N_1054,N_986,N_932);
nand U1055 (N_1055,N_877,N_803);
nor U1056 (N_1056,N_807,N_978);
nand U1057 (N_1057,N_816,N_906);
or U1058 (N_1058,N_908,N_814);
or U1059 (N_1059,N_939,N_997);
or U1060 (N_1060,N_834,N_857);
nand U1061 (N_1061,N_910,N_995);
or U1062 (N_1062,N_896,N_879);
nor U1063 (N_1063,N_848,N_971);
xnor U1064 (N_1064,N_976,N_996);
and U1065 (N_1065,N_844,N_975);
and U1066 (N_1066,N_887,N_968);
xnor U1067 (N_1067,N_821,N_817);
nor U1068 (N_1068,N_813,N_806);
xor U1069 (N_1069,N_983,N_989);
and U1070 (N_1070,N_865,N_853);
xnor U1071 (N_1071,N_944,N_829);
and U1072 (N_1072,N_942,N_915);
and U1073 (N_1073,N_840,N_805);
or U1074 (N_1074,N_985,N_890);
or U1075 (N_1075,N_833,N_845);
or U1076 (N_1076,N_929,N_802);
nand U1077 (N_1077,N_907,N_899);
nand U1078 (N_1078,N_921,N_964);
nor U1079 (N_1079,N_878,N_946);
xnor U1080 (N_1080,N_937,N_949);
nand U1081 (N_1081,N_832,N_894);
nor U1082 (N_1082,N_841,N_861);
nand U1083 (N_1083,N_810,N_889);
or U1084 (N_1084,N_916,N_947);
nand U1085 (N_1085,N_808,N_862);
xor U1086 (N_1086,N_873,N_858);
xnor U1087 (N_1087,N_843,N_855);
or U1088 (N_1088,N_866,N_902);
and U1089 (N_1089,N_859,N_904);
or U1090 (N_1090,N_927,N_981);
or U1091 (N_1091,N_972,N_864);
xnor U1092 (N_1092,N_815,N_925);
and U1093 (N_1093,N_988,N_874);
xor U1094 (N_1094,N_973,N_885);
xor U1095 (N_1095,N_922,N_905);
xor U1096 (N_1096,N_969,N_970);
nand U1097 (N_1097,N_912,N_924);
or U1098 (N_1098,N_936,N_941);
xor U1099 (N_1099,N_895,N_800);
and U1100 (N_1100,N_860,N_882);
and U1101 (N_1101,N_878,N_922);
and U1102 (N_1102,N_866,N_826);
nand U1103 (N_1103,N_868,N_867);
nor U1104 (N_1104,N_952,N_850);
nor U1105 (N_1105,N_999,N_867);
nor U1106 (N_1106,N_982,N_899);
nand U1107 (N_1107,N_875,N_907);
and U1108 (N_1108,N_885,N_803);
and U1109 (N_1109,N_913,N_929);
or U1110 (N_1110,N_840,N_995);
nand U1111 (N_1111,N_891,N_903);
nand U1112 (N_1112,N_923,N_974);
nand U1113 (N_1113,N_937,N_962);
xor U1114 (N_1114,N_993,N_971);
nand U1115 (N_1115,N_923,N_808);
and U1116 (N_1116,N_837,N_867);
and U1117 (N_1117,N_935,N_839);
nand U1118 (N_1118,N_900,N_993);
nand U1119 (N_1119,N_884,N_974);
or U1120 (N_1120,N_820,N_938);
nor U1121 (N_1121,N_964,N_816);
and U1122 (N_1122,N_946,N_929);
and U1123 (N_1123,N_884,N_858);
or U1124 (N_1124,N_994,N_874);
or U1125 (N_1125,N_937,N_822);
or U1126 (N_1126,N_822,N_961);
or U1127 (N_1127,N_959,N_883);
and U1128 (N_1128,N_892,N_933);
xnor U1129 (N_1129,N_998,N_865);
nor U1130 (N_1130,N_923,N_986);
nand U1131 (N_1131,N_844,N_983);
nand U1132 (N_1132,N_850,N_890);
and U1133 (N_1133,N_992,N_945);
or U1134 (N_1134,N_809,N_802);
nand U1135 (N_1135,N_993,N_807);
xor U1136 (N_1136,N_896,N_923);
nor U1137 (N_1137,N_962,N_977);
nand U1138 (N_1138,N_861,N_883);
or U1139 (N_1139,N_888,N_802);
nand U1140 (N_1140,N_998,N_931);
nor U1141 (N_1141,N_860,N_880);
or U1142 (N_1142,N_833,N_972);
nor U1143 (N_1143,N_843,N_952);
nand U1144 (N_1144,N_920,N_882);
nor U1145 (N_1145,N_853,N_856);
nor U1146 (N_1146,N_916,N_927);
or U1147 (N_1147,N_962,N_840);
nand U1148 (N_1148,N_906,N_855);
and U1149 (N_1149,N_833,N_848);
nor U1150 (N_1150,N_921,N_945);
or U1151 (N_1151,N_808,N_996);
xnor U1152 (N_1152,N_938,N_809);
nor U1153 (N_1153,N_872,N_850);
nand U1154 (N_1154,N_930,N_944);
xnor U1155 (N_1155,N_916,N_905);
nand U1156 (N_1156,N_863,N_875);
or U1157 (N_1157,N_921,N_850);
or U1158 (N_1158,N_916,N_811);
nor U1159 (N_1159,N_925,N_814);
and U1160 (N_1160,N_824,N_823);
and U1161 (N_1161,N_962,N_975);
nor U1162 (N_1162,N_822,N_869);
nor U1163 (N_1163,N_917,N_989);
nand U1164 (N_1164,N_960,N_934);
or U1165 (N_1165,N_924,N_955);
or U1166 (N_1166,N_900,N_946);
nand U1167 (N_1167,N_846,N_925);
nand U1168 (N_1168,N_987,N_909);
and U1169 (N_1169,N_800,N_848);
or U1170 (N_1170,N_887,N_903);
nand U1171 (N_1171,N_842,N_968);
or U1172 (N_1172,N_970,N_872);
or U1173 (N_1173,N_967,N_817);
nand U1174 (N_1174,N_887,N_959);
nand U1175 (N_1175,N_802,N_988);
and U1176 (N_1176,N_960,N_949);
nor U1177 (N_1177,N_987,N_975);
and U1178 (N_1178,N_809,N_912);
nor U1179 (N_1179,N_928,N_848);
nand U1180 (N_1180,N_982,N_957);
and U1181 (N_1181,N_854,N_962);
nor U1182 (N_1182,N_886,N_969);
nand U1183 (N_1183,N_999,N_969);
or U1184 (N_1184,N_844,N_984);
or U1185 (N_1185,N_932,N_822);
xnor U1186 (N_1186,N_901,N_955);
or U1187 (N_1187,N_921,N_829);
nor U1188 (N_1188,N_998,N_905);
xor U1189 (N_1189,N_982,N_935);
nand U1190 (N_1190,N_891,N_993);
and U1191 (N_1191,N_906,N_896);
or U1192 (N_1192,N_843,N_936);
and U1193 (N_1193,N_916,N_989);
or U1194 (N_1194,N_941,N_921);
or U1195 (N_1195,N_985,N_995);
nor U1196 (N_1196,N_875,N_858);
and U1197 (N_1197,N_906,N_872);
nand U1198 (N_1198,N_940,N_816);
and U1199 (N_1199,N_820,N_870);
nand U1200 (N_1200,N_1049,N_1152);
or U1201 (N_1201,N_1051,N_1039);
nand U1202 (N_1202,N_1158,N_1025);
xnor U1203 (N_1203,N_1035,N_1074);
and U1204 (N_1204,N_1069,N_1160);
xnor U1205 (N_1205,N_1161,N_1080);
nand U1206 (N_1206,N_1113,N_1064);
xor U1207 (N_1207,N_1185,N_1166);
and U1208 (N_1208,N_1001,N_1148);
nor U1209 (N_1209,N_1055,N_1177);
nor U1210 (N_1210,N_1184,N_1193);
or U1211 (N_1211,N_1116,N_1014);
xor U1212 (N_1212,N_1156,N_1186);
nand U1213 (N_1213,N_1173,N_1151);
nor U1214 (N_1214,N_1023,N_1136);
nand U1215 (N_1215,N_1190,N_1098);
or U1216 (N_1216,N_1128,N_1005);
and U1217 (N_1217,N_1092,N_1077);
and U1218 (N_1218,N_1149,N_1171);
and U1219 (N_1219,N_1181,N_1018);
nor U1220 (N_1220,N_1119,N_1107);
nand U1221 (N_1221,N_1199,N_1118);
or U1222 (N_1222,N_1006,N_1110);
xor U1223 (N_1223,N_1137,N_1115);
xor U1224 (N_1224,N_1143,N_1083);
or U1225 (N_1225,N_1062,N_1026);
or U1226 (N_1226,N_1078,N_1093);
nand U1227 (N_1227,N_1060,N_1102);
and U1228 (N_1228,N_1042,N_1073);
and U1229 (N_1229,N_1129,N_1157);
xnor U1230 (N_1230,N_1163,N_1133);
nand U1231 (N_1231,N_1033,N_1147);
nor U1232 (N_1232,N_1135,N_1013);
nand U1233 (N_1233,N_1031,N_1117);
and U1234 (N_1234,N_1121,N_1086);
nor U1235 (N_1235,N_1144,N_1057);
nand U1236 (N_1236,N_1141,N_1027);
xor U1237 (N_1237,N_1139,N_1187);
and U1238 (N_1238,N_1179,N_1066);
or U1239 (N_1239,N_1071,N_1021);
or U1240 (N_1240,N_1132,N_1089);
and U1241 (N_1241,N_1094,N_1159);
nor U1242 (N_1242,N_1038,N_1106);
nor U1243 (N_1243,N_1036,N_1032);
and U1244 (N_1244,N_1088,N_1154);
and U1245 (N_1245,N_1120,N_1097);
nor U1246 (N_1246,N_1010,N_1056);
xor U1247 (N_1247,N_1146,N_1020);
nand U1248 (N_1248,N_1114,N_1198);
and U1249 (N_1249,N_1180,N_1170);
or U1250 (N_1250,N_1101,N_1046);
xnor U1251 (N_1251,N_1048,N_1167);
nor U1252 (N_1252,N_1007,N_1168);
or U1253 (N_1253,N_1019,N_1029);
or U1254 (N_1254,N_1075,N_1095);
and U1255 (N_1255,N_1124,N_1043);
or U1256 (N_1256,N_1068,N_1105);
and U1257 (N_1257,N_1002,N_1197);
nor U1258 (N_1258,N_1053,N_1090);
nand U1259 (N_1259,N_1155,N_1150);
nand U1260 (N_1260,N_1194,N_1134);
or U1261 (N_1261,N_1003,N_1126);
and U1262 (N_1262,N_1065,N_1070);
nor U1263 (N_1263,N_1131,N_1008);
or U1264 (N_1264,N_1153,N_1044);
nor U1265 (N_1265,N_1176,N_1047);
xor U1266 (N_1266,N_1028,N_1109);
nor U1267 (N_1267,N_1175,N_1045);
or U1268 (N_1268,N_1054,N_1063);
nand U1269 (N_1269,N_1082,N_1041);
nor U1270 (N_1270,N_1091,N_1059);
or U1271 (N_1271,N_1081,N_1191);
nand U1272 (N_1272,N_1112,N_1084);
and U1273 (N_1273,N_1009,N_1079);
nand U1274 (N_1274,N_1192,N_1122);
nand U1275 (N_1275,N_1174,N_1030);
or U1276 (N_1276,N_1016,N_1172);
and U1277 (N_1277,N_1015,N_1164);
nand U1278 (N_1278,N_1024,N_1058);
and U1279 (N_1279,N_1096,N_1076);
and U1280 (N_1280,N_1145,N_1012);
xor U1281 (N_1281,N_1034,N_1104);
or U1282 (N_1282,N_1138,N_1188);
nand U1283 (N_1283,N_1189,N_1085);
nand U1284 (N_1284,N_1142,N_1127);
nor U1285 (N_1285,N_1037,N_1011);
nor U1286 (N_1286,N_1140,N_1162);
or U1287 (N_1287,N_1072,N_1040);
or U1288 (N_1288,N_1123,N_1050);
nor U1289 (N_1289,N_1108,N_1111);
xor U1290 (N_1290,N_1004,N_1100);
nor U1291 (N_1291,N_1195,N_1125);
and U1292 (N_1292,N_1182,N_1183);
xor U1293 (N_1293,N_1165,N_1087);
nand U1294 (N_1294,N_1178,N_1052);
nor U1295 (N_1295,N_1017,N_1099);
nand U1296 (N_1296,N_1130,N_1061);
and U1297 (N_1297,N_1196,N_1022);
nor U1298 (N_1298,N_1169,N_1000);
or U1299 (N_1299,N_1103,N_1067);
nand U1300 (N_1300,N_1000,N_1007);
nor U1301 (N_1301,N_1075,N_1023);
nor U1302 (N_1302,N_1119,N_1148);
or U1303 (N_1303,N_1199,N_1197);
or U1304 (N_1304,N_1061,N_1111);
xnor U1305 (N_1305,N_1062,N_1141);
or U1306 (N_1306,N_1091,N_1008);
nor U1307 (N_1307,N_1051,N_1050);
xor U1308 (N_1308,N_1139,N_1010);
or U1309 (N_1309,N_1038,N_1012);
or U1310 (N_1310,N_1193,N_1095);
nand U1311 (N_1311,N_1174,N_1042);
nor U1312 (N_1312,N_1093,N_1198);
nor U1313 (N_1313,N_1090,N_1004);
and U1314 (N_1314,N_1010,N_1008);
nand U1315 (N_1315,N_1191,N_1041);
or U1316 (N_1316,N_1192,N_1121);
nand U1317 (N_1317,N_1092,N_1154);
nor U1318 (N_1318,N_1075,N_1051);
or U1319 (N_1319,N_1125,N_1047);
nor U1320 (N_1320,N_1111,N_1066);
or U1321 (N_1321,N_1061,N_1042);
or U1322 (N_1322,N_1012,N_1029);
nor U1323 (N_1323,N_1002,N_1096);
nor U1324 (N_1324,N_1005,N_1074);
nor U1325 (N_1325,N_1185,N_1189);
nor U1326 (N_1326,N_1078,N_1046);
or U1327 (N_1327,N_1055,N_1000);
nand U1328 (N_1328,N_1032,N_1113);
or U1329 (N_1329,N_1044,N_1081);
nand U1330 (N_1330,N_1067,N_1094);
or U1331 (N_1331,N_1050,N_1120);
nor U1332 (N_1332,N_1013,N_1181);
nand U1333 (N_1333,N_1172,N_1165);
and U1334 (N_1334,N_1181,N_1031);
nand U1335 (N_1335,N_1131,N_1109);
nor U1336 (N_1336,N_1182,N_1164);
and U1337 (N_1337,N_1109,N_1162);
and U1338 (N_1338,N_1137,N_1107);
and U1339 (N_1339,N_1117,N_1197);
or U1340 (N_1340,N_1071,N_1133);
and U1341 (N_1341,N_1134,N_1083);
nand U1342 (N_1342,N_1129,N_1195);
and U1343 (N_1343,N_1106,N_1050);
nand U1344 (N_1344,N_1130,N_1018);
nor U1345 (N_1345,N_1136,N_1078);
nand U1346 (N_1346,N_1077,N_1005);
or U1347 (N_1347,N_1097,N_1059);
nand U1348 (N_1348,N_1172,N_1002);
nor U1349 (N_1349,N_1188,N_1106);
and U1350 (N_1350,N_1144,N_1190);
nand U1351 (N_1351,N_1128,N_1150);
or U1352 (N_1352,N_1132,N_1164);
nand U1353 (N_1353,N_1014,N_1007);
xnor U1354 (N_1354,N_1002,N_1133);
nor U1355 (N_1355,N_1023,N_1183);
nor U1356 (N_1356,N_1195,N_1032);
nor U1357 (N_1357,N_1197,N_1086);
or U1358 (N_1358,N_1168,N_1125);
or U1359 (N_1359,N_1004,N_1000);
nor U1360 (N_1360,N_1052,N_1050);
nor U1361 (N_1361,N_1041,N_1061);
xor U1362 (N_1362,N_1198,N_1146);
nand U1363 (N_1363,N_1036,N_1011);
nand U1364 (N_1364,N_1150,N_1070);
nand U1365 (N_1365,N_1041,N_1071);
xnor U1366 (N_1366,N_1134,N_1106);
nor U1367 (N_1367,N_1185,N_1089);
xor U1368 (N_1368,N_1117,N_1006);
nand U1369 (N_1369,N_1002,N_1081);
nor U1370 (N_1370,N_1114,N_1011);
nand U1371 (N_1371,N_1008,N_1004);
and U1372 (N_1372,N_1020,N_1025);
nor U1373 (N_1373,N_1155,N_1099);
or U1374 (N_1374,N_1125,N_1147);
and U1375 (N_1375,N_1052,N_1180);
xnor U1376 (N_1376,N_1091,N_1193);
nor U1377 (N_1377,N_1140,N_1148);
xor U1378 (N_1378,N_1168,N_1105);
nand U1379 (N_1379,N_1162,N_1185);
and U1380 (N_1380,N_1036,N_1171);
nand U1381 (N_1381,N_1184,N_1133);
nor U1382 (N_1382,N_1120,N_1139);
nand U1383 (N_1383,N_1174,N_1018);
or U1384 (N_1384,N_1180,N_1128);
and U1385 (N_1385,N_1079,N_1156);
xor U1386 (N_1386,N_1087,N_1126);
or U1387 (N_1387,N_1137,N_1076);
nor U1388 (N_1388,N_1140,N_1113);
nand U1389 (N_1389,N_1053,N_1040);
and U1390 (N_1390,N_1190,N_1177);
nor U1391 (N_1391,N_1059,N_1136);
xnor U1392 (N_1392,N_1148,N_1126);
nand U1393 (N_1393,N_1033,N_1110);
nand U1394 (N_1394,N_1123,N_1129);
nor U1395 (N_1395,N_1005,N_1033);
and U1396 (N_1396,N_1031,N_1198);
nor U1397 (N_1397,N_1198,N_1079);
xnor U1398 (N_1398,N_1057,N_1086);
or U1399 (N_1399,N_1087,N_1121);
nand U1400 (N_1400,N_1275,N_1224);
or U1401 (N_1401,N_1237,N_1351);
nor U1402 (N_1402,N_1213,N_1214);
and U1403 (N_1403,N_1359,N_1203);
nor U1404 (N_1404,N_1290,N_1233);
or U1405 (N_1405,N_1315,N_1368);
xnor U1406 (N_1406,N_1232,N_1243);
nand U1407 (N_1407,N_1209,N_1329);
and U1408 (N_1408,N_1254,N_1376);
nor U1409 (N_1409,N_1255,N_1364);
or U1410 (N_1410,N_1378,N_1317);
nand U1411 (N_1411,N_1305,N_1377);
nand U1412 (N_1412,N_1325,N_1216);
and U1413 (N_1413,N_1231,N_1293);
or U1414 (N_1414,N_1393,N_1373);
or U1415 (N_1415,N_1353,N_1263);
nor U1416 (N_1416,N_1265,N_1370);
nand U1417 (N_1417,N_1306,N_1331);
and U1418 (N_1418,N_1271,N_1355);
nor U1419 (N_1419,N_1383,N_1308);
nand U1420 (N_1420,N_1215,N_1225);
or U1421 (N_1421,N_1205,N_1270);
and U1422 (N_1422,N_1350,N_1365);
or U1423 (N_1423,N_1294,N_1330);
and U1424 (N_1424,N_1202,N_1210);
or U1425 (N_1425,N_1357,N_1391);
nor U1426 (N_1426,N_1399,N_1288);
nor U1427 (N_1427,N_1261,N_1274);
nor U1428 (N_1428,N_1312,N_1234);
and U1429 (N_1429,N_1239,N_1256);
nor U1430 (N_1430,N_1249,N_1314);
and U1431 (N_1431,N_1278,N_1208);
nand U1432 (N_1432,N_1387,N_1379);
or U1433 (N_1433,N_1339,N_1301);
or U1434 (N_1434,N_1326,N_1321);
and U1435 (N_1435,N_1366,N_1386);
nand U1436 (N_1436,N_1276,N_1253);
and U1437 (N_1437,N_1228,N_1303);
and U1438 (N_1438,N_1269,N_1240);
or U1439 (N_1439,N_1217,N_1259);
nor U1440 (N_1440,N_1338,N_1250);
nor U1441 (N_1441,N_1211,N_1349);
and U1442 (N_1442,N_1299,N_1251);
or U1443 (N_1443,N_1367,N_1374);
nor U1444 (N_1444,N_1345,N_1246);
and U1445 (N_1445,N_1398,N_1252);
or U1446 (N_1446,N_1392,N_1340);
and U1447 (N_1447,N_1284,N_1333);
nand U1448 (N_1448,N_1323,N_1341);
and U1449 (N_1449,N_1328,N_1244);
and U1450 (N_1450,N_1375,N_1313);
nand U1451 (N_1451,N_1226,N_1336);
xor U1452 (N_1452,N_1227,N_1298);
and U1453 (N_1453,N_1322,N_1230);
or U1454 (N_1454,N_1236,N_1277);
nand U1455 (N_1455,N_1245,N_1337);
xor U1456 (N_1456,N_1356,N_1334);
and U1457 (N_1457,N_1267,N_1382);
nor U1458 (N_1458,N_1319,N_1266);
and U1459 (N_1459,N_1289,N_1218);
nor U1460 (N_1460,N_1324,N_1384);
or U1461 (N_1461,N_1371,N_1248);
nand U1462 (N_1462,N_1343,N_1388);
or U1463 (N_1463,N_1242,N_1260);
nor U1464 (N_1464,N_1381,N_1396);
nor U1465 (N_1465,N_1241,N_1268);
nor U1466 (N_1466,N_1212,N_1332);
nor U1467 (N_1467,N_1354,N_1206);
nor U1468 (N_1468,N_1335,N_1297);
nand U1469 (N_1469,N_1258,N_1264);
nand U1470 (N_1470,N_1279,N_1280);
nor U1471 (N_1471,N_1307,N_1309);
nand U1472 (N_1472,N_1273,N_1281);
nand U1473 (N_1473,N_1296,N_1204);
or U1474 (N_1474,N_1229,N_1362);
and U1475 (N_1475,N_1344,N_1394);
nand U1476 (N_1476,N_1272,N_1347);
nor U1477 (N_1477,N_1286,N_1310);
or U1478 (N_1478,N_1395,N_1287);
xnor U1479 (N_1479,N_1300,N_1223);
nor U1480 (N_1480,N_1222,N_1257);
nor U1481 (N_1481,N_1295,N_1302);
nor U1482 (N_1482,N_1207,N_1363);
nand U1483 (N_1483,N_1358,N_1352);
and U1484 (N_1484,N_1235,N_1200);
nand U1485 (N_1485,N_1380,N_1348);
or U1486 (N_1486,N_1361,N_1282);
or U1487 (N_1487,N_1369,N_1262);
xnor U1488 (N_1488,N_1327,N_1247);
nand U1489 (N_1489,N_1318,N_1316);
nor U1490 (N_1490,N_1372,N_1304);
and U1491 (N_1491,N_1220,N_1346);
and U1492 (N_1492,N_1320,N_1360);
xor U1493 (N_1493,N_1342,N_1397);
nand U1494 (N_1494,N_1291,N_1285);
nor U1495 (N_1495,N_1238,N_1201);
or U1496 (N_1496,N_1385,N_1390);
nor U1497 (N_1497,N_1283,N_1292);
xnor U1498 (N_1498,N_1389,N_1219);
nand U1499 (N_1499,N_1221,N_1311);
or U1500 (N_1500,N_1221,N_1224);
nand U1501 (N_1501,N_1352,N_1217);
xnor U1502 (N_1502,N_1253,N_1228);
nor U1503 (N_1503,N_1346,N_1338);
and U1504 (N_1504,N_1262,N_1264);
and U1505 (N_1505,N_1238,N_1289);
or U1506 (N_1506,N_1351,N_1346);
or U1507 (N_1507,N_1342,N_1341);
or U1508 (N_1508,N_1249,N_1240);
and U1509 (N_1509,N_1256,N_1330);
xor U1510 (N_1510,N_1287,N_1267);
and U1511 (N_1511,N_1379,N_1310);
nand U1512 (N_1512,N_1235,N_1313);
nor U1513 (N_1513,N_1292,N_1399);
nand U1514 (N_1514,N_1387,N_1373);
nand U1515 (N_1515,N_1313,N_1303);
or U1516 (N_1516,N_1260,N_1206);
nand U1517 (N_1517,N_1285,N_1394);
nand U1518 (N_1518,N_1377,N_1320);
or U1519 (N_1519,N_1327,N_1221);
and U1520 (N_1520,N_1354,N_1279);
xnor U1521 (N_1521,N_1388,N_1332);
nor U1522 (N_1522,N_1289,N_1395);
nand U1523 (N_1523,N_1324,N_1357);
and U1524 (N_1524,N_1306,N_1227);
nor U1525 (N_1525,N_1345,N_1208);
nand U1526 (N_1526,N_1224,N_1388);
nand U1527 (N_1527,N_1353,N_1340);
xnor U1528 (N_1528,N_1210,N_1330);
and U1529 (N_1529,N_1287,N_1200);
nor U1530 (N_1530,N_1323,N_1329);
nand U1531 (N_1531,N_1302,N_1386);
and U1532 (N_1532,N_1281,N_1361);
or U1533 (N_1533,N_1231,N_1297);
and U1534 (N_1534,N_1279,N_1336);
or U1535 (N_1535,N_1384,N_1275);
nor U1536 (N_1536,N_1208,N_1313);
and U1537 (N_1537,N_1277,N_1373);
nand U1538 (N_1538,N_1217,N_1271);
and U1539 (N_1539,N_1270,N_1201);
nor U1540 (N_1540,N_1344,N_1288);
nand U1541 (N_1541,N_1347,N_1264);
or U1542 (N_1542,N_1324,N_1332);
nand U1543 (N_1543,N_1343,N_1200);
and U1544 (N_1544,N_1291,N_1215);
and U1545 (N_1545,N_1299,N_1203);
nor U1546 (N_1546,N_1297,N_1223);
nor U1547 (N_1547,N_1337,N_1326);
and U1548 (N_1548,N_1368,N_1281);
or U1549 (N_1549,N_1261,N_1322);
or U1550 (N_1550,N_1238,N_1343);
nor U1551 (N_1551,N_1212,N_1323);
nor U1552 (N_1552,N_1266,N_1388);
nor U1553 (N_1553,N_1276,N_1386);
nand U1554 (N_1554,N_1290,N_1382);
and U1555 (N_1555,N_1378,N_1286);
nand U1556 (N_1556,N_1212,N_1257);
nor U1557 (N_1557,N_1349,N_1311);
and U1558 (N_1558,N_1330,N_1262);
nor U1559 (N_1559,N_1222,N_1369);
nor U1560 (N_1560,N_1349,N_1382);
or U1561 (N_1561,N_1253,N_1377);
nor U1562 (N_1562,N_1250,N_1213);
or U1563 (N_1563,N_1269,N_1234);
and U1564 (N_1564,N_1337,N_1311);
nand U1565 (N_1565,N_1243,N_1397);
nand U1566 (N_1566,N_1315,N_1376);
and U1567 (N_1567,N_1247,N_1364);
or U1568 (N_1568,N_1368,N_1305);
xnor U1569 (N_1569,N_1283,N_1333);
nor U1570 (N_1570,N_1201,N_1317);
and U1571 (N_1571,N_1393,N_1361);
or U1572 (N_1572,N_1237,N_1332);
nand U1573 (N_1573,N_1308,N_1259);
nor U1574 (N_1574,N_1265,N_1315);
xnor U1575 (N_1575,N_1333,N_1259);
or U1576 (N_1576,N_1388,N_1207);
or U1577 (N_1577,N_1342,N_1214);
nor U1578 (N_1578,N_1280,N_1354);
nor U1579 (N_1579,N_1387,N_1300);
nor U1580 (N_1580,N_1241,N_1327);
and U1581 (N_1581,N_1242,N_1203);
nor U1582 (N_1582,N_1352,N_1331);
nand U1583 (N_1583,N_1201,N_1374);
nor U1584 (N_1584,N_1286,N_1380);
nand U1585 (N_1585,N_1204,N_1279);
nand U1586 (N_1586,N_1246,N_1230);
nor U1587 (N_1587,N_1324,N_1257);
xor U1588 (N_1588,N_1348,N_1204);
nand U1589 (N_1589,N_1337,N_1247);
nor U1590 (N_1590,N_1395,N_1320);
nor U1591 (N_1591,N_1274,N_1311);
and U1592 (N_1592,N_1387,N_1213);
nor U1593 (N_1593,N_1283,N_1374);
or U1594 (N_1594,N_1244,N_1287);
or U1595 (N_1595,N_1306,N_1337);
nor U1596 (N_1596,N_1399,N_1277);
nor U1597 (N_1597,N_1289,N_1247);
nand U1598 (N_1598,N_1366,N_1368);
nand U1599 (N_1599,N_1296,N_1376);
xnor U1600 (N_1600,N_1553,N_1448);
nor U1601 (N_1601,N_1402,N_1541);
nor U1602 (N_1602,N_1521,N_1539);
and U1603 (N_1603,N_1488,N_1540);
nor U1604 (N_1604,N_1595,N_1430);
nand U1605 (N_1605,N_1431,N_1561);
nand U1606 (N_1606,N_1442,N_1492);
and U1607 (N_1607,N_1481,N_1412);
xor U1608 (N_1608,N_1475,N_1422);
nor U1609 (N_1609,N_1571,N_1554);
nand U1610 (N_1610,N_1477,N_1400);
xnor U1611 (N_1611,N_1415,N_1580);
or U1612 (N_1612,N_1457,N_1545);
nor U1613 (N_1613,N_1567,N_1570);
or U1614 (N_1614,N_1487,N_1591);
nand U1615 (N_1615,N_1516,N_1432);
nor U1616 (N_1616,N_1537,N_1526);
and U1617 (N_1617,N_1417,N_1564);
nand U1618 (N_1618,N_1505,N_1584);
and U1619 (N_1619,N_1520,N_1445);
nor U1620 (N_1620,N_1529,N_1440);
and U1621 (N_1621,N_1557,N_1597);
or U1622 (N_1622,N_1522,N_1453);
xnor U1623 (N_1623,N_1456,N_1506);
nand U1624 (N_1624,N_1588,N_1474);
nor U1625 (N_1625,N_1427,N_1579);
nor U1626 (N_1626,N_1424,N_1425);
and U1627 (N_1627,N_1443,N_1414);
xnor U1628 (N_1628,N_1490,N_1444);
nor U1629 (N_1629,N_1573,N_1596);
or U1630 (N_1630,N_1583,N_1433);
or U1631 (N_1631,N_1404,N_1519);
or U1632 (N_1632,N_1503,N_1403);
nor U1633 (N_1633,N_1578,N_1501);
nand U1634 (N_1634,N_1439,N_1507);
and U1635 (N_1635,N_1418,N_1484);
and U1636 (N_1636,N_1437,N_1461);
and U1637 (N_1637,N_1462,N_1426);
nor U1638 (N_1638,N_1502,N_1435);
nor U1639 (N_1639,N_1464,N_1500);
or U1640 (N_1640,N_1528,N_1480);
or U1641 (N_1641,N_1458,N_1574);
or U1642 (N_1642,N_1509,N_1504);
and U1643 (N_1643,N_1548,N_1586);
nand U1644 (N_1644,N_1550,N_1482);
nand U1645 (N_1645,N_1486,N_1568);
nand U1646 (N_1646,N_1441,N_1581);
xor U1647 (N_1647,N_1410,N_1523);
xor U1648 (N_1648,N_1423,N_1562);
and U1649 (N_1649,N_1429,N_1483);
and U1650 (N_1650,N_1473,N_1498);
nand U1651 (N_1651,N_1447,N_1497);
and U1652 (N_1652,N_1534,N_1416);
nand U1653 (N_1653,N_1585,N_1589);
nand U1654 (N_1654,N_1552,N_1547);
or U1655 (N_1655,N_1555,N_1476);
and U1656 (N_1656,N_1560,N_1434);
nand U1657 (N_1657,N_1599,N_1544);
nor U1658 (N_1658,N_1405,N_1499);
or U1659 (N_1659,N_1489,N_1452);
nor U1660 (N_1660,N_1408,N_1455);
nand U1661 (N_1661,N_1590,N_1470);
nor U1662 (N_1662,N_1546,N_1517);
and U1663 (N_1663,N_1469,N_1536);
nand U1664 (N_1664,N_1575,N_1446);
and U1665 (N_1665,N_1420,N_1438);
and U1666 (N_1666,N_1479,N_1496);
nand U1667 (N_1667,N_1592,N_1563);
and U1668 (N_1668,N_1511,N_1594);
and U1669 (N_1669,N_1454,N_1485);
nand U1670 (N_1670,N_1450,N_1530);
nor U1671 (N_1671,N_1508,N_1472);
xor U1672 (N_1672,N_1465,N_1510);
nand U1673 (N_1673,N_1524,N_1538);
nand U1674 (N_1674,N_1466,N_1535);
and U1675 (N_1675,N_1593,N_1569);
or U1676 (N_1676,N_1467,N_1478);
xor U1677 (N_1677,N_1542,N_1468);
nand U1678 (N_1678,N_1566,N_1471);
nor U1679 (N_1679,N_1577,N_1525);
or U1680 (N_1680,N_1436,N_1419);
nor U1681 (N_1681,N_1551,N_1543);
and U1682 (N_1682,N_1559,N_1518);
nor U1683 (N_1683,N_1532,N_1463);
or U1684 (N_1684,N_1406,N_1576);
or U1685 (N_1685,N_1598,N_1533);
nand U1686 (N_1686,N_1401,N_1582);
nor U1687 (N_1687,N_1411,N_1459);
nor U1688 (N_1688,N_1556,N_1587);
or U1689 (N_1689,N_1460,N_1558);
nand U1690 (N_1690,N_1565,N_1495);
nor U1691 (N_1691,N_1549,N_1513);
xnor U1692 (N_1692,N_1413,N_1531);
nor U1693 (N_1693,N_1493,N_1449);
or U1694 (N_1694,N_1512,N_1572);
nor U1695 (N_1695,N_1515,N_1409);
and U1696 (N_1696,N_1491,N_1428);
nor U1697 (N_1697,N_1527,N_1494);
nor U1698 (N_1698,N_1514,N_1451);
and U1699 (N_1699,N_1421,N_1407);
nor U1700 (N_1700,N_1535,N_1438);
or U1701 (N_1701,N_1574,N_1468);
nor U1702 (N_1702,N_1528,N_1401);
and U1703 (N_1703,N_1541,N_1453);
nor U1704 (N_1704,N_1540,N_1558);
and U1705 (N_1705,N_1432,N_1444);
nor U1706 (N_1706,N_1518,N_1599);
nand U1707 (N_1707,N_1413,N_1479);
or U1708 (N_1708,N_1584,N_1554);
nand U1709 (N_1709,N_1413,N_1597);
nor U1710 (N_1710,N_1526,N_1481);
nand U1711 (N_1711,N_1415,N_1491);
nor U1712 (N_1712,N_1434,N_1562);
nand U1713 (N_1713,N_1515,N_1456);
nand U1714 (N_1714,N_1529,N_1485);
nor U1715 (N_1715,N_1467,N_1432);
and U1716 (N_1716,N_1465,N_1505);
nor U1717 (N_1717,N_1470,N_1413);
nand U1718 (N_1718,N_1446,N_1544);
nor U1719 (N_1719,N_1468,N_1505);
xnor U1720 (N_1720,N_1533,N_1453);
and U1721 (N_1721,N_1420,N_1491);
or U1722 (N_1722,N_1482,N_1418);
or U1723 (N_1723,N_1452,N_1410);
or U1724 (N_1724,N_1543,N_1456);
nand U1725 (N_1725,N_1401,N_1520);
nor U1726 (N_1726,N_1553,N_1478);
or U1727 (N_1727,N_1459,N_1498);
nor U1728 (N_1728,N_1571,N_1458);
nand U1729 (N_1729,N_1515,N_1433);
nor U1730 (N_1730,N_1466,N_1534);
and U1731 (N_1731,N_1419,N_1476);
nor U1732 (N_1732,N_1598,N_1559);
and U1733 (N_1733,N_1401,N_1564);
nand U1734 (N_1734,N_1508,N_1494);
or U1735 (N_1735,N_1516,N_1565);
nand U1736 (N_1736,N_1589,N_1411);
nand U1737 (N_1737,N_1473,N_1574);
nand U1738 (N_1738,N_1525,N_1503);
nand U1739 (N_1739,N_1412,N_1485);
and U1740 (N_1740,N_1478,N_1534);
and U1741 (N_1741,N_1458,N_1506);
nand U1742 (N_1742,N_1598,N_1561);
or U1743 (N_1743,N_1494,N_1439);
nand U1744 (N_1744,N_1451,N_1527);
and U1745 (N_1745,N_1491,N_1439);
and U1746 (N_1746,N_1590,N_1485);
nand U1747 (N_1747,N_1438,N_1575);
nand U1748 (N_1748,N_1476,N_1499);
xnor U1749 (N_1749,N_1547,N_1580);
nand U1750 (N_1750,N_1558,N_1409);
and U1751 (N_1751,N_1561,N_1569);
xor U1752 (N_1752,N_1523,N_1541);
nor U1753 (N_1753,N_1483,N_1572);
or U1754 (N_1754,N_1484,N_1572);
nand U1755 (N_1755,N_1585,N_1530);
nand U1756 (N_1756,N_1400,N_1519);
xnor U1757 (N_1757,N_1545,N_1419);
or U1758 (N_1758,N_1409,N_1505);
and U1759 (N_1759,N_1489,N_1479);
nor U1760 (N_1760,N_1520,N_1428);
xnor U1761 (N_1761,N_1464,N_1538);
xor U1762 (N_1762,N_1580,N_1516);
nand U1763 (N_1763,N_1577,N_1540);
and U1764 (N_1764,N_1530,N_1461);
nor U1765 (N_1765,N_1472,N_1422);
or U1766 (N_1766,N_1507,N_1556);
or U1767 (N_1767,N_1491,N_1551);
or U1768 (N_1768,N_1489,N_1424);
xnor U1769 (N_1769,N_1555,N_1578);
nand U1770 (N_1770,N_1446,N_1579);
nor U1771 (N_1771,N_1424,N_1478);
and U1772 (N_1772,N_1562,N_1447);
or U1773 (N_1773,N_1484,N_1459);
nor U1774 (N_1774,N_1491,N_1587);
or U1775 (N_1775,N_1400,N_1501);
nand U1776 (N_1776,N_1476,N_1444);
nand U1777 (N_1777,N_1565,N_1533);
and U1778 (N_1778,N_1563,N_1515);
nand U1779 (N_1779,N_1495,N_1551);
nor U1780 (N_1780,N_1453,N_1587);
and U1781 (N_1781,N_1532,N_1497);
nor U1782 (N_1782,N_1483,N_1597);
or U1783 (N_1783,N_1548,N_1468);
and U1784 (N_1784,N_1565,N_1446);
nor U1785 (N_1785,N_1589,N_1497);
or U1786 (N_1786,N_1464,N_1430);
nand U1787 (N_1787,N_1402,N_1436);
xor U1788 (N_1788,N_1495,N_1406);
nand U1789 (N_1789,N_1503,N_1504);
nor U1790 (N_1790,N_1566,N_1432);
nand U1791 (N_1791,N_1451,N_1463);
or U1792 (N_1792,N_1582,N_1513);
or U1793 (N_1793,N_1425,N_1554);
or U1794 (N_1794,N_1575,N_1523);
nand U1795 (N_1795,N_1588,N_1485);
and U1796 (N_1796,N_1411,N_1406);
and U1797 (N_1797,N_1411,N_1543);
nand U1798 (N_1798,N_1488,N_1444);
or U1799 (N_1799,N_1534,N_1596);
or U1800 (N_1800,N_1621,N_1722);
and U1801 (N_1801,N_1764,N_1692);
nor U1802 (N_1802,N_1627,N_1626);
or U1803 (N_1803,N_1675,N_1618);
nor U1804 (N_1804,N_1700,N_1744);
or U1805 (N_1805,N_1754,N_1645);
nand U1806 (N_1806,N_1688,N_1625);
or U1807 (N_1807,N_1767,N_1638);
and U1808 (N_1808,N_1710,N_1765);
nand U1809 (N_1809,N_1720,N_1619);
and U1810 (N_1810,N_1676,N_1751);
nand U1811 (N_1811,N_1707,N_1745);
or U1812 (N_1812,N_1736,N_1723);
nand U1813 (N_1813,N_1602,N_1662);
or U1814 (N_1814,N_1795,N_1660);
or U1815 (N_1815,N_1622,N_1652);
nor U1816 (N_1816,N_1641,N_1709);
nor U1817 (N_1817,N_1642,N_1646);
or U1818 (N_1818,N_1636,N_1753);
and U1819 (N_1819,N_1718,N_1682);
or U1820 (N_1820,N_1649,N_1631);
nor U1821 (N_1821,N_1686,N_1677);
and U1822 (N_1822,N_1726,N_1609);
xnor U1823 (N_1823,N_1670,N_1797);
xnor U1824 (N_1824,N_1773,N_1613);
and U1825 (N_1825,N_1712,N_1724);
nor U1826 (N_1826,N_1664,N_1655);
or U1827 (N_1827,N_1721,N_1786);
or U1828 (N_1828,N_1766,N_1789);
nand U1829 (N_1829,N_1693,N_1635);
xor U1830 (N_1830,N_1787,N_1782);
or U1831 (N_1831,N_1615,N_1672);
nor U1832 (N_1832,N_1762,N_1623);
or U1833 (N_1833,N_1630,N_1796);
nor U1834 (N_1834,N_1603,N_1794);
nand U1835 (N_1835,N_1772,N_1757);
and U1836 (N_1836,N_1737,N_1654);
and U1837 (N_1837,N_1628,N_1756);
or U1838 (N_1838,N_1759,N_1705);
nand U1839 (N_1839,N_1774,N_1658);
nand U1840 (N_1840,N_1616,N_1763);
nor U1841 (N_1841,N_1606,N_1699);
nor U1842 (N_1842,N_1634,N_1768);
nor U1843 (N_1843,N_1777,N_1637);
and U1844 (N_1844,N_1708,N_1743);
nand U1845 (N_1845,N_1632,N_1650);
nor U1846 (N_1846,N_1669,N_1730);
nor U1847 (N_1847,N_1780,N_1758);
xnor U1848 (N_1848,N_1680,N_1770);
nand U1849 (N_1849,N_1716,N_1776);
or U1850 (N_1850,N_1704,N_1719);
or U1851 (N_1851,N_1694,N_1798);
or U1852 (N_1852,N_1614,N_1760);
or U1853 (N_1853,N_1701,N_1728);
nand U1854 (N_1854,N_1746,N_1689);
nand U1855 (N_1855,N_1741,N_1799);
nand U1856 (N_1856,N_1775,N_1729);
or U1857 (N_1857,N_1666,N_1706);
nor U1858 (N_1858,N_1752,N_1749);
xnor U1859 (N_1859,N_1792,N_1674);
nor U1860 (N_1860,N_1715,N_1713);
nand U1861 (N_1861,N_1673,N_1651);
or U1862 (N_1862,N_1617,N_1633);
nor U1863 (N_1863,N_1656,N_1604);
and U1864 (N_1864,N_1717,N_1690);
nor U1865 (N_1865,N_1600,N_1734);
xnor U1866 (N_1866,N_1607,N_1711);
and U1867 (N_1867,N_1608,N_1648);
nand U1868 (N_1868,N_1769,N_1755);
and U1869 (N_1869,N_1647,N_1747);
nand U1870 (N_1870,N_1742,N_1684);
nor U1871 (N_1871,N_1748,N_1731);
nor U1872 (N_1872,N_1791,N_1643);
or U1873 (N_1873,N_1653,N_1702);
nand U1874 (N_1874,N_1668,N_1685);
or U1875 (N_1875,N_1679,N_1629);
nor U1876 (N_1876,N_1624,N_1659);
and U1877 (N_1877,N_1605,N_1620);
or U1878 (N_1878,N_1683,N_1783);
or U1879 (N_1879,N_1714,N_1644);
nor U1880 (N_1880,N_1771,N_1739);
nand U1881 (N_1881,N_1703,N_1778);
nor U1882 (N_1882,N_1667,N_1678);
and U1883 (N_1883,N_1725,N_1698);
nand U1884 (N_1884,N_1639,N_1695);
xnor U1885 (N_1885,N_1732,N_1750);
and U1886 (N_1886,N_1611,N_1697);
or U1887 (N_1887,N_1671,N_1681);
nand U1888 (N_1888,N_1665,N_1610);
and U1889 (N_1889,N_1687,N_1761);
nor U1890 (N_1890,N_1691,N_1784);
nor U1891 (N_1891,N_1612,N_1785);
nor U1892 (N_1892,N_1661,N_1640);
and U1893 (N_1893,N_1779,N_1781);
xnor U1894 (N_1894,N_1727,N_1738);
nor U1895 (N_1895,N_1663,N_1733);
and U1896 (N_1896,N_1735,N_1740);
nor U1897 (N_1897,N_1601,N_1696);
nand U1898 (N_1898,N_1790,N_1657);
or U1899 (N_1899,N_1793,N_1788);
nand U1900 (N_1900,N_1704,N_1663);
nand U1901 (N_1901,N_1635,N_1773);
or U1902 (N_1902,N_1725,N_1798);
or U1903 (N_1903,N_1650,N_1765);
or U1904 (N_1904,N_1651,N_1674);
and U1905 (N_1905,N_1721,N_1755);
nand U1906 (N_1906,N_1626,N_1695);
nor U1907 (N_1907,N_1693,N_1637);
nand U1908 (N_1908,N_1702,N_1776);
and U1909 (N_1909,N_1617,N_1720);
nor U1910 (N_1910,N_1710,N_1689);
nor U1911 (N_1911,N_1738,N_1695);
or U1912 (N_1912,N_1734,N_1751);
and U1913 (N_1913,N_1610,N_1614);
nand U1914 (N_1914,N_1694,N_1685);
nand U1915 (N_1915,N_1672,N_1610);
or U1916 (N_1916,N_1635,N_1654);
and U1917 (N_1917,N_1776,N_1650);
and U1918 (N_1918,N_1715,N_1780);
nor U1919 (N_1919,N_1704,N_1645);
and U1920 (N_1920,N_1736,N_1700);
and U1921 (N_1921,N_1656,N_1658);
nor U1922 (N_1922,N_1747,N_1704);
xnor U1923 (N_1923,N_1623,N_1726);
nor U1924 (N_1924,N_1618,N_1773);
xnor U1925 (N_1925,N_1767,N_1749);
nor U1926 (N_1926,N_1691,N_1641);
and U1927 (N_1927,N_1646,N_1782);
and U1928 (N_1928,N_1611,N_1733);
or U1929 (N_1929,N_1633,N_1793);
nand U1930 (N_1930,N_1752,N_1775);
or U1931 (N_1931,N_1609,N_1719);
nor U1932 (N_1932,N_1629,N_1796);
and U1933 (N_1933,N_1758,N_1655);
and U1934 (N_1934,N_1662,N_1734);
and U1935 (N_1935,N_1708,N_1676);
and U1936 (N_1936,N_1648,N_1774);
nor U1937 (N_1937,N_1778,N_1646);
or U1938 (N_1938,N_1738,N_1735);
or U1939 (N_1939,N_1627,N_1642);
nand U1940 (N_1940,N_1797,N_1697);
nand U1941 (N_1941,N_1604,N_1677);
or U1942 (N_1942,N_1671,N_1636);
nor U1943 (N_1943,N_1798,N_1742);
and U1944 (N_1944,N_1700,N_1651);
nor U1945 (N_1945,N_1606,N_1739);
nand U1946 (N_1946,N_1652,N_1618);
nand U1947 (N_1947,N_1728,N_1744);
or U1948 (N_1948,N_1625,N_1779);
nor U1949 (N_1949,N_1795,N_1748);
and U1950 (N_1950,N_1606,N_1717);
nand U1951 (N_1951,N_1747,N_1612);
nand U1952 (N_1952,N_1757,N_1764);
or U1953 (N_1953,N_1691,N_1740);
or U1954 (N_1954,N_1667,N_1798);
nand U1955 (N_1955,N_1732,N_1655);
or U1956 (N_1956,N_1779,N_1602);
nand U1957 (N_1957,N_1727,N_1669);
nand U1958 (N_1958,N_1635,N_1797);
xor U1959 (N_1959,N_1612,N_1780);
or U1960 (N_1960,N_1638,N_1666);
nand U1961 (N_1961,N_1687,N_1633);
nand U1962 (N_1962,N_1739,N_1633);
or U1963 (N_1963,N_1695,N_1629);
or U1964 (N_1964,N_1603,N_1720);
and U1965 (N_1965,N_1632,N_1754);
nand U1966 (N_1966,N_1725,N_1740);
nand U1967 (N_1967,N_1643,N_1776);
and U1968 (N_1968,N_1773,N_1711);
nand U1969 (N_1969,N_1648,N_1750);
nor U1970 (N_1970,N_1604,N_1636);
and U1971 (N_1971,N_1768,N_1690);
nand U1972 (N_1972,N_1655,N_1603);
and U1973 (N_1973,N_1624,N_1765);
nor U1974 (N_1974,N_1752,N_1687);
xor U1975 (N_1975,N_1612,N_1649);
nand U1976 (N_1976,N_1793,N_1680);
nor U1977 (N_1977,N_1708,N_1668);
nand U1978 (N_1978,N_1686,N_1627);
xor U1979 (N_1979,N_1600,N_1683);
xor U1980 (N_1980,N_1613,N_1679);
nor U1981 (N_1981,N_1763,N_1769);
nor U1982 (N_1982,N_1604,N_1719);
or U1983 (N_1983,N_1625,N_1642);
or U1984 (N_1984,N_1664,N_1761);
xor U1985 (N_1985,N_1687,N_1629);
nor U1986 (N_1986,N_1780,N_1602);
or U1987 (N_1987,N_1637,N_1764);
nand U1988 (N_1988,N_1766,N_1760);
nor U1989 (N_1989,N_1650,N_1761);
or U1990 (N_1990,N_1781,N_1709);
or U1991 (N_1991,N_1672,N_1775);
xnor U1992 (N_1992,N_1654,N_1796);
nand U1993 (N_1993,N_1680,N_1724);
nand U1994 (N_1994,N_1694,N_1678);
nor U1995 (N_1995,N_1706,N_1633);
nor U1996 (N_1996,N_1669,N_1742);
nand U1997 (N_1997,N_1713,N_1698);
nor U1998 (N_1998,N_1688,N_1796);
or U1999 (N_1999,N_1766,N_1660);
and U2000 (N_2000,N_1822,N_1951);
and U2001 (N_2001,N_1840,N_1863);
nor U2002 (N_2002,N_1967,N_1828);
and U2003 (N_2003,N_1804,N_1809);
nand U2004 (N_2004,N_1979,N_1976);
nand U2005 (N_2005,N_1986,N_1875);
nand U2006 (N_2006,N_1850,N_1854);
nor U2007 (N_2007,N_1958,N_1920);
and U2008 (N_2008,N_1930,N_1907);
nand U2009 (N_2009,N_1855,N_1818);
nor U2010 (N_2010,N_1945,N_1836);
nor U2011 (N_2011,N_1996,N_1857);
or U2012 (N_2012,N_1905,N_1862);
or U2013 (N_2013,N_1974,N_1977);
or U2014 (N_2014,N_1948,N_1807);
xnor U2015 (N_2015,N_1995,N_1894);
nor U2016 (N_2016,N_1903,N_1889);
or U2017 (N_2017,N_1975,N_1802);
or U2018 (N_2018,N_1832,N_1801);
nor U2019 (N_2019,N_1871,N_1960);
nor U2020 (N_2020,N_1914,N_1987);
xor U2021 (N_2021,N_1901,N_1962);
xnor U2022 (N_2022,N_1963,N_1815);
nor U2023 (N_2023,N_1848,N_1806);
nor U2024 (N_2024,N_1814,N_1938);
nand U2025 (N_2025,N_1965,N_1800);
nor U2026 (N_2026,N_1844,N_1819);
or U2027 (N_2027,N_1829,N_1919);
or U2028 (N_2028,N_1912,N_1821);
nand U2029 (N_2029,N_1851,N_1849);
nand U2030 (N_2030,N_1830,N_1865);
nand U2031 (N_2031,N_1913,N_1908);
nand U2032 (N_2032,N_1954,N_1937);
or U2033 (N_2033,N_1994,N_1939);
nand U2034 (N_2034,N_1956,N_1825);
or U2035 (N_2035,N_1856,N_1918);
nand U2036 (N_2036,N_1959,N_1992);
nor U2037 (N_2037,N_1893,N_1877);
nand U2038 (N_2038,N_1989,N_1916);
nor U2039 (N_2039,N_1973,N_1860);
or U2040 (N_2040,N_1833,N_1980);
nor U2041 (N_2041,N_1805,N_1926);
nor U2042 (N_2042,N_1872,N_1892);
or U2043 (N_2043,N_1928,N_1941);
and U2044 (N_2044,N_1891,N_1887);
xnor U2045 (N_2045,N_1881,N_1924);
nor U2046 (N_2046,N_1895,N_1882);
xnor U2047 (N_2047,N_1886,N_1846);
nand U2048 (N_2048,N_1988,N_1985);
nand U2049 (N_2049,N_1803,N_1869);
or U2050 (N_2050,N_1972,N_1834);
nand U2051 (N_2051,N_1880,N_1983);
or U2052 (N_2052,N_1904,N_1861);
xnor U2053 (N_2053,N_1971,N_1837);
nor U2054 (N_2054,N_1969,N_1816);
or U2055 (N_2055,N_1839,N_1957);
nor U2056 (N_2056,N_1981,N_1993);
nand U2057 (N_2057,N_1847,N_1921);
nand U2058 (N_2058,N_1978,N_1858);
and U2059 (N_2059,N_1922,N_1842);
or U2060 (N_2060,N_1934,N_1812);
or U2061 (N_2061,N_1852,N_1823);
or U2062 (N_2062,N_1838,N_1883);
and U2063 (N_2063,N_1824,N_1884);
or U2064 (N_2064,N_1929,N_1933);
xor U2065 (N_2065,N_1931,N_1935);
xor U2066 (N_2066,N_1911,N_1946);
nand U2067 (N_2067,N_1947,N_1866);
nand U2068 (N_2068,N_1990,N_1902);
or U2069 (N_2069,N_1864,N_1888);
xnor U2070 (N_2070,N_1917,N_1909);
or U2071 (N_2071,N_1898,N_1870);
nand U2072 (N_2072,N_1997,N_1874);
xnor U2073 (N_2073,N_1953,N_1915);
nand U2074 (N_2074,N_1900,N_1876);
and U2075 (N_2075,N_1923,N_1817);
and U2076 (N_2076,N_1925,N_1897);
nand U2077 (N_2077,N_1955,N_1991);
or U2078 (N_2078,N_1813,N_1999);
nor U2079 (N_2079,N_1932,N_1873);
or U2080 (N_2080,N_1982,N_1984);
or U2081 (N_2081,N_1968,N_1936);
and U2082 (N_2082,N_1906,N_1961);
xor U2083 (N_2083,N_1808,N_1868);
and U2084 (N_2084,N_1899,N_1879);
nand U2085 (N_2085,N_1843,N_1827);
or U2086 (N_2086,N_1966,N_1885);
xnor U2087 (N_2087,N_1896,N_1943);
nand U2088 (N_2088,N_1970,N_1998);
nand U2089 (N_2089,N_1944,N_1853);
and U2090 (N_2090,N_1952,N_1845);
or U2091 (N_2091,N_1811,N_1964);
nor U2092 (N_2092,N_1910,N_1867);
nor U2093 (N_2093,N_1927,N_1950);
xnor U2094 (N_2094,N_1820,N_1835);
nand U2095 (N_2095,N_1810,N_1890);
and U2096 (N_2096,N_1841,N_1831);
and U2097 (N_2097,N_1878,N_1942);
nor U2098 (N_2098,N_1949,N_1826);
or U2099 (N_2099,N_1859,N_1940);
or U2100 (N_2100,N_1878,N_1968);
nand U2101 (N_2101,N_1929,N_1908);
or U2102 (N_2102,N_1898,N_1979);
nor U2103 (N_2103,N_1995,N_1878);
xor U2104 (N_2104,N_1986,N_1974);
or U2105 (N_2105,N_1889,N_1855);
xor U2106 (N_2106,N_1846,N_1858);
or U2107 (N_2107,N_1959,N_1982);
nor U2108 (N_2108,N_1995,N_1970);
nor U2109 (N_2109,N_1826,N_1932);
nand U2110 (N_2110,N_1955,N_1939);
xor U2111 (N_2111,N_1912,N_1835);
xor U2112 (N_2112,N_1963,N_1949);
or U2113 (N_2113,N_1986,N_1804);
and U2114 (N_2114,N_1873,N_1874);
or U2115 (N_2115,N_1936,N_1873);
xor U2116 (N_2116,N_1857,N_1964);
nand U2117 (N_2117,N_1856,N_1808);
nor U2118 (N_2118,N_1940,N_1982);
xor U2119 (N_2119,N_1944,N_1907);
or U2120 (N_2120,N_1993,N_1961);
and U2121 (N_2121,N_1806,N_1800);
or U2122 (N_2122,N_1897,N_1961);
or U2123 (N_2123,N_1870,N_1858);
nand U2124 (N_2124,N_1840,N_1929);
or U2125 (N_2125,N_1955,N_1822);
nor U2126 (N_2126,N_1986,N_1939);
and U2127 (N_2127,N_1816,N_1819);
nand U2128 (N_2128,N_1930,N_1857);
xor U2129 (N_2129,N_1917,N_1925);
nand U2130 (N_2130,N_1940,N_1975);
nor U2131 (N_2131,N_1969,N_1940);
and U2132 (N_2132,N_1837,N_1832);
and U2133 (N_2133,N_1890,N_1909);
nand U2134 (N_2134,N_1826,N_1911);
xor U2135 (N_2135,N_1965,N_1967);
and U2136 (N_2136,N_1914,N_1850);
or U2137 (N_2137,N_1814,N_1874);
xnor U2138 (N_2138,N_1922,N_1999);
nand U2139 (N_2139,N_1996,N_1803);
xor U2140 (N_2140,N_1954,N_1862);
or U2141 (N_2141,N_1960,N_1952);
nand U2142 (N_2142,N_1815,N_1875);
nand U2143 (N_2143,N_1808,N_1981);
nand U2144 (N_2144,N_1895,N_1819);
nor U2145 (N_2145,N_1830,N_1952);
or U2146 (N_2146,N_1904,N_1834);
and U2147 (N_2147,N_1811,N_1861);
nand U2148 (N_2148,N_1920,N_1911);
xor U2149 (N_2149,N_1825,N_1936);
nand U2150 (N_2150,N_1865,N_1940);
xor U2151 (N_2151,N_1870,N_1861);
or U2152 (N_2152,N_1938,N_1909);
and U2153 (N_2153,N_1981,N_1965);
or U2154 (N_2154,N_1827,N_1962);
nand U2155 (N_2155,N_1985,N_1924);
nor U2156 (N_2156,N_1827,N_1805);
nor U2157 (N_2157,N_1889,N_1827);
nand U2158 (N_2158,N_1922,N_1945);
xnor U2159 (N_2159,N_1926,N_1813);
nand U2160 (N_2160,N_1964,N_1941);
or U2161 (N_2161,N_1927,N_1870);
and U2162 (N_2162,N_1827,N_1954);
and U2163 (N_2163,N_1906,N_1837);
or U2164 (N_2164,N_1881,N_1956);
nand U2165 (N_2165,N_1986,N_1821);
nand U2166 (N_2166,N_1827,N_1882);
and U2167 (N_2167,N_1878,N_1836);
or U2168 (N_2168,N_1825,N_1937);
and U2169 (N_2169,N_1906,N_1894);
and U2170 (N_2170,N_1923,N_1994);
nor U2171 (N_2171,N_1969,N_1882);
and U2172 (N_2172,N_1919,N_1806);
xnor U2173 (N_2173,N_1800,N_1861);
and U2174 (N_2174,N_1836,N_1865);
nand U2175 (N_2175,N_1871,N_1915);
or U2176 (N_2176,N_1996,N_1938);
nand U2177 (N_2177,N_1800,N_1907);
or U2178 (N_2178,N_1911,N_1863);
nand U2179 (N_2179,N_1889,N_1823);
and U2180 (N_2180,N_1913,N_1849);
xnor U2181 (N_2181,N_1831,N_1994);
nand U2182 (N_2182,N_1824,N_1900);
nand U2183 (N_2183,N_1805,N_1806);
nor U2184 (N_2184,N_1905,N_1928);
and U2185 (N_2185,N_1844,N_1889);
and U2186 (N_2186,N_1822,N_1829);
or U2187 (N_2187,N_1906,N_1905);
and U2188 (N_2188,N_1958,N_1932);
nand U2189 (N_2189,N_1995,N_1842);
or U2190 (N_2190,N_1804,N_1852);
nor U2191 (N_2191,N_1874,N_1894);
xnor U2192 (N_2192,N_1898,N_1807);
nor U2193 (N_2193,N_1864,N_1839);
nor U2194 (N_2194,N_1872,N_1966);
and U2195 (N_2195,N_1837,N_1855);
and U2196 (N_2196,N_1863,N_1892);
and U2197 (N_2197,N_1835,N_1995);
nand U2198 (N_2198,N_1921,N_1901);
or U2199 (N_2199,N_1879,N_1821);
nand U2200 (N_2200,N_2172,N_2052);
nor U2201 (N_2201,N_2154,N_2046);
or U2202 (N_2202,N_2058,N_2074);
nor U2203 (N_2203,N_2160,N_2105);
or U2204 (N_2204,N_2121,N_2128);
nand U2205 (N_2205,N_2008,N_2125);
nor U2206 (N_2206,N_2187,N_2186);
nor U2207 (N_2207,N_2049,N_2112);
or U2208 (N_2208,N_2048,N_2053);
xor U2209 (N_2209,N_2155,N_2095);
or U2210 (N_2210,N_2163,N_2101);
and U2211 (N_2211,N_2098,N_2152);
nand U2212 (N_2212,N_2017,N_2004);
nand U2213 (N_2213,N_2142,N_2035);
nor U2214 (N_2214,N_2018,N_2060);
nor U2215 (N_2215,N_2119,N_2036);
xor U2216 (N_2216,N_2088,N_2159);
nand U2217 (N_2217,N_2113,N_2042);
nand U2218 (N_2218,N_2020,N_2059);
nand U2219 (N_2219,N_2100,N_2199);
nand U2220 (N_2220,N_2037,N_2136);
or U2221 (N_2221,N_2115,N_2151);
and U2222 (N_2222,N_2044,N_2065);
nand U2223 (N_2223,N_2179,N_2009);
and U2224 (N_2224,N_2024,N_2068);
and U2225 (N_2225,N_2080,N_2034);
and U2226 (N_2226,N_2056,N_2062);
or U2227 (N_2227,N_2064,N_2073);
and U2228 (N_2228,N_2176,N_2000);
or U2229 (N_2229,N_2093,N_2021);
and U2230 (N_2230,N_2012,N_2120);
nor U2231 (N_2231,N_2003,N_2149);
nor U2232 (N_2232,N_2026,N_2013);
nor U2233 (N_2233,N_2180,N_2097);
nand U2234 (N_2234,N_2072,N_2107);
and U2235 (N_2235,N_2178,N_2085);
nand U2236 (N_2236,N_2051,N_2092);
nand U2237 (N_2237,N_2019,N_2143);
or U2238 (N_2238,N_2185,N_2130);
nand U2239 (N_2239,N_2114,N_2027);
xor U2240 (N_2240,N_2116,N_2127);
nor U2241 (N_2241,N_2165,N_2045);
nand U2242 (N_2242,N_2040,N_2134);
nor U2243 (N_2243,N_2031,N_2108);
nand U2244 (N_2244,N_2129,N_2188);
nand U2245 (N_2245,N_2023,N_2123);
or U2246 (N_2246,N_2171,N_2099);
nor U2247 (N_2247,N_2041,N_2150);
or U2248 (N_2248,N_2096,N_2194);
nor U2249 (N_2249,N_2139,N_2190);
nor U2250 (N_2250,N_2167,N_2109);
nor U2251 (N_2251,N_2032,N_2077);
nor U2252 (N_2252,N_2066,N_2078);
or U2253 (N_2253,N_2137,N_2104);
and U2254 (N_2254,N_2182,N_2039);
or U2255 (N_2255,N_2195,N_2054);
and U2256 (N_2256,N_2089,N_2164);
nor U2257 (N_2257,N_2161,N_2166);
or U2258 (N_2258,N_2168,N_2030);
nor U2259 (N_2259,N_2087,N_2083);
xor U2260 (N_2260,N_2156,N_2086);
and U2261 (N_2261,N_2175,N_2090);
nor U2262 (N_2262,N_2010,N_2197);
nor U2263 (N_2263,N_2144,N_2135);
or U2264 (N_2264,N_2147,N_2082);
and U2265 (N_2265,N_2069,N_2061);
nor U2266 (N_2266,N_2001,N_2181);
and U2267 (N_2267,N_2091,N_2131);
nor U2268 (N_2268,N_2157,N_2140);
nand U2269 (N_2269,N_2084,N_2124);
nor U2270 (N_2270,N_2103,N_2015);
or U2271 (N_2271,N_2005,N_2141);
nand U2272 (N_2272,N_2192,N_2076);
and U2273 (N_2273,N_2148,N_2106);
and U2274 (N_2274,N_2153,N_2183);
and U2275 (N_2275,N_2133,N_2170);
or U2276 (N_2276,N_2173,N_2025);
nor U2277 (N_2277,N_2022,N_2029);
or U2278 (N_2278,N_2145,N_2158);
nor U2279 (N_2279,N_2193,N_2110);
or U2280 (N_2280,N_2043,N_2033);
and U2281 (N_2281,N_2007,N_2102);
and U2282 (N_2282,N_2014,N_2028);
nand U2283 (N_2283,N_2177,N_2075);
or U2284 (N_2284,N_2071,N_2122);
and U2285 (N_2285,N_2081,N_2079);
nor U2286 (N_2286,N_2011,N_2070);
or U2287 (N_2287,N_2050,N_2047);
or U2288 (N_2288,N_2189,N_2002);
xnor U2289 (N_2289,N_2055,N_2126);
and U2290 (N_2290,N_2016,N_2094);
and U2291 (N_2291,N_2174,N_2184);
and U2292 (N_2292,N_2196,N_2057);
or U2293 (N_2293,N_2146,N_2117);
nor U2294 (N_2294,N_2191,N_2198);
or U2295 (N_2295,N_2063,N_2138);
or U2296 (N_2296,N_2132,N_2111);
or U2297 (N_2297,N_2038,N_2162);
nor U2298 (N_2298,N_2169,N_2006);
nor U2299 (N_2299,N_2067,N_2118);
nand U2300 (N_2300,N_2105,N_2010);
xnor U2301 (N_2301,N_2192,N_2158);
nand U2302 (N_2302,N_2127,N_2081);
or U2303 (N_2303,N_2064,N_2163);
nand U2304 (N_2304,N_2190,N_2106);
and U2305 (N_2305,N_2190,N_2129);
nor U2306 (N_2306,N_2176,N_2081);
or U2307 (N_2307,N_2042,N_2080);
or U2308 (N_2308,N_2174,N_2164);
or U2309 (N_2309,N_2072,N_2014);
nor U2310 (N_2310,N_2177,N_2034);
and U2311 (N_2311,N_2167,N_2009);
nor U2312 (N_2312,N_2138,N_2126);
nor U2313 (N_2313,N_2052,N_2011);
and U2314 (N_2314,N_2187,N_2064);
nand U2315 (N_2315,N_2107,N_2102);
and U2316 (N_2316,N_2100,N_2172);
nand U2317 (N_2317,N_2010,N_2167);
nor U2318 (N_2318,N_2100,N_2003);
and U2319 (N_2319,N_2187,N_2053);
nand U2320 (N_2320,N_2141,N_2121);
and U2321 (N_2321,N_2070,N_2006);
nand U2322 (N_2322,N_2186,N_2084);
xnor U2323 (N_2323,N_2184,N_2086);
nor U2324 (N_2324,N_2034,N_2161);
and U2325 (N_2325,N_2103,N_2025);
xor U2326 (N_2326,N_2157,N_2162);
and U2327 (N_2327,N_2156,N_2035);
xor U2328 (N_2328,N_2099,N_2184);
nand U2329 (N_2329,N_2184,N_2071);
nand U2330 (N_2330,N_2121,N_2181);
or U2331 (N_2331,N_2010,N_2190);
or U2332 (N_2332,N_2024,N_2176);
and U2333 (N_2333,N_2152,N_2011);
nor U2334 (N_2334,N_2009,N_2047);
nor U2335 (N_2335,N_2100,N_2113);
and U2336 (N_2336,N_2155,N_2064);
nor U2337 (N_2337,N_2031,N_2053);
or U2338 (N_2338,N_2073,N_2137);
or U2339 (N_2339,N_2067,N_2193);
nor U2340 (N_2340,N_2059,N_2117);
nor U2341 (N_2341,N_2160,N_2097);
or U2342 (N_2342,N_2195,N_2125);
nand U2343 (N_2343,N_2153,N_2048);
nor U2344 (N_2344,N_2144,N_2031);
nor U2345 (N_2345,N_2042,N_2156);
and U2346 (N_2346,N_2188,N_2031);
or U2347 (N_2347,N_2073,N_2103);
nand U2348 (N_2348,N_2004,N_2108);
nand U2349 (N_2349,N_2113,N_2155);
and U2350 (N_2350,N_2187,N_2131);
and U2351 (N_2351,N_2099,N_2158);
nand U2352 (N_2352,N_2050,N_2014);
and U2353 (N_2353,N_2038,N_2023);
nand U2354 (N_2354,N_2055,N_2062);
and U2355 (N_2355,N_2021,N_2006);
nor U2356 (N_2356,N_2064,N_2170);
nand U2357 (N_2357,N_2165,N_2086);
and U2358 (N_2358,N_2151,N_2080);
xnor U2359 (N_2359,N_2148,N_2085);
or U2360 (N_2360,N_2058,N_2020);
and U2361 (N_2361,N_2006,N_2142);
xor U2362 (N_2362,N_2172,N_2110);
nor U2363 (N_2363,N_2007,N_2019);
and U2364 (N_2364,N_2189,N_2027);
nand U2365 (N_2365,N_2086,N_2149);
or U2366 (N_2366,N_2097,N_2183);
nor U2367 (N_2367,N_2022,N_2060);
nand U2368 (N_2368,N_2027,N_2132);
xor U2369 (N_2369,N_2097,N_2147);
xor U2370 (N_2370,N_2062,N_2084);
nor U2371 (N_2371,N_2071,N_2069);
and U2372 (N_2372,N_2152,N_2135);
nor U2373 (N_2373,N_2123,N_2097);
nand U2374 (N_2374,N_2165,N_2149);
and U2375 (N_2375,N_2096,N_2029);
nor U2376 (N_2376,N_2031,N_2128);
and U2377 (N_2377,N_2069,N_2199);
nand U2378 (N_2378,N_2092,N_2080);
nand U2379 (N_2379,N_2145,N_2096);
and U2380 (N_2380,N_2152,N_2048);
or U2381 (N_2381,N_2051,N_2193);
nand U2382 (N_2382,N_2168,N_2043);
or U2383 (N_2383,N_2168,N_2153);
or U2384 (N_2384,N_2060,N_2082);
nor U2385 (N_2385,N_2074,N_2171);
nor U2386 (N_2386,N_2029,N_2190);
xor U2387 (N_2387,N_2029,N_2164);
or U2388 (N_2388,N_2167,N_2133);
nand U2389 (N_2389,N_2126,N_2079);
or U2390 (N_2390,N_2036,N_2159);
nor U2391 (N_2391,N_2025,N_2033);
nand U2392 (N_2392,N_2001,N_2144);
nand U2393 (N_2393,N_2187,N_2070);
nand U2394 (N_2394,N_2058,N_2072);
and U2395 (N_2395,N_2103,N_2191);
or U2396 (N_2396,N_2164,N_2106);
and U2397 (N_2397,N_2176,N_2027);
nand U2398 (N_2398,N_2070,N_2164);
xor U2399 (N_2399,N_2167,N_2149);
or U2400 (N_2400,N_2352,N_2388);
nand U2401 (N_2401,N_2264,N_2303);
nand U2402 (N_2402,N_2355,N_2260);
and U2403 (N_2403,N_2381,N_2208);
nor U2404 (N_2404,N_2350,N_2202);
nand U2405 (N_2405,N_2266,N_2293);
xor U2406 (N_2406,N_2326,N_2257);
nor U2407 (N_2407,N_2325,N_2201);
nand U2408 (N_2408,N_2270,N_2313);
and U2409 (N_2409,N_2343,N_2216);
or U2410 (N_2410,N_2390,N_2254);
and U2411 (N_2411,N_2375,N_2327);
and U2412 (N_2412,N_2275,N_2247);
nor U2413 (N_2413,N_2203,N_2278);
or U2414 (N_2414,N_2320,N_2356);
and U2415 (N_2415,N_2259,N_2358);
nor U2416 (N_2416,N_2206,N_2217);
or U2417 (N_2417,N_2359,N_2287);
and U2418 (N_2418,N_2398,N_2305);
or U2419 (N_2419,N_2207,N_2237);
nand U2420 (N_2420,N_2339,N_2221);
xnor U2421 (N_2421,N_2240,N_2280);
and U2422 (N_2422,N_2276,N_2252);
or U2423 (N_2423,N_2291,N_2351);
xnor U2424 (N_2424,N_2328,N_2300);
nor U2425 (N_2425,N_2330,N_2226);
or U2426 (N_2426,N_2397,N_2304);
nand U2427 (N_2427,N_2379,N_2360);
nor U2428 (N_2428,N_2246,N_2384);
nor U2429 (N_2429,N_2363,N_2211);
and U2430 (N_2430,N_2210,N_2357);
nand U2431 (N_2431,N_2367,N_2277);
nand U2432 (N_2432,N_2376,N_2393);
and U2433 (N_2433,N_2310,N_2329);
and U2434 (N_2434,N_2315,N_2228);
nand U2435 (N_2435,N_2253,N_2336);
nand U2436 (N_2436,N_2340,N_2338);
nor U2437 (N_2437,N_2285,N_2213);
or U2438 (N_2438,N_2392,N_2324);
and U2439 (N_2439,N_2225,N_2235);
or U2440 (N_2440,N_2321,N_2238);
nor U2441 (N_2441,N_2265,N_2395);
and U2442 (N_2442,N_2364,N_2374);
nor U2443 (N_2443,N_2200,N_2289);
or U2444 (N_2444,N_2284,N_2349);
nand U2445 (N_2445,N_2382,N_2233);
or U2446 (N_2446,N_2241,N_2378);
xnor U2447 (N_2447,N_2319,N_2337);
or U2448 (N_2448,N_2295,N_2348);
nand U2449 (N_2449,N_2244,N_2236);
and U2450 (N_2450,N_2204,N_2281);
nand U2451 (N_2451,N_2368,N_2333);
nor U2452 (N_2452,N_2250,N_2383);
nor U2453 (N_2453,N_2262,N_2373);
nor U2454 (N_2454,N_2209,N_2279);
and U2455 (N_2455,N_2298,N_2361);
and U2456 (N_2456,N_2261,N_2269);
xor U2457 (N_2457,N_2248,N_2387);
nor U2458 (N_2458,N_2322,N_2258);
or U2459 (N_2459,N_2370,N_2286);
or U2460 (N_2460,N_2239,N_2385);
or U2461 (N_2461,N_2371,N_2314);
nand U2462 (N_2462,N_2288,N_2222);
nor U2463 (N_2463,N_2341,N_2218);
nand U2464 (N_2464,N_2317,N_2212);
or U2465 (N_2465,N_2292,N_2214);
and U2466 (N_2466,N_2342,N_2308);
nand U2467 (N_2467,N_2227,N_2345);
xnor U2468 (N_2468,N_2273,N_2294);
and U2469 (N_2469,N_2231,N_2334);
or U2470 (N_2470,N_2311,N_2309);
xor U2471 (N_2471,N_2386,N_2224);
nand U2472 (N_2472,N_2312,N_2223);
nor U2473 (N_2473,N_2274,N_2307);
and U2474 (N_2474,N_2263,N_2220);
and U2475 (N_2475,N_2283,N_2272);
or U2476 (N_2476,N_2380,N_2399);
and U2477 (N_2477,N_2369,N_2302);
or U2478 (N_2478,N_2249,N_2296);
and U2479 (N_2479,N_2344,N_2396);
and U2480 (N_2480,N_2323,N_2256);
nor U2481 (N_2481,N_2271,N_2299);
xnor U2482 (N_2482,N_2372,N_2316);
nand U2483 (N_2483,N_2267,N_2229);
nor U2484 (N_2484,N_2335,N_2251);
xnor U2485 (N_2485,N_2282,N_2354);
and U2486 (N_2486,N_2205,N_2243);
nor U2487 (N_2487,N_2245,N_2389);
nor U2488 (N_2488,N_2230,N_2290);
nor U2489 (N_2489,N_2391,N_2366);
or U2490 (N_2490,N_2234,N_2377);
nand U2491 (N_2491,N_2306,N_2232);
or U2492 (N_2492,N_2365,N_2353);
and U2493 (N_2493,N_2347,N_2332);
nand U2494 (N_2494,N_2219,N_2242);
nor U2495 (N_2495,N_2394,N_2318);
nor U2496 (N_2496,N_2268,N_2331);
or U2497 (N_2497,N_2301,N_2362);
nand U2498 (N_2498,N_2255,N_2215);
or U2499 (N_2499,N_2297,N_2346);
and U2500 (N_2500,N_2316,N_2377);
xnor U2501 (N_2501,N_2293,N_2274);
and U2502 (N_2502,N_2305,N_2219);
nand U2503 (N_2503,N_2248,N_2234);
nor U2504 (N_2504,N_2259,N_2340);
or U2505 (N_2505,N_2362,N_2212);
and U2506 (N_2506,N_2306,N_2275);
nand U2507 (N_2507,N_2320,N_2258);
nand U2508 (N_2508,N_2284,N_2316);
nand U2509 (N_2509,N_2317,N_2238);
nor U2510 (N_2510,N_2320,N_2303);
and U2511 (N_2511,N_2276,N_2381);
and U2512 (N_2512,N_2355,N_2338);
xnor U2513 (N_2513,N_2376,N_2347);
and U2514 (N_2514,N_2334,N_2322);
nor U2515 (N_2515,N_2204,N_2369);
nor U2516 (N_2516,N_2385,N_2285);
and U2517 (N_2517,N_2268,N_2240);
or U2518 (N_2518,N_2364,N_2259);
nor U2519 (N_2519,N_2202,N_2234);
or U2520 (N_2520,N_2268,N_2297);
nor U2521 (N_2521,N_2323,N_2301);
nor U2522 (N_2522,N_2227,N_2330);
nand U2523 (N_2523,N_2348,N_2271);
nand U2524 (N_2524,N_2287,N_2300);
nor U2525 (N_2525,N_2381,N_2233);
nand U2526 (N_2526,N_2384,N_2371);
or U2527 (N_2527,N_2356,N_2331);
nor U2528 (N_2528,N_2260,N_2306);
nand U2529 (N_2529,N_2299,N_2376);
and U2530 (N_2530,N_2248,N_2349);
nand U2531 (N_2531,N_2202,N_2227);
nor U2532 (N_2532,N_2298,N_2397);
or U2533 (N_2533,N_2222,N_2342);
or U2534 (N_2534,N_2232,N_2298);
xor U2535 (N_2535,N_2398,N_2377);
nor U2536 (N_2536,N_2345,N_2224);
or U2537 (N_2537,N_2303,N_2348);
nand U2538 (N_2538,N_2368,N_2326);
xnor U2539 (N_2539,N_2311,N_2252);
and U2540 (N_2540,N_2293,N_2330);
nor U2541 (N_2541,N_2303,N_2209);
or U2542 (N_2542,N_2315,N_2212);
nand U2543 (N_2543,N_2293,N_2259);
xnor U2544 (N_2544,N_2357,N_2355);
nand U2545 (N_2545,N_2302,N_2286);
nor U2546 (N_2546,N_2365,N_2241);
and U2547 (N_2547,N_2239,N_2246);
xnor U2548 (N_2548,N_2250,N_2265);
nor U2549 (N_2549,N_2297,N_2323);
and U2550 (N_2550,N_2306,N_2383);
or U2551 (N_2551,N_2293,N_2378);
nor U2552 (N_2552,N_2395,N_2235);
nor U2553 (N_2553,N_2284,N_2226);
and U2554 (N_2554,N_2209,N_2339);
nand U2555 (N_2555,N_2312,N_2365);
or U2556 (N_2556,N_2377,N_2347);
or U2557 (N_2557,N_2364,N_2340);
nor U2558 (N_2558,N_2295,N_2212);
or U2559 (N_2559,N_2321,N_2333);
and U2560 (N_2560,N_2202,N_2284);
and U2561 (N_2561,N_2328,N_2237);
and U2562 (N_2562,N_2368,N_2218);
nor U2563 (N_2563,N_2247,N_2375);
nand U2564 (N_2564,N_2325,N_2209);
nand U2565 (N_2565,N_2258,N_2372);
nand U2566 (N_2566,N_2260,N_2284);
nand U2567 (N_2567,N_2397,N_2305);
nor U2568 (N_2568,N_2243,N_2374);
and U2569 (N_2569,N_2220,N_2396);
nand U2570 (N_2570,N_2279,N_2281);
xnor U2571 (N_2571,N_2317,N_2314);
or U2572 (N_2572,N_2334,N_2227);
xor U2573 (N_2573,N_2334,N_2271);
xnor U2574 (N_2574,N_2238,N_2326);
nor U2575 (N_2575,N_2259,N_2271);
and U2576 (N_2576,N_2364,N_2215);
nand U2577 (N_2577,N_2376,N_2398);
or U2578 (N_2578,N_2382,N_2399);
nor U2579 (N_2579,N_2220,N_2207);
nor U2580 (N_2580,N_2335,N_2327);
or U2581 (N_2581,N_2353,N_2264);
xnor U2582 (N_2582,N_2286,N_2352);
and U2583 (N_2583,N_2261,N_2380);
or U2584 (N_2584,N_2355,N_2283);
nor U2585 (N_2585,N_2240,N_2266);
or U2586 (N_2586,N_2301,N_2244);
and U2587 (N_2587,N_2394,N_2355);
nor U2588 (N_2588,N_2306,N_2218);
nor U2589 (N_2589,N_2327,N_2369);
nor U2590 (N_2590,N_2214,N_2237);
and U2591 (N_2591,N_2275,N_2323);
xor U2592 (N_2592,N_2255,N_2337);
and U2593 (N_2593,N_2250,N_2330);
and U2594 (N_2594,N_2283,N_2375);
nor U2595 (N_2595,N_2215,N_2377);
nor U2596 (N_2596,N_2352,N_2350);
and U2597 (N_2597,N_2203,N_2225);
xnor U2598 (N_2598,N_2369,N_2386);
nor U2599 (N_2599,N_2248,N_2307);
and U2600 (N_2600,N_2486,N_2506);
nand U2601 (N_2601,N_2537,N_2505);
or U2602 (N_2602,N_2508,N_2568);
nand U2603 (N_2603,N_2498,N_2532);
or U2604 (N_2604,N_2494,N_2533);
nor U2605 (N_2605,N_2493,N_2558);
and U2606 (N_2606,N_2567,N_2466);
and U2607 (N_2607,N_2473,N_2502);
and U2608 (N_2608,N_2546,N_2513);
or U2609 (N_2609,N_2481,N_2531);
and U2610 (N_2610,N_2431,N_2455);
nand U2611 (N_2611,N_2402,N_2582);
or U2612 (N_2612,N_2422,N_2413);
and U2613 (N_2613,N_2564,N_2515);
or U2614 (N_2614,N_2523,N_2427);
or U2615 (N_2615,N_2459,N_2565);
or U2616 (N_2616,N_2511,N_2593);
nand U2617 (N_2617,N_2577,N_2530);
or U2618 (N_2618,N_2425,N_2501);
nand U2619 (N_2619,N_2550,N_2424);
and U2620 (N_2620,N_2405,N_2461);
or U2621 (N_2621,N_2433,N_2518);
nand U2622 (N_2622,N_2599,N_2578);
nand U2623 (N_2623,N_2416,N_2432);
and U2624 (N_2624,N_2529,N_2591);
nor U2625 (N_2625,N_2544,N_2426);
nor U2626 (N_2626,N_2576,N_2587);
xor U2627 (N_2627,N_2504,N_2517);
or U2628 (N_2628,N_2509,N_2480);
xor U2629 (N_2629,N_2476,N_2468);
nor U2630 (N_2630,N_2454,N_2419);
nand U2631 (N_2631,N_2542,N_2430);
or U2632 (N_2632,N_2421,N_2453);
and U2633 (N_2633,N_2445,N_2474);
nand U2634 (N_2634,N_2470,N_2477);
or U2635 (N_2635,N_2536,N_2446);
xnor U2636 (N_2636,N_2524,N_2574);
nand U2637 (N_2637,N_2525,N_2566);
or U2638 (N_2638,N_2541,N_2503);
or U2639 (N_2639,N_2436,N_2545);
nor U2640 (N_2640,N_2540,N_2451);
and U2641 (N_2641,N_2572,N_2490);
nor U2642 (N_2642,N_2527,N_2557);
nand U2643 (N_2643,N_2435,N_2594);
nor U2644 (N_2644,N_2534,N_2483);
nor U2645 (N_2645,N_2596,N_2448);
nand U2646 (N_2646,N_2495,N_2479);
xor U2647 (N_2647,N_2588,N_2584);
or U2648 (N_2648,N_2450,N_2583);
nand U2649 (N_2649,N_2528,N_2561);
nand U2650 (N_2650,N_2553,N_2575);
and U2651 (N_2651,N_2428,N_2520);
or U2652 (N_2652,N_2535,N_2485);
nand U2653 (N_2653,N_2581,N_2595);
nor U2654 (N_2654,N_2547,N_2560);
and U2655 (N_2655,N_2403,N_2487);
and U2656 (N_2656,N_2482,N_2437);
or U2657 (N_2657,N_2423,N_2438);
and U2658 (N_2658,N_2496,N_2463);
nand U2659 (N_2659,N_2456,N_2439);
xor U2660 (N_2660,N_2514,N_2415);
xnor U2661 (N_2661,N_2548,N_2400);
and U2662 (N_2662,N_2447,N_2491);
and U2663 (N_2663,N_2510,N_2590);
xnor U2664 (N_2664,N_2406,N_2418);
or U2665 (N_2665,N_2579,N_2420);
or U2666 (N_2666,N_2440,N_2571);
xnor U2667 (N_2667,N_2460,N_2462);
nor U2668 (N_2668,N_2526,N_2555);
nand U2669 (N_2669,N_2484,N_2589);
and U2670 (N_2670,N_2443,N_2556);
xnor U2671 (N_2671,N_2489,N_2441);
and U2672 (N_2672,N_2580,N_2408);
xor U2673 (N_2673,N_2586,N_2497);
nand U2674 (N_2674,N_2411,N_2507);
and U2675 (N_2675,N_2598,N_2442);
or U2676 (N_2676,N_2457,N_2407);
xor U2677 (N_2677,N_2538,N_2414);
or U2678 (N_2678,N_2562,N_2554);
nand U2679 (N_2679,N_2409,N_2452);
nand U2680 (N_2680,N_2478,N_2472);
or U2681 (N_2681,N_2551,N_2475);
nor U2682 (N_2682,N_2492,N_2410);
xor U2683 (N_2683,N_2429,N_2521);
nand U2684 (N_2684,N_2467,N_2585);
nor U2685 (N_2685,N_2464,N_2543);
and U2686 (N_2686,N_2499,N_2401);
and U2687 (N_2687,N_2549,N_2465);
nor U2688 (N_2688,N_2539,N_2488);
or U2689 (N_2689,N_2471,N_2569);
nor U2690 (N_2690,N_2519,N_2469);
xnor U2691 (N_2691,N_2434,N_2592);
nand U2692 (N_2692,N_2573,N_2444);
nor U2693 (N_2693,N_2570,N_2559);
xnor U2694 (N_2694,N_2522,N_2500);
xnor U2695 (N_2695,N_2512,N_2412);
and U2696 (N_2696,N_2417,N_2449);
nor U2697 (N_2697,N_2516,N_2458);
nor U2698 (N_2698,N_2563,N_2552);
and U2699 (N_2699,N_2597,N_2404);
xor U2700 (N_2700,N_2505,N_2577);
and U2701 (N_2701,N_2575,N_2479);
nor U2702 (N_2702,N_2578,N_2410);
or U2703 (N_2703,N_2594,N_2496);
nor U2704 (N_2704,N_2406,N_2467);
nor U2705 (N_2705,N_2573,N_2536);
and U2706 (N_2706,N_2562,N_2445);
or U2707 (N_2707,N_2551,N_2490);
nor U2708 (N_2708,N_2542,N_2565);
or U2709 (N_2709,N_2570,N_2590);
xor U2710 (N_2710,N_2545,N_2520);
and U2711 (N_2711,N_2441,N_2572);
nor U2712 (N_2712,N_2498,N_2500);
nor U2713 (N_2713,N_2516,N_2555);
nor U2714 (N_2714,N_2485,N_2532);
nor U2715 (N_2715,N_2459,N_2463);
nor U2716 (N_2716,N_2426,N_2532);
nor U2717 (N_2717,N_2562,N_2433);
or U2718 (N_2718,N_2556,N_2417);
nor U2719 (N_2719,N_2490,N_2578);
and U2720 (N_2720,N_2596,N_2524);
or U2721 (N_2721,N_2599,N_2515);
xor U2722 (N_2722,N_2459,N_2556);
xnor U2723 (N_2723,N_2549,N_2486);
nor U2724 (N_2724,N_2586,N_2568);
nand U2725 (N_2725,N_2551,N_2592);
nand U2726 (N_2726,N_2473,N_2427);
nand U2727 (N_2727,N_2497,N_2440);
and U2728 (N_2728,N_2552,N_2500);
nand U2729 (N_2729,N_2529,N_2432);
and U2730 (N_2730,N_2553,N_2571);
and U2731 (N_2731,N_2519,N_2582);
nand U2732 (N_2732,N_2426,N_2562);
or U2733 (N_2733,N_2403,N_2560);
nor U2734 (N_2734,N_2557,N_2439);
or U2735 (N_2735,N_2419,N_2575);
nand U2736 (N_2736,N_2471,N_2593);
or U2737 (N_2737,N_2507,N_2522);
nor U2738 (N_2738,N_2532,N_2548);
and U2739 (N_2739,N_2580,N_2572);
and U2740 (N_2740,N_2414,N_2555);
nor U2741 (N_2741,N_2478,N_2509);
and U2742 (N_2742,N_2471,N_2488);
and U2743 (N_2743,N_2468,N_2543);
nand U2744 (N_2744,N_2429,N_2571);
nand U2745 (N_2745,N_2432,N_2541);
and U2746 (N_2746,N_2438,N_2596);
nor U2747 (N_2747,N_2497,N_2487);
nand U2748 (N_2748,N_2456,N_2519);
nor U2749 (N_2749,N_2530,N_2506);
and U2750 (N_2750,N_2556,N_2500);
nand U2751 (N_2751,N_2487,N_2588);
or U2752 (N_2752,N_2459,N_2542);
xnor U2753 (N_2753,N_2429,N_2480);
nand U2754 (N_2754,N_2524,N_2404);
nand U2755 (N_2755,N_2523,N_2479);
or U2756 (N_2756,N_2558,N_2504);
and U2757 (N_2757,N_2405,N_2482);
nor U2758 (N_2758,N_2533,N_2404);
or U2759 (N_2759,N_2405,N_2411);
nor U2760 (N_2760,N_2400,N_2433);
nand U2761 (N_2761,N_2594,N_2555);
nor U2762 (N_2762,N_2558,N_2521);
nor U2763 (N_2763,N_2594,N_2445);
or U2764 (N_2764,N_2502,N_2438);
nor U2765 (N_2765,N_2496,N_2486);
and U2766 (N_2766,N_2493,N_2454);
xnor U2767 (N_2767,N_2494,N_2496);
and U2768 (N_2768,N_2468,N_2498);
and U2769 (N_2769,N_2518,N_2404);
and U2770 (N_2770,N_2417,N_2472);
or U2771 (N_2771,N_2573,N_2492);
nor U2772 (N_2772,N_2469,N_2557);
nor U2773 (N_2773,N_2599,N_2577);
and U2774 (N_2774,N_2592,N_2407);
xor U2775 (N_2775,N_2493,N_2584);
nor U2776 (N_2776,N_2568,N_2419);
and U2777 (N_2777,N_2431,N_2457);
or U2778 (N_2778,N_2451,N_2504);
and U2779 (N_2779,N_2496,N_2512);
nand U2780 (N_2780,N_2400,N_2562);
xnor U2781 (N_2781,N_2446,N_2564);
nor U2782 (N_2782,N_2478,N_2452);
nand U2783 (N_2783,N_2569,N_2453);
or U2784 (N_2784,N_2422,N_2523);
or U2785 (N_2785,N_2430,N_2437);
or U2786 (N_2786,N_2526,N_2491);
nor U2787 (N_2787,N_2482,N_2473);
and U2788 (N_2788,N_2533,N_2408);
and U2789 (N_2789,N_2469,N_2410);
and U2790 (N_2790,N_2478,N_2532);
nor U2791 (N_2791,N_2552,N_2549);
or U2792 (N_2792,N_2451,N_2520);
nor U2793 (N_2793,N_2595,N_2538);
xor U2794 (N_2794,N_2419,N_2468);
or U2795 (N_2795,N_2466,N_2571);
and U2796 (N_2796,N_2575,N_2443);
nand U2797 (N_2797,N_2440,N_2574);
nor U2798 (N_2798,N_2448,N_2432);
or U2799 (N_2799,N_2588,N_2590);
xor U2800 (N_2800,N_2617,N_2624);
nand U2801 (N_2801,N_2766,N_2775);
xor U2802 (N_2802,N_2735,N_2725);
nor U2803 (N_2803,N_2686,N_2785);
nand U2804 (N_2804,N_2791,N_2759);
nand U2805 (N_2805,N_2777,N_2632);
or U2806 (N_2806,N_2622,N_2752);
or U2807 (N_2807,N_2690,N_2607);
or U2808 (N_2808,N_2745,N_2664);
nand U2809 (N_2809,N_2732,N_2693);
xor U2810 (N_2810,N_2730,N_2653);
or U2811 (N_2811,N_2659,N_2712);
nor U2812 (N_2812,N_2729,N_2675);
nand U2813 (N_2813,N_2701,N_2610);
and U2814 (N_2814,N_2741,N_2630);
and U2815 (N_2815,N_2756,N_2644);
nand U2816 (N_2816,N_2788,N_2746);
xor U2817 (N_2817,N_2660,N_2736);
and U2818 (N_2818,N_2799,N_2709);
nand U2819 (N_2819,N_2606,N_2683);
nand U2820 (N_2820,N_2749,N_2681);
or U2821 (N_2821,N_2688,N_2600);
nor U2822 (N_2822,N_2718,N_2768);
nor U2823 (N_2823,N_2760,N_2792);
nand U2824 (N_2824,N_2774,N_2783);
or U2825 (N_2825,N_2757,N_2793);
and U2826 (N_2826,N_2704,N_2784);
nor U2827 (N_2827,N_2685,N_2639);
or U2828 (N_2828,N_2739,N_2773);
xor U2829 (N_2829,N_2671,N_2682);
xnor U2830 (N_2830,N_2765,N_2723);
and U2831 (N_2831,N_2790,N_2636);
nand U2832 (N_2832,N_2738,N_2615);
nor U2833 (N_2833,N_2669,N_2798);
and U2834 (N_2834,N_2770,N_2706);
nor U2835 (N_2835,N_2654,N_2710);
and U2836 (N_2836,N_2795,N_2692);
nand U2837 (N_2837,N_2623,N_2713);
nand U2838 (N_2838,N_2769,N_2734);
or U2839 (N_2839,N_2767,N_2680);
nor U2840 (N_2840,N_2626,N_2667);
and U2841 (N_2841,N_2646,N_2689);
nor U2842 (N_2842,N_2780,N_2611);
xnor U2843 (N_2843,N_2789,N_2628);
and U2844 (N_2844,N_2715,N_2740);
and U2845 (N_2845,N_2695,N_2668);
and U2846 (N_2846,N_2676,N_2649);
or U2847 (N_2847,N_2678,N_2707);
nor U2848 (N_2848,N_2641,N_2684);
xor U2849 (N_2849,N_2743,N_2763);
nor U2850 (N_2850,N_2724,N_2609);
nand U2851 (N_2851,N_2705,N_2674);
and U2852 (N_2852,N_2782,N_2612);
nor U2853 (N_2853,N_2634,N_2754);
and U2854 (N_2854,N_2702,N_2666);
and U2855 (N_2855,N_2778,N_2751);
nor U2856 (N_2856,N_2779,N_2605);
nor U2857 (N_2857,N_2733,N_2656);
xor U2858 (N_2858,N_2651,N_2744);
nand U2859 (N_2859,N_2670,N_2629);
and U2860 (N_2860,N_2771,N_2647);
and U2861 (N_2861,N_2662,N_2711);
nand U2862 (N_2862,N_2677,N_2665);
and U2863 (N_2863,N_2750,N_2691);
and U2864 (N_2864,N_2726,N_2764);
nand U2865 (N_2865,N_2635,N_2794);
or U2866 (N_2866,N_2672,N_2643);
and U2867 (N_2867,N_2797,N_2620);
or U2868 (N_2868,N_2772,N_2758);
nand U2869 (N_2869,N_2645,N_2755);
or U2870 (N_2870,N_2618,N_2721);
nor U2871 (N_2871,N_2700,N_2603);
xnor U2872 (N_2872,N_2716,N_2673);
or U2873 (N_2873,N_2601,N_2753);
nor U2874 (N_2874,N_2638,N_2722);
and U2875 (N_2875,N_2742,N_2796);
nor U2876 (N_2876,N_2699,N_2637);
or U2877 (N_2877,N_2650,N_2625);
nor U2878 (N_2878,N_2687,N_2633);
or U2879 (N_2879,N_2719,N_2731);
and U2880 (N_2880,N_2608,N_2640);
or U2881 (N_2881,N_2776,N_2694);
nor U2882 (N_2882,N_2696,N_2613);
and U2883 (N_2883,N_2781,N_2747);
and U2884 (N_2884,N_2661,N_2642);
xor U2885 (N_2885,N_2679,N_2602);
nor U2886 (N_2886,N_2663,N_2614);
or U2887 (N_2887,N_2631,N_2714);
nand U2888 (N_2888,N_2648,N_2786);
nand U2889 (N_2889,N_2762,N_2787);
nand U2890 (N_2890,N_2761,N_2703);
and U2891 (N_2891,N_2616,N_2708);
xnor U2892 (N_2892,N_2658,N_2619);
nor U2893 (N_2893,N_2698,N_2728);
nor U2894 (N_2894,N_2717,N_2727);
nand U2895 (N_2895,N_2720,N_2737);
and U2896 (N_2896,N_2652,N_2657);
nand U2897 (N_2897,N_2621,N_2604);
nor U2898 (N_2898,N_2748,N_2697);
nor U2899 (N_2899,N_2627,N_2655);
nand U2900 (N_2900,N_2647,N_2629);
nor U2901 (N_2901,N_2690,N_2602);
and U2902 (N_2902,N_2696,N_2642);
nand U2903 (N_2903,N_2776,N_2750);
nand U2904 (N_2904,N_2639,N_2758);
and U2905 (N_2905,N_2681,N_2606);
or U2906 (N_2906,N_2751,N_2609);
or U2907 (N_2907,N_2623,N_2696);
xnor U2908 (N_2908,N_2686,N_2688);
nor U2909 (N_2909,N_2756,N_2795);
xnor U2910 (N_2910,N_2661,N_2600);
and U2911 (N_2911,N_2726,N_2773);
nor U2912 (N_2912,N_2657,N_2791);
nor U2913 (N_2913,N_2610,N_2608);
nand U2914 (N_2914,N_2638,N_2627);
and U2915 (N_2915,N_2792,N_2703);
or U2916 (N_2916,N_2710,N_2777);
nor U2917 (N_2917,N_2607,N_2693);
nor U2918 (N_2918,N_2684,N_2783);
nand U2919 (N_2919,N_2784,N_2713);
and U2920 (N_2920,N_2698,N_2727);
and U2921 (N_2921,N_2769,N_2782);
nand U2922 (N_2922,N_2610,N_2615);
or U2923 (N_2923,N_2731,N_2751);
xor U2924 (N_2924,N_2636,N_2717);
and U2925 (N_2925,N_2657,N_2631);
nand U2926 (N_2926,N_2675,N_2695);
and U2927 (N_2927,N_2620,N_2747);
and U2928 (N_2928,N_2677,N_2718);
and U2929 (N_2929,N_2746,N_2675);
xnor U2930 (N_2930,N_2778,N_2643);
or U2931 (N_2931,N_2622,N_2761);
or U2932 (N_2932,N_2705,N_2766);
xnor U2933 (N_2933,N_2680,N_2610);
or U2934 (N_2934,N_2761,N_2677);
nand U2935 (N_2935,N_2726,N_2766);
or U2936 (N_2936,N_2609,N_2652);
nand U2937 (N_2937,N_2753,N_2751);
or U2938 (N_2938,N_2677,N_2780);
or U2939 (N_2939,N_2681,N_2724);
and U2940 (N_2940,N_2701,N_2695);
xnor U2941 (N_2941,N_2758,N_2765);
nor U2942 (N_2942,N_2729,N_2701);
nand U2943 (N_2943,N_2723,N_2653);
xor U2944 (N_2944,N_2729,N_2747);
nand U2945 (N_2945,N_2725,N_2656);
or U2946 (N_2946,N_2681,N_2642);
and U2947 (N_2947,N_2794,N_2709);
nand U2948 (N_2948,N_2763,N_2676);
nand U2949 (N_2949,N_2677,N_2632);
nor U2950 (N_2950,N_2773,N_2638);
nand U2951 (N_2951,N_2624,N_2757);
nor U2952 (N_2952,N_2666,N_2607);
nor U2953 (N_2953,N_2611,N_2687);
and U2954 (N_2954,N_2651,N_2629);
nand U2955 (N_2955,N_2621,N_2779);
nand U2956 (N_2956,N_2786,N_2731);
nand U2957 (N_2957,N_2691,N_2696);
nor U2958 (N_2958,N_2713,N_2667);
nor U2959 (N_2959,N_2604,N_2697);
or U2960 (N_2960,N_2711,N_2779);
xnor U2961 (N_2961,N_2619,N_2776);
and U2962 (N_2962,N_2669,N_2726);
or U2963 (N_2963,N_2626,N_2780);
and U2964 (N_2964,N_2743,N_2679);
nand U2965 (N_2965,N_2775,N_2623);
and U2966 (N_2966,N_2664,N_2783);
xor U2967 (N_2967,N_2651,N_2669);
nand U2968 (N_2968,N_2772,N_2787);
or U2969 (N_2969,N_2793,N_2799);
or U2970 (N_2970,N_2735,N_2688);
xnor U2971 (N_2971,N_2640,N_2618);
nor U2972 (N_2972,N_2749,N_2778);
nand U2973 (N_2973,N_2782,N_2716);
nand U2974 (N_2974,N_2668,N_2682);
or U2975 (N_2975,N_2767,N_2661);
nand U2976 (N_2976,N_2684,N_2628);
nand U2977 (N_2977,N_2749,N_2636);
nor U2978 (N_2978,N_2759,N_2748);
or U2979 (N_2979,N_2653,N_2639);
or U2980 (N_2980,N_2750,N_2795);
nand U2981 (N_2981,N_2692,N_2625);
or U2982 (N_2982,N_2780,N_2732);
nor U2983 (N_2983,N_2607,N_2699);
nand U2984 (N_2984,N_2614,N_2691);
nor U2985 (N_2985,N_2715,N_2769);
or U2986 (N_2986,N_2793,N_2641);
nor U2987 (N_2987,N_2794,N_2748);
nand U2988 (N_2988,N_2626,N_2738);
or U2989 (N_2989,N_2634,N_2663);
nand U2990 (N_2990,N_2786,N_2686);
xnor U2991 (N_2991,N_2726,N_2630);
nand U2992 (N_2992,N_2787,N_2620);
or U2993 (N_2993,N_2791,N_2678);
or U2994 (N_2994,N_2669,N_2658);
or U2995 (N_2995,N_2677,N_2765);
xnor U2996 (N_2996,N_2640,N_2606);
nor U2997 (N_2997,N_2604,N_2625);
nor U2998 (N_2998,N_2674,N_2706);
xor U2999 (N_2999,N_2686,N_2716);
or U3000 (N_3000,N_2876,N_2916);
nand U3001 (N_3001,N_2977,N_2878);
nand U3002 (N_3002,N_2854,N_2870);
and U3003 (N_3003,N_2840,N_2936);
nor U3004 (N_3004,N_2990,N_2868);
nand U3005 (N_3005,N_2901,N_2995);
nand U3006 (N_3006,N_2938,N_2985);
or U3007 (N_3007,N_2869,N_2902);
nor U3008 (N_3008,N_2927,N_2818);
or U3009 (N_3009,N_2867,N_2893);
nor U3010 (N_3010,N_2826,N_2863);
nor U3011 (N_3011,N_2883,N_2884);
and U3012 (N_3012,N_2871,N_2802);
nor U3013 (N_3013,N_2856,N_2830);
nor U3014 (N_3014,N_2887,N_2941);
and U3015 (N_3015,N_2843,N_2973);
or U3016 (N_3016,N_2807,N_2858);
nand U3017 (N_3017,N_2874,N_2851);
nor U3018 (N_3018,N_2993,N_2958);
or U3019 (N_3019,N_2957,N_2945);
or U3020 (N_3020,N_2805,N_2821);
and U3021 (N_3021,N_2994,N_2906);
or U3022 (N_3022,N_2837,N_2862);
nor U3023 (N_3023,N_2976,N_2801);
nor U3024 (N_3024,N_2815,N_2888);
and U3025 (N_3025,N_2865,N_2980);
or U3026 (N_3026,N_2953,N_2829);
and U3027 (N_3027,N_2820,N_2929);
nor U3028 (N_3028,N_2983,N_2895);
nor U3029 (N_3029,N_2924,N_2838);
nand U3030 (N_3030,N_2951,N_2948);
nand U3031 (N_3031,N_2885,N_2882);
nor U3032 (N_3032,N_2986,N_2970);
nand U3033 (N_3033,N_2839,N_2812);
nand U3034 (N_3034,N_2825,N_2959);
or U3035 (N_3035,N_2930,N_2928);
nor U3036 (N_3036,N_2920,N_2833);
or U3037 (N_3037,N_2956,N_2900);
or U3038 (N_3038,N_2947,N_2940);
or U3039 (N_3039,N_2914,N_2824);
nand U3040 (N_3040,N_2831,N_2817);
and U3041 (N_3041,N_2827,N_2890);
nand U3042 (N_3042,N_2964,N_2909);
nor U3043 (N_3043,N_2861,N_2923);
or U3044 (N_3044,N_2905,N_2939);
and U3045 (N_3045,N_2999,N_2960);
and U3046 (N_3046,N_2950,N_2992);
or U3047 (N_3047,N_2850,N_2955);
nor U3048 (N_3048,N_2849,N_2808);
nand U3049 (N_3049,N_2859,N_2896);
nand U3050 (N_3050,N_2918,N_2919);
and U3051 (N_3051,N_2915,N_2813);
or U3052 (N_3052,N_2847,N_2907);
nand U3053 (N_3053,N_2917,N_2879);
or U3054 (N_3054,N_2963,N_2889);
nand U3055 (N_3055,N_2968,N_2877);
nand U3056 (N_3056,N_2969,N_2962);
nand U3057 (N_3057,N_2800,N_2943);
nand U3058 (N_3058,N_2966,N_2855);
nand U3059 (N_3059,N_2810,N_2875);
nand U3060 (N_3060,N_2903,N_2809);
nand U3061 (N_3061,N_2848,N_2997);
xnor U3062 (N_3062,N_2832,N_2897);
and U3063 (N_3063,N_2836,N_2845);
or U3064 (N_3064,N_2921,N_2841);
nor U3065 (N_3065,N_2996,N_2816);
nor U3066 (N_3066,N_2908,N_2844);
xnor U3067 (N_3067,N_2852,N_2864);
nor U3068 (N_3068,N_2981,N_2819);
and U3069 (N_3069,N_2881,N_2892);
nand U3070 (N_3070,N_2931,N_2811);
nor U3071 (N_3071,N_2926,N_2835);
and U3072 (N_3072,N_2942,N_2842);
and U3073 (N_3073,N_2911,N_2971);
nor U3074 (N_3074,N_2934,N_2922);
nand U3075 (N_3075,N_2944,N_2873);
nor U3076 (N_3076,N_2972,N_2822);
nor U3077 (N_3077,N_2899,N_2967);
and U3078 (N_3078,N_2932,N_2946);
nand U3079 (N_3079,N_2952,N_2828);
nand U3080 (N_3080,N_2978,N_2898);
nor U3081 (N_3081,N_2806,N_2857);
nor U3082 (N_3082,N_2886,N_2974);
and U3083 (N_3083,N_2912,N_2987);
and U3084 (N_3084,N_2803,N_2880);
nor U3085 (N_3085,N_2979,N_2834);
nor U3086 (N_3086,N_2975,N_2988);
or U3087 (N_3087,N_2853,N_2991);
and U3088 (N_3088,N_2823,N_2814);
nor U3089 (N_3089,N_2846,N_2910);
or U3090 (N_3090,N_2984,N_2935);
xor U3091 (N_3091,N_2866,N_2933);
and U3092 (N_3092,N_2891,N_2937);
or U3093 (N_3093,N_2913,N_2904);
nor U3094 (N_3094,N_2860,N_2804);
nor U3095 (N_3095,N_2998,N_2894);
or U3096 (N_3096,N_2989,N_2872);
xnor U3097 (N_3097,N_2961,N_2982);
nor U3098 (N_3098,N_2925,N_2954);
xor U3099 (N_3099,N_2965,N_2949);
nand U3100 (N_3100,N_2893,N_2970);
and U3101 (N_3101,N_2903,N_2901);
and U3102 (N_3102,N_2805,N_2951);
and U3103 (N_3103,N_2943,N_2903);
nand U3104 (N_3104,N_2803,N_2834);
and U3105 (N_3105,N_2879,N_2866);
nor U3106 (N_3106,N_2880,N_2929);
and U3107 (N_3107,N_2896,N_2989);
and U3108 (N_3108,N_2916,N_2897);
nand U3109 (N_3109,N_2942,N_2831);
and U3110 (N_3110,N_2921,N_2886);
nor U3111 (N_3111,N_2869,N_2814);
nor U3112 (N_3112,N_2851,N_2833);
nand U3113 (N_3113,N_2829,N_2841);
and U3114 (N_3114,N_2928,N_2839);
nand U3115 (N_3115,N_2915,N_2889);
nand U3116 (N_3116,N_2933,N_2872);
nor U3117 (N_3117,N_2942,N_2976);
or U3118 (N_3118,N_2876,N_2817);
nand U3119 (N_3119,N_2867,N_2908);
and U3120 (N_3120,N_2913,N_2989);
nand U3121 (N_3121,N_2825,N_2921);
and U3122 (N_3122,N_2894,N_2912);
nor U3123 (N_3123,N_2970,N_2957);
or U3124 (N_3124,N_2827,N_2843);
or U3125 (N_3125,N_2919,N_2986);
xor U3126 (N_3126,N_2929,N_2802);
or U3127 (N_3127,N_2875,N_2842);
and U3128 (N_3128,N_2971,N_2886);
or U3129 (N_3129,N_2860,N_2993);
or U3130 (N_3130,N_2988,N_2867);
and U3131 (N_3131,N_2974,N_2888);
nand U3132 (N_3132,N_2843,N_2896);
and U3133 (N_3133,N_2846,N_2872);
or U3134 (N_3134,N_2976,N_2805);
nand U3135 (N_3135,N_2909,N_2919);
nand U3136 (N_3136,N_2849,N_2844);
or U3137 (N_3137,N_2994,N_2940);
or U3138 (N_3138,N_2824,N_2897);
or U3139 (N_3139,N_2995,N_2823);
nand U3140 (N_3140,N_2928,N_2912);
or U3141 (N_3141,N_2857,N_2912);
nor U3142 (N_3142,N_2800,N_2878);
nand U3143 (N_3143,N_2899,N_2837);
nor U3144 (N_3144,N_2933,N_2948);
nand U3145 (N_3145,N_2913,N_2884);
or U3146 (N_3146,N_2893,N_2877);
or U3147 (N_3147,N_2907,N_2868);
or U3148 (N_3148,N_2910,N_2993);
or U3149 (N_3149,N_2810,N_2876);
or U3150 (N_3150,N_2872,N_2807);
nand U3151 (N_3151,N_2980,N_2928);
nand U3152 (N_3152,N_2995,N_2824);
nor U3153 (N_3153,N_2909,N_2984);
or U3154 (N_3154,N_2973,N_2977);
nand U3155 (N_3155,N_2805,N_2964);
and U3156 (N_3156,N_2974,N_2934);
and U3157 (N_3157,N_2981,N_2921);
or U3158 (N_3158,N_2908,N_2883);
nand U3159 (N_3159,N_2872,N_2811);
or U3160 (N_3160,N_2841,N_2803);
nand U3161 (N_3161,N_2813,N_2812);
or U3162 (N_3162,N_2826,N_2911);
and U3163 (N_3163,N_2978,N_2963);
or U3164 (N_3164,N_2920,N_2883);
xor U3165 (N_3165,N_2914,N_2935);
xnor U3166 (N_3166,N_2928,N_2823);
nand U3167 (N_3167,N_2869,N_2995);
nand U3168 (N_3168,N_2864,N_2887);
nor U3169 (N_3169,N_2853,N_2910);
nand U3170 (N_3170,N_2861,N_2941);
nor U3171 (N_3171,N_2815,N_2933);
nor U3172 (N_3172,N_2956,N_2892);
and U3173 (N_3173,N_2977,N_2871);
xor U3174 (N_3174,N_2911,N_2864);
or U3175 (N_3175,N_2833,N_2820);
and U3176 (N_3176,N_2901,N_2866);
and U3177 (N_3177,N_2931,N_2978);
nand U3178 (N_3178,N_2907,N_2953);
or U3179 (N_3179,N_2887,N_2953);
and U3180 (N_3180,N_2987,N_2891);
or U3181 (N_3181,N_2933,N_2914);
and U3182 (N_3182,N_2957,N_2946);
nor U3183 (N_3183,N_2878,N_2838);
nand U3184 (N_3184,N_2840,N_2905);
nand U3185 (N_3185,N_2916,N_2804);
nand U3186 (N_3186,N_2983,N_2911);
nand U3187 (N_3187,N_2956,N_2835);
or U3188 (N_3188,N_2938,N_2997);
nor U3189 (N_3189,N_2944,N_2990);
nand U3190 (N_3190,N_2954,N_2834);
nor U3191 (N_3191,N_2840,N_2985);
and U3192 (N_3192,N_2894,N_2839);
nor U3193 (N_3193,N_2921,N_2917);
nand U3194 (N_3194,N_2807,N_2913);
xor U3195 (N_3195,N_2961,N_2888);
nor U3196 (N_3196,N_2924,N_2920);
nand U3197 (N_3197,N_2927,N_2807);
and U3198 (N_3198,N_2816,N_2832);
nand U3199 (N_3199,N_2863,N_2985);
xor U3200 (N_3200,N_3040,N_3126);
and U3201 (N_3201,N_3020,N_3085);
or U3202 (N_3202,N_3194,N_3180);
and U3203 (N_3203,N_3129,N_3139);
nand U3204 (N_3204,N_3113,N_3197);
nor U3205 (N_3205,N_3029,N_3012);
xor U3206 (N_3206,N_3195,N_3140);
nor U3207 (N_3207,N_3125,N_3080);
nand U3208 (N_3208,N_3013,N_3193);
and U3209 (N_3209,N_3145,N_3004);
xnor U3210 (N_3210,N_3019,N_3042);
nand U3211 (N_3211,N_3107,N_3133);
or U3212 (N_3212,N_3101,N_3088);
and U3213 (N_3213,N_3167,N_3161);
nor U3214 (N_3214,N_3196,N_3064);
or U3215 (N_3215,N_3060,N_3141);
nand U3216 (N_3216,N_3175,N_3168);
nor U3217 (N_3217,N_3047,N_3059);
xor U3218 (N_3218,N_3044,N_3084);
or U3219 (N_3219,N_3138,N_3031);
or U3220 (N_3220,N_3137,N_3028);
and U3221 (N_3221,N_3102,N_3067);
or U3222 (N_3222,N_3186,N_3163);
or U3223 (N_3223,N_3049,N_3151);
or U3224 (N_3224,N_3165,N_3043);
nand U3225 (N_3225,N_3173,N_3035);
nor U3226 (N_3226,N_3018,N_3053);
nand U3227 (N_3227,N_3144,N_3191);
nor U3228 (N_3228,N_3000,N_3070);
nor U3229 (N_3229,N_3025,N_3094);
nor U3230 (N_3230,N_3002,N_3091);
and U3231 (N_3231,N_3150,N_3009);
and U3232 (N_3232,N_3072,N_3066);
nand U3233 (N_3233,N_3117,N_3081);
and U3234 (N_3234,N_3185,N_3045);
or U3235 (N_3235,N_3065,N_3055);
nand U3236 (N_3236,N_3082,N_3164);
and U3237 (N_3237,N_3152,N_3007);
or U3238 (N_3238,N_3179,N_3112);
nor U3239 (N_3239,N_3127,N_3003);
xor U3240 (N_3240,N_3100,N_3036);
nor U3241 (N_3241,N_3011,N_3052);
nor U3242 (N_3242,N_3027,N_3010);
nand U3243 (N_3243,N_3083,N_3069);
xor U3244 (N_3244,N_3178,N_3098);
xor U3245 (N_3245,N_3030,N_3132);
or U3246 (N_3246,N_3021,N_3177);
nand U3247 (N_3247,N_3130,N_3014);
nand U3248 (N_3248,N_3038,N_3170);
nand U3249 (N_3249,N_3001,N_3147);
or U3250 (N_3250,N_3162,N_3048);
and U3251 (N_3251,N_3041,N_3099);
nor U3252 (N_3252,N_3121,N_3017);
or U3253 (N_3253,N_3093,N_3058);
nor U3254 (N_3254,N_3056,N_3149);
and U3255 (N_3255,N_3096,N_3192);
and U3256 (N_3256,N_3166,N_3181);
nor U3257 (N_3257,N_3057,N_3157);
nand U3258 (N_3258,N_3115,N_3090);
xnor U3259 (N_3259,N_3171,N_3135);
nor U3260 (N_3260,N_3148,N_3054);
and U3261 (N_3261,N_3119,N_3037);
xnor U3262 (N_3262,N_3160,N_3079);
or U3263 (N_3263,N_3199,N_3134);
nor U3264 (N_3264,N_3187,N_3077);
nand U3265 (N_3265,N_3174,N_3032);
and U3266 (N_3266,N_3154,N_3189);
nand U3267 (N_3267,N_3024,N_3095);
nor U3268 (N_3268,N_3097,N_3172);
or U3269 (N_3269,N_3155,N_3026);
and U3270 (N_3270,N_3122,N_3153);
nor U3271 (N_3271,N_3076,N_3022);
or U3272 (N_3272,N_3190,N_3087);
or U3273 (N_3273,N_3128,N_3078);
nor U3274 (N_3274,N_3075,N_3184);
or U3275 (N_3275,N_3016,N_3183);
nor U3276 (N_3276,N_3063,N_3061);
nand U3277 (N_3277,N_3131,N_3074);
nand U3278 (N_3278,N_3062,N_3106);
nand U3279 (N_3279,N_3023,N_3089);
and U3280 (N_3280,N_3086,N_3123);
nand U3281 (N_3281,N_3092,N_3008);
nor U3282 (N_3282,N_3110,N_3159);
nand U3283 (N_3283,N_3182,N_3033);
and U3284 (N_3284,N_3118,N_3142);
nor U3285 (N_3285,N_3111,N_3105);
and U3286 (N_3286,N_3198,N_3104);
or U3287 (N_3287,N_3176,N_3120);
and U3288 (N_3288,N_3108,N_3051);
and U3289 (N_3289,N_3039,N_3071);
and U3290 (N_3290,N_3109,N_3116);
or U3291 (N_3291,N_3103,N_3114);
or U3292 (N_3292,N_3143,N_3136);
and U3293 (N_3293,N_3146,N_3050);
nand U3294 (N_3294,N_3034,N_3006);
or U3295 (N_3295,N_3156,N_3073);
nand U3296 (N_3296,N_3158,N_3124);
or U3297 (N_3297,N_3169,N_3068);
or U3298 (N_3298,N_3005,N_3188);
and U3299 (N_3299,N_3015,N_3046);
nand U3300 (N_3300,N_3002,N_3104);
and U3301 (N_3301,N_3095,N_3129);
xor U3302 (N_3302,N_3002,N_3123);
or U3303 (N_3303,N_3159,N_3064);
nor U3304 (N_3304,N_3045,N_3064);
nor U3305 (N_3305,N_3021,N_3017);
nand U3306 (N_3306,N_3028,N_3030);
or U3307 (N_3307,N_3164,N_3108);
nor U3308 (N_3308,N_3016,N_3126);
nor U3309 (N_3309,N_3099,N_3151);
or U3310 (N_3310,N_3175,N_3045);
nor U3311 (N_3311,N_3176,N_3024);
and U3312 (N_3312,N_3021,N_3175);
nand U3313 (N_3313,N_3166,N_3084);
nor U3314 (N_3314,N_3122,N_3198);
or U3315 (N_3315,N_3072,N_3084);
nand U3316 (N_3316,N_3040,N_3080);
nand U3317 (N_3317,N_3095,N_3195);
nor U3318 (N_3318,N_3159,N_3183);
and U3319 (N_3319,N_3148,N_3012);
or U3320 (N_3320,N_3029,N_3147);
and U3321 (N_3321,N_3139,N_3101);
and U3322 (N_3322,N_3159,N_3111);
and U3323 (N_3323,N_3019,N_3105);
nand U3324 (N_3324,N_3145,N_3156);
and U3325 (N_3325,N_3025,N_3064);
or U3326 (N_3326,N_3010,N_3032);
or U3327 (N_3327,N_3074,N_3077);
nor U3328 (N_3328,N_3071,N_3145);
and U3329 (N_3329,N_3197,N_3058);
nor U3330 (N_3330,N_3199,N_3027);
or U3331 (N_3331,N_3102,N_3095);
nor U3332 (N_3332,N_3144,N_3078);
nand U3333 (N_3333,N_3092,N_3080);
nand U3334 (N_3334,N_3000,N_3199);
nor U3335 (N_3335,N_3101,N_3168);
nand U3336 (N_3336,N_3090,N_3100);
or U3337 (N_3337,N_3066,N_3012);
nand U3338 (N_3338,N_3164,N_3025);
or U3339 (N_3339,N_3139,N_3175);
nand U3340 (N_3340,N_3154,N_3042);
or U3341 (N_3341,N_3128,N_3055);
and U3342 (N_3342,N_3164,N_3154);
or U3343 (N_3343,N_3078,N_3037);
nor U3344 (N_3344,N_3191,N_3060);
nor U3345 (N_3345,N_3198,N_3133);
nor U3346 (N_3346,N_3001,N_3057);
nor U3347 (N_3347,N_3051,N_3052);
nor U3348 (N_3348,N_3039,N_3152);
or U3349 (N_3349,N_3032,N_3012);
and U3350 (N_3350,N_3007,N_3098);
xnor U3351 (N_3351,N_3029,N_3129);
or U3352 (N_3352,N_3106,N_3001);
or U3353 (N_3353,N_3191,N_3169);
nand U3354 (N_3354,N_3117,N_3143);
nand U3355 (N_3355,N_3043,N_3054);
nor U3356 (N_3356,N_3011,N_3149);
xnor U3357 (N_3357,N_3058,N_3045);
and U3358 (N_3358,N_3169,N_3129);
or U3359 (N_3359,N_3188,N_3101);
and U3360 (N_3360,N_3113,N_3062);
and U3361 (N_3361,N_3171,N_3176);
and U3362 (N_3362,N_3016,N_3146);
or U3363 (N_3363,N_3089,N_3019);
nor U3364 (N_3364,N_3041,N_3172);
and U3365 (N_3365,N_3003,N_3077);
and U3366 (N_3366,N_3023,N_3000);
nor U3367 (N_3367,N_3159,N_3002);
and U3368 (N_3368,N_3075,N_3003);
and U3369 (N_3369,N_3071,N_3033);
and U3370 (N_3370,N_3146,N_3176);
nor U3371 (N_3371,N_3199,N_3014);
or U3372 (N_3372,N_3050,N_3111);
nor U3373 (N_3373,N_3013,N_3022);
xor U3374 (N_3374,N_3036,N_3033);
or U3375 (N_3375,N_3151,N_3169);
nor U3376 (N_3376,N_3135,N_3165);
nand U3377 (N_3377,N_3074,N_3092);
nor U3378 (N_3378,N_3109,N_3035);
nand U3379 (N_3379,N_3026,N_3014);
xnor U3380 (N_3380,N_3138,N_3084);
or U3381 (N_3381,N_3066,N_3195);
nor U3382 (N_3382,N_3064,N_3053);
nor U3383 (N_3383,N_3010,N_3067);
or U3384 (N_3384,N_3145,N_3104);
nand U3385 (N_3385,N_3146,N_3128);
nor U3386 (N_3386,N_3069,N_3000);
and U3387 (N_3387,N_3127,N_3147);
and U3388 (N_3388,N_3106,N_3025);
nor U3389 (N_3389,N_3107,N_3199);
or U3390 (N_3390,N_3175,N_3186);
or U3391 (N_3391,N_3066,N_3032);
nand U3392 (N_3392,N_3178,N_3090);
and U3393 (N_3393,N_3177,N_3013);
or U3394 (N_3394,N_3124,N_3099);
nand U3395 (N_3395,N_3045,N_3133);
nor U3396 (N_3396,N_3039,N_3043);
nor U3397 (N_3397,N_3173,N_3086);
nor U3398 (N_3398,N_3021,N_3132);
xnor U3399 (N_3399,N_3039,N_3189);
nor U3400 (N_3400,N_3227,N_3262);
or U3401 (N_3401,N_3337,N_3317);
or U3402 (N_3402,N_3360,N_3283);
nor U3403 (N_3403,N_3391,N_3326);
or U3404 (N_3404,N_3387,N_3381);
and U3405 (N_3405,N_3269,N_3295);
or U3406 (N_3406,N_3256,N_3340);
nor U3407 (N_3407,N_3257,N_3341);
nor U3408 (N_3408,N_3253,N_3325);
or U3409 (N_3409,N_3343,N_3298);
nor U3410 (N_3410,N_3372,N_3225);
xor U3411 (N_3411,N_3328,N_3280);
nand U3412 (N_3412,N_3264,N_3393);
nor U3413 (N_3413,N_3357,N_3306);
or U3414 (N_3414,N_3375,N_3263);
or U3415 (N_3415,N_3378,N_3331);
and U3416 (N_3416,N_3338,N_3354);
and U3417 (N_3417,N_3274,N_3207);
and U3418 (N_3418,N_3273,N_3202);
or U3419 (N_3419,N_3342,N_3254);
and U3420 (N_3420,N_3310,N_3228);
nand U3421 (N_3421,N_3349,N_3388);
and U3422 (N_3422,N_3235,N_3332);
nand U3423 (N_3423,N_3327,N_3287);
or U3424 (N_3424,N_3292,N_3397);
or U3425 (N_3425,N_3311,N_3205);
nor U3426 (N_3426,N_3308,N_3284);
or U3427 (N_3427,N_3210,N_3245);
nor U3428 (N_3428,N_3209,N_3282);
nand U3429 (N_3429,N_3222,N_3290);
nor U3430 (N_3430,N_3220,N_3203);
and U3431 (N_3431,N_3250,N_3398);
and U3432 (N_3432,N_3322,N_3335);
and U3433 (N_3433,N_3318,N_3352);
nand U3434 (N_3434,N_3217,N_3286);
nand U3435 (N_3435,N_3334,N_3214);
nand U3436 (N_3436,N_3396,N_3383);
nor U3437 (N_3437,N_3297,N_3369);
nand U3438 (N_3438,N_3353,N_3305);
nor U3439 (N_3439,N_3304,N_3293);
nor U3440 (N_3440,N_3336,N_3278);
nor U3441 (N_3441,N_3246,N_3277);
nor U3442 (N_3442,N_3365,N_3260);
nor U3443 (N_3443,N_3316,N_3212);
xor U3444 (N_3444,N_3265,N_3211);
or U3445 (N_3445,N_3233,N_3301);
and U3446 (N_3446,N_3309,N_3392);
nor U3447 (N_3447,N_3348,N_3276);
nor U3448 (N_3448,N_3355,N_3275);
nor U3449 (N_3449,N_3288,N_3359);
nor U3450 (N_3450,N_3386,N_3314);
and U3451 (N_3451,N_3270,N_3201);
or U3452 (N_3452,N_3339,N_3234);
and U3453 (N_3453,N_3279,N_3204);
and U3454 (N_3454,N_3226,N_3267);
nand U3455 (N_3455,N_3307,N_3266);
xnor U3456 (N_3456,N_3313,N_3382);
or U3457 (N_3457,N_3380,N_3200);
or U3458 (N_3458,N_3320,N_3206);
or U3459 (N_3459,N_3368,N_3244);
nor U3460 (N_3460,N_3347,N_3376);
nand U3461 (N_3461,N_3224,N_3239);
or U3462 (N_3462,N_3231,N_3315);
nor U3463 (N_3463,N_3370,N_3251);
nor U3464 (N_3464,N_3259,N_3361);
and U3465 (N_3465,N_3249,N_3285);
nand U3466 (N_3466,N_3216,N_3364);
and U3467 (N_3467,N_3367,N_3242);
nor U3468 (N_3468,N_3300,N_3268);
nor U3469 (N_3469,N_3356,N_3241);
or U3470 (N_3470,N_3296,N_3255);
or U3471 (N_3471,N_3243,N_3344);
xnor U3472 (N_3472,N_3321,N_3333);
and U3473 (N_3473,N_3351,N_3399);
and U3474 (N_3474,N_3261,N_3395);
or U3475 (N_3475,N_3384,N_3248);
xor U3476 (N_3476,N_3294,N_3358);
nand U3477 (N_3477,N_3236,N_3299);
nor U3478 (N_3478,N_3363,N_3346);
and U3479 (N_3479,N_3208,N_3330);
and U3480 (N_3480,N_3329,N_3390);
and U3481 (N_3481,N_3394,N_3221);
and U3482 (N_3482,N_3366,N_3324);
or U3483 (N_3483,N_3223,N_3232);
nor U3484 (N_3484,N_3272,N_3350);
or U3485 (N_3485,N_3389,N_3215);
and U3486 (N_3486,N_3291,N_3385);
nor U3487 (N_3487,N_3312,N_3362);
and U3488 (N_3488,N_3379,N_3237);
nand U3489 (N_3489,N_3374,N_3252);
and U3490 (N_3490,N_3218,N_3258);
nand U3491 (N_3491,N_3213,N_3377);
or U3492 (N_3492,N_3281,N_3303);
nor U3493 (N_3493,N_3323,N_3240);
xor U3494 (N_3494,N_3271,N_3371);
and U3495 (N_3495,N_3219,N_3302);
and U3496 (N_3496,N_3345,N_3373);
xor U3497 (N_3497,N_3238,N_3247);
and U3498 (N_3498,N_3229,N_3230);
nor U3499 (N_3499,N_3319,N_3289);
and U3500 (N_3500,N_3208,N_3352);
or U3501 (N_3501,N_3256,N_3234);
nor U3502 (N_3502,N_3358,N_3263);
or U3503 (N_3503,N_3206,N_3299);
nand U3504 (N_3504,N_3381,N_3237);
or U3505 (N_3505,N_3329,N_3260);
and U3506 (N_3506,N_3333,N_3366);
nand U3507 (N_3507,N_3319,N_3251);
nor U3508 (N_3508,N_3248,N_3366);
nor U3509 (N_3509,N_3372,N_3300);
nand U3510 (N_3510,N_3334,N_3215);
nor U3511 (N_3511,N_3339,N_3329);
and U3512 (N_3512,N_3351,N_3380);
xnor U3513 (N_3513,N_3315,N_3212);
nand U3514 (N_3514,N_3258,N_3344);
nor U3515 (N_3515,N_3318,N_3229);
xor U3516 (N_3516,N_3306,N_3313);
nor U3517 (N_3517,N_3343,N_3276);
nand U3518 (N_3518,N_3285,N_3246);
or U3519 (N_3519,N_3353,N_3385);
nor U3520 (N_3520,N_3397,N_3337);
nor U3521 (N_3521,N_3280,N_3300);
xor U3522 (N_3522,N_3270,N_3215);
nand U3523 (N_3523,N_3262,N_3250);
and U3524 (N_3524,N_3296,N_3320);
or U3525 (N_3525,N_3367,N_3310);
nand U3526 (N_3526,N_3347,N_3266);
or U3527 (N_3527,N_3371,N_3335);
or U3528 (N_3528,N_3314,N_3270);
xnor U3529 (N_3529,N_3345,N_3330);
or U3530 (N_3530,N_3281,N_3302);
nand U3531 (N_3531,N_3346,N_3289);
nor U3532 (N_3532,N_3378,N_3353);
xnor U3533 (N_3533,N_3313,N_3384);
or U3534 (N_3534,N_3341,N_3356);
or U3535 (N_3535,N_3202,N_3314);
nor U3536 (N_3536,N_3283,N_3355);
or U3537 (N_3537,N_3233,N_3365);
nand U3538 (N_3538,N_3356,N_3319);
nand U3539 (N_3539,N_3297,N_3232);
and U3540 (N_3540,N_3390,N_3342);
nand U3541 (N_3541,N_3208,N_3262);
and U3542 (N_3542,N_3329,N_3203);
nor U3543 (N_3543,N_3342,N_3292);
nand U3544 (N_3544,N_3382,N_3256);
nand U3545 (N_3545,N_3379,N_3280);
xor U3546 (N_3546,N_3240,N_3338);
and U3547 (N_3547,N_3247,N_3366);
or U3548 (N_3548,N_3315,N_3301);
nand U3549 (N_3549,N_3238,N_3275);
nor U3550 (N_3550,N_3278,N_3354);
nor U3551 (N_3551,N_3228,N_3244);
and U3552 (N_3552,N_3294,N_3216);
xor U3553 (N_3553,N_3355,N_3202);
or U3554 (N_3554,N_3264,N_3367);
nor U3555 (N_3555,N_3248,N_3219);
and U3556 (N_3556,N_3375,N_3388);
nor U3557 (N_3557,N_3213,N_3229);
nand U3558 (N_3558,N_3334,N_3381);
or U3559 (N_3559,N_3394,N_3378);
or U3560 (N_3560,N_3302,N_3265);
nand U3561 (N_3561,N_3271,N_3348);
or U3562 (N_3562,N_3289,N_3339);
nor U3563 (N_3563,N_3376,N_3299);
and U3564 (N_3564,N_3320,N_3310);
nand U3565 (N_3565,N_3395,N_3348);
or U3566 (N_3566,N_3364,N_3396);
nand U3567 (N_3567,N_3305,N_3349);
and U3568 (N_3568,N_3316,N_3230);
nand U3569 (N_3569,N_3214,N_3259);
nand U3570 (N_3570,N_3298,N_3294);
and U3571 (N_3571,N_3231,N_3368);
nor U3572 (N_3572,N_3384,N_3319);
nor U3573 (N_3573,N_3271,N_3370);
and U3574 (N_3574,N_3382,N_3311);
or U3575 (N_3575,N_3295,N_3381);
or U3576 (N_3576,N_3378,N_3308);
and U3577 (N_3577,N_3222,N_3301);
xnor U3578 (N_3578,N_3398,N_3272);
and U3579 (N_3579,N_3242,N_3386);
xnor U3580 (N_3580,N_3375,N_3361);
or U3581 (N_3581,N_3218,N_3381);
and U3582 (N_3582,N_3292,N_3336);
nand U3583 (N_3583,N_3282,N_3291);
nor U3584 (N_3584,N_3364,N_3320);
or U3585 (N_3585,N_3347,N_3285);
and U3586 (N_3586,N_3231,N_3320);
and U3587 (N_3587,N_3214,N_3349);
or U3588 (N_3588,N_3346,N_3247);
nand U3589 (N_3589,N_3285,N_3254);
nand U3590 (N_3590,N_3372,N_3343);
or U3591 (N_3591,N_3278,N_3357);
or U3592 (N_3592,N_3336,N_3265);
nand U3593 (N_3593,N_3308,N_3265);
nand U3594 (N_3594,N_3398,N_3303);
nor U3595 (N_3595,N_3356,N_3266);
nor U3596 (N_3596,N_3393,N_3278);
xnor U3597 (N_3597,N_3231,N_3211);
nor U3598 (N_3598,N_3385,N_3395);
nor U3599 (N_3599,N_3322,N_3246);
xnor U3600 (N_3600,N_3521,N_3553);
or U3601 (N_3601,N_3468,N_3580);
nor U3602 (N_3602,N_3448,N_3484);
and U3603 (N_3603,N_3482,N_3545);
nor U3604 (N_3604,N_3587,N_3466);
or U3605 (N_3605,N_3523,N_3538);
nor U3606 (N_3606,N_3568,N_3530);
nand U3607 (N_3607,N_3428,N_3502);
nor U3608 (N_3608,N_3411,N_3571);
nor U3609 (N_3609,N_3589,N_3418);
or U3610 (N_3610,N_3540,N_3500);
and U3611 (N_3611,N_3499,N_3507);
or U3612 (N_3612,N_3429,N_3597);
nand U3613 (N_3613,N_3401,N_3400);
or U3614 (N_3614,N_3457,N_3599);
nand U3615 (N_3615,N_3410,N_3470);
xor U3616 (N_3616,N_3539,N_3434);
nor U3617 (N_3617,N_3556,N_3471);
nor U3618 (N_3618,N_3460,N_3421);
xnor U3619 (N_3619,N_3464,N_3423);
nand U3620 (N_3620,N_3406,N_3592);
nor U3621 (N_3621,N_3476,N_3550);
or U3622 (N_3622,N_3497,N_3433);
nand U3623 (N_3623,N_3488,N_3560);
xor U3624 (N_3624,N_3583,N_3420);
or U3625 (N_3625,N_3442,N_3524);
nand U3626 (N_3626,N_3478,N_3426);
nand U3627 (N_3627,N_3537,N_3505);
and U3628 (N_3628,N_3572,N_3472);
or U3629 (N_3629,N_3512,N_3474);
or U3630 (N_3630,N_3573,N_3508);
xnor U3631 (N_3631,N_3593,N_3590);
nor U3632 (N_3632,N_3408,N_3456);
nand U3633 (N_3633,N_3407,N_3437);
nand U3634 (N_3634,N_3492,N_3449);
nand U3635 (N_3635,N_3503,N_3535);
or U3636 (N_3636,N_3419,N_3479);
xor U3637 (N_3637,N_3402,N_3458);
nor U3638 (N_3638,N_3465,N_3447);
and U3639 (N_3639,N_3547,N_3432);
and U3640 (N_3640,N_3534,N_3519);
or U3641 (N_3641,N_3412,N_3588);
and U3642 (N_3642,N_3494,N_3493);
nand U3643 (N_3643,N_3528,N_3529);
nor U3644 (N_3644,N_3452,N_3566);
nor U3645 (N_3645,N_3511,N_3517);
or U3646 (N_3646,N_3549,N_3454);
nor U3647 (N_3647,N_3473,N_3513);
or U3648 (N_3648,N_3565,N_3491);
and U3649 (N_3649,N_3532,N_3489);
or U3650 (N_3650,N_3440,N_3467);
or U3651 (N_3651,N_3595,N_3533);
nor U3652 (N_3652,N_3480,N_3563);
nand U3653 (N_3653,N_3579,N_3515);
xor U3654 (N_3654,N_3561,N_3469);
nand U3655 (N_3655,N_3496,N_3463);
nor U3656 (N_3656,N_3504,N_3430);
or U3657 (N_3657,N_3557,N_3527);
nor U3658 (N_3658,N_3438,N_3541);
and U3659 (N_3659,N_3462,N_3578);
and U3660 (N_3660,N_3435,N_3591);
or U3661 (N_3661,N_3425,N_3436);
nand U3662 (N_3662,N_3575,N_3594);
nor U3663 (N_3663,N_3552,N_3554);
and U3664 (N_3664,N_3481,N_3439);
and U3665 (N_3665,N_3427,N_3431);
nor U3666 (N_3666,N_3567,N_3516);
and U3667 (N_3667,N_3441,N_3586);
xnor U3668 (N_3668,N_3405,N_3558);
nand U3669 (N_3669,N_3510,N_3443);
xor U3670 (N_3670,N_3577,N_3461);
nand U3671 (N_3671,N_3451,N_3446);
nand U3672 (N_3672,N_3555,N_3548);
or U3673 (N_3673,N_3498,N_3551);
or U3674 (N_3674,N_3455,N_3414);
or U3675 (N_3675,N_3409,N_3520);
and U3676 (N_3676,N_3485,N_3486);
and U3677 (N_3677,N_3596,N_3450);
nor U3678 (N_3678,N_3417,N_3584);
nand U3679 (N_3679,N_3444,N_3576);
and U3680 (N_3680,N_3475,N_3542);
xnor U3681 (N_3681,N_3536,N_3526);
or U3682 (N_3682,N_3582,N_3559);
and U3683 (N_3683,N_3403,N_3514);
and U3684 (N_3684,N_3501,N_3509);
and U3685 (N_3685,N_3490,N_3525);
nor U3686 (N_3686,N_3531,N_3562);
nand U3687 (N_3687,N_3422,N_3483);
nor U3688 (N_3688,N_3487,N_3416);
nand U3689 (N_3689,N_3598,N_3413);
and U3690 (N_3690,N_3564,N_3570);
nor U3691 (N_3691,N_3522,N_3544);
nand U3692 (N_3692,N_3518,N_3585);
nand U3693 (N_3693,N_3546,N_3445);
nor U3694 (N_3694,N_3404,N_3424);
nor U3695 (N_3695,N_3569,N_3506);
nand U3696 (N_3696,N_3415,N_3477);
nor U3697 (N_3697,N_3453,N_3574);
nand U3698 (N_3698,N_3581,N_3543);
and U3699 (N_3699,N_3495,N_3459);
or U3700 (N_3700,N_3410,N_3506);
nor U3701 (N_3701,N_3413,N_3561);
or U3702 (N_3702,N_3530,N_3441);
and U3703 (N_3703,N_3528,N_3442);
nand U3704 (N_3704,N_3502,N_3499);
and U3705 (N_3705,N_3430,N_3507);
xnor U3706 (N_3706,N_3472,N_3577);
nor U3707 (N_3707,N_3572,N_3570);
nor U3708 (N_3708,N_3470,N_3404);
or U3709 (N_3709,N_3521,N_3412);
nor U3710 (N_3710,N_3480,N_3457);
or U3711 (N_3711,N_3419,N_3579);
or U3712 (N_3712,N_3500,N_3412);
nor U3713 (N_3713,N_3441,N_3584);
nand U3714 (N_3714,N_3560,N_3522);
nor U3715 (N_3715,N_3570,N_3579);
or U3716 (N_3716,N_3530,N_3492);
nor U3717 (N_3717,N_3520,N_3503);
or U3718 (N_3718,N_3523,N_3435);
and U3719 (N_3719,N_3551,N_3572);
xor U3720 (N_3720,N_3493,N_3423);
and U3721 (N_3721,N_3501,N_3550);
nand U3722 (N_3722,N_3453,N_3458);
or U3723 (N_3723,N_3510,N_3436);
nor U3724 (N_3724,N_3470,N_3500);
or U3725 (N_3725,N_3420,N_3431);
and U3726 (N_3726,N_3533,N_3568);
nand U3727 (N_3727,N_3441,N_3513);
nand U3728 (N_3728,N_3491,N_3553);
or U3729 (N_3729,N_3461,N_3588);
or U3730 (N_3730,N_3516,N_3491);
or U3731 (N_3731,N_3489,N_3575);
and U3732 (N_3732,N_3566,N_3464);
xnor U3733 (N_3733,N_3508,N_3549);
nand U3734 (N_3734,N_3558,N_3406);
and U3735 (N_3735,N_3487,N_3438);
nand U3736 (N_3736,N_3575,N_3496);
and U3737 (N_3737,N_3572,N_3491);
and U3738 (N_3738,N_3481,N_3446);
or U3739 (N_3739,N_3495,N_3461);
nor U3740 (N_3740,N_3585,N_3524);
and U3741 (N_3741,N_3473,N_3594);
nand U3742 (N_3742,N_3499,N_3540);
and U3743 (N_3743,N_3558,N_3569);
and U3744 (N_3744,N_3599,N_3446);
nand U3745 (N_3745,N_3577,N_3436);
nand U3746 (N_3746,N_3551,N_3427);
nor U3747 (N_3747,N_3598,N_3541);
nor U3748 (N_3748,N_3556,N_3453);
nand U3749 (N_3749,N_3473,N_3521);
or U3750 (N_3750,N_3457,N_3525);
nand U3751 (N_3751,N_3506,N_3583);
and U3752 (N_3752,N_3481,N_3470);
nand U3753 (N_3753,N_3462,N_3409);
and U3754 (N_3754,N_3525,N_3439);
nand U3755 (N_3755,N_3490,N_3491);
xnor U3756 (N_3756,N_3540,N_3558);
nand U3757 (N_3757,N_3572,N_3586);
xor U3758 (N_3758,N_3455,N_3556);
and U3759 (N_3759,N_3458,N_3432);
or U3760 (N_3760,N_3416,N_3529);
and U3761 (N_3761,N_3474,N_3487);
nor U3762 (N_3762,N_3576,N_3438);
and U3763 (N_3763,N_3543,N_3433);
nor U3764 (N_3764,N_3567,N_3528);
xnor U3765 (N_3765,N_3566,N_3543);
nor U3766 (N_3766,N_3452,N_3555);
and U3767 (N_3767,N_3479,N_3554);
nand U3768 (N_3768,N_3403,N_3470);
nor U3769 (N_3769,N_3491,N_3498);
or U3770 (N_3770,N_3589,N_3467);
and U3771 (N_3771,N_3414,N_3516);
and U3772 (N_3772,N_3506,N_3522);
and U3773 (N_3773,N_3482,N_3592);
xor U3774 (N_3774,N_3406,N_3400);
or U3775 (N_3775,N_3509,N_3489);
nor U3776 (N_3776,N_3496,N_3412);
nand U3777 (N_3777,N_3493,N_3405);
or U3778 (N_3778,N_3521,N_3424);
and U3779 (N_3779,N_3547,N_3412);
nor U3780 (N_3780,N_3444,N_3547);
nor U3781 (N_3781,N_3583,N_3466);
and U3782 (N_3782,N_3570,N_3560);
nand U3783 (N_3783,N_3434,N_3547);
or U3784 (N_3784,N_3518,N_3515);
or U3785 (N_3785,N_3549,N_3542);
and U3786 (N_3786,N_3444,N_3455);
or U3787 (N_3787,N_3523,N_3431);
and U3788 (N_3788,N_3554,N_3417);
or U3789 (N_3789,N_3462,N_3522);
nand U3790 (N_3790,N_3478,N_3524);
nand U3791 (N_3791,N_3552,N_3422);
nor U3792 (N_3792,N_3516,N_3475);
nand U3793 (N_3793,N_3556,N_3412);
and U3794 (N_3794,N_3434,N_3413);
and U3795 (N_3795,N_3566,N_3451);
or U3796 (N_3796,N_3490,N_3447);
nand U3797 (N_3797,N_3553,N_3443);
or U3798 (N_3798,N_3511,N_3461);
nand U3799 (N_3799,N_3504,N_3439);
or U3800 (N_3800,N_3772,N_3638);
nand U3801 (N_3801,N_3687,N_3719);
or U3802 (N_3802,N_3686,N_3761);
and U3803 (N_3803,N_3624,N_3621);
nor U3804 (N_3804,N_3737,N_3727);
or U3805 (N_3805,N_3721,N_3648);
xnor U3806 (N_3806,N_3789,N_3739);
or U3807 (N_3807,N_3752,N_3629);
or U3808 (N_3808,N_3601,N_3705);
and U3809 (N_3809,N_3707,N_3650);
nand U3810 (N_3810,N_3765,N_3643);
nand U3811 (N_3811,N_3791,N_3672);
or U3812 (N_3812,N_3794,N_3763);
or U3813 (N_3813,N_3704,N_3665);
nor U3814 (N_3814,N_3699,N_3793);
and U3815 (N_3815,N_3682,N_3634);
xnor U3816 (N_3816,N_3792,N_3779);
nand U3817 (N_3817,N_3742,N_3776);
nor U3818 (N_3818,N_3647,N_3735);
or U3819 (N_3819,N_3733,N_3713);
and U3820 (N_3820,N_3741,N_3784);
and U3821 (N_3821,N_3639,N_3782);
nand U3822 (N_3822,N_3659,N_3731);
xor U3823 (N_3823,N_3669,N_3680);
and U3824 (N_3824,N_3612,N_3717);
or U3825 (N_3825,N_3736,N_3746);
or U3826 (N_3826,N_3773,N_3732);
or U3827 (N_3827,N_3745,N_3694);
nand U3828 (N_3828,N_3786,N_3653);
nor U3829 (N_3829,N_3652,N_3649);
nor U3830 (N_3830,N_3718,N_3766);
nor U3831 (N_3831,N_3703,N_3693);
xor U3832 (N_3832,N_3657,N_3754);
nand U3833 (N_3833,N_3750,N_3645);
nand U3834 (N_3834,N_3668,N_3614);
nand U3835 (N_3835,N_3684,N_3767);
and U3836 (N_3836,N_3681,N_3613);
nand U3837 (N_3837,N_3799,N_3607);
or U3838 (N_3838,N_3685,N_3642);
nor U3839 (N_3839,N_3770,N_3637);
or U3840 (N_3840,N_3714,N_3683);
nand U3841 (N_3841,N_3723,N_3666);
nor U3842 (N_3842,N_3738,N_3603);
nor U3843 (N_3843,N_3796,N_3795);
and U3844 (N_3844,N_3679,N_3762);
nand U3845 (N_3845,N_3798,N_3768);
and U3846 (N_3846,N_3749,N_3744);
nor U3847 (N_3847,N_3753,N_3640);
and U3848 (N_3848,N_3774,N_3617);
and U3849 (N_3849,N_3604,N_3620);
nand U3850 (N_3850,N_3641,N_3778);
xnor U3851 (N_3851,N_3696,N_3663);
nor U3852 (N_3852,N_3654,N_3716);
nor U3853 (N_3853,N_3622,N_3726);
xor U3854 (N_3854,N_3671,N_3695);
nand U3855 (N_3855,N_3781,N_3655);
or U3856 (N_3856,N_3712,N_3709);
or U3857 (N_3857,N_3691,N_3673);
nor U3858 (N_3858,N_3698,N_3644);
or U3859 (N_3859,N_3785,N_3636);
nor U3860 (N_3860,N_3771,N_3780);
nor U3861 (N_3861,N_3783,N_3747);
nand U3862 (N_3862,N_3610,N_3740);
xnor U3863 (N_3863,N_3748,N_3720);
nor U3864 (N_3864,N_3700,N_3627);
nand U3865 (N_3865,N_3619,N_3674);
nand U3866 (N_3866,N_3630,N_3692);
and U3867 (N_3867,N_3715,N_3670);
nand U3868 (N_3868,N_3729,N_3600);
xnor U3869 (N_3869,N_3651,N_3758);
nor U3870 (N_3870,N_3756,N_3777);
or U3871 (N_3871,N_3608,N_3702);
or U3872 (N_3872,N_3730,N_3662);
nand U3873 (N_3873,N_3690,N_3743);
nor U3874 (N_3874,N_3646,N_3615);
nor U3875 (N_3875,N_3676,N_3759);
nand U3876 (N_3876,N_3701,N_3728);
or U3877 (N_3877,N_3688,N_3631);
or U3878 (N_3878,N_3618,N_3656);
and U3879 (N_3879,N_3769,N_3722);
or U3880 (N_3880,N_3626,N_3675);
and U3881 (N_3881,N_3788,N_3734);
xor U3882 (N_3882,N_3678,N_3706);
nor U3883 (N_3883,N_3664,N_3757);
nand U3884 (N_3884,N_3661,N_3724);
nand U3885 (N_3885,N_3611,N_3632);
or U3886 (N_3886,N_3797,N_3725);
or U3887 (N_3887,N_3606,N_3633);
xor U3888 (N_3888,N_3658,N_3764);
nand U3889 (N_3889,N_3635,N_3751);
or U3890 (N_3890,N_3697,N_3760);
and U3891 (N_3891,N_3625,N_3711);
or U3892 (N_3892,N_3628,N_3609);
nor U3893 (N_3893,N_3623,N_3708);
xnor U3894 (N_3894,N_3667,N_3755);
and U3895 (N_3895,N_3616,N_3605);
nor U3896 (N_3896,N_3677,N_3710);
nand U3897 (N_3897,N_3660,N_3775);
or U3898 (N_3898,N_3790,N_3602);
and U3899 (N_3899,N_3689,N_3787);
nand U3900 (N_3900,N_3618,N_3706);
nand U3901 (N_3901,N_3790,N_3631);
xnor U3902 (N_3902,N_3665,N_3768);
nor U3903 (N_3903,N_3723,N_3771);
and U3904 (N_3904,N_3713,N_3745);
nand U3905 (N_3905,N_3684,N_3668);
nor U3906 (N_3906,N_3713,N_3731);
or U3907 (N_3907,N_3692,N_3703);
or U3908 (N_3908,N_3631,N_3774);
or U3909 (N_3909,N_3715,N_3761);
nor U3910 (N_3910,N_3663,N_3642);
nor U3911 (N_3911,N_3712,N_3792);
or U3912 (N_3912,N_3771,N_3624);
nor U3913 (N_3913,N_3722,N_3611);
and U3914 (N_3914,N_3673,N_3767);
nand U3915 (N_3915,N_3646,N_3658);
and U3916 (N_3916,N_3716,N_3605);
and U3917 (N_3917,N_3756,N_3635);
or U3918 (N_3918,N_3697,N_3676);
and U3919 (N_3919,N_3615,N_3654);
nor U3920 (N_3920,N_3764,N_3627);
xnor U3921 (N_3921,N_3610,N_3675);
nand U3922 (N_3922,N_3632,N_3751);
and U3923 (N_3923,N_3751,N_3604);
or U3924 (N_3924,N_3677,N_3649);
and U3925 (N_3925,N_3778,N_3695);
nor U3926 (N_3926,N_3666,N_3663);
and U3927 (N_3927,N_3679,N_3670);
nand U3928 (N_3928,N_3791,N_3751);
nor U3929 (N_3929,N_3686,N_3649);
xnor U3930 (N_3930,N_3633,N_3784);
and U3931 (N_3931,N_3663,N_3619);
and U3932 (N_3932,N_3730,N_3796);
xor U3933 (N_3933,N_3782,N_3788);
nor U3934 (N_3934,N_3761,N_3792);
or U3935 (N_3935,N_3751,N_3731);
or U3936 (N_3936,N_3614,N_3636);
nand U3937 (N_3937,N_3796,N_3698);
nand U3938 (N_3938,N_3744,N_3659);
or U3939 (N_3939,N_3622,N_3699);
nor U3940 (N_3940,N_3652,N_3677);
nand U3941 (N_3941,N_3725,N_3778);
and U3942 (N_3942,N_3662,N_3750);
nor U3943 (N_3943,N_3609,N_3692);
and U3944 (N_3944,N_3710,N_3728);
and U3945 (N_3945,N_3715,N_3604);
and U3946 (N_3946,N_3642,N_3627);
nor U3947 (N_3947,N_3646,N_3766);
or U3948 (N_3948,N_3622,N_3646);
or U3949 (N_3949,N_3626,N_3750);
and U3950 (N_3950,N_3713,N_3786);
nand U3951 (N_3951,N_3601,N_3618);
xor U3952 (N_3952,N_3748,N_3753);
or U3953 (N_3953,N_3706,N_3717);
and U3954 (N_3954,N_3679,N_3629);
and U3955 (N_3955,N_3643,N_3695);
nor U3956 (N_3956,N_3702,N_3609);
nor U3957 (N_3957,N_3650,N_3636);
and U3958 (N_3958,N_3792,N_3737);
xnor U3959 (N_3959,N_3657,N_3760);
and U3960 (N_3960,N_3757,N_3632);
and U3961 (N_3961,N_3740,N_3778);
nand U3962 (N_3962,N_3646,N_3731);
nand U3963 (N_3963,N_3664,N_3792);
nand U3964 (N_3964,N_3752,N_3616);
or U3965 (N_3965,N_3733,N_3672);
or U3966 (N_3966,N_3672,N_3623);
nand U3967 (N_3967,N_3799,N_3786);
nor U3968 (N_3968,N_3708,N_3681);
and U3969 (N_3969,N_3740,N_3774);
and U3970 (N_3970,N_3729,N_3614);
nand U3971 (N_3971,N_3711,N_3795);
nand U3972 (N_3972,N_3647,N_3644);
or U3973 (N_3973,N_3776,N_3622);
or U3974 (N_3974,N_3708,N_3612);
or U3975 (N_3975,N_3719,N_3747);
nor U3976 (N_3976,N_3661,N_3670);
or U3977 (N_3977,N_3655,N_3784);
nor U3978 (N_3978,N_3729,N_3640);
nor U3979 (N_3979,N_3643,N_3769);
nor U3980 (N_3980,N_3631,N_3679);
xor U3981 (N_3981,N_3749,N_3748);
nand U3982 (N_3982,N_3799,N_3722);
nand U3983 (N_3983,N_3625,N_3719);
nor U3984 (N_3984,N_3672,N_3764);
nor U3985 (N_3985,N_3679,N_3613);
or U3986 (N_3986,N_3634,N_3749);
and U3987 (N_3987,N_3692,N_3684);
or U3988 (N_3988,N_3725,N_3670);
xor U3989 (N_3989,N_3681,N_3772);
nor U3990 (N_3990,N_3616,N_3700);
xnor U3991 (N_3991,N_3634,N_3778);
and U3992 (N_3992,N_3658,N_3779);
nand U3993 (N_3993,N_3648,N_3639);
xor U3994 (N_3994,N_3745,N_3692);
nor U3995 (N_3995,N_3642,N_3680);
or U3996 (N_3996,N_3686,N_3764);
nor U3997 (N_3997,N_3619,N_3754);
nor U3998 (N_3998,N_3687,N_3675);
nand U3999 (N_3999,N_3716,N_3639);
and U4000 (N_4000,N_3926,N_3897);
or U4001 (N_4001,N_3902,N_3915);
and U4002 (N_4002,N_3824,N_3983);
or U4003 (N_4003,N_3998,N_3858);
and U4004 (N_4004,N_3910,N_3865);
nor U4005 (N_4005,N_3900,N_3924);
or U4006 (N_4006,N_3906,N_3842);
or U4007 (N_4007,N_3934,N_3957);
or U4008 (N_4008,N_3937,N_3996);
nor U4009 (N_4009,N_3823,N_3953);
and U4010 (N_4010,N_3965,N_3839);
xor U4011 (N_4011,N_3829,N_3942);
nor U4012 (N_4012,N_3801,N_3978);
nor U4013 (N_4013,N_3859,N_3972);
and U4014 (N_4014,N_3994,N_3853);
nand U4015 (N_4015,N_3833,N_3952);
nand U4016 (N_4016,N_3964,N_3875);
xnor U4017 (N_4017,N_3886,N_3907);
and U4018 (N_4018,N_3830,N_3800);
nand U4019 (N_4019,N_3916,N_3845);
nand U4020 (N_4020,N_3922,N_3832);
or U4021 (N_4021,N_3914,N_3899);
and U4022 (N_4022,N_3966,N_3960);
and U4023 (N_4023,N_3822,N_3923);
xor U4024 (N_4024,N_3861,N_3955);
and U4025 (N_4025,N_3940,N_3939);
or U4026 (N_4026,N_3951,N_3993);
nor U4027 (N_4027,N_3873,N_3895);
or U4028 (N_4028,N_3918,N_3913);
and U4029 (N_4029,N_3811,N_3834);
nand U4030 (N_4030,N_3870,N_3809);
nand U4031 (N_4031,N_3981,N_3948);
and U4032 (N_4032,N_3864,N_3869);
xor U4033 (N_4033,N_3929,N_3888);
nand U4034 (N_4034,N_3896,N_3813);
and U4035 (N_4035,N_3825,N_3831);
nor U4036 (N_4036,N_3881,N_3961);
or U4037 (N_4037,N_3871,N_3905);
and U4038 (N_4038,N_3944,N_3962);
nor U4039 (N_4039,N_3927,N_3843);
xor U4040 (N_4040,N_3890,N_3912);
xnor U4041 (N_4041,N_3930,N_3821);
and U4042 (N_4042,N_3982,N_3936);
or U4043 (N_4043,N_3885,N_3959);
nand U4044 (N_4044,N_3874,N_3876);
xnor U4045 (N_4045,N_3815,N_3908);
and U4046 (N_4046,N_3851,N_3891);
and U4047 (N_4047,N_3928,N_3878);
nand U4048 (N_4048,N_3999,N_3806);
nor U4049 (N_4049,N_3904,N_3932);
or U4050 (N_4050,N_3975,N_3812);
and U4051 (N_4051,N_3894,N_3958);
nor U4052 (N_4052,N_3803,N_3956);
nor U4053 (N_4053,N_3986,N_3802);
nor U4054 (N_4054,N_3884,N_3849);
and U4055 (N_4055,N_3840,N_3992);
nor U4056 (N_4056,N_3968,N_3987);
nor U4057 (N_4057,N_3827,N_3826);
and U4058 (N_4058,N_3847,N_3893);
xor U4059 (N_4059,N_3921,N_3971);
nor U4060 (N_4060,N_3963,N_3804);
nor U4061 (N_4061,N_3938,N_3828);
or U4062 (N_4062,N_3855,N_3985);
nand U4063 (N_4063,N_3898,N_3860);
or U4064 (N_4064,N_3988,N_3920);
xnor U4065 (N_4065,N_3941,N_3903);
nand U4066 (N_4066,N_3950,N_3817);
and U4067 (N_4067,N_3933,N_3877);
nor U4068 (N_4068,N_3969,N_3814);
and U4069 (N_4069,N_3970,N_3967);
nand U4070 (N_4070,N_3810,N_3846);
and U4071 (N_4071,N_3889,N_3883);
and U4072 (N_4072,N_3838,N_3977);
nand U4073 (N_4073,N_3837,N_3819);
or U4074 (N_4074,N_3880,N_3945);
or U4075 (N_4075,N_3867,N_3989);
and U4076 (N_4076,N_3997,N_3820);
nor U4077 (N_4077,N_3863,N_3943);
nand U4078 (N_4078,N_3807,N_3974);
or U4079 (N_4079,N_3879,N_3976);
nor U4080 (N_4080,N_3946,N_3841);
or U4081 (N_4081,N_3844,N_3835);
or U4082 (N_4082,N_3995,N_3954);
nor U4083 (N_4083,N_3808,N_3836);
and U4084 (N_4084,N_3991,N_3848);
nor U4085 (N_4085,N_3850,N_3949);
nand U4086 (N_4086,N_3917,N_3892);
nand U4087 (N_4087,N_3980,N_3857);
and U4088 (N_4088,N_3852,N_3947);
nor U4089 (N_4089,N_3856,N_3911);
xnor U4090 (N_4090,N_3901,N_3925);
xor U4091 (N_4091,N_3872,N_3935);
and U4092 (N_4092,N_3862,N_3816);
or U4093 (N_4093,N_3984,N_3931);
and U4094 (N_4094,N_3919,N_3990);
xnor U4095 (N_4095,N_3887,N_3973);
and U4096 (N_4096,N_3805,N_3854);
xnor U4097 (N_4097,N_3979,N_3882);
nand U4098 (N_4098,N_3868,N_3866);
nor U4099 (N_4099,N_3818,N_3909);
nor U4100 (N_4100,N_3849,N_3853);
nand U4101 (N_4101,N_3832,N_3816);
and U4102 (N_4102,N_3899,N_3950);
or U4103 (N_4103,N_3865,N_3813);
nand U4104 (N_4104,N_3946,N_3807);
or U4105 (N_4105,N_3885,N_3900);
nand U4106 (N_4106,N_3818,N_3978);
or U4107 (N_4107,N_3867,N_3962);
nand U4108 (N_4108,N_3927,N_3920);
or U4109 (N_4109,N_3843,N_3975);
and U4110 (N_4110,N_3854,N_3912);
and U4111 (N_4111,N_3981,N_3970);
or U4112 (N_4112,N_3897,N_3854);
or U4113 (N_4113,N_3942,N_3884);
nand U4114 (N_4114,N_3948,N_3852);
and U4115 (N_4115,N_3881,N_3885);
nand U4116 (N_4116,N_3830,N_3959);
xor U4117 (N_4117,N_3929,N_3850);
and U4118 (N_4118,N_3924,N_3995);
nand U4119 (N_4119,N_3886,N_3964);
and U4120 (N_4120,N_3830,N_3813);
nand U4121 (N_4121,N_3955,N_3939);
or U4122 (N_4122,N_3940,N_3834);
nor U4123 (N_4123,N_3958,N_3839);
nor U4124 (N_4124,N_3808,N_3943);
xor U4125 (N_4125,N_3803,N_3889);
and U4126 (N_4126,N_3938,N_3870);
and U4127 (N_4127,N_3840,N_3963);
nand U4128 (N_4128,N_3821,N_3807);
and U4129 (N_4129,N_3927,N_3959);
nor U4130 (N_4130,N_3926,N_3816);
nand U4131 (N_4131,N_3970,N_3937);
xnor U4132 (N_4132,N_3959,N_3812);
nand U4133 (N_4133,N_3988,N_3899);
nand U4134 (N_4134,N_3912,N_3866);
and U4135 (N_4135,N_3827,N_3942);
and U4136 (N_4136,N_3908,N_3904);
nor U4137 (N_4137,N_3951,N_3994);
or U4138 (N_4138,N_3876,N_3858);
and U4139 (N_4139,N_3833,N_3894);
nand U4140 (N_4140,N_3946,N_3842);
and U4141 (N_4141,N_3850,N_3864);
nand U4142 (N_4142,N_3883,N_3870);
or U4143 (N_4143,N_3803,N_3918);
or U4144 (N_4144,N_3849,N_3938);
nand U4145 (N_4145,N_3892,N_3925);
nand U4146 (N_4146,N_3983,N_3942);
nand U4147 (N_4147,N_3936,N_3887);
nor U4148 (N_4148,N_3910,N_3971);
xor U4149 (N_4149,N_3811,N_3868);
nand U4150 (N_4150,N_3836,N_3956);
or U4151 (N_4151,N_3814,N_3911);
xor U4152 (N_4152,N_3952,N_3899);
xor U4153 (N_4153,N_3852,N_3963);
nand U4154 (N_4154,N_3821,N_3819);
nand U4155 (N_4155,N_3855,N_3931);
xor U4156 (N_4156,N_3887,N_3874);
nand U4157 (N_4157,N_3853,N_3851);
nor U4158 (N_4158,N_3899,N_3922);
or U4159 (N_4159,N_3960,N_3888);
or U4160 (N_4160,N_3911,N_3969);
nor U4161 (N_4161,N_3919,N_3878);
or U4162 (N_4162,N_3983,N_3982);
nand U4163 (N_4163,N_3955,N_3953);
or U4164 (N_4164,N_3859,N_3839);
nor U4165 (N_4165,N_3950,N_3900);
xnor U4166 (N_4166,N_3986,N_3899);
and U4167 (N_4167,N_3846,N_3844);
or U4168 (N_4168,N_3846,N_3907);
and U4169 (N_4169,N_3819,N_3964);
nand U4170 (N_4170,N_3802,N_3809);
or U4171 (N_4171,N_3977,N_3856);
and U4172 (N_4172,N_3892,N_3883);
and U4173 (N_4173,N_3883,N_3962);
and U4174 (N_4174,N_3901,N_3942);
and U4175 (N_4175,N_3870,N_3810);
nand U4176 (N_4176,N_3966,N_3930);
and U4177 (N_4177,N_3844,N_3916);
and U4178 (N_4178,N_3857,N_3806);
nand U4179 (N_4179,N_3918,N_3819);
nor U4180 (N_4180,N_3844,N_3994);
nand U4181 (N_4181,N_3920,N_3917);
nor U4182 (N_4182,N_3894,N_3943);
nand U4183 (N_4183,N_3834,N_3977);
xor U4184 (N_4184,N_3933,N_3880);
nor U4185 (N_4185,N_3890,N_3913);
nand U4186 (N_4186,N_3960,N_3997);
nand U4187 (N_4187,N_3911,N_3888);
or U4188 (N_4188,N_3817,N_3887);
or U4189 (N_4189,N_3850,N_3966);
xnor U4190 (N_4190,N_3908,N_3828);
or U4191 (N_4191,N_3894,N_3851);
nand U4192 (N_4192,N_3981,N_3846);
or U4193 (N_4193,N_3881,N_3934);
and U4194 (N_4194,N_3963,N_3901);
nand U4195 (N_4195,N_3911,N_3980);
or U4196 (N_4196,N_3936,N_3832);
or U4197 (N_4197,N_3881,N_3827);
nand U4198 (N_4198,N_3872,N_3850);
or U4199 (N_4199,N_3932,N_3906);
and U4200 (N_4200,N_4105,N_4034);
xnor U4201 (N_4201,N_4019,N_4135);
xor U4202 (N_4202,N_4077,N_4024);
and U4203 (N_4203,N_4130,N_4061);
and U4204 (N_4204,N_4088,N_4147);
nor U4205 (N_4205,N_4154,N_4109);
and U4206 (N_4206,N_4094,N_4033);
or U4207 (N_4207,N_4055,N_4100);
or U4208 (N_4208,N_4184,N_4148);
nand U4209 (N_4209,N_4045,N_4058);
nand U4210 (N_4210,N_4008,N_4004);
nand U4211 (N_4211,N_4095,N_4129);
and U4212 (N_4212,N_4062,N_4196);
nor U4213 (N_4213,N_4082,N_4149);
nor U4214 (N_4214,N_4025,N_4028);
and U4215 (N_4215,N_4066,N_4150);
nor U4216 (N_4216,N_4153,N_4116);
and U4217 (N_4217,N_4040,N_4132);
nand U4218 (N_4218,N_4039,N_4113);
or U4219 (N_4219,N_4070,N_4133);
and U4220 (N_4220,N_4178,N_4051);
nand U4221 (N_4221,N_4089,N_4050);
nand U4222 (N_4222,N_4111,N_4176);
or U4223 (N_4223,N_4097,N_4117);
nor U4224 (N_4224,N_4092,N_4005);
and U4225 (N_4225,N_4120,N_4106);
nand U4226 (N_4226,N_4158,N_4027);
nand U4227 (N_4227,N_4191,N_4142);
nand U4228 (N_4228,N_4122,N_4166);
nor U4229 (N_4229,N_4143,N_4084);
nor U4230 (N_4230,N_4074,N_4046);
nand U4231 (N_4231,N_4198,N_4096);
nand U4232 (N_4232,N_4038,N_4003);
xnor U4233 (N_4233,N_4169,N_4114);
nand U4234 (N_4234,N_4014,N_4128);
xnor U4235 (N_4235,N_4190,N_4011);
nand U4236 (N_4236,N_4110,N_4002);
xnor U4237 (N_4237,N_4031,N_4118);
xnor U4238 (N_4238,N_4192,N_4049);
nand U4239 (N_4239,N_4020,N_4104);
nand U4240 (N_4240,N_4081,N_4163);
and U4241 (N_4241,N_4021,N_4013);
or U4242 (N_4242,N_4199,N_4015);
or U4243 (N_4243,N_4182,N_4123);
nor U4244 (N_4244,N_4065,N_4093);
and U4245 (N_4245,N_4102,N_4072);
nand U4246 (N_4246,N_4187,N_4141);
and U4247 (N_4247,N_4175,N_4159);
and U4248 (N_4248,N_4193,N_4168);
and U4249 (N_4249,N_4060,N_4157);
nand U4250 (N_4250,N_4010,N_4047);
and U4251 (N_4251,N_4054,N_4037);
and U4252 (N_4252,N_4006,N_4181);
nand U4253 (N_4253,N_4016,N_4067);
or U4254 (N_4254,N_4185,N_4017);
xor U4255 (N_4255,N_4155,N_4091);
nand U4256 (N_4256,N_4108,N_4156);
and U4257 (N_4257,N_4085,N_4167);
and U4258 (N_4258,N_4194,N_4195);
nand U4259 (N_4259,N_4151,N_4023);
nor U4260 (N_4260,N_4101,N_4022);
xnor U4261 (N_4261,N_4087,N_4057);
and U4262 (N_4262,N_4107,N_4145);
or U4263 (N_4263,N_4090,N_4086);
nor U4264 (N_4264,N_4007,N_4030);
nand U4265 (N_4265,N_4121,N_4079);
nand U4266 (N_4266,N_4165,N_4078);
and U4267 (N_4267,N_4140,N_4063);
and U4268 (N_4268,N_4146,N_4075);
xnor U4269 (N_4269,N_4161,N_4009);
or U4270 (N_4270,N_4173,N_4071);
and U4271 (N_4271,N_4069,N_4152);
nand U4272 (N_4272,N_4127,N_4180);
nor U4273 (N_4273,N_4026,N_4197);
nand U4274 (N_4274,N_4174,N_4125);
xnor U4275 (N_4275,N_4001,N_4043);
or U4276 (N_4276,N_4183,N_4073);
nand U4277 (N_4277,N_4018,N_4172);
nand U4278 (N_4278,N_4000,N_4144);
xnor U4279 (N_4279,N_4080,N_4126);
and U4280 (N_4280,N_4056,N_4099);
and U4281 (N_4281,N_4068,N_4032);
xnor U4282 (N_4282,N_4171,N_4137);
nor U4283 (N_4283,N_4083,N_4115);
nor U4284 (N_4284,N_4136,N_4124);
or U4285 (N_4285,N_4138,N_4012);
nand U4286 (N_4286,N_4042,N_4064);
nor U4287 (N_4287,N_4131,N_4052);
nand U4288 (N_4288,N_4162,N_4053);
nand U4289 (N_4289,N_4188,N_4164);
or U4290 (N_4290,N_4029,N_4035);
nor U4291 (N_4291,N_4177,N_4160);
or U4292 (N_4292,N_4076,N_4036);
or U4293 (N_4293,N_4059,N_4041);
nor U4294 (N_4294,N_4098,N_4048);
xnor U4295 (N_4295,N_4170,N_4189);
and U4296 (N_4296,N_4134,N_4112);
nand U4297 (N_4297,N_4119,N_4139);
nor U4298 (N_4298,N_4103,N_4186);
nand U4299 (N_4299,N_4179,N_4044);
nor U4300 (N_4300,N_4082,N_4061);
and U4301 (N_4301,N_4089,N_4083);
and U4302 (N_4302,N_4122,N_4198);
xnor U4303 (N_4303,N_4006,N_4081);
nand U4304 (N_4304,N_4084,N_4064);
and U4305 (N_4305,N_4171,N_4186);
nor U4306 (N_4306,N_4199,N_4050);
nand U4307 (N_4307,N_4173,N_4043);
nand U4308 (N_4308,N_4158,N_4016);
or U4309 (N_4309,N_4038,N_4184);
nor U4310 (N_4310,N_4039,N_4121);
or U4311 (N_4311,N_4129,N_4134);
xnor U4312 (N_4312,N_4067,N_4132);
nand U4313 (N_4313,N_4064,N_4153);
nand U4314 (N_4314,N_4095,N_4167);
nand U4315 (N_4315,N_4150,N_4127);
or U4316 (N_4316,N_4059,N_4132);
nand U4317 (N_4317,N_4048,N_4198);
or U4318 (N_4318,N_4044,N_4174);
nand U4319 (N_4319,N_4126,N_4043);
or U4320 (N_4320,N_4105,N_4179);
or U4321 (N_4321,N_4070,N_4180);
and U4322 (N_4322,N_4082,N_4064);
xnor U4323 (N_4323,N_4046,N_4050);
xnor U4324 (N_4324,N_4162,N_4035);
or U4325 (N_4325,N_4024,N_4110);
and U4326 (N_4326,N_4082,N_4035);
nand U4327 (N_4327,N_4192,N_4104);
nor U4328 (N_4328,N_4118,N_4122);
nor U4329 (N_4329,N_4086,N_4183);
or U4330 (N_4330,N_4195,N_4116);
nand U4331 (N_4331,N_4128,N_4079);
nor U4332 (N_4332,N_4149,N_4133);
nor U4333 (N_4333,N_4040,N_4009);
nand U4334 (N_4334,N_4004,N_4022);
or U4335 (N_4335,N_4124,N_4097);
nand U4336 (N_4336,N_4065,N_4146);
or U4337 (N_4337,N_4140,N_4170);
nand U4338 (N_4338,N_4061,N_4014);
and U4339 (N_4339,N_4058,N_4101);
or U4340 (N_4340,N_4163,N_4024);
xnor U4341 (N_4341,N_4072,N_4132);
nor U4342 (N_4342,N_4148,N_4155);
and U4343 (N_4343,N_4126,N_4026);
and U4344 (N_4344,N_4001,N_4057);
and U4345 (N_4345,N_4105,N_4092);
nor U4346 (N_4346,N_4182,N_4190);
nand U4347 (N_4347,N_4005,N_4032);
or U4348 (N_4348,N_4165,N_4144);
nand U4349 (N_4349,N_4194,N_4052);
nand U4350 (N_4350,N_4194,N_4111);
nor U4351 (N_4351,N_4029,N_4092);
or U4352 (N_4352,N_4173,N_4136);
and U4353 (N_4353,N_4111,N_4007);
and U4354 (N_4354,N_4122,N_4026);
nor U4355 (N_4355,N_4096,N_4187);
or U4356 (N_4356,N_4038,N_4082);
nor U4357 (N_4357,N_4195,N_4020);
nor U4358 (N_4358,N_4157,N_4175);
or U4359 (N_4359,N_4142,N_4037);
or U4360 (N_4360,N_4151,N_4165);
nor U4361 (N_4361,N_4084,N_4187);
nor U4362 (N_4362,N_4075,N_4041);
or U4363 (N_4363,N_4170,N_4116);
and U4364 (N_4364,N_4123,N_4098);
or U4365 (N_4365,N_4134,N_4000);
xor U4366 (N_4366,N_4173,N_4036);
or U4367 (N_4367,N_4164,N_4127);
and U4368 (N_4368,N_4031,N_4040);
nor U4369 (N_4369,N_4089,N_4173);
or U4370 (N_4370,N_4142,N_4107);
or U4371 (N_4371,N_4085,N_4029);
nor U4372 (N_4372,N_4040,N_4120);
or U4373 (N_4373,N_4011,N_4161);
and U4374 (N_4374,N_4139,N_4164);
nor U4375 (N_4375,N_4075,N_4130);
and U4376 (N_4376,N_4127,N_4183);
xor U4377 (N_4377,N_4128,N_4091);
and U4378 (N_4378,N_4057,N_4050);
nor U4379 (N_4379,N_4069,N_4161);
nand U4380 (N_4380,N_4091,N_4081);
or U4381 (N_4381,N_4109,N_4085);
nand U4382 (N_4382,N_4082,N_4012);
and U4383 (N_4383,N_4000,N_4087);
nor U4384 (N_4384,N_4176,N_4135);
nand U4385 (N_4385,N_4153,N_4107);
or U4386 (N_4386,N_4028,N_4111);
nand U4387 (N_4387,N_4033,N_4104);
and U4388 (N_4388,N_4172,N_4081);
or U4389 (N_4389,N_4040,N_4057);
and U4390 (N_4390,N_4039,N_4125);
nand U4391 (N_4391,N_4093,N_4000);
nand U4392 (N_4392,N_4089,N_4121);
xor U4393 (N_4393,N_4041,N_4032);
nand U4394 (N_4394,N_4164,N_4198);
nand U4395 (N_4395,N_4045,N_4071);
nor U4396 (N_4396,N_4177,N_4133);
and U4397 (N_4397,N_4185,N_4035);
nor U4398 (N_4398,N_4177,N_4060);
or U4399 (N_4399,N_4113,N_4189);
and U4400 (N_4400,N_4269,N_4260);
nor U4401 (N_4401,N_4369,N_4388);
or U4402 (N_4402,N_4257,N_4237);
nand U4403 (N_4403,N_4389,N_4392);
xor U4404 (N_4404,N_4292,N_4227);
nand U4405 (N_4405,N_4295,N_4353);
nor U4406 (N_4406,N_4359,N_4309);
nor U4407 (N_4407,N_4219,N_4299);
xor U4408 (N_4408,N_4396,N_4391);
nor U4409 (N_4409,N_4339,N_4221);
xnor U4410 (N_4410,N_4246,N_4349);
nand U4411 (N_4411,N_4267,N_4297);
nor U4412 (N_4412,N_4387,N_4384);
nand U4413 (N_4413,N_4264,N_4208);
nor U4414 (N_4414,N_4371,N_4254);
nand U4415 (N_4415,N_4215,N_4320);
or U4416 (N_4416,N_4271,N_4235);
nor U4417 (N_4417,N_4212,N_4368);
nand U4418 (N_4418,N_4285,N_4201);
nand U4419 (N_4419,N_4251,N_4231);
nor U4420 (N_4420,N_4335,N_4329);
or U4421 (N_4421,N_4307,N_4274);
nor U4422 (N_4422,N_4317,N_4358);
and U4423 (N_4423,N_4310,N_4284);
nor U4424 (N_4424,N_4261,N_4362);
nor U4425 (N_4425,N_4318,N_4398);
nand U4426 (N_4426,N_4298,N_4390);
or U4427 (N_4427,N_4313,N_4345);
nand U4428 (N_4428,N_4370,N_4289);
or U4429 (N_4429,N_4355,N_4294);
nor U4430 (N_4430,N_4203,N_4346);
xnor U4431 (N_4431,N_4375,N_4385);
nor U4432 (N_4432,N_4305,N_4393);
or U4433 (N_4433,N_4249,N_4342);
xor U4434 (N_4434,N_4331,N_4250);
nand U4435 (N_4435,N_4248,N_4364);
nor U4436 (N_4436,N_4363,N_4340);
or U4437 (N_4437,N_4236,N_4281);
nand U4438 (N_4438,N_4334,N_4316);
nand U4439 (N_4439,N_4376,N_4347);
nor U4440 (N_4440,N_4226,N_4330);
nand U4441 (N_4441,N_4399,N_4224);
nand U4442 (N_4442,N_4210,N_4296);
or U4443 (N_4443,N_4379,N_4301);
or U4444 (N_4444,N_4366,N_4277);
nor U4445 (N_4445,N_4238,N_4360);
or U4446 (N_4446,N_4243,N_4397);
and U4447 (N_4447,N_4252,N_4288);
nor U4448 (N_4448,N_4382,N_4328);
and U4449 (N_4449,N_4381,N_4282);
and U4450 (N_4450,N_4365,N_4314);
nor U4451 (N_4451,N_4200,N_4280);
nand U4452 (N_4452,N_4202,N_4325);
and U4453 (N_4453,N_4265,N_4279);
nor U4454 (N_4454,N_4204,N_4290);
nor U4455 (N_4455,N_4270,N_4321);
nand U4456 (N_4456,N_4256,N_4312);
and U4457 (N_4457,N_4278,N_4383);
or U4458 (N_4458,N_4259,N_4332);
nor U4459 (N_4459,N_4268,N_4263);
nor U4460 (N_4460,N_4209,N_4293);
or U4461 (N_4461,N_4344,N_4300);
nor U4462 (N_4462,N_4239,N_4304);
nor U4463 (N_4463,N_4234,N_4386);
and U4464 (N_4464,N_4374,N_4218);
and U4465 (N_4465,N_4241,N_4242);
xor U4466 (N_4466,N_4306,N_4354);
nand U4467 (N_4467,N_4207,N_4222);
nor U4468 (N_4468,N_4205,N_4244);
nor U4469 (N_4469,N_4394,N_4333);
xnor U4470 (N_4470,N_4327,N_4258);
nor U4471 (N_4471,N_4230,N_4276);
and U4472 (N_4472,N_4367,N_4395);
nor U4473 (N_4473,N_4211,N_4377);
nor U4474 (N_4474,N_4273,N_4206);
or U4475 (N_4475,N_4357,N_4351);
nand U4476 (N_4476,N_4315,N_4233);
nand U4477 (N_4477,N_4380,N_4308);
xor U4478 (N_4478,N_4240,N_4286);
or U4479 (N_4479,N_4223,N_4356);
and U4480 (N_4480,N_4266,N_4303);
xor U4481 (N_4481,N_4361,N_4378);
and U4482 (N_4482,N_4311,N_4228);
and U4483 (N_4483,N_4275,N_4336);
and U4484 (N_4484,N_4287,N_4319);
nand U4485 (N_4485,N_4341,N_4372);
nand U4486 (N_4486,N_4283,N_4220);
and U4487 (N_4487,N_4216,N_4302);
and U4488 (N_4488,N_4350,N_4291);
or U4489 (N_4489,N_4338,N_4255);
and U4490 (N_4490,N_4229,N_4373);
and U4491 (N_4491,N_4245,N_4326);
and U4492 (N_4492,N_4214,N_4322);
nand U4493 (N_4493,N_4232,N_4343);
nor U4494 (N_4494,N_4272,N_4348);
nand U4495 (N_4495,N_4262,N_4253);
nor U4496 (N_4496,N_4213,N_4217);
and U4497 (N_4497,N_4337,N_4225);
or U4498 (N_4498,N_4323,N_4324);
nor U4499 (N_4499,N_4352,N_4247);
xnor U4500 (N_4500,N_4385,N_4337);
and U4501 (N_4501,N_4364,N_4305);
and U4502 (N_4502,N_4351,N_4290);
or U4503 (N_4503,N_4231,N_4254);
nor U4504 (N_4504,N_4255,N_4217);
or U4505 (N_4505,N_4294,N_4335);
and U4506 (N_4506,N_4344,N_4271);
and U4507 (N_4507,N_4329,N_4320);
nor U4508 (N_4508,N_4281,N_4274);
and U4509 (N_4509,N_4331,N_4278);
and U4510 (N_4510,N_4298,N_4273);
and U4511 (N_4511,N_4200,N_4370);
or U4512 (N_4512,N_4287,N_4282);
and U4513 (N_4513,N_4203,N_4359);
or U4514 (N_4514,N_4334,N_4222);
nor U4515 (N_4515,N_4308,N_4328);
nor U4516 (N_4516,N_4356,N_4261);
nor U4517 (N_4517,N_4343,N_4200);
nand U4518 (N_4518,N_4351,N_4307);
or U4519 (N_4519,N_4271,N_4338);
nand U4520 (N_4520,N_4204,N_4296);
nand U4521 (N_4521,N_4272,N_4358);
nand U4522 (N_4522,N_4302,N_4256);
xor U4523 (N_4523,N_4387,N_4353);
xor U4524 (N_4524,N_4201,N_4207);
or U4525 (N_4525,N_4341,N_4274);
or U4526 (N_4526,N_4228,N_4232);
and U4527 (N_4527,N_4374,N_4303);
or U4528 (N_4528,N_4252,N_4306);
and U4529 (N_4529,N_4285,N_4394);
nand U4530 (N_4530,N_4365,N_4306);
or U4531 (N_4531,N_4336,N_4292);
nor U4532 (N_4532,N_4367,N_4365);
or U4533 (N_4533,N_4222,N_4244);
nand U4534 (N_4534,N_4251,N_4233);
xnor U4535 (N_4535,N_4221,N_4280);
nand U4536 (N_4536,N_4266,N_4260);
nand U4537 (N_4537,N_4349,N_4279);
or U4538 (N_4538,N_4385,N_4267);
nor U4539 (N_4539,N_4246,N_4260);
and U4540 (N_4540,N_4231,N_4220);
nor U4541 (N_4541,N_4292,N_4229);
or U4542 (N_4542,N_4340,N_4389);
nor U4543 (N_4543,N_4382,N_4393);
and U4544 (N_4544,N_4213,N_4392);
nand U4545 (N_4545,N_4215,N_4255);
nor U4546 (N_4546,N_4265,N_4344);
nor U4547 (N_4547,N_4372,N_4232);
nor U4548 (N_4548,N_4338,N_4254);
nand U4549 (N_4549,N_4397,N_4364);
xnor U4550 (N_4550,N_4393,N_4392);
nor U4551 (N_4551,N_4262,N_4377);
or U4552 (N_4552,N_4207,N_4232);
nor U4553 (N_4553,N_4291,N_4264);
nor U4554 (N_4554,N_4206,N_4326);
and U4555 (N_4555,N_4201,N_4366);
and U4556 (N_4556,N_4295,N_4304);
xnor U4557 (N_4557,N_4201,N_4264);
nand U4558 (N_4558,N_4237,N_4287);
nand U4559 (N_4559,N_4324,N_4357);
or U4560 (N_4560,N_4399,N_4203);
nand U4561 (N_4561,N_4250,N_4370);
nand U4562 (N_4562,N_4306,N_4231);
nand U4563 (N_4563,N_4341,N_4394);
nor U4564 (N_4564,N_4281,N_4336);
and U4565 (N_4565,N_4284,N_4210);
and U4566 (N_4566,N_4312,N_4391);
nand U4567 (N_4567,N_4236,N_4367);
or U4568 (N_4568,N_4274,N_4378);
nand U4569 (N_4569,N_4325,N_4205);
xor U4570 (N_4570,N_4362,N_4274);
nand U4571 (N_4571,N_4288,N_4243);
and U4572 (N_4572,N_4271,N_4239);
nand U4573 (N_4573,N_4206,N_4237);
or U4574 (N_4574,N_4375,N_4242);
or U4575 (N_4575,N_4328,N_4359);
nor U4576 (N_4576,N_4282,N_4380);
and U4577 (N_4577,N_4324,N_4222);
or U4578 (N_4578,N_4263,N_4221);
nand U4579 (N_4579,N_4382,N_4325);
xor U4580 (N_4580,N_4256,N_4200);
nand U4581 (N_4581,N_4330,N_4218);
nand U4582 (N_4582,N_4202,N_4223);
nor U4583 (N_4583,N_4363,N_4253);
and U4584 (N_4584,N_4385,N_4380);
nand U4585 (N_4585,N_4328,N_4237);
xor U4586 (N_4586,N_4235,N_4357);
and U4587 (N_4587,N_4219,N_4354);
nor U4588 (N_4588,N_4309,N_4274);
nand U4589 (N_4589,N_4236,N_4387);
xor U4590 (N_4590,N_4324,N_4361);
nor U4591 (N_4591,N_4368,N_4375);
xnor U4592 (N_4592,N_4370,N_4237);
xnor U4593 (N_4593,N_4284,N_4389);
and U4594 (N_4594,N_4202,N_4347);
or U4595 (N_4595,N_4285,N_4211);
and U4596 (N_4596,N_4375,N_4224);
or U4597 (N_4597,N_4317,N_4379);
xor U4598 (N_4598,N_4303,N_4313);
nand U4599 (N_4599,N_4262,N_4280);
nor U4600 (N_4600,N_4414,N_4513);
nor U4601 (N_4601,N_4444,N_4450);
nor U4602 (N_4602,N_4406,N_4562);
nor U4603 (N_4603,N_4595,N_4531);
or U4604 (N_4604,N_4544,N_4465);
and U4605 (N_4605,N_4476,N_4539);
nor U4606 (N_4606,N_4434,N_4564);
or U4607 (N_4607,N_4578,N_4538);
xnor U4608 (N_4608,N_4587,N_4400);
or U4609 (N_4609,N_4556,N_4520);
or U4610 (N_4610,N_4479,N_4448);
nor U4611 (N_4611,N_4483,N_4436);
nor U4612 (N_4612,N_4557,N_4464);
nor U4613 (N_4613,N_4484,N_4472);
nand U4614 (N_4614,N_4516,N_4559);
or U4615 (N_4615,N_4519,N_4521);
nand U4616 (N_4616,N_4478,N_4586);
xor U4617 (N_4617,N_4552,N_4443);
or U4618 (N_4618,N_4504,N_4423);
nor U4619 (N_4619,N_4553,N_4439);
nor U4620 (N_4620,N_4433,N_4402);
or U4621 (N_4621,N_4512,N_4525);
nand U4622 (N_4622,N_4575,N_4583);
nor U4623 (N_4623,N_4530,N_4452);
or U4624 (N_4624,N_4473,N_4415);
nor U4625 (N_4625,N_4574,N_4487);
nor U4626 (N_4626,N_4593,N_4486);
nand U4627 (N_4627,N_4485,N_4580);
and U4628 (N_4628,N_4555,N_4458);
xnor U4629 (N_4629,N_4418,N_4515);
nand U4630 (N_4630,N_4475,N_4568);
or U4631 (N_4631,N_4505,N_4528);
and U4632 (N_4632,N_4427,N_4592);
nand U4633 (N_4633,N_4577,N_4469);
nand U4634 (N_4634,N_4529,N_4491);
xnor U4635 (N_4635,N_4492,N_4554);
and U4636 (N_4636,N_4503,N_4590);
nor U4637 (N_4637,N_4569,N_4498);
nand U4638 (N_4638,N_4488,N_4417);
and U4639 (N_4639,N_4468,N_4424);
and U4640 (N_4640,N_4445,N_4596);
or U4641 (N_4641,N_4548,N_4533);
nand U4642 (N_4642,N_4407,N_4409);
and U4643 (N_4643,N_4584,N_4566);
xor U4644 (N_4644,N_4496,N_4435);
and U4645 (N_4645,N_4411,N_4534);
and U4646 (N_4646,N_4489,N_4514);
or U4647 (N_4647,N_4510,N_4535);
and U4648 (N_4648,N_4573,N_4471);
xnor U4649 (N_4649,N_4536,N_4599);
or U4650 (N_4650,N_4502,N_4432);
or U4651 (N_4651,N_4522,N_4412);
xor U4652 (N_4652,N_4497,N_4560);
or U4653 (N_4653,N_4511,N_4563);
nand U4654 (N_4654,N_4466,N_4547);
nand U4655 (N_4655,N_4526,N_4565);
and U4656 (N_4656,N_4572,N_4570);
or U4657 (N_4657,N_4426,N_4542);
nand U4658 (N_4658,N_4591,N_4493);
and U4659 (N_4659,N_4405,N_4500);
and U4660 (N_4660,N_4431,N_4550);
and U4661 (N_4661,N_4518,N_4567);
xor U4662 (N_4662,N_4545,N_4467);
nor U4663 (N_4663,N_4410,N_4437);
and U4664 (N_4664,N_4480,N_4456);
nor U4665 (N_4665,N_4549,N_4442);
or U4666 (N_4666,N_4527,N_4541);
or U4667 (N_4667,N_4585,N_4453);
nor U4668 (N_4668,N_4546,N_4509);
nand U4669 (N_4669,N_4455,N_4447);
and U4670 (N_4670,N_4576,N_4501);
or U4671 (N_4671,N_4579,N_4451);
or U4672 (N_4672,N_4462,N_4499);
nor U4673 (N_4673,N_4446,N_4403);
or U4674 (N_4674,N_4532,N_4494);
nor U4675 (N_4675,N_4428,N_4598);
and U4676 (N_4676,N_4463,N_4477);
or U4677 (N_4677,N_4495,N_4401);
and U4678 (N_4678,N_4408,N_4440);
nand U4679 (N_4679,N_4419,N_4507);
nor U4680 (N_4680,N_4438,N_4490);
and U4681 (N_4681,N_4404,N_4508);
nor U4682 (N_4682,N_4537,N_4416);
or U4683 (N_4683,N_4430,N_4524);
nor U4684 (N_4684,N_4459,N_4594);
and U4685 (N_4685,N_4589,N_4581);
nor U4686 (N_4686,N_4481,N_4454);
and U4687 (N_4687,N_4470,N_4429);
nand U4688 (N_4688,N_4597,N_4457);
or U4689 (N_4689,N_4517,N_4543);
nor U4690 (N_4690,N_4482,N_4441);
nand U4691 (N_4691,N_4474,N_4540);
and U4692 (N_4692,N_4461,N_4551);
xor U4693 (N_4693,N_4425,N_4561);
nand U4694 (N_4694,N_4420,N_4413);
or U4695 (N_4695,N_4571,N_4506);
nor U4696 (N_4696,N_4449,N_4588);
nand U4697 (N_4697,N_4460,N_4421);
nor U4698 (N_4698,N_4582,N_4422);
nor U4699 (N_4699,N_4523,N_4558);
and U4700 (N_4700,N_4461,N_4451);
nor U4701 (N_4701,N_4488,N_4434);
or U4702 (N_4702,N_4468,N_4576);
and U4703 (N_4703,N_4558,N_4408);
and U4704 (N_4704,N_4591,N_4557);
xor U4705 (N_4705,N_4543,N_4575);
or U4706 (N_4706,N_4591,N_4597);
and U4707 (N_4707,N_4434,N_4539);
nand U4708 (N_4708,N_4483,N_4453);
nand U4709 (N_4709,N_4557,N_4588);
and U4710 (N_4710,N_4480,N_4522);
or U4711 (N_4711,N_4587,N_4427);
nand U4712 (N_4712,N_4554,N_4592);
nor U4713 (N_4713,N_4542,N_4447);
nand U4714 (N_4714,N_4563,N_4575);
nor U4715 (N_4715,N_4531,N_4448);
or U4716 (N_4716,N_4493,N_4447);
nand U4717 (N_4717,N_4567,N_4457);
or U4718 (N_4718,N_4583,N_4419);
and U4719 (N_4719,N_4577,N_4437);
nor U4720 (N_4720,N_4435,N_4527);
nand U4721 (N_4721,N_4551,N_4510);
and U4722 (N_4722,N_4426,N_4469);
nor U4723 (N_4723,N_4486,N_4462);
nand U4724 (N_4724,N_4598,N_4402);
nand U4725 (N_4725,N_4416,N_4583);
nand U4726 (N_4726,N_4502,N_4451);
and U4727 (N_4727,N_4528,N_4551);
and U4728 (N_4728,N_4563,N_4488);
nor U4729 (N_4729,N_4461,N_4548);
nand U4730 (N_4730,N_4497,N_4495);
and U4731 (N_4731,N_4439,N_4463);
nor U4732 (N_4732,N_4501,N_4479);
nand U4733 (N_4733,N_4596,N_4487);
and U4734 (N_4734,N_4466,N_4469);
or U4735 (N_4735,N_4519,N_4502);
nand U4736 (N_4736,N_4583,N_4570);
nand U4737 (N_4737,N_4454,N_4472);
nand U4738 (N_4738,N_4461,N_4410);
nor U4739 (N_4739,N_4504,N_4492);
and U4740 (N_4740,N_4596,N_4506);
and U4741 (N_4741,N_4511,N_4582);
or U4742 (N_4742,N_4480,N_4504);
and U4743 (N_4743,N_4403,N_4474);
and U4744 (N_4744,N_4427,N_4539);
nor U4745 (N_4745,N_4501,N_4450);
or U4746 (N_4746,N_4452,N_4406);
nand U4747 (N_4747,N_4596,N_4453);
or U4748 (N_4748,N_4485,N_4428);
and U4749 (N_4749,N_4587,N_4591);
nor U4750 (N_4750,N_4570,N_4462);
and U4751 (N_4751,N_4414,N_4554);
and U4752 (N_4752,N_4486,N_4406);
and U4753 (N_4753,N_4414,N_4523);
and U4754 (N_4754,N_4432,N_4542);
nand U4755 (N_4755,N_4498,N_4538);
nand U4756 (N_4756,N_4484,N_4423);
nand U4757 (N_4757,N_4562,N_4480);
or U4758 (N_4758,N_4559,N_4474);
nand U4759 (N_4759,N_4464,N_4426);
or U4760 (N_4760,N_4510,N_4531);
nor U4761 (N_4761,N_4564,N_4408);
nand U4762 (N_4762,N_4447,N_4581);
and U4763 (N_4763,N_4539,N_4496);
nor U4764 (N_4764,N_4594,N_4547);
xnor U4765 (N_4765,N_4465,N_4551);
nor U4766 (N_4766,N_4408,N_4452);
and U4767 (N_4767,N_4436,N_4594);
nand U4768 (N_4768,N_4416,N_4419);
nor U4769 (N_4769,N_4490,N_4549);
nand U4770 (N_4770,N_4488,N_4485);
nand U4771 (N_4771,N_4423,N_4401);
or U4772 (N_4772,N_4500,N_4411);
or U4773 (N_4773,N_4521,N_4467);
and U4774 (N_4774,N_4464,N_4478);
nand U4775 (N_4775,N_4445,N_4440);
or U4776 (N_4776,N_4404,N_4498);
or U4777 (N_4777,N_4472,N_4567);
nand U4778 (N_4778,N_4504,N_4525);
xnor U4779 (N_4779,N_4514,N_4459);
nor U4780 (N_4780,N_4524,N_4474);
or U4781 (N_4781,N_4423,N_4549);
nor U4782 (N_4782,N_4567,N_4559);
nor U4783 (N_4783,N_4453,N_4415);
and U4784 (N_4784,N_4503,N_4593);
nand U4785 (N_4785,N_4438,N_4478);
nor U4786 (N_4786,N_4404,N_4501);
nand U4787 (N_4787,N_4514,N_4506);
and U4788 (N_4788,N_4418,N_4431);
nand U4789 (N_4789,N_4531,N_4532);
nand U4790 (N_4790,N_4436,N_4519);
or U4791 (N_4791,N_4525,N_4406);
and U4792 (N_4792,N_4568,N_4558);
or U4793 (N_4793,N_4502,N_4596);
nand U4794 (N_4794,N_4588,N_4427);
or U4795 (N_4795,N_4498,N_4495);
or U4796 (N_4796,N_4563,N_4516);
or U4797 (N_4797,N_4552,N_4452);
or U4798 (N_4798,N_4410,N_4586);
nor U4799 (N_4799,N_4465,N_4427);
nand U4800 (N_4800,N_4684,N_4687);
nor U4801 (N_4801,N_4726,N_4685);
or U4802 (N_4802,N_4609,N_4771);
xor U4803 (N_4803,N_4749,N_4743);
nor U4804 (N_4804,N_4733,N_4678);
nand U4805 (N_4805,N_4746,N_4706);
xor U4806 (N_4806,N_4671,N_4797);
nor U4807 (N_4807,N_4623,N_4646);
or U4808 (N_4808,N_4773,N_4638);
and U4809 (N_4809,N_4704,N_4738);
or U4810 (N_4810,N_4636,N_4673);
xor U4811 (N_4811,N_4770,N_4703);
nor U4812 (N_4812,N_4754,N_4748);
and U4813 (N_4813,N_4639,N_4651);
and U4814 (N_4814,N_4735,N_4731);
or U4815 (N_4815,N_4669,N_4697);
nor U4816 (N_4816,N_4653,N_4760);
or U4817 (N_4817,N_4634,N_4615);
and U4818 (N_4818,N_4790,N_4766);
or U4819 (N_4819,N_4739,N_4755);
or U4820 (N_4820,N_4781,N_4768);
nand U4821 (N_4821,N_4605,N_4788);
or U4822 (N_4822,N_4759,N_4649);
nand U4823 (N_4823,N_4747,N_4780);
nor U4824 (N_4824,N_4689,N_4719);
or U4825 (N_4825,N_4796,N_4789);
nand U4826 (N_4826,N_4660,N_4787);
nand U4827 (N_4827,N_4705,N_4715);
or U4828 (N_4828,N_4792,N_4799);
or U4829 (N_4829,N_4690,N_4745);
or U4830 (N_4830,N_4741,N_4722);
nand U4831 (N_4831,N_4647,N_4682);
or U4832 (N_4832,N_4778,N_4620);
nor U4833 (N_4833,N_4717,N_4603);
or U4834 (N_4834,N_4652,N_4712);
nor U4835 (N_4835,N_4751,N_4650);
nor U4836 (N_4836,N_4737,N_4718);
and U4837 (N_4837,N_4711,N_4798);
nand U4838 (N_4838,N_4645,N_4723);
nor U4839 (N_4839,N_4698,N_4602);
or U4840 (N_4840,N_4765,N_4606);
nor U4841 (N_4841,N_4707,N_4693);
xor U4842 (N_4842,N_4661,N_4728);
nand U4843 (N_4843,N_4643,N_4710);
and U4844 (N_4844,N_4648,N_4637);
or U4845 (N_4845,N_4656,N_4607);
and U4846 (N_4846,N_4720,N_4694);
and U4847 (N_4847,N_4785,N_4665);
or U4848 (N_4848,N_4696,N_4794);
or U4849 (N_4849,N_4667,N_4672);
and U4850 (N_4850,N_4692,N_4608);
nor U4851 (N_4851,N_4627,N_4763);
or U4852 (N_4852,N_4662,N_4752);
nor U4853 (N_4853,N_4611,N_4625);
nand U4854 (N_4854,N_4757,N_4612);
and U4855 (N_4855,N_4716,N_4688);
xnor U4856 (N_4856,N_4680,N_4644);
nand U4857 (N_4857,N_4736,N_4708);
and U4858 (N_4858,N_4633,N_4668);
nor U4859 (N_4859,N_4730,N_4774);
nand U4860 (N_4860,N_4775,N_4756);
nor U4861 (N_4861,N_4664,N_4626);
and U4862 (N_4862,N_4630,N_4721);
nand U4863 (N_4863,N_4655,N_4740);
nand U4864 (N_4864,N_4622,N_4617);
nand U4865 (N_4865,N_4679,N_4786);
and U4866 (N_4866,N_4695,N_4795);
nor U4867 (N_4867,N_4629,N_4610);
nand U4868 (N_4868,N_4742,N_4691);
or U4869 (N_4869,N_4714,N_4729);
or U4870 (N_4870,N_4621,N_4784);
nor U4871 (N_4871,N_4724,N_4744);
xnor U4872 (N_4872,N_4631,N_4663);
xor U4873 (N_4873,N_4761,N_4642);
xor U4874 (N_4874,N_4659,N_4614);
or U4875 (N_4875,N_4783,N_4750);
and U4876 (N_4876,N_4699,N_4793);
nor U4877 (N_4877,N_4686,N_4734);
nor U4878 (N_4878,N_4777,N_4628);
or U4879 (N_4879,N_4675,N_4624);
and U4880 (N_4880,N_4758,N_4658);
nor U4881 (N_4881,N_4613,N_4676);
and U4882 (N_4882,N_4701,N_4791);
and U4883 (N_4883,N_4635,N_4725);
nor U4884 (N_4884,N_4601,N_4674);
nand U4885 (N_4885,N_4713,N_4619);
xnor U4886 (N_4886,N_4641,N_4666);
or U4887 (N_4887,N_4670,N_4782);
nand U4888 (N_4888,N_4618,N_4769);
and U4889 (N_4889,N_4764,N_4753);
or U4890 (N_4890,N_4677,N_4657);
and U4891 (N_4891,N_4776,N_4762);
or U4892 (N_4892,N_4632,N_4767);
or U4893 (N_4893,N_4683,N_4654);
nand U4894 (N_4894,N_4732,N_4600);
xor U4895 (N_4895,N_4700,N_4727);
nand U4896 (N_4896,N_4709,N_4604);
nor U4897 (N_4897,N_4772,N_4616);
nand U4898 (N_4898,N_4640,N_4681);
nand U4899 (N_4899,N_4779,N_4702);
nand U4900 (N_4900,N_4707,N_4776);
or U4901 (N_4901,N_4692,N_4753);
nand U4902 (N_4902,N_4774,N_4605);
xor U4903 (N_4903,N_4737,N_4708);
and U4904 (N_4904,N_4743,N_4622);
and U4905 (N_4905,N_4620,N_4610);
nand U4906 (N_4906,N_4739,N_4757);
or U4907 (N_4907,N_4647,N_4792);
nand U4908 (N_4908,N_4626,N_4778);
or U4909 (N_4909,N_4765,N_4777);
nor U4910 (N_4910,N_4685,N_4784);
and U4911 (N_4911,N_4601,N_4787);
nand U4912 (N_4912,N_4717,N_4797);
and U4913 (N_4913,N_4602,N_4650);
xnor U4914 (N_4914,N_4653,N_4736);
nand U4915 (N_4915,N_4675,N_4704);
nor U4916 (N_4916,N_4603,N_4624);
nor U4917 (N_4917,N_4792,N_4727);
and U4918 (N_4918,N_4781,N_4791);
xor U4919 (N_4919,N_4755,N_4749);
nand U4920 (N_4920,N_4755,N_4673);
or U4921 (N_4921,N_4715,N_4778);
nor U4922 (N_4922,N_4610,N_4750);
and U4923 (N_4923,N_4794,N_4763);
nand U4924 (N_4924,N_4630,N_4725);
nand U4925 (N_4925,N_4670,N_4781);
and U4926 (N_4926,N_4791,N_4604);
nor U4927 (N_4927,N_4792,N_4644);
nor U4928 (N_4928,N_4742,N_4740);
nand U4929 (N_4929,N_4775,N_4768);
nand U4930 (N_4930,N_4612,N_4754);
or U4931 (N_4931,N_4648,N_4773);
nor U4932 (N_4932,N_4772,N_4643);
or U4933 (N_4933,N_4665,N_4754);
and U4934 (N_4934,N_4686,N_4755);
xor U4935 (N_4935,N_4788,N_4779);
nand U4936 (N_4936,N_4764,N_4629);
xnor U4937 (N_4937,N_4656,N_4686);
or U4938 (N_4938,N_4764,N_4744);
xnor U4939 (N_4939,N_4690,N_4766);
and U4940 (N_4940,N_4697,N_4671);
xor U4941 (N_4941,N_4600,N_4752);
nor U4942 (N_4942,N_4661,N_4679);
or U4943 (N_4943,N_4687,N_4732);
nor U4944 (N_4944,N_4778,N_4783);
and U4945 (N_4945,N_4617,N_4654);
xor U4946 (N_4946,N_4780,N_4785);
xnor U4947 (N_4947,N_4688,N_4694);
and U4948 (N_4948,N_4719,N_4644);
nand U4949 (N_4949,N_4754,N_4668);
xor U4950 (N_4950,N_4771,N_4799);
nor U4951 (N_4951,N_4689,N_4678);
and U4952 (N_4952,N_4747,N_4797);
nand U4953 (N_4953,N_4625,N_4674);
nand U4954 (N_4954,N_4713,N_4695);
nand U4955 (N_4955,N_4629,N_4754);
nor U4956 (N_4956,N_4620,N_4784);
or U4957 (N_4957,N_4717,N_4739);
and U4958 (N_4958,N_4739,N_4770);
nor U4959 (N_4959,N_4764,N_4715);
or U4960 (N_4960,N_4681,N_4728);
nor U4961 (N_4961,N_4785,N_4784);
xor U4962 (N_4962,N_4770,N_4783);
nor U4963 (N_4963,N_4623,N_4686);
or U4964 (N_4964,N_4764,N_4738);
or U4965 (N_4965,N_4697,N_4782);
nand U4966 (N_4966,N_4618,N_4652);
xnor U4967 (N_4967,N_4667,N_4650);
nor U4968 (N_4968,N_4664,N_4658);
nand U4969 (N_4969,N_4629,N_4795);
nand U4970 (N_4970,N_4606,N_4770);
and U4971 (N_4971,N_4664,N_4762);
and U4972 (N_4972,N_4617,N_4718);
nand U4973 (N_4973,N_4712,N_4698);
or U4974 (N_4974,N_4771,N_4662);
nor U4975 (N_4975,N_4641,N_4786);
and U4976 (N_4976,N_4770,N_4759);
xnor U4977 (N_4977,N_4697,N_4682);
nor U4978 (N_4978,N_4797,N_4658);
and U4979 (N_4979,N_4762,N_4623);
nor U4980 (N_4980,N_4789,N_4756);
nor U4981 (N_4981,N_4668,N_4650);
or U4982 (N_4982,N_4771,N_4781);
nand U4983 (N_4983,N_4649,N_4774);
nand U4984 (N_4984,N_4736,N_4738);
nor U4985 (N_4985,N_4675,N_4671);
or U4986 (N_4986,N_4645,N_4772);
nand U4987 (N_4987,N_4763,N_4758);
nand U4988 (N_4988,N_4716,N_4663);
and U4989 (N_4989,N_4768,N_4680);
nor U4990 (N_4990,N_4772,N_4681);
and U4991 (N_4991,N_4652,N_4776);
and U4992 (N_4992,N_4617,N_4669);
and U4993 (N_4993,N_4633,N_4725);
and U4994 (N_4994,N_4706,N_4781);
and U4995 (N_4995,N_4669,N_4645);
nand U4996 (N_4996,N_4628,N_4603);
or U4997 (N_4997,N_4773,N_4694);
or U4998 (N_4998,N_4673,N_4679);
nand U4999 (N_4999,N_4718,N_4658);
and UO_0 (O_0,N_4937,N_4883);
and UO_1 (O_1,N_4886,N_4849);
nand UO_2 (O_2,N_4943,N_4839);
and UO_3 (O_3,N_4820,N_4963);
and UO_4 (O_4,N_4955,N_4959);
or UO_5 (O_5,N_4928,N_4854);
xnor UO_6 (O_6,N_4816,N_4958);
nor UO_7 (O_7,N_4973,N_4826);
nand UO_8 (O_8,N_4867,N_4814);
nor UO_9 (O_9,N_4843,N_4862);
or UO_10 (O_10,N_4819,N_4805);
and UO_11 (O_11,N_4813,N_4914);
xnor UO_12 (O_12,N_4897,N_4803);
xor UO_13 (O_13,N_4917,N_4994);
nand UO_14 (O_14,N_4919,N_4988);
nand UO_15 (O_15,N_4865,N_4936);
nand UO_16 (O_16,N_4868,N_4837);
or UO_17 (O_17,N_4829,N_4907);
nand UO_18 (O_18,N_4881,N_4991);
and UO_19 (O_19,N_4824,N_4930);
nand UO_20 (O_20,N_4961,N_4836);
and UO_21 (O_21,N_4845,N_4817);
or UO_22 (O_22,N_4896,N_4864);
nand UO_23 (O_23,N_4890,N_4997);
nor UO_24 (O_24,N_4835,N_4978);
nand UO_25 (O_25,N_4894,N_4893);
or UO_26 (O_26,N_4982,N_4830);
nor UO_27 (O_27,N_4898,N_4832);
nand UO_28 (O_28,N_4987,N_4840);
nand UO_29 (O_29,N_4852,N_4825);
or UO_30 (O_30,N_4876,N_4884);
or UO_31 (O_31,N_4815,N_4934);
nor UO_32 (O_32,N_4915,N_4960);
nor UO_33 (O_33,N_4810,N_4941);
and UO_34 (O_34,N_4892,N_4861);
nand UO_35 (O_35,N_4956,N_4908);
and UO_36 (O_36,N_4850,N_4834);
nand UO_37 (O_37,N_4828,N_4831);
and UO_38 (O_38,N_4848,N_4906);
or UO_39 (O_39,N_4935,N_4980);
and UO_40 (O_40,N_4913,N_4900);
xor UO_41 (O_41,N_4986,N_4841);
and UO_42 (O_42,N_4860,N_4968);
nand UO_43 (O_43,N_4871,N_4899);
nor UO_44 (O_44,N_4844,N_4995);
or UO_45 (O_45,N_4911,N_4838);
nor UO_46 (O_46,N_4891,N_4903);
or UO_47 (O_47,N_4802,N_4901);
or UO_48 (O_48,N_4969,N_4947);
nor UO_49 (O_49,N_4990,N_4909);
nor UO_50 (O_50,N_4926,N_4873);
xor UO_51 (O_51,N_4921,N_4944);
xnor UO_52 (O_52,N_4869,N_4853);
and UO_53 (O_53,N_4974,N_4940);
nor UO_54 (O_54,N_4938,N_4927);
and UO_55 (O_55,N_4957,N_4954);
nor UO_56 (O_56,N_4970,N_4847);
and UO_57 (O_57,N_4823,N_4976);
and UO_58 (O_58,N_4812,N_4916);
nor UO_59 (O_59,N_4939,N_4851);
xor UO_60 (O_60,N_4855,N_4999);
or UO_61 (O_61,N_4967,N_4932);
or UO_62 (O_62,N_4842,N_4910);
and UO_63 (O_63,N_4889,N_4931);
or UO_64 (O_64,N_4822,N_4993);
and UO_65 (O_65,N_4858,N_4918);
nor UO_66 (O_66,N_4964,N_4981);
or UO_67 (O_67,N_4996,N_4952);
nand UO_68 (O_68,N_4818,N_4821);
nand UO_69 (O_69,N_4965,N_4902);
nor UO_70 (O_70,N_4863,N_4972);
or UO_71 (O_71,N_4827,N_4998);
nor UO_72 (O_72,N_4923,N_4946);
and UO_73 (O_73,N_4888,N_4962);
and UO_74 (O_74,N_4833,N_4880);
and UO_75 (O_75,N_4945,N_4875);
nand UO_76 (O_76,N_4887,N_4992);
and UO_77 (O_77,N_4800,N_4951);
nand UO_78 (O_78,N_4895,N_4971);
or UO_79 (O_79,N_4804,N_4977);
or UO_80 (O_80,N_4933,N_4929);
or UO_81 (O_81,N_4966,N_4882);
or UO_82 (O_82,N_4948,N_4950);
nor UO_83 (O_83,N_4885,N_4846);
or UO_84 (O_84,N_4984,N_4922);
nand UO_85 (O_85,N_4979,N_4801);
xnor UO_86 (O_86,N_4859,N_4989);
nand UO_87 (O_87,N_4878,N_4866);
nor UO_88 (O_88,N_4857,N_4949);
nand UO_89 (O_89,N_4874,N_4925);
nand UO_90 (O_90,N_4808,N_4953);
or UO_91 (O_91,N_4870,N_4879);
xor UO_92 (O_92,N_4807,N_4904);
or UO_93 (O_93,N_4920,N_4924);
and UO_94 (O_94,N_4811,N_4872);
nor UO_95 (O_95,N_4985,N_4877);
nand UO_96 (O_96,N_4806,N_4983);
nand UO_97 (O_97,N_4942,N_4809);
nand UO_98 (O_98,N_4856,N_4975);
xor UO_99 (O_99,N_4912,N_4905);
or UO_100 (O_100,N_4829,N_4850);
nand UO_101 (O_101,N_4872,N_4807);
or UO_102 (O_102,N_4834,N_4821);
and UO_103 (O_103,N_4964,N_4968);
nand UO_104 (O_104,N_4992,N_4866);
or UO_105 (O_105,N_4971,N_4960);
nand UO_106 (O_106,N_4891,N_4816);
and UO_107 (O_107,N_4942,N_4978);
nor UO_108 (O_108,N_4937,N_4979);
and UO_109 (O_109,N_4851,N_4865);
nor UO_110 (O_110,N_4890,N_4911);
and UO_111 (O_111,N_4852,N_4978);
xor UO_112 (O_112,N_4890,N_4917);
or UO_113 (O_113,N_4809,N_4832);
and UO_114 (O_114,N_4997,N_4999);
nor UO_115 (O_115,N_4947,N_4978);
and UO_116 (O_116,N_4845,N_4857);
nand UO_117 (O_117,N_4960,N_4959);
nor UO_118 (O_118,N_4906,N_4958);
or UO_119 (O_119,N_4988,N_4817);
or UO_120 (O_120,N_4952,N_4835);
nand UO_121 (O_121,N_4895,N_4869);
and UO_122 (O_122,N_4873,N_4903);
or UO_123 (O_123,N_4861,N_4994);
or UO_124 (O_124,N_4939,N_4961);
or UO_125 (O_125,N_4971,N_4996);
nor UO_126 (O_126,N_4973,N_4832);
nand UO_127 (O_127,N_4844,N_4959);
and UO_128 (O_128,N_4967,N_4976);
or UO_129 (O_129,N_4813,N_4905);
and UO_130 (O_130,N_4939,N_4805);
and UO_131 (O_131,N_4816,N_4920);
nand UO_132 (O_132,N_4926,N_4943);
or UO_133 (O_133,N_4997,N_4936);
nand UO_134 (O_134,N_4953,N_4820);
nand UO_135 (O_135,N_4930,N_4951);
or UO_136 (O_136,N_4904,N_4890);
nand UO_137 (O_137,N_4868,N_4977);
nor UO_138 (O_138,N_4898,N_4810);
nand UO_139 (O_139,N_4814,N_4907);
nor UO_140 (O_140,N_4881,N_4822);
nand UO_141 (O_141,N_4900,N_4808);
nor UO_142 (O_142,N_4825,N_4960);
nor UO_143 (O_143,N_4873,N_4846);
or UO_144 (O_144,N_4906,N_4930);
or UO_145 (O_145,N_4879,N_4846);
and UO_146 (O_146,N_4964,N_4840);
nand UO_147 (O_147,N_4982,N_4889);
and UO_148 (O_148,N_4850,N_4904);
xnor UO_149 (O_149,N_4843,N_4901);
nand UO_150 (O_150,N_4934,N_4886);
nand UO_151 (O_151,N_4972,N_4916);
xor UO_152 (O_152,N_4860,N_4832);
xnor UO_153 (O_153,N_4833,N_4903);
and UO_154 (O_154,N_4818,N_4910);
and UO_155 (O_155,N_4838,N_4933);
nand UO_156 (O_156,N_4870,N_4891);
nand UO_157 (O_157,N_4835,N_4956);
nand UO_158 (O_158,N_4864,N_4868);
and UO_159 (O_159,N_4863,N_4988);
nor UO_160 (O_160,N_4925,N_4918);
xor UO_161 (O_161,N_4871,N_4930);
xnor UO_162 (O_162,N_4997,N_4896);
xnor UO_163 (O_163,N_4831,N_4909);
nand UO_164 (O_164,N_4803,N_4814);
nand UO_165 (O_165,N_4936,N_4885);
or UO_166 (O_166,N_4971,N_4867);
or UO_167 (O_167,N_4814,N_4948);
nand UO_168 (O_168,N_4842,N_4801);
and UO_169 (O_169,N_4941,N_4813);
xor UO_170 (O_170,N_4854,N_4806);
or UO_171 (O_171,N_4982,N_4901);
or UO_172 (O_172,N_4974,N_4886);
or UO_173 (O_173,N_4980,N_4967);
or UO_174 (O_174,N_4940,N_4857);
xor UO_175 (O_175,N_4973,N_4933);
nand UO_176 (O_176,N_4872,N_4959);
nand UO_177 (O_177,N_4996,N_4800);
nand UO_178 (O_178,N_4809,N_4826);
nand UO_179 (O_179,N_4979,N_4902);
nand UO_180 (O_180,N_4803,N_4935);
nor UO_181 (O_181,N_4947,N_4856);
nand UO_182 (O_182,N_4828,N_4986);
nor UO_183 (O_183,N_4985,N_4954);
xnor UO_184 (O_184,N_4887,N_4934);
nor UO_185 (O_185,N_4934,N_4875);
nand UO_186 (O_186,N_4848,N_4897);
or UO_187 (O_187,N_4985,N_4901);
nand UO_188 (O_188,N_4856,N_4960);
nand UO_189 (O_189,N_4850,N_4935);
nor UO_190 (O_190,N_4993,N_4878);
nand UO_191 (O_191,N_4934,N_4944);
nand UO_192 (O_192,N_4921,N_4804);
and UO_193 (O_193,N_4891,N_4832);
or UO_194 (O_194,N_4932,N_4863);
nor UO_195 (O_195,N_4880,N_4950);
or UO_196 (O_196,N_4860,N_4826);
and UO_197 (O_197,N_4811,N_4963);
and UO_198 (O_198,N_4858,N_4950);
or UO_199 (O_199,N_4989,N_4992);
xor UO_200 (O_200,N_4900,N_4873);
xor UO_201 (O_201,N_4958,N_4883);
and UO_202 (O_202,N_4890,N_4928);
nor UO_203 (O_203,N_4960,N_4854);
or UO_204 (O_204,N_4979,N_4863);
and UO_205 (O_205,N_4972,N_4872);
nand UO_206 (O_206,N_4876,N_4885);
nor UO_207 (O_207,N_4891,N_4960);
nand UO_208 (O_208,N_4813,N_4879);
xor UO_209 (O_209,N_4827,N_4988);
and UO_210 (O_210,N_4966,N_4899);
nor UO_211 (O_211,N_4953,N_4836);
and UO_212 (O_212,N_4814,N_4801);
or UO_213 (O_213,N_4937,N_4893);
nand UO_214 (O_214,N_4909,N_4951);
or UO_215 (O_215,N_4808,N_4846);
nand UO_216 (O_216,N_4979,N_4875);
or UO_217 (O_217,N_4873,N_4806);
nor UO_218 (O_218,N_4861,N_4925);
nand UO_219 (O_219,N_4966,N_4839);
nand UO_220 (O_220,N_4804,N_4848);
nand UO_221 (O_221,N_4920,N_4994);
nand UO_222 (O_222,N_4913,N_4857);
or UO_223 (O_223,N_4803,N_4860);
nand UO_224 (O_224,N_4845,N_4979);
or UO_225 (O_225,N_4800,N_4845);
or UO_226 (O_226,N_4897,N_4869);
or UO_227 (O_227,N_4915,N_4905);
nand UO_228 (O_228,N_4999,N_4875);
nor UO_229 (O_229,N_4816,N_4979);
or UO_230 (O_230,N_4859,N_4925);
and UO_231 (O_231,N_4989,N_4811);
or UO_232 (O_232,N_4885,N_4891);
and UO_233 (O_233,N_4828,N_4981);
and UO_234 (O_234,N_4831,N_4904);
and UO_235 (O_235,N_4992,N_4991);
or UO_236 (O_236,N_4895,N_4948);
xor UO_237 (O_237,N_4843,N_4915);
and UO_238 (O_238,N_4912,N_4985);
or UO_239 (O_239,N_4961,N_4986);
or UO_240 (O_240,N_4907,N_4944);
nor UO_241 (O_241,N_4908,N_4826);
or UO_242 (O_242,N_4989,N_4922);
and UO_243 (O_243,N_4974,N_4807);
or UO_244 (O_244,N_4940,N_4812);
or UO_245 (O_245,N_4923,N_4956);
or UO_246 (O_246,N_4951,N_4979);
xnor UO_247 (O_247,N_4951,N_4995);
nand UO_248 (O_248,N_4813,N_4955);
or UO_249 (O_249,N_4857,N_4887);
nand UO_250 (O_250,N_4905,N_4998);
or UO_251 (O_251,N_4949,N_4892);
nand UO_252 (O_252,N_4854,N_4995);
and UO_253 (O_253,N_4980,N_4837);
or UO_254 (O_254,N_4812,N_4887);
or UO_255 (O_255,N_4879,N_4853);
or UO_256 (O_256,N_4848,N_4968);
or UO_257 (O_257,N_4809,N_4804);
nor UO_258 (O_258,N_4815,N_4846);
xnor UO_259 (O_259,N_4980,N_4819);
and UO_260 (O_260,N_4971,N_4952);
nand UO_261 (O_261,N_4837,N_4865);
nor UO_262 (O_262,N_4846,N_4868);
nand UO_263 (O_263,N_4839,N_4823);
nor UO_264 (O_264,N_4925,N_4990);
nor UO_265 (O_265,N_4903,N_4976);
nor UO_266 (O_266,N_4815,N_4919);
nor UO_267 (O_267,N_4974,N_4818);
and UO_268 (O_268,N_4822,N_4809);
nand UO_269 (O_269,N_4813,N_4802);
or UO_270 (O_270,N_4889,N_4938);
or UO_271 (O_271,N_4938,N_4906);
or UO_272 (O_272,N_4843,N_4952);
and UO_273 (O_273,N_4847,N_4916);
nor UO_274 (O_274,N_4890,N_4990);
nand UO_275 (O_275,N_4931,N_4972);
or UO_276 (O_276,N_4954,N_4916);
and UO_277 (O_277,N_4856,N_4986);
nor UO_278 (O_278,N_4956,N_4902);
and UO_279 (O_279,N_4935,N_4921);
and UO_280 (O_280,N_4930,N_4912);
nand UO_281 (O_281,N_4948,N_4981);
and UO_282 (O_282,N_4983,N_4870);
nor UO_283 (O_283,N_4945,N_4873);
and UO_284 (O_284,N_4977,N_4875);
or UO_285 (O_285,N_4828,N_4940);
nand UO_286 (O_286,N_4893,N_4960);
xnor UO_287 (O_287,N_4818,N_4846);
xnor UO_288 (O_288,N_4948,N_4890);
nand UO_289 (O_289,N_4916,N_4803);
xor UO_290 (O_290,N_4938,N_4987);
nor UO_291 (O_291,N_4926,N_4944);
nor UO_292 (O_292,N_4841,N_4976);
or UO_293 (O_293,N_4967,N_4987);
or UO_294 (O_294,N_4880,N_4809);
and UO_295 (O_295,N_4962,N_4802);
nand UO_296 (O_296,N_4976,N_4845);
nor UO_297 (O_297,N_4985,N_4979);
and UO_298 (O_298,N_4951,N_4906);
or UO_299 (O_299,N_4806,N_4835);
nor UO_300 (O_300,N_4940,N_4849);
or UO_301 (O_301,N_4965,N_4858);
nor UO_302 (O_302,N_4976,N_4872);
nor UO_303 (O_303,N_4888,N_4929);
nor UO_304 (O_304,N_4974,N_4993);
xnor UO_305 (O_305,N_4873,N_4841);
xor UO_306 (O_306,N_4906,N_4814);
nor UO_307 (O_307,N_4836,N_4891);
nand UO_308 (O_308,N_4877,N_4853);
or UO_309 (O_309,N_4845,N_4809);
or UO_310 (O_310,N_4975,N_4878);
nand UO_311 (O_311,N_4850,N_4818);
nand UO_312 (O_312,N_4981,N_4935);
or UO_313 (O_313,N_4893,N_4987);
and UO_314 (O_314,N_4824,N_4819);
nor UO_315 (O_315,N_4856,N_4911);
nor UO_316 (O_316,N_4993,N_4871);
and UO_317 (O_317,N_4837,N_4895);
nand UO_318 (O_318,N_4968,N_4950);
nand UO_319 (O_319,N_4959,N_4866);
and UO_320 (O_320,N_4897,N_4823);
xor UO_321 (O_321,N_4951,N_4908);
nor UO_322 (O_322,N_4836,N_4998);
xnor UO_323 (O_323,N_4929,N_4871);
nor UO_324 (O_324,N_4984,N_4901);
or UO_325 (O_325,N_4836,N_4937);
or UO_326 (O_326,N_4994,N_4992);
and UO_327 (O_327,N_4901,N_4916);
nand UO_328 (O_328,N_4967,N_4950);
nand UO_329 (O_329,N_4950,N_4925);
and UO_330 (O_330,N_4880,N_4832);
or UO_331 (O_331,N_4821,N_4838);
and UO_332 (O_332,N_4862,N_4810);
nor UO_333 (O_333,N_4923,N_4895);
nand UO_334 (O_334,N_4838,N_4982);
xor UO_335 (O_335,N_4841,N_4974);
nand UO_336 (O_336,N_4936,N_4948);
and UO_337 (O_337,N_4899,N_4819);
or UO_338 (O_338,N_4857,N_4876);
and UO_339 (O_339,N_4839,N_4846);
xor UO_340 (O_340,N_4820,N_4983);
nand UO_341 (O_341,N_4936,N_4903);
or UO_342 (O_342,N_4923,N_4861);
xnor UO_343 (O_343,N_4810,N_4992);
nor UO_344 (O_344,N_4879,N_4823);
and UO_345 (O_345,N_4960,N_4812);
or UO_346 (O_346,N_4885,N_4941);
nor UO_347 (O_347,N_4934,N_4903);
xnor UO_348 (O_348,N_4983,N_4884);
or UO_349 (O_349,N_4913,N_4823);
or UO_350 (O_350,N_4811,N_4842);
or UO_351 (O_351,N_4822,N_4843);
xor UO_352 (O_352,N_4807,N_4962);
xnor UO_353 (O_353,N_4858,N_4966);
or UO_354 (O_354,N_4888,N_4954);
and UO_355 (O_355,N_4920,N_4859);
xor UO_356 (O_356,N_4817,N_4927);
nand UO_357 (O_357,N_4899,N_4974);
nand UO_358 (O_358,N_4999,N_4949);
nor UO_359 (O_359,N_4938,N_4994);
and UO_360 (O_360,N_4839,N_4932);
nor UO_361 (O_361,N_4838,N_4802);
and UO_362 (O_362,N_4838,N_4985);
and UO_363 (O_363,N_4885,N_4985);
and UO_364 (O_364,N_4895,N_4831);
nand UO_365 (O_365,N_4981,N_4908);
and UO_366 (O_366,N_4916,N_4825);
nor UO_367 (O_367,N_4916,N_4969);
nand UO_368 (O_368,N_4872,N_4836);
nand UO_369 (O_369,N_4963,N_4841);
and UO_370 (O_370,N_4882,N_4845);
nand UO_371 (O_371,N_4917,N_4871);
nand UO_372 (O_372,N_4873,N_4891);
nor UO_373 (O_373,N_4873,N_4961);
xnor UO_374 (O_374,N_4953,N_4982);
nor UO_375 (O_375,N_4992,N_4891);
nand UO_376 (O_376,N_4923,N_4818);
nand UO_377 (O_377,N_4824,N_4920);
or UO_378 (O_378,N_4986,N_4901);
or UO_379 (O_379,N_4863,N_4913);
and UO_380 (O_380,N_4940,N_4844);
nand UO_381 (O_381,N_4853,N_4999);
or UO_382 (O_382,N_4801,N_4873);
and UO_383 (O_383,N_4944,N_4918);
and UO_384 (O_384,N_4926,N_4912);
and UO_385 (O_385,N_4809,N_4829);
nand UO_386 (O_386,N_4878,N_4885);
xnor UO_387 (O_387,N_4817,N_4915);
xor UO_388 (O_388,N_4976,N_4906);
or UO_389 (O_389,N_4911,N_4827);
xor UO_390 (O_390,N_4847,N_4893);
nand UO_391 (O_391,N_4815,N_4907);
and UO_392 (O_392,N_4886,N_4912);
or UO_393 (O_393,N_4888,N_4987);
or UO_394 (O_394,N_4834,N_4911);
or UO_395 (O_395,N_4869,N_4832);
nor UO_396 (O_396,N_4828,N_4894);
nor UO_397 (O_397,N_4976,N_4826);
nor UO_398 (O_398,N_4943,N_4921);
nand UO_399 (O_399,N_4969,N_4920);
nand UO_400 (O_400,N_4895,N_4935);
nor UO_401 (O_401,N_4807,N_4997);
nor UO_402 (O_402,N_4855,N_4993);
nand UO_403 (O_403,N_4994,N_4928);
xor UO_404 (O_404,N_4902,N_4898);
nand UO_405 (O_405,N_4827,N_4885);
nand UO_406 (O_406,N_4843,N_4821);
or UO_407 (O_407,N_4845,N_4973);
nand UO_408 (O_408,N_4847,N_4815);
or UO_409 (O_409,N_4875,N_4840);
and UO_410 (O_410,N_4842,N_4802);
nand UO_411 (O_411,N_4838,N_4803);
and UO_412 (O_412,N_4872,N_4856);
xor UO_413 (O_413,N_4904,N_4953);
or UO_414 (O_414,N_4813,N_4931);
and UO_415 (O_415,N_4828,N_4857);
nand UO_416 (O_416,N_4854,N_4857);
or UO_417 (O_417,N_4941,N_4884);
or UO_418 (O_418,N_4816,N_4824);
nand UO_419 (O_419,N_4837,N_4952);
or UO_420 (O_420,N_4877,N_4929);
or UO_421 (O_421,N_4995,N_4984);
nand UO_422 (O_422,N_4825,N_4971);
and UO_423 (O_423,N_4833,N_4993);
nor UO_424 (O_424,N_4903,N_4827);
nor UO_425 (O_425,N_4969,N_4911);
nor UO_426 (O_426,N_4938,N_4807);
nor UO_427 (O_427,N_4983,N_4833);
and UO_428 (O_428,N_4813,N_4814);
nand UO_429 (O_429,N_4937,N_4948);
and UO_430 (O_430,N_4816,N_4840);
and UO_431 (O_431,N_4912,N_4808);
or UO_432 (O_432,N_4938,N_4806);
nor UO_433 (O_433,N_4994,N_4918);
or UO_434 (O_434,N_4951,N_4961);
or UO_435 (O_435,N_4951,N_4859);
and UO_436 (O_436,N_4924,N_4838);
nor UO_437 (O_437,N_4810,N_4848);
nor UO_438 (O_438,N_4984,N_4953);
and UO_439 (O_439,N_4815,N_4971);
xor UO_440 (O_440,N_4873,N_4929);
nand UO_441 (O_441,N_4895,N_4822);
nor UO_442 (O_442,N_4822,N_4896);
nand UO_443 (O_443,N_4986,N_4992);
and UO_444 (O_444,N_4929,N_4886);
xnor UO_445 (O_445,N_4914,N_4803);
nor UO_446 (O_446,N_4850,N_4800);
nor UO_447 (O_447,N_4908,N_4857);
nor UO_448 (O_448,N_4877,N_4816);
xor UO_449 (O_449,N_4852,N_4903);
or UO_450 (O_450,N_4904,N_4800);
and UO_451 (O_451,N_4837,N_4964);
nand UO_452 (O_452,N_4962,N_4960);
and UO_453 (O_453,N_4907,N_4986);
and UO_454 (O_454,N_4852,N_4921);
and UO_455 (O_455,N_4968,N_4919);
nor UO_456 (O_456,N_4836,N_4874);
or UO_457 (O_457,N_4954,N_4822);
and UO_458 (O_458,N_4925,N_4977);
nor UO_459 (O_459,N_4820,N_4821);
nand UO_460 (O_460,N_4880,N_4873);
nand UO_461 (O_461,N_4870,N_4985);
and UO_462 (O_462,N_4839,N_4879);
nor UO_463 (O_463,N_4851,N_4981);
nand UO_464 (O_464,N_4994,N_4860);
and UO_465 (O_465,N_4973,N_4996);
and UO_466 (O_466,N_4847,N_4858);
nand UO_467 (O_467,N_4847,N_4826);
nor UO_468 (O_468,N_4864,N_4821);
and UO_469 (O_469,N_4835,N_4977);
xnor UO_470 (O_470,N_4906,N_4819);
or UO_471 (O_471,N_4849,N_4867);
or UO_472 (O_472,N_4882,N_4993);
nor UO_473 (O_473,N_4959,N_4890);
and UO_474 (O_474,N_4971,N_4941);
nor UO_475 (O_475,N_4805,N_4904);
nor UO_476 (O_476,N_4801,N_4892);
nor UO_477 (O_477,N_4933,N_4980);
nand UO_478 (O_478,N_4947,N_4844);
nor UO_479 (O_479,N_4881,N_4895);
and UO_480 (O_480,N_4834,N_4895);
nor UO_481 (O_481,N_4974,N_4871);
and UO_482 (O_482,N_4947,N_4906);
nor UO_483 (O_483,N_4864,N_4838);
nor UO_484 (O_484,N_4894,N_4838);
or UO_485 (O_485,N_4921,N_4862);
or UO_486 (O_486,N_4956,N_4850);
nand UO_487 (O_487,N_4803,N_4863);
or UO_488 (O_488,N_4822,N_4933);
nand UO_489 (O_489,N_4889,N_4848);
and UO_490 (O_490,N_4857,N_4912);
and UO_491 (O_491,N_4940,N_4984);
nand UO_492 (O_492,N_4911,N_4909);
and UO_493 (O_493,N_4832,N_4909);
nor UO_494 (O_494,N_4861,N_4845);
xor UO_495 (O_495,N_4870,N_4945);
nor UO_496 (O_496,N_4998,N_4812);
nand UO_497 (O_497,N_4852,N_4948);
or UO_498 (O_498,N_4948,N_4953);
xnor UO_499 (O_499,N_4962,N_4939);
nor UO_500 (O_500,N_4958,N_4987);
nor UO_501 (O_501,N_4914,N_4825);
nor UO_502 (O_502,N_4854,N_4977);
or UO_503 (O_503,N_4939,N_4890);
or UO_504 (O_504,N_4942,N_4955);
or UO_505 (O_505,N_4813,N_4857);
nor UO_506 (O_506,N_4986,N_4940);
or UO_507 (O_507,N_4854,N_4931);
and UO_508 (O_508,N_4946,N_4948);
xor UO_509 (O_509,N_4970,N_4892);
and UO_510 (O_510,N_4868,N_4870);
and UO_511 (O_511,N_4996,N_4899);
nand UO_512 (O_512,N_4835,N_4850);
or UO_513 (O_513,N_4839,N_4909);
nor UO_514 (O_514,N_4908,N_4823);
and UO_515 (O_515,N_4943,N_4918);
nand UO_516 (O_516,N_4841,N_4985);
or UO_517 (O_517,N_4867,N_4848);
nand UO_518 (O_518,N_4988,N_4823);
and UO_519 (O_519,N_4812,N_4835);
nor UO_520 (O_520,N_4992,N_4840);
or UO_521 (O_521,N_4809,N_4860);
nor UO_522 (O_522,N_4877,N_4978);
or UO_523 (O_523,N_4942,N_4895);
nand UO_524 (O_524,N_4927,N_4963);
xor UO_525 (O_525,N_4955,N_4838);
xnor UO_526 (O_526,N_4883,N_4851);
nand UO_527 (O_527,N_4812,N_4833);
or UO_528 (O_528,N_4862,N_4889);
and UO_529 (O_529,N_4959,N_4829);
nor UO_530 (O_530,N_4883,N_4918);
nor UO_531 (O_531,N_4973,N_4846);
and UO_532 (O_532,N_4933,N_4808);
and UO_533 (O_533,N_4804,N_4938);
nor UO_534 (O_534,N_4934,N_4938);
and UO_535 (O_535,N_4895,N_4952);
nand UO_536 (O_536,N_4842,N_4876);
or UO_537 (O_537,N_4824,N_4845);
nand UO_538 (O_538,N_4850,N_4937);
and UO_539 (O_539,N_4983,N_4914);
and UO_540 (O_540,N_4990,N_4864);
nor UO_541 (O_541,N_4930,N_4933);
nand UO_542 (O_542,N_4804,N_4811);
or UO_543 (O_543,N_4984,N_4868);
or UO_544 (O_544,N_4997,N_4987);
or UO_545 (O_545,N_4983,N_4839);
xnor UO_546 (O_546,N_4894,N_4854);
nand UO_547 (O_547,N_4991,N_4960);
nand UO_548 (O_548,N_4810,N_4958);
or UO_549 (O_549,N_4990,N_4845);
nand UO_550 (O_550,N_4997,N_4924);
nand UO_551 (O_551,N_4831,N_4811);
xor UO_552 (O_552,N_4951,N_4851);
xnor UO_553 (O_553,N_4816,N_4861);
or UO_554 (O_554,N_4881,N_4925);
and UO_555 (O_555,N_4876,N_4921);
or UO_556 (O_556,N_4946,N_4996);
and UO_557 (O_557,N_4986,N_4932);
and UO_558 (O_558,N_4902,N_4976);
and UO_559 (O_559,N_4983,N_4952);
nand UO_560 (O_560,N_4995,N_4910);
nor UO_561 (O_561,N_4878,N_4914);
nor UO_562 (O_562,N_4979,N_4859);
nor UO_563 (O_563,N_4872,N_4964);
nand UO_564 (O_564,N_4884,N_4808);
and UO_565 (O_565,N_4972,N_4816);
nor UO_566 (O_566,N_4987,N_4899);
and UO_567 (O_567,N_4821,N_4970);
xnor UO_568 (O_568,N_4984,N_4895);
nand UO_569 (O_569,N_4994,N_4945);
xor UO_570 (O_570,N_4918,N_4989);
or UO_571 (O_571,N_4888,N_4975);
and UO_572 (O_572,N_4942,N_4967);
or UO_573 (O_573,N_4985,N_4821);
nand UO_574 (O_574,N_4978,N_4963);
xnor UO_575 (O_575,N_4931,N_4857);
or UO_576 (O_576,N_4971,N_4841);
and UO_577 (O_577,N_4866,N_4875);
nor UO_578 (O_578,N_4924,N_4821);
xnor UO_579 (O_579,N_4808,N_4968);
nor UO_580 (O_580,N_4984,N_4931);
nand UO_581 (O_581,N_4896,N_4853);
and UO_582 (O_582,N_4801,N_4935);
or UO_583 (O_583,N_4865,N_4947);
xnor UO_584 (O_584,N_4904,N_4971);
or UO_585 (O_585,N_4928,N_4807);
or UO_586 (O_586,N_4854,N_4913);
or UO_587 (O_587,N_4966,N_4832);
nor UO_588 (O_588,N_4988,N_4894);
nor UO_589 (O_589,N_4977,N_4929);
or UO_590 (O_590,N_4826,N_4959);
nor UO_591 (O_591,N_4975,N_4934);
nor UO_592 (O_592,N_4805,N_4806);
and UO_593 (O_593,N_4908,N_4852);
or UO_594 (O_594,N_4854,N_4838);
nand UO_595 (O_595,N_4938,N_4830);
nor UO_596 (O_596,N_4986,N_4922);
nor UO_597 (O_597,N_4893,N_4826);
nand UO_598 (O_598,N_4934,N_4939);
xnor UO_599 (O_599,N_4975,N_4858);
and UO_600 (O_600,N_4949,N_4910);
nand UO_601 (O_601,N_4917,N_4918);
and UO_602 (O_602,N_4840,N_4869);
or UO_603 (O_603,N_4822,N_4989);
nor UO_604 (O_604,N_4986,N_4991);
and UO_605 (O_605,N_4971,N_4958);
nand UO_606 (O_606,N_4917,N_4862);
and UO_607 (O_607,N_4886,N_4970);
nand UO_608 (O_608,N_4800,N_4843);
or UO_609 (O_609,N_4960,N_4920);
and UO_610 (O_610,N_4895,N_4824);
xnor UO_611 (O_611,N_4960,N_4918);
or UO_612 (O_612,N_4802,N_4984);
or UO_613 (O_613,N_4821,N_4993);
or UO_614 (O_614,N_4979,N_4898);
nor UO_615 (O_615,N_4878,N_4933);
or UO_616 (O_616,N_4886,N_4910);
nand UO_617 (O_617,N_4912,N_4866);
or UO_618 (O_618,N_4866,N_4867);
nand UO_619 (O_619,N_4928,N_4880);
nor UO_620 (O_620,N_4982,N_4948);
and UO_621 (O_621,N_4865,N_4970);
nand UO_622 (O_622,N_4963,N_4985);
xor UO_623 (O_623,N_4858,N_4921);
nand UO_624 (O_624,N_4816,N_4976);
nand UO_625 (O_625,N_4976,N_4969);
nor UO_626 (O_626,N_4858,N_4803);
nor UO_627 (O_627,N_4831,N_4880);
and UO_628 (O_628,N_4988,N_4929);
nor UO_629 (O_629,N_4929,N_4906);
nand UO_630 (O_630,N_4887,N_4837);
and UO_631 (O_631,N_4870,N_4850);
or UO_632 (O_632,N_4962,N_4857);
and UO_633 (O_633,N_4942,N_4987);
or UO_634 (O_634,N_4895,N_4943);
nand UO_635 (O_635,N_4882,N_4940);
nor UO_636 (O_636,N_4863,N_4964);
nand UO_637 (O_637,N_4827,N_4826);
or UO_638 (O_638,N_4923,N_4968);
or UO_639 (O_639,N_4994,N_4834);
nand UO_640 (O_640,N_4861,N_4912);
or UO_641 (O_641,N_4840,N_4893);
nor UO_642 (O_642,N_4880,N_4823);
and UO_643 (O_643,N_4982,N_4907);
xnor UO_644 (O_644,N_4812,N_4963);
and UO_645 (O_645,N_4878,N_4893);
nor UO_646 (O_646,N_4847,N_4886);
nor UO_647 (O_647,N_4836,N_4809);
or UO_648 (O_648,N_4958,N_4823);
or UO_649 (O_649,N_4913,N_4931);
or UO_650 (O_650,N_4991,N_4847);
nand UO_651 (O_651,N_4931,N_4906);
nand UO_652 (O_652,N_4823,N_4974);
nand UO_653 (O_653,N_4990,N_4984);
nand UO_654 (O_654,N_4941,N_4867);
nand UO_655 (O_655,N_4845,N_4904);
nand UO_656 (O_656,N_4852,N_4935);
nand UO_657 (O_657,N_4841,N_4936);
nand UO_658 (O_658,N_4951,N_4986);
nand UO_659 (O_659,N_4835,N_4992);
nor UO_660 (O_660,N_4893,N_4839);
or UO_661 (O_661,N_4974,N_4824);
and UO_662 (O_662,N_4898,N_4994);
and UO_663 (O_663,N_4983,N_4867);
xor UO_664 (O_664,N_4856,N_4870);
or UO_665 (O_665,N_4878,N_4855);
nand UO_666 (O_666,N_4828,N_4971);
nor UO_667 (O_667,N_4889,N_4970);
and UO_668 (O_668,N_4948,N_4934);
and UO_669 (O_669,N_4919,N_4848);
nand UO_670 (O_670,N_4886,N_4807);
nand UO_671 (O_671,N_4994,N_4961);
and UO_672 (O_672,N_4888,N_4953);
or UO_673 (O_673,N_4906,N_4884);
and UO_674 (O_674,N_4930,N_4929);
and UO_675 (O_675,N_4988,N_4862);
xnor UO_676 (O_676,N_4801,N_4871);
and UO_677 (O_677,N_4815,N_4962);
nor UO_678 (O_678,N_4954,N_4932);
and UO_679 (O_679,N_4904,N_4942);
and UO_680 (O_680,N_4922,N_4952);
or UO_681 (O_681,N_4864,N_4938);
or UO_682 (O_682,N_4866,N_4851);
nand UO_683 (O_683,N_4921,N_4805);
nand UO_684 (O_684,N_4803,N_4800);
or UO_685 (O_685,N_4861,N_4971);
nand UO_686 (O_686,N_4836,N_4972);
or UO_687 (O_687,N_4985,N_4941);
and UO_688 (O_688,N_4832,N_4933);
or UO_689 (O_689,N_4994,N_4950);
or UO_690 (O_690,N_4991,N_4851);
nor UO_691 (O_691,N_4811,N_4886);
nor UO_692 (O_692,N_4937,N_4831);
nand UO_693 (O_693,N_4924,N_4958);
nor UO_694 (O_694,N_4828,N_4923);
and UO_695 (O_695,N_4848,N_4869);
nor UO_696 (O_696,N_4800,N_4896);
xnor UO_697 (O_697,N_4804,N_4933);
or UO_698 (O_698,N_4848,N_4862);
nor UO_699 (O_699,N_4913,N_4969);
and UO_700 (O_700,N_4995,N_4903);
nor UO_701 (O_701,N_4859,N_4863);
nor UO_702 (O_702,N_4918,N_4971);
and UO_703 (O_703,N_4864,N_4870);
xnor UO_704 (O_704,N_4847,N_4902);
and UO_705 (O_705,N_4880,N_4917);
and UO_706 (O_706,N_4940,N_4806);
nor UO_707 (O_707,N_4944,N_4873);
and UO_708 (O_708,N_4903,N_4928);
nor UO_709 (O_709,N_4994,N_4971);
and UO_710 (O_710,N_4951,N_4914);
nor UO_711 (O_711,N_4952,N_4871);
nand UO_712 (O_712,N_4921,N_4934);
or UO_713 (O_713,N_4890,N_4992);
nand UO_714 (O_714,N_4941,N_4998);
nor UO_715 (O_715,N_4888,N_4980);
or UO_716 (O_716,N_4807,N_4987);
xnor UO_717 (O_717,N_4923,N_4856);
nand UO_718 (O_718,N_4966,N_4954);
and UO_719 (O_719,N_4907,N_4935);
and UO_720 (O_720,N_4865,N_4803);
nor UO_721 (O_721,N_4824,N_4809);
nand UO_722 (O_722,N_4941,N_4833);
nor UO_723 (O_723,N_4888,N_4834);
nor UO_724 (O_724,N_4819,N_4907);
xnor UO_725 (O_725,N_4835,N_4999);
xor UO_726 (O_726,N_4819,N_4826);
xor UO_727 (O_727,N_4888,N_4880);
and UO_728 (O_728,N_4923,N_4853);
or UO_729 (O_729,N_4884,N_4852);
or UO_730 (O_730,N_4890,N_4953);
nand UO_731 (O_731,N_4961,N_4912);
nand UO_732 (O_732,N_4894,N_4866);
or UO_733 (O_733,N_4926,N_4820);
nor UO_734 (O_734,N_4839,N_4990);
nor UO_735 (O_735,N_4913,N_4902);
nor UO_736 (O_736,N_4945,N_4913);
and UO_737 (O_737,N_4917,N_4970);
and UO_738 (O_738,N_4938,N_4854);
xor UO_739 (O_739,N_4804,N_4889);
and UO_740 (O_740,N_4879,N_4948);
nor UO_741 (O_741,N_4954,N_4912);
nand UO_742 (O_742,N_4969,N_4902);
nor UO_743 (O_743,N_4957,N_4898);
nor UO_744 (O_744,N_4844,N_4910);
nor UO_745 (O_745,N_4836,N_4973);
nand UO_746 (O_746,N_4824,N_4889);
nand UO_747 (O_747,N_4851,N_4856);
nor UO_748 (O_748,N_4959,N_4931);
or UO_749 (O_749,N_4962,N_4970);
and UO_750 (O_750,N_4812,N_4995);
nand UO_751 (O_751,N_4810,N_4938);
nor UO_752 (O_752,N_4942,N_4856);
or UO_753 (O_753,N_4856,N_4944);
and UO_754 (O_754,N_4997,N_4815);
nand UO_755 (O_755,N_4864,N_4911);
xor UO_756 (O_756,N_4915,N_4940);
and UO_757 (O_757,N_4826,N_4939);
nor UO_758 (O_758,N_4920,N_4817);
nand UO_759 (O_759,N_4867,N_4973);
and UO_760 (O_760,N_4866,N_4983);
or UO_761 (O_761,N_4922,N_4966);
nand UO_762 (O_762,N_4877,N_4846);
nor UO_763 (O_763,N_4972,N_4874);
nor UO_764 (O_764,N_4888,N_4991);
nand UO_765 (O_765,N_4973,N_4966);
and UO_766 (O_766,N_4935,N_4944);
and UO_767 (O_767,N_4919,N_4832);
nor UO_768 (O_768,N_4946,N_4859);
and UO_769 (O_769,N_4911,N_4866);
xnor UO_770 (O_770,N_4869,N_4940);
nor UO_771 (O_771,N_4943,N_4966);
nand UO_772 (O_772,N_4934,N_4894);
xor UO_773 (O_773,N_4924,N_4902);
and UO_774 (O_774,N_4839,N_4986);
and UO_775 (O_775,N_4846,N_4882);
or UO_776 (O_776,N_4914,N_4957);
nand UO_777 (O_777,N_4967,N_4838);
and UO_778 (O_778,N_4823,N_4977);
nor UO_779 (O_779,N_4875,N_4838);
or UO_780 (O_780,N_4930,N_4823);
nor UO_781 (O_781,N_4820,N_4976);
nor UO_782 (O_782,N_4802,N_4866);
and UO_783 (O_783,N_4802,N_4879);
nand UO_784 (O_784,N_4809,N_4801);
nor UO_785 (O_785,N_4877,N_4984);
and UO_786 (O_786,N_4827,N_4955);
xnor UO_787 (O_787,N_4876,N_4908);
and UO_788 (O_788,N_4806,N_4834);
and UO_789 (O_789,N_4972,N_4840);
or UO_790 (O_790,N_4969,N_4989);
nand UO_791 (O_791,N_4910,N_4987);
nor UO_792 (O_792,N_4869,N_4854);
and UO_793 (O_793,N_4997,N_4931);
or UO_794 (O_794,N_4943,N_4950);
or UO_795 (O_795,N_4967,N_4943);
and UO_796 (O_796,N_4802,N_4846);
nand UO_797 (O_797,N_4944,N_4883);
nand UO_798 (O_798,N_4925,N_4988);
and UO_799 (O_799,N_4891,N_4880);
or UO_800 (O_800,N_4992,N_4955);
or UO_801 (O_801,N_4919,N_4938);
nand UO_802 (O_802,N_4898,N_4999);
nand UO_803 (O_803,N_4825,N_4910);
or UO_804 (O_804,N_4903,N_4953);
nor UO_805 (O_805,N_4987,N_4990);
and UO_806 (O_806,N_4923,N_4951);
nor UO_807 (O_807,N_4806,N_4880);
and UO_808 (O_808,N_4993,N_4881);
xor UO_809 (O_809,N_4860,N_4834);
or UO_810 (O_810,N_4820,N_4959);
or UO_811 (O_811,N_4879,N_4969);
or UO_812 (O_812,N_4820,N_4814);
or UO_813 (O_813,N_4946,N_4911);
and UO_814 (O_814,N_4843,N_4949);
nand UO_815 (O_815,N_4922,N_4851);
nor UO_816 (O_816,N_4991,N_4877);
and UO_817 (O_817,N_4968,N_4889);
or UO_818 (O_818,N_4866,N_4842);
or UO_819 (O_819,N_4859,N_4806);
nor UO_820 (O_820,N_4828,N_4987);
nand UO_821 (O_821,N_4966,N_4850);
xor UO_822 (O_822,N_4992,N_4956);
nand UO_823 (O_823,N_4937,N_4935);
nand UO_824 (O_824,N_4850,N_4916);
nand UO_825 (O_825,N_4819,N_4894);
xnor UO_826 (O_826,N_4962,N_4957);
and UO_827 (O_827,N_4883,N_4888);
nand UO_828 (O_828,N_4956,N_4851);
nand UO_829 (O_829,N_4840,N_4970);
nor UO_830 (O_830,N_4946,N_4902);
xnor UO_831 (O_831,N_4818,N_4988);
xor UO_832 (O_832,N_4909,N_4876);
nand UO_833 (O_833,N_4938,N_4867);
nor UO_834 (O_834,N_4848,N_4895);
nand UO_835 (O_835,N_4915,N_4933);
nor UO_836 (O_836,N_4875,N_4860);
nand UO_837 (O_837,N_4823,N_4901);
nand UO_838 (O_838,N_4805,N_4860);
or UO_839 (O_839,N_4941,N_4891);
and UO_840 (O_840,N_4825,N_4972);
or UO_841 (O_841,N_4839,N_4967);
or UO_842 (O_842,N_4983,N_4894);
or UO_843 (O_843,N_4991,N_4970);
nand UO_844 (O_844,N_4827,N_4874);
nor UO_845 (O_845,N_4815,N_4996);
or UO_846 (O_846,N_4951,N_4832);
nor UO_847 (O_847,N_4876,N_4940);
nor UO_848 (O_848,N_4830,N_4851);
or UO_849 (O_849,N_4924,N_4806);
nor UO_850 (O_850,N_4888,N_4822);
nand UO_851 (O_851,N_4854,N_4804);
and UO_852 (O_852,N_4800,N_4837);
nand UO_853 (O_853,N_4910,N_4885);
nor UO_854 (O_854,N_4969,N_4867);
nand UO_855 (O_855,N_4887,N_4823);
nand UO_856 (O_856,N_4909,N_4966);
nor UO_857 (O_857,N_4975,N_4890);
and UO_858 (O_858,N_4914,N_4910);
or UO_859 (O_859,N_4852,N_4920);
nor UO_860 (O_860,N_4984,N_4847);
or UO_861 (O_861,N_4866,N_4975);
nand UO_862 (O_862,N_4878,N_4806);
nand UO_863 (O_863,N_4884,N_4847);
and UO_864 (O_864,N_4823,N_4972);
nand UO_865 (O_865,N_4910,N_4951);
and UO_866 (O_866,N_4909,N_4897);
nand UO_867 (O_867,N_4945,N_4839);
or UO_868 (O_868,N_4805,N_4861);
nor UO_869 (O_869,N_4891,N_4848);
and UO_870 (O_870,N_4809,N_4948);
or UO_871 (O_871,N_4812,N_4951);
nor UO_872 (O_872,N_4865,N_4987);
nand UO_873 (O_873,N_4806,N_4910);
or UO_874 (O_874,N_4984,N_4897);
nand UO_875 (O_875,N_4891,N_4863);
or UO_876 (O_876,N_4830,N_4800);
and UO_877 (O_877,N_4974,N_4844);
nor UO_878 (O_878,N_4871,N_4953);
nor UO_879 (O_879,N_4806,N_4852);
or UO_880 (O_880,N_4870,N_4845);
nor UO_881 (O_881,N_4834,N_4813);
and UO_882 (O_882,N_4987,N_4909);
nor UO_883 (O_883,N_4918,N_4968);
xnor UO_884 (O_884,N_4937,N_4874);
nor UO_885 (O_885,N_4997,N_4939);
or UO_886 (O_886,N_4951,N_4852);
xnor UO_887 (O_887,N_4859,N_4963);
nor UO_888 (O_888,N_4858,N_4825);
nor UO_889 (O_889,N_4807,N_4923);
nand UO_890 (O_890,N_4913,N_4963);
nand UO_891 (O_891,N_4935,N_4906);
nor UO_892 (O_892,N_4845,N_4827);
xor UO_893 (O_893,N_4831,N_4974);
nor UO_894 (O_894,N_4991,N_4841);
nor UO_895 (O_895,N_4816,N_4854);
nand UO_896 (O_896,N_4815,N_4880);
nor UO_897 (O_897,N_4839,N_4980);
and UO_898 (O_898,N_4984,N_4842);
nor UO_899 (O_899,N_4918,N_4879);
and UO_900 (O_900,N_4848,N_4923);
or UO_901 (O_901,N_4852,N_4819);
nand UO_902 (O_902,N_4927,N_4907);
nor UO_903 (O_903,N_4972,N_4895);
nor UO_904 (O_904,N_4933,N_4959);
or UO_905 (O_905,N_4832,N_4988);
nand UO_906 (O_906,N_4841,N_4807);
and UO_907 (O_907,N_4949,N_4903);
nand UO_908 (O_908,N_4880,N_4818);
or UO_909 (O_909,N_4929,N_4862);
or UO_910 (O_910,N_4808,N_4849);
nand UO_911 (O_911,N_4866,N_4834);
or UO_912 (O_912,N_4804,N_4928);
nor UO_913 (O_913,N_4901,N_4997);
nor UO_914 (O_914,N_4918,N_4981);
or UO_915 (O_915,N_4859,N_4883);
nor UO_916 (O_916,N_4899,N_4892);
nand UO_917 (O_917,N_4984,N_4967);
or UO_918 (O_918,N_4840,N_4863);
nand UO_919 (O_919,N_4967,N_4814);
and UO_920 (O_920,N_4988,N_4971);
and UO_921 (O_921,N_4846,N_4862);
and UO_922 (O_922,N_4879,N_4937);
nand UO_923 (O_923,N_4880,N_4990);
nand UO_924 (O_924,N_4820,N_4800);
nor UO_925 (O_925,N_4801,N_4879);
and UO_926 (O_926,N_4924,N_4820);
and UO_927 (O_927,N_4838,N_4832);
nand UO_928 (O_928,N_4838,N_4810);
nor UO_929 (O_929,N_4914,N_4915);
or UO_930 (O_930,N_4935,N_4986);
nor UO_931 (O_931,N_4892,N_4833);
or UO_932 (O_932,N_4842,N_4874);
or UO_933 (O_933,N_4860,N_4864);
and UO_934 (O_934,N_4929,N_4834);
and UO_935 (O_935,N_4845,N_4865);
nand UO_936 (O_936,N_4921,N_4976);
nand UO_937 (O_937,N_4996,N_4858);
or UO_938 (O_938,N_4970,N_4998);
nand UO_939 (O_939,N_4959,N_4954);
or UO_940 (O_940,N_4881,N_4974);
or UO_941 (O_941,N_4928,N_4916);
nor UO_942 (O_942,N_4928,N_4861);
or UO_943 (O_943,N_4956,N_4870);
xor UO_944 (O_944,N_4819,N_4878);
or UO_945 (O_945,N_4816,N_4814);
nor UO_946 (O_946,N_4981,N_4934);
and UO_947 (O_947,N_4900,N_4977);
nand UO_948 (O_948,N_4894,N_4974);
or UO_949 (O_949,N_4937,N_4812);
nor UO_950 (O_950,N_4929,N_4903);
and UO_951 (O_951,N_4940,N_4890);
or UO_952 (O_952,N_4965,N_4933);
and UO_953 (O_953,N_4918,N_4875);
xor UO_954 (O_954,N_4920,N_4971);
nor UO_955 (O_955,N_4867,N_4823);
nand UO_956 (O_956,N_4938,N_4905);
and UO_957 (O_957,N_4932,N_4907);
or UO_958 (O_958,N_4903,N_4947);
and UO_959 (O_959,N_4988,N_4950);
and UO_960 (O_960,N_4857,N_4827);
and UO_961 (O_961,N_4825,N_4990);
xor UO_962 (O_962,N_4936,N_4822);
nand UO_963 (O_963,N_4931,N_4837);
and UO_964 (O_964,N_4825,N_4833);
nand UO_965 (O_965,N_4869,N_4894);
and UO_966 (O_966,N_4807,N_4881);
nor UO_967 (O_967,N_4979,N_4810);
nand UO_968 (O_968,N_4864,N_4969);
and UO_969 (O_969,N_4814,N_4954);
xor UO_970 (O_970,N_4857,N_4801);
xor UO_971 (O_971,N_4852,N_4802);
and UO_972 (O_972,N_4930,N_4975);
nor UO_973 (O_973,N_4891,N_4811);
nor UO_974 (O_974,N_4924,N_4935);
nor UO_975 (O_975,N_4995,N_4889);
nand UO_976 (O_976,N_4968,N_4858);
or UO_977 (O_977,N_4961,N_4922);
nand UO_978 (O_978,N_4924,N_4848);
xnor UO_979 (O_979,N_4932,N_4809);
nor UO_980 (O_980,N_4945,N_4894);
xor UO_981 (O_981,N_4867,N_4846);
nor UO_982 (O_982,N_4926,N_4806);
nand UO_983 (O_983,N_4975,N_4892);
or UO_984 (O_984,N_4890,N_4808);
nand UO_985 (O_985,N_4962,N_4980);
nand UO_986 (O_986,N_4922,N_4943);
xnor UO_987 (O_987,N_4882,N_4925);
xnor UO_988 (O_988,N_4857,N_4921);
or UO_989 (O_989,N_4820,N_4862);
nand UO_990 (O_990,N_4887,N_4941);
xnor UO_991 (O_991,N_4996,N_4804);
or UO_992 (O_992,N_4965,N_4841);
or UO_993 (O_993,N_4931,N_4881);
nor UO_994 (O_994,N_4847,N_4963);
nor UO_995 (O_995,N_4958,N_4814);
xnor UO_996 (O_996,N_4806,N_4908);
or UO_997 (O_997,N_4862,N_4976);
nor UO_998 (O_998,N_4886,N_4865);
nand UO_999 (O_999,N_4862,N_4874);
endmodule