module basic_1500_15000_2000_3_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10010,N_10011,N_10012,N_10014,N_10016,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10026,N_10027,N_10028,N_10029,N_10031,N_10032,N_10033,N_10034,N_10035,N_10038,N_10039,N_10040,N_10041,N_10043,N_10044,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10088,N_10090,N_10091,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10100,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10118,N_10119,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10134,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10143,N_10144,N_10145,N_10147,N_10148,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10159,N_10160,N_10161,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10192,N_10193,N_10194,N_10196,N_10198,N_10199,N_10200,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10226,N_10228,N_10230,N_10231,N_10232,N_10233,N_10235,N_10236,N_10237,N_10238,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10251,N_10252,N_10254,N_10256,N_10257,N_10259,N_10261,N_10265,N_10266,N_10267,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10304,N_10306,N_10307,N_10309,N_10310,N_10312,N_10313,N_10315,N_10316,N_10317,N_10318,N_10319,N_10321,N_10322,N_10323,N_10324,N_10326,N_10327,N_10329,N_10330,N_10332,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10355,N_10356,N_10357,N_10359,N_10360,N_10361,N_10362,N_10363,N_10365,N_10368,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10381,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10391,N_10392,N_10393,N_10394,N_10396,N_10397,N_10398,N_10400,N_10402,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10419,N_10420,N_10421,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10447,N_10451,N_10452,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10464,N_10466,N_10467,N_10468,N_10469,N_10471,N_10472,N_10473,N_10474,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10488,N_10489,N_10490,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10518,N_10520,N_10521,N_10522,N_10523,N_10524,N_10527,N_10528,N_10530,N_10531,N_10535,N_10536,N_10537,N_10538,N_10539,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10551,N_10552,N_10553,N_10555,N_10557,N_10558,N_10560,N_10561,N_10562,N_10563,N_10564,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10588,N_10589,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10629,N_10630,N_10632,N_10633,N_10635,N_10637,N_10638,N_10640,N_10641,N_10642,N_10643,N_10644,N_10646,N_10648,N_10650,N_10652,N_10653,N_10654,N_10655,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10677,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10687,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10697,N_10698,N_10699,N_10701,N_10703,N_10704,N_10705,N_10706,N_10707,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10762,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10778,N_10779,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10793,N_10794,N_10796,N_10798,N_10799,N_10800,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10819,N_10820,N_10821,N_10822,N_10823,N_10825,N_10826,N_10827,N_10828,N_10829,N_10831,N_10832,N_10833,N_10834,N_10835,N_10838,N_10839,N_10840,N_10841,N_10842,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10858,N_10859,N_10860,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10878,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10891,N_10892,N_10893,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10934,N_10935,N_10937,N_10938,N_10939,N_10940,N_10942,N_10943,N_10945,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10969,N_10970,N_10971,N_10973,N_10974,N_10975,N_10976,N_10977,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10987,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10997,N_10998,N_10999,N_11000,N_11002,N_11003,N_11004,N_11006,N_11007,N_11008,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11021,N_11024,N_11025,N_11026,N_11027,N_11029,N_11030,N_11031,N_11032,N_11033,N_11035,N_11036,N_11037,N_11039,N_11040,N_11041,N_11043,N_11044,N_11046,N_11047,N_11049,N_11050,N_11051,N_11052,N_11053,N_11055,N_11056,N_11057,N_11058,N_11059,N_11062,N_11063,N_11064,N_11065,N_11067,N_11068,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11077,N_11078,N_11079,N_11080,N_11083,N_11084,N_11085,N_11086,N_11087,N_11090,N_11091,N_11093,N_11094,N_11095,N_11098,N_11099,N_11100,N_11101,N_11103,N_11104,N_11105,N_11106,N_11107,N_11110,N_11111,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11134,N_11136,N_11137,N_11139,N_11140,N_11141,N_11142,N_11144,N_11145,N_11147,N_11149,N_11152,N_11153,N_11154,N_11155,N_11157,N_11158,N_11159,N_11161,N_11162,N_11163,N_11164,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11190,N_11191,N_11192,N_11194,N_11197,N_11198,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11207,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11230,N_11231,N_11232,N_11234,N_11235,N_11236,N_11240,N_11241,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11251,N_11252,N_11253,N_11254,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11263,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11303,N_11304,N_11305,N_11306,N_11307,N_11309,N_11311,N_11312,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11326,N_11327,N_11328,N_11330,N_11331,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11343,N_11344,N_11345,N_11346,N_11349,N_11350,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11360,N_11361,N_11362,N_11363,N_11365,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11393,N_11394,N_11395,N_11396,N_11398,N_11399,N_11400,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11419,N_11421,N_11422,N_11423,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11443,N_11444,N_11445,N_11447,N_11449,N_11451,N_11452,N_11453,N_11454,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11469,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11479,N_11481,N_11482,N_11483,N_11484,N_11485,N_11487,N_11488,N_11489,N_11490,N_11492,N_11494,N_11495,N_11496,N_11498,N_11499,N_11500,N_11501,N_11502,N_11504,N_11505,N_11506,N_11507,N_11509,N_11510,N_11511,N_11513,N_11515,N_11516,N_11518,N_11519,N_11522,N_11524,N_11525,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11536,N_11537,N_11538,N_11542,N_11544,N_11545,N_11546,N_11548,N_11549,N_11551,N_11552,N_11555,N_11556,N_11557,N_11558,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11570,N_11571,N_11572,N_11573,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11593,N_11594,N_11595,N_11596,N_11598,N_11599,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11619,N_11621,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11648,N_11649,N_11650,N_11652,N_11653,N_11655,N_11656,N_11658,N_11659,N_11660,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11685,N_11686,N_11690,N_11692,N_11693,N_11694,N_11695,N_11696,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11723,N_11724,N_11725,N_11726,N_11727,N_11729,N_11731,N_11732,N_11733,N_11734,N_11736,N_11737,N_11738,N_11739,N_11740,N_11743,N_11745,N_11746,N_11747,N_11749,N_11750,N_11752,N_11753,N_11754,N_11755,N_11756,N_11758,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11780,N_11781,N_11782,N_11783,N_11784,N_11786,N_11787,N_11788,N_11789,N_11790,N_11793,N_11794,N_11800,N_11801,N_11802,N_11803,N_11804,N_11808,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11818,N_11819,N_11820,N_11822,N_11823,N_11824,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11834,N_11835,N_11837,N_11839,N_11840,N_11841,N_11842,N_11844,N_11846,N_11847,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11883,N_11884,N_11886,N_11887,N_11888,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11915,N_11917,N_11919,N_11920,N_11921,N_11922,N_11924,N_11925,N_11926,N_11927,N_11928,N_11930,N_11931,N_11932,N_11934,N_11935,N_11936,N_11937,N_11938,N_11940,N_11941,N_11942,N_11943,N_11945,N_11946,N_11947,N_11950,N_11951,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11969,N_11971,N_11972,N_11973,N_11974,N_11975,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11985,N_11986,N_11987,N_11989,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12011,N_12012,N_12013,N_12015,N_12017,N_12018,N_12019,N_12021,N_12023,N_12024,N_12027,N_12029,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12059,N_12060,N_12061,N_12062,N_12064,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12075,N_12076,N_12077,N_12078,N_12079,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12100,N_12101,N_12103,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12112,N_12113,N_12115,N_12117,N_12118,N_12119,N_12120,N_12121,N_12123,N_12124,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12134,N_12136,N_12137,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12157,N_12158,N_12159,N_12160,N_12163,N_12164,N_12166,N_12167,N_12168,N_12170,N_12172,N_12173,N_12174,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12188,N_12189,N_12191,N_12192,N_12193,N_12194,N_12195,N_12197,N_12198,N_12199,N_12200,N_12202,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12216,N_12217,N_12218,N_12219,N_12221,N_12222,N_12224,N_12225,N_12227,N_12228,N_12229,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12247,N_12248,N_12249,N_12250,N_12252,N_12254,N_12256,N_12257,N_12259,N_12260,N_12262,N_12263,N_12264,N_12266,N_12267,N_12268,N_12269,N_12271,N_12272,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12282,N_12283,N_12285,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12305,N_12306,N_12307,N_12308,N_12310,N_12311,N_12312,N_12313,N_12314,N_12316,N_12317,N_12319,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12329,N_12330,N_12332,N_12333,N_12335,N_12337,N_12338,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12347,N_12348,N_12349,N_12350,N_12352,N_12354,N_12356,N_12357,N_12358,N_12359,N_12360,N_12363,N_12364,N_12365,N_12366,N_12369,N_12371,N_12372,N_12373,N_12374,N_12377,N_12378,N_12380,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12396,N_12397,N_12398,N_12400,N_12401,N_12402,N_12403,N_12404,N_12406,N_12407,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12428,N_12430,N_12432,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12446,N_12447,N_12449,N_12450,N_12451,N_12452,N_12454,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12481,N_12482,N_12484,N_12486,N_12488,N_12490,N_12493,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12525,N_12526,N_12527,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12542,N_12543,N_12544,N_12546,N_12547,N_12548,N_12549,N_12551,N_12552,N_12553,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12566,N_12567,N_12568,N_12570,N_12571,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12593,N_12594,N_12595,N_12598,N_12599,N_12600,N_12601,N_12602,N_12604,N_12605,N_12607,N_12608,N_12609,N_12610,N_12611,N_12613,N_12614,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12626,N_12627,N_12628,N_12631,N_12632,N_12633,N_12634,N_12635,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12670,N_12672,N_12673,N_12674,N_12675,N_12676,N_12678,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12690,N_12692,N_12693,N_12694,N_12695,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12718,N_12719,N_12720,N_12721,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12732,N_12733,N_12734,N_12735,N_12737,N_12738,N_12739,N_12740,N_12741,N_12743,N_12744,N_12745,N_12746,N_12748,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12766,N_12768,N_12769,N_12770,N_12771,N_12772,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12801,N_12803,N_12804,N_12805,N_12807,N_12809,N_12810,N_12812,N_12813,N_12815,N_12816,N_12817,N_12818,N_12819,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12857,N_12858,N_12859,N_12861,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12872,N_12873,N_12874,N_12875,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12889,N_12890,N_12891,N_12892,N_12893,N_12895,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12934,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12945,N_12946,N_12947,N_12948,N_12950,N_12951,N_12954,N_12955,N_12956,N_12957,N_12958,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12972,N_12973,N_12974,N_12975,N_12976,N_12978,N_12979,N_12980,N_12981,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12994,N_12995,N_12997,N_12999,N_13000,N_13001,N_13002,N_13004,N_13005,N_13006,N_13007,N_13008,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13030,N_13032,N_13033,N_13035,N_13036,N_13037,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13061,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13090,N_13092,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13135,N_13137,N_13138,N_13139,N_13140,N_13143,N_13144,N_13145,N_13147,N_13148,N_13149,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13166,N_13167,N_13168,N_13170,N_13171,N_13172,N_13173,N_13174,N_13176,N_13178,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13190,N_13191,N_13192,N_13193,N_13194,N_13197,N_13198,N_13199,N_13200,N_13201,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13216,N_13217,N_13219,N_13220,N_13222,N_13223,N_13224,N_13225,N_13227,N_13228,N_13229,N_13230,N_13232,N_13233,N_13234,N_13235,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13251,N_13252,N_13253,N_13254,N_13255,N_13257,N_13258,N_13259,N_13260,N_13261,N_13264,N_13265,N_13266,N_13267,N_13268,N_13270,N_13271,N_13274,N_13275,N_13276,N_13277,N_13278,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13300,N_13302,N_13303,N_13304,N_13305,N_13306,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13317,N_13318,N_13319,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13332,N_13334,N_13335,N_13338,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13351,N_13352,N_13354,N_13355,N_13357,N_13360,N_13361,N_13362,N_13364,N_13365,N_13366,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13376,N_13377,N_13378,N_13379,N_13380,N_13382,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13406,N_13407,N_13408,N_13409,N_13410,N_13412,N_13413,N_13414,N_13415,N_13416,N_13418,N_13419,N_13421,N_13422,N_13424,N_13425,N_13426,N_13427,N_13429,N_13430,N_13432,N_13433,N_13434,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13453,N_13454,N_13455,N_13457,N_13458,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13482,N_13483,N_13484,N_13485,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13500,N_13502,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13536,N_13537,N_13538,N_13539,N_13540,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13560,N_13562,N_13565,N_13566,N_13567,N_13568,N_13571,N_13572,N_13573,N_13575,N_13576,N_13577,N_13578,N_13579,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13589,N_13590,N_13591,N_13593,N_13594,N_13596,N_13597,N_13598,N_13600,N_13601,N_13602,N_13603,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13625,N_13626,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13637,N_13638,N_13639,N_13640,N_13641,N_13644,N_13645,N_13647,N_13648,N_13649,N_13651,N_13652,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13679,N_13680,N_13681,N_13683,N_13684,N_13685,N_13686,N_13687,N_13689,N_13691,N_13692,N_13694,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13714,N_13717,N_13718,N_13719,N_13721,N_13722,N_13723,N_13724,N_13725,N_13727,N_13728,N_13729,N_13733,N_13734,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13748,N_13749,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13766,N_13767,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13791,N_13792,N_13794,N_13796,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13829,N_13831,N_13832,N_13833,N_13835,N_13836,N_13838,N_13839,N_13840,N_13841,N_13842,N_13847,N_13848,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13864,N_13865,N_13867,N_13868,N_13870,N_13871,N_13872,N_13874,N_13875,N_13876,N_13878,N_13879,N_13880,N_13881,N_13882,N_13886,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13897,N_13898,N_13900,N_13902,N_13904,N_13905,N_13906,N_13907,N_13910,N_13911,N_13912,N_13913,N_13914,N_13916,N_13917,N_13918,N_13920,N_13921,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13939,N_13940,N_13941,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13963,N_13964,N_13967,N_13968,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13977,N_13978,N_13979,N_13980,N_13981,N_13983,N_13984,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13995,N_13996,N_13997,N_13999,N_14000,N_14001,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14022,N_14024,N_14025,N_14026,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14039,N_14040,N_14041,N_14043,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14053,N_14054,N_14057,N_14058,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14075,N_14077,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14090,N_14092,N_14093,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14120,N_14121,N_14122,N_14123,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14135,N_14136,N_14140,N_14141,N_14142,N_14144,N_14145,N_14146,N_14147,N_14149,N_14150,N_14152,N_14153,N_14155,N_14156,N_14158,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14183,N_14184,N_14185,N_14186,N_14189,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14206,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14218,N_14219,N_14221,N_14223,N_14224,N_14225,N_14226,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14238,N_14239,N_14240,N_14242,N_14243,N_14244,N_14247,N_14249,N_14250,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14260,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14272,N_14273,N_14274,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14288,N_14289,N_14290,N_14291,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14307,N_14308,N_14309,N_14310,N_14311,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14327,N_14328,N_14329,N_14330,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14339,N_14340,N_14341,N_14343,N_14344,N_14345,N_14346,N_14347,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14365,N_14368,N_14369,N_14370,N_14371,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14400,N_14402,N_14404,N_14405,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14416,N_14417,N_14418,N_14419,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14442,N_14443,N_14445,N_14448,N_14449,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14458,N_14459,N_14460,N_14461,N_14463,N_14464,N_14465,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14474,N_14476,N_14478,N_14479,N_14480,N_14481,N_14482,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14491,N_14492,N_14493,N_14494,N_14497,N_14499,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14509,N_14510,N_14511,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14531,N_14532,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14544,N_14545,N_14546,N_14547,N_14549,N_14551,N_14552,N_14553,N_14554,N_14556,N_14557,N_14558,N_14559,N_14561,N_14562,N_14563,N_14565,N_14566,N_14567,N_14568,N_14569,N_14571,N_14572,N_14573,N_14574,N_14577,N_14579,N_14581,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14589,N_14590,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14600,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14613,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14627,N_14629,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14643,N_14644,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14656,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14665,N_14666,N_14667,N_14668,N_14669,N_14672,N_14673,N_14674,N_14675,N_14677,N_14678,N_14679,N_14680,N_14681,N_14683,N_14684,N_14685,N_14686,N_14687,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14749,N_14750,N_14751,N_14752,N_14753,N_14755,N_14756,N_14757,N_14758,N_14760,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14773,N_14774,N_14775,N_14776,N_14777,N_14779,N_14780,N_14781,N_14782,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14792,N_14793,N_14794,N_14795,N_14796,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14806,N_14807,N_14809,N_14810,N_14812,N_14814,N_14815,N_14816,N_14817,N_14819,N_14820,N_14821,N_14825,N_14828,N_14829,N_14832,N_14833,N_14834,N_14835,N_14836,N_14838,N_14839,N_14840,N_14841,N_14842,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14853,N_14855,N_14856,N_14857,N_14858,N_14861,N_14862,N_14863,N_14864,N_14867,N_14869,N_14870,N_14871,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14902,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14925,N_14926,N_14928,N_14929,N_14931,N_14933,N_14935,N_14936,N_14938,N_14940,N_14941,N_14942,N_14944,N_14945,N_14946,N_14947,N_14948,N_14950,N_14951,N_14952,N_14953,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14965,N_14967,N_14968,N_14969,N_14970,N_14972,N_14974,N_14975,N_14976,N_14977,N_14980,N_14982,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_282,In_1332);
nand U1 (N_1,In_778,In_803);
and U2 (N_2,In_1109,In_110);
nand U3 (N_3,In_574,In_1015);
and U4 (N_4,In_1327,In_1044);
and U5 (N_5,In_203,In_1482);
and U6 (N_6,In_1423,In_664);
or U7 (N_7,In_1008,In_1091);
and U8 (N_8,In_908,In_169);
or U9 (N_9,In_504,In_1235);
nand U10 (N_10,In_1020,In_997);
and U11 (N_11,In_1284,In_724);
or U12 (N_12,In_1022,In_103);
xor U13 (N_13,In_928,In_1282);
nand U14 (N_14,In_660,In_1037);
nand U15 (N_15,In_880,In_335);
nor U16 (N_16,In_1182,In_1442);
and U17 (N_17,In_1330,In_460);
nor U18 (N_18,In_349,In_693);
nand U19 (N_19,In_108,In_590);
and U20 (N_20,In_163,In_999);
or U21 (N_21,In_210,In_632);
nand U22 (N_22,In_1036,In_1387);
nor U23 (N_23,In_1280,In_529);
and U24 (N_24,In_1033,In_856);
or U25 (N_25,In_961,In_1121);
nand U26 (N_26,In_1093,In_909);
or U27 (N_27,In_937,In_1353);
or U28 (N_28,In_1427,In_138);
nand U29 (N_29,In_618,In_600);
nand U30 (N_30,In_1187,In_742);
or U31 (N_31,In_982,In_1207);
nor U32 (N_32,In_17,In_1127);
nand U33 (N_33,In_1231,In_76);
nor U34 (N_34,In_667,In_125);
nand U35 (N_35,In_1463,In_881);
nand U36 (N_36,In_415,In_680);
nand U37 (N_37,In_1276,In_53);
nor U38 (N_38,In_1234,In_1339);
nand U39 (N_39,In_967,In_554);
or U40 (N_40,In_261,In_508);
nand U41 (N_41,In_551,In_850);
or U42 (N_42,In_95,In_863);
and U43 (N_43,In_20,In_388);
and U44 (N_44,In_309,In_322);
or U45 (N_45,In_440,In_1081);
or U46 (N_46,In_375,In_1270);
nand U47 (N_47,In_932,In_283);
nand U48 (N_48,In_1242,In_1324);
and U49 (N_49,In_621,In_754);
or U50 (N_50,In_289,In_100);
nor U51 (N_51,In_740,In_1341);
nand U52 (N_52,In_1023,In_979);
and U53 (N_53,In_1455,In_66);
nor U54 (N_54,In_264,In_1135);
or U55 (N_55,In_1138,In_1417);
and U56 (N_56,In_471,In_109);
nor U57 (N_57,In_528,In_1106);
nor U58 (N_58,In_720,In_1201);
nor U59 (N_59,In_511,In_1254);
or U60 (N_60,In_185,In_1205);
nor U61 (N_61,In_338,In_614);
nor U62 (N_62,In_1085,In_479);
nand U63 (N_63,In_1185,In_1489);
or U64 (N_64,In_1397,In_844);
xor U65 (N_65,In_975,In_430);
nor U66 (N_66,In_1395,In_780);
and U67 (N_67,In_313,In_966);
or U68 (N_68,In_382,In_73);
or U69 (N_69,In_944,In_256);
and U70 (N_70,In_752,In_358);
or U71 (N_71,In_1351,In_924);
nor U72 (N_72,In_1074,In_1133);
or U73 (N_73,In_790,In_955);
or U74 (N_74,In_348,In_1487);
and U75 (N_75,In_80,In_535);
or U76 (N_76,In_1035,In_336);
nor U77 (N_77,In_232,In_903);
and U78 (N_78,In_635,In_643);
nand U79 (N_79,In_1082,In_570);
nor U80 (N_80,In_1291,In_324);
nor U81 (N_81,In_1173,In_1430);
or U82 (N_82,In_917,In_836);
nor U83 (N_83,In_82,In_534);
and U84 (N_84,In_1272,In_1249);
nand U85 (N_85,In_255,In_821);
nand U86 (N_86,In_1010,In_1088);
or U87 (N_87,In_1432,In_211);
and U88 (N_88,In_25,In_670);
nor U89 (N_89,In_902,In_1203);
and U90 (N_90,In_661,In_68);
and U91 (N_91,In_716,In_709);
nor U92 (N_92,In_1123,In_747);
nand U93 (N_93,In_1244,In_330);
nand U94 (N_94,In_225,In_1004);
nor U95 (N_95,In_1319,In_1027);
nor U96 (N_96,In_1105,In_1401);
nand U97 (N_97,In_870,In_146);
and U98 (N_98,In_810,In_1306);
nor U99 (N_99,In_391,In_706);
nor U100 (N_100,In_1388,In_369);
nand U101 (N_101,In_353,In_875);
nand U102 (N_102,In_81,In_1287);
nand U103 (N_103,In_963,In_927);
nor U104 (N_104,In_450,In_29);
and U105 (N_105,In_978,In_459);
nor U106 (N_106,In_1099,In_804);
nor U107 (N_107,In_695,In_719);
and U108 (N_108,In_419,In_1084);
or U109 (N_109,In_187,In_1011);
xnor U110 (N_110,In_47,In_1331);
or U111 (N_111,In_594,In_265);
nand U112 (N_112,In_767,In_507);
or U113 (N_113,In_853,In_623);
and U114 (N_114,In_129,In_1160);
nand U115 (N_115,In_973,In_363);
and U116 (N_116,In_1475,In_300);
or U117 (N_117,In_320,In_646);
nor U118 (N_118,In_243,In_654);
nand U119 (N_119,In_253,In_735);
nor U120 (N_120,In_974,In_984);
nand U121 (N_121,In_1454,In_591);
nor U122 (N_122,In_140,In_698);
or U123 (N_123,In_1453,In_295);
and U124 (N_124,In_768,In_1025);
or U125 (N_125,In_1316,In_481);
nor U126 (N_126,In_1232,In_0);
and U127 (N_127,In_1309,In_372);
nor U128 (N_128,In_990,In_628);
and U129 (N_129,In_468,In_377);
nand U130 (N_130,In_565,In_123);
nand U131 (N_131,In_1165,In_820);
nor U132 (N_132,In_285,In_866);
or U133 (N_133,In_1342,In_1003);
nor U134 (N_134,In_30,In_732);
and U135 (N_135,In_823,In_241);
or U136 (N_136,In_16,In_1061);
nor U137 (N_137,In_704,In_659);
or U138 (N_138,In_5,In_23);
or U139 (N_139,In_1153,In_121);
and U140 (N_140,In_1265,In_387);
nand U141 (N_141,In_556,In_429);
nand U142 (N_142,In_173,In_687);
nor U143 (N_143,In_1223,In_354);
and U144 (N_144,In_1005,In_729);
nand U145 (N_145,In_128,In_311);
and U146 (N_146,In_1190,In_1134);
or U147 (N_147,In_819,In_452);
nand U148 (N_148,In_1049,In_1041);
and U149 (N_149,In_222,In_718);
nand U150 (N_150,In_1217,In_730);
or U151 (N_151,In_41,In_615);
nor U152 (N_152,In_1474,In_1269);
and U153 (N_153,In_1126,In_1066);
nand U154 (N_154,In_342,In_885);
nand U155 (N_155,In_624,In_35);
and U156 (N_156,In_1046,In_1381);
and U157 (N_157,In_931,In_1399);
nor U158 (N_158,In_956,In_1470);
or U159 (N_159,In_1363,In_22);
nand U160 (N_160,In_1458,In_1128);
or U161 (N_161,In_65,In_142);
nor U162 (N_162,In_492,In_52);
nand U163 (N_163,In_580,In_364);
nor U164 (N_164,In_1278,In_672);
nor U165 (N_165,In_217,In_1224);
or U166 (N_166,In_447,In_421);
and U167 (N_167,In_1444,In_287);
and U168 (N_168,In_1295,In_1189);
nand U169 (N_169,In_748,In_874);
and U170 (N_170,In_1259,In_1079);
or U171 (N_171,In_1334,In_708);
or U172 (N_172,In_1169,In_1415);
nor U173 (N_173,In_86,In_189);
or U174 (N_174,In_1196,In_784);
and U175 (N_175,In_425,In_200);
or U176 (N_176,In_948,In_1273);
or U177 (N_177,In_1321,In_51);
or U178 (N_178,In_1416,In_878);
or U179 (N_179,In_764,In_1021);
nand U180 (N_180,In_1043,In_1293);
nand U181 (N_181,In_1107,In_1304);
or U182 (N_182,In_43,In_689);
and U183 (N_183,In_872,In_1492);
nor U184 (N_184,In_1343,In_858);
or U185 (N_185,In_278,In_692);
or U186 (N_186,In_1494,In_521);
and U187 (N_187,In_861,In_1053);
and U188 (N_188,In_463,In_549);
nand U189 (N_189,In_94,In_770);
and U190 (N_190,In_734,In_470);
and U191 (N_191,In_912,In_525);
nor U192 (N_192,In_947,In_454);
or U193 (N_193,In_771,In_1132);
and U194 (N_194,In_1443,In_490);
and U195 (N_195,In_299,In_416);
and U196 (N_196,In_906,In_677);
nand U197 (N_197,In_325,In_1446);
and U198 (N_198,In_33,In_393);
or U199 (N_199,In_604,In_40);
nor U200 (N_200,In_207,In_464);
nand U201 (N_201,In_1400,In_188);
or U202 (N_202,In_88,In_276);
nand U203 (N_203,In_582,In_1377);
nor U204 (N_204,In_1407,In_1409);
nand U205 (N_205,In_316,In_18);
nor U206 (N_206,In_1239,In_376);
nand U207 (N_207,In_1420,In_1226);
nor U208 (N_208,In_157,In_321);
or U209 (N_209,In_337,In_250);
or U210 (N_210,In_1448,In_36);
and U211 (N_211,In_550,In_1083);
nand U212 (N_212,In_845,In_1472);
nor U213 (N_213,In_1161,In_1411);
nand U214 (N_214,In_352,In_736);
nor U215 (N_215,In_1250,In_1002);
and U216 (N_216,In_238,In_402);
nand U217 (N_217,In_964,In_114);
xnor U218 (N_218,In_487,In_559);
nor U219 (N_219,In_1001,In_512);
and U220 (N_220,In_1206,In_343);
nand U221 (N_221,In_763,In_1271);
and U222 (N_222,In_132,In_616);
or U223 (N_223,In_150,In_1118);
and U224 (N_224,In_294,In_45);
nand U225 (N_225,In_789,In_921);
nor U226 (N_226,In_894,In_1108);
and U227 (N_227,In_996,In_977);
or U228 (N_228,In_674,In_1092);
and U229 (N_229,In_260,In_972);
nand U230 (N_230,In_562,In_331);
and U231 (N_231,In_1275,In_1335);
and U232 (N_232,In_777,In_1318);
or U233 (N_233,In_603,In_1240);
and U234 (N_234,In_746,In_830);
nor U235 (N_235,In_539,In_523);
and U236 (N_236,In_236,In_1302);
and U237 (N_237,In_650,In_1426);
and U238 (N_238,In_543,In_758);
nor U239 (N_239,In_1499,In_705);
or U240 (N_240,In_1452,In_153);
and U241 (N_241,In_597,In_1016);
or U242 (N_242,In_1243,In_1218);
nand U243 (N_243,In_293,In_1398);
and U244 (N_244,In_1439,In_892);
nand U245 (N_245,In_8,In_1345);
and U246 (N_246,In_1204,In_1305);
nand U247 (N_247,In_514,In_398);
and U248 (N_248,In_1264,In_914);
nand U249 (N_249,In_1166,In_969);
or U250 (N_250,In_957,In_1054);
and U251 (N_251,In_801,In_254);
or U252 (N_252,In_195,In_658);
nand U253 (N_253,In_449,In_433);
and U254 (N_254,In_198,In_587);
and U255 (N_255,In_496,In_1300);
nor U256 (N_256,In_71,In_346);
nand U257 (N_257,In_531,In_945);
nor U258 (N_258,In_572,In_905);
or U259 (N_259,In_405,In_1373);
nand U260 (N_260,In_373,In_1137);
nand U261 (N_261,In_1157,In_1198);
nand U262 (N_262,In_808,In_141);
nand U263 (N_263,In_1122,In_782);
nand U264 (N_264,In_394,In_542);
nor U265 (N_265,In_831,In_893);
nand U266 (N_266,In_537,In_759);
nand U267 (N_267,In_149,In_249);
and U268 (N_268,In_31,In_179);
nand U269 (N_269,In_783,In_867);
nor U270 (N_270,In_196,In_133);
xor U271 (N_271,In_1298,In_351);
nand U272 (N_272,In_599,In_1145);
nor U273 (N_273,In_1063,In_1466);
or U274 (N_274,In_1119,In_569);
nand U275 (N_275,In_929,In_818);
and U276 (N_276,In_710,In_1162);
nor U277 (N_277,In_682,In_798);
or U278 (N_278,In_242,In_1140);
nand U279 (N_279,In_446,In_1155);
nand U280 (N_280,In_292,In_87);
or U281 (N_281,In_949,In_315);
and U282 (N_282,In_883,In_988);
and U283 (N_283,In_1315,In_381);
nand U284 (N_284,In_1497,In_199);
nor U285 (N_285,In_205,In_50);
nand U286 (N_286,In_77,In_291);
and U287 (N_287,In_923,In_1404);
and U288 (N_288,In_1178,In_1307);
nand U289 (N_289,In_1,In_1195);
and U290 (N_290,In_1357,In_715);
nor U291 (N_291,In_1139,In_1013);
nor U292 (N_292,In_700,In_319);
or U293 (N_293,In_1480,In_1086);
or U294 (N_294,In_466,In_1256);
and U295 (N_295,In_1104,In_1263);
nor U296 (N_296,In_1051,In_467);
nand U297 (N_297,In_1422,In_474);
or U298 (N_298,In_1467,In_506);
and U299 (N_299,In_105,In_448);
or U300 (N_300,In_1247,In_1418);
nor U301 (N_301,In_1285,In_1210);
nand U302 (N_302,In_613,In_1113);
and U303 (N_303,In_378,In_575);
and U304 (N_304,In_443,In_428);
or U305 (N_305,In_1148,In_1485);
and U306 (N_306,In_277,In_1253);
nor U307 (N_307,In_1125,In_1116);
nand U308 (N_308,In_145,In_1212);
or U309 (N_309,In_432,In_965);
and U310 (N_310,In_439,In_655);
nand U311 (N_311,In_1228,In_156);
or U312 (N_312,In_773,In_1386);
or U313 (N_313,In_802,In_234);
or U314 (N_314,In_395,In_829);
or U315 (N_315,In_161,In_28);
nand U316 (N_316,In_794,In_476);
or U317 (N_317,In_608,In_1481);
nor U318 (N_318,In_1486,In_606);
nand U319 (N_319,In_540,In_1170);
and U320 (N_320,In_548,In_832);
nand U321 (N_321,In_1055,In_744);
and U322 (N_322,In_1344,In_517);
nor U323 (N_323,In_279,In_334);
and U324 (N_324,In_1408,In_1478);
or U325 (N_325,In_898,In_852);
or U326 (N_326,In_1255,In_1057);
and U327 (N_327,In_204,In_314);
nor U328 (N_328,In_745,In_491);
nor U329 (N_329,In_9,In_427);
and U330 (N_330,In_1364,In_183);
nand U331 (N_331,In_323,In_1413);
and U332 (N_332,In_1208,In_389);
nand U333 (N_333,In_318,In_115);
nand U334 (N_334,In_610,In_1246);
or U335 (N_335,In_805,In_411);
or U336 (N_336,In_270,In_916);
and U337 (N_337,In_135,In_126);
nor U338 (N_338,In_1156,In_669);
or U339 (N_339,In_34,In_544);
and U340 (N_340,In_1347,In_882);
and U341 (N_341,In_456,In_1031);
nand U342 (N_342,In_1009,In_175);
nor U343 (N_343,In_101,In_1117);
and U344 (N_344,In_926,In_1183);
nand U345 (N_345,In_202,In_130);
or U346 (N_346,In_1460,In_940);
nand U347 (N_347,In_873,In_647);
nor U348 (N_348,In_812,In_13);
and U349 (N_349,In_738,In_686);
nor U350 (N_350,In_939,In_879);
and U351 (N_351,In_558,In_1112);
or U352 (N_352,In_769,In_79);
nor U353 (N_353,In_1267,In_1469);
and U354 (N_354,In_557,In_953);
or U355 (N_355,In_843,In_1461);
and U356 (N_356,In_656,In_578);
or U357 (N_357,In_99,In_345);
nor U358 (N_358,In_855,In_1471);
and U359 (N_359,In_326,In_397);
nor U360 (N_360,In_530,In_1087);
or U361 (N_361,In_489,In_714);
and U362 (N_362,In_339,In_106);
nor U363 (N_363,In_365,In_159);
nand U364 (N_364,In_118,In_1392);
and U365 (N_365,In_438,In_968);
and U366 (N_366,In_1371,In_233);
nand U367 (N_367,In_1248,In_743);
nand U368 (N_368,In_596,In_685);
and U369 (N_369,In_403,In_1314);
or U370 (N_370,In_44,In_849);
or U371 (N_371,In_1152,In_435);
nand U372 (N_372,In_633,In_1167);
nor U373 (N_373,In_679,In_221);
nand U374 (N_374,In_1098,In_1177);
nand U375 (N_375,In_1312,In_987);
and U376 (N_376,In_1076,In_1144);
nor U377 (N_377,In_181,In_1360);
or U378 (N_378,In_703,In_1359);
nor U379 (N_379,In_116,In_1236);
and U380 (N_380,In_757,In_1361);
nor U381 (N_381,In_56,In_648);
or U382 (N_382,In_1019,In_341);
or U383 (N_383,In_1356,In_46);
nand U384 (N_384,In_1329,In_465);
or U385 (N_385,In_317,In_792);
and U386 (N_386,In_526,In_119);
or U387 (N_387,In_1496,In_785);
and U388 (N_388,In_174,In_1340);
nor U389 (N_389,In_148,In_1445);
or U390 (N_390,In_97,In_329);
or U391 (N_391,In_107,In_1065);
nor U392 (N_392,In_694,In_598);
nor U393 (N_393,In_1090,In_257);
or U394 (N_394,In_228,In_611);
and U395 (N_395,In_848,In_486);
and U396 (N_396,In_1326,In_359);
nand U397 (N_397,In_942,In_919);
nand U398 (N_398,In_756,In_1393);
nor U399 (N_399,In_122,In_64);
and U400 (N_400,In_824,In_859);
or U401 (N_401,In_1292,In_1241);
and U402 (N_402,In_1070,In_11);
or U403 (N_403,In_631,In_91);
nand U404 (N_404,In_1154,In_515);
nor U405 (N_405,In_884,In_147);
nor U406 (N_406,In_1096,In_1131);
nand U407 (N_407,In_1048,In_2);
nand U408 (N_408,In_407,In_1483);
or U409 (N_409,In_209,In_223);
and U410 (N_410,In_485,In_248);
or U411 (N_411,In_833,In_561);
and U412 (N_412,In_500,In_941);
nor U413 (N_413,In_1039,In_1143);
or U414 (N_414,In_431,In_842);
nor U415 (N_415,In_567,In_713);
nor U416 (N_416,In_347,In_98);
and U417 (N_417,In_1465,In_38);
nor U418 (N_418,In_568,In_208);
or U419 (N_419,In_946,In_192);
nand U420 (N_420,In_312,In_922);
nand U421 (N_421,In_627,In_665);
or U422 (N_422,In_246,In_1369);
nand U423 (N_423,In_214,In_1073);
nor U424 (N_424,In_595,In_838);
nand U425 (N_425,In_834,In_104);
nor U426 (N_426,In_1389,In_1110);
nor U427 (N_427,In_62,In_712);
and U428 (N_428,In_1075,In_1464);
nor U429 (N_429,In_612,In_1440);
xnor U430 (N_430,In_976,In_1336);
and U431 (N_431,In_418,In_1366);
or U432 (N_432,In_619,In_1493);
and U433 (N_433,In_536,In_136);
and U434 (N_434,In_96,In_1308);
nand U435 (N_435,In_482,In_268);
or U436 (N_436,In_1346,In_1078);
nand U437 (N_437,In_1017,In_641);
nor U438 (N_438,In_502,In_327);
nand U439 (N_439,In_781,In_907);
nand U440 (N_440,In_1310,In_26);
and U441 (N_441,In_721,In_1479);
nand U442 (N_442,In_304,In_1390);
or U443 (N_443,In_822,In_12);
nand U444 (N_444,In_588,In_576);
or U445 (N_445,In_1394,In_751);
nand U446 (N_446,In_642,In_305);
nor U447 (N_447,In_400,In_472);
and U448 (N_448,In_226,In_1274);
or U449 (N_449,In_1414,In_37);
or U450 (N_450,In_728,In_333);
and U451 (N_451,In_451,In_816);
nor U452 (N_452,In_112,In_176);
or U453 (N_453,In_1313,In_901);
nor U454 (N_454,In_652,In_1375);
nand U455 (N_455,In_553,In_620);
nor U456 (N_456,In_58,In_1000);
and U457 (N_457,In_671,In_281);
or U458 (N_458,In_237,In_1194);
or U459 (N_459,In_1103,In_994);
nor U460 (N_460,In_518,In_441);
or U461 (N_461,In_950,In_1114);
nor U462 (N_462,In_1338,In_298);
nor U463 (N_463,In_1214,In_1337);
nand U464 (N_464,In_144,In_899);
and U465 (N_465,In_1498,In_1402);
nor U466 (N_466,In_1333,In_1007);
and U467 (N_467,In_1193,In_379);
nor U468 (N_468,In_678,In_733);
nor U469 (N_469,In_1355,In_840);
nand U470 (N_470,In_1289,In_683);
and U471 (N_471,In_920,In_1262);
nor U472 (N_472,In_1026,In_930);
nor U473 (N_473,In_252,In_960);
nand U474 (N_474,In_1362,In_462);
and U475 (N_475,In_178,In_275);
or U476 (N_476,In_811,In_589);
and U477 (N_477,In_1006,In_609);
and U478 (N_478,In_1266,In_865);
nand U479 (N_479,In_868,In_90);
or U480 (N_480,In_760,In_453);
nand U481 (N_481,In_1163,In_442);
nand U482 (N_482,In_1219,In_933);
nor U483 (N_483,In_839,In_1370);
nor U484 (N_484,In_1045,In_753);
and U485 (N_485,In_1186,In_420);
and U486 (N_486,In_497,In_269);
and U487 (N_487,In_1077,In_1457);
nand U488 (N_488,In_60,In_488);
nor U489 (N_489,In_288,In_1322);
or U490 (N_490,In_871,In_800);
or U491 (N_491,In_1238,In_1376);
and U492 (N_492,In_1245,In_1225);
nor U493 (N_493,In_555,In_6);
or U494 (N_494,In_478,In_1438);
and U495 (N_495,In_900,In_1192);
nor U496 (N_496,In_513,In_172);
nor U497 (N_497,In_986,In_847);
nand U498 (N_498,In_306,In_1383);
or U499 (N_499,In_697,In_191);
nor U500 (N_500,In_1261,In_137);
nand U501 (N_501,In_533,In_328);
and U502 (N_502,In_374,In_247);
nor U503 (N_503,In_581,In_15);
nand U504 (N_504,In_59,In_1473);
nor U505 (N_505,In_1089,In_813);
nand U506 (N_506,In_1447,In_1350);
nor U507 (N_507,In_290,In_1468);
and U508 (N_508,In_1456,In_1260);
nand U509 (N_509,In_688,In_284);
or U510 (N_510,In_1072,In_201);
and U511 (N_511,In_1382,In_1428);
nor U512 (N_512,In_524,In_1251);
nor U513 (N_513,In_731,In_869);
or U514 (N_514,In_1258,In_484);
nand U515 (N_515,In_573,In_227);
nor U516 (N_516,In_399,In_1111);
nand U517 (N_517,In_1436,In_367);
nand U518 (N_518,In_1191,In_954);
or U519 (N_519,In_1252,In_131);
nor U520 (N_520,In_886,In_970);
nand U521 (N_521,In_1323,In_925);
nand U522 (N_522,In_971,In_1094);
nand U523 (N_523,In_213,In_699);
and U524 (N_524,In_980,In_61);
nor U525 (N_525,In_286,In_725);
and U526 (N_526,In_340,In_263);
nand U527 (N_527,In_444,In_1211);
or U528 (N_528,In_1188,In_552);
nor U529 (N_529,In_14,In_749);
or U530 (N_530,In_1171,In_951);
nand U531 (N_531,In_1014,In_495);
and U532 (N_532,In_739,In_846);
or U533 (N_533,In_422,In_424);
or U534 (N_534,In_1147,In_139);
and U535 (N_535,In_1213,In_83);
and U536 (N_536,In_934,In_995);
or U537 (N_537,In_190,In_1233);
or U538 (N_538,In_814,In_1024);
or U539 (N_539,In_887,In_775);
nor U540 (N_540,In_390,In_162);
and U541 (N_541,In_1095,In_1100);
nand U542 (N_542,In_538,In_897);
nand U543 (N_543,In_54,In_1491);
nor U544 (N_544,In_936,In_547);
and U545 (N_545,In_206,In_585);
nor U546 (N_546,In_1229,In_1050);
or U547 (N_547,In_1281,In_409);
nor U548 (N_548,In_958,In_644);
or U549 (N_549,In_1179,In_1146);
and U550 (N_550,In_579,In_1450);
nor U551 (N_551,In_297,In_640);
and U552 (N_552,In_498,In_630);
or U553 (N_553,In_170,In_308);
or U554 (N_554,In_584,In_992);
nand U555 (N_555,In_637,In_85);
xor U556 (N_556,In_197,In_571);
nor U557 (N_557,In_1449,In_151);
nor U558 (N_558,In_841,In_935);
nor U559 (N_559,In_1290,In_1130);
or U560 (N_560,In_350,In_605);
nand U561 (N_561,In_155,In_164);
and U562 (N_562,In_239,In_494);
nand U563 (N_563,In_1372,In_741);
or U564 (N_564,In_622,In_357);
nor U565 (N_565,In_651,In_1038);
nor U566 (N_566,In_617,In_49);
or U567 (N_567,In_891,In_634);
and U568 (N_568,In_1320,In_1080);
or U569 (N_569,In_684,In_1412);
nand U570 (N_570,In_943,In_1405);
nor U571 (N_571,In_1215,In_1429);
and U572 (N_572,In_436,In_653);
or U573 (N_573,In_918,In_1286);
and U574 (N_574,In_1257,In_301);
nor U575 (N_575,In_864,In_602);
nand U576 (N_576,In_1385,In_21);
and U577 (N_577,In_410,In_480);
or U578 (N_578,In_70,In_1164);
or U579 (N_579,In_434,In_952);
and U580 (N_580,In_1477,In_127);
nor U581 (N_581,In_1180,In_1230);
and U582 (N_582,In_267,In_113);
nor U583 (N_583,In_1368,In_1101);
and U584 (N_584,In_457,In_519);
nor U585 (N_585,In_404,In_1425);
nor U586 (N_586,In_1068,In_55);
nand U587 (N_587,In_837,In_1476);
nor U588 (N_588,In_1294,In_1056);
or U589 (N_589,In_408,In_564);
xnor U590 (N_590,In_828,In_1197);
nor U591 (N_591,In_1071,In_1040);
or U592 (N_592,In_1222,In_681);
or U593 (N_593,In_860,In_1034);
and U594 (N_594,In_366,In_786);
or U595 (N_595,In_303,In_505);
or U596 (N_596,In_1012,In_406);
or U597 (N_597,In_913,In_186);
nor U598 (N_598,In_509,In_160);
or U599 (N_599,In_593,In_522);
or U600 (N_600,In_171,In_1352);
nor U601 (N_601,In_1047,In_177);
or U602 (N_602,In_827,In_1296);
and U603 (N_603,In_445,In_663);
nor U604 (N_604,In_1209,In_1028);
and U605 (N_605,In_493,In_1158);
nand U606 (N_606,In_796,In_92);
nand U607 (N_607,In_154,In_332);
or U608 (N_608,In_475,In_696);
or U609 (N_609,In_1437,In_39);
nand U610 (N_610,In_1151,In_657);
nand U611 (N_611,In_74,In_75);
or U612 (N_612,In_1279,In_251);
or U613 (N_613,In_702,In_273);
nor U614 (N_614,In_1184,In_499);
and U615 (N_615,In_985,In_645);
nor U616 (N_616,In_862,In_461);
nor U617 (N_617,In_412,In_962);
nand U618 (N_618,In_216,In_607);
nor U619 (N_619,In_1431,In_854);
and U620 (N_620,In_910,In_19);
or U621 (N_621,In_220,In_67);
nand U622 (N_622,In_1488,In_638);
or U623 (N_623,In_809,In_194);
nor U624 (N_624,In_244,In_1018);
and U625 (N_625,In_560,In_1150);
or U626 (N_626,In_835,In_1142);
and U627 (N_627,In_1384,In_826);
or U628 (N_628,In_601,In_1419);
and U629 (N_629,In_1490,In_455);
nor U630 (N_630,In_662,In_1462);
nand U631 (N_631,In_673,In_370);
or U632 (N_632,In_501,In_701);
and U633 (N_633,In_959,In_896);
nand U634 (N_634,In_1379,In_361);
and U635 (N_635,In_307,In_1299);
nand U636 (N_636,In_1484,In_675);
nand U637 (N_637,In_27,In_258);
xor U638 (N_638,In_134,In_392);
or U639 (N_639,In_707,In_274);
and U640 (N_640,In_1200,In_78);
or U641 (N_641,In_57,In_414);
or U642 (N_642,In_1199,In_143);
nor U643 (N_643,In_1102,In_215);
and U644 (N_644,In_368,In_636);
nor U645 (N_645,In_676,In_158);
or U646 (N_646,In_815,In_42);
nand U647 (N_647,In_541,In_1459);
nor U648 (N_648,In_355,In_1221);
or U649 (N_649,In_1042,In_516);
nor U650 (N_650,In_1424,In_1062);
or U651 (N_651,In_386,In_360);
nand U652 (N_652,In_69,In_266);
nor U653 (N_653,In_1328,In_1433);
nor U654 (N_654,In_1403,In_772);
or U655 (N_655,In_1227,In_851);
or U656 (N_656,In_779,In_356);
nor U657 (N_657,In_24,In_520);
nand U658 (N_658,In_1434,In_888);
or U659 (N_659,In_1374,In_727);
nor U660 (N_660,In_527,In_231);
and U661 (N_661,In_229,In_991);
or U662 (N_662,In_120,In_1378);
and U663 (N_663,In_1124,In_344);
nor U664 (N_664,In_1175,In_1325);
nor U665 (N_665,In_473,In_362);
nand U666 (N_666,In_795,In_1030);
nand U667 (N_667,In_629,In_235);
and U668 (N_668,In_1396,In_212);
nor U669 (N_669,In_722,In_417);
and U670 (N_670,In_280,In_666);
nand U671 (N_671,In_691,In_1220);
and U672 (N_672,In_793,In_219);
nor U673 (N_673,In_1237,In_690);
nand U674 (N_674,In_396,In_583);
nor U675 (N_675,In_426,In_890);
and U676 (N_676,In_168,In_532);
nor U677 (N_677,In_761,In_981);
and U678 (N_678,In_371,In_938);
and U679 (N_679,In_787,In_797);
or U680 (N_680,In_1406,In_766);
or U681 (N_681,In_152,In_423);
nand U682 (N_682,In_877,In_1120);
nor U683 (N_683,In_1311,In_271);
nor U684 (N_684,In_240,In_3);
nor U685 (N_685,In_649,In_904);
or U686 (N_686,In_563,In_117);
or U687 (N_687,In_1052,In_1348);
or U688 (N_688,In_1136,In_807);
or U689 (N_689,In_165,In_737);
or U690 (N_690,In_7,In_817);
nand U691 (N_691,In_93,In_124);
and U692 (N_692,In_1115,In_1060);
nand U693 (N_693,In_503,In_63);
nor U694 (N_694,In_726,In_983);
or U695 (N_695,In_296,In_102);
or U696 (N_696,In_895,In_1202);
and U697 (N_697,In_1410,In_32);
nand U698 (N_698,In_1435,In_1149);
nand U699 (N_699,In_1391,In_230);
or U700 (N_700,In_1421,In_546);
nor U701 (N_701,In_245,In_791);
nand U702 (N_702,In_180,In_1176);
nor U703 (N_703,In_1441,In_755);
or U704 (N_704,In_1380,In_1283);
or U705 (N_705,In_218,In_1354);
nand U706 (N_706,In_1168,In_72);
and U707 (N_707,In_310,In_723);
and U708 (N_708,In_401,In_545);
or U709 (N_709,In_48,In_1495);
nor U710 (N_710,In_1129,In_167);
and U711 (N_711,In_1064,In_302);
and U712 (N_712,In_1067,In_224);
nand U713 (N_713,In_383,In_84);
or U714 (N_714,In_825,In_774);
or U715 (N_715,In_788,In_385);
nor U716 (N_716,In_889,In_458);
nand U717 (N_717,In_989,In_89);
nand U718 (N_718,In_750,In_1058);
nand U719 (N_719,In_1159,In_4);
or U720 (N_720,In_380,In_1303);
xnor U721 (N_721,In_806,In_577);
nand U722 (N_722,In_182,In_166);
and U723 (N_723,In_1097,In_111);
nor U724 (N_724,In_1032,In_1268);
or U725 (N_725,In_876,In_765);
and U726 (N_726,In_1367,In_1365);
or U727 (N_727,In_857,In_799);
nor U728 (N_728,In_1317,In_1216);
and U729 (N_729,In_413,In_776);
and U730 (N_730,In_1069,In_1277);
and U731 (N_731,In_262,In_998);
nor U732 (N_732,In_1349,In_1029);
or U733 (N_733,In_911,In_711);
or U734 (N_734,In_1297,In_483);
nand U735 (N_735,In_272,In_477);
nor U736 (N_736,In_384,In_469);
and U737 (N_737,In_1288,In_626);
or U738 (N_738,In_639,In_762);
nor U739 (N_739,In_566,In_1451);
and U740 (N_740,In_437,In_1181);
and U741 (N_741,In_510,In_1301);
nor U742 (N_742,In_717,In_915);
and U743 (N_743,In_586,In_1172);
and U744 (N_744,In_1174,In_1141);
or U745 (N_745,In_259,In_993);
or U746 (N_746,In_668,In_1358);
nand U747 (N_747,In_10,In_184);
nand U748 (N_748,In_1059,In_193);
or U749 (N_749,In_592,In_625);
and U750 (N_750,In_291,In_567);
nor U751 (N_751,In_601,In_1294);
or U752 (N_752,In_135,In_1005);
nor U753 (N_753,In_1077,In_1365);
nand U754 (N_754,In_597,In_677);
nand U755 (N_755,In_798,In_845);
nand U756 (N_756,In_805,In_1205);
and U757 (N_757,In_904,In_873);
nor U758 (N_758,In_490,In_784);
and U759 (N_759,In_771,In_389);
nor U760 (N_760,In_798,In_758);
nand U761 (N_761,In_1137,In_996);
nor U762 (N_762,In_1126,In_17);
and U763 (N_763,In_92,In_1098);
or U764 (N_764,In_286,In_185);
and U765 (N_765,In_1353,In_367);
nand U766 (N_766,In_1062,In_222);
nand U767 (N_767,In_1403,In_467);
nor U768 (N_768,In_1190,In_59);
nand U769 (N_769,In_142,In_362);
nor U770 (N_770,In_629,In_339);
nor U771 (N_771,In_1116,In_1323);
and U772 (N_772,In_400,In_624);
or U773 (N_773,In_568,In_593);
or U774 (N_774,In_88,In_76);
and U775 (N_775,In_812,In_77);
nand U776 (N_776,In_1371,In_1480);
or U777 (N_777,In_731,In_17);
nand U778 (N_778,In_858,In_792);
or U779 (N_779,In_1158,In_863);
or U780 (N_780,In_1397,In_320);
nor U781 (N_781,In_313,In_50);
nand U782 (N_782,In_1334,In_1489);
nor U783 (N_783,In_1065,In_771);
or U784 (N_784,In_492,In_529);
nor U785 (N_785,In_1427,In_130);
nor U786 (N_786,In_1225,In_940);
nor U787 (N_787,In_838,In_321);
nor U788 (N_788,In_1413,In_1156);
nor U789 (N_789,In_278,In_1226);
or U790 (N_790,In_53,In_911);
and U791 (N_791,In_654,In_587);
and U792 (N_792,In_348,In_289);
nand U793 (N_793,In_994,In_590);
nor U794 (N_794,In_1184,In_604);
nand U795 (N_795,In_221,In_999);
and U796 (N_796,In_811,In_781);
and U797 (N_797,In_794,In_7);
nand U798 (N_798,In_1181,In_1469);
nand U799 (N_799,In_377,In_140);
or U800 (N_800,In_364,In_807);
nor U801 (N_801,In_240,In_641);
and U802 (N_802,In_467,In_382);
or U803 (N_803,In_795,In_1303);
and U804 (N_804,In_259,In_49);
and U805 (N_805,In_233,In_1314);
nand U806 (N_806,In_1237,In_1084);
and U807 (N_807,In_582,In_931);
or U808 (N_808,In_579,In_218);
nand U809 (N_809,In_2,In_902);
or U810 (N_810,In_411,In_1158);
or U811 (N_811,In_325,In_69);
nor U812 (N_812,In_271,In_230);
or U813 (N_813,In_1379,In_442);
nor U814 (N_814,In_291,In_1261);
nand U815 (N_815,In_913,In_1267);
nor U816 (N_816,In_1023,In_106);
or U817 (N_817,In_824,In_172);
nand U818 (N_818,In_821,In_535);
or U819 (N_819,In_37,In_1157);
and U820 (N_820,In_1260,In_415);
nand U821 (N_821,In_873,In_1342);
nor U822 (N_822,In_246,In_697);
and U823 (N_823,In_1042,In_1291);
nand U824 (N_824,In_349,In_779);
nor U825 (N_825,In_120,In_411);
nor U826 (N_826,In_1100,In_202);
nand U827 (N_827,In_673,In_1269);
xor U828 (N_828,In_1321,In_256);
nor U829 (N_829,In_1229,In_1059);
and U830 (N_830,In_1393,In_923);
nand U831 (N_831,In_622,In_621);
nand U832 (N_832,In_1313,In_766);
nand U833 (N_833,In_362,In_1035);
or U834 (N_834,In_803,In_1107);
nor U835 (N_835,In_524,In_1482);
and U836 (N_836,In_114,In_134);
or U837 (N_837,In_200,In_237);
nor U838 (N_838,In_910,In_271);
and U839 (N_839,In_348,In_1432);
or U840 (N_840,In_824,In_1243);
and U841 (N_841,In_407,In_573);
nand U842 (N_842,In_782,In_776);
nor U843 (N_843,In_489,In_1203);
xnor U844 (N_844,In_200,In_1454);
nand U845 (N_845,In_931,In_490);
nor U846 (N_846,In_958,In_290);
and U847 (N_847,In_1137,In_1251);
or U848 (N_848,In_1425,In_1370);
nand U849 (N_849,In_379,In_103);
nor U850 (N_850,In_512,In_1447);
nor U851 (N_851,In_953,In_734);
nor U852 (N_852,In_1343,In_895);
nand U853 (N_853,In_295,In_1130);
nor U854 (N_854,In_1409,In_792);
and U855 (N_855,In_927,In_646);
or U856 (N_856,In_1209,In_161);
or U857 (N_857,In_1012,In_547);
nor U858 (N_858,In_141,In_815);
nand U859 (N_859,In_1184,In_449);
or U860 (N_860,In_1086,In_310);
nand U861 (N_861,In_1381,In_1382);
or U862 (N_862,In_411,In_673);
or U863 (N_863,In_923,In_138);
nor U864 (N_864,In_506,In_951);
or U865 (N_865,In_1,In_568);
or U866 (N_866,In_1374,In_226);
and U867 (N_867,In_263,In_655);
nand U868 (N_868,In_22,In_785);
nand U869 (N_869,In_352,In_111);
and U870 (N_870,In_840,In_25);
or U871 (N_871,In_428,In_609);
xnor U872 (N_872,In_1333,In_468);
nand U873 (N_873,In_229,In_476);
nand U874 (N_874,In_47,In_384);
nor U875 (N_875,In_1458,In_681);
or U876 (N_876,In_588,In_124);
and U877 (N_877,In_747,In_689);
or U878 (N_878,In_863,In_778);
or U879 (N_879,In_360,In_1005);
and U880 (N_880,In_462,In_1239);
or U881 (N_881,In_1435,In_277);
nor U882 (N_882,In_819,In_1045);
nand U883 (N_883,In_743,In_623);
nand U884 (N_884,In_1064,In_212);
and U885 (N_885,In_803,In_714);
or U886 (N_886,In_806,In_853);
and U887 (N_887,In_876,In_1235);
nand U888 (N_888,In_1272,In_1498);
and U889 (N_889,In_93,In_322);
nor U890 (N_890,In_695,In_1005);
and U891 (N_891,In_1366,In_1320);
and U892 (N_892,In_300,In_669);
and U893 (N_893,In_505,In_337);
or U894 (N_894,In_1399,In_887);
nor U895 (N_895,In_1123,In_935);
or U896 (N_896,In_416,In_312);
nor U897 (N_897,In_371,In_467);
nor U898 (N_898,In_1313,In_1416);
nor U899 (N_899,In_364,In_442);
nor U900 (N_900,In_255,In_702);
nand U901 (N_901,In_968,In_240);
or U902 (N_902,In_1438,In_1198);
or U903 (N_903,In_71,In_985);
and U904 (N_904,In_1337,In_99);
nor U905 (N_905,In_1371,In_303);
or U906 (N_906,In_1134,In_167);
nand U907 (N_907,In_54,In_426);
or U908 (N_908,In_874,In_334);
nand U909 (N_909,In_822,In_568);
nor U910 (N_910,In_902,In_1003);
and U911 (N_911,In_784,In_1398);
or U912 (N_912,In_1118,In_500);
or U913 (N_913,In_991,In_89);
nand U914 (N_914,In_538,In_969);
nand U915 (N_915,In_364,In_1387);
nor U916 (N_916,In_431,In_697);
nor U917 (N_917,In_661,In_56);
or U918 (N_918,In_85,In_1052);
or U919 (N_919,In_246,In_980);
nand U920 (N_920,In_1451,In_200);
or U921 (N_921,In_410,In_858);
nand U922 (N_922,In_640,In_1091);
nor U923 (N_923,In_1126,In_1078);
or U924 (N_924,In_129,In_204);
or U925 (N_925,In_591,In_1257);
and U926 (N_926,In_422,In_1472);
or U927 (N_927,In_842,In_223);
nand U928 (N_928,In_411,In_663);
and U929 (N_929,In_896,In_678);
or U930 (N_930,In_1133,In_1315);
nor U931 (N_931,In_1234,In_16);
and U932 (N_932,In_710,In_1084);
nand U933 (N_933,In_471,In_994);
nor U934 (N_934,In_923,In_1465);
nor U935 (N_935,In_180,In_782);
nor U936 (N_936,In_960,In_921);
nand U937 (N_937,In_1113,In_901);
and U938 (N_938,In_695,In_2);
or U939 (N_939,In_1186,In_284);
nor U940 (N_940,In_725,In_858);
or U941 (N_941,In_1478,In_1433);
or U942 (N_942,In_284,In_224);
or U943 (N_943,In_292,In_1303);
nor U944 (N_944,In_534,In_518);
nand U945 (N_945,In_1229,In_214);
nand U946 (N_946,In_363,In_462);
or U947 (N_947,In_1106,In_453);
nand U948 (N_948,In_821,In_1131);
or U949 (N_949,In_45,In_111);
and U950 (N_950,In_430,In_587);
nand U951 (N_951,In_1271,In_1178);
and U952 (N_952,In_688,In_205);
and U953 (N_953,In_1283,In_1346);
and U954 (N_954,In_1101,In_717);
nor U955 (N_955,In_498,In_898);
nand U956 (N_956,In_394,In_1487);
nand U957 (N_957,In_86,In_239);
or U958 (N_958,In_637,In_846);
and U959 (N_959,In_674,In_367);
or U960 (N_960,In_918,In_309);
and U961 (N_961,In_1258,In_185);
or U962 (N_962,In_873,In_1334);
nor U963 (N_963,In_503,In_292);
nor U964 (N_964,In_5,In_257);
nand U965 (N_965,In_781,In_1364);
nand U966 (N_966,In_153,In_1232);
nor U967 (N_967,In_1104,In_1266);
or U968 (N_968,In_1188,In_1418);
or U969 (N_969,In_607,In_818);
nor U970 (N_970,In_873,In_888);
nand U971 (N_971,In_135,In_1475);
or U972 (N_972,In_65,In_1358);
or U973 (N_973,In_1127,In_726);
nand U974 (N_974,In_609,In_497);
and U975 (N_975,In_1157,In_671);
or U976 (N_976,In_232,In_1443);
or U977 (N_977,In_797,In_415);
and U978 (N_978,In_313,In_121);
nand U979 (N_979,In_89,In_409);
or U980 (N_980,In_674,In_1400);
nor U981 (N_981,In_574,In_144);
nor U982 (N_982,In_512,In_34);
nor U983 (N_983,In_962,In_1265);
or U984 (N_984,In_865,In_1496);
and U985 (N_985,In_869,In_1122);
and U986 (N_986,In_783,In_925);
nand U987 (N_987,In_1143,In_1320);
or U988 (N_988,In_855,In_1168);
nand U989 (N_989,In_581,In_1228);
or U990 (N_990,In_474,In_1469);
or U991 (N_991,In_982,In_1467);
nor U992 (N_992,In_657,In_659);
and U993 (N_993,In_257,In_1359);
nor U994 (N_994,In_610,In_1197);
or U995 (N_995,In_1329,In_7);
nand U996 (N_996,In_1036,In_60);
nor U997 (N_997,In_1215,In_464);
nand U998 (N_998,In_1450,In_344);
nor U999 (N_999,In_23,In_1248);
or U1000 (N_1000,In_927,In_518);
or U1001 (N_1001,In_507,In_376);
nand U1002 (N_1002,In_583,In_78);
and U1003 (N_1003,In_349,In_1028);
nor U1004 (N_1004,In_864,In_701);
nor U1005 (N_1005,In_906,In_1166);
nor U1006 (N_1006,In_1041,In_19);
nand U1007 (N_1007,In_1340,In_516);
nor U1008 (N_1008,In_344,In_886);
or U1009 (N_1009,In_570,In_1253);
or U1010 (N_1010,In_1172,In_1448);
or U1011 (N_1011,In_294,In_49);
or U1012 (N_1012,In_160,In_833);
and U1013 (N_1013,In_1450,In_1007);
nand U1014 (N_1014,In_16,In_981);
nand U1015 (N_1015,In_463,In_214);
or U1016 (N_1016,In_1432,In_500);
and U1017 (N_1017,In_115,In_1367);
nor U1018 (N_1018,In_1467,In_757);
or U1019 (N_1019,In_1127,In_679);
and U1020 (N_1020,In_945,In_104);
nand U1021 (N_1021,In_671,In_228);
and U1022 (N_1022,In_1004,In_537);
nand U1023 (N_1023,In_71,In_61);
nand U1024 (N_1024,In_1499,In_238);
nor U1025 (N_1025,In_787,In_1169);
nand U1026 (N_1026,In_1110,In_1224);
or U1027 (N_1027,In_33,In_64);
nand U1028 (N_1028,In_150,In_1443);
nor U1029 (N_1029,In_1343,In_1121);
or U1030 (N_1030,In_356,In_337);
nand U1031 (N_1031,In_1094,In_229);
nand U1032 (N_1032,In_583,In_491);
nor U1033 (N_1033,In_1293,In_79);
nand U1034 (N_1034,In_289,In_379);
nor U1035 (N_1035,In_1465,In_504);
and U1036 (N_1036,In_904,In_894);
nand U1037 (N_1037,In_1069,In_931);
nand U1038 (N_1038,In_541,In_25);
and U1039 (N_1039,In_1226,In_916);
nand U1040 (N_1040,In_1104,In_1248);
and U1041 (N_1041,In_1074,In_1249);
nor U1042 (N_1042,In_750,In_763);
nand U1043 (N_1043,In_1152,In_905);
or U1044 (N_1044,In_394,In_1056);
and U1045 (N_1045,In_871,In_532);
and U1046 (N_1046,In_1185,In_548);
nor U1047 (N_1047,In_753,In_489);
and U1048 (N_1048,In_432,In_754);
nand U1049 (N_1049,In_882,In_769);
and U1050 (N_1050,In_207,In_990);
or U1051 (N_1051,In_1244,In_797);
and U1052 (N_1052,In_1109,In_1119);
or U1053 (N_1053,In_1192,In_1030);
or U1054 (N_1054,In_130,In_27);
and U1055 (N_1055,In_1462,In_1373);
nor U1056 (N_1056,In_1033,In_1384);
nor U1057 (N_1057,In_519,In_16);
nand U1058 (N_1058,In_721,In_1396);
or U1059 (N_1059,In_954,In_58);
nand U1060 (N_1060,In_878,In_222);
nand U1061 (N_1061,In_305,In_1363);
nand U1062 (N_1062,In_347,In_352);
nor U1063 (N_1063,In_1422,In_576);
or U1064 (N_1064,In_794,In_630);
nand U1065 (N_1065,In_385,In_935);
nor U1066 (N_1066,In_770,In_1410);
nor U1067 (N_1067,In_234,In_698);
or U1068 (N_1068,In_446,In_1244);
and U1069 (N_1069,In_654,In_47);
or U1070 (N_1070,In_804,In_47);
or U1071 (N_1071,In_81,In_66);
nand U1072 (N_1072,In_1411,In_735);
and U1073 (N_1073,In_476,In_1444);
nand U1074 (N_1074,In_254,In_1278);
or U1075 (N_1075,In_1242,In_792);
nand U1076 (N_1076,In_541,In_1105);
or U1077 (N_1077,In_1131,In_1120);
nor U1078 (N_1078,In_274,In_62);
or U1079 (N_1079,In_60,In_432);
nand U1080 (N_1080,In_510,In_743);
nor U1081 (N_1081,In_625,In_60);
and U1082 (N_1082,In_289,In_802);
or U1083 (N_1083,In_1046,In_611);
nor U1084 (N_1084,In_523,In_278);
nor U1085 (N_1085,In_295,In_490);
nor U1086 (N_1086,In_815,In_1194);
and U1087 (N_1087,In_337,In_456);
or U1088 (N_1088,In_1434,In_1433);
or U1089 (N_1089,In_187,In_997);
nand U1090 (N_1090,In_737,In_329);
nand U1091 (N_1091,In_368,In_53);
nand U1092 (N_1092,In_430,In_507);
and U1093 (N_1093,In_1318,In_504);
and U1094 (N_1094,In_655,In_637);
nand U1095 (N_1095,In_85,In_651);
and U1096 (N_1096,In_643,In_931);
nand U1097 (N_1097,In_404,In_1376);
and U1098 (N_1098,In_729,In_1258);
xor U1099 (N_1099,In_1064,In_664);
nand U1100 (N_1100,In_248,In_43);
or U1101 (N_1101,In_1301,In_305);
and U1102 (N_1102,In_897,In_281);
or U1103 (N_1103,In_963,In_1153);
and U1104 (N_1104,In_243,In_1337);
nand U1105 (N_1105,In_180,In_1291);
nand U1106 (N_1106,In_414,In_764);
and U1107 (N_1107,In_1333,In_1492);
and U1108 (N_1108,In_243,In_868);
nor U1109 (N_1109,In_1364,In_72);
or U1110 (N_1110,In_756,In_1344);
or U1111 (N_1111,In_1264,In_504);
and U1112 (N_1112,In_923,In_137);
or U1113 (N_1113,In_35,In_555);
nor U1114 (N_1114,In_863,In_40);
nor U1115 (N_1115,In_498,In_18);
and U1116 (N_1116,In_223,In_1004);
nor U1117 (N_1117,In_447,In_504);
nor U1118 (N_1118,In_9,In_535);
or U1119 (N_1119,In_454,In_684);
nor U1120 (N_1120,In_590,In_394);
and U1121 (N_1121,In_1307,In_1089);
and U1122 (N_1122,In_535,In_217);
or U1123 (N_1123,In_1099,In_1143);
nand U1124 (N_1124,In_1313,In_158);
nand U1125 (N_1125,In_612,In_240);
and U1126 (N_1126,In_1466,In_956);
nand U1127 (N_1127,In_1079,In_806);
and U1128 (N_1128,In_726,In_1483);
or U1129 (N_1129,In_1454,In_1329);
and U1130 (N_1130,In_288,In_544);
or U1131 (N_1131,In_839,In_234);
nand U1132 (N_1132,In_719,In_661);
nand U1133 (N_1133,In_1183,In_807);
nor U1134 (N_1134,In_776,In_829);
and U1135 (N_1135,In_890,In_611);
and U1136 (N_1136,In_753,In_806);
and U1137 (N_1137,In_1229,In_400);
nor U1138 (N_1138,In_1460,In_726);
nand U1139 (N_1139,In_937,In_1241);
nor U1140 (N_1140,In_360,In_779);
nand U1141 (N_1141,In_443,In_52);
and U1142 (N_1142,In_1445,In_567);
or U1143 (N_1143,In_59,In_1189);
nor U1144 (N_1144,In_1248,In_129);
nand U1145 (N_1145,In_450,In_276);
nor U1146 (N_1146,In_425,In_669);
nor U1147 (N_1147,In_1444,In_173);
nor U1148 (N_1148,In_84,In_313);
or U1149 (N_1149,In_1160,In_332);
nor U1150 (N_1150,In_707,In_1075);
or U1151 (N_1151,In_51,In_287);
nor U1152 (N_1152,In_1488,In_481);
nor U1153 (N_1153,In_1,In_591);
or U1154 (N_1154,In_612,In_1158);
nand U1155 (N_1155,In_263,In_685);
nor U1156 (N_1156,In_1116,In_1425);
and U1157 (N_1157,In_214,In_499);
nand U1158 (N_1158,In_1043,In_1342);
nor U1159 (N_1159,In_351,In_521);
nor U1160 (N_1160,In_1324,In_642);
nand U1161 (N_1161,In_873,In_1036);
or U1162 (N_1162,In_972,In_1105);
or U1163 (N_1163,In_423,In_827);
nand U1164 (N_1164,In_1058,In_916);
and U1165 (N_1165,In_967,In_1448);
and U1166 (N_1166,In_1368,In_508);
or U1167 (N_1167,In_1033,In_748);
nor U1168 (N_1168,In_1021,In_590);
or U1169 (N_1169,In_533,In_1310);
and U1170 (N_1170,In_895,In_453);
nand U1171 (N_1171,In_449,In_1257);
or U1172 (N_1172,In_820,In_571);
or U1173 (N_1173,In_534,In_1292);
or U1174 (N_1174,In_69,In_574);
nand U1175 (N_1175,In_1494,In_856);
nor U1176 (N_1176,In_75,In_1205);
nor U1177 (N_1177,In_443,In_336);
and U1178 (N_1178,In_261,In_1459);
or U1179 (N_1179,In_1453,In_1273);
and U1180 (N_1180,In_108,In_712);
nor U1181 (N_1181,In_833,In_1460);
and U1182 (N_1182,In_1209,In_768);
and U1183 (N_1183,In_1332,In_440);
nand U1184 (N_1184,In_748,In_1211);
nor U1185 (N_1185,In_1083,In_12);
nand U1186 (N_1186,In_75,In_979);
nand U1187 (N_1187,In_1091,In_1335);
and U1188 (N_1188,In_251,In_634);
or U1189 (N_1189,In_400,In_825);
xor U1190 (N_1190,In_816,In_865);
and U1191 (N_1191,In_208,In_672);
or U1192 (N_1192,In_1423,In_364);
and U1193 (N_1193,In_760,In_1204);
nor U1194 (N_1194,In_962,In_98);
or U1195 (N_1195,In_841,In_1490);
nor U1196 (N_1196,In_826,In_1243);
nand U1197 (N_1197,In_1483,In_945);
and U1198 (N_1198,In_1087,In_882);
nor U1199 (N_1199,In_452,In_700);
and U1200 (N_1200,In_1159,In_1428);
and U1201 (N_1201,In_291,In_124);
nand U1202 (N_1202,In_987,In_407);
and U1203 (N_1203,In_125,In_541);
or U1204 (N_1204,In_430,In_746);
nand U1205 (N_1205,In_1452,In_1203);
nor U1206 (N_1206,In_154,In_934);
nand U1207 (N_1207,In_1109,In_1444);
or U1208 (N_1208,In_476,In_95);
nor U1209 (N_1209,In_390,In_93);
or U1210 (N_1210,In_1365,In_774);
or U1211 (N_1211,In_911,In_537);
nand U1212 (N_1212,In_87,In_148);
nand U1213 (N_1213,In_1178,In_874);
nand U1214 (N_1214,In_1302,In_1383);
nor U1215 (N_1215,In_103,In_51);
and U1216 (N_1216,In_841,In_1278);
nor U1217 (N_1217,In_15,In_268);
or U1218 (N_1218,In_1019,In_1148);
nor U1219 (N_1219,In_1487,In_609);
and U1220 (N_1220,In_835,In_329);
or U1221 (N_1221,In_480,In_727);
nand U1222 (N_1222,In_1325,In_1150);
or U1223 (N_1223,In_1258,In_1004);
and U1224 (N_1224,In_1486,In_1369);
nor U1225 (N_1225,In_965,In_298);
or U1226 (N_1226,In_395,In_21);
or U1227 (N_1227,In_842,In_133);
nand U1228 (N_1228,In_1128,In_153);
and U1229 (N_1229,In_579,In_296);
nor U1230 (N_1230,In_501,In_1494);
nor U1231 (N_1231,In_1331,In_1428);
or U1232 (N_1232,In_1318,In_1487);
and U1233 (N_1233,In_874,In_259);
nand U1234 (N_1234,In_346,In_1452);
xor U1235 (N_1235,In_804,In_445);
nand U1236 (N_1236,In_1337,In_678);
nor U1237 (N_1237,In_1300,In_1202);
or U1238 (N_1238,In_1227,In_406);
nand U1239 (N_1239,In_90,In_733);
or U1240 (N_1240,In_1012,In_629);
or U1241 (N_1241,In_822,In_856);
nand U1242 (N_1242,In_348,In_427);
nor U1243 (N_1243,In_1280,In_695);
or U1244 (N_1244,In_1388,In_992);
nor U1245 (N_1245,In_179,In_848);
or U1246 (N_1246,In_728,In_498);
nand U1247 (N_1247,In_1007,In_291);
nand U1248 (N_1248,In_1354,In_965);
or U1249 (N_1249,In_627,In_750);
nand U1250 (N_1250,In_1347,In_1351);
nor U1251 (N_1251,In_1372,In_896);
or U1252 (N_1252,In_1015,In_930);
nand U1253 (N_1253,In_1170,In_428);
nand U1254 (N_1254,In_1127,In_208);
nor U1255 (N_1255,In_999,In_700);
and U1256 (N_1256,In_1463,In_869);
or U1257 (N_1257,In_1452,In_551);
nand U1258 (N_1258,In_1277,In_57);
nand U1259 (N_1259,In_1259,In_477);
or U1260 (N_1260,In_999,In_26);
nor U1261 (N_1261,In_205,In_93);
nor U1262 (N_1262,In_862,In_882);
and U1263 (N_1263,In_1194,In_205);
or U1264 (N_1264,In_1413,In_1485);
nand U1265 (N_1265,In_220,In_1368);
nor U1266 (N_1266,In_1429,In_1075);
nor U1267 (N_1267,In_322,In_516);
nand U1268 (N_1268,In_547,In_324);
or U1269 (N_1269,In_836,In_199);
nand U1270 (N_1270,In_302,In_962);
or U1271 (N_1271,In_1003,In_476);
nand U1272 (N_1272,In_1388,In_320);
nand U1273 (N_1273,In_179,In_212);
nor U1274 (N_1274,In_155,In_668);
nor U1275 (N_1275,In_820,In_367);
and U1276 (N_1276,In_968,In_541);
nand U1277 (N_1277,In_723,In_386);
nand U1278 (N_1278,In_818,In_523);
nor U1279 (N_1279,In_948,In_837);
nand U1280 (N_1280,In_902,In_1111);
nand U1281 (N_1281,In_1271,In_51);
nor U1282 (N_1282,In_495,In_1029);
or U1283 (N_1283,In_686,In_773);
or U1284 (N_1284,In_331,In_1078);
and U1285 (N_1285,In_1397,In_1108);
and U1286 (N_1286,In_127,In_772);
and U1287 (N_1287,In_229,In_220);
nand U1288 (N_1288,In_865,In_744);
nand U1289 (N_1289,In_894,In_479);
or U1290 (N_1290,In_1068,In_750);
and U1291 (N_1291,In_1439,In_237);
nor U1292 (N_1292,In_823,In_1456);
nand U1293 (N_1293,In_776,In_871);
nand U1294 (N_1294,In_253,In_685);
nor U1295 (N_1295,In_376,In_216);
or U1296 (N_1296,In_1282,In_472);
nor U1297 (N_1297,In_699,In_177);
nand U1298 (N_1298,In_944,In_132);
nand U1299 (N_1299,In_716,In_425);
and U1300 (N_1300,In_304,In_175);
and U1301 (N_1301,In_385,In_644);
or U1302 (N_1302,In_118,In_877);
and U1303 (N_1303,In_181,In_1064);
nand U1304 (N_1304,In_704,In_923);
nand U1305 (N_1305,In_515,In_686);
or U1306 (N_1306,In_608,In_320);
or U1307 (N_1307,In_994,In_1072);
and U1308 (N_1308,In_903,In_1025);
or U1309 (N_1309,In_136,In_1391);
or U1310 (N_1310,In_703,In_489);
nor U1311 (N_1311,In_836,In_1008);
nor U1312 (N_1312,In_1324,In_701);
nand U1313 (N_1313,In_111,In_467);
or U1314 (N_1314,In_185,In_363);
and U1315 (N_1315,In_1006,In_799);
nor U1316 (N_1316,In_987,In_890);
or U1317 (N_1317,In_30,In_670);
nand U1318 (N_1318,In_1402,In_112);
nand U1319 (N_1319,In_1082,In_1438);
nand U1320 (N_1320,In_451,In_158);
xor U1321 (N_1321,In_1398,In_1210);
or U1322 (N_1322,In_636,In_551);
and U1323 (N_1323,In_794,In_1434);
and U1324 (N_1324,In_29,In_1102);
or U1325 (N_1325,In_249,In_775);
and U1326 (N_1326,In_30,In_951);
or U1327 (N_1327,In_1300,In_330);
or U1328 (N_1328,In_812,In_540);
nor U1329 (N_1329,In_653,In_421);
nor U1330 (N_1330,In_157,In_408);
and U1331 (N_1331,In_1088,In_931);
nor U1332 (N_1332,In_95,In_753);
or U1333 (N_1333,In_169,In_674);
xor U1334 (N_1334,In_51,In_1241);
and U1335 (N_1335,In_595,In_1288);
nand U1336 (N_1336,In_1377,In_14);
or U1337 (N_1337,In_1236,In_1369);
nor U1338 (N_1338,In_327,In_1143);
and U1339 (N_1339,In_1022,In_819);
nor U1340 (N_1340,In_1497,In_384);
or U1341 (N_1341,In_183,In_1436);
or U1342 (N_1342,In_987,In_420);
nand U1343 (N_1343,In_548,In_362);
and U1344 (N_1344,In_160,In_890);
or U1345 (N_1345,In_649,In_37);
and U1346 (N_1346,In_728,In_169);
nor U1347 (N_1347,In_1183,In_1008);
nor U1348 (N_1348,In_893,In_1030);
or U1349 (N_1349,In_951,In_864);
and U1350 (N_1350,In_49,In_1340);
nor U1351 (N_1351,In_741,In_1169);
and U1352 (N_1352,In_198,In_1452);
and U1353 (N_1353,In_906,In_903);
or U1354 (N_1354,In_392,In_163);
nor U1355 (N_1355,In_456,In_70);
or U1356 (N_1356,In_682,In_340);
nand U1357 (N_1357,In_1364,In_463);
nand U1358 (N_1358,In_499,In_16);
nor U1359 (N_1359,In_1324,In_1369);
nor U1360 (N_1360,In_1009,In_1442);
nand U1361 (N_1361,In_1197,In_1391);
or U1362 (N_1362,In_82,In_539);
nor U1363 (N_1363,In_762,In_1215);
and U1364 (N_1364,In_870,In_1008);
nand U1365 (N_1365,In_1210,In_1255);
or U1366 (N_1366,In_742,In_718);
nand U1367 (N_1367,In_1469,In_539);
nand U1368 (N_1368,In_678,In_137);
nand U1369 (N_1369,In_304,In_1228);
or U1370 (N_1370,In_1369,In_851);
or U1371 (N_1371,In_682,In_1355);
and U1372 (N_1372,In_346,In_352);
nor U1373 (N_1373,In_426,In_798);
and U1374 (N_1374,In_432,In_982);
nand U1375 (N_1375,In_415,In_1078);
nor U1376 (N_1376,In_111,In_30);
nor U1377 (N_1377,In_1285,In_813);
nand U1378 (N_1378,In_1414,In_250);
nand U1379 (N_1379,In_33,In_1322);
nand U1380 (N_1380,In_38,In_697);
nand U1381 (N_1381,In_934,In_1076);
nor U1382 (N_1382,In_239,In_101);
and U1383 (N_1383,In_1039,In_188);
and U1384 (N_1384,In_237,In_627);
and U1385 (N_1385,In_422,In_664);
nand U1386 (N_1386,In_459,In_877);
or U1387 (N_1387,In_1349,In_4);
and U1388 (N_1388,In_832,In_607);
and U1389 (N_1389,In_1157,In_784);
and U1390 (N_1390,In_985,In_827);
and U1391 (N_1391,In_1472,In_1295);
nor U1392 (N_1392,In_1491,In_1060);
nand U1393 (N_1393,In_78,In_104);
nor U1394 (N_1394,In_941,In_873);
nand U1395 (N_1395,In_31,In_852);
or U1396 (N_1396,In_988,In_804);
nand U1397 (N_1397,In_14,In_219);
or U1398 (N_1398,In_1333,In_908);
or U1399 (N_1399,In_513,In_1098);
nor U1400 (N_1400,In_62,In_370);
nand U1401 (N_1401,In_1316,In_88);
nand U1402 (N_1402,In_1350,In_878);
nor U1403 (N_1403,In_621,In_967);
nand U1404 (N_1404,In_732,In_1056);
nand U1405 (N_1405,In_1429,In_254);
nor U1406 (N_1406,In_211,In_1135);
and U1407 (N_1407,In_492,In_1251);
nor U1408 (N_1408,In_1002,In_127);
nor U1409 (N_1409,In_1190,In_650);
nand U1410 (N_1410,In_38,In_62);
nor U1411 (N_1411,In_812,In_1135);
or U1412 (N_1412,In_1140,In_1086);
or U1413 (N_1413,In_458,In_1171);
nand U1414 (N_1414,In_674,In_1140);
or U1415 (N_1415,In_428,In_1355);
and U1416 (N_1416,In_730,In_784);
nand U1417 (N_1417,In_188,In_632);
nand U1418 (N_1418,In_1201,In_130);
nor U1419 (N_1419,In_1323,In_1348);
nor U1420 (N_1420,In_56,In_335);
or U1421 (N_1421,In_1423,In_189);
nor U1422 (N_1422,In_163,In_487);
nor U1423 (N_1423,In_759,In_46);
nor U1424 (N_1424,In_1284,In_689);
nor U1425 (N_1425,In_498,In_745);
nand U1426 (N_1426,In_350,In_227);
and U1427 (N_1427,In_582,In_1192);
and U1428 (N_1428,In_117,In_1001);
nand U1429 (N_1429,In_1150,In_759);
and U1430 (N_1430,In_133,In_1185);
or U1431 (N_1431,In_906,In_497);
nand U1432 (N_1432,In_1368,In_1471);
or U1433 (N_1433,In_1047,In_414);
nand U1434 (N_1434,In_1286,In_307);
and U1435 (N_1435,In_836,In_1391);
nand U1436 (N_1436,In_782,In_1129);
and U1437 (N_1437,In_1253,In_50);
xnor U1438 (N_1438,In_581,In_1154);
and U1439 (N_1439,In_559,In_657);
nand U1440 (N_1440,In_373,In_5);
or U1441 (N_1441,In_126,In_695);
and U1442 (N_1442,In_204,In_104);
nand U1443 (N_1443,In_488,In_838);
nand U1444 (N_1444,In_1372,In_643);
nand U1445 (N_1445,In_1434,In_466);
or U1446 (N_1446,In_244,In_195);
nand U1447 (N_1447,In_227,In_1367);
nor U1448 (N_1448,In_689,In_1147);
and U1449 (N_1449,In_245,In_674);
and U1450 (N_1450,In_41,In_874);
or U1451 (N_1451,In_0,In_1054);
and U1452 (N_1452,In_1482,In_479);
and U1453 (N_1453,In_919,In_499);
nor U1454 (N_1454,In_933,In_1373);
nor U1455 (N_1455,In_1465,In_795);
and U1456 (N_1456,In_899,In_912);
or U1457 (N_1457,In_295,In_640);
nor U1458 (N_1458,In_723,In_1144);
or U1459 (N_1459,In_933,In_209);
and U1460 (N_1460,In_363,In_538);
nor U1461 (N_1461,In_306,In_1196);
and U1462 (N_1462,In_667,In_364);
and U1463 (N_1463,In_738,In_1053);
or U1464 (N_1464,In_580,In_1098);
nand U1465 (N_1465,In_367,In_312);
or U1466 (N_1466,In_366,In_500);
or U1467 (N_1467,In_654,In_1212);
nand U1468 (N_1468,In_1152,In_571);
nand U1469 (N_1469,In_505,In_831);
xor U1470 (N_1470,In_34,In_391);
or U1471 (N_1471,In_466,In_604);
and U1472 (N_1472,In_1252,In_1368);
and U1473 (N_1473,In_342,In_687);
nor U1474 (N_1474,In_660,In_1435);
nor U1475 (N_1475,In_492,In_765);
nand U1476 (N_1476,In_891,In_1077);
xor U1477 (N_1477,In_595,In_317);
nand U1478 (N_1478,In_1133,In_584);
or U1479 (N_1479,In_465,In_476);
nand U1480 (N_1480,In_114,In_642);
and U1481 (N_1481,In_1418,In_1140);
and U1482 (N_1482,In_6,In_1409);
nor U1483 (N_1483,In_528,In_481);
nand U1484 (N_1484,In_1371,In_499);
nand U1485 (N_1485,In_1481,In_689);
or U1486 (N_1486,In_520,In_182);
nand U1487 (N_1487,In_1072,In_494);
and U1488 (N_1488,In_612,In_3);
and U1489 (N_1489,In_794,In_1173);
nor U1490 (N_1490,In_69,In_747);
and U1491 (N_1491,In_1382,In_253);
and U1492 (N_1492,In_435,In_796);
or U1493 (N_1493,In_614,In_948);
nor U1494 (N_1494,In_857,In_1174);
and U1495 (N_1495,In_779,In_49);
nor U1496 (N_1496,In_1045,In_1038);
nor U1497 (N_1497,In_373,In_767);
or U1498 (N_1498,In_1233,In_181);
or U1499 (N_1499,In_656,In_1118);
nand U1500 (N_1500,In_52,In_170);
nor U1501 (N_1501,In_1057,In_784);
nand U1502 (N_1502,In_552,In_360);
nor U1503 (N_1503,In_260,In_77);
or U1504 (N_1504,In_371,In_244);
or U1505 (N_1505,In_112,In_233);
and U1506 (N_1506,In_905,In_1227);
nand U1507 (N_1507,In_1251,In_712);
nor U1508 (N_1508,In_595,In_371);
nand U1509 (N_1509,In_1279,In_1215);
nand U1510 (N_1510,In_299,In_1024);
or U1511 (N_1511,In_196,In_979);
or U1512 (N_1512,In_1493,In_656);
nor U1513 (N_1513,In_827,In_957);
xnor U1514 (N_1514,In_601,In_719);
nor U1515 (N_1515,In_1304,In_769);
nand U1516 (N_1516,In_631,In_1027);
nor U1517 (N_1517,In_73,In_1130);
nand U1518 (N_1518,In_49,In_396);
nor U1519 (N_1519,In_839,In_890);
nor U1520 (N_1520,In_424,In_502);
nand U1521 (N_1521,In_897,In_972);
nand U1522 (N_1522,In_1234,In_585);
nand U1523 (N_1523,In_1285,In_1277);
nor U1524 (N_1524,In_853,In_582);
and U1525 (N_1525,In_800,In_1475);
nand U1526 (N_1526,In_425,In_102);
nor U1527 (N_1527,In_87,In_419);
nor U1528 (N_1528,In_744,In_1467);
and U1529 (N_1529,In_76,In_821);
or U1530 (N_1530,In_1373,In_825);
nand U1531 (N_1531,In_1129,In_506);
nor U1532 (N_1532,In_775,In_828);
or U1533 (N_1533,In_168,In_894);
or U1534 (N_1534,In_607,In_480);
nor U1535 (N_1535,In_857,In_207);
nand U1536 (N_1536,In_635,In_456);
or U1537 (N_1537,In_356,In_759);
and U1538 (N_1538,In_400,In_528);
or U1539 (N_1539,In_733,In_1141);
and U1540 (N_1540,In_279,In_744);
nor U1541 (N_1541,In_904,In_1026);
or U1542 (N_1542,In_152,In_113);
or U1543 (N_1543,In_539,In_1457);
nor U1544 (N_1544,In_95,In_80);
nor U1545 (N_1545,In_1271,In_1304);
nand U1546 (N_1546,In_146,In_187);
or U1547 (N_1547,In_410,In_1355);
or U1548 (N_1548,In_1493,In_768);
nor U1549 (N_1549,In_1415,In_1459);
nor U1550 (N_1550,In_413,In_274);
and U1551 (N_1551,In_1366,In_538);
nand U1552 (N_1552,In_1464,In_486);
nor U1553 (N_1553,In_407,In_736);
nand U1554 (N_1554,In_1325,In_68);
xor U1555 (N_1555,In_1485,In_120);
nor U1556 (N_1556,In_554,In_843);
nor U1557 (N_1557,In_208,In_944);
nand U1558 (N_1558,In_333,In_1244);
nor U1559 (N_1559,In_982,In_887);
nand U1560 (N_1560,In_1252,In_91);
nor U1561 (N_1561,In_1274,In_766);
nand U1562 (N_1562,In_465,In_641);
xor U1563 (N_1563,In_222,In_2);
or U1564 (N_1564,In_154,In_523);
nand U1565 (N_1565,In_24,In_1044);
nand U1566 (N_1566,In_613,In_1126);
nor U1567 (N_1567,In_860,In_1243);
and U1568 (N_1568,In_817,In_648);
nand U1569 (N_1569,In_1015,In_252);
or U1570 (N_1570,In_575,In_766);
or U1571 (N_1571,In_1001,In_716);
nor U1572 (N_1572,In_1421,In_295);
nor U1573 (N_1573,In_351,In_985);
nand U1574 (N_1574,In_631,In_1325);
and U1575 (N_1575,In_29,In_198);
or U1576 (N_1576,In_1313,In_630);
nor U1577 (N_1577,In_546,In_290);
nand U1578 (N_1578,In_153,In_559);
nor U1579 (N_1579,In_103,In_130);
nor U1580 (N_1580,In_1256,In_718);
nor U1581 (N_1581,In_785,In_212);
and U1582 (N_1582,In_1149,In_399);
nand U1583 (N_1583,In_930,In_84);
nand U1584 (N_1584,In_665,In_1097);
nor U1585 (N_1585,In_111,In_1224);
or U1586 (N_1586,In_1347,In_1280);
nor U1587 (N_1587,In_804,In_422);
nand U1588 (N_1588,In_1231,In_981);
and U1589 (N_1589,In_292,In_1232);
nand U1590 (N_1590,In_870,In_549);
xor U1591 (N_1591,In_147,In_65);
nor U1592 (N_1592,In_1024,In_1372);
xor U1593 (N_1593,In_1315,In_143);
and U1594 (N_1594,In_144,In_1148);
nand U1595 (N_1595,In_836,In_232);
nor U1596 (N_1596,In_701,In_1139);
and U1597 (N_1597,In_1235,In_558);
xnor U1598 (N_1598,In_223,In_970);
nor U1599 (N_1599,In_516,In_830);
nor U1600 (N_1600,In_359,In_1114);
and U1601 (N_1601,In_1190,In_1410);
and U1602 (N_1602,In_50,In_851);
nand U1603 (N_1603,In_419,In_576);
xnor U1604 (N_1604,In_379,In_628);
nor U1605 (N_1605,In_211,In_868);
nand U1606 (N_1606,In_48,In_134);
nand U1607 (N_1607,In_473,In_70);
and U1608 (N_1608,In_627,In_466);
nor U1609 (N_1609,In_522,In_224);
nor U1610 (N_1610,In_852,In_1123);
and U1611 (N_1611,In_945,In_573);
or U1612 (N_1612,In_1342,In_237);
and U1613 (N_1613,In_1280,In_1107);
nand U1614 (N_1614,In_1196,In_1326);
nor U1615 (N_1615,In_37,In_1331);
nand U1616 (N_1616,In_1108,In_780);
nor U1617 (N_1617,In_759,In_1186);
nor U1618 (N_1618,In_391,In_1490);
and U1619 (N_1619,In_79,In_449);
or U1620 (N_1620,In_996,In_1383);
nand U1621 (N_1621,In_1071,In_1226);
or U1622 (N_1622,In_548,In_195);
and U1623 (N_1623,In_1262,In_1001);
or U1624 (N_1624,In_1420,In_1023);
or U1625 (N_1625,In_1350,In_908);
and U1626 (N_1626,In_11,In_419);
or U1627 (N_1627,In_1310,In_711);
or U1628 (N_1628,In_1312,In_1266);
or U1629 (N_1629,In_387,In_763);
and U1630 (N_1630,In_779,In_669);
or U1631 (N_1631,In_399,In_1472);
nand U1632 (N_1632,In_271,In_630);
nand U1633 (N_1633,In_1113,In_668);
or U1634 (N_1634,In_468,In_1288);
or U1635 (N_1635,In_807,In_817);
nor U1636 (N_1636,In_1329,In_511);
or U1637 (N_1637,In_767,In_1003);
nand U1638 (N_1638,In_501,In_1249);
or U1639 (N_1639,In_769,In_638);
and U1640 (N_1640,In_961,In_61);
and U1641 (N_1641,In_894,In_1372);
and U1642 (N_1642,In_458,In_327);
or U1643 (N_1643,In_1458,In_282);
nand U1644 (N_1644,In_1496,In_1469);
and U1645 (N_1645,In_1375,In_1058);
and U1646 (N_1646,In_155,In_1241);
or U1647 (N_1647,In_1271,In_1452);
nor U1648 (N_1648,In_977,In_306);
and U1649 (N_1649,In_283,In_1412);
or U1650 (N_1650,In_404,In_44);
nand U1651 (N_1651,In_1228,In_357);
nor U1652 (N_1652,In_187,In_877);
and U1653 (N_1653,In_127,In_1337);
nand U1654 (N_1654,In_230,In_885);
and U1655 (N_1655,In_1174,In_846);
nor U1656 (N_1656,In_983,In_1276);
nand U1657 (N_1657,In_245,In_904);
or U1658 (N_1658,In_253,In_1100);
nor U1659 (N_1659,In_376,In_1313);
and U1660 (N_1660,In_689,In_62);
and U1661 (N_1661,In_1411,In_1325);
or U1662 (N_1662,In_1292,In_911);
nand U1663 (N_1663,In_620,In_1367);
and U1664 (N_1664,In_1168,In_1113);
nor U1665 (N_1665,In_147,In_333);
or U1666 (N_1666,In_1222,In_368);
or U1667 (N_1667,In_602,In_488);
nand U1668 (N_1668,In_930,In_1453);
or U1669 (N_1669,In_1069,In_1183);
nor U1670 (N_1670,In_895,In_62);
nor U1671 (N_1671,In_475,In_87);
nor U1672 (N_1672,In_1254,In_444);
and U1673 (N_1673,In_783,In_14);
or U1674 (N_1674,In_1293,In_405);
or U1675 (N_1675,In_1368,In_790);
and U1676 (N_1676,In_1001,In_38);
or U1677 (N_1677,In_612,In_1466);
nor U1678 (N_1678,In_1108,In_1484);
nand U1679 (N_1679,In_668,In_144);
and U1680 (N_1680,In_84,In_277);
and U1681 (N_1681,In_1364,In_750);
or U1682 (N_1682,In_991,In_389);
nor U1683 (N_1683,In_1126,In_1074);
or U1684 (N_1684,In_1321,In_1044);
nand U1685 (N_1685,In_100,In_1236);
nand U1686 (N_1686,In_414,In_1071);
nand U1687 (N_1687,In_69,In_511);
or U1688 (N_1688,In_338,In_951);
nor U1689 (N_1689,In_1278,In_1463);
nand U1690 (N_1690,In_492,In_358);
or U1691 (N_1691,In_410,In_892);
and U1692 (N_1692,In_769,In_309);
nor U1693 (N_1693,In_1022,In_1086);
and U1694 (N_1694,In_117,In_144);
nor U1695 (N_1695,In_673,In_270);
nand U1696 (N_1696,In_426,In_465);
nor U1697 (N_1697,In_529,In_660);
or U1698 (N_1698,In_1193,In_213);
and U1699 (N_1699,In_170,In_1260);
or U1700 (N_1700,In_251,In_138);
or U1701 (N_1701,In_558,In_1499);
or U1702 (N_1702,In_672,In_541);
nor U1703 (N_1703,In_1158,In_323);
and U1704 (N_1704,In_136,In_405);
nor U1705 (N_1705,In_854,In_54);
nand U1706 (N_1706,In_1066,In_590);
nand U1707 (N_1707,In_1470,In_671);
or U1708 (N_1708,In_878,In_1115);
nand U1709 (N_1709,In_704,In_1145);
nor U1710 (N_1710,In_1106,In_1286);
nor U1711 (N_1711,In_1052,In_1332);
and U1712 (N_1712,In_554,In_28);
or U1713 (N_1713,In_221,In_419);
nor U1714 (N_1714,In_1367,In_885);
and U1715 (N_1715,In_832,In_628);
nand U1716 (N_1716,In_515,In_699);
nand U1717 (N_1717,In_848,In_476);
nand U1718 (N_1718,In_400,In_1476);
or U1719 (N_1719,In_1309,In_1494);
or U1720 (N_1720,In_1135,In_1184);
nand U1721 (N_1721,In_96,In_279);
and U1722 (N_1722,In_516,In_157);
and U1723 (N_1723,In_56,In_1347);
nand U1724 (N_1724,In_1465,In_854);
and U1725 (N_1725,In_1025,In_1210);
nand U1726 (N_1726,In_839,In_1247);
nand U1727 (N_1727,In_253,In_963);
and U1728 (N_1728,In_1419,In_315);
nor U1729 (N_1729,In_434,In_646);
nor U1730 (N_1730,In_551,In_1106);
and U1731 (N_1731,In_460,In_337);
or U1732 (N_1732,In_64,In_1427);
nand U1733 (N_1733,In_435,In_650);
or U1734 (N_1734,In_981,In_501);
nor U1735 (N_1735,In_916,In_510);
nand U1736 (N_1736,In_442,In_775);
nand U1737 (N_1737,In_1279,In_453);
nor U1738 (N_1738,In_347,In_819);
nor U1739 (N_1739,In_306,In_345);
nand U1740 (N_1740,In_1341,In_37);
and U1741 (N_1741,In_722,In_783);
nor U1742 (N_1742,In_345,In_1019);
nor U1743 (N_1743,In_1178,In_1297);
and U1744 (N_1744,In_621,In_207);
and U1745 (N_1745,In_867,In_412);
nor U1746 (N_1746,In_1262,In_1225);
nand U1747 (N_1747,In_1263,In_1037);
nor U1748 (N_1748,In_662,In_1394);
nand U1749 (N_1749,In_1230,In_711);
and U1750 (N_1750,In_630,In_593);
or U1751 (N_1751,In_688,In_1220);
nand U1752 (N_1752,In_385,In_369);
or U1753 (N_1753,In_850,In_1377);
and U1754 (N_1754,In_1239,In_1182);
or U1755 (N_1755,In_527,In_88);
or U1756 (N_1756,In_347,In_215);
nor U1757 (N_1757,In_1130,In_267);
nand U1758 (N_1758,In_931,In_1223);
nor U1759 (N_1759,In_634,In_843);
nand U1760 (N_1760,In_1348,In_953);
nor U1761 (N_1761,In_277,In_1037);
nor U1762 (N_1762,In_1285,In_527);
or U1763 (N_1763,In_860,In_888);
nor U1764 (N_1764,In_1413,In_1167);
or U1765 (N_1765,In_996,In_459);
or U1766 (N_1766,In_43,In_1179);
nor U1767 (N_1767,In_299,In_816);
or U1768 (N_1768,In_484,In_715);
and U1769 (N_1769,In_1471,In_1130);
and U1770 (N_1770,In_597,In_572);
nor U1771 (N_1771,In_619,In_309);
nand U1772 (N_1772,In_1095,In_367);
or U1773 (N_1773,In_50,In_746);
and U1774 (N_1774,In_582,In_772);
nor U1775 (N_1775,In_309,In_96);
nor U1776 (N_1776,In_51,In_294);
or U1777 (N_1777,In_1050,In_689);
or U1778 (N_1778,In_83,In_1251);
or U1779 (N_1779,In_75,In_294);
or U1780 (N_1780,In_1235,In_399);
and U1781 (N_1781,In_312,In_896);
nand U1782 (N_1782,In_1406,In_395);
and U1783 (N_1783,In_600,In_751);
nor U1784 (N_1784,In_721,In_182);
or U1785 (N_1785,In_916,In_1021);
nand U1786 (N_1786,In_512,In_788);
and U1787 (N_1787,In_936,In_1255);
or U1788 (N_1788,In_540,In_289);
nand U1789 (N_1789,In_853,In_1035);
nor U1790 (N_1790,In_702,In_1346);
and U1791 (N_1791,In_579,In_279);
nor U1792 (N_1792,In_387,In_866);
nand U1793 (N_1793,In_1145,In_341);
nor U1794 (N_1794,In_570,In_688);
and U1795 (N_1795,In_235,In_1352);
nor U1796 (N_1796,In_155,In_624);
and U1797 (N_1797,In_600,In_1325);
nand U1798 (N_1798,In_351,In_1242);
and U1799 (N_1799,In_217,In_407);
nor U1800 (N_1800,In_994,In_642);
and U1801 (N_1801,In_705,In_342);
nand U1802 (N_1802,In_997,In_420);
nor U1803 (N_1803,In_761,In_946);
nand U1804 (N_1804,In_344,In_1192);
nor U1805 (N_1805,In_672,In_486);
nor U1806 (N_1806,In_1348,In_261);
or U1807 (N_1807,In_1479,In_1279);
or U1808 (N_1808,In_714,In_1281);
and U1809 (N_1809,In_1460,In_635);
nor U1810 (N_1810,In_599,In_441);
or U1811 (N_1811,In_775,In_462);
nor U1812 (N_1812,In_801,In_895);
nor U1813 (N_1813,In_738,In_30);
or U1814 (N_1814,In_1188,In_1265);
or U1815 (N_1815,In_139,In_576);
or U1816 (N_1816,In_1245,In_1257);
nor U1817 (N_1817,In_1393,In_625);
and U1818 (N_1818,In_1335,In_1072);
or U1819 (N_1819,In_966,In_644);
or U1820 (N_1820,In_48,In_1256);
or U1821 (N_1821,In_414,In_145);
nand U1822 (N_1822,In_897,In_551);
nand U1823 (N_1823,In_165,In_1170);
nor U1824 (N_1824,In_1388,In_252);
nand U1825 (N_1825,In_399,In_252);
and U1826 (N_1826,In_1139,In_977);
nor U1827 (N_1827,In_1470,In_1386);
or U1828 (N_1828,In_1053,In_128);
or U1829 (N_1829,In_1112,In_1309);
and U1830 (N_1830,In_877,In_154);
nor U1831 (N_1831,In_745,In_867);
xor U1832 (N_1832,In_994,In_1373);
or U1833 (N_1833,In_1382,In_601);
or U1834 (N_1834,In_899,In_1075);
nor U1835 (N_1835,In_782,In_117);
nor U1836 (N_1836,In_355,In_924);
nor U1837 (N_1837,In_866,In_404);
and U1838 (N_1838,In_761,In_339);
and U1839 (N_1839,In_1194,In_654);
nand U1840 (N_1840,In_31,In_210);
or U1841 (N_1841,In_576,In_922);
and U1842 (N_1842,In_574,In_749);
nor U1843 (N_1843,In_933,In_33);
and U1844 (N_1844,In_914,In_469);
nor U1845 (N_1845,In_1025,In_1199);
and U1846 (N_1846,In_825,In_1353);
nor U1847 (N_1847,In_375,In_673);
nand U1848 (N_1848,In_1460,In_1033);
nand U1849 (N_1849,In_123,In_757);
or U1850 (N_1850,In_866,In_781);
or U1851 (N_1851,In_169,In_1038);
nor U1852 (N_1852,In_947,In_1093);
or U1853 (N_1853,In_545,In_466);
and U1854 (N_1854,In_846,In_1237);
nand U1855 (N_1855,In_409,In_1156);
nand U1856 (N_1856,In_280,In_52);
and U1857 (N_1857,In_581,In_1025);
and U1858 (N_1858,In_1062,In_510);
nand U1859 (N_1859,In_1021,In_1209);
or U1860 (N_1860,In_263,In_1263);
nor U1861 (N_1861,In_729,In_1392);
or U1862 (N_1862,In_1190,In_316);
nand U1863 (N_1863,In_749,In_919);
or U1864 (N_1864,In_156,In_1180);
or U1865 (N_1865,In_1420,In_159);
and U1866 (N_1866,In_1189,In_1261);
nand U1867 (N_1867,In_1419,In_889);
nand U1868 (N_1868,In_546,In_1412);
nand U1869 (N_1869,In_1188,In_674);
and U1870 (N_1870,In_457,In_1248);
nand U1871 (N_1871,In_459,In_8);
and U1872 (N_1872,In_702,In_1120);
nand U1873 (N_1873,In_96,In_1427);
and U1874 (N_1874,In_317,In_873);
nand U1875 (N_1875,In_702,In_500);
or U1876 (N_1876,In_179,In_908);
nand U1877 (N_1877,In_185,In_338);
nor U1878 (N_1878,In_686,In_580);
or U1879 (N_1879,In_334,In_355);
nor U1880 (N_1880,In_846,In_1345);
nor U1881 (N_1881,In_496,In_625);
nor U1882 (N_1882,In_1456,In_330);
or U1883 (N_1883,In_85,In_698);
nand U1884 (N_1884,In_1371,In_502);
or U1885 (N_1885,In_0,In_680);
and U1886 (N_1886,In_366,In_1183);
and U1887 (N_1887,In_1477,In_501);
nand U1888 (N_1888,In_1241,In_1052);
nor U1889 (N_1889,In_954,In_1183);
or U1890 (N_1890,In_487,In_737);
xor U1891 (N_1891,In_55,In_1352);
nand U1892 (N_1892,In_274,In_580);
or U1893 (N_1893,In_928,In_843);
or U1894 (N_1894,In_581,In_559);
and U1895 (N_1895,In_812,In_914);
or U1896 (N_1896,In_976,In_522);
or U1897 (N_1897,In_1315,In_648);
and U1898 (N_1898,In_1198,In_1456);
nand U1899 (N_1899,In_811,In_5);
and U1900 (N_1900,In_1245,In_783);
nand U1901 (N_1901,In_317,In_218);
or U1902 (N_1902,In_579,In_930);
nor U1903 (N_1903,In_750,In_1490);
nor U1904 (N_1904,In_262,In_516);
nand U1905 (N_1905,In_1448,In_1375);
or U1906 (N_1906,In_441,In_629);
nand U1907 (N_1907,In_181,In_858);
nand U1908 (N_1908,In_460,In_1476);
nor U1909 (N_1909,In_965,In_250);
nor U1910 (N_1910,In_677,In_792);
and U1911 (N_1911,In_472,In_1201);
or U1912 (N_1912,In_633,In_686);
nand U1913 (N_1913,In_826,In_1283);
nor U1914 (N_1914,In_831,In_476);
nor U1915 (N_1915,In_1126,In_1003);
or U1916 (N_1916,In_1255,In_167);
and U1917 (N_1917,In_1329,In_464);
and U1918 (N_1918,In_904,In_771);
nand U1919 (N_1919,In_748,In_491);
or U1920 (N_1920,In_1218,In_1464);
and U1921 (N_1921,In_1439,In_917);
and U1922 (N_1922,In_517,In_1286);
or U1923 (N_1923,In_1139,In_1317);
nand U1924 (N_1924,In_115,In_147);
nor U1925 (N_1925,In_209,In_1109);
nor U1926 (N_1926,In_360,In_1184);
and U1927 (N_1927,In_1079,In_699);
and U1928 (N_1928,In_451,In_1356);
or U1929 (N_1929,In_583,In_974);
nand U1930 (N_1930,In_116,In_703);
nand U1931 (N_1931,In_950,In_450);
nor U1932 (N_1932,In_122,In_938);
nor U1933 (N_1933,In_804,In_1194);
nand U1934 (N_1934,In_785,In_517);
nand U1935 (N_1935,In_424,In_319);
nor U1936 (N_1936,In_493,In_732);
nor U1937 (N_1937,In_469,In_305);
nor U1938 (N_1938,In_806,In_72);
or U1939 (N_1939,In_303,In_490);
nand U1940 (N_1940,In_1473,In_533);
nor U1941 (N_1941,In_1300,In_853);
nand U1942 (N_1942,In_1371,In_1403);
nand U1943 (N_1943,In_42,In_531);
nor U1944 (N_1944,In_906,In_1402);
or U1945 (N_1945,In_174,In_244);
or U1946 (N_1946,In_1400,In_856);
nor U1947 (N_1947,In_1114,In_0);
and U1948 (N_1948,In_1344,In_954);
and U1949 (N_1949,In_723,In_978);
nor U1950 (N_1950,In_708,In_772);
and U1951 (N_1951,In_52,In_1475);
nand U1952 (N_1952,In_1260,In_578);
and U1953 (N_1953,In_1330,In_1302);
nor U1954 (N_1954,In_1134,In_475);
and U1955 (N_1955,In_1201,In_317);
nand U1956 (N_1956,In_420,In_1313);
or U1957 (N_1957,In_135,In_917);
nor U1958 (N_1958,In_369,In_968);
and U1959 (N_1959,In_63,In_703);
nand U1960 (N_1960,In_333,In_646);
xor U1961 (N_1961,In_1350,In_649);
and U1962 (N_1962,In_964,In_546);
nand U1963 (N_1963,In_342,In_52);
or U1964 (N_1964,In_236,In_47);
or U1965 (N_1965,In_208,In_1110);
or U1966 (N_1966,In_552,In_595);
or U1967 (N_1967,In_872,In_192);
or U1968 (N_1968,In_75,In_157);
nor U1969 (N_1969,In_215,In_998);
nand U1970 (N_1970,In_63,In_1227);
xor U1971 (N_1971,In_1024,In_707);
nor U1972 (N_1972,In_14,In_305);
nand U1973 (N_1973,In_298,In_859);
and U1974 (N_1974,In_788,In_22);
nor U1975 (N_1975,In_789,In_186);
and U1976 (N_1976,In_656,In_1099);
and U1977 (N_1977,In_662,In_49);
nor U1978 (N_1978,In_276,In_1303);
nand U1979 (N_1979,In_391,In_337);
and U1980 (N_1980,In_980,In_683);
and U1981 (N_1981,In_826,In_913);
nor U1982 (N_1982,In_908,In_6);
or U1983 (N_1983,In_24,In_723);
and U1984 (N_1984,In_1282,In_1350);
nand U1985 (N_1985,In_445,In_470);
and U1986 (N_1986,In_176,In_621);
nand U1987 (N_1987,In_1330,In_1232);
nor U1988 (N_1988,In_1258,In_481);
nor U1989 (N_1989,In_32,In_357);
nand U1990 (N_1990,In_187,In_756);
nor U1991 (N_1991,In_126,In_1248);
or U1992 (N_1992,In_931,In_663);
and U1993 (N_1993,In_581,In_1028);
nand U1994 (N_1994,In_830,In_831);
and U1995 (N_1995,In_1388,In_501);
nor U1996 (N_1996,In_238,In_200);
nand U1997 (N_1997,In_1489,In_884);
and U1998 (N_1998,In_700,In_843);
or U1999 (N_1999,In_1108,In_850);
and U2000 (N_2000,In_896,In_690);
and U2001 (N_2001,In_343,In_198);
and U2002 (N_2002,In_839,In_382);
or U2003 (N_2003,In_1420,In_1022);
nor U2004 (N_2004,In_938,In_1029);
nor U2005 (N_2005,In_1074,In_404);
nor U2006 (N_2006,In_56,In_1493);
and U2007 (N_2007,In_193,In_1390);
and U2008 (N_2008,In_1281,In_1120);
or U2009 (N_2009,In_330,In_660);
or U2010 (N_2010,In_1128,In_1246);
and U2011 (N_2011,In_1258,In_765);
nand U2012 (N_2012,In_97,In_1113);
nor U2013 (N_2013,In_216,In_1184);
nand U2014 (N_2014,In_206,In_989);
nand U2015 (N_2015,In_1347,In_138);
nor U2016 (N_2016,In_1473,In_445);
nor U2017 (N_2017,In_434,In_8);
nor U2018 (N_2018,In_256,In_1177);
nor U2019 (N_2019,In_1133,In_150);
nor U2020 (N_2020,In_596,In_515);
nor U2021 (N_2021,In_430,In_1247);
nor U2022 (N_2022,In_332,In_1203);
nor U2023 (N_2023,In_130,In_1145);
or U2024 (N_2024,In_1420,In_209);
or U2025 (N_2025,In_363,In_800);
and U2026 (N_2026,In_532,In_1343);
and U2027 (N_2027,In_1235,In_1026);
nand U2028 (N_2028,In_15,In_660);
or U2029 (N_2029,In_1169,In_931);
nor U2030 (N_2030,In_1355,In_866);
or U2031 (N_2031,In_488,In_1043);
or U2032 (N_2032,In_294,In_514);
nor U2033 (N_2033,In_907,In_1080);
nor U2034 (N_2034,In_753,In_1268);
nand U2035 (N_2035,In_515,In_1373);
or U2036 (N_2036,In_526,In_578);
and U2037 (N_2037,In_152,In_238);
nor U2038 (N_2038,In_879,In_636);
nor U2039 (N_2039,In_1379,In_366);
and U2040 (N_2040,In_912,In_1132);
nor U2041 (N_2041,In_1468,In_53);
and U2042 (N_2042,In_687,In_572);
or U2043 (N_2043,In_457,In_62);
nand U2044 (N_2044,In_751,In_501);
or U2045 (N_2045,In_1326,In_103);
or U2046 (N_2046,In_384,In_775);
nor U2047 (N_2047,In_509,In_873);
nor U2048 (N_2048,In_442,In_940);
and U2049 (N_2049,In_93,In_105);
nand U2050 (N_2050,In_604,In_1065);
nor U2051 (N_2051,In_160,In_296);
and U2052 (N_2052,In_543,In_142);
or U2053 (N_2053,In_1273,In_61);
nand U2054 (N_2054,In_878,In_651);
and U2055 (N_2055,In_676,In_179);
nor U2056 (N_2056,In_1410,In_799);
nor U2057 (N_2057,In_1177,In_1330);
nand U2058 (N_2058,In_90,In_112);
nor U2059 (N_2059,In_190,In_174);
and U2060 (N_2060,In_400,In_334);
xor U2061 (N_2061,In_885,In_1243);
or U2062 (N_2062,In_1164,In_1086);
and U2063 (N_2063,In_723,In_1478);
nand U2064 (N_2064,In_922,In_626);
nand U2065 (N_2065,In_400,In_804);
nor U2066 (N_2066,In_101,In_266);
nor U2067 (N_2067,In_505,In_1047);
nand U2068 (N_2068,In_553,In_1204);
and U2069 (N_2069,In_893,In_692);
nand U2070 (N_2070,In_867,In_262);
and U2071 (N_2071,In_1390,In_1123);
or U2072 (N_2072,In_451,In_426);
or U2073 (N_2073,In_800,In_1479);
nand U2074 (N_2074,In_305,In_1423);
nand U2075 (N_2075,In_1244,In_116);
or U2076 (N_2076,In_836,In_782);
nand U2077 (N_2077,In_1470,In_1049);
nor U2078 (N_2078,In_280,In_200);
and U2079 (N_2079,In_1113,In_571);
and U2080 (N_2080,In_1191,In_797);
or U2081 (N_2081,In_863,In_569);
and U2082 (N_2082,In_1371,In_197);
xnor U2083 (N_2083,In_24,In_546);
and U2084 (N_2084,In_280,In_1255);
or U2085 (N_2085,In_326,In_1001);
and U2086 (N_2086,In_944,In_1397);
or U2087 (N_2087,In_938,In_788);
or U2088 (N_2088,In_1459,In_1092);
nand U2089 (N_2089,In_1122,In_1130);
nor U2090 (N_2090,In_297,In_958);
and U2091 (N_2091,In_1257,In_294);
or U2092 (N_2092,In_353,In_1496);
or U2093 (N_2093,In_507,In_139);
nor U2094 (N_2094,In_1111,In_254);
xor U2095 (N_2095,In_1276,In_595);
nand U2096 (N_2096,In_791,In_6);
and U2097 (N_2097,In_532,In_270);
nor U2098 (N_2098,In_1488,In_166);
and U2099 (N_2099,In_101,In_842);
nor U2100 (N_2100,In_981,In_1232);
and U2101 (N_2101,In_1317,In_1056);
nor U2102 (N_2102,In_100,In_1330);
or U2103 (N_2103,In_482,In_1129);
or U2104 (N_2104,In_1347,In_1328);
nand U2105 (N_2105,In_900,In_1257);
nand U2106 (N_2106,In_818,In_1338);
nand U2107 (N_2107,In_241,In_1288);
or U2108 (N_2108,In_947,In_1225);
nand U2109 (N_2109,In_1426,In_1462);
and U2110 (N_2110,In_679,In_365);
and U2111 (N_2111,In_498,In_1483);
and U2112 (N_2112,In_726,In_1078);
and U2113 (N_2113,In_1326,In_227);
nand U2114 (N_2114,In_1362,In_1280);
nor U2115 (N_2115,In_1319,In_367);
nor U2116 (N_2116,In_1461,In_614);
nor U2117 (N_2117,In_1040,In_78);
or U2118 (N_2118,In_300,In_1091);
and U2119 (N_2119,In_20,In_1366);
or U2120 (N_2120,In_1216,In_1328);
nand U2121 (N_2121,In_265,In_848);
or U2122 (N_2122,In_1075,In_264);
or U2123 (N_2123,In_45,In_1086);
and U2124 (N_2124,In_23,In_641);
or U2125 (N_2125,In_1414,In_643);
nand U2126 (N_2126,In_430,In_482);
nand U2127 (N_2127,In_1172,In_156);
and U2128 (N_2128,In_30,In_513);
and U2129 (N_2129,In_1376,In_1471);
nand U2130 (N_2130,In_158,In_1338);
nor U2131 (N_2131,In_312,In_1084);
and U2132 (N_2132,In_475,In_405);
nor U2133 (N_2133,In_549,In_1139);
or U2134 (N_2134,In_1139,In_881);
or U2135 (N_2135,In_1343,In_708);
nand U2136 (N_2136,In_1004,In_863);
nand U2137 (N_2137,In_1103,In_701);
nor U2138 (N_2138,In_541,In_1054);
nor U2139 (N_2139,In_266,In_1207);
or U2140 (N_2140,In_895,In_1009);
or U2141 (N_2141,In_1373,In_553);
or U2142 (N_2142,In_241,In_870);
nand U2143 (N_2143,In_203,In_14);
nand U2144 (N_2144,In_1224,In_440);
nor U2145 (N_2145,In_575,In_384);
nor U2146 (N_2146,In_648,In_892);
nor U2147 (N_2147,In_1323,In_1357);
or U2148 (N_2148,In_265,In_885);
or U2149 (N_2149,In_198,In_820);
nor U2150 (N_2150,In_783,In_921);
nand U2151 (N_2151,In_1131,In_1128);
nand U2152 (N_2152,In_858,In_1314);
nor U2153 (N_2153,In_797,In_1107);
nand U2154 (N_2154,In_1247,In_555);
and U2155 (N_2155,In_495,In_163);
xor U2156 (N_2156,In_543,In_1355);
or U2157 (N_2157,In_1358,In_888);
nor U2158 (N_2158,In_754,In_668);
nor U2159 (N_2159,In_109,In_1489);
nand U2160 (N_2160,In_627,In_930);
nor U2161 (N_2161,In_640,In_1385);
or U2162 (N_2162,In_1124,In_798);
nor U2163 (N_2163,In_1000,In_948);
nor U2164 (N_2164,In_295,In_1116);
nand U2165 (N_2165,In_1,In_1449);
nor U2166 (N_2166,In_1208,In_579);
nand U2167 (N_2167,In_537,In_499);
nand U2168 (N_2168,In_839,In_194);
or U2169 (N_2169,In_1121,In_749);
or U2170 (N_2170,In_551,In_1072);
nor U2171 (N_2171,In_22,In_1015);
nand U2172 (N_2172,In_1214,In_1021);
and U2173 (N_2173,In_1384,In_1055);
and U2174 (N_2174,In_675,In_711);
nor U2175 (N_2175,In_574,In_1312);
or U2176 (N_2176,In_975,In_314);
nor U2177 (N_2177,In_74,In_1050);
nand U2178 (N_2178,In_814,In_515);
and U2179 (N_2179,In_124,In_703);
and U2180 (N_2180,In_643,In_360);
or U2181 (N_2181,In_345,In_1096);
nand U2182 (N_2182,In_53,In_713);
or U2183 (N_2183,In_293,In_1270);
nand U2184 (N_2184,In_316,In_1046);
or U2185 (N_2185,In_769,In_1048);
nor U2186 (N_2186,In_966,In_518);
xor U2187 (N_2187,In_998,In_769);
and U2188 (N_2188,In_478,In_744);
and U2189 (N_2189,In_1157,In_346);
nor U2190 (N_2190,In_840,In_1386);
nand U2191 (N_2191,In_1135,In_127);
or U2192 (N_2192,In_849,In_1403);
and U2193 (N_2193,In_605,In_875);
nor U2194 (N_2194,In_1074,In_294);
and U2195 (N_2195,In_604,In_859);
nand U2196 (N_2196,In_1309,In_434);
nor U2197 (N_2197,In_54,In_800);
nand U2198 (N_2198,In_685,In_169);
nand U2199 (N_2199,In_90,In_665);
and U2200 (N_2200,In_65,In_186);
and U2201 (N_2201,In_415,In_1084);
nand U2202 (N_2202,In_1225,In_661);
and U2203 (N_2203,In_457,In_546);
and U2204 (N_2204,In_38,In_480);
nand U2205 (N_2205,In_334,In_276);
nor U2206 (N_2206,In_9,In_613);
nor U2207 (N_2207,In_966,In_714);
nand U2208 (N_2208,In_364,In_950);
nor U2209 (N_2209,In_1492,In_257);
or U2210 (N_2210,In_1010,In_554);
and U2211 (N_2211,In_290,In_1095);
or U2212 (N_2212,In_991,In_385);
nor U2213 (N_2213,In_216,In_75);
or U2214 (N_2214,In_1215,In_758);
and U2215 (N_2215,In_1159,In_1258);
nand U2216 (N_2216,In_1480,In_380);
nor U2217 (N_2217,In_320,In_796);
or U2218 (N_2218,In_1083,In_1218);
or U2219 (N_2219,In_417,In_99);
nand U2220 (N_2220,In_95,In_106);
or U2221 (N_2221,In_654,In_1146);
or U2222 (N_2222,In_113,In_1057);
nor U2223 (N_2223,In_1354,In_1281);
or U2224 (N_2224,In_939,In_1155);
xor U2225 (N_2225,In_162,In_1075);
or U2226 (N_2226,In_900,In_745);
nor U2227 (N_2227,In_425,In_499);
or U2228 (N_2228,In_370,In_1085);
nor U2229 (N_2229,In_160,In_1321);
nor U2230 (N_2230,In_159,In_1038);
nor U2231 (N_2231,In_352,In_873);
nand U2232 (N_2232,In_309,In_559);
xor U2233 (N_2233,In_178,In_594);
nor U2234 (N_2234,In_947,In_1339);
nor U2235 (N_2235,In_158,In_236);
and U2236 (N_2236,In_634,In_112);
nor U2237 (N_2237,In_1311,In_923);
nor U2238 (N_2238,In_823,In_322);
or U2239 (N_2239,In_1377,In_449);
nand U2240 (N_2240,In_977,In_1440);
nor U2241 (N_2241,In_613,In_1047);
nand U2242 (N_2242,In_1180,In_498);
or U2243 (N_2243,In_1483,In_736);
nor U2244 (N_2244,In_502,In_1392);
nor U2245 (N_2245,In_1245,In_535);
or U2246 (N_2246,In_319,In_1482);
or U2247 (N_2247,In_278,In_287);
nor U2248 (N_2248,In_140,In_767);
and U2249 (N_2249,In_470,In_877);
nor U2250 (N_2250,In_453,In_1027);
nand U2251 (N_2251,In_108,In_1251);
and U2252 (N_2252,In_178,In_608);
and U2253 (N_2253,In_960,In_1065);
or U2254 (N_2254,In_946,In_879);
nor U2255 (N_2255,In_789,In_1402);
nand U2256 (N_2256,In_1043,In_709);
nor U2257 (N_2257,In_574,In_1202);
or U2258 (N_2258,In_965,In_1391);
or U2259 (N_2259,In_1023,In_1488);
and U2260 (N_2260,In_258,In_1241);
nor U2261 (N_2261,In_1429,In_871);
nand U2262 (N_2262,In_571,In_736);
and U2263 (N_2263,In_344,In_1375);
nor U2264 (N_2264,In_108,In_507);
nand U2265 (N_2265,In_769,In_525);
and U2266 (N_2266,In_1455,In_482);
nand U2267 (N_2267,In_1079,In_1411);
nor U2268 (N_2268,In_375,In_1328);
or U2269 (N_2269,In_1001,In_1339);
nand U2270 (N_2270,In_1242,In_1463);
nor U2271 (N_2271,In_196,In_229);
nand U2272 (N_2272,In_1160,In_37);
nor U2273 (N_2273,In_1092,In_125);
or U2274 (N_2274,In_1009,In_991);
and U2275 (N_2275,In_428,In_1177);
nand U2276 (N_2276,In_113,In_1433);
and U2277 (N_2277,In_169,In_1290);
or U2278 (N_2278,In_56,In_505);
nand U2279 (N_2279,In_238,In_1136);
and U2280 (N_2280,In_607,In_555);
and U2281 (N_2281,In_1303,In_1015);
or U2282 (N_2282,In_732,In_252);
or U2283 (N_2283,In_128,In_1329);
nor U2284 (N_2284,In_1359,In_76);
or U2285 (N_2285,In_1048,In_60);
nor U2286 (N_2286,In_185,In_621);
or U2287 (N_2287,In_1150,In_1468);
nand U2288 (N_2288,In_90,In_1338);
nor U2289 (N_2289,In_48,In_96);
and U2290 (N_2290,In_1029,In_48);
nand U2291 (N_2291,In_352,In_756);
nor U2292 (N_2292,In_914,In_24);
nor U2293 (N_2293,In_677,In_313);
nor U2294 (N_2294,In_1422,In_1217);
or U2295 (N_2295,In_629,In_508);
and U2296 (N_2296,In_611,In_566);
nor U2297 (N_2297,In_1491,In_798);
or U2298 (N_2298,In_849,In_911);
or U2299 (N_2299,In_638,In_217);
or U2300 (N_2300,In_634,In_41);
nor U2301 (N_2301,In_554,In_1125);
nand U2302 (N_2302,In_756,In_1082);
and U2303 (N_2303,In_1241,In_461);
and U2304 (N_2304,In_1069,In_230);
or U2305 (N_2305,In_289,In_678);
xor U2306 (N_2306,In_428,In_1218);
nand U2307 (N_2307,In_1220,In_1420);
or U2308 (N_2308,In_1361,In_989);
nand U2309 (N_2309,In_542,In_1002);
nand U2310 (N_2310,In_330,In_1162);
or U2311 (N_2311,In_362,In_1388);
and U2312 (N_2312,In_8,In_1398);
and U2313 (N_2313,In_386,In_256);
or U2314 (N_2314,In_964,In_1362);
nand U2315 (N_2315,In_1092,In_345);
nand U2316 (N_2316,In_907,In_1187);
nand U2317 (N_2317,In_1251,In_30);
and U2318 (N_2318,In_816,In_113);
or U2319 (N_2319,In_431,In_193);
or U2320 (N_2320,In_550,In_1247);
nor U2321 (N_2321,In_133,In_1024);
nand U2322 (N_2322,In_234,In_1200);
nand U2323 (N_2323,In_206,In_914);
nand U2324 (N_2324,In_997,In_505);
nor U2325 (N_2325,In_932,In_170);
or U2326 (N_2326,In_34,In_640);
xnor U2327 (N_2327,In_141,In_188);
and U2328 (N_2328,In_877,In_847);
and U2329 (N_2329,In_912,In_1443);
nor U2330 (N_2330,In_23,In_1255);
nor U2331 (N_2331,In_1314,In_1013);
or U2332 (N_2332,In_1439,In_377);
or U2333 (N_2333,In_1186,In_647);
nand U2334 (N_2334,In_790,In_1028);
and U2335 (N_2335,In_744,In_1251);
and U2336 (N_2336,In_1359,In_1022);
nand U2337 (N_2337,In_1351,In_1102);
or U2338 (N_2338,In_40,In_1309);
nor U2339 (N_2339,In_598,In_27);
or U2340 (N_2340,In_252,In_1479);
and U2341 (N_2341,In_143,In_912);
nand U2342 (N_2342,In_1251,In_1260);
nand U2343 (N_2343,In_992,In_52);
nor U2344 (N_2344,In_910,In_819);
nand U2345 (N_2345,In_970,In_406);
and U2346 (N_2346,In_1058,In_995);
or U2347 (N_2347,In_26,In_1366);
and U2348 (N_2348,In_1484,In_1175);
or U2349 (N_2349,In_1074,In_581);
nor U2350 (N_2350,In_1463,In_1024);
or U2351 (N_2351,In_660,In_517);
nand U2352 (N_2352,In_290,In_620);
nand U2353 (N_2353,In_55,In_836);
nor U2354 (N_2354,In_774,In_1076);
nor U2355 (N_2355,In_392,In_1444);
or U2356 (N_2356,In_256,In_1200);
or U2357 (N_2357,In_254,In_921);
nand U2358 (N_2358,In_436,In_152);
xnor U2359 (N_2359,In_1244,In_368);
nor U2360 (N_2360,In_900,In_1322);
or U2361 (N_2361,In_383,In_958);
or U2362 (N_2362,In_108,In_686);
nand U2363 (N_2363,In_996,In_806);
or U2364 (N_2364,In_213,In_697);
nand U2365 (N_2365,In_824,In_1444);
nor U2366 (N_2366,In_115,In_24);
and U2367 (N_2367,In_831,In_218);
nor U2368 (N_2368,In_245,In_938);
and U2369 (N_2369,In_290,In_219);
xnor U2370 (N_2370,In_1236,In_766);
nand U2371 (N_2371,In_361,In_1362);
nand U2372 (N_2372,In_1252,In_1223);
and U2373 (N_2373,In_303,In_1283);
nor U2374 (N_2374,In_1434,In_1279);
nand U2375 (N_2375,In_1457,In_1093);
and U2376 (N_2376,In_570,In_829);
nand U2377 (N_2377,In_1492,In_1225);
and U2378 (N_2378,In_165,In_933);
nand U2379 (N_2379,In_78,In_179);
or U2380 (N_2380,In_715,In_1005);
and U2381 (N_2381,In_895,In_644);
nand U2382 (N_2382,In_466,In_678);
nor U2383 (N_2383,In_99,In_1314);
nor U2384 (N_2384,In_444,In_1409);
or U2385 (N_2385,In_1164,In_242);
nor U2386 (N_2386,In_228,In_1343);
nand U2387 (N_2387,In_647,In_805);
and U2388 (N_2388,In_571,In_445);
xnor U2389 (N_2389,In_1241,In_1145);
nor U2390 (N_2390,In_1104,In_1196);
nand U2391 (N_2391,In_221,In_387);
and U2392 (N_2392,In_327,In_536);
nor U2393 (N_2393,In_539,In_1264);
nor U2394 (N_2394,In_121,In_1116);
nand U2395 (N_2395,In_484,In_707);
nor U2396 (N_2396,In_612,In_741);
or U2397 (N_2397,In_342,In_573);
nor U2398 (N_2398,In_1433,In_89);
or U2399 (N_2399,In_210,In_350);
nand U2400 (N_2400,In_175,In_1031);
and U2401 (N_2401,In_4,In_1232);
and U2402 (N_2402,In_891,In_1221);
nand U2403 (N_2403,In_179,In_553);
nor U2404 (N_2404,In_1340,In_616);
nand U2405 (N_2405,In_1181,In_1473);
nor U2406 (N_2406,In_1318,In_1209);
nor U2407 (N_2407,In_112,In_970);
nor U2408 (N_2408,In_90,In_796);
nand U2409 (N_2409,In_265,In_977);
or U2410 (N_2410,In_1131,In_1172);
xor U2411 (N_2411,In_1466,In_992);
nor U2412 (N_2412,In_54,In_1445);
nor U2413 (N_2413,In_862,In_1323);
or U2414 (N_2414,In_302,In_1099);
and U2415 (N_2415,In_63,In_928);
nand U2416 (N_2416,In_1164,In_1298);
or U2417 (N_2417,In_445,In_644);
nand U2418 (N_2418,In_994,In_1018);
and U2419 (N_2419,In_1494,In_1456);
nand U2420 (N_2420,In_1320,In_1157);
or U2421 (N_2421,In_1207,In_363);
nor U2422 (N_2422,In_1271,In_468);
nor U2423 (N_2423,In_263,In_1199);
nor U2424 (N_2424,In_1009,In_1477);
nor U2425 (N_2425,In_145,In_17);
and U2426 (N_2426,In_1132,In_495);
or U2427 (N_2427,In_1295,In_897);
nand U2428 (N_2428,In_285,In_732);
nand U2429 (N_2429,In_143,In_342);
nor U2430 (N_2430,In_485,In_619);
or U2431 (N_2431,In_1077,In_1010);
or U2432 (N_2432,In_1260,In_887);
and U2433 (N_2433,In_1497,In_739);
or U2434 (N_2434,In_1068,In_1214);
nand U2435 (N_2435,In_234,In_926);
nand U2436 (N_2436,In_1026,In_380);
nor U2437 (N_2437,In_973,In_238);
nand U2438 (N_2438,In_492,In_227);
or U2439 (N_2439,In_710,In_785);
nor U2440 (N_2440,In_1026,In_526);
and U2441 (N_2441,In_666,In_1287);
and U2442 (N_2442,In_1000,In_878);
nor U2443 (N_2443,In_1256,In_400);
nand U2444 (N_2444,In_269,In_1262);
and U2445 (N_2445,In_1100,In_32);
nor U2446 (N_2446,In_237,In_4);
or U2447 (N_2447,In_70,In_1428);
or U2448 (N_2448,In_244,In_1221);
or U2449 (N_2449,In_1442,In_766);
nand U2450 (N_2450,In_616,In_698);
nand U2451 (N_2451,In_1167,In_919);
nand U2452 (N_2452,In_449,In_929);
or U2453 (N_2453,In_209,In_237);
nor U2454 (N_2454,In_526,In_1349);
nor U2455 (N_2455,In_214,In_675);
and U2456 (N_2456,In_239,In_642);
nor U2457 (N_2457,In_185,In_158);
nand U2458 (N_2458,In_549,In_744);
or U2459 (N_2459,In_8,In_1285);
nor U2460 (N_2460,In_1284,In_509);
nand U2461 (N_2461,In_108,In_320);
or U2462 (N_2462,In_131,In_592);
or U2463 (N_2463,In_52,In_92);
and U2464 (N_2464,In_1491,In_849);
nand U2465 (N_2465,In_629,In_921);
nor U2466 (N_2466,In_221,In_352);
nor U2467 (N_2467,In_251,In_115);
and U2468 (N_2468,In_429,In_630);
nand U2469 (N_2469,In_990,In_215);
nand U2470 (N_2470,In_831,In_1431);
nand U2471 (N_2471,In_788,In_77);
nand U2472 (N_2472,In_262,In_804);
nand U2473 (N_2473,In_282,In_702);
or U2474 (N_2474,In_273,In_158);
and U2475 (N_2475,In_1274,In_1220);
or U2476 (N_2476,In_226,In_779);
nand U2477 (N_2477,In_275,In_712);
and U2478 (N_2478,In_362,In_1471);
or U2479 (N_2479,In_135,In_926);
and U2480 (N_2480,In_236,In_381);
nand U2481 (N_2481,In_266,In_625);
nor U2482 (N_2482,In_1288,In_252);
nor U2483 (N_2483,In_284,In_1008);
and U2484 (N_2484,In_93,In_1224);
nand U2485 (N_2485,In_422,In_967);
nor U2486 (N_2486,In_1174,In_1393);
nor U2487 (N_2487,In_944,In_1348);
or U2488 (N_2488,In_453,In_688);
nand U2489 (N_2489,In_328,In_1135);
nand U2490 (N_2490,In_851,In_1427);
nand U2491 (N_2491,In_1403,In_636);
nand U2492 (N_2492,In_305,In_1262);
nand U2493 (N_2493,In_1240,In_376);
nand U2494 (N_2494,In_1384,In_999);
and U2495 (N_2495,In_65,In_978);
nand U2496 (N_2496,In_264,In_885);
nor U2497 (N_2497,In_1238,In_183);
xor U2498 (N_2498,In_929,In_1108);
or U2499 (N_2499,In_1066,In_784);
nand U2500 (N_2500,In_280,In_1368);
or U2501 (N_2501,In_528,In_1067);
and U2502 (N_2502,In_248,In_397);
and U2503 (N_2503,In_1468,In_1242);
or U2504 (N_2504,In_86,In_934);
nor U2505 (N_2505,In_102,In_383);
or U2506 (N_2506,In_918,In_504);
nand U2507 (N_2507,In_1132,In_1231);
and U2508 (N_2508,In_1158,In_94);
or U2509 (N_2509,In_685,In_1271);
or U2510 (N_2510,In_1131,In_69);
or U2511 (N_2511,In_438,In_284);
nand U2512 (N_2512,In_429,In_1169);
and U2513 (N_2513,In_440,In_1149);
nand U2514 (N_2514,In_463,In_830);
nor U2515 (N_2515,In_957,In_1445);
nand U2516 (N_2516,In_1178,In_200);
and U2517 (N_2517,In_682,In_452);
nor U2518 (N_2518,In_1185,In_1458);
and U2519 (N_2519,In_735,In_928);
nor U2520 (N_2520,In_742,In_782);
and U2521 (N_2521,In_79,In_187);
nor U2522 (N_2522,In_1427,In_1493);
or U2523 (N_2523,In_1309,In_1455);
nand U2524 (N_2524,In_1238,In_545);
and U2525 (N_2525,In_462,In_63);
or U2526 (N_2526,In_145,In_104);
and U2527 (N_2527,In_133,In_94);
nor U2528 (N_2528,In_1323,In_1289);
or U2529 (N_2529,In_1000,In_886);
nor U2530 (N_2530,In_727,In_1464);
nand U2531 (N_2531,In_170,In_1200);
or U2532 (N_2532,In_1093,In_684);
nor U2533 (N_2533,In_935,In_1285);
nand U2534 (N_2534,In_507,In_1271);
nand U2535 (N_2535,In_586,In_990);
nor U2536 (N_2536,In_297,In_558);
nand U2537 (N_2537,In_966,In_1104);
nand U2538 (N_2538,In_1298,In_687);
nand U2539 (N_2539,In_1409,In_437);
nor U2540 (N_2540,In_1356,In_1233);
and U2541 (N_2541,In_1432,In_1114);
nor U2542 (N_2542,In_395,In_806);
and U2543 (N_2543,In_560,In_1388);
or U2544 (N_2544,In_1057,In_421);
or U2545 (N_2545,In_1279,In_1246);
nand U2546 (N_2546,In_1483,In_350);
nand U2547 (N_2547,In_31,In_1348);
nand U2548 (N_2548,In_512,In_1270);
nand U2549 (N_2549,In_296,In_1054);
nor U2550 (N_2550,In_1157,In_762);
nor U2551 (N_2551,In_305,In_588);
nor U2552 (N_2552,In_490,In_1490);
or U2553 (N_2553,In_1313,In_198);
or U2554 (N_2554,In_547,In_785);
and U2555 (N_2555,In_1243,In_1131);
nor U2556 (N_2556,In_270,In_250);
nor U2557 (N_2557,In_480,In_418);
or U2558 (N_2558,In_1208,In_25);
nor U2559 (N_2559,In_1200,In_335);
nand U2560 (N_2560,In_777,In_1047);
or U2561 (N_2561,In_812,In_1161);
or U2562 (N_2562,In_1498,In_1366);
nand U2563 (N_2563,In_710,In_1081);
and U2564 (N_2564,In_1362,In_796);
or U2565 (N_2565,In_677,In_732);
and U2566 (N_2566,In_149,In_1238);
and U2567 (N_2567,In_1079,In_1206);
nand U2568 (N_2568,In_978,In_379);
nor U2569 (N_2569,In_1088,In_1497);
or U2570 (N_2570,In_1089,In_1359);
nor U2571 (N_2571,In_268,In_1471);
or U2572 (N_2572,In_466,In_488);
nor U2573 (N_2573,In_254,In_427);
and U2574 (N_2574,In_812,In_1271);
xor U2575 (N_2575,In_1308,In_1191);
nor U2576 (N_2576,In_1466,In_26);
nand U2577 (N_2577,In_1103,In_341);
or U2578 (N_2578,In_363,In_1085);
or U2579 (N_2579,In_640,In_203);
and U2580 (N_2580,In_861,In_942);
or U2581 (N_2581,In_874,In_145);
and U2582 (N_2582,In_713,In_317);
nor U2583 (N_2583,In_1231,In_1055);
nand U2584 (N_2584,In_1040,In_634);
nand U2585 (N_2585,In_362,In_343);
nor U2586 (N_2586,In_1054,In_1168);
nand U2587 (N_2587,In_1440,In_485);
nand U2588 (N_2588,In_422,In_988);
nor U2589 (N_2589,In_1074,In_299);
nor U2590 (N_2590,In_659,In_831);
or U2591 (N_2591,In_440,In_391);
or U2592 (N_2592,In_1067,In_584);
nor U2593 (N_2593,In_991,In_622);
nand U2594 (N_2594,In_284,In_1395);
nand U2595 (N_2595,In_121,In_383);
xor U2596 (N_2596,In_881,In_87);
nor U2597 (N_2597,In_1174,In_859);
and U2598 (N_2598,In_319,In_537);
nand U2599 (N_2599,In_752,In_582);
nor U2600 (N_2600,In_312,In_73);
or U2601 (N_2601,In_1421,In_1467);
or U2602 (N_2602,In_422,In_907);
xnor U2603 (N_2603,In_1124,In_1327);
nor U2604 (N_2604,In_259,In_178);
nor U2605 (N_2605,In_511,In_1164);
and U2606 (N_2606,In_241,In_1418);
nor U2607 (N_2607,In_897,In_106);
nor U2608 (N_2608,In_902,In_1373);
or U2609 (N_2609,In_472,In_1085);
or U2610 (N_2610,In_1059,In_636);
or U2611 (N_2611,In_1477,In_1189);
and U2612 (N_2612,In_131,In_1048);
nor U2613 (N_2613,In_1031,In_642);
and U2614 (N_2614,In_1325,In_1338);
nor U2615 (N_2615,In_1472,In_503);
and U2616 (N_2616,In_105,In_239);
or U2617 (N_2617,In_1369,In_1446);
or U2618 (N_2618,In_355,In_1358);
nand U2619 (N_2619,In_442,In_1017);
and U2620 (N_2620,In_1046,In_162);
nor U2621 (N_2621,In_1170,In_67);
and U2622 (N_2622,In_1270,In_1403);
nor U2623 (N_2623,In_265,In_165);
nand U2624 (N_2624,In_1331,In_1373);
or U2625 (N_2625,In_149,In_814);
and U2626 (N_2626,In_1005,In_937);
nand U2627 (N_2627,In_523,In_312);
nand U2628 (N_2628,In_154,In_169);
or U2629 (N_2629,In_826,In_489);
nor U2630 (N_2630,In_1227,In_144);
nor U2631 (N_2631,In_922,In_1039);
nor U2632 (N_2632,In_30,In_1189);
or U2633 (N_2633,In_889,In_136);
or U2634 (N_2634,In_384,In_1294);
nor U2635 (N_2635,In_862,In_1001);
nand U2636 (N_2636,In_518,In_806);
and U2637 (N_2637,In_321,In_1198);
and U2638 (N_2638,In_716,In_1493);
nor U2639 (N_2639,In_1391,In_453);
nor U2640 (N_2640,In_251,In_734);
nor U2641 (N_2641,In_1205,In_1411);
and U2642 (N_2642,In_613,In_1258);
and U2643 (N_2643,In_521,In_240);
nor U2644 (N_2644,In_1031,In_1278);
and U2645 (N_2645,In_933,In_994);
xnor U2646 (N_2646,In_484,In_1126);
nor U2647 (N_2647,In_1049,In_1473);
and U2648 (N_2648,In_473,In_89);
and U2649 (N_2649,In_303,In_881);
and U2650 (N_2650,In_1299,In_408);
nand U2651 (N_2651,In_1271,In_1497);
nor U2652 (N_2652,In_1454,In_1212);
nand U2653 (N_2653,In_1327,In_766);
or U2654 (N_2654,In_542,In_240);
and U2655 (N_2655,In_1268,In_450);
and U2656 (N_2656,In_657,In_907);
or U2657 (N_2657,In_743,In_174);
nand U2658 (N_2658,In_871,In_910);
nor U2659 (N_2659,In_1272,In_381);
xor U2660 (N_2660,In_1448,In_66);
and U2661 (N_2661,In_47,In_287);
and U2662 (N_2662,In_424,In_699);
nand U2663 (N_2663,In_886,In_869);
and U2664 (N_2664,In_936,In_420);
or U2665 (N_2665,In_267,In_1309);
or U2666 (N_2666,In_209,In_413);
or U2667 (N_2667,In_224,In_1459);
nor U2668 (N_2668,In_359,In_1458);
or U2669 (N_2669,In_620,In_315);
nand U2670 (N_2670,In_636,In_1378);
nand U2671 (N_2671,In_12,In_240);
nand U2672 (N_2672,In_945,In_386);
or U2673 (N_2673,In_21,In_685);
and U2674 (N_2674,In_1058,In_341);
and U2675 (N_2675,In_695,In_486);
nor U2676 (N_2676,In_1146,In_518);
nand U2677 (N_2677,In_1063,In_6);
nand U2678 (N_2678,In_1415,In_335);
and U2679 (N_2679,In_639,In_660);
or U2680 (N_2680,In_807,In_352);
nand U2681 (N_2681,In_1492,In_1056);
and U2682 (N_2682,In_756,In_471);
nand U2683 (N_2683,In_318,In_1398);
nor U2684 (N_2684,In_497,In_125);
nand U2685 (N_2685,In_370,In_1202);
nor U2686 (N_2686,In_1272,In_132);
nand U2687 (N_2687,In_339,In_917);
or U2688 (N_2688,In_847,In_639);
nand U2689 (N_2689,In_1182,In_712);
nor U2690 (N_2690,In_1338,In_643);
or U2691 (N_2691,In_619,In_86);
or U2692 (N_2692,In_387,In_779);
nand U2693 (N_2693,In_817,In_1476);
nor U2694 (N_2694,In_275,In_264);
and U2695 (N_2695,In_160,In_534);
nor U2696 (N_2696,In_1305,In_405);
and U2697 (N_2697,In_271,In_955);
nand U2698 (N_2698,In_1168,In_216);
and U2699 (N_2699,In_1477,In_174);
nor U2700 (N_2700,In_14,In_1392);
and U2701 (N_2701,In_189,In_633);
and U2702 (N_2702,In_223,In_0);
nand U2703 (N_2703,In_1087,In_1080);
nand U2704 (N_2704,In_103,In_561);
or U2705 (N_2705,In_61,In_679);
nand U2706 (N_2706,In_857,In_337);
and U2707 (N_2707,In_613,In_679);
or U2708 (N_2708,In_50,In_277);
or U2709 (N_2709,In_658,In_1428);
nor U2710 (N_2710,In_1311,In_1416);
nor U2711 (N_2711,In_42,In_449);
xnor U2712 (N_2712,In_1308,In_849);
and U2713 (N_2713,In_236,In_336);
xor U2714 (N_2714,In_1296,In_1109);
and U2715 (N_2715,In_725,In_1321);
and U2716 (N_2716,In_339,In_1447);
nor U2717 (N_2717,In_515,In_461);
nand U2718 (N_2718,In_1264,In_1049);
or U2719 (N_2719,In_287,In_870);
or U2720 (N_2720,In_760,In_529);
nand U2721 (N_2721,In_216,In_1467);
nand U2722 (N_2722,In_1332,In_304);
and U2723 (N_2723,In_1390,In_1339);
and U2724 (N_2724,In_449,In_1137);
nand U2725 (N_2725,In_1289,In_287);
nand U2726 (N_2726,In_263,In_235);
or U2727 (N_2727,In_1273,In_1103);
nand U2728 (N_2728,In_1399,In_35);
nor U2729 (N_2729,In_444,In_1063);
nand U2730 (N_2730,In_504,In_682);
or U2731 (N_2731,In_332,In_279);
xor U2732 (N_2732,In_57,In_1297);
nor U2733 (N_2733,In_1013,In_153);
nor U2734 (N_2734,In_1020,In_1494);
nand U2735 (N_2735,In_572,In_246);
or U2736 (N_2736,In_309,In_645);
nand U2737 (N_2737,In_1387,In_913);
or U2738 (N_2738,In_681,In_1483);
nor U2739 (N_2739,In_994,In_373);
nand U2740 (N_2740,In_958,In_1015);
nand U2741 (N_2741,In_951,In_890);
nand U2742 (N_2742,In_1465,In_290);
and U2743 (N_2743,In_667,In_1429);
and U2744 (N_2744,In_911,In_1360);
nand U2745 (N_2745,In_741,In_572);
nand U2746 (N_2746,In_821,In_1145);
nor U2747 (N_2747,In_1132,In_656);
and U2748 (N_2748,In_301,In_1463);
nand U2749 (N_2749,In_1148,In_1488);
nor U2750 (N_2750,In_1100,In_655);
nand U2751 (N_2751,In_448,In_310);
or U2752 (N_2752,In_910,In_406);
xnor U2753 (N_2753,In_611,In_881);
nand U2754 (N_2754,In_142,In_582);
nand U2755 (N_2755,In_752,In_0);
and U2756 (N_2756,In_188,In_663);
nor U2757 (N_2757,In_419,In_967);
nand U2758 (N_2758,In_735,In_348);
or U2759 (N_2759,In_1061,In_923);
nand U2760 (N_2760,In_312,In_645);
nand U2761 (N_2761,In_1392,In_31);
nand U2762 (N_2762,In_695,In_234);
nor U2763 (N_2763,In_947,In_91);
nand U2764 (N_2764,In_839,In_112);
nand U2765 (N_2765,In_78,In_425);
nand U2766 (N_2766,In_157,In_559);
nor U2767 (N_2767,In_524,In_958);
nor U2768 (N_2768,In_1386,In_388);
nor U2769 (N_2769,In_195,In_482);
or U2770 (N_2770,In_1240,In_282);
and U2771 (N_2771,In_508,In_145);
or U2772 (N_2772,In_1020,In_829);
and U2773 (N_2773,In_700,In_1100);
and U2774 (N_2774,In_498,In_928);
and U2775 (N_2775,In_872,In_474);
or U2776 (N_2776,In_1480,In_408);
nand U2777 (N_2777,In_308,In_173);
and U2778 (N_2778,In_507,In_1402);
nor U2779 (N_2779,In_15,In_97);
and U2780 (N_2780,In_1095,In_1175);
and U2781 (N_2781,In_420,In_1140);
nand U2782 (N_2782,In_775,In_132);
nor U2783 (N_2783,In_447,In_89);
nand U2784 (N_2784,In_847,In_693);
and U2785 (N_2785,In_448,In_178);
nand U2786 (N_2786,In_609,In_375);
nand U2787 (N_2787,In_793,In_493);
or U2788 (N_2788,In_460,In_1333);
or U2789 (N_2789,In_1391,In_827);
nor U2790 (N_2790,In_1297,In_407);
or U2791 (N_2791,In_1001,In_1164);
and U2792 (N_2792,In_275,In_1143);
and U2793 (N_2793,In_929,In_1352);
or U2794 (N_2794,In_493,In_964);
or U2795 (N_2795,In_135,In_318);
or U2796 (N_2796,In_319,In_937);
nand U2797 (N_2797,In_387,In_164);
nor U2798 (N_2798,In_338,In_32);
or U2799 (N_2799,In_565,In_820);
nor U2800 (N_2800,In_161,In_866);
nor U2801 (N_2801,In_1122,In_537);
nor U2802 (N_2802,In_633,In_445);
and U2803 (N_2803,In_808,In_880);
nor U2804 (N_2804,In_1203,In_1234);
or U2805 (N_2805,In_1228,In_162);
or U2806 (N_2806,In_518,In_256);
nor U2807 (N_2807,In_353,In_540);
and U2808 (N_2808,In_551,In_642);
and U2809 (N_2809,In_1177,In_685);
or U2810 (N_2810,In_391,In_501);
and U2811 (N_2811,In_649,In_937);
nand U2812 (N_2812,In_1283,In_686);
and U2813 (N_2813,In_1136,In_378);
or U2814 (N_2814,In_220,In_791);
nand U2815 (N_2815,In_329,In_1213);
and U2816 (N_2816,In_1483,In_272);
nand U2817 (N_2817,In_1308,In_1388);
nor U2818 (N_2818,In_1093,In_598);
or U2819 (N_2819,In_1258,In_1319);
nand U2820 (N_2820,In_1337,In_1434);
nand U2821 (N_2821,In_573,In_689);
nand U2822 (N_2822,In_463,In_344);
or U2823 (N_2823,In_350,In_700);
or U2824 (N_2824,In_416,In_962);
nand U2825 (N_2825,In_88,In_1231);
nor U2826 (N_2826,In_906,In_682);
and U2827 (N_2827,In_1114,In_854);
nand U2828 (N_2828,In_151,In_322);
nand U2829 (N_2829,In_984,In_239);
nand U2830 (N_2830,In_1103,In_1073);
and U2831 (N_2831,In_450,In_30);
and U2832 (N_2832,In_679,In_618);
and U2833 (N_2833,In_474,In_1218);
or U2834 (N_2834,In_922,In_322);
nor U2835 (N_2835,In_1123,In_521);
or U2836 (N_2836,In_602,In_405);
nor U2837 (N_2837,In_280,In_38);
or U2838 (N_2838,In_12,In_3);
nand U2839 (N_2839,In_311,In_547);
xor U2840 (N_2840,In_1153,In_1039);
nor U2841 (N_2841,In_1232,In_681);
nand U2842 (N_2842,In_1427,In_1254);
nand U2843 (N_2843,In_491,In_926);
and U2844 (N_2844,In_659,In_605);
and U2845 (N_2845,In_1313,In_205);
nand U2846 (N_2846,In_655,In_681);
nand U2847 (N_2847,In_45,In_692);
or U2848 (N_2848,In_941,In_990);
nand U2849 (N_2849,In_1342,In_1109);
nor U2850 (N_2850,In_222,In_1466);
and U2851 (N_2851,In_148,In_1157);
nor U2852 (N_2852,In_269,In_1208);
nand U2853 (N_2853,In_83,In_1464);
and U2854 (N_2854,In_199,In_748);
nand U2855 (N_2855,In_705,In_1254);
nor U2856 (N_2856,In_385,In_330);
nand U2857 (N_2857,In_1007,In_446);
nand U2858 (N_2858,In_1038,In_1207);
or U2859 (N_2859,In_781,In_1016);
or U2860 (N_2860,In_1171,In_1430);
and U2861 (N_2861,In_679,In_1466);
and U2862 (N_2862,In_272,In_1423);
nand U2863 (N_2863,In_976,In_1437);
nand U2864 (N_2864,In_1287,In_239);
nand U2865 (N_2865,In_763,In_715);
or U2866 (N_2866,In_969,In_799);
or U2867 (N_2867,In_1285,In_400);
or U2868 (N_2868,In_1092,In_356);
or U2869 (N_2869,In_425,In_1413);
and U2870 (N_2870,In_1066,In_528);
nor U2871 (N_2871,In_536,In_130);
or U2872 (N_2872,In_938,In_1353);
nor U2873 (N_2873,In_733,In_587);
nor U2874 (N_2874,In_669,In_1174);
nand U2875 (N_2875,In_1492,In_928);
nand U2876 (N_2876,In_1313,In_1232);
nand U2877 (N_2877,In_1402,In_916);
and U2878 (N_2878,In_1407,In_1154);
nor U2879 (N_2879,In_1496,In_1168);
nor U2880 (N_2880,In_80,In_47);
nor U2881 (N_2881,In_838,In_1230);
or U2882 (N_2882,In_589,In_347);
nor U2883 (N_2883,In_201,In_1177);
or U2884 (N_2884,In_1133,In_569);
nand U2885 (N_2885,In_1270,In_306);
nand U2886 (N_2886,In_998,In_1406);
and U2887 (N_2887,In_1023,In_819);
nand U2888 (N_2888,In_705,In_951);
nor U2889 (N_2889,In_976,In_64);
nand U2890 (N_2890,In_661,In_626);
nor U2891 (N_2891,In_754,In_571);
nor U2892 (N_2892,In_1213,In_620);
or U2893 (N_2893,In_1308,In_688);
nor U2894 (N_2894,In_1472,In_976);
and U2895 (N_2895,In_488,In_464);
or U2896 (N_2896,In_92,In_928);
or U2897 (N_2897,In_1394,In_726);
and U2898 (N_2898,In_840,In_174);
nor U2899 (N_2899,In_550,In_335);
nor U2900 (N_2900,In_199,In_405);
nand U2901 (N_2901,In_1245,In_682);
nor U2902 (N_2902,In_912,In_778);
and U2903 (N_2903,In_1404,In_1164);
nor U2904 (N_2904,In_1375,In_793);
and U2905 (N_2905,In_876,In_772);
nand U2906 (N_2906,In_772,In_283);
nor U2907 (N_2907,In_815,In_598);
and U2908 (N_2908,In_1248,In_426);
or U2909 (N_2909,In_170,In_1096);
nor U2910 (N_2910,In_1078,In_1337);
nor U2911 (N_2911,In_563,In_298);
nand U2912 (N_2912,In_376,In_789);
and U2913 (N_2913,In_1092,In_1445);
and U2914 (N_2914,In_828,In_904);
nor U2915 (N_2915,In_377,In_832);
or U2916 (N_2916,In_1407,In_598);
and U2917 (N_2917,In_241,In_1414);
and U2918 (N_2918,In_749,In_974);
nand U2919 (N_2919,In_1149,In_1301);
nor U2920 (N_2920,In_1262,In_52);
nor U2921 (N_2921,In_545,In_502);
nand U2922 (N_2922,In_1216,In_402);
or U2923 (N_2923,In_336,In_106);
or U2924 (N_2924,In_354,In_875);
and U2925 (N_2925,In_160,In_1152);
nor U2926 (N_2926,In_1477,In_411);
and U2927 (N_2927,In_1076,In_995);
nor U2928 (N_2928,In_1301,In_176);
nand U2929 (N_2929,In_1250,In_1071);
nand U2930 (N_2930,In_889,In_407);
or U2931 (N_2931,In_777,In_354);
nor U2932 (N_2932,In_899,In_197);
nor U2933 (N_2933,In_1334,In_1026);
and U2934 (N_2934,In_414,In_1476);
or U2935 (N_2935,In_491,In_1426);
and U2936 (N_2936,In_549,In_701);
or U2937 (N_2937,In_75,In_1156);
nor U2938 (N_2938,In_214,In_44);
nand U2939 (N_2939,In_424,In_254);
and U2940 (N_2940,In_780,In_1481);
nor U2941 (N_2941,In_441,In_133);
and U2942 (N_2942,In_937,In_304);
and U2943 (N_2943,In_304,In_1120);
or U2944 (N_2944,In_1167,In_75);
nand U2945 (N_2945,In_162,In_849);
and U2946 (N_2946,In_1237,In_1381);
nor U2947 (N_2947,In_1185,In_657);
and U2948 (N_2948,In_915,In_448);
nor U2949 (N_2949,In_127,In_46);
nor U2950 (N_2950,In_1080,In_1242);
or U2951 (N_2951,In_672,In_1139);
or U2952 (N_2952,In_14,In_268);
or U2953 (N_2953,In_376,In_1499);
or U2954 (N_2954,In_1160,In_546);
nand U2955 (N_2955,In_1051,In_659);
nand U2956 (N_2956,In_719,In_727);
nor U2957 (N_2957,In_452,In_991);
nand U2958 (N_2958,In_655,In_1471);
or U2959 (N_2959,In_988,In_741);
nand U2960 (N_2960,In_73,In_1446);
nor U2961 (N_2961,In_1,In_1103);
or U2962 (N_2962,In_1086,In_1079);
nand U2963 (N_2963,In_957,In_305);
xor U2964 (N_2964,In_58,In_560);
nand U2965 (N_2965,In_542,In_653);
nor U2966 (N_2966,In_1405,In_1221);
nand U2967 (N_2967,In_694,In_263);
or U2968 (N_2968,In_36,In_1140);
nor U2969 (N_2969,In_124,In_103);
or U2970 (N_2970,In_153,In_1281);
or U2971 (N_2971,In_513,In_94);
nand U2972 (N_2972,In_827,In_783);
nor U2973 (N_2973,In_969,In_390);
or U2974 (N_2974,In_641,In_1425);
nor U2975 (N_2975,In_443,In_2);
and U2976 (N_2976,In_1259,In_1054);
or U2977 (N_2977,In_60,In_25);
nor U2978 (N_2978,In_768,In_1141);
or U2979 (N_2979,In_1244,In_1093);
and U2980 (N_2980,In_1162,In_806);
or U2981 (N_2981,In_135,In_183);
and U2982 (N_2982,In_1489,In_881);
nand U2983 (N_2983,In_68,In_1148);
or U2984 (N_2984,In_535,In_852);
nand U2985 (N_2985,In_1310,In_1458);
nor U2986 (N_2986,In_125,In_1061);
and U2987 (N_2987,In_1369,In_703);
and U2988 (N_2988,In_836,In_155);
or U2989 (N_2989,In_214,In_368);
and U2990 (N_2990,In_1354,In_574);
and U2991 (N_2991,In_516,In_513);
or U2992 (N_2992,In_858,In_742);
nor U2993 (N_2993,In_1353,In_894);
and U2994 (N_2994,In_271,In_864);
or U2995 (N_2995,In_512,In_1242);
and U2996 (N_2996,In_755,In_205);
and U2997 (N_2997,In_1040,In_31);
nand U2998 (N_2998,In_1411,In_586);
or U2999 (N_2999,In_1472,In_1493);
and U3000 (N_3000,In_809,In_624);
or U3001 (N_3001,In_939,In_811);
or U3002 (N_3002,In_1399,In_238);
nor U3003 (N_3003,In_387,In_1126);
nand U3004 (N_3004,In_151,In_1173);
nand U3005 (N_3005,In_393,In_111);
nor U3006 (N_3006,In_452,In_184);
or U3007 (N_3007,In_802,In_1427);
and U3008 (N_3008,In_1023,In_63);
nor U3009 (N_3009,In_1118,In_1042);
nor U3010 (N_3010,In_777,In_708);
nor U3011 (N_3011,In_474,In_701);
nand U3012 (N_3012,In_924,In_1331);
and U3013 (N_3013,In_1363,In_535);
or U3014 (N_3014,In_1369,In_715);
or U3015 (N_3015,In_666,In_1240);
or U3016 (N_3016,In_129,In_351);
nor U3017 (N_3017,In_1190,In_60);
and U3018 (N_3018,In_615,In_274);
or U3019 (N_3019,In_750,In_1015);
and U3020 (N_3020,In_809,In_304);
nor U3021 (N_3021,In_971,In_683);
and U3022 (N_3022,In_835,In_1220);
or U3023 (N_3023,In_1105,In_347);
nor U3024 (N_3024,In_86,In_618);
nand U3025 (N_3025,In_1214,In_688);
nand U3026 (N_3026,In_847,In_308);
nor U3027 (N_3027,In_431,In_921);
and U3028 (N_3028,In_1157,In_1490);
or U3029 (N_3029,In_1222,In_928);
or U3030 (N_3030,In_779,In_659);
or U3031 (N_3031,In_1055,In_988);
nor U3032 (N_3032,In_255,In_1345);
nor U3033 (N_3033,In_868,In_706);
or U3034 (N_3034,In_1186,In_103);
nand U3035 (N_3035,In_1075,In_940);
nand U3036 (N_3036,In_903,In_1007);
nand U3037 (N_3037,In_251,In_1163);
or U3038 (N_3038,In_351,In_1194);
nor U3039 (N_3039,In_4,In_1052);
nand U3040 (N_3040,In_1303,In_200);
and U3041 (N_3041,In_429,In_953);
and U3042 (N_3042,In_310,In_312);
nand U3043 (N_3043,In_290,In_418);
or U3044 (N_3044,In_809,In_1169);
or U3045 (N_3045,In_54,In_1070);
or U3046 (N_3046,In_1310,In_389);
or U3047 (N_3047,In_1288,In_972);
nand U3048 (N_3048,In_282,In_766);
and U3049 (N_3049,In_724,In_1203);
or U3050 (N_3050,In_333,In_1371);
nor U3051 (N_3051,In_490,In_92);
or U3052 (N_3052,In_297,In_401);
nand U3053 (N_3053,In_1455,In_604);
nand U3054 (N_3054,In_182,In_1384);
or U3055 (N_3055,In_285,In_1026);
nand U3056 (N_3056,In_1000,In_163);
nand U3057 (N_3057,In_108,In_1017);
nor U3058 (N_3058,In_903,In_1323);
and U3059 (N_3059,In_295,In_1067);
or U3060 (N_3060,In_204,In_1299);
and U3061 (N_3061,In_646,In_295);
and U3062 (N_3062,In_982,In_25);
and U3063 (N_3063,In_921,In_1309);
and U3064 (N_3064,In_41,In_354);
nand U3065 (N_3065,In_179,In_428);
nor U3066 (N_3066,In_1127,In_134);
and U3067 (N_3067,In_1108,In_859);
xor U3068 (N_3068,In_28,In_1191);
nor U3069 (N_3069,In_397,In_351);
nor U3070 (N_3070,In_499,In_1376);
nand U3071 (N_3071,In_346,In_749);
nand U3072 (N_3072,In_312,In_636);
nand U3073 (N_3073,In_1289,In_32);
nand U3074 (N_3074,In_1446,In_481);
and U3075 (N_3075,In_474,In_1499);
and U3076 (N_3076,In_441,In_1318);
and U3077 (N_3077,In_146,In_726);
or U3078 (N_3078,In_874,In_1091);
and U3079 (N_3079,In_1023,In_715);
nand U3080 (N_3080,In_860,In_1453);
nor U3081 (N_3081,In_172,In_929);
or U3082 (N_3082,In_612,In_1391);
xor U3083 (N_3083,In_739,In_303);
xnor U3084 (N_3084,In_1044,In_1272);
nor U3085 (N_3085,In_382,In_1024);
nand U3086 (N_3086,In_537,In_495);
or U3087 (N_3087,In_286,In_84);
nor U3088 (N_3088,In_544,In_437);
nand U3089 (N_3089,In_1475,In_620);
nor U3090 (N_3090,In_413,In_1083);
nor U3091 (N_3091,In_1458,In_470);
nor U3092 (N_3092,In_1159,In_871);
and U3093 (N_3093,In_1026,In_7);
and U3094 (N_3094,In_492,In_1384);
and U3095 (N_3095,In_1091,In_1407);
nand U3096 (N_3096,In_1386,In_1483);
nor U3097 (N_3097,In_1050,In_1060);
and U3098 (N_3098,In_72,In_191);
or U3099 (N_3099,In_118,In_554);
or U3100 (N_3100,In_236,In_135);
nor U3101 (N_3101,In_477,In_1486);
or U3102 (N_3102,In_1485,In_793);
or U3103 (N_3103,In_536,In_519);
nor U3104 (N_3104,In_1336,In_1093);
nor U3105 (N_3105,In_525,In_1378);
and U3106 (N_3106,In_1054,In_545);
or U3107 (N_3107,In_240,In_898);
and U3108 (N_3108,In_684,In_1386);
or U3109 (N_3109,In_379,In_1343);
and U3110 (N_3110,In_361,In_1309);
or U3111 (N_3111,In_99,In_1017);
and U3112 (N_3112,In_217,In_366);
or U3113 (N_3113,In_1233,In_982);
nor U3114 (N_3114,In_793,In_1025);
and U3115 (N_3115,In_1229,In_1150);
nor U3116 (N_3116,In_1426,In_1320);
nand U3117 (N_3117,In_730,In_1015);
and U3118 (N_3118,In_338,In_141);
nand U3119 (N_3119,In_609,In_1387);
nor U3120 (N_3120,In_640,In_530);
nand U3121 (N_3121,In_742,In_9);
or U3122 (N_3122,In_1119,In_1393);
nand U3123 (N_3123,In_1198,In_1395);
and U3124 (N_3124,In_33,In_1433);
and U3125 (N_3125,In_12,In_812);
and U3126 (N_3126,In_249,In_239);
nand U3127 (N_3127,In_430,In_539);
nor U3128 (N_3128,In_1222,In_1437);
xnor U3129 (N_3129,In_211,In_449);
and U3130 (N_3130,In_91,In_300);
nor U3131 (N_3131,In_484,In_680);
nor U3132 (N_3132,In_985,In_616);
nor U3133 (N_3133,In_1408,In_295);
nand U3134 (N_3134,In_1017,In_337);
or U3135 (N_3135,In_887,In_555);
and U3136 (N_3136,In_765,In_737);
or U3137 (N_3137,In_960,In_708);
nand U3138 (N_3138,In_382,In_1418);
nand U3139 (N_3139,In_151,In_944);
or U3140 (N_3140,In_1097,In_1060);
nor U3141 (N_3141,In_398,In_294);
and U3142 (N_3142,In_1309,In_811);
and U3143 (N_3143,In_914,In_1346);
or U3144 (N_3144,In_790,In_923);
nor U3145 (N_3145,In_698,In_206);
nand U3146 (N_3146,In_1462,In_208);
nand U3147 (N_3147,In_1019,In_1249);
or U3148 (N_3148,In_945,In_131);
or U3149 (N_3149,In_341,In_93);
and U3150 (N_3150,In_604,In_865);
nor U3151 (N_3151,In_441,In_652);
or U3152 (N_3152,In_1244,In_865);
and U3153 (N_3153,In_385,In_1483);
nand U3154 (N_3154,In_203,In_306);
nand U3155 (N_3155,In_637,In_1387);
and U3156 (N_3156,In_1310,In_1377);
or U3157 (N_3157,In_221,In_724);
nor U3158 (N_3158,In_274,In_1142);
and U3159 (N_3159,In_135,In_15);
or U3160 (N_3160,In_1018,In_151);
nand U3161 (N_3161,In_1081,In_1041);
nand U3162 (N_3162,In_63,In_108);
nand U3163 (N_3163,In_887,In_592);
or U3164 (N_3164,In_913,In_977);
nor U3165 (N_3165,In_496,In_716);
nor U3166 (N_3166,In_1069,In_1495);
and U3167 (N_3167,In_906,In_40);
and U3168 (N_3168,In_1263,In_550);
or U3169 (N_3169,In_1098,In_276);
nand U3170 (N_3170,In_439,In_199);
and U3171 (N_3171,In_1060,In_84);
and U3172 (N_3172,In_416,In_1229);
xnor U3173 (N_3173,In_1365,In_46);
nand U3174 (N_3174,In_689,In_490);
or U3175 (N_3175,In_726,In_690);
nor U3176 (N_3176,In_290,In_250);
and U3177 (N_3177,In_1449,In_1045);
and U3178 (N_3178,In_554,In_392);
or U3179 (N_3179,In_1258,In_206);
and U3180 (N_3180,In_631,In_1439);
nor U3181 (N_3181,In_1251,In_899);
nor U3182 (N_3182,In_544,In_1396);
or U3183 (N_3183,In_1339,In_556);
nand U3184 (N_3184,In_1322,In_773);
nor U3185 (N_3185,In_1353,In_466);
nand U3186 (N_3186,In_665,In_167);
nor U3187 (N_3187,In_668,In_1145);
nor U3188 (N_3188,In_1081,In_136);
nor U3189 (N_3189,In_131,In_356);
or U3190 (N_3190,In_626,In_276);
or U3191 (N_3191,In_633,In_892);
or U3192 (N_3192,In_526,In_16);
nor U3193 (N_3193,In_498,In_238);
nand U3194 (N_3194,In_418,In_1273);
or U3195 (N_3195,In_879,In_41);
nor U3196 (N_3196,In_859,In_315);
nor U3197 (N_3197,In_396,In_12);
and U3198 (N_3198,In_1248,In_527);
and U3199 (N_3199,In_178,In_387);
and U3200 (N_3200,In_1254,In_1383);
nand U3201 (N_3201,In_651,In_1280);
nor U3202 (N_3202,In_1089,In_1118);
nand U3203 (N_3203,In_789,In_1481);
nor U3204 (N_3204,In_235,In_1227);
nand U3205 (N_3205,In_736,In_822);
nand U3206 (N_3206,In_225,In_221);
nand U3207 (N_3207,In_192,In_1229);
nand U3208 (N_3208,In_546,In_311);
and U3209 (N_3209,In_795,In_976);
nor U3210 (N_3210,In_9,In_138);
and U3211 (N_3211,In_855,In_1478);
or U3212 (N_3212,In_339,In_901);
nor U3213 (N_3213,In_189,In_498);
and U3214 (N_3214,In_556,In_932);
nand U3215 (N_3215,In_95,In_1419);
or U3216 (N_3216,In_1335,In_740);
nor U3217 (N_3217,In_510,In_251);
and U3218 (N_3218,In_640,In_238);
nand U3219 (N_3219,In_811,In_488);
nor U3220 (N_3220,In_674,In_807);
nor U3221 (N_3221,In_1178,In_738);
nand U3222 (N_3222,In_96,In_126);
and U3223 (N_3223,In_275,In_401);
or U3224 (N_3224,In_300,In_740);
or U3225 (N_3225,In_939,In_1042);
nor U3226 (N_3226,In_49,In_1470);
and U3227 (N_3227,In_1251,In_1428);
and U3228 (N_3228,In_724,In_483);
and U3229 (N_3229,In_389,In_971);
or U3230 (N_3230,In_583,In_773);
or U3231 (N_3231,In_503,In_29);
or U3232 (N_3232,In_1494,In_419);
and U3233 (N_3233,In_587,In_995);
or U3234 (N_3234,In_799,In_1235);
or U3235 (N_3235,In_377,In_25);
nand U3236 (N_3236,In_912,In_701);
nor U3237 (N_3237,In_649,In_266);
or U3238 (N_3238,In_907,In_625);
and U3239 (N_3239,In_184,In_339);
nor U3240 (N_3240,In_1113,In_825);
or U3241 (N_3241,In_206,In_1453);
xor U3242 (N_3242,In_825,In_225);
or U3243 (N_3243,In_870,In_1304);
and U3244 (N_3244,In_1022,In_477);
and U3245 (N_3245,In_316,In_534);
and U3246 (N_3246,In_1048,In_122);
nor U3247 (N_3247,In_218,In_731);
and U3248 (N_3248,In_804,In_943);
nand U3249 (N_3249,In_1284,In_586);
nand U3250 (N_3250,In_1175,In_828);
nand U3251 (N_3251,In_596,In_1162);
nand U3252 (N_3252,In_728,In_239);
or U3253 (N_3253,In_1372,In_560);
and U3254 (N_3254,In_246,In_930);
and U3255 (N_3255,In_1285,In_281);
nand U3256 (N_3256,In_542,In_178);
nor U3257 (N_3257,In_475,In_778);
nor U3258 (N_3258,In_194,In_1233);
or U3259 (N_3259,In_160,In_281);
xor U3260 (N_3260,In_943,In_672);
or U3261 (N_3261,In_1129,In_1388);
and U3262 (N_3262,In_27,In_644);
or U3263 (N_3263,In_697,In_793);
and U3264 (N_3264,In_217,In_795);
and U3265 (N_3265,In_695,In_237);
or U3266 (N_3266,In_40,In_544);
and U3267 (N_3267,In_54,In_576);
nand U3268 (N_3268,In_257,In_1376);
nor U3269 (N_3269,In_153,In_1187);
nand U3270 (N_3270,In_1017,In_1459);
and U3271 (N_3271,In_1361,In_921);
or U3272 (N_3272,In_1330,In_1047);
nor U3273 (N_3273,In_149,In_1375);
and U3274 (N_3274,In_322,In_407);
or U3275 (N_3275,In_533,In_780);
nor U3276 (N_3276,In_1146,In_781);
or U3277 (N_3277,In_367,In_58);
nor U3278 (N_3278,In_22,In_1025);
or U3279 (N_3279,In_713,In_215);
nand U3280 (N_3280,In_441,In_906);
nor U3281 (N_3281,In_906,In_650);
and U3282 (N_3282,In_921,In_808);
nor U3283 (N_3283,In_375,In_634);
or U3284 (N_3284,In_1405,In_908);
nand U3285 (N_3285,In_1459,In_832);
nor U3286 (N_3286,In_413,In_107);
nor U3287 (N_3287,In_382,In_191);
or U3288 (N_3288,In_4,In_35);
nor U3289 (N_3289,In_343,In_601);
and U3290 (N_3290,In_301,In_945);
and U3291 (N_3291,In_1258,In_1396);
nand U3292 (N_3292,In_1187,In_362);
and U3293 (N_3293,In_443,In_378);
nand U3294 (N_3294,In_336,In_1361);
nand U3295 (N_3295,In_233,In_1042);
nand U3296 (N_3296,In_1457,In_806);
nand U3297 (N_3297,In_1211,In_485);
nand U3298 (N_3298,In_674,In_1435);
nor U3299 (N_3299,In_808,In_217);
or U3300 (N_3300,In_264,In_1295);
and U3301 (N_3301,In_127,In_759);
and U3302 (N_3302,In_390,In_1439);
or U3303 (N_3303,In_1305,In_325);
or U3304 (N_3304,In_1170,In_941);
or U3305 (N_3305,In_1432,In_1127);
and U3306 (N_3306,In_179,In_521);
nand U3307 (N_3307,In_943,In_420);
nand U3308 (N_3308,In_712,In_303);
or U3309 (N_3309,In_1257,In_1110);
and U3310 (N_3310,In_626,In_225);
and U3311 (N_3311,In_1271,In_722);
nand U3312 (N_3312,In_1035,In_784);
nor U3313 (N_3313,In_761,In_689);
nor U3314 (N_3314,In_1015,In_144);
or U3315 (N_3315,In_821,In_1386);
nor U3316 (N_3316,In_901,In_1196);
or U3317 (N_3317,In_284,In_960);
and U3318 (N_3318,In_1281,In_260);
and U3319 (N_3319,In_157,In_1445);
nand U3320 (N_3320,In_1134,In_1168);
and U3321 (N_3321,In_1126,In_1353);
and U3322 (N_3322,In_382,In_686);
or U3323 (N_3323,In_353,In_73);
nand U3324 (N_3324,In_911,In_917);
or U3325 (N_3325,In_1482,In_1084);
nor U3326 (N_3326,In_134,In_500);
and U3327 (N_3327,In_208,In_1244);
or U3328 (N_3328,In_1285,In_916);
or U3329 (N_3329,In_530,In_708);
or U3330 (N_3330,In_340,In_404);
or U3331 (N_3331,In_1095,In_1016);
nor U3332 (N_3332,In_35,In_402);
nor U3333 (N_3333,In_653,In_1428);
or U3334 (N_3334,In_94,In_1247);
nand U3335 (N_3335,In_27,In_388);
and U3336 (N_3336,In_353,In_1235);
or U3337 (N_3337,In_1283,In_526);
nand U3338 (N_3338,In_605,In_804);
nand U3339 (N_3339,In_318,In_765);
nor U3340 (N_3340,In_173,In_1119);
or U3341 (N_3341,In_801,In_709);
nor U3342 (N_3342,In_789,In_453);
and U3343 (N_3343,In_187,In_519);
nand U3344 (N_3344,In_600,In_172);
nand U3345 (N_3345,In_968,In_698);
nand U3346 (N_3346,In_792,In_736);
xnor U3347 (N_3347,In_487,In_400);
nand U3348 (N_3348,In_1352,In_753);
nor U3349 (N_3349,In_1195,In_1243);
or U3350 (N_3350,In_284,In_982);
and U3351 (N_3351,In_177,In_706);
nand U3352 (N_3352,In_519,In_1074);
or U3353 (N_3353,In_64,In_1041);
and U3354 (N_3354,In_635,In_61);
nor U3355 (N_3355,In_633,In_283);
and U3356 (N_3356,In_1364,In_1238);
or U3357 (N_3357,In_1477,In_913);
nand U3358 (N_3358,In_1133,In_708);
or U3359 (N_3359,In_266,In_466);
nor U3360 (N_3360,In_592,In_1450);
and U3361 (N_3361,In_400,In_287);
or U3362 (N_3362,In_1496,In_562);
nand U3363 (N_3363,In_737,In_725);
nand U3364 (N_3364,In_194,In_660);
or U3365 (N_3365,In_1016,In_1067);
or U3366 (N_3366,In_884,In_354);
nor U3367 (N_3367,In_1155,In_525);
or U3368 (N_3368,In_686,In_1296);
or U3369 (N_3369,In_1429,In_1291);
or U3370 (N_3370,In_1153,In_799);
and U3371 (N_3371,In_1004,In_1091);
and U3372 (N_3372,In_19,In_804);
or U3373 (N_3373,In_184,In_671);
nand U3374 (N_3374,In_731,In_837);
nor U3375 (N_3375,In_1471,In_501);
nand U3376 (N_3376,In_1374,In_54);
or U3377 (N_3377,In_570,In_405);
or U3378 (N_3378,In_222,In_282);
and U3379 (N_3379,In_1020,In_353);
or U3380 (N_3380,In_1065,In_259);
nand U3381 (N_3381,In_581,In_319);
nor U3382 (N_3382,In_694,In_1026);
and U3383 (N_3383,In_1108,In_787);
and U3384 (N_3384,In_538,In_1153);
and U3385 (N_3385,In_807,In_190);
nor U3386 (N_3386,In_625,In_740);
nand U3387 (N_3387,In_827,In_905);
and U3388 (N_3388,In_1374,In_1431);
and U3389 (N_3389,In_743,In_982);
or U3390 (N_3390,In_1251,In_1297);
nor U3391 (N_3391,In_872,In_801);
nand U3392 (N_3392,In_469,In_740);
and U3393 (N_3393,In_970,In_647);
and U3394 (N_3394,In_1422,In_561);
and U3395 (N_3395,In_483,In_530);
and U3396 (N_3396,In_1443,In_1048);
and U3397 (N_3397,In_321,In_687);
or U3398 (N_3398,In_933,In_450);
nand U3399 (N_3399,In_744,In_652);
nand U3400 (N_3400,In_1194,In_759);
or U3401 (N_3401,In_266,In_127);
nor U3402 (N_3402,In_487,In_15);
nor U3403 (N_3403,In_1193,In_1388);
nand U3404 (N_3404,In_160,In_1011);
or U3405 (N_3405,In_1164,In_947);
nor U3406 (N_3406,In_619,In_1087);
and U3407 (N_3407,In_269,In_1168);
nand U3408 (N_3408,In_661,In_227);
or U3409 (N_3409,In_840,In_1429);
or U3410 (N_3410,In_863,In_1060);
or U3411 (N_3411,In_978,In_1418);
nor U3412 (N_3412,In_1010,In_508);
nor U3413 (N_3413,In_165,In_911);
and U3414 (N_3414,In_648,In_658);
or U3415 (N_3415,In_62,In_1274);
or U3416 (N_3416,In_401,In_185);
nand U3417 (N_3417,In_165,In_107);
and U3418 (N_3418,In_844,In_429);
and U3419 (N_3419,In_125,In_794);
and U3420 (N_3420,In_1470,In_1497);
nand U3421 (N_3421,In_759,In_750);
or U3422 (N_3422,In_436,In_392);
or U3423 (N_3423,In_564,In_1125);
or U3424 (N_3424,In_252,In_1083);
or U3425 (N_3425,In_921,In_209);
nand U3426 (N_3426,In_800,In_1150);
and U3427 (N_3427,In_50,In_884);
and U3428 (N_3428,In_1465,In_1375);
nand U3429 (N_3429,In_744,In_1089);
and U3430 (N_3430,In_134,In_877);
nand U3431 (N_3431,In_1004,In_408);
or U3432 (N_3432,In_726,In_894);
nor U3433 (N_3433,In_188,In_1372);
nor U3434 (N_3434,In_22,In_331);
nand U3435 (N_3435,In_204,In_1454);
nor U3436 (N_3436,In_1008,In_1244);
nand U3437 (N_3437,In_156,In_1077);
or U3438 (N_3438,In_416,In_1368);
and U3439 (N_3439,In_1182,In_209);
and U3440 (N_3440,In_770,In_1054);
and U3441 (N_3441,In_297,In_1237);
nor U3442 (N_3442,In_292,In_1452);
or U3443 (N_3443,In_354,In_1059);
nor U3444 (N_3444,In_1023,In_873);
xnor U3445 (N_3445,In_118,In_622);
and U3446 (N_3446,In_696,In_612);
and U3447 (N_3447,In_564,In_637);
or U3448 (N_3448,In_1417,In_93);
and U3449 (N_3449,In_1492,In_1250);
nand U3450 (N_3450,In_265,In_1225);
or U3451 (N_3451,In_661,In_7);
nor U3452 (N_3452,In_281,In_1013);
nor U3453 (N_3453,In_416,In_352);
nand U3454 (N_3454,In_987,In_120);
and U3455 (N_3455,In_1421,In_460);
nor U3456 (N_3456,In_740,In_637);
or U3457 (N_3457,In_179,In_961);
nand U3458 (N_3458,In_1165,In_1426);
nand U3459 (N_3459,In_1022,In_817);
or U3460 (N_3460,In_64,In_720);
nor U3461 (N_3461,In_839,In_609);
nor U3462 (N_3462,In_1195,In_961);
nor U3463 (N_3463,In_499,In_1213);
or U3464 (N_3464,In_994,In_1422);
or U3465 (N_3465,In_733,In_1387);
and U3466 (N_3466,In_1113,In_81);
nor U3467 (N_3467,In_1170,In_1007);
and U3468 (N_3468,In_42,In_897);
or U3469 (N_3469,In_90,In_1483);
nor U3470 (N_3470,In_28,In_795);
or U3471 (N_3471,In_635,In_947);
and U3472 (N_3472,In_770,In_907);
and U3473 (N_3473,In_1426,In_1336);
nor U3474 (N_3474,In_142,In_1123);
or U3475 (N_3475,In_875,In_272);
and U3476 (N_3476,In_790,In_385);
nand U3477 (N_3477,In_751,In_1093);
and U3478 (N_3478,In_1004,In_359);
nor U3479 (N_3479,In_567,In_1082);
nor U3480 (N_3480,In_944,In_322);
nor U3481 (N_3481,In_342,In_1128);
or U3482 (N_3482,In_821,In_721);
nand U3483 (N_3483,In_724,In_259);
nor U3484 (N_3484,In_1465,In_478);
and U3485 (N_3485,In_570,In_225);
xnor U3486 (N_3486,In_1001,In_376);
or U3487 (N_3487,In_641,In_921);
nor U3488 (N_3488,In_166,In_71);
nor U3489 (N_3489,In_220,In_816);
or U3490 (N_3490,In_403,In_1489);
and U3491 (N_3491,In_889,In_875);
or U3492 (N_3492,In_381,In_1354);
or U3493 (N_3493,In_1399,In_1013);
nor U3494 (N_3494,In_710,In_16);
nand U3495 (N_3495,In_401,In_500);
and U3496 (N_3496,In_273,In_465);
or U3497 (N_3497,In_1374,In_998);
and U3498 (N_3498,In_704,In_737);
nor U3499 (N_3499,In_238,In_1089);
nand U3500 (N_3500,In_1364,In_547);
nand U3501 (N_3501,In_1193,In_875);
nor U3502 (N_3502,In_156,In_340);
xor U3503 (N_3503,In_1480,In_111);
nand U3504 (N_3504,In_243,In_1347);
or U3505 (N_3505,In_676,In_1388);
nor U3506 (N_3506,In_949,In_891);
or U3507 (N_3507,In_330,In_110);
and U3508 (N_3508,In_708,In_1413);
or U3509 (N_3509,In_504,In_430);
nand U3510 (N_3510,In_247,In_341);
and U3511 (N_3511,In_156,In_1069);
or U3512 (N_3512,In_297,In_929);
nand U3513 (N_3513,In_1413,In_137);
nand U3514 (N_3514,In_1415,In_254);
or U3515 (N_3515,In_1390,In_1389);
nand U3516 (N_3516,In_645,In_291);
nand U3517 (N_3517,In_795,In_1054);
or U3518 (N_3518,In_188,In_526);
and U3519 (N_3519,In_918,In_960);
nand U3520 (N_3520,In_1310,In_1066);
and U3521 (N_3521,In_729,In_740);
and U3522 (N_3522,In_925,In_752);
nand U3523 (N_3523,In_1,In_1061);
and U3524 (N_3524,In_684,In_1357);
xnor U3525 (N_3525,In_801,In_284);
and U3526 (N_3526,In_990,In_1149);
and U3527 (N_3527,In_150,In_857);
and U3528 (N_3528,In_46,In_113);
and U3529 (N_3529,In_439,In_1234);
xnor U3530 (N_3530,In_523,In_866);
and U3531 (N_3531,In_1080,In_616);
nand U3532 (N_3532,In_506,In_1128);
or U3533 (N_3533,In_1405,In_568);
nand U3534 (N_3534,In_741,In_338);
nor U3535 (N_3535,In_595,In_698);
nand U3536 (N_3536,In_244,In_1461);
xnor U3537 (N_3537,In_209,In_925);
or U3538 (N_3538,In_1388,In_989);
or U3539 (N_3539,In_717,In_1229);
nand U3540 (N_3540,In_782,In_806);
nor U3541 (N_3541,In_1472,In_301);
xor U3542 (N_3542,In_960,In_732);
or U3543 (N_3543,In_1009,In_1179);
nand U3544 (N_3544,In_463,In_26);
or U3545 (N_3545,In_608,In_854);
nand U3546 (N_3546,In_1369,In_326);
or U3547 (N_3547,In_552,In_311);
and U3548 (N_3548,In_1246,In_464);
and U3549 (N_3549,In_1077,In_606);
and U3550 (N_3550,In_1341,In_72);
nor U3551 (N_3551,In_609,In_672);
and U3552 (N_3552,In_659,In_1027);
nor U3553 (N_3553,In_557,In_669);
or U3554 (N_3554,In_331,In_884);
nor U3555 (N_3555,In_536,In_56);
nor U3556 (N_3556,In_537,In_436);
nor U3557 (N_3557,In_656,In_1052);
and U3558 (N_3558,In_1240,In_1072);
or U3559 (N_3559,In_1127,In_1288);
or U3560 (N_3560,In_1362,In_548);
and U3561 (N_3561,In_99,In_1376);
or U3562 (N_3562,In_564,In_487);
or U3563 (N_3563,In_1019,In_1214);
and U3564 (N_3564,In_1181,In_1047);
nand U3565 (N_3565,In_426,In_1467);
or U3566 (N_3566,In_1432,In_47);
nor U3567 (N_3567,In_1325,In_650);
and U3568 (N_3568,In_87,In_994);
or U3569 (N_3569,In_1293,In_1140);
nand U3570 (N_3570,In_666,In_173);
nor U3571 (N_3571,In_1153,In_1341);
nand U3572 (N_3572,In_199,In_232);
and U3573 (N_3573,In_751,In_508);
or U3574 (N_3574,In_381,In_1198);
and U3575 (N_3575,In_293,In_1229);
nor U3576 (N_3576,In_319,In_934);
or U3577 (N_3577,In_68,In_190);
nand U3578 (N_3578,In_582,In_496);
and U3579 (N_3579,In_715,In_536);
nor U3580 (N_3580,In_1458,In_1280);
nand U3581 (N_3581,In_97,In_541);
nand U3582 (N_3582,In_789,In_283);
nor U3583 (N_3583,In_886,In_343);
nand U3584 (N_3584,In_297,In_864);
and U3585 (N_3585,In_112,In_1239);
nor U3586 (N_3586,In_1164,In_458);
nand U3587 (N_3587,In_24,In_477);
or U3588 (N_3588,In_106,In_1489);
nor U3589 (N_3589,In_966,In_217);
nor U3590 (N_3590,In_35,In_288);
nand U3591 (N_3591,In_50,In_96);
and U3592 (N_3592,In_832,In_711);
and U3593 (N_3593,In_589,In_291);
or U3594 (N_3594,In_1270,In_806);
nand U3595 (N_3595,In_493,In_782);
nand U3596 (N_3596,In_1403,In_1296);
nor U3597 (N_3597,In_1081,In_139);
nor U3598 (N_3598,In_692,In_213);
and U3599 (N_3599,In_1393,In_853);
and U3600 (N_3600,In_611,In_96);
nor U3601 (N_3601,In_1252,In_19);
and U3602 (N_3602,In_1205,In_714);
or U3603 (N_3603,In_1015,In_1008);
nand U3604 (N_3604,In_1159,In_151);
nor U3605 (N_3605,In_1443,In_1);
or U3606 (N_3606,In_1356,In_1471);
and U3607 (N_3607,In_618,In_45);
nand U3608 (N_3608,In_1372,In_517);
or U3609 (N_3609,In_83,In_288);
nand U3610 (N_3610,In_1080,In_335);
or U3611 (N_3611,In_544,In_123);
and U3612 (N_3612,In_788,In_665);
and U3613 (N_3613,In_551,In_686);
nand U3614 (N_3614,In_1167,In_1259);
nor U3615 (N_3615,In_329,In_1308);
nor U3616 (N_3616,In_233,In_248);
nor U3617 (N_3617,In_514,In_792);
and U3618 (N_3618,In_1176,In_1387);
nor U3619 (N_3619,In_1306,In_181);
nand U3620 (N_3620,In_1034,In_973);
or U3621 (N_3621,In_1280,In_7);
nor U3622 (N_3622,In_595,In_228);
and U3623 (N_3623,In_1236,In_615);
nor U3624 (N_3624,In_305,In_790);
or U3625 (N_3625,In_524,In_1157);
and U3626 (N_3626,In_1076,In_1301);
or U3627 (N_3627,In_1284,In_632);
or U3628 (N_3628,In_367,In_722);
or U3629 (N_3629,In_91,In_1272);
and U3630 (N_3630,In_1331,In_1202);
and U3631 (N_3631,In_83,In_715);
nor U3632 (N_3632,In_175,In_132);
or U3633 (N_3633,In_1258,In_1191);
or U3634 (N_3634,In_1143,In_190);
nand U3635 (N_3635,In_598,In_1392);
nor U3636 (N_3636,In_1024,In_508);
nand U3637 (N_3637,In_317,In_347);
nand U3638 (N_3638,In_1212,In_1426);
or U3639 (N_3639,In_1185,In_895);
or U3640 (N_3640,In_569,In_582);
nand U3641 (N_3641,In_310,In_526);
nor U3642 (N_3642,In_588,In_1478);
or U3643 (N_3643,In_597,In_809);
nand U3644 (N_3644,In_157,In_861);
nand U3645 (N_3645,In_92,In_1268);
nand U3646 (N_3646,In_1172,In_1259);
nor U3647 (N_3647,In_67,In_569);
nor U3648 (N_3648,In_581,In_530);
or U3649 (N_3649,In_1099,In_1251);
or U3650 (N_3650,In_59,In_1130);
nand U3651 (N_3651,In_1042,In_749);
nor U3652 (N_3652,In_1479,In_573);
nor U3653 (N_3653,In_1364,In_229);
nand U3654 (N_3654,In_1448,In_917);
and U3655 (N_3655,In_1028,In_701);
or U3656 (N_3656,In_394,In_890);
nand U3657 (N_3657,In_1177,In_355);
and U3658 (N_3658,In_279,In_280);
nand U3659 (N_3659,In_1424,In_387);
and U3660 (N_3660,In_1116,In_357);
nor U3661 (N_3661,In_1292,In_1362);
and U3662 (N_3662,In_255,In_753);
and U3663 (N_3663,In_601,In_214);
nand U3664 (N_3664,In_68,In_537);
and U3665 (N_3665,In_1487,In_487);
or U3666 (N_3666,In_792,In_1329);
nor U3667 (N_3667,In_1192,In_494);
or U3668 (N_3668,In_1462,In_1318);
nand U3669 (N_3669,In_774,In_453);
and U3670 (N_3670,In_148,In_1171);
nor U3671 (N_3671,In_1318,In_1061);
or U3672 (N_3672,In_1488,In_727);
and U3673 (N_3673,In_175,In_1456);
and U3674 (N_3674,In_1386,In_730);
and U3675 (N_3675,In_1171,In_741);
and U3676 (N_3676,In_1287,In_1295);
or U3677 (N_3677,In_214,In_784);
nand U3678 (N_3678,In_334,In_914);
nor U3679 (N_3679,In_1412,In_1328);
or U3680 (N_3680,In_1460,In_1248);
nand U3681 (N_3681,In_33,In_1357);
or U3682 (N_3682,In_819,In_988);
or U3683 (N_3683,In_488,In_965);
nor U3684 (N_3684,In_257,In_208);
nand U3685 (N_3685,In_639,In_705);
nand U3686 (N_3686,In_1087,In_685);
nand U3687 (N_3687,In_964,In_530);
nand U3688 (N_3688,In_1464,In_35);
nand U3689 (N_3689,In_307,In_1051);
and U3690 (N_3690,In_230,In_206);
and U3691 (N_3691,In_499,In_1017);
nor U3692 (N_3692,In_576,In_287);
and U3693 (N_3693,In_520,In_584);
and U3694 (N_3694,In_1238,In_431);
and U3695 (N_3695,In_126,In_1246);
or U3696 (N_3696,In_452,In_1467);
and U3697 (N_3697,In_640,In_1268);
or U3698 (N_3698,In_536,In_1456);
nand U3699 (N_3699,In_1206,In_1034);
or U3700 (N_3700,In_490,In_472);
or U3701 (N_3701,In_1357,In_450);
nor U3702 (N_3702,In_1105,In_630);
nor U3703 (N_3703,In_827,In_1221);
nand U3704 (N_3704,In_791,In_742);
or U3705 (N_3705,In_16,In_847);
nand U3706 (N_3706,In_1039,In_382);
or U3707 (N_3707,In_2,In_1377);
nand U3708 (N_3708,In_1006,In_1045);
nor U3709 (N_3709,In_976,In_207);
nand U3710 (N_3710,In_1210,In_155);
and U3711 (N_3711,In_1345,In_854);
or U3712 (N_3712,In_371,In_438);
or U3713 (N_3713,In_1418,In_1350);
or U3714 (N_3714,In_1077,In_656);
nor U3715 (N_3715,In_863,In_1104);
nand U3716 (N_3716,In_878,In_1261);
nor U3717 (N_3717,In_352,In_907);
nand U3718 (N_3718,In_717,In_846);
and U3719 (N_3719,In_883,In_796);
nand U3720 (N_3720,In_929,In_921);
nor U3721 (N_3721,In_9,In_769);
and U3722 (N_3722,In_758,In_1421);
nor U3723 (N_3723,In_1435,In_169);
nand U3724 (N_3724,In_702,In_1330);
nand U3725 (N_3725,In_1205,In_57);
and U3726 (N_3726,In_1011,In_93);
or U3727 (N_3727,In_1273,In_1023);
nor U3728 (N_3728,In_531,In_146);
or U3729 (N_3729,In_1109,In_1194);
nor U3730 (N_3730,In_1074,In_919);
nor U3731 (N_3731,In_560,In_1076);
and U3732 (N_3732,In_1016,In_803);
nor U3733 (N_3733,In_181,In_761);
nor U3734 (N_3734,In_482,In_633);
or U3735 (N_3735,In_236,In_811);
and U3736 (N_3736,In_868,In_904);
or U3737 (N_3737,In_1195,In_927);
and U3738 (N_3738,In_1414,In_638);
nor U3739 (N_3739,In_1486,In_1233);
or U3740 (N_3740,In_905,In_1417);
nand U3741 (N_3741,In_1479,In_1243);
and U3742 (N_3742,In_101,In_796);
xnor U3743 (N_3743,In_345,In_626);
nand U3744 (N_3744,In_1060,In_807);
nor U3745 (N_3745,In_66,In_76);
or U3746 (N_3746,In_1262,In_1411);
or U3747 (N_3747,In_788,In_1233);
nor U3748 (N_3748,In_1184,In_18);
and U3749 (N_3749,In_718,In_889);
or U3750 (N_3750,In_1477,In_186);
nor U3751 (N_3751,In_890,In_1290);
and U3752 (N_3752,In_320,In_1187);
nand U3753 (N_3753,In_1216,In_1199);
nor U3754 (N_3754,In_804,In_1146);
nand U3755 (N_3755,In_291,In_1219);
and U3756 (N_3756,In_220,In_88);
nor U3757 (N_3757,In_328,In_1383);
nand U3758 (N_3758,In_535,In_882);
nand U3759 (N_3759,In_1206,In_834);
or U3760 (N_3760,In_1034,In_747);
or U3761 (N_3761,In_791,In_1314);
or U3762 (N_3762,In_507,In_438);
and U3763 (N_3763,In_1054,In_10);
and U3764 (N_3764,In_515,In_1085);
and U3765 (N_3765,In_670,In_517);
nor U3766 (N_3766,In_139,In_1451);
and U3767 (N_3767,In_1100,In_833);
nor U3768 (N_3768,In_517,In_1305);
or U3769 (N_3769,In_1428,In_964);
nor U3770 (N_3770,In_705,In_807);
or U3771 (N_3771,In_1140,In_470);
or U3772 (N_3772,In_805,In_1180);
nand U3773 (N_3773,In_679,In_1161);
and U3774 (N_3774,In_516,In_673);
nor U3775 (N_3775,In_652,In_1346);
nor U3776 (N_3776,In_233,In_443);
nand U3777 (N_3777,In_600,In_385);
or U3778 (N_3778,In_62,In_1238);
nor U3779 (N_3779,In_1126,In_505);
nand U3780 (N_3780,In_1461,In_140);
and U3781 (N_3781,In_308,In_362);
or U3782 (N_3782,In_993,In_69);
nand U3783 (N_3783,In_331,In_818);
and U3784 (N_3784,In_1140,In_561);
nand U3785 (N_3785,In_1277,In_1396);
or U3786 (N_3786,In_945,In_1016);
and U3787 (N_3787,In_458,In_765);
nor U3788 (N_3788,In_641,In_620);
and U3789 (N_3789,In_204,In_17);
and U3790 (N_3790,In_182,In_362);
nor U3791 (N_3791,In_1090,In_725);
nor U3792 (N_3792,In_497,In_430);
nand U3793 (N_3793,In_854,In_165);
and U3794 (N_3794,In_224,In_476);
nand U3795 (N_3795,In_656,In_260);
or U3796 (N_3796,In_684,In_225);
and U3797 (N_3797,In_1196,In_1078);
nor U3798 (N_3798,In_221,In_1247);
nor U3799 (N_3799,In_283,In_1428);
or U3800 (N_3800,In_219,In_298);
nor U3801 (N_3801,In_947,In_1446);
nor U3802 (N_3802,In_1124,In_1000);
and U3803 (N_3803,In_1168,In_781);
and U3804 (N_3804,In_750,In_381);
and U3805 (N_3805,In_820,In_34);
nand U3806 (N_3806,In_1282,In_1333);
and U3807 (N_3807,In_1054,In_1409);
or U3808 (N_3808,In_248,In_167);
or U3809 (N_3809,In_1486,In_1110);
or U3810 (N_3810,In_1065,In_247);
or U3811 (N_3811,In_841,In_339);
or U3812 (N_3812,In_136,In_730);
nor U3813 (N_3813,In_1263,In_156);
or U3814 (N_3814,In_787,In_1298);
nand U3815 (N_3815,In_56,In_204);
nor U3816 (N_3816,In_1045,In_724);
and U3817 (N_3817,In_1444,In_857);
or U3818 (N_3818,In_417,In_52);
nand U3819 (N_3819,In_1139,In_45);
and U3820 (N_3820,In_501,In_1211);
and U3821 (N_3821,In_1123,In_1292);
and U3822 (N_3822,In_1363,In_956);
nor U3823 (N_3823,In_1176,In_1287);
or U3824 (N_3824,In_585,In_456);
and U3825 (N_3825,In_507,In_1043);
or U3826 (N_3826,In_554,In_637);
nor U3827 (N_3827,In_1473,In_1078);
nor U3828 (N_3828,In_218,In_1038);
and U3829 (N_3829,In_200,In_1163);
nor U3830 (N_3830,In_484,In_335);
nand U3831 (N_3831,In_891,In_1086);
and U3832 (N_3832,In_1369,In_1329);
xor U3833 (N_3833,In_226,In_83);
nand U3834 (N_3834,In_291,In_1273);
nand U3835 (N_3835,In_937,In_451);
and U3836 (N_3836,In_6,In_1055);
nor U3837 (N_3837,In_1273,In_116);
nand U3838 (N_3838,In_71,In_517);
nor U3839 (N_3839,In_1280,In_96);
nand U3840 (N_3840,In_761,In_55);
nand U3841 (N_3841,In_1152,In_267);
nand U3842 (N_3842,In_1070,In_167);
or U3843 (N_3843,In_320,In_1002);
and U3844 (N_3844,In_1202,In_310);
nor U3845 (N_3845,In_1112,In_465);
nand U3846 (N_3846,In_187,In_1306);
nor U3847 (N_3847,In_503,In_1041);
nand U3848 (N_3848,In_1427,In_918);
and U3849 (N_3849,In_150,In_1411);
nor U3850 (N_3850,In_359,In_1013);
or U3851 (N_3851,In_693,In_1464);
nand U3852 (N_3852,In_85,In_1136);
nand U3853 (N_3853,In_859,In_988);
and U3854 (N_3854,In_473,In_111);
nor U3855 (N_3855,In_667,In_1160);
or U3856 (N_3856,In_444,In_734);
or U3857 (N_3857,In_142,In_499);
nand U3858 (N_3858,In_317,In_1300);
and U3859 (N_3859,In_89,In_1176);
nand U3860 (N_3860,In_77,In_679);
and U3861 (N_3861,In_912,In_1237);
or U3862 (N_3862,In_736,In_252);
nor U3863 (N_3863,In_1108,In_572);
and U3864 (N_3864,In_1399,In_1303);
nand U3865 (N_3865,In_188,In_1394);
or U3866 (N_3866,In_863,In_971);
or U3867 (N_3867,In_1437,In_61);
nor U3868 (N_3868,In_937,In_1212);
and U3869 (N_3869,In_520,In_175);
nand U3870 (N_3870,In_1081,In_992);
or U3871 (N_3871,In_1178,In_76);
nor U3872 (N_3872,In_1437,In_987);
nand U3873 (N_3873,In_978,In_1084);
or U3874 (N_3874,In_1048,In_484);
xor U3875 (N_3875,In_285,In_1416);
or U3876 (N_3876,In_1264,In_413);
and U3877 (N_3877,In_54,In_1305);
and U3878 (N_3878,In_1441,In_145);
nor U3879 (N_3879,In_116,In_674);
and U3880 (N_3880,In_68,In_728);
nand U3881 (N_3881,In_865,In_338);
nor U3882 (N_3882,In_717,In_1401);
nand U3883 (N_3883,In_1249,In_108);
xor U3884 (N_3884,In_1494,In_1364);
or U3885 (N_3885,In_631,In_227);
and U3886 (N_3886,In_812,In_493);
or U3887 (N_3887,In_209,In_1191);
nand U3888 (N_3888,In_1076,In_1336);
and U3889 (N_3889,In_304,In_1107);
and U3890 (N_3890,In_399,In_1154);
and U3891 (N_3891,In_1386,In_55);
or U3892 (N_3892,In_1411,In_1027);
nand U3893 (N_3893,In_1428,In_1347);
or U3894 (N_3894,In_1471,In_883);
and U3895 (N_3895,In_1169,In_419);
nor U3896 (N_3896,In_307,In_1151);
nand U3897 (N_3897,In_107,In_1058);
and U3898 (N_3898,In_378,In_557);
and U3899 (N_3899,In_1404,In_1474);
nand U3900 (N_3900,In_269,In_537);
nor U3901 (N_3901,In_1467,In_954);
or U3902 (N_3902,In_1264,In_434);
nand U3903 (N_3903,In_831,In_439);
nor U3904 (N_3904,In_159,In_1066);
nand U3905 (N_3905,In_694,In_1203);
or U3906 (N_3906,In_923,In_328);
nand U3907 (N_3907,In_707,In_977);
nand U3908 (N_3908,In_818,In_996);
and U3909 (N_3909,In_1316,In_858);
or U3910 (N_3910,In_1403,In_1416);
or U3911 (N_3911,In_1204,In_1350);
nor U3912 (N_3912,In_1104,In_1455);
nand U3913 (N_3913,In_643,In_1047);
or U3914 (N_3914,In_551,In_1236);
nor U3915 (N_3915,In_678,In_1328);
and U3916 (N_3916,In_304,In_1404);
or U3917 (N_3917,In_925,In_759);
nand U3918 (N_3918,In_108,In_662);
or U3919 (N_3919,In_564,In_414);
and U3920 (N_3920,In_140,In_419);
and U3921 (N_3921,In_346,In_1032);
nor U3922 (N_3922,In_1263,In_1024);
and U3923 (N_3923,In_358,In_48);
or U3924 (N_3924,In_678,In_717);
and U3925 (N_3925,In_1327,In_1050);
and U3926 (N_3926,In_144,In_1470);
or U3927 (N_3927,In_550,In_35);
nor U3928 (N_3928,In_900,In_936);
nor U3929 (N_3929,In_592,In_866);
and U3930 (N_3930,In_874,In_1475);
nand U3931 (N_3931,In_998,In_129);
or U3932 (N_3932,In_836,In_1113);
or U3933 (N_3933,In_742,In_766);
and U3934 (N_3934,In_694,In_906);
or U3935 (N_3935,In_473,In_297);
nor U3936 (N_3936,In_913,In_552);
nand U3937 (N_3937,In_437,In_938);
nand U3938 (N_3938,In_1368,In_196);
and U3939 (N_3939,In_550,In_841);
nand U3940 (N_3940,In_1464,In_534);
nor U3941 (N_3941,In_1260,In_10);
or U3942 (N_3942,In_327,In_276);
nor U3943 (N_3943,In_1442,In_862);
and U3944 (N_3944,In_253,In_1001);
or U3945 (N_3945,In_281,In_1181);
and U3946 (N_3946,In_59,In_557);
and U3947 (N_3947,In_1476,In_516);
nand U3948 (N_3948,In_1104,In_478);
nand U3949 (N_3949,In_704,In_638);
and U3950 (N_3950,In_964,In_1118);
or U3951 (N_3951,In_437,In_1113);
and U3952 (N_3952,In_1383,In_726);
nor U3953 (N_3953,In_450,In_510);
and U3954 (N_3954,In_1207,In_262);
or U3955 (N_3955,In_280,In_1265);
and U3956 (N_3956,In_200,In_983);
and U3957 (N_3957,In_895,In_566);
nor U3958 (N_3958,In_449,In_804);
nand U3959 (N_3959,In_1270,In_1289);
nor U3960 (N_3960,In_1320,In_1065);
nor U3961 (N_3961,In_1055,In_636);
and U3962 (N_3962,In_779,In_771);
or U3963 (N_3963,In_1169,In_1483);
or U3964 (N_3964,In_1186,In_958);
and U3965 (N_3965,In_341,In_1082);
nand U3966 (N_3966,In_1340,In_173);
and U3967 (N_3967,In_887,In_190);
or U3968 (N_3968,In_1180,In_887);
nand U3969 (N_3969,In_880,In_1417);
nand U3970 (N_3970,In_901,In_968);
or U3971 (N_3971,In_766,In_86);
nor U3972 (N_3972,In_1499,In_1076);
or U3973 (N_3973,In_806,In_250);
nor U3974 (N_3974,In_1498,In_606);
nand U3975 (N_3975,In_136,In_1426);
or U3976 (N_3976,In_1220,In_114);
or U3977 (N_3977,In_1045,In_649);
and U3978 (N_3978,In_1195,In_672);
nor U3979 (N_3979,In_29,In_328);
and U3980 (N_3980,In_1301,In_1370);
nand U3981 (N_3981,In_510,In_390);
nor U3982 (N_3982,In_1411,In_985);
nor U3983 (N_3983,In_629,In_170);
and U3984 (N_3984,In_356,In_13);
nor U3985 (N_3985,In_1317,In_1229);
nor U3986 (N_3986,In_108,In_1340);
and U3987 (N_3987,In_1154,In_601);
nor U3988 (N_3988,In_660,In_281);
nand U3989 (N_3989,In_210,In_1364);
or U3990 (N_3990,In_7,In_946);
nand U3991 (N_3991,In_417,In_955);
nor U3992 (N_3992,In_221,In_507);
and U3993 (N_3993,In_847,In_1143);
nand U3994 (N_3994,In_416,In_1014);
and U3995 (N_3995,In_45,In_16);
and U3996 (N_3996,In_776,In_89);
nand U3997 (N_3997,In_1171,In_506);
nand U3998 (N_3998,In_348,In_878);
xor U3999 (N_3999,In_474,In_292);
or U4000 (N_4000,In_1023,In_42);
nand U4001 (N_4001,In_473,In_10);
and U4002 (N_4002,In_887,In_1232);
nor U4003 (N_4003,In_989,In_600);
or U4004 (N_4004,In_492,In_719);
nor U4005 (N_4005,In_60,In_423);
nor U4006 (N_4006,In_282,In_409);
nand U4007 (N_4007,In_1475,In_335);
nor U4008 (N_4008,In_231,In_617);
and U4009 (N_4009,In_944,In_1435);
and U4010 (N_4010,In_870,In_840);
nand U4011 (N_4011,In_1449,In_888);
nor U4012 (N_4012,In_1402,In_1370);
or U4013 (N_4013,In_317,In_1057);
and U4014 (N_4014,In_563,In_888);
nor U4015 (N_4015,In_1395,In_790);
or U4016 (N_4016,In_324,In_1061);
or U4017 (N_4017,In_559,In_3);
nor U4018 (N_4018,In_1061,In_1009);
or U4019 (N_4019,In_768,In_1286);
and U4020 (N_4020,In_104,In_726);
nand U4021 (N_4021,In_773,In_54);
nand U4022 (N_4022,In_1448,In_391);
or U4023 (N_4023,In_472,In_19);
or U4024 (N_4024,In_633,In_1132);
and U4025 (N_4025,In_1420,In_1111);
nor U4026 (N_4026,In_1265,In_1454);
nand U4027 (N_4027,In_1071,In_438);
and U4028 (N_4028,In_1121,In_91);
nand U4029 (N_4029,In_725,In_479);
or U4030 (N_4030,In_863,In_659);
nor U4031 (N_4031,In_840,In_156);
and U4032 (N_4032,In_656,In_804);
nand U4033 (N_4033,In_1492,In_1171);
and U4034 (N_4034,In_875,In_828);
nand U4035 (N_4035,In_423,In_1118);
nand U4036 (N_4036,In_1309,In_55);
nand U4037 (N_4037,In_1441,In_1461);
or U4038 (N_4038,In_194,In_1139);
nor U4039 (N_4039,In_1228,In_33);
and U4040 (N_4040,In_818,In_890);
nand U4041 (N_4041,In_505,In_446);
and U4042 (N_4042,In_589,In_1104);
nor U4043 (N_4043,In_523,In_342);
and U4044 (N_4044,In_1072,In_1337);
nand U4045 (N_4045,In_626,In_351);
and U4046 (N_4046,In_618,In_1493);
or U4047 (N_4047,In_689,In_869);
or U4048 (N_4048,In_1106,In_63);
or U4049 (N_4049,In_562,In_635);
or U4050 (N_4050,In_1421,In_144);
and U4051 (N_4051,In_464,In_358);
and U4052 (N_4052,In_1412,In_278);
nor U4053 (N_4053,In_333,In_175);
or U4054 (N_4054,In_1235,In_253);
nand U4055 (N_4055,In_1476,In_518);
or U4056 (N_4056,In_194,In_1116);
nand U4057 (N_4057,In_98,In_1211);
nor U4058 (N_4058,In_936,In_457);
nand U4059 (N_4059,In_1381,In_737);
nand U4060 (N_4060,In_337,In_11);
or U4061 (N_4061,In_567,In_1192);
or U4062 (N_4062,In_961,In_1241);
nor U4063 (N_4063,In_1017,In_546);
nor U4064 (N_4064,In_1275,In_901);
and U4065 (N_4065,In_1031,In_1004);
and U4066 (N_4066,In_834,In_183);
and U4067 (N_4067,In_1185,In_787);
nand U4068 (N_4068,In_505,In_1145);
nand U4069 (N_4069,In_125,In_301);
and U4070 (N_4070,In_817,In_834);
nor U4071 (N_4071,In_763,In_856);
xor U4072 (N_4072,In_51,In_1393);
and U4073 (N_4073,In_1139,In_498);
and U4074 (N_4074,In_960,In_135);
or U4075 (N_4075,In_963,In_344);
nor U4076 (N_4076,In_1378,In_1111);
nor U4077 (N_4077,In_554,In_622);
or U4078 (N_4078,In_573,In_1126);
nor U4079 (N_4079,In_455,In_997);
nand U4080 (N_4080,In_107,In_476);
and U4081 (N_4081,In_1465,In_557);
and U4082 (N_4082,In_564,In_1303);
nor U4083 (N_4083,In_1314,In_1158);
nor U4084 (N_4084,In_585,In_87);
or U4085 (N_4085,In_1455,In_155);
and U4086 (N_4086,In_619,In_738);
nand U4087 (N_4087,In_450,In_607);
nand U4088 (N_4088,In_179,In_230);
and U4089 (N_4089,In_450,In_519);
nor U4090 (N_4090,In_209,In_797);
and U4091 (N_4091,In_1025,In_598);
nor U4092 (N_4092,In_998,In_1371);
nand U4093 (N_4093,In_1393,In_537);
or U4094 (N_4094,In_1498,In_90);
nand U4095 (N_4095,In_1092,In_1330);
nor U4096 (N_4096,In_387,In_1062);
nand U4097 (N_4097,In_221,In_1027);
or U4098 (N_4098,In_852,In_1287);
or U4099 (N_4099,In_1428,In_798);
and U4100 (N_4100,In_392,In_896);
or U4101 (N_4101,In_403,In_1363);
and U4102 (N_4102,In_578,In_810);
and U4103 (N_4103,In_1496,In_300);
or U4104 (N_4104,In_858,In_1153);
and U4105 (N_4105,In_1411,In_378);
nor U4106 (N_4106,In_570,In_46);
and U4107 (N_4107,In_1260,In_864);
nand U4108 (N_4108,In_1401,In_351);
nor U4109 (N_4109,In_388,In_257);
nand U4110 (N_4110,In_1246,In_1314);
xnor U4111 (N_4111,In_171,In_727);
nor U4112 (N_4112,In_948,In_760);
or U4113 (N_4113,In_474,In_607);
and U4114 (N_4114,In_1400,In_1164);
and U4115 (N_4115,In_517,In_108);
and U4116 (N_4116,In_1221,In_991);
and U4117 (N_4117,In_728,In_1037);
or U4118 (N_4118,In_1466,In_533);
nand U4119 (N_4119,In_501,In_193);
nand U4120 (N_4120,In_1021,In_547);
and U4121 (N_4121,In_212,In_290);
nand U4122 (N_4122,In_1462,In_511);
nor U4123 (N_4123,In_1267,In_1140);
nor U4124 (N_4124,In_928,In_1283);
nor U4125 (N_4125,In_1193,In_1070);
nand U4126 (N_4126,In_260,In_8);
nand U4127 (N_4127,In_836,In_537);
or U4128 (N_4128,In_1318,In_73);
nor U4129 (N_4129,In_765,In_1334);
xnor U4130 (N_4130,In_362,In_862);
nand U4131 (N_4131,In_1398,In_560);
nand U4132 (N_4132,In_1343,In_770);
or U4133 (N_4133,In_170,In_345);
nor U4134 (N_4134,In_246,In_1070);
or U4135 (N_4135,In_437,In_1373);
or U4136 (N_4136,In_381,In_1478);
nor U4137 (N_4137,In_1389,In_1446);
nand U4138 (N_4138,In_976,In_442);
nor U4139 (N_4139,In_109,In_1107);
nand U4140 (N_4140,In_48,In_602);
nor U4141 (N_4141,In_293,In_1376);
and U4142 (N_4142,In_301,In_722);
nand U4143 (N_4143,In_846,In_853);
nor U4144 (N_4144,In_727,In_989);
nor U4145 (N_4145,In_1136,In_648);
nor U4146 (N_4146,In_144,In_211);
and U4147 (N_4147,In_712,In_203);
nor U4148 (N_4148,In_216,In_520);
nor U4149 (N_4149,In_1340,In_406);
nor U4150 (N_4150,In_345,In_935);
or U4151 (N_4151,In_147,In_808);
and U4152 (N_4152,In_210,In_995);
and U4153 (N_4153,In_668,In_628);
and U4154 (N_4154,In_1192,In_965);
or U4155 (N_4155,In_772,In_836);
nand U4156 (N_4156,In_509,In_1433);
nand U4157 (N_4157,In_1061,In_615);
or U4158 (N_4158,In_628,In_256);
nor U4159 (N_4159,In_14,In_112);
and U4160 (N_4160,In_1334,In_448);
nor U4161 (N_4161,In_825,In_322);
and U4162 (N_4162,In_1198,In_965);
or U4163 (N_4163,In_1068,In_822);
nor U4164 (N_4164,In_110,In_925);
nor U4165 (N_4165,In_1371,In_862);
and U4166 (N_4166,In_1343,In_1431);
or U4167 (N_4167,In_1456,In_1341);
and U4168 (N_4168,In_69,In_158);
or U4169 (N_4169,In_298,In_1360);
nand U4170 (N_4170,In_1465,In_880);
nor U4171 (N_4171,In_1336,In_346);
nor U4172 (N_4172,In_652,In_258);
nand U4173 (N_4173,In_92,In_1406);
nand U4174 (N_4174,In_327,In_1018);
or U4175 (N_4175,In_1307,In_956);
nand U4176 (N_4176,In_995,In_541);
nand U4177 (N_4177,In_343,In_165);
and U4178 (N_4178,In_390,In_1148);
or U4179 (N_4179,In_1395,In_652);
and U4180 (N_4180,In_435,In_185);
or U4181 (N_4181,In_1,In_249);
nor U4182 (N_4182,In_368,In_238);
or U4183 (N_4183,In_218,In_191);
and U4184 (N_4184,In_465,In_512);
nand U4185 (N_4185,In_1029,In_1304);
and U4186 (N_4186,In_1250,In_617);
nor U4187 (N_4187,In_395,In_43);
nor U4188 (N_4188,In_354,In_1273);
and U4189 (N_4189,In_843,In_1091);
nor U4190 (N_4190,In_1138,In_141);
nor U4191 (N_4191,In_832,In_1356);
or U4192 (N_4192,In_1447,In_1142);
and U4193 (N_4193,In_1375,In_59);
and U4194 (N_4194,In_913,In_1086);
nand U4195 (N_4195,In_813,In_442);
or U4196 (N_4196,In_1489,In_1058);
nor U4197 (N_4197,In_1040,In_1104);
nor U4198 (N_4198,In_739,In_833);
nor U4199 (N_4199,In_937,In_522);
and U4200 (N_4200,In_654,In_503);
nor U4201 (N_4201,In_184,In_263);
nand U4202 (N_4202,In_723,In_656);
nand U4203 (N_4203,In_64,In_100);
nand U4204 (N_4204,In_370,In_1023);
and U4205 (N_4205,In_165,In_1002);
nor U4206 (N_4206,In_314,In_446);
nand U4207 (N_4207,In_198,In_421);
and U4208 (N_4208,In_690,In_1299);
nand U4209 (N_4209,In_796,In_1365);
nand U4210 (N_4210,In_15,In_1179);
nor U4211 (N_4211,In_468,In_968);
nand U4212 (N_4212,In_892,In_176);
nand U4213 (N_4213,In_1098,In_309);
and U4214 (N_4214,In_1095,In_626);
and U4215 (N_4215,In_12,In_610);
nor U4216 (N_4216,In_896,In_578);
or U4217 (N_4217,In_987,In_1241);
nor U4218 (N_4218,In_365,In_58);
nor U4219 (N_4219,In_1123,In_257);
nand U4220 (N_4220,In_110,In_531);
and U4221 (N_4221,In_1463,In_815);
and U4222 (N_4222,In_354,In_509);
or U4223 (N_4223,In_1411,In_768);
nor U4224 (N_4224,In_631,In_1480);
nor U4225 (N_4225,In_1205,In_218);
or U4226 (N_4226,In_1158,In_1475);
and U4227 (N_4227,In_128,In_1192);
nor U4228 (N_4228,In_1392,In_645);
nand U4229 (N_4229,In_498,In_406);
and U4230 (N_4230,In_988,In_1288);
nor U4231 (N_4231,In_443,In_962);
nor U4232 (N_4232,In_467,In_1060);
nand U4233 (N_4233,In_932,In_1262);
nand U4234 (N_4234,In_619,In_967);
nand U4235 (N_4235,In_592,In_1243);
and U4236 (N_4236,In_719,In_1324);
and U4237 (N_4237,In_268,In_872);
nor U4238 (N_4238,In_273,In_145);
or U4239 (N_4239,In_1331,In_10);
nor U4240 (N_4240,In_114,In_901);
or U4241 (N_4241,In_53,In_1498);
and U4242 (N_4242,In_812,In_859);
or U4243 (N_4243,In_58,In_211);
or U4244 (N_4244,In_309,In_656);
nor U4245 (N_4245,In_1331,In_61);
or U4246 (N_4246,In_933,In_428);
nand U4247 (N_4247,In_1495,In_823);
or U4248 (N_4248,In_890,In_621);
nor U4249 (N_4249,In_1384,In_1028);
nand U4250 (N_4250,In_406,In_162);
nand U4251 (N_4251,In_1440,In_408);
nor U4252 (N_4252,In_636,In_393);
or U4253 (N_4253,In_871,In_437);
nand U4254 (N_4254,In_1343,In_39);
nand U4255 (N_4255,In_142,In_1067);
nand U4256 (N_4256,In_394,In_1184);
nand U4257 (N_4257,In_117,In_1430);
or U4258 (N_4258,In_325,In_1079);
or U4259 (N_4259,In_426,In_1);
or U4260 (N_4260,In_1366,In_65);
and U4261 (N_4261,In_1097,In_843);
nor U4262 (N_4262,In_1327,In_270);
and U4263 (N_4263,In_418,In_1275);
or U4264 (N_4264,In_1247,In_859);
nand U4265 (N_4265,In_823,In_1259);
and U4266 (N_4266,In_1265,In_756);
and U4267 (N_4267,In_552,In_410);
nand U4268 (N_4268,In_1279,In_744);
or U4269 (N_4269,In_1253,In_602);
and U4270 (N_4270,In_1249,In_368);
and U4271 (N_4271,In_889,In_546);
nor U4272 (N_4272,In_607,In_400);
nand U4273 (N_4273,In_303,In_138);
and U4274 (N_4274,In_809,In_394);
xor U4275 (N_4275,In_840,In_469);
or U4276 (N_4276,In_845,In_85);
nor U4277 (N_4277,In_1177,In_1091);
and U4278 (N_4278,In_1034,In_169);
nand U4279 (N_4279,In_1419,In_1213);
and U4280 (N_4280,In_619,In_144);
nand U4281 (N_4281,In_1405,In_1429);
nand U4282 (N_4282,In_1197,In_65);
nor U4283 (N_4283,In_534,In_1082);
or U4284 (N_4284,In_67,In_877);
nand U4285 (N_4285,In_410,In_894);
nand U4286 (N_4286,In_484,In_235);
or U4287 (N_4287,In_1397,In_873);
nand U4288 (N_4288,In_857,In_239);
and U4289 (N_4289,In_1140,In_456);
nor U4290 (N_4290,In_32,In_947);
nor U4291 (N_4291,In_690,In_63);
or U4292 (N_4292,In_47,In_230);
nor U4293 (N_4293,In_903,In_1131);
or U4294 (N_4294,In_1032,In_553);
or U4295 (N_4295,In_613,In_1261);
nor U4296 (N_4296,In_1386,In_979);
nand U4297 (N_4297,In_815,In_234);
nand U4298 (N_4298,In_1133,In_1085);
nor U4299 (N_4299,In_81,In_71);
and U4300 (N_4300,In_1153,In_438);
or U4301 (N_4301,In_990,In_517);
nand U4302 (N_4302,In_1154,In_256);
or U4303 (N_4303,In_70,In_338);
and U4304 (N_4304,In_1241,In_282);
nand U4305 (N_4305,In_3,In_978);
nor U4306 (N_4306,In_809,In_319);
nand U4307 (N_4307,In_978,In_861);
and U4308 (N_4308,In_293,In_551);
nor U4309 (N_4309,In_1016,In_702);
and U4310 (N_4310,In_556,In_282);
and U4311 (N_4311,In_556,In_1155);
nor U4312 (N_4312,In_891,In_415);
nand U4313 (N_4313,In_522,In_871);
nand U4314 (N_4314,In_1341,In_179);
and U4315 (N_4315,In_883,In_1476);
or U4316 (N_4316,In_1250,In_899);
nor U4317 (N_4317,In_332,In_144);
nand U4318 (N_4318,In_190,In_919);
nand U4319 (N_4319,In_275,In_463);
nor U4320 (N_4320,In_260,In_1361);
nor U4321 (N_4321,In_693,In_832);
nor U4322 (N_4322,In_85,In_614);
nor U4323 (N_4323,In_732,In_445);
nand U4324 (N_4324,In_1256,In_771);
nor U4325 (N_4325,In_230,In_403);
nand U4326 (N_4326,In_1112,In_559);
and U4327 (N_4327,In_437,In_855);
and U4328 (N_4328,In_653,In_1349);
and U4329 (N_4329,In_651,In_1161);
nor U4330 (N_4330,In_1293,In_1231);
nand U4331 (N_4331,In_24,In_458);
nand U4332 (N_4332,In_310,In_655);
nand U4333 (N_4333,In_403,In_1077);
or U4334 (N_4334,In_234,In_476);
nor U4335 (N_4335,In_374,In_1351);
nand U4336 (N_4336,In_1157,In_63);
or U4337 (N_4337,In_347,In_820);
or U4338 (N_4338,In_1076,In_538);
and U4339 (N_4339,In_138,In_1316);
or U4340 (N_4340,In_33,In_927);
and U4341 (N_4341,In_1148,In_210);
and U4342 (N_4342,In_528,In_417);
and U4343 (N_4343,In_834,In_865);
and U4344 (N_4344,In_310,In_787);
and U4345 (N_4345,In_989,In_1325);
xnor U4346 (N_4346,In_868,In_163);
nand U4347 (N_4347,In_669,In_486);
or U4348 (N_4348,In_772,In_1377);
and U4349 (N_4349,In_792,In_1075);
nor U4350 (N_4350,In_613,In_168);
nor U4351 (N_4351,In_527,In_1055);
nor U4352 (N_4352,In_1068,In_1399);
nand U4353 (N_4353,In_867,In_772);
and U4354 (N_4354,In_958,In_570);
and U4355 (N_4355,In_676,In_1405);
or U4356 (N_4356,In_1088,In_1474);
and U4357 (N_4357,In_680,In_1303);
or U4358 (N_4358,In_570,In_381);
nor U4359 (N_4359,In_671,In_764);
nor U4360 (N_4360,In_435,In_938);
and U4361 (N_4361,In_1004,In_1155);
and U4362 (N_4362,In_690,In_1298);
nand U4363 (N_4363,In_1374,In_241);
nor U4364 (N_4364,In_976,In_921);
nand U4365 (N_4365,In_1418,In_928);
or U4366 (N_4366,In_1221,In_1297);
nand U4367 (N_4367,In_1400,In_516);
nor U4368 (N_4368,In_1120,In_1118);
nor U4369 (N_4369,In_456,In_1231);
and U4370 (N_4370,In_1404,In_553);
and U4371 (N_4371,In_208,In_1194);
and U4372 (N_4372,In_55,In_225);
and U4373 (N_4373,In_134,In_478);
nor U4374 (N_4374,In_7,In_1198);
or U4375 (N_4375,In_342,In_318);
nor U4376 (N_4376,In_271,In_1401);
or U4377 (N_4377,In_602,In_1463);
nor U4378 (N_4378,In_1460,In_902);
and U4379 (N_4379,In_1047,In_1224);
nand U4380 (N_4380,In_308,In_46);
and U4381 (N_4381,In_125,In_77);
nor U4382 (N_4382,In_246,In_870);
or U4383 (N_4383,In_1208,In_1196);
or U4384 (N_4384,In_1371,In_19);
and U4385 (N_4385,In_634,In_1059);
or U4386 (N_4386,In_1249,In_497);
nand U4387 (N_4387,In_24,In_1204);
nor U4388 (N_4388,In_73,In_297);
and U4389 (N_4389,In_947,In_787);
nor U4390 (N_4390,In_168,In_405);
or U4391 (N_4391,In_1295,In_992);
nand U4392 (N_4392,In_857,In_54);
nand U4393 (N_4393,In_1166,In_307);
or U4394 (N_4394,In_1283,In_1399);
nor U4395 (N_4395,In_193,In_1156);
or U4396 (N_4396,In_3,In_691);
and U4397 (N_4397,In_302,In_1239);
nand U4398 (N_4398,In_519,In_1174);
nor U4399 (N_4399,In_213,In_1010);
nor U4400 (N_4400,In_117,In_312);
nor U4401 (N_4401,In_1418,In_312);
nand U4402 (N_4402,In_1442,In_471);
nor U4403 (N_4403,In_124,In_1301);
nand U4404 (N_4404,In_563,In_468);
and U4405 (N_4405,In_614,In_517);
or U4406 (N_4406,In_231,In_594);
nor U4407 (N_4407,In_747,In_299);
or U4408 (N_4408,In_18,In_1073);
and U4409 (N_4409,In_1303,In_93);
or U4410 (N_4410,In_1131,In_1382);
nor U4411 (N_4411,In_1065,In_939);
and U4412 (N_4412,In_1491,In_289);
nand U4413 (N_4413,In_457,In_915);
nor U4414 (N_4414,In_343,In_62);
or U4415 (N_4415,In_902,In_167);
and U4416 (N_4416,In_681,In_173);
or U4417 (N_4417,In_941,In_1249);
and U4418 (N_4418,In_933,In_879);
nor U4419 (N_4419,In_349,In_453);
or U4420 (N_4420,In_1039,In_1360);
nor U4421 (N_4421,In_818,In_1144);
and U4422 (N_4422,In_1208,In_906);
or U4423 (N_4423,In_1470,In_765);
and U4424 (N_4424,In_504,In_26);
nor U4425 (N_4425,In_853,In_763);
or U4426 (N_4426,In_511,In_1324);
nor U4427 (N_4427,In_992,In_291);
nor U4428 (N_4428,In_1120,In_1262);
nor U4429 (N_4429,In_1274,In_158);
nor U4430 (N_4430,In_1076,In_1426);
and U4431 (N_4431,In_629,In_1215);
nand U4432 (N_4432,In_983,In_1309);
nand U4433 (N_4433,In_963,In_71);
and U4434 (N_4434,In_596,In_1225);
nor U4435 (N_4435,In_245,In_51);
nand U4436 (N_4436,In_400,In_1045);
nand U4437 (N_4437,In_439,In_816);
nor U4438 (N_4438,In_43,In_1135);
xor U4439 (N_4439,In_1415,In_1058);
nor U4440 (N_4440,In_449,In_469);
xnor U4441 (N_4441,In_478,In_590);
nor U4442 (N_4442,In_1435,In_1086);
and U4443 (N_4443,In_1394,In_107);
nand U4444 (N_4444,In_1060,In_340);
nand U4445 (N_4445,In_1420,In_799);
nor U4446 (N_4446,In_963,In_916);
and U4447 (N_4447,In_915,In_786);
and U4448 (N_4448,In_656,In_1179);
nor U4449 (N_4449,In_1019,In_1297);
or U4450 (N_4450,In_958,In_703);
or U4451 (N_4451,In_105,In_494);
nand U4452 (N_4452,In_1048,In_280);
and U4453 (N_4453,In_1156,In_816);
nor U4454 (N_4454,In_293,In_930);
or U4455 (N_4455,In_1205,In_542);
or U4456 (N_4456,In_1108,In_1115);
nand U4457 (N_4457,In_1280,In_798);
or U4458 (N_4458,In_1440,In_1420);
nand U4459 (N_4459,In_328,In_131);
nor U4460 (N_4460,In_988,In_1325);
or U4461 (N_4461,In_1466,In_9);
nand U4462 (N_4462,In_158,In_232);
xnor U4463 (N_4463,In_545,In_1242);
nor U4464 (N_4464,In_252,In_1104);
nand U4465 (N_4465,In_1360,In_259);
or U4466 (N_4466,In_461,In_1387);
nand U4467 (N_4467,In_360,In_1322);
nor U4468 (N_4468,In_715,In_1009);
nand U4469 (N_4469,In_142,In_987);
nand U4470 (N_4470,In_1196,In_10);
nand U4471 (N_4471,In_132,In_69);
and U4472 (N_4472,In_1308,In_1244);
and U4473 (N_4473,In_1245,In_1492);
and U4474 (N_4474,In_429,In_621);
nand U4475 (N_4475,In_647,In_365);
nor U4476 (N_4476,In_1355,In_1016);
and U4477 (N_4477,In_1139,In_902);
and U4478 (N_4478,In_74,In_727);
nand U4479 (N_4479,In_1029,In_631);
and U4480 (N_4480,In_268,In_373);
nor U4481 (N_4481,In_254,In_419);
nor U4482 (N_4482,In_1292,In_254);
or U4483 (N_4483,In_203,In_678);
and U4484 (N_4484,In_1353,In_1167);
and U4485 (N_4485,In_604,In_1086);
nor U4486 (N_4486,In_1025,In_1331);
nor U4487 (N_4487,In_210,In_627);
and U4488 (N_4488,In_530,In_703);
and U4489 (N_4489,In_79,In_451);
nand U4490 (N_4490,In_384,In_224);
and U4491 (N_4491,In_345,In_297);
and U4492 (N_4492,In_1364,In_1115);
nor U4493 (N_4493,In_1333,In_581);
nand U4494 (N_4494,In_985,In_854);
or U4495 (N_4495,In_1080,In_1404);
nand U4496 (N_4496,In_291,In_1205);
and U4497 (N_4497,In_635,In_982);
xnor U4498 (N_4498,In_462,In_1021);
or U4499 (N_4499,In_1456,In_351);
and U4500 (N_4500,In_761,In_1493);
and U4501 (N_4501,In_1043,In_1471);
nor U4502 (N_4502,In_1467,In_443);
or U4503 (N_4503,In_39,In_1061);
and U4504 (N_4504,In_829,In_293);
nor U4505 (N_4505,In_1416,In_1088);
or U4506 (N_4506,In_516,In_1205);
nor U4507 (N_4507,In_563,In_1441);
and U4508 (N_4508,In_203,In_155);
nand U4509 (N_4509,In_1300,In_45);
nor U4510 (N_4510,In_1481,In_931);
xor U4511 (N_4511,In_318,In_191);
and U4512 (N_4512,In_520,In_550);
or U4513 (N_4513,In_1437,In_985);
nand U4514 (N_4514,In_1436,In_171);
nor U4515 (N_4515,In_47,In_108);
or U4516 (N_4516,In_189,In_699);
xor U4517 (N_4517,In_937,In_885);
nand U4518 (N_4518,In_1449,In_93);
or U4519 (N_4519,In_956,In_656);
nand U4520 (N_4520,In_879,In_808);
and U4521 (N_4521,In_1267,In_297);
and U4522 (N_4522,In_1003,In_1299);
and U4523 (N_4523,In_535,In_496);
nand U4524 (N_4524,In_803,In_336);
or U4525 (N_4525,In_378,In_937);
or U4526 (N_4526,In_1295,In_295);
or U4527 (N_4527,In_1474,In_1283);
or U4528 (N_4528,In_35,In_416);
or U4529 (N_4529,In_303,In_920);
and U4530 (N_4530,In_1173,In_679);
nand U4531 (N_4531,In_571,In_612);
and U4532 (N_4532,In_1482,In_1126);
xor U4533 (N_4533,In_414,In_1445);
xor U4534 (N_4534,In_1302,In_35);
or U4535 (N_4535,In_668,In_1009);
or U4536 (N_4536,In_698,In_597);
nand U4537 (N_4537,In_605,In_369);
and U4538 (N_4538,In_85,In_1312);
or U4539 (N_4539,In_1286,In_526);
nand U4540 (N_4540,In_669,In_1169);
nand U4541 (N_4541,In_576,In_278);
or U4542 (N_4542,In_769,In_707);
nor U4543 (N_4543,In_539,In_877);
nor U4544 (N_4544,In_614,In_1465);
and U4545 (N_4545,In_1333,In_127);
or U4546 (N_4546,In_320,In_66);
nand U4547 (N_4547,In_871,In_1127);
or U4548 (N_4548,In_567,In_68);
nand U4549 (N_4549,In_282,In_814);
nor U4550 (N_4550,In_232,In_600);
and U4551 (N_4551,In_904,In_762);
nor U4552 (N_4552,In_215,In_1354);
nand U4553 (N_4553,In_1150,In_1065);
or U4554 (N_4554,In_545,In_585);
nor U4555 (N_4555,In_906,In_788);
xnor U4556 (N_4556,In_182,In_895);
nand U4557 (N_4557,In_1336,In_1044);
nor U4558 (N_4558,In_1029,In_187);
nand U4559 (N_4559,In_1265,In_60);
nand U4560 (N_4560,In_1119,In_89);
or U4561 (N_4561,In_136,In_395);
nand U4562 (N_4562,In_871,In_819);
or U4563 (N_4563,In_443,In_679);
nand U4564 (N_4564,In_1066,In_1288);
and U4565 (N_4565,In_930,In_703);
and U4566 (N_4566,In_1127,In_1495);
nor U4567 (N_4567,In_806,In_924);
and U4568 (N_4568,In_793,In_1212);
or U4569 (N_4569,In_1190,In_1138);
and U4570 (N_4570,In_1131,In_1431);
nor U4571 (N_4571,In_330,In_1332);
nor U4572 (N_4572,In_1227,In_1099);
nor U4573 (N_4573,In_1159,In_1486);
or U4574 (N_4574,In_1207,In_301);
or U4575 (N_4575,In_1354,In_484);
or U4576 (N_4576,In_802,In_878);
and U4577 (N_4577,In_588,In_624);
nor U4578 (N_4578,In_1197,In_1265);
nand U4579 (N_4579,In_223,In_257);
nand U4580 (N_4580,In_1462,In_1023);
nand U4581 (N_4581,In_893,In_1496);
nand U4582 (N_4582,In_4,In_1217);
nand U4583 (N_4583,In_121,In_1031);
or U4584 (N_4584,In_15,In_1225);
nand U4585 (N_4585,In_1199,In_373);
nand U4586 (N_4586,In_1461,In_415);
or U4587 (N_4587,In_137,In_1485);
nand U4588 (N_4588,In_1408,In_686);
nor U4589 (N_4589,In_440,In_99);
nor U4590 (N_4590,In_953,In_1143);
nor U4591 (N_4591,In_78,In_842);
nand U4592 (N_4592,In_949,In_734);
nand U4593 (N_4593,In_1478,In_690);
or U4594 (N_4594,In_462,In_900);
and U4595 (N_4595,In_413,In_1456);
xnor U4596 (N_4596,In_658,In_1351);
and U4597 (N_4597,In_1093,In_969);
or U4598 (N_4598,In_906,In_766);
or U4599 (N_4599,In_672,In_1401);
and U4600 (N_4600,In_1498,In_945);
and U4601 (N_4601,In_1380,In_221);
and U4602 (N_4602,In_980,In_619);
and U4603 (N_4603,In_226,In_862);
or U4604 (N_4604,In_688,In_1110);
xor U4605 (N_4605,In_377,In_984);
nand U4606 (N_4606,In_1106,In_367);
and U4607 (N_4607,In_472,In_445);
or U4608 (N_4608,In_1406,In_417);
or U4609 (N_4609,In_71,In_1305);
or U4610 (N_4610,In_1279,In_107);
or U4611 (N_4611,In_125,In_36);
or U4612 (N_4612,In_722,In_580);
and U4613 (N_4613,In_1268,In_1105);
and U4614 (N_4614,In_354,In_1214);
or U4615 (N_4615,In_288,In_832);
or U4616 (N_4616,In_650,In_143);
nor U4617 (N_4617,In_432,In_890);
or U4618 (N_4618,In_1004,In_1089);
and U4619 (N_4619,In_705,In_1135);
nand U4620 (N_4620,In_388,In_972);
nor U4621 (N_4621,In_200,In_1482);
and U4622 (N_4622,In_1011,In_440);
xor U4623 (N_4623,In_1363,In_1496);
and U4624 (N_4624,In_660,In_1045);
and U4625 (N_4625,In_42,In_575);
or U4626 (N_4626,In_771,In_290);
and U4627 (N_4627,In_227,In_1388);
nand U4628 (N_4628,In_1347,In_493);
and U4629 (N_4629,In_302,In_1009);
or U4630 (N_4630,In_1192,In_16);
nor U4631 (N_4631,In_1418,In_511);
or U4632 (N_4632,In_576,In_1498);
and U4633 (N_4633,In_1394,In_958);
nor U4634 (N_4634,In_71,In_1492);
nor U4635 (N_4635,In_768,In_30);
nor U4636 (N_4636,In_1419,In_147);
and U4637 (N_4637,In_1284,In_1382);
or U4638 (N_4638,In_779,In_74);
nor U4639 (N_4639,In_920,In_768);
or U4640 (N_4640,In_69,In_62);
nand U4641 (N_4641,In_1216,In_795);
or U4642 (N_4642,In_441,In_1003);
and U4643 (N_4643,In_793,In_1424);
and U4644 (N_4644,In_267,In_684);
nand U4645 (N_4645,In_298,In_801);
nand U4646 (N_4646,In_1337,In_44);
nor U4647 (N_4647,In_346,In_349);
nand U4648 (N_4648,In_603,In_1328);
or U4649 (N_4649,In_1158,In_1291);
xnor U4650 (N_4650,In_204,In_192);
and U4651 (N_4651,In_1148,In_543);
and U4652 (N_4652,In_157,In_1050);
nor U4653 (N_4653,In_916,In_411);
or U4654 (N_4654,In_982,In_44);
nor U4655 (N_4655,In_104,In_203);
nor U4656 (N_4656,In_1463,In_1479);
or U4657 (N_4657,In_1398,In_179);
nand U4658 (N_4658,In_888,In_198);
nand U4659 (N_4659,In_30,In_166);
nor U4660 (N_4660,In_557,In_1203);
nand U4661 (N_4661,In_1077,In_570);
or U4662 (N_4662,In_210,In_988);
or U4663 (N_4663,In_1151,In_1161);
nand U4664 (N_4664,In_247,In_0);
nand U4665 (N_4665,In_219,In_488);
nand U4666 (N_4666,In_415,In_145);
or U4667 (N_4667,In_945,In_276);
and U4668 (N_4668,In_579,In_233);
nor U4669 (N_4669,In_788,In_1400);
nor U4670 (N_4670,In_1250,In_711);
nand U4671 (N_4671,In_794,In_1279);
and U4672 (N_4672,In_309,In_1291);
nor U4673 (N_4673,In_257,In_654);
and U4674 (N_4674,In_943,In_91);
xor U4675 (N_4675,In_1243,In_33);
nand U4676 (N_4676,In_579,In_1233);
and U4677 (N_4677,In_610,In_814);
nand U4678 (N_4678,In_633,In_1032);
or U4679 (N_4679,In_557,In_50);
and U4680 (N_4680,In_67,In_926);
nand U4681 (N_4681,In_55,In_444);
nand U4682 (N_4682,In_1484,In_703);
nor U4683 (N_4683,In_500,In_298);
or U4684 (N_4684,In_463,In_705);
and U4685 (N_4685,In_750,In_1003);
nand U4686 (N_4686,In_361,In_137);
or U4687 (N_4687,In_64,In_397);
and U4688 (N_4688,In_264,In_223);
nand U4689 (N_4689,In_354,In_503);
or U4690 (N_4690,In_359,In_1430);
and U4691 (N_4691,In_233,In_51);
nand U4692 (N_4692,In_177,In_436);
nand U4693 (N_4693,In_1450,In_813);
and U4694 (N_4694,In_1358,In_1136);
or U4695 (N_4695,In_722,In_796);
nand U4696 (N_4696,In_292,In_1365);
nand U4697 (N_4697,In_563,In_1217);
nand U4698 (N_4698,In_4,In_1321);
or U4699 (N_4699,In_942,In_640);
nand U4700 (N_4700,In_1457,In_715);
nand U4701 (N_4701,In_522,In_298);
nor U4702 (N_4702,In_625,In_135);
or U4703 (N_4703,In_1269,In_215);
xnor U4704 (N_4704,In_240,In_1244);
nand U4705 (N_4705,In_1046,In_422);
and U4706 (N_4706,In_929,In_838);
nor U4707 (N_4707,In_1087,In_1140);
or U4708 (N_4708,In_91,In_451);
nor U4709 (N_4709,In_633,In_386);
nand U4710 (N_4710,In_147,In_57);
nor U4711 (N_4711,In_747,In_1050);
and U4712 (N_4712,In_526,In_1337);
and U4713 (N_4713,In_863,In_884);
and U4714 (N_4714,In_481,In_116);
or U4715 (N_4715,In_836,In_458);
nor U4716 (N_4716,In_1170,In_73);
or U4717 (N_4717,In_1477,In_1180);
or U4718 (N_4718,In_351,In_66);
and U4719 (N_4719,In_1019,In_106);
or U4720 (N_4720,In_978,In_255);
nand U4721 (N_4721,In_560,In_599);
or U4722 (N_4722,In_83,In_1499);
nor U4723 (N_4723,In_699,In_596);
nand U4724 (N_4724,In_949,In_1147);
or U4725 (N_4725,In_338,In_83);
or U4726 (N_4726,In_1146,In_215);
and U4727 (N_4727,In_1062,In_1010);
or U4728 (N_4728,In_1233,In_165);
nand U4729 (N_4729,In_102,In_798);
nand U4730 (N_4730,In_490,In_754);
or U4731 (N_4731,In_76,In_784);
nor U4732 (N_4732,In_244,In_1455);
nand U4733 (N_4733,In_430,In_835);
nor U4734 (N_4734,In_727,In_1287);
or U4735 (N_4735,In_162,In_869);
nor U4736 (N_4736,In_950,In_472);
nand U4737 (N_4737,In_1250,In_60);
nor U4738 (N_4738,In_317,In_510);
nand U4739 (N_4739,In_1057,In_292);
nand U4740 (N_4740,In_522,In_217);
nor U4741 (N_4741,In_149,In_490);
nor U4742 (N_4742,In_462,In_693);
or U4743 (N_4743,In_1299,In_1099);
nand U4744 (N_4744,In_77,In_1033);
and U4745 (N_4745,In_951,In_350);
or U4746 (N_4746,In_301,In_850);
and U4747 (N_4747,In_1336,In_1153);
nand U4748 (N_4748,In_560,In_572);
and U4749 (N_4749,In_752,In_978);
and U4750 (N_4750,In_1180,In_71);
and U4751 (N_4751,In_263,In_1304);
or U4752 (N_4752,In_1312,In_1383);
and U4753 (N_4753,In_1239,In_396);
nor U4754 (N_4754,In_598,In_632);
or U4755 (N_4755,In_352,In_524);
nor U4756 (N_4756,In_131,In_909);
or U4757 (N_4757,In_1440,In_769);
and U4758 (N_4758,In_1299,In_1100);
nor U4759 (N_4759,In_1364,In_1343);
nand U4760 (N_4760,In_579,In_578);
and U4761 (N_4761,In_1094,In_751);
or U4762 (N_4762,In_1184,In_48);
and U4763 (N_4763,In_1179,In_321);
nor U4764 (N_4764,In_977,In_366);
or U4765 (N_4765,In_854,In_698);
nor U4766 (N_4766,In_496,In_871);
and U4767 (N_4767,In_827,In_1187);
and U4768 (N_4768,In_193,In_1223);
nor U4769 (N_4769,In_684,In_247);
nor U4770 (N_4770,In_1212,In_573);
nor U4771 (N_4771,In_793,In_990);
nand U4772 (N_4772,In_640,In_709);
nand U4773 (N_4773,In_60,In_65);
or U4774 (N_4774,In_983,In_398);
xor U4775 (N_4775,In_1351,In_1017);
nor U4776 (N_4776,In_1487,In_961);
and U4777 (N_4777,In_1291,In_200);
nand U4778 (N_4778,In_1422,In_59);
or U4779 (N_4779,In_103,In_689);
or U4780 (N_4780,In_964,In_173);
nor U4781 (N_4781,In_680,In_458);
and U4782 (N_4782,In_757,In_845);
and U4783 (N_4783,In_1348,In_1478);
nand U4784 (N_4784,In_1222,In_183);
nor U4785 (N_4785,In_446,In_982);
nand U4786 (N_4786,In_716,In_1179);
and U4787 (N_4787,In_400,In_1202);
nor U4788 (N_4788,In_485,In_1118);
nor U4789 (N_4789,In_441,In_912);
and U4790 (N_4790,In_1080,In_781);
nand U4791 (N_4791,In_1072,In_739);
or U4792 (N_4792,In_383,In_1363);
nor U4793 (N_4793,In_1467,In_1172);
and U4794 (N_4794,In_1023,In_445);
nor U4795 (N_4795,In_701,In_600);
or U4796 (N_4796,In_748,In_1221);
and U4797 (N_4797,In_0,In_171);
and U4798 (N_4798,In_1383,In_912);
nor U4799 (N_4799,In_322,In_789);
or U4800 (N_4800,In_1120,In_1145);
nor U4801 (N_4801,In_286,In_291);
or U4802 (N_4802,In_858,In_1176);
nor U4803 (N_4803,In_1457,In_1260);
or U4804 (N_4804,In_754,In_1221);
nand U4805 (N_4805,In_713,In_267);
or U4806 (N_4806,In_107,In_965);
or U4807 (N_4807,In_1100,In_378);
and U4808 (N_4808,In_668,In_765);
nand U4809 (N_4809,In_797,In_1355);
and U4810 (N_4810,In_1033,In_1477);
nand U4811 (N_4811,In_373,In_1387);
nor U4812 (N_4812,In_1324,In_942);
nand U4813 (N_4813,In_1251,In_788);
nor U4814 (N_4814,In_621,In_715);
nand U4815 (N_4815,In_439,In_140);
or U4816 (N_4816,In_1439,In_246);
or U4817 (N_4817,In_733,In_1052);
and U4818 (N_4818,In_1107,In_396);
nand U4819 (N_4819,In_538,In_22);
or U4820 (N_4820,In_1385,In_179);
or U4821 (N_4821,In_8,In_634);
or U4822 (N_4822,In_234,In_256);
or U4823 (N_4823,In_833,In_499);
nand U4824 (N_4824,In_1104,In_1315);
or U4825 (N_4825,In_611,In_644);
and U4826 (N_4826,In_498,In_1417);
nor U4827 (N_4827,In_228,In_1388);
nor U4828 (N_4828,In_162,In_739);
and U4829 (N_4829,In_1020,In_434);
nand U4830 (N_4830,In_674,In_26);
nor U4831 (N_4831,In_1156,In_536);
and U4832 (N_4832,In_1417,In_1392);
and U4833 (N_4833,In_136,In_1225);
and U4834 (N_4834,In_332,In_1273);
nand U4835 (N_4835,In_329,In_730);
xnor U4836 (N_4836,In_532,In_676);
or U4837 (N_4837,In_1116,In_238);
and U4838 (N_4838,In_902,In_698);
nor U4839 (N_4839,In_267,In_714);
nor U4840 (N_4840,In_44,In_838);
and U4841 (N_4841,In_763,In_6);
and U4842 (N_4842,In_320,In_124);
and U4843 (N_4843,In_1154,In_263);
and U4844 (N_4844,In_996,In_809);
and U4845 (N_4845,In_923,In_72);
or U4846 (N_4846,In_1469,In_1021);
nor U4847 (N_4847,In_132,In_66);
nand U4848 (N_4848,In_248,In_720);
nand U4849 (N_4849,In_13,In_230);
nor U4850 (N_4850,In_1241,In_1489);
nor U4851 (N_4851,In_478,In_1142);
and U4852 (N_4852,In_179,In_438);
and U4853 (N_4853,In_867,In_420);
and U4854 (N_4854,In_1006,In_217);
nor U4855 (N_4855,In_475,In_1458);
nor U4856 (N_4856,In_1398,In_450);
nand U4857 (N_4857,In_58,In_1026);
nand U4858 (N_4858,In_1139,In_1029);
xnor U4859 (N_4859,In_463,In_580);
or U4860 (N_4860,In_785,In_1189);
or U4861 (N_4861,In_201,In_978);
or U4862 (N_4862,In_1399,In_839);
nor U4863 (N_4863,In_716,In_420);
nor U4864 (N_4864,In_1410,In_747);
or U4865 (N_4865,In_1180,In_1087);
or U4866 (N_4866,In_295,In_714);
and U4867 (N_4867,In_224,In_176);
and U4868 (N_4868,In_32,In_350);
or U4869 (N_4869,In_341,In_1094);
or U4870 (N_4870,In_1057,In_949);
nor U4871 (N_4871,In_743,In_65);
nand U4872 (N_4872,In_983,In_593);
and U4873 (N_4873,In_171,In_972);
nor U4874 (N_4874,In_1128,In_1015);
nor U4875 (N_4875,In_1090,In_1261);
nor U4876 (N_4876,In_812,In_1017);
or U4877 (N_4877,In_925,In_1056);
nand U4878 (N_4878,In_1438,In_1093);
and U4879 (N_4879,In_1247,In_150);
and U4880 (N_4880,In_710,In_393);
and U4881 (N_4881,In_1461,In_1124);
nor U4882 (N_4882,In_1176,In_776);
or U4883 (N_4883,In_500,In_486);
nand U4884 (N_4884,In_1305,In_842);
nor U4885 (N_4885,In_656,In_26);
nor U4886 (N_4886,In_1117,In_485);
or U4887 (N_4887,In_564,In_386);
or U4888 (N_4888,In_933,In_781);
nand U4889 (N_4889,In_1464,In_345);
nor U4890 (N_4890,In_1233,In_1187);
or U4891 (N_4891,In_980,In_1419);
and U4892 (N_4892,In_1160,In_1354);
nand U4893 (N_4893,In_927,In_219);
and U4894 (N_4894,In_302,In_1300);
nand U4895 (N_4895,In_1193,In_641);
or U4896 (N_4896,In_689,In_95);
nor U4897 (N_4897,In_537,In_1031);
and U4898 (N_4898,In_917,In_284);
and U4899 (N_4899,In_707,In_401);
and U4900 (N_4900,In_507,In_1197);
nor U4901 (N_4901,In_1174,In_95);
or U4902 (N_4902,In_1069,In_101);
nand U4903 (N_4903,In_717,In_293);
nand U4904 (N_4904,In_89,In_913);
nand U4905 (N_4905,In_432,In_650);
and U4906 (N_4906,In_504,In_940);
nand U4907 (N_4907,In_1388,In_283);
or U4908 (N_4908,In_1132,In_245);
nand U4909 (N_4909,In_1478,In_922);
or U4910 (N_4910,In_1278,In_1030);
and U4911 (N_4911,In_1005,In_262);
and U4912 (N_4912,In_1372,In_762);
and U4913 (N_4913,In_864,In_208);
nand U4914 (N_4914,In_1073,In_975);
and U4915 (N_4915,In_210,In_680);
and U4916 (N_4916,In_1457,In_342);
nand U4917 (N_4917,In_561,In_323);
nand U4918 (N_4918,In_1051,In_888);
or U4919 (N_4919,In_1466,In_255);
nand U4920 (N_4920,In_460,In_135);
or U4921 (N_4921,In_323,In_611);
nand U4922 (N_4922,In_1134,In_461);
and U4923 (N_4923,In_1323,In_198);
nand U4924 (N_4924,In_899,In_648);
nand U4925 (N_4925,In_537,In_1370);
nand U4926 (N_4926,In_33,In_241);
and U4927 (N_4927,In_1316,In_120);
nand U4928 (N_4928,In_291,In_44);
nand U4929 (N_4929,In_281,In_626);
or U4930 (N_4930,In_879,In_47);
nor U4931 (N_4931,In_995,In_224);
nor U4932 (N_4932,In_1414,In_1330);
or U4933 (N_4933,In_1393,In_1449);
and U4934 (N_4934,In_782,In_568);
nor U4935 (N_4935,In_373,In_723);
or U4936 (N_4936,In_402,In_73);
nand U4937 (N_4937,In_676,In_49);
nand U4938 (N_4938,In_1002,In_867);
nor U4939 (N_4939,In_524,In_121);
nand U4940 (N_4940,In_1301,In_1446);
and U4941 (N_4941,In_1179,In_323);
or U4942 (N_4942,In_1428,In_892);
nor U4943 (N_4943,In_791,In_978);
and U4944 (N_4944,In_169,In_307);
or U4945 (N_4945,In_1271,In_567);
and U4946 (N_4946,In_10,In_490);
nor U4947 (N_4947,In_858,In_1228);
and U4948 (N_4948,In_1267,In_309);
or U4949 (N_4949,In_1110,In_562);
and U4950 (N_4950,In_913,In_1139);
or U4951 (N_4951,In_1410,In_1044);
nand U4952 (N_4952,In_1046,In_402);
nor U4953 (N_4953,In_1454,In_806);
nor U4954 (N_4954,In_1086,In_840);
nor U4955 (N_4955,In_1340,In_184);
nor U4956 (N_4956,In_1271,In_914);
nor U4957 (N_4957,In_875,In_713);
or U4958 (N_4958,In_405,In_983);
nand U4959 (N_4959,In_1042,In_1172);
and U4960 (N_4960,In_955,In_531);
or U4961 (N_4961,In_1463,In_649);
and U4962 (N_4962,In_1078,In_955);
nand U4963 (N_4963,In_973,In_700);
nor U4964 (N_4964,In_270,In_1390);
nor U4965 (N_4965,In_810,In_73);
nand U4966 (N_4966,In_934,In_81);
and U4967 (N_4967,In_1336,In_48);
nand U4968 (N_4968,In_605,In_207);
nor U4969 (N_4969,In_1062,In_907);
and U4970 (N_4970,In_1027,In_939);
nor U4971 (N_4971,In_79,In_12);
and U4972 (N_4972,In_462,In_601);
nand U4973 (N_4973,In_1145,In_40);
nand U4974 (N_4974,In_1166,In_1070);
or U4975 (N_4975,In_1403,In_851);
nor U4976 (N_4976,In_203,In_312);
nor U4977 (N_4977,In_1122,In_1165);
and U4978 (N_4978,In_1103,In_416);
or U4979 (N_4979,In_1055,In_1162);
and U4980 (N_4980,In_1325,In_686);
or U4981 (N_4981,In_279,In_630);
nand U4982 (N_4982,In_1082,In_1208);
nand U4983 (N_4983,In_958,In_1481);
and U4984 (N_4984,In_696,In_681);
and U4985 (N_4985,In_1017,In_827);
nor U4986 (N_4986,In_976,In_449);
or U4987 (N_4987,In_1365,In_1072);
and U4988 (N_4988,In_1050,In_1052);
and U4989 (N_4989,In_280,In_509);
nand U4990 (N_4990,In_403,In_709);
nand U4991 (N_4991,In_926,In_222);
and U4992 (N_4992,In_1236,In_1058);
or U4993 (N_4993,In_1152,In_171);
and U4994 (N_4994,In_622,In_757);
nand U4995 (N_4995,In_991,In_1289);
nor U4996 (N_4996,In_707,In_720);
or U4997 (N_4997,In_297,In_259);
nand U4998 (N_4998,In_1183,In_39);
nand U4999 (N_4999,In_444,In_125);
nand U5000 (N_5000,N_39,N_3216);
or U5001 (N_5001,N_2112,N_2612);
or U5002 (N_5002,N_3855,N_547);
nor U5003 (N_5003,N_868,N_4403);
nand U5004 (N_5004,N_2330,N_518);
nor U5005 (N_5005,N_3009,N_3564);
nand U5006 (N_5006,N_4012,N_1401);
or U5007 (N_5007,N_4010,N_1872);
or U5008 (N_5008,N_630,N_3360);
and U5009 (N_5009,N_4570,N_186);
nor U5010 (N_5010,N_914,N_2278);
or U5011 (N_5011,N_3272,N_1357);
nand U5012 (N_5012,N_309,N_3132);
and U5013 (N_5013,N_2656,N_2782);
or U5014 (N_5014,N_2650,N_610);
and U5015 (N_5015,N_784,N_626);
nor U5016 (N_5016,N_4406,N_877);
and U5017 (N_5017,N_2897,N_3143);
and U5018 (N_5018,N_4522,N_1721);
or U5019 (N_5019,N_1536,N_4722);
or U5020 (N_5020,N_4930,N_3575);
nand U5021 (N_5021,N_75,N_1430);
and U5022 (N_5022,N_3354,N_1085);
and U5023 (N_5023,N_4299,N_4230);
or U5024 (N_5024,N_4197,N_223);
and U5025 (N_5025,N_1834,N_3805);
nand U5026 (N_5026,N_1545,N_1528);
or U5027 (N_5027,N_4467,N_2580);
and U5028 (N_5028,N_1628,N_4666);
nor U5029 (N_5029,N_2424,N_1347);
and U5030 (N_5030,N_1437,N_3246);
or U5031 (N_5031,N_2592,N_3980);
nand U5032 (N_5032,N_1622,N_1425);
or U5033 (N_5033,N_632,N_2118);
nand U5034 (N_5034,N_3638,N_4645);
nor U5035 (N_5035,N_362,N_3522);
or U5036 (N_5036,N_2039,N_3134);
and U5037 (N_5037,N_4983,N_1658);
nand U5038 (N_5038,N_1514,N_1712);
and U5039 (N_5039,N_2637,N_4968);
and U5040 (N_5040,N_4946,N_915);
or U5041 (N_5041,N_664,N_3932);
and U5042 (N_5042,N_3150,N_1144);
or U5043 (N_5043,N_2335,N_2326);
nor U5044 (N_5044,N_4650,N_1064);
and U5045 (N_5045,N_4380,N_1975);
or U5046 (N_5046,N_3,N_2657);
and U5047 (N_5047,N_1250,N_974);
and U5048 (N_5048,N_1125,N_3944);
and U5049 (N_5049,N_4066,N_2715);
or U5050 (N_5050,N_4778,N_1949);
or U5051 (N_5051,N_1923,N_3118);
or U5052 (N_5052,N_4411,N_2953);
and U5053 (N_5053,N_708,N_1606);
and U5054 (N_5054,N_3733,N_2887);
or U5055 (N_5055,N_4875,N_2395);
and U5056 (N_5056,N_2261,N_3352);
and U5057 (N_5057,N_4783,N_3356);
or U5058 (N_5058,N_3102,N_3481);
or U5059 (N_5059,N_2375,N_652);
or U5060 (N_5060,N_4312,N_4508);
nand U5061 (N_5061,N_1393,N_710);
xor U5062 (N_5062,N_4557,N_4539);
nor U5063 (N_5063,N_1461,N_2783);
and U5064 (N_5064,N_2538,N_3124);
nand U5065 (N_5065,N_4042,N_4428);
nand U5066 (N_5066,N_3683,N_3346);
and U5067 (N_5067,N_1753,N_529);
nor U5068 (N_5068,N_544,N_929);
and U5069 (N_5069,N_1392,N_3204);
and U5070 (N_5070,N_3223,N_2381);
and U5071 (N_5071,N_1568,N_3446);
nor U5072 (N_5072,N_4372,N_2463);
nor U5073 (N_5073,N_2271,N_3402);
nor U5074 (N_5074,N_4479,N_1871);
and U5075 (N_5075,N_4785,N_4268);
nand U5076 (N_5076,N_2960,N_4888);
xnor U5077 (N_5077,N_2111,N_1459);
nand U5078 (N_5078,N_3913,N_4914);
nand U5079 (N_5079,N_2927,N_3533);
and U5080 (N_5080,N_365,N_1876);
or U5081 (N_5081,N_3770,N_1657);
nand U5082 (N_5082,N_3478,N_4473);
or U5083 (N_5083,N_1413,N_2459);
nor U5084 (N_5084,N_2990,N_1724);
nor U5085 (N_5085,N_1601,N_4697);
and U5086 (N_5086,N_2037,N_4512);
and U5087 (N_5087,N_4300,N_72);
or U5088 (N_5088,N_3235,N_2382);
and U5089 (N_5089,N_2033,N_3562);
and U5090 (N_5090,N_4103,N_3985);
nand U5091 (N_5091,N_2251,N_4366);
and U5092 (N_5092,N_1207,N_4152);
nor U5093 (N_5093,N_1690,N_2041);
nor U5094 (N_5094,N_2687,N_470);
nand U5095 (N_5095,N_2473,N_4409);
or U5096 (N_5096,N_198,N_2460);
nand U5097 (N_5097,N_3295,N_508);
or U5098 (N_5098,N_4381,N_1932);
nor U5099 (N_5099,N_3852,N_2408);
nand U5100 (N_5100,N_538,N_826);
or U5101 (N_5101,N_4279,N_3858);
nand U5102 (N_5102,N_2167,N_3826);
nor U5103 (N_5103,N_3109,N_1056);
nand U5104 (N_5104,N_1277,N_1020);
or U5105 (N_5105,N_2400,N_4593);
nand U5106 (N_5106,N_2920,N_54);
or U5107 (N_5107,N_4863,N_4905);
and U5108 (N_5108,N_1443,N_3008);
nand U5109 (N_5109,N_723,N_1643);
or U5110 (N_5110,N_3623,N_788);
and U5111 (N_5111,N_278,N_918);
and U5112 (N_5112,N_2841,N_903);
nand U5113 (N_5113,N_1473,N_711);
or U5114 (N_5114,N_410,N_2055);
nor U5115 (N_5115,N_34,N_1880);
or U5116 (N_5116,N_284,N_3798);
and U5117 (N_5117,N_855,N_1363);
nor U5118 (N_5118,N_4080,N_4390);
nand U5119 (N_5119,N_900,N_957);
nor U5120 (N_5120,N_404,N_2994);
nor U5121 (N_5121,N_2232,N_4965);
xnor U5122 (N_5122,N_3513,N_2120);
nand U5123 (N_5123,N_1229,N_913);
nor U5124 (N_5124,N_3397,N_4639);
or U5125 (N_5125,N_3382,N_1798);
nand U5126 (N_5126,N_421,N_4681);
or U5127 (N_5127,N_4034,N_4215);
and U5128 (N_5128,N_3987,N_2038);
or U5129 (N_5129,N_2601,N_3656);
or U5130 (N_5130,N_4611,N_4980);
or U5131 (N_5131,N_2652,N_422);
nand U5132 (N_5132,N_3393,N_3471);
or U5133 (N_5133,N_3276,N_4347);
nor U5134 (N_5134,N_1318,N_3037);
nor U5135 (N_5135,N_4736,N_3129);
and U5136 (N_5136,N_2341,N_3467);
or U5137 (N_5137,N_1300,N_1692);
xnor U5138 (N_5138,N_4089,N_3563);
or U5139 (N_5139,N_820,N_3810);
nand U5140 (N_5140,N_4072,N_4961);
nand U5141 (N_5141,N_59,N_2478);
and U5142 (N_5142,N_681,N_1426);
or U5143 (N_5143,N_563,N_3018);
or U5144 (N_5144,N_4928,N_3064);
and U5145 (N_5145,N_1043,N_3054);
nor U5146 (N_5146,N_2329,N_0);
and U5147 (N_5147,N_3297,N_2632);
nand U5148 (N_5148,N_2756,N_4146);
nor U5149 (N_5149,N_2258,N_2540);
nor U5150 (N_5150,N_4203,N_3293);
nand U5151 (N_5151,N_133,N_9);
nor U5152 (N_5152,N_1799,N_3399);
nor U5153 (N_5153,N_4500,N_1626);
and U5154 (N_5154,N_3709,N_35);
nand U5155 (N_5155,N_3141,N_3797);
and U5156 (N_5156,N_156,N_1581);
or U5157 (N_5157,N_3470,N_3166);
nor U5158 (N_5158,N_2061,N_2587);
nand U5159 (N_5159,N_477,N_2048);
or U5160 (N_5160,N_670,N_67);
or U5161 (N_5161,N_1902,N_4504);
or U5162 (N_5162,N_2978,N_2529);
nor U5163 (N_5163,N_3576,N_174);
and U5164 (N_5164,N_675,N_1794);
nor U5165 (N_5165,N_2136,N_4936);
or U5166 (N_5166,N_2688,N_3909);
and U5167 (N_5167,N_2233,N_1711);
xor U5168 (N_5168,N_3714,N_3344);
or U5169 (N_5169,N_245,N_3973);
and U5170 (N_5170,N_4092,N_4290);
or U5171 (N_5171,N_3574,N_3867);
nand U5172 (N_5172,N_1491,N_1398);
and U5173 (N_5173,N_3396,N_986);
nor U5174 (N_5174,N_4664,N_897);
xor U5175 (N_5175,N_2918,N_1573);
nand U5176 (N_5176,N_3773,N_3818);
nor U5177 (N_5177,N_2151,N_2230);
nand U5178 (N_5178,N_2524,N_481);
or U5179 (N_5179,N_3946,N_377);
nor U5180 (N_5180,N_642,N_4569);
nand U5181 (N_5181,N_2647,N_3322);
or U5182 (N_5182,N_2757,N_2397);
nor U5183 (N_5183,N_1041,N_3047);
and U5184 (N_5184,N_1050,N_4741);
nor U5185 (N_5185,N_1620,N_1727);
or U5186 (N_5186,N_2586,N_1676);
nor U5187 (N_5187,N_1265,N_591);
and U5188 (N_5188,N_3260,N_2496);
nor U5189 (N_5189,N_1122,N_4046);
nand U5190 (N_5190,N_1939,N_1731);
nand U5191 (N_5191,N_2740,N_3903);
or U5192 (N_5192,N_4809,N_2822);
or U5193 (N_5193,N_110,N_715);
and U5194 (N_5194,N_3831,N_2682);
or U5195 (N_5195,N_4458,N_4418);
nand U5196 (N_5196,N_205,N_3571);
and U5197 (N_5197,N_2186,N_2217);
or U5198 (N_5198,N_3219,N_3299);
and U5199 (N_5199,N_968,N_2116);
nor U5200 (N_5200,N_696,N_3924);
or U5201 (N_5201,N_976,N_3658);
and U5202 (N_5202,N_4180,N_2380);
nor U5203 (N_5203,N_1844,N_3560);
nand U5204 (N_5204,N_4449,N_1533);
or U5205 (N_5205,N_23,N_4261);
or U5206 (N_5206,N_2807,N_1890);
or U5207 (N_5207,N_3572,N_4813);
and U5208 (N_5208,N_2317,N_4478);
and U5209 (N_5209,N_535,N_2215);
nor U5210 (N_5210,N_3937,N_275);
and U5211 (N_5211,N_1380,N_1675);
nor U5212 (N_5212,N_3310,N_1184);
and U5213 (N_5213,N_1191,N_1947);
or U5214 (N_5214,N_2670,N_4594);
nor U5215 (N_5215,N_348,N_962);
or U5216 (N_5216,N_3547,N_1935);
or U5217 (N_5217,N_2816,N_4963);
and U5218 (N_5218,N_4748,N_465);
or U5219 (N_5219,N_460,N_1320);
and U5220 (N_5220,N_241,N_2651);
nand U5221 (N_5221,N_2805,N_532);
nand U5222 (N_5222,N_2311,N_744);
nand U5223 (N_5223,N_3370,N_4790);
nand U5224 (N_5224,N_1295,N_327);
or U5225 (N_5225,N_4059,N_3596);
or U5226 (N_5226,N_844,N_4618);
and U5227 (N_5227,N_4388,N_2253);
nand U5228 (N_5228,N_1354,N_3390);
nand U5229 (N_5229,N_1789,N_1176);
xor U5230 (N_5230,N_1506,N_679);
nor U5231 (N_5231,N_227,N_2596);
and U5232 (N_5232,N_3379,N_995);
nand U5233 (N_5233,N_1351,N_2158);
nand U5234 (N_5234,N_282,N_1924);
and U5235 (N_5235,N_1544,N_4002);
and U5236 (N_5236,N_1817,N_2210);
nor U5237 (N_5237,N_3080,N_288);
nand U5238 (N_5238,N_2152,N_1014);
and U5239 (N_5239,N_1030,N_4257);
or U5240 (N_5240,N_11,N_46);
and U5241 (N_5241,N_4604,N_1781);
nand U5242 (N_5242,N_2624,N_1463);
and U5243 (N_5243,N_3180,N_3318);
or U5244 (N_5244,N_182,N_2778);
and U5245 (N_5245,N_2083,N_526);
or U5246 (N_5246,N_2906,N_3633);
nor U5247 (N_5247,N_673,N_395);
and U5248 (N_5248,N_4538,N_4891);
nand U5249 (N_5249,N_2803,N_2338);
or U5250 (N_5250,N_2826,N_3104);
nand U5251 (N_5251,N_4139,N_1726);
and U5252 (N_5252,N_2200,N_1499);
nand U5253 (N_5253,N_3215,N_2537);
nor U5254 (N_5254,N_3965,N_3463);
nand U5255 (N_5255,N_4584,N_1057);
and U5256 (N_5256,N_1080,N_2367);
nand U5257 (N_5257,N_611,N_4029);
and U5258 (N_5258,N_2628,N_1460);
and U5259 (N_5259,N_3445,N_1126);
nor U5260 (N_5260,N_4796,N_1655);
nor U5261 (N_5261,N_3271,N_302);
or U5262 (N_5262,N_4601,N_2535);
nand U5263 (N_5263,N_265,N_3169);
and U5264 (N_5264,N_4142,N_1369);
nor U5265 (N_5265,N_3569,N_2159);
or U5266 (N_5266,N_3435,N_4025);
and U5267 (N_5267,N_3545,N_121);
nor U5268 (N_5268,N_2594,N_2570);
nor U5269 (N_5269,N_2323,N_1151);
and U5270 (N_5270,N_129,N_506);
nand U5271 (N_5271,N_2372,N_1964);
xnor U5272 (N_5272,N_2679,N_3464);
and U5273 (N_5273,N_3282,N_2800);
nand U5274 (N_5274,N_1329,N_2267);
and U5275 (N_5275,N_2823,N_3094);
and U5276 (N_5276,N_2842,N_2391);
nand U5277 (N_5277,N_3962,N_707);
nand U5278 (N_5278,N_1303,N_3898);
or U5279 (N_5279,N_651,N_1774);
or U5280 (N_5280,N_3044,N_644);
nand U5281 (N_5281,N_1879,N_1034);
nor U5282 (N_5282,N_1173,N_2925);
nor U5283 (N_5283,N_127,N_3558);
nor U5284 (N_5284,N_3431,N_1747);
and U5285 (N_5285,N_4067,N_4063);
nor U5286 (N_5286,N_91,N_3253);
nand U5287 (N_5287,N_326,N_1023);
and U5288 (N_5288,N_4466,N_1679);
nor U5289 (N_5289,N_3388,N_12);
nand U5290 (N_5290,N_4709,N_4082);
nand U5291 (N_5291,N_2465,N_2820);
nor U5292 (N_5292,N_4942,N_3305);
nor U5293 (N_5293,N_2222,N_7);
and U5294 (N_5294,N_4629,N_3391);
or U5295 (N_5295,N_4459,N_2074);
nand U5296 (N_5296,N_249,N_2436);
nor U5297 (N_5297,N_2172,N_416);
nor U5298 (N_5298,N_3320,N_2684);
and U5299 (N_5299,N_3438,N_1495);
or U5300 (N_5300,N_2458,N_1878);
or U5301 (N_5301,N_3873,N_2533);
nand U5302 (N_5302,N_1217,N_4669);
nor U5303 (N_5303,N_4859,N_1886);
nor U5304 (N_5304,N_3043,N_4583);
or U5305 (N_5305,N_4143,N_3686);
and U5306 (N_5306,N_4858,N_4693);
nand U5307 (N_5307,N_836,N_3784);
nor U5308 (N_5308,N_2451,N_2543);
and U5309 (N_5309,N_1139,N_3025);
nor U5310 (N_5310,N_2057,N_1042);
and U5311 (N_5311,N_4958,N_2471);
or U5312 (N_5312,N_2815,N_2228);
nand U5313 (N_5313,N_1367,N_4114);
nand U5314 (N_5314,N_2640,N_1252);
and U5315 (N_5315,N_1504,N_2623);
nor U5316 (N_5316,N_414,N_2991);
nand U5317 (N_5317,N_2494,N_2646);
or U5318 (N_5318,N_2551,N_586);
or U5319 (N_5319,N_3042,N_276);
nor U5320 (N_5320,N_301,N_297);
nand U5321 (N_5321,N_925,N_2928);
nand U5322 (N_5322,N_3398,N_135);
nand U5323 (N_5323,N_2195,N_4781);
and U5324 (N_5324,N_285,N_3230);
or U5325 (N_5325,N_2699,N_1513);
and U5326 (N_5326,N_1293,N_961);
and U5327 (N_5327,N_4079,N_943);
or U5328 (N_5328,N_77,N_1732);
and U5329 (N_5329,N_2618,N_3177);
nor U5330 (N_5330,N_4433,N_2910);
or U5331 (N_5331,N_1447,N_4084);
or U5332 (N_5332,N_1467,N_4281);
nand U5333 (N_5333,N_768,N_498);
and U5334 (N_5334,N_1400,N_1331);
or U5335 (N_5335,N_4670,N_3959);
nor U5336 (N_5336,N_2087,N_2641);
nor U5337 (N_5337,N_1859,N_1756);
or U5338 (N_5338,N_360,N_1596);
nor U5339 (N_5339,N_257,N_4019);
nor U5340 (N_5340,N_1296,N_4149);
nand U5341 (N_5341,N_2536,N_4646);
nand U5342 (N_5342,N_1966,N_4673);
nand U5343 (N_5343,N_1240,N_2418);
nor U5344 (N_5344,N_4075,N_4386);
or U5345 (N_5345,N_1740,N_175);
nor U5346 (N_5346,N_4043,N_1275);
or U5347 (N_5347,N_3786,N_1739);
and U5348 (N_5348,N_2903,N_543);
nand U5349 (N_5349,N_3030,N_4581);
nor U5350 (N_5350,N_592,N_3990);
nor U5351 (N_5351,N_2742,N_3364);
and U5352 (N_5352,N_4582,N_1607);
or U5353 (N_5353,N_3535,N_4493);
and U5354 (N_5354,N_4022,N_1807);
nand U5355 (N_5355,N_2435,N_1550);
nor U5356 (N_5356,N_3525,N_4295);
nor U5357 (N_5357,N_3688,N_3872);
nand U5358 (N_5358,N_1847,N_274);
or U5359 (N_5359,N_493,N_3474);
nand U5360 (N_5360,N_4689,N_3750);
or U5361 (N_5361,N_3184,N_61);
nor U5362 (N_5362,N_1019,N_2550);
nand U5363 (N_5363,N_3549,N_1471);
and U5364 (N_5364,N_3103,N_277);
nand U5365 (N_5365,N_3775,N_3776);
or U5366 (N_5366,N_3365,N_1306);
and U5367 (N_5367,N_310,N_238);
or U5368 (N_5368,N_1082,N_1999);
and U5369 (N_5369,N_874,N_507);
nor U5370 (N_5370,N_4249,N_3306);
or U5371 (N_5371,N_2930,N_1666);
nand U5372 (N_5372,N_1507,N_4305);
and U5373 (N_5373,N_3880,N_3268);
nand U5374 (N_5374,N_4396,N_4608);
or U5375 (N_5375,N_558,N_2515);
nand U5376 (N_5376,N_4714,N_393);
or U5377 (N_5377,N_1309,N_2293);
or U5378 (N_5378,N_1206,N_1083);
or U5379 (N_5379,N_4941,N_4110);
nor U5380 (N_5380,N_2598,N_3274);
nor U5381 (N_5381,N_371,N_4560);
and U5382 (N_5382,N_298,N_1686);
nor U5383 (N_5383,N_4940,N_3617);
nand U5384 (N_5384,N_3294,N_3774);
and U5385 (N_5385,N_1073,N_1772);
nor U5386 (N_5386,N_1917,N_4763);
nand U5387 (N_5387,N_4461,N_2100);
nor U5388 (N_5388,N_2649,N_668);
and U5389 (N_5389,N_1382,N_1600);
or U5390 (N_5390,N_3512,N_1813);
and U5391 (N_5391,N_290,N_2683);
nand U5392 (N_5392,N_2089,N_596);
nand U5393 (N_5393,N_1728,N_27);
nor U5394 (N_5394,N_4031,N_2104);
or U5395 (N_5395,N_2208,N_4823);
nor U5396 (N_5396,N_239,N_4797);
or U5397 (N_5397,N_1431,N_737);
or U5398 (N_5398,N_3874,N_1375);
and U5399 (N_5399,N_2553,N_3527);
or U5400 (N_5400,N_1040,N_803);
nand U5401 (N_5401,N_3579,N_2310);
or U5402 (N_5402,N_1232,N_2593);
nor U5403 (N_5403,N_1809,N_4827);
nand U5404 (N_5404,N_727,N_4545);
or U5405 (N_5405,N_502,N_2140);
nor U5406 (N_5406,N_3105,N_3748);
nand U5407 (N_5407,N_689,N_998);
nand U5408 (N_5408,N_952,N_2563);
nand U5409 (N_5409,N_4271,N_2838);
nand U5410 (N_5410,N_2702,N_4216);
and U5411 (N_5411,N_1412,N_3259);
nor U5412 (N_5412,N_1362,N_3144);
and U5413 (N_5413,N_147,N_108);
or U5414 (N_5414,N_323,N_4705);
nor U5415 (N_5415,N_3347,N_4527);
nand U5416 (N_5416,N_1142,N_143);
nand U5417 (N_5417,N_1560,N_3367);
nand U5418 (N_5418,N_318,N_4549);
nor U5419 (N_5419,N_427,N_1895);
nor U5420 (N_5420,N_2958,N_990);
nor U5421 (N_5421,N_1365,N_3436);
nand U5422 (N_5422,N_4925,N_3803);
nor U5423 (N_5423,N_1285,N_2668);
or U5424 (N_5424,N_4158,N_2781);
xor U5425 (N_5425,N_4678,N_4169);
and U5426 (N_5426,N_4625,N_4990);
nor U5427 (N_5427,N_2901,N_4463);
and U5428 (N_5428,N_636,N_1960);
xor U5429 (N_5429,N_1314,N_647);
nor U5430 (N_5430,N_3062,N_1830);
nand U5431 (N_5431,N_4306,N_3842);
nand U5432 (N_5432,N_686,N_2739);
nand U5433 (N_5433,N_4,N_1591);
nor U5434 (N_5434,N_2517,N_4050);
nand U5435 (N_5435,N_3082,N_838);
or U5436 (N_5436,N_2813,N_793);
and U5437 (N_5437,N_2491,N_4760);
or U5438 (N_5438,N_4647,N_2933);
and U5439 (N_5439,N_24,N_2448);
and U5440 (N_5440,N_3136,N_4655);
or U5441 (N_5441,N_2401,N_1705);
and U5442 (N_5442,N_4931,N_3785);
or U5443 (N_5443,N_3956,N_705);
nand U5444 (N_5444,N_4932,N_312);
or U5445 (N_5445,N_951,N_3926);
xnor U5446 (N_5446,N_3619,N_1084);
nand U5447 (N_5447,N_3366,N_4016);
and U5448 (N_5448,N_3416,N_2212);
and U5449 (N_5449,N_2327,N_802);
nand U5450 (N_5450,N_3553,N_1103);
nor U5451 (N_5451,N_985,N_3920);
or U5452 (N_5452,N_4897,N_1337);
nor U5453 (N_5453,N_4324,N_1108);
nor U5454 (N_5454,N_317,N_3114);
and U5455 (N_5455,N_444,N_894);
nor U5456 (N_5456,N_1520,N_3466);
and U5457 (N_5457,N_4971,N_937);
and U5458 (N_5458,N_740,N_1166);
nand U5459 (N_5459,N_761,N_627);
and U5460 (N_5460,N_819,N_1963);
nor U5461 (N_5461,N_4124,N_2528);
nand U5462 (N_5462,N_3779,N_2404);
nor U5463 (N_5463,N_1755,N_4145);
nor U5464 (N_5464,N_20,N_633);
or U5465 (N_5465,N_3531,N_3639);
nor U5466 (N_5466,N_1266,N_1067);
and U5467 (N_5467,N_105,N_478);
or U5468 (N_5468,N_3741,N_3964);
nand U5469 (N_5469,N_1282,N_4865);
and U5470 (N_5470,N_4755,N_1332);
nand U5471 (N_5471,N_4294,N_577);
nand U5472 (N_5472,N_2804,N_4830);
nor U5473 (N_5473,N_1647,N_717);
or U5474 (N_5474,N_397,N_2211);
nand U5475 (N_5475,N_4571,N_4472);
and U5476 (N_5476,N_682,N_4615);
nand U5477 (N_5477,N_4652,N_1933);
or U5478 (N_5478,N_3460,N_4534);
nand U5479 (N_5479,N_3529,N_3999);
nand U5480 (N_5480,N_2749,N_2472);
or U5481 (N_5481,N_455,N_2125);
nor U5482 (N_5482,N_2560,N_4619);
or U5483 (N_5483,N_4917,N_3745);
nor U5484 (N_5484,N_839,N_2464);
or U5485 (N_5485,N_1381,N_2452);
and U5486 (N_5486,N_247,N_1819);
nand U5487 (N_5487,N_3743,N_2312);
and U5488 (N_5488,N_2824,N_620);
and U5489 (N_5489,N_2274,N_594);
or U5490 (N_5490,N_1714,N_2706);
nand U5491 (N_5491,N_1328,N_1353);
nor U5492 (N_5492,N_805,N_2081);
nand U5493 (N_5493,N_4754,N_2578);
or U5494 (N_5494,N_2664,N_3736);
or U5495 (N_5495,N_1595,N_3884);
and U5496 (N_5496,N_3634,N_3283);
and U5497 (N_5497,N_429,N_4464);
or U5498 (N_5498,N_1782,N_471);
nor U5499 (N_5499,N_2872,N_1190);
nor U5500 (N_5500,N_415,N_1047);
and U5501 (N_5501,N_2655,N_4501);
or U5502 (N_5502,N_2434,N_83);
or U5503 (N_5503,N_1095,N_2772);
or U5504 (N_5504,N_413,N_462);
or U5505 (N_5505,N_3500,N_1012);
nand U5506 (N_5506,N_2028,N_2738);
and U5507 (N_5507,N_3954,N_3304);
nor U5508 (N_5508,N_2879,N_4984);
or U5509 (N_5509,N_437,N_2429);
nand U5510 (N_5510,N_2874,N_3640);
or U5511 (N_5511,N_4235,N_2997);
or U5512 (N_5512,N_3162,N_2345);
nand U5513 (N_5513,N_1671,N_4273);
nand U5514 (N_5514,N_3725,N_1909);
or U5515 (N_5515,N_2676,N_3765);
nand U5516 (N_5516,N_4543,N_3063);
or U5517 (N_5517,N_4400,N_4240);
nor U5518 (N_5518,N_3655,N_3326);
nor U5519 (N_5519,N_3910,N_3314);
or U5520 (N_5520,N_452,N_1336);
nand U5521 (N_5521,N_1893,N_4982);
or U5522 (N_5522,N_3731,N_4335);
nand U5523 (N_5523,N_858,N_2453);
nand U5524 (N_5524,N_2965,N_1632);
and U5525 (N_5525,N_2082,N_3394);
nor U5526 (N_5526,N_4605,N_1498);
and U5527 (N_5527,N_1765,N_4060);
and U5528 (N_5528,N_3667,N_2753);
or U5529 (N_5529,N_4732,N_2970);
nand U5530 (N_5530,N_3298,N_356);
and U5531 (N_5531,N_3694,N_2294);
nor U5532 (N_5532,N_4374,N_865);
nor U5533 (N_5533,N_2245,N_1575);
nand U5534 (N_5534,N_2180,N_3705);
and U5535 (N_5535,N_3419,N_2270);
and U5536 (N_5536,N_875,N_4480);
or U5537 (N_5537,N_3300,N_496);
or U5538 (N_5538,N_3877,N_4804);
nand U5539 (N_5539,N_1851,N_1927);
and U5540 (N_5540,N_1298,N_1132);
or U5541 (N_5541,N_4743,N_2108);
xor U5542 (N_5542,N_4630,N_1280);
and U5543 (N_5543,N_4272,N_1662);
and U5544 (N_5544,N_492,N_665);
or U5545 (N_5545,N_4731,N_3612);
nand U5546 (N_5546,N_3040,N_2328);
nor U5547 (N_5547,N_841,N_3796);
and U5548 (N_5548,N_3280,N_2192);
and U5549 (N_5549,N_4762,N_2493);
nor U5550 (N_5550,N_1841,N_2669);
nand U5551 (N_5551,N_4270,N_847);
or U5552 (N_5552,N_3830,N_319);
nand U5553 (N_5553,N_2221,N_3893);
nand U5554 (N_5554,N_2387,N_4179);
nand U5555 (N_5555,N_3224,N_263);
and U5556 (N_5556,N_762,N_2846);
nand U5557 (N_5557,N_1484,N_3395);
and U5558 (N_5558,N_2495,N_2727);
nor U5559 (N_5559,N_1355,N_1215);
and U5560 (N_5560,N_619,N_4219);
nand U5561 (N_5561,N_4727,N_4246);
nor U5562 (N_5562,N_1253,N_1610);
or U5563 (N_5563,N_179,N_4443);
nor U5564 (N_5564,N_3723,N_1599);
nor U5565 (N_5565,N_3241,N_3591);
or U5566 (N_5566,N_2248,N_4590);
nor U5567 (N_5567,N_4108,N_3122);
or U5568 (N_5568,N_4892,N_3163);
or U5569 (N_5569,N_1592,N_4384);
or U5570 (N_5570,N_2921,N_3998);
nand U5571 (N_5571,N_1957,N_3887);
nand U5572 (N_5572,N_2356,N_917);
or U5573 (N_5573,N_810,N_3505);
or U5574 (N_5574,N_345,N_4711);
or U5575 (N_5575,N_3252,N_1029);
or U5576 (N_5576,N_2922,N_1107);
xor U5577 (N_5577,N_1797,N_1723);
and U5578 (N_5578,N_3142,N_3707);
nand U5579 (N_5579,N_942,N_41);
nand U5580 (N_5580,N_4712,N_1405);
and U5581 (N_5581,N_438,N_814);
nand U5582 (N_5582,N_154,N_1861);
or U5583 (N_5583,N_823,N_895);
nor U5584 (N_5584,N_4354,N_3096);
nor U5585 (N_5585,N_4364,N_4383);
or U5586 (N_5586,N_4879,N_1360);
nand U5587 (N_5587,N_4038,N_2863);
xnor U5588 (N_5588,N_4779,N_4451);
nand U5589 (N_5589,N_4227,N_273);
or U5590 (N_5590,N_2091,N_4187);
or U5591 (N_5591,N_749,N_916);
nor U5592 (N_5592,N_1980,N_1684);
nor U5593 (N_5593,N_3716,N_1004);
and U5594 (N_5594,N_2394,N_1776);
nand U5595 (N_5595,N_2132,N_4163);
nand U5596 (N_5596,N_1334,N_3468);
or U5597 (N_5597,N_40,N_2056);
or U5598 (N_5598,N_3302,N_1419);
or U5599 (N_5599,N_3482,N_4144);
nand U5600 (N_5600,N_568,N_607);
nor U5601 (N_5601,N_240,N_3088);
nand U5602 (N_5602,N_1652,N_2325);
nand U5603 (N_5603,N_4955,N_385);
nand U5604 (N_5604,N_106,N_617);
nor U5605 (N_5605,N_1673,N_4536);
or U5606 (N_5606,N_2486,N_1865);
and U5607 (N_5607,N_388,N_1477);
nand U5608 (N_5608,N_550,N_1518);
and U5609 (N_5609,N_3698,N_2617);
and U5610 (N_5610,N_3342,N_4636);
and U5611 (N_5611,N_1302,N_2575);
nor U5612 (N_5612,N_1875,N_1625);
nand U5613 (N_5613,N_1704,N_485);
or U5614 (N_5614,N_2516,N_3503);
and U5615 (N_5615,N_4359,N_4017);
nand U5616 (N_5616,N_1887,N_2224);
nand U5617 (N_5617,N_1154,N_4419);
or U5618 (N_5618,N_2142,N_3012);
nor U5619 (N_5619,N_4435,N_849);
nand U5620 (N_5620,N_801,N_2468);
and U5621 (N_5621,N_4173,N_4405);
and U5622 (N_5622,N_3936,N_928);
or U5623 (N_5623,N_3487,N_2888);
nor U5624 (N_5624,N_2996,N_4292);
and U5625 (N_5625,N_2830,N_3941);
or U5626 (N_5626,N_4414,N_3488);
nor U5627 (N_5627,N_1961,N_3751);
and U5628 (N_5628,N_1315,N_562);
nor U5629 (N_5629,N_1045,N_1446);
nand U5630 (N_5630,N_4953,N_3135);
or U5631 (N_5631,N_1356,N_3782);
nand U5632 (N_5632,N_4018,N_799);
and U5633 (N_5633,N_4319,N_181);
and U5634 (N_5634,N_1286,N_2181);
or U5635 (N_5635,N_3894,N_3111);
nor U5636 (N_5636,N_4808,N_1340);
xor U5637 (N_5637,N_3170,N_1445);
nor U5638 (N_5638,N_2145,N_2698);
or U5639 (N_5639,N_2269,N_3629);
nor U5640 (N_5640,N_1574,N_780);
nand U5641 (N_5641,N_3410,N_37);
and U5642 (N_5642,N_653,N_2276);
and U5643 (N_5643,N_3628,N_417);
nor U5644 (N_5644,N_3413,N_975);
nor U5645 (N_5645,N_1542,N_1754);
nand U5646 (N_5646,N_1197,N_4412);
and U5647 (N_5647,N_1186,N_2962);
nand U5648 (N_5648,N_4469,N_835);
and U5649 (N_5649,N_2725,N_4951);
nor U5650 (N_5650,N_1399,N_1906);
nor U5651 (N_5651,N_1667,N_2643);
and U5652 (N_5652,N_3155,N_2712);
nor U5653 (N_5653,N_536,N_2777);
or U5654 (N_5654,N_1646,N_4127);
and U5655 (N_5655,N_4998,N_1245);
and U5656 (N_5656,N_2525,N_1395);
nor U5657 (N_5657,N_3070,N_1811);
and U5658 (N_5658,N_221,N_2036);
nor U5659 (N_5659,N_3159,N_1976);
or U5660 (N_5660,N_1842,N_267);
nor U5661 (N_5661,N_4098,N_3710);
nor U5662 (N_5662,N_4657,N_605);
or U5663 (N_5663,N_3422,N_1200);
and U5664 (N_5664,N_4171,N_4541);
xnor U5665 (N_5665,N_1541,N_1535);
nand U5666 (N_5666,N_4233,N_2883);
xor U5667 (N_5667,N_3506,N_880);
nor U5668 (N_5668,N_4402,N_2557);
and U5669 (N_5669,N_96,N_2257);
nand U5670 (N_5670,N_3644,N_2357);
or U5671 (N_5671,N_2018,N_1670);
nand U5672 (N_5672,N_4170,N_695);
or U5673 (N_5673,N_811,N_3450);
nand U5674 (N_5674,N_2876,N_3205);
nand U5675 (N_5675,N_3516,N_4119);
and U5676 (N_5676,N_1182,N_783);
nand U5677 (N_5677,N_268,N_1039);
nor U5678 (N_5678,N_2148,N_950);
nor U5679 (N_5679,N_403,N_2678);
nor U5680 (N_5680,N_320,N_654);
nand U5681 (N_5681,N_2207,N_3138);
nor U5682 (N_5682,N_1060,N_3663);
or U5683 (N_5683,N_3981,N_3409);
nand U5684 (N_5684,N_2539,N_4908);
or U5685 (N_5685,N_2793,N_2030);
or U5686 (N_5686,N_1508,N_69);
and U5687 (N_5687,N_4323,N_3739);
nor U5688 (N_5688,N_128,N_4413);
nand U5689 (N_5689,N_4814,N_4475);
and U5690 (N_5690,N_4313,N_4429);
nor U5691 (N_5691,N_66,N_1048);
nor U5692 (N_5692,N_1105,N_3957);
nor U5693 (N_5693,N_1391,N_3036);
or U5694 (N_5694,N_3679,N_3006);
nor U5695 (N_5695,N_871,N_2406);
or U5696 (N_5696,N_842,N_3199);
xnor U5697 (N_5697,N_548,N_1984);
or U5698 (N_5698,N_1489,N_3301);
and U5699 (N_5699,N_3179,N_3387);
nand U5700 (N_5700,N_2234,N_1580);
and U5701 (N_5701,N_4438,N_2981);
nand U5702 (N_5702,N_3130,N_4922);
nor U5703 (N_5703,N_4175,N_4289);
or U5704 (N_5704,N_2289,N_4004);
nand U5705 (N_5705,N_1651,N_2069);
nand U5706 (N_5706,N_1198,N_2787);
and U5707 (N_5707,N_3154,N_2754);
and U5708 (N_5708,N_1326,N_4453);
or U5709 (N_5709,N_3443,N_3048);
or U5710 (N_5710,N_2574,N_2878);
and U5711 (N_5711,N_4027,N_2919);
xor U5712 (N_5712,N_1072,N_1517);
and U5713 (N_5713,N_2847,N_1335);
or U5714 (N_5714,N_4104,N_2737);
nand U5715 (N_5715,N_1911,N_3333);
and U5716 (N_5716,N_4439,N_3238);
nor U5717 (N_5717,N_1235,N_691);
or U5718 (N_5718,N_4759,N_1321);
and U5719 (N_5719,N_119,N_4254);
and U5720 (N_5720,N_270,N_4724);
nand U5721 (N_5721,N_3383,N_4902);
or U5722 (N_5722,N_1579,N_1702);
and U5723 (N_5723,N_4764,N_2915);
nand U5724 (N_5724,N_4490,N_1611);
and U5725 (N_5725,N_177,N_2964);
nor U5726 (N_5726,N_731,N_1572);
and U5727 (N_5727,N_3381,N_401);
and U5728 (N_5728,N_2561,N_3835);
or U5729 (N_5729,N_1005,N_645);
or U5730 (N_5730,N_2576,N_4220);
nor U5731 (N_5731,N_833,N_4515);
and U5732 (N_5732,N_4805,N_2833);
and U5733 (N_5733,N_2789,N_4242);
nand U5734 (N_5734,N_4446,N_3996);
nand U5735 (N_5735,N_2032,N_2109);
and U5736 (N_5736,N_2487,N_90);
and U5737 (N_5737,N_1522,N_4924);
or U5738 (N_5738,N_1133,N_898);
nand U5739 (N_5739,N_4873,N_184);
and U5740 (N_5740,N_2771,N_1221);
nor U5741 (N_5741,N_2681,N_4120);
nand U5742 (N_5742,N_3097,N_2791);
or U5743 (N_5743,N_4000,N_2658);
and U5744 (N_5744,N_4130,N_4880);
nand U5745 (N_5745,N_4314,N_1954);
or U5746 (N_5746,N_3757,N_3914);
nor U5747 (N_5747,N_2165,N_4710);
nor U5748 (N_5748,N_1571,N_55);
and U5749 (N_5749,N_2526,N_116);
nand U5750 (N_5750,N_4214,N_4634);
and U5751 (N_5751,N_3859,N_447);
nand U5752 (N_5752,N_2806,N_4696);
nor U5753 (N_5753,N_4342,N_2073);
nand U5754 (N_5754,N_3081,N_4658);
nor U5755 (N_5755,N_2203,N_322);
and U5756 (N_5756,N_1301,N_882);
nor U5757 (N_5757,N_584,N_1339);
nand U5758 (N_5758,N_203,N_2810);
and U5759 (N_5759,N_378,N_4816);
and U5760 (N_5760,N_4668,N_2971);
nor U5761 (N_5761,N_559,N_2389);
and U5762 (N_5762,N_3507,N_2590);
nor U5763 (N_5763,N_3889,N_1833);
nor U5764 (N_5764,N_4026,N_3760);
and U5765 (N_5765,N_4766,N_2047);
nor U5766 (N_5766,N_623,N_2045);
nor U5767 (N_5767,N_2016,N_4430);
nor U5768 (N_5768,N_2541,N_1824);
nor U5769 (N_5769,N_65,N_4699);
or U5770 (N_5770,N_3793,N_4445);
and U5771 (N_5771,N_4415,N_2243);
and U5772 (N_5772,N_2281,N_949);
nand U5773 (N_5773,N_2220,N_666);
nand U5774 (N_5774,N_2610,N_1701);
and U5775 (N_5775,N_2088,N_4252);
nor U5776 (N_5776,N_3581,N_808);
nand U5777 (N_5777,N_183,N_2319);
nand U5778 (N_5778,N_1874,N_753);
or U5779 (N_5779,N_292,N_767);
and U5780 (N_5780,N_13,N_4969);
nand U5781 (N_5781,N_1212,N_53);
or U5782 (N_5782,N_4592,N_1377);
nor U5783 (N_5783,N_2760,N_4794);
nand U5784 (N_5784,N_3107,N_4269);
or U5785 (N_5785,N_165,N_85);
nor U5786 (N_5786,N_4795,N_3110);
and U5787 (N_5787,N_1889,N_1642);
and U5788 (N_5788,N_3992,N_1304);
nand U5789 (N_5789,N_4167,N_3139);
nand U5790 (N_5790,N_4015,N_3039);
nor U5791 (N_5791,N_4265,N_4622);
or U5792 (N_5792,N_2568,N_1470);
and U5793 (N_5793,N_4850,N_4083);
and U5794 (N_5794,N_4994,N_1979);
or U5795 (N_5795,N_3227,N_1862);
nor U5796 (N_5796,N_698,N_1294);
and U5797 (N_5797,N_2107,N_4340);
or U5798 (N_5798,N_2860,N_3925);
and U5799 (N_5799,N_693,N_2349);
nor U5800 (N_5800,N_904,N_722);
and U5801 (N_5801,N_1908,N_1766);
and U5802 (N_5802,N_1974,N_3133);
or U5803 (N_5803,N_4837,N_4728);
and U5804 (N_5804,N_4221,N_2374);
or U5805 (N_5805,N_2343,N_978);
nand U5806 (N_5806,N_2619,N_4944);
nor U5807 (N_5807,N_3087,N_4116);
nand U5808 (N_5808,N_4974,N_883);
nand U5809 (N_5809,N_843,N_1032);
or U5810 (N_5810,N_557,N_4155);
and U5811 (N_5811,N_688,N_1995);
nor U5812 (N_5812,N_2333,N_4424);
nand U5813 (N_5813,N_3544,N_1900);
or U5814 (N_5814,N_3161,N_587);
nand U5815 (N_5815,N_353,N_4822);
nand U5816 (N_5816,N_4024,N_807);
and U5817 (N_5817,N_759,N_3029);
and U5818 (N_5818,N_4899,N_1760);
nand U5819 (N_5819,N_4327,N_4665);
and U5820 (N_5820,N_2912,N_2114);
or U5821 (N_5821,N_1697,N_420);
or U5822 (N_5822,N_1187,N_3789);
and U5823 (N_5823,N_1803,N_4053);
or U5824 (N_5824,N_3868,N_969);
and U5825 (N_5825,N_3790,N_367);
nand U5826 (N_5826,N_3524,N_637);
or U5827 (N_5827,N_1674,N_2266);
and U5828 (N_5828,N_4803,N_3787);
nor U5829 (N_5829,N_1539,N_4245);
or U5830 (N_5830,N_2607,N_433);
nor U5831 (N_5831,N_4920,N_1174);
and U5832 (N_5832,N_3498,N_1468);
nand U5833 (N_5833,N_1269,N_89);
or U5834 (N_5834,N_4420,N_2857);
nor U5835 (N_5835,N_63,N_4185);
and U5836 (N_5836,N_987,N_4126);
nor U5837 (N_5837,N_2348,N_3190);
and U5838 (N_5838,N_2106,N_2161);
and U5839 (N_5839,N_2183,N_4172);
or U5840 (N_5840,N_3430,N_2673);
nand U5841 (N_5841,N_3401,N_3192);
nand U5842 (N_5842,N_3191,N_4460);
or U5843 (N_5843,N_4006,N_2614);
nor U5844 (N_5844,N_4194,N_1515);
and U5845 (N_5845,N_1421,N_3338);
nor U5846 (N_5846,N_3072,N_2851);
nand U5847 (N_5847,N_2784,N_1147);
or U5848 (N_5848,N_2392,N_718);
or U5849 (N_5849,N_4062,N_2701);
and U5850 (N_5850,N_2966,N_1525);
and U5851 (N_5851,N_1534,N_1482);
and U5852 (N_5852,N_4744,N_4909);
nand U5853 (N_5853,N_4224,N_1031);
nor U5854 (N_5854,N_463,N_2924);
nor U5855 (N_5855,N_4286,N_4777);
nand U5856 (N_5856,N_2377,N_222);
or U5857 (N_5857,N_4317,N_3670);
nand U5858 (N_5858,N_948,N_3677);
nor U5859 (N_5859,N_1942,N_2667);
or U5860 (N_5860,N_1761,N_1457);
or U5861 (N_5861,N_2945,N_2884);
nand U5862 (N_5862,N_1305,N_3620);
nand U5863 (N_5863,N_3479,N_4131);
nand U5864 (N_5864,N_3207,N_720);
and U5865 (N_5865,N_892,N_4357);
nand U5866 (N_5866,N_1183,N_1837);
nand U5867 (N_5867,N_3551,N_2746);
and U5868 (N_5868,N_683,N_2239);
nand U5869 (N_5869,N_1532,N_3519);
nor U5870 (N_5870,N_2340,N_2513);
nand U5871 (N_5871,N_1623,N_3989);
nand U5872 (N_5872,N_1053,N_391);
nor U5873 (N_5873,N_1219,N_3489);
or U5874 (N_5874,N_3439,N_4486);
nor U5875 (N_5875,N_4526,N_3024);
nand U5876 (N_5876,N_1648,N_1868);
and U5877 (N_5877,N_4703,N_2146);
nor U5878 (N_5878,N_3475,N_1836);
nor U5879 (N_5879,N_374,N_1021);
nand U5880 (N_5880,N_1649,N_4883);
and U5881 (N_5881,N_2144,N_520);
nand U5882 (N_5882,N_2811,N_781);
nor U5883 (N_5883,N_207,N_2332);
nand U5884 (N_5884,N_4112,N_4421);
and U5885 (N_5885,N_1637,N_2322);
nand U5886 (N_5886,N_3019,N_2062);
or U5887 (N_5887,N_1741,N_4524);
or U5888 (N_5888,N_2839,N_583);
nor U5889 (N_5889,N_1453,N_2989);
and U5890 (N_5890,N_2384,N_381);
and U5891 (N_5891,N_1617,N_2728);
nand U5892 (N_5892,N_4135,N_3611);
and U5893 (N_5893,N_4566,N_3239);
nand U5894 (N_5894,N_955,N_3350);
nand U5895 (N_5895,N_3486,N_3501);
nor U5896 (N_5896,N_1993,N_195);
nor U5897 (N_5897,N_1846,N_4923);
nor U5898 (N_5898,N_2873,N_2029);
or U5899 (N_5899,N_1903,N_1587);
nor U5900 (N_5900,N_4895,N_2713);
nand U5901 (N_5901,N_4841,N_1009);
or U5902 (N_5902,N_589,N_4903);
nand U5903 (N_5903,N_1160,N_2581);
or U5904 (N_5904,N_4761,N_531);
nor U5905 (N_5905,N_2985,N_4498);
and U5906 (N_5906,N_2121,N_2065);
or U5907 (N_5907,N_2219,N_3552);
nand U5908 (N_5908,N_1130,N_482);
and U5909 (N_5909,N_4603,N_2431);
nand U5910 (N_5910,N_4885,N_2808);
nor U5911 (N_5911,N_1124,N_3032);
nor U5912 (N_5912,N_1098,N_2365);
nor U5913 (N_5913,N_187,N_3213);
and U5914 (N_5914,N_1458,N_4918);
nand U5915 (N_5915,N_851,N_1715);
nor U5916 (N_5916,N_4248,N_4013);
or U5917 (N_5917,N_1475,N_4447);
or U5918 (N_5918,N_4045,N_3820);
and U5919 (N_5919,N_3938,N_49);
or U5920 (N_5920,N_2755,N_1348);
or U5921 (N_5921,N_979,N_3613);
nor U5922 (N_5922,N_2254,N_4353);
nor U5923 (N_5923,N_384,N_4656);
nor U5924 (N_5924,N_1563,N_3806);
nand U5925 (N_5925,N_2794,N_1823);
nor U5926 (N_5926,N_231,N_2714);
nor U5927 (N_5927,N_1584,N_2287);
and U5928 (N_5928,N_3511,N_4195);
nor U5929 (N_5929,N_3188,N_3022);
nand U5930 (N_5930,N_684,N_4481);
nor U5931 (N_5931,N_4970,N_4857);
and U5932 (N_5932,N_4437,N_2198);
or U5933 (N_5933,N_180,N_1680);
nand U5934 (N_5934,N_3137,N_1260);
nor U5935 (N_5935,N_3055,N_2440);
nor U5936 (N_5936,N_1929,N_3504);
and U5937 (N_5937,N_4842,N_3747);
nand U5938 (N_5938,N_1892,N_2764);
and U5939 (N_5939,N_631,N_2015);
nor U5940 (N_5940,N_3079,N_1156);
nand U5941 (N_5941,N_2986,N_3727);
nand U5942 (N_5942,N_3934,N_436);
nand U5943 (N_5943,N_2042,N_3151);
or U5944 (N_5944,N_1244,N_2954);
nand U5945 (N_5945,N_379,N_1218);
or U5946 (N_5946,N_3945,N_4768);
or U5947 (N_5947,N_4196,N_2892);
or U5948 (N_5948,N_2415,N_2307);
and U5949 (N_5949,N_225,N_702);
nand U5950 (N_5950,N_4090,N_158);
or U5951 (N_5951,N_3495,N_260);
and U5952 (N_5952,N_2748,N_213);
and U5953 (N_5953,N_3871,N_488);
or U5954 (N_5954,N_2184,N_1722);
and U5955 (N_5955,N_3448,N_1914);
or U5956 (N_5956,N_3000,N_4208);
and U5957 (N_5957,N_4349,N_2174);
nor U5958 (N_5958,N_1243,N_2188);
nand U5959 (N_5959,N_1002,N_4362);
or U5960 (N_5960,N_996,N_2170);
nor U5961 (N_5961,N_2900,N_4091);
or U5962 (N_5962,N_1414,N_909);
and U5963 (N_5963,N_2941,N_940);
or U5964 (N_5964,N_1719,N_782);
nand U5965 (N_5965,N_3026,N_1236);
nand U5966 (N_5966,N_2209,N_1969);
or U5967 (N_5967,N_4117,N_3583);
nand U5968 (N_5968,N_1858,N_934);
nand U5969 (N_5969,N_1237,N_609);
nand U5970 (N_5970,N_86,N_4977);
nand U5971 (N_5971,N_1808,N_2359);
and U5972 (N_5972,N_2731,N_2636);
and U5973 (N_5973,N_101,N_1444);
nand U5974 (N_5974,N_3876,N_99);
nor U5975 (N_5975,N_4151,N_4621);
nor U5976 (N_5976,N_1919,N_3257);
nand U5977 (N_5977,N_4189,N_4561);
nand U5978 (N_5978,N_1058,N_2868);
and U5979 (N_5979,N_3328,N_1588);
nor U5980 (N_5980,N_4852,N_4910);
and U5981 (N_5981,N_264,N_4577);
nor U5982 (N_5982,N_4654,N_4713);
or U5983 (N_5983,N_512,N_1028);
nor U5984 (N_5984,N_1069,N_1910);
or U5985 (N_5985,N_2388,N_1668);
and U5986 (N_5986,N_95,N_4236);
or U5987 (N_5987,N_4692,N_3007);
and U5988 (N_5988,N_2864,N_1555);
and U5989 (N_5989,N_1230,N_3377);
nor U5990 (N_5990,N_4301,N_3963);
nor U5991 (N_5991,N_4348,N_2767);
xor U5992 (N_5992,N_3057,N_1519);
nor U5993 (N_5993,N_139,N_4878);
and U5994 (N_5994,N_4884,N_476);
nand U5995 (N_5995,N_1901,N_2476);
nor U5996 (N_5996,N_1055,N_2829);
or U5997 (N_5997,N_1462,N_1251);
and U5998 (N_5998,N_3254,N_580);
nand U5999 (N_5999,N_504,N_3860);
and U6000 (N_6000,N_4514,N_2609);
or U6001 (N_6001,N_1157,N_3657);
and U6002 (N_6002,N_2818,N_1543);
nand U6003 (N_6003,N_2393,N_329);
and U6004 (N_6004,N_4860,N_4981);
or U6005 (N_6005,N_1619,N_3746);
and U6006 (N_6006,N_1877,N_864);
nor U6007 (N_6007,N_2155,N_4685);
and U6008 (N_6008,N_1324,N_3113);
nand U6009 (N_6009,N_770,N_4280);
nor U6010 (N_6010,N_1239,N_1989);
nand U6011 (N_6011,N_1113,N_4416);
or U6012 (N_6012,N_2013,N_2890);
and U6013 (N_6013,N_2225,N_3546);
nor U6014 (N_6014,N_411,N_4361);
nand U6015 (N_6015,N_1109,N_1330);
nor U6016 (N_6016,N_3908,N_3834);
nand U6017 (N_6017,N_1757,N_2943);
or U6018 (N_6018,N_3578,N_4820);
or U6019 (N_6019,N_1793,N_3149);
and U6020 (N_6020,N_3832,N_1283);
nor U6021 (N_6021,N_3324,N_3323);
nor U6022 (N_6022,N_4929,N_3210);
and U6023 (N_6023,N_4192,N_2371);
xnor U6024 (N_6024,N_1227,N_2376);
nand U6025 (N_6025,N_2573,N_1435);
nor U6026 (N_6026,N_3247,N_4202);
or U6027 (N_6027,N_2169,N_1992);
nor U6028 (N_6028,N_522,N_430);
and U6029 (N_6029,N_51,N_4427);
nand U6030 (N_6030,N_424,N_4989);
nand U6031 (N_6031,N_3816,N_3691);
nand U6032 (N_6032,N_2638,N_4377);
and U6033 (N_6033,N_3212,N_1299);
or U6034 (N_6034,N_1636,N_501);
or U6035 (N_6035,N_4876,N_618);
nor U6036 (N_6036,N_2862,N_2011);
nor U6037 (N_6037,N_1614,N_2792);
and U6038 (N_6038,N_2769,N_3521);
and U6039 (N_6039,N_382,N_3955);
and U6040 (N_6040,N_4262,N_661);
nand U6041 (N_6041,N_3002,N_2127);
and U6042 (N_6042,N_1297,N_1135);
nand U6043 (N_6043,N_3472,N_336);
or U6044 (N_6044,N_4575,N_445);
and U6045 (N_6045,N_2692,N_4510);
nor U6046 (N_6046,N_1943,N_999);
or U6047 (N_6047,N_4182,N_3695);
nand U6048 (N_6048,N_60,N_2331);
nor U6049 (N_6049,N_2799,N_4506);
nand U6050 (N_6050,N_373,N_4422);
or U6051 (N_6051,N_4398,N_1106);
nor U6052 (N_6052,N_189,N_4496);
and U6053 (N_6053,N_2410,N_1863);
nor U6054 (N_6054,N_4529,N_2475);
or U6055 (N_6055,N_314,N_4540);
nand U6056 (N_6056,N_725,N_3221);
and U6057 (N_6057,N_2414,N_2277);
and U6058 (N_6058,N_1268,N_972);
nand U6059 (N_6059,N_2660,N_2370);
nand U6060 (N_6060,N_3185,N_357);
or U6061 (N_6061,N_578,N_625);
nand U6062 (N_6062,N_2730,N_4455);
or U6063 (N_6063,N_3158,N_2084);
or U6064 (N_6064,N_2665,N_303);
xor U6065 (N_6065,N_1566,N_585);
or U6066 (N_6066,N_4553,N_4602);
and U6067 (N_6067,N_2732,N_509);
or U6068 (N_6068,N_4159,N_79);
nor U6069 (N_6069,N_1111,N_2765);
or U6070 (N_6070,N_1247,N_3631);
and U6071 (N_6071,N_4343,N_1792);
or U6072 (N_6072,N_1449,N_261);
and U6073 (N_6073,N_846,N_4877);
or U6074 (N_6074,N_853,N_4845);
nand U6075 (N_6075,N_443,N_1423);
nand U6076 (N_6076,N_1991,N_2238);
nor U6077 (N_6077,N_1422,N_2296);
nor U6078 (N_6078,N_97,N_1930);
and U6079 (N_6079,N_848,N_4776);
and U6080 (N_6080,N_3808,N_3075);
xnor U6081 (N_6081,N_2700,N_3194);
or U6082 (N_6082,N_510,N_2115);
xnor U6083 (N_6083,N_1713,N_3229);
nor U6084 (N_6084,N_2190,N_4483);
and U6085 (N_6085,N_287,N_1849);
or U6086 (N_6086,N_3510,N_3942);
nor U6087 (N_6087,N_2983,N_3892);
nor U6088 (N_6088,N_1729,N_3664);
nand U6089 (N_6089,N_1523,N_2785);
and U6090 (N_6090,N_2674,N_4992);
and U6091 (N_6091,N_3120,N_1850);
or U6092 (N_6092,N_2511,N_3802);
or U6093 (N_6093,N_4912,N_2993);
nand U6094 (N_6094,N_4106,N_2123);
nand U6095 (N_6095,N_383,N_3827);
nor U6096 (N_6096,N_2729,N_4952);
nor U6097 (N_6097,N_988,N_1089);
or U6098 (N_6098,N_4229,N_2802);
or U6099 (N_6099,N_4141,N_3250);
nand U6100 (N_6100,N_4828,N_2518);
or U6101 (N_6101,N_1681,N_1529);
and U6102 (N_6102,N_902,N_1784);
or U6103 (N_6103,N_73,N_4640);
or U6104 (N_6104,N_758,N_1261);
nand U6105 (N_6105,N_3334,N_2236);
and U6106 (N_6106,N_4288,N_3735);
and U6107 (N_6107,N_745,N_2763);
nor U6108 (N_6108,N_201,N_22);
or U6109 (N_6109,N_1650,N_1442);
nor U6110 (N_6110,N_3766,N_3588);
nor U6111 (N_6111,N_4468,N_1433);
nand U6112 (N_6112,N_1178,N_712);
or U6113 (N_6113,N_3804,N_368);
nand U6114 (N_6114,N_889,N_714);
nor U6115 (N_6115,N_3841,N_1209);
and U6116 (N_6116,N_3939,N_4638);
nor U6117 (N_6117,N_3555,N_1167);
and U6118 (N_6118,N_1469,N_74);
nand U6119 (N_6119,N_2014,N_2631);
nor U6120 (N_6120,N_3348,N_3345);
nor U6121 (N_6121,N_4166,N_2179);
or U6122 (N_6122,N_4789,N_1152);
nand U6123 (N_6123,N_763,N_1603);
and U6124 (N_6124,N_824,N_2242);
nand U6125 (N_6125,N_1389,N_4078);
nor U6126 (N_6126,N_3844,N_676);
nor U6127 (N_6127,N_3598,N_4087);
or U6128 (N_6128,N_2474,N_852);
nor U6129 (N_6129,N_4502,N_380);
or U6130 (N_6130,N_2898,N_3799);
nor U6131 (N_6131,N_3917,N_332);
nor U6132 (N_6132,N_4769,N_2446);
and U6133 (N_6133,N_3684,N_2361);
or U6134 (N_6134,N_1778,N_2321);
and U6135 (N_6135,N_4544,N_554);
and U6136 (N_6136,N_2137,N_3233);
nand U6137 (N_6137,N_490,N_3532);
nor U6138 (N_6138,N_872,N_4617);
or U6139 (N_6139,N_571,N_4825);
nand U6140 (N_6140,N_1170,N_1748);
nor U6141 (N_6141,N_2193,N_338);
nand U6142 (N_6142,N_3618,N_3819);
or U6143 (N_6143,N_4906,N_3469);
nor U6144 (N_6144,N_21,N_3195);
or U6145 (N_6145,N_146,N_3378);
and U6146 (N_6146,N_4274,N_3726);
nor U6147 (N_6147,N_2044,N_2812);
or U6148 (N_6148,N_2059,N_4454);
and U6149 (N_6149,N_3100,N_3586);
or U6150 (N_6150,N_2616,N_795);
and U6151 (N_6151,N_4210,N_1627);
nor U6152 (N_6152,N_448,N_235);
and U6153 (N_6153,N_4315,N_4730);
or U6154 (N_6154,N_2096,N_4391);
nor U6155 (N_6155,N_2716,N_3123);
nand U6156 (N_6156,N_4485,N_4734);
or U6157 (N_6157,N_2035,N_3567);
nor U6158 (N_6158,N_405,N_796);
nand U6159 (N_6159,N_4868,N_1148);
and U6160 (N_6160,N_1361,N_18);
and U6161 (N_6161,N_3718,N_2334);
nor U6162 (N_6162,N_980,N_3630);
nor U6163 (N_6163,N_612,N_608);
nor U6164 (N_6164,N_4183,N_4168);
or U6165 (N_6165,N_1127,N_2138);
and U6166 (N_6166,N_1492,N_4378);
or U6167 (N_6167,N_2354,N_1669);
nor U6168 (N_6168,N_1410,N_330);
nor U6169 (N_6169,N_2724,N_4788);
nor U6170 (N_6170,N_347,N_4350);
nor U6171 (N_6171,N_2130,N_4408);
or U6172 (N_6172,N_604,N_1070);
nand U6173 (N_6173,N_1466,N_4266);
nor U6174 (N_6174,N_2430,N_2008);
nor U6175 (N_6175,N_2718,N_1869);
nand U6176 (N_6176,N_2743,N_3662);
nand U6177 (N_6177,N_2711,N_1791);
or U6178 (N_6178,N_140,N_1561);
or U6179 (N_6179,N_4069,N_2426);
nor U6180 (N_6180,N_2103,N_4122);
or U6181 (N_6181,N_30,N_1385);
or U6182 (N_6182,N_4579,N_3256);
or U6183 (N_6183,N_2095,N_4847);
nor U6184 (N_6184,N_2399,N_4470);
nand U6185 (N_6185,N_1749,N_2523);
nand U6186 (N_6186,N_2292,N_4684);
nor U6187 (N_6187,N_64,N_2454);
nor U6188 (N_6188,N_3284,N_4954);
nor U6189 (N_6189,N_4174,N_3997);
or U6190 (N_6190,N_3312,N_2129);
nor U6191 (N_6191,N_3557,N_2500);
and U6192 (N_6192,N_2175,N_1501);
nand U6193 (N_6193,N_3815,N_920);
or U6194 (N_6194,N_487,N_3290);
and U6195 (N_6195,N_4733,N_2490);
nor U6196 (N_6196,N_3485,N_2423);
and U6197 (N_6197,N_1289,N_1978);
and U6198 (N_6198,N_466,N_104);
nor U6199 (N_6199,N_1956,N_4871);
or U6200 (N_6200,N_590,N_2218);
or U6201 (N_6201,N_4751,N_1856);
and U6202 (N_6202,N_1786,N_3752);
or U6203 (N_6203,N_3690,N_2735);
nor U6204 (N_6204,N_2202,N_1102);
and U6205 (N_6205,N_3437,N_102);
nor U6206 (N_6206,N_1845,N_528);
nand U6207 (N_6207,N_4576,N_1853);
nor U6208 (N_6208,N_3311,N_4831);
nor U6209 (N_6209,N_3682,N_912);
and U6210 (N_6210,N_166,N_2902);
nand U6211 (N_6211,N_3780,N_2832);
and U6212 (N_6212,N_3896,N_4904);
or U6213 (N_6213,N_283,N_1589);
nand U6214 (N_6214,N_964,N_4118);
nor U6215 (N_6215,N_4259,N_4663);
nor U6216 (N_6216,N_4471,N_224);
and U6217 (N_6217,N_1428,N_4973);
nand U6218 (N_6218,N_3308,N_3121);
nand U6219 (N_6219,N_78,N_4644);
and U6220 (N_6220,N_2480,N_1046);
nor U6221 (N_6221,N_394,N_2201);
nand U6222 (N_6222,N_742,N_254);
nand U6223 (N_6223,N_130,N_4365);
or U6224 (N_6224,N_2853,N_4368);
or U6225 (N_6225,N_2588,N_3897);
nand U6226 (N_6226,N_1530,N_2639);
and U6227 (N_6227,N_3053,N_830);
or U6228 (N_6228,N_1396,N_648);
and U6229 (N_6229,N_334,N_2836);
and U6230 (N_6230,N_3706,N_3108);
nand U6231 (N_6231,N_2955,N_4991);
nand U6232 (N_6232,N_3119,N_475);
and U6233 (N_6233,N_1621,N_4094);
or U6234 (N_6234,N_2135,N_878);
or U6235 (N_6235,N_2591,N_1531);
or U6236 (N_6236,N_1119,N_3483);
nand U6237 (N_6237,N_4371,N_4519);
and U6238 (N_6238,N_2762,N_2131);
nor U6239 (N_6239,N_4616,N_4334);
nor U6240 (N_6240,N_1383,N_4005);
or U6241 (N_6241,N_1371,N_2606);
and U6242 (N_6242,N_337,N_941);
xor U6243 (N_6243,N_4567,N_511);
xnor U6244 (N_6244,N_4753,N_1717);
or U6245 (N_6245,N_199,N_1292);
and U6246 (N_6246,N_3604,N_3839);
nor U6247 (N_6247,N_428,N_1511);
or U6248 (N_6248,N_1898,N_3953);
nor U6249 (N_6249,N_4745,N_3590);
and U6250 (N_6250,N_3454,N_480);
and U6251 (N_6251,N_2385,N_4102);
and U6252 (N_6252,N_4870,N_2522);
or U6253 (N_6253,N_114,N_3979);
or U6254 (N_6254,N_4578,N_4107);
and U6255 (N_6255,N_4599,N_36);
nor U6256 (N_6256,N_1472,N_406);
xnor U6257 (N_6257,N_1884,N_4887);
nand U6258 (N_6258,N_1913,N_1323);
and U6259 (N_6259,N_831,N_2024);
nand U6260 (N_6260,N_111,N_1832);
nor U6261 (N_6261,N_1730,N_441);
and U6262 (N_6262,N_3704,N_743);
nand U6263 (N_6263,N_2510,N_1264);
and U6264 (N_6264,N_1796,N_3369);
or U6265 (N_6265,N_3279,N_1931);
nand U6266 (N_6266,N_1145,N_1915);
or U6267 (N_6267,N_2076,N_2704);
and U6268 (N_6268,N_3708,N_1624);
and U6269 (N_6269,N_4721,N_656);
nor U6270 (N_6270,N_1079,N_3967);
xor U6271 (N_6271,N_176,N_2880);
nor U6272 (N_6272,N_1718,N_2886);
nor U6273 (N_6273,N_115,N_3361);
and U6274 (N_6274,N_419,N_4113);
nor U6275 (N_6275,N_2944,N_214);
nor U6276 (N_6276,N_3988,N_4134);
or U6277 (N_6277,N_4784,N_1883);
and U6278 (N_6278,N_3508,N_3637);
or U6279 (N_6279,N_3829,N_3661);
or U6280 (N_6280,N_863,N_4251);
and U6281 (N_6281,N_3407,N_2889);
or U6282 (N_6282,N_4133,N_4283);
nor U6283 (N_6283,N_4966,N_2934);
nand U6284 (N_6284,N_4311,N_983);
or U6285 (N_6285,N_2545,N_1695);
and U6286 (N_6286,N_3228,N_1866);
nor U6287 (N_6287,N_4856,N_1465);
or U6288 (N_6288,N_3160,N_3033);
or U6289 (N_6289,N_3115,N_4806);
and U6290 (N_6290,N_4255,N_3768);
and U6291 (N_6291,N_4874,N_4488);
and U6292 (N_6292,N_1359,N_893);
nor U6293 (N_6293,N_4030,N_3477);
nand U6294 (N_6294,N_457,N_185);
nand U6295 (N_6295,N_1770,N_3993);
nand U6296 (N_6296,N_3315,N_1270);
nor U6297 (N_6297,N_3556,N_2569);
nand U6298 (N_6298,N_792,N_14);
and U6299 (N_6299,N_1262,N_1093);
and U6300 (N_6300,N_4959,N_152);
nor U6301 (N_6301,N_1738,N_1242);
nand U6302 (N_6302,N_2946,N_4740);
nand U6303 (N_6303,N_4154,N_4756);
or U6304 (N_6304,N_534,N_3791);
and U6305 (N_6305,N_4358,N_3335);
xnor U6306 (N_6306,N_3972,N_3589);
and U6307 (N_6307,N_1168,N_3854);
and U6308 (N_6308,N_2324,N_1564);
nand U6309 (N_6309,N_4200,N_1703);
nor U6310 (N_6310,N_1276,N_4369);
nor U6311 (N_6311,N_4835,N_3078);
nor U6312 (N_6312,N_2882,N_638);
nor U6313 (N_6313,N_2433,N_2940);
nand U6314 (N_6314,N_3949,N_2871);
nand U6315 (N_6315,N_324,N_4564);
nand U6316 (N_6316,N_1759,N_4125);
nor U6317 (N_6317,N_1455,N_1509);
or U6318 (N_6318,N_2850,N_1608);
xnor U6319 (N_6319,N_2690,N_3209);
or U6320 (N_6320,N_4780,N_355);
nor U6321 (N_6321,N_271,N_2558);
or U6322 (N_6322,N_15,N_2259);
nand U6323 (N_6323,N_3017,N_3881);
and U6324 (N_6324,N_4285,N_1559);
or U6325 (N_6325,N_3888,N_887);
or U6326 (N_6326,N_4425,N_4105);
or U6327 (N_6327,N_1970,N_2633);
nor U6328 (N_6328,N_4052,N_2726);
or U6329 (N_6329,N_3603,N_3172);
and U6330 (N_6330,N_4967,N_4565);
and U6331 (N_6331,N_752,N_570);
nor U6332 (N_6332,N_4309,N_1241);
or U6333 (N_6333,N_614,N_1024);
and U6334 (N_6334,N_671,N_869);
and U6335 (N_6335,N_32,N_1100);
and U6336 (N_6336,N_1254,N_821);
nor U6337 (N_6337,N_2968,N_773);
nand U6338 (N_6338,N_2666,N_2917);
and U6339 (N_6339,N_3313,N_1612);
nor U6340 (N_6340,N_1417,N_560);
and U6341 (N_6341,N_3737,N_4898);
nor U6342 (N_6342,N_746,N_3245);
nand U6343 (N_6343,N_1386,N_2022);
nand U6344 (N_6344,N_3277,N_2780);
and U6345 (N_6345,N_1117,N_2814);
and U6346 (N_6346,N_812,N_1424);
nand U6347 (N_6347,N_2546,N_151);
or U6348 (N_6348,N_3781,N_1333);
and U6349 (N_6349,N_1758,N_87);
nor U6350 (N_6350,N_1752,N_876);
and U6351 (N_6351,N_3052,N_3292);
nand U6352 (N_6352,N_3355,N_2295);
or U6353 (N_6353,N_2622,N_2600);
nor U6354 (N_6354,N_923,N_2744);
or U6355 (N_6355,N_3051,N_4345);
or U6356 (N_6356,N_2654,N_2026);
or U6357 (N_6357,N_2508,N_237);
and U6358 (N_6358,N_2425,N_50);
nand U6359 (N_6359,N_4886,N_1656);
nor U6360 (N_6360,N_1767,N_2066);
or U6361 (N_6361,N_1211,N_3794);
and U6362 (N_6362,N_1578,N_1456);
and U6363 (N_6363,N_1694,N_1736);
nor U6364 (N_6364,N_3570,N_4793);
nor U6365 (N_6365,N_1815,N_3231);
and U6366 (N_6366,N_2300,N_667);
and U6367 (N_6367,N_1615,N_4786);
nand U6368 (N_6368,N_236,N_1408);
nor U6369 (N_6369,N_4945,N_1101);
nand U6370 (N_6370,N_4975,N_2947);
nand U6371 (N_6371,N_4296,N_3198);
or U6372 (N_6372,N_573,N_3693);
and U6373 (N_6373,N_2980,N_3189);
nor U6374 (N_6374,N_2316,N_2907);
and U6375 (N_6375,N_1407,N_4950);
and U6376 (N_6376,N_760,N_1272);
nand U6377 (N_6377,N_574,N_3461);
nand U6378 (N_6378,N_26,N_3838);
nor U6379 (N_6379,N_4694,N_3561);
nor U6380 (N_6380,N_1720,N_1420);
xor U6381 (N_6381,N_118,N_3289);
nand U6382 (N_6382,N_1146,N_4838);
nand U6383 (N_6383,N_4260,N_519);
and U6384 (N_6384,N_1775,N_306);
or U6385 (N_6385,N_3966,N_3597);
nand U6386 (N_6386,N_1548,N_4792);
nor U6387 (N_6387,N_4287,N_1313);
nor U6388 (N_6388,N_2534,N_3173);
nor U6389 (N_6389,N_4735,N_1274);
nor U6390 (N_6390,N_1051,N_840);
nand U6391 (N_6391,N_4212,N_2204);
and U6392 (N_6392,N_1881,N_1136);
nor U6393 (N_6393,N_3046,N_2484);
nand U6394 (N_6394,N_1941,N_3425);
nand U6395 (N_6395,N_1537,N_4531);
and U6396 (N_6396,N_4198,N_545);
nor U6397 (N_6397,N_3242,N_4225);
or U6398 (N_6398,N_2009,N_624);
and U6399 (N_6399,N_1202,N_3899);
and U6400 (N_6400,N_3056,N_124);
or U6401 (N_6401,N_4770,N_4720);
or U6402 (N_6402,N_2049,N_3412);
nor U6403 (N_6403,N_1593,N_1885);
nand U6404 (N_6404,N_3148,N_4588);
and U6405 (N_6405,N_191,N_2913);
and U6406 (N_6406,N_3991,N_4044);
nand U6407 (N_6407,N_2840,N_3031);
and U6408 (N_6408,N_209,N_3005);
nor U6409 (N_6409,N_3865,N_1972);
or U6410 (N_6410,N_2286,N_2723);
or U6411 (N_6411,N_4586,N_4263);
nand U6412 (N_6412,N_2747,N_1439);
nand U6413 (N_6413,N_4389,N_250);
or U6414 (N_6414,N_3875,N_3339);
nor U6415 (N_6415,N_2680,N_1912);
nor U6416 (N_6416,N_4231,N_1743);
or U6417 (N_6417,N_4162,N_2027);
or U6418 (N_6418,N_3343,N_3912);
xor U6419 (N_6419,N_112,N_4297);
nor U6420 (N_6420,N_3577,N_4055);
and U6421 (N_6421,N_1569,N_2896);
and U6422 (N_6422,N_3864,N_1918);
or U6423 (N_6423,N_2992,N_4333);
and U6424 (N_6424,N_4081,N_4277);
nor U6425 (N_6425,N_364,N_3208);
nand U6426 (N_6426,N_1521,N_1556);
nor U6427 (N_6427,N_4211,N_3843);
nand U6428 (N_6428,N_1982,N_3968);
and U6429 (N_6429,N_3821,N_2894);
nand U6430 (N_6430,N_3648,N_3462);
nand U6431 (N_6431,N_3645,N_4707);
nor U6432 (N_6432,N_4927,N_4773);
and U6433 (N_6433,N_1016,N_2952);
or U6434 (N_6434,N_3336,N_2931);
nor U6435 (N_6435,N_4056,N_634);
or U6436 (N_6436,N_2360,N_3484);
or U6437 (N_6437,N_2584,N_2020);
or U6438 (N_6438,N_2644,N_1986);
nor U6439 (N_6439,N_1677,N_3376);
nand U6440 (N_6440,N_1325,N_4232);
nand U6441 (N_6441,N_1087,N_602);
nor U6442 (N_6442,N_1213,N_120);
nand U6443 (N_6443,N_685,N_136);
nand U6444 (N_6444,N_2364,N_4431);
and U6445 (N_6445,N_1864,N_2346);
nand U6446 (N_6446,N_1411,N_3174);
and U6447 (N_6447,N_3671,N_4774);
or U6448 (N_6448,N_2422,N_4633);
and U6449 (N_6449,N_4329,N_4833);
nor U6450 (N_6450,N_2386,N_777);
nor U6451 (N_6451,N_4985,N_1155);
nand U6452 (N_6452,N_2355,N_1737);
or U6453 (N_6453,N_4036,N_1228);
and U6454 (N_6454,N_3389,N_137);
nor U6455 (N_6455,N_3003,N_1783);
nand U6456 (N_6456,N_1271,N_3919);
or U6457 (N_6457,N_2413,N_1583);
nand U6458 (N_6458,N_2998,N_2507);
and U6459 (N_6459,N_1077,N_4129);
nand U6460 (N_6460,N_1955,N_29);
nand U6461 (N_6461,N_2445,N_2554);
nor U6462 (N_6462,N_4041,N_2939);
or U6463 (N_6463,N_3627,N_3232);
and U6464 (N_6464,N_1804,N_2717);
and U6465 (N_6465,N_4492,N_862);
or U6466 (N_6466,N_2244,N_4771);
nor U6467 (N_6467,N_1554,N_1317);
or U6468 (N_6468,N_3902,N_2695);
and U6469 (N_6469,N_4613,N_6);
and U6470 (N_6470,N_188,N_3262);
or U6471 (N_6471,N_3905,N_1602);
and U6472 (N_6472,N_3303,N_4979);
nand U6473 (N_6473,N_464,N_4643);
or U6474 (N_6474,N_4465,N_4011);
xor U6475 (N_6475,N_704,N_2834);
or U6476 (N_6476,N_4676,N_1116);
or U6477 (N_6477,N_4507,N_4037);
and U6478 (N_6478,N_2092,N_4815);
nor U6479 (N_6479,N_2301,N_1855);
nand U6480 (N_6480,N_1099,N_1936);
or U6481 (N_6481,N_1750,N_1576);
or U6482 (N_6482,N_2975,N_769);
and U6483 (N_6483,N_4385,N_4826);
nand U6484 (N_6484,N_3984,N_4737);
or U6485 (N_6485,N_561,N_1483);
and U6486 (N_6486,N_1278,N_4516);
or U6487 (N_6487,N_228,N_3582);
or U6488 (N_6488,N_931,N_751);
or U6489 (N_6489,N_1308,N_4900);
or U6490 (N_6490,N_451,N_1000);
or U6491 (N_6491,N_3117,N_4726);
nand U6492 (N_6492,N_4649,N_1474);
xnor U6493 (N_6493,N_1577,N_1480);
and U6494 (N_6494,N_1609,N_293);
and U6495 (N_6495,N_1540,N_109);
and U6496 (N_6496,N_2078,N_741);
and U6497 (N_6497,N_1476,N_1860);
or U6498 (N_6498,N_690,N_4558);
nand U6499 (N_6499,N_1693,N_3660);
and U6500 (N_6500,N_1193,N_4695);
and U6501 (N_6501,N_2858,N_3050);
nor U6502 (N_6502,N_3983,N_3641);
and U6503 (N_6503,N_1981,N_3330);
or U6504 (N_6504,N_3459,N_503);
or U6505 (N_6505,N_739,N_754);
or U6506 (N_6506,N_3550,N_1450);
nand U6507 (N_6507,N_2852,N_251);
nor U6508 (N_6508,N_3846,N_4671);
and U6509 (N_6509,N_439,N_3666);
nor U6510 (N_6510,N_514,N_4866);
and U6511 (N_6511,N_4161,N_867);
nand U6512 (N_6512,N_4568,N_341);
and U6513 (N_6513,N_1888,N_3824);
and U6514 (N_6514,N_1352,N_4344);
nand U6515 (N_6515,N_1672,N_196);
nor U6516 (N_6516,N_1368,N_3004);
and U6517 (N_6517,N_359,N_1091);
and U6518 (N_6518,N_724,N_4585);
nor U6519 (N_6519,N_3175,N_4612);
or U6520 (N_6520,N_3952,N_4680);
nor U6521 (N_6521,N_2642,N_2488);
nor U6522 (N_6522,N_3665,N_43);
nor U6523 (N_6523,N_2671,N_3891);
nand U6524 (N_6524,N_3164,N_1505);
nor U6525 (N_6525,N_4843,N_639);
and U6526 (N_6526,N_1814,N_3647);
or U6527 (N_6527,N_3237,N_333);
and U6528 (N_6528,N_709,N_3699);
and U6529 (N_6529,N_4057,N_1653);
nand U6530 (N_6530,N_2285,N_921);
xnor U6531 (N_6531,N_3721,N_2128);
nor U6532 (N_6532,N_4432,N_2213);
nor U6533 (N_6533,N_870,N_3878);
and U6534 (N_6534,N_3801,N_1454);
or U6535 (N_6535,N_539,N_3197);
nand U6536 (N_6536,N_4798,N_1707);
nor U6537 (N_6537,N_3028,N_70);
nand U6538 (N_6538,N_2462,N_1502);
nand U6539 (N_6539,N_45,N_2870);
or U6540 (N_6540,N_3523,N_982);
and U6541 (N_6541,N_622,N_3995);
nand U6542 (N_6542,N_1968,N_3650);
or U6543 (N_6543,N_4546,N_3255);
nor U6544 (N_6544,N_600,N_499);
nand U6545 (N_6545,N_4363,N_646);
nand U6546 (N_6546,N_197,N_1496);
nand U6547 (N_6547,N_960,N_2105);
and U6548 (N_6548,N_2113,N_552);
nand U6549 (N_6549,N_3813,N_616);
and U6550 (N_6550,N_1181,N_211);
or U6551 (N_6551,N_1951,N_3526);
nor U6552 (N_6552,N_1255,N_3234);
nand U6553 (N_6553,N_4244,N_1149);
nand U6554 (N_6554,N_2416,N_572);
nand U6555 (N_6555,N_4738,N_687);
nor U6556 (N_6556,N_2223,N_1661);
or U6557 (N_6557,N_3536,N_4450);
or U6558 (N_6558,N_3548,N_3730);
nand U6559 (N_6559,N_2969,N_4020);
and U6560 (N_6560,N_4637,N_3248);
nand U6561 (N_6561,N_2071,N_3822);
nor U6562 (N_6562,N_474,N_2398);
and U6563 (N_6563,N_1038,N_3442);
and U6564 (N_6564,N_549,N_342);
nand U6565 (N_6565,N_1944,N_3918);
nand U6566 (N_6566,N_1344,N_266);
nor U6567 (N_6567,N_2189,N_168);
or U6568 (N_6568,N_1092,N_4752);
nor U6569 (N_6569,N_2166,N_2976);
nand U6570 (N_6570,N_2268,N_2283);
and U6571 (N_6571,N_1631,N_1946);
or U6572 (N_6572,N_2758,N_2708);
or U6573 (N_6573,N_2961,N_1171);
and U6574 (N_6574,N_3083,N_2441);
or U6575 (N_6575,N_418,N_2844);
and U6576 (N_6576,N_1780,N_3817);
or U6577 (N_6577,N_2867,N_1950);
nor U6578 (N_6578,N_291,N_2974);
nor U6579 (N_6579,N_4937,N_1746);
nor U6580 (N_6580,N_2110,N_4661);
xor U6581 (N_6581,N_1164,N_3065);
or U6582 (N_6582,N_4495,N_1075);
or U6583 (N_6583,N_640,N_2949);
and U6584 (N_6584,N_3261,N_4033);
or U6585 (N_6585,N_1725,N_3359);
and U6586 (N_6586,N_1358,N_2562);
nand U6587 (N_6587,N_1665,N_2291);
and U6588 (N_6588,N_2409,N_4758);
or U6589 (N_6589,N_2308,N_2337);
or U6590 (N_6590,N_3534,N_94);
and U6591 (N_6591,N_2191,N_52);
or U6592 (N_6592,N_2122,N_1962);
and U6593 (N_6593,N_2043,N_4128);
nand U6594 (N_6594,N_1699,N_2865);
nor U6595 (N_6595,N_825,N_3222);
or U6596 (N_6596,N_517,N_1432);
and U6597 (N_6597,N_1104,N_4258);
or U6598 (N_6598,N_4218,N_3636);
nor U6599 (N_6599,N_3853,N_3895);
and U6600 (N_6600,N_4864,N_2653);
nor U6601 (N_6601,N_398,N_4533);
and U6602 (N_6602,N_366,N_4476);
and U6603 (N_6603,N_4851,N_806);
nor U6604 (N_6604,N_541,N_2173);
and U6605 (N_6605,N_733,N_160);
nand U6606 (N_6606,N_3434,N_906);
or U6607 (N_6607,N_1452,N_2006);
nand U6608 (N_6608,N_3236,N_4150);
nand U6609 (N_6609,N_2379,N_2703);
nand U6610 (N_6610,N_2097,N_1820);
nand U6611 (N_6611,N_190,N_1494);
nor U6612 (N_6612,N_1816,N_3672);
nand U6613 (N_6613,N_126,N_3976);
nor U6614 (N_6614,N_3411,N_2604);
nand U6615 (N_6615,N_3187,N_3101);
nand U6616 (N_6616,N_947,N_1322);
nor U6617 (N_6617,N_4310,N_2497);
or U6618 (N_6618,N_2347,N_372);
nand U6619 (N_6619,N_3375,N_4308);
and U6620 (N_6620,N_1279,N_1049);
and U6621 (N_6621,N_4962,N_649);
or U6622 (N_6622,N_2058,N_1273);
or U6623 (N_6623,N_1192,N_4704);
and U6624 (N_6624,N_907,N_4548);
nand U6625 (N_6625,N_3167,N_412);
and U6626 (N_6626,N_305,N_4848);
nand U6627 (N_6627,N_4913,N_361);
nor U6628 (N_6628,N_748,N_2521);
nand U6629 (N_6629,N_4610,N_3600);
nand U6630 (N_6630,N_3711,N_3703);
nand U6631 (N_6631,N_161,N_3994);
or U6632 (N_6632,N_33,N_351);
or U6633 (N_6633,N_3738,N_3719);
and U6634 (N_6634,N_4376,N_248);
and U6635 (N_6635,N_2362,N_1246);
nand U6636 (N_6636,N_2645,N_726);
nand U6637 (N_6637,N_426,N_2835);
and U6638 (N_6638,N_2363,N_944);
or U6639 (N_6639,N_1953,N_2532);
nor U6640 (N_6640,N_3349,N_2339);
nand U6641 (N_6641,N_2505,N_76);
nand U6642 (N_6642,N_1441,N_1709);
nand U6643 (N_6643,N_272,N_103);
or U6644 (N_6644,N_4651,N_3807);
nor U6645 (N_6645,N_4239,N_4893);
nor U6646 (N_6646,N_3606,N_3753);
nand U6647 (N_6647,N_1052,N_1451);
nand U6648 (N_6648,N_1605,N_2821);
and U6649 (N_6649,N_3541,N_2779);
or U6650 (N_6650,N_4076,N_4987);
nor U6651 (N_6651,N_3432,N_757);
and U6652 (N_6652,N_1288,N_3116);
nor U6653 (N_6653,N_4137,N_1188);
and U6654 (N_6654,N_1403,N_1081);
and U6655 (N_6655,N_4373,N_2555);
nor U6656 (N_6656,N_3668,N_815);
nor U6657 (N_6657,N_3595,N_3126);
and U6658 (N_6658,N_62,N_4264);
or U6659 (N_6659,N_3023,N_98);
and U6660 (N_6660,N_706,N_1683);
and U6661 (N_6661,N_728,N_4523);
nor U6662 (N_6662,N_2150,N_2025);
nand U6663 (N_6663,N_4542,N_131);
xnor U6664 (N_6664,N_390,N_2761);
and U6665 (N_6665,N_3862,N_755);
nand U6666 (N_6666,N_1618,N_3093);
and U6667 (N_6667,N_2648,N_1973);
nand U6668 (N_6668,N_4717,N_1598);
nand U6669 (N_6669,N_3935,N_2094);
and U6670 (N_6670,N_4824,N_598);
and U6671 (N_6671,N_2625,N_1210);
nand U6672 (N_6672,N_2417,N_1848);
nand U6673 (N_6673,N_446,N_3734);
nand U6674 (N_6674,N_860,N_2736);
and U6675 (N_6675,N_4935,N_1008);
or U6676 (N_6676,N_1645,N_4367);
nand U6677 (N_6677,N_1035,N_1478);
or U6678 (N_6678,N_3408,N_286);
nor U6679 (N_6679,N_3267,N_4307);
or U6680 (N_6680,N_672,N_1464);
nor U6681 (N_6681,N_262,N_2519);
nor U6682 (N_6682,N_1013,N_4068);
nor U6683 (N_6683,N_4085,N_1263);
and U6684 (N_6684,N_2205,N_1129);
or U6685 (N_6685,N_313,N_1137);
nor U6686 (N_6686,N_486,N_1497);
or U6687 (N_6687,N_3982,N_4836);
nor U6688 (N_6688,N_1063,N_845);
or U6689 (N_6689,N_4716,N_4452);
nand U6690 (N_6690,N_1068,N_2187);
nand U6691 (N_6691,N_3341,N_4562);
and U6692 (N_6692,N_716,N_4988);
nor U6693 (N_6693,N_3414,N_4589);
and U6694 (N_6694,N_3769,N_3514);
nor U6695 (N_6695,N_4986,N_2881);
and U6696 (N_6696,N_1764,N_3157);
and U6697 (N_6697,N_4093,N_771);
nand U6698 (N_6698,N_3316,N_468);
or U6699 (N_6699,N_2050,N_2246);
or U6700 (N_6700,N_3673,N_2866);
and U6701 (N_6701,N_1826,N_4503);
nor U6702 (N_6702,N_3307,N_316);
or U6703 (N_6703,N_2265,N_3265);
nand U6704 (N_6704,N_299,N_4291);
or U6705 (N_6705,N_4620,N_1843);
and U6706 (N_6706,N_4303,N_4520);
and U6707 (N_6707,N_516,N_331);
nor U6708 (N_6708,N_1882,N_4001);
and U6709 (N_6709,N_1256,N_2582);
or U6710 (N_6710,N_4121,N_2766);
nor U6711 (N_6711,N_981,N_581);
or U6712 (N_6712,N_2801,N_4691);
nand U6713 (N_6713,N_2119,N_1248);
nand U6714 (N_6714,N_1565,N_2314);
or U6715 (N_6715,N_150,N_1017);
nand U6716 (N_6716,N_3368,N_729);
nand U6717 (N_6717,N_1777,N_3041);
nor U6718 (N_6718,N_2875,N_2284);
or U6719 (N_6719,N_829,N_1613);
and U6720 (N_6720,N_100,N_3427);
nand U6721 (N_6721,N_4206,N_1201);
nor U6722 (N_6722,N_4679,N_2855);
and U6723 (N_6723,N_1821,N_3869);
nand U6724 (N_6724,N_315,N_2419);
or U6725 (N_6725,N_1788,N_200);
nor U6726 (N_6726,N_2620,N_2449);
nand U6727 (N_6727,N_3152,N_4123);
or U6728 (N_6728,N_4223,N_3625);
nand U6729 (N_6729,N_4739,N_734);
or U6730 (N_6730,N_4659,N_4960);
nor U6731 (N_6731,N_4316,N_3060);
or U6732 (N_6732,N_138,N_2214);
nor U6733 (N_6733,N_1698,N_1224);
nor U6734 (N_6734,N_1418,N_3362);
xor U6735 (N_6735,N_2003,N_3849);
nor U6736 (N_6736,N_2390,N_294);
and U6737 (N_6737,N_4077,N_2275);
nand U6738 (N_6738,N_1948,N_3465);
and U6739 (N_6739,N_2959,N_2603);
nor U6740 (N_6740,N_192,N_3724);
or U6741 (N_6741,N_1311,N_1429);
nor U6742 (N_6742,N_3883,N_1952);
and U6743 (N_6743,N_4782,N_1744);
or U6744 (N_6744,N_3014,N_2751);
or U6745 (N_6745,N_3720,N_1378);
and U6746 (N_6746,N_1708,N_4896);
and U6747 (N_6747,N_3777,N_2421);
nand U6748 (N_6748,N_2935,N_713);
and U6749 (N_6749,N_938,N_4095);
nor U6750 (N_6750,N_2182,N_2427);
nor U6751 (N_6751,N_4138,N_2530);
nor U6752 (N_6752,N_926,N_756);
or U6753 (N_6753,N_1691,N_349);
nand U6754 (N_6754,N_246,N_4934);
and U6755 (N_6755,N_817,N_2694);
and U6756 (N_6756,N_4642,N_1546);
nand U6757 (N_6757,N_2509,N_1988);
or U6758 (N_6758,N_3016,N_2877);
nand U6759 (N_6759,N_3125,N_3901);
nor U6760 (N_6760,N_1310,N_832);
and U6761 (N_6761,N_3214,N_3069);
nand U6762 (N_6762,N_3226,N_3493);
or U6763 (N_6763,N_4040,N_3950);
nor U6764 (N_6764,N_4819,N_932);
nor U6765 (N_6765,N_1700,N_4181);
nor U6766 (N_6766,N_4007,N_3217);
and U6767 (N_6767,N_1806,N_2466);
or U6768 (N_6768,N_88,N_4241);
and U6769 (N_6769,N_4800,N_2412);
nand U6770 (N_6770,N_4184,N_4547);
and U6771 (N_6771,N_1937,N_4115);
nand U6772 (N_6772,N_3473,N_3659);
and U6773 (N_6773,N_3763,N_4397);
or U6774 (N_6774,N_4051,N_1409);
and U6775 (N_6775,N_495,N_3196);
and U6776 (N_6776,N_2263,N_953);
or U6777 (N_6777,N_597,N_1934);
nand U6778 (N_6778,N_3021,N_1597);
or U6779 (N_6779,N_3911,N_1486);
and U6780 (N_6780,N_1131,N_2457);
nand U6781 (N_6781,N_4550,N_3958);
nor U6782 (N_6782,N_4100,N_1379);
nor U6783 (N_6783,N_3977,N_3772);
nor U6784 (N_6784,N_92,N_4499);
or U6785 (N_6785,N_2101,N_2383);
or U6786 (N_6786,N_2752,N_3833);
and U6787 (N_6787,N_4775,N_2280);
nor U6788 (N_6788,N_2023,N_1696);
nand U6789 (N_6789,N_2527,N_4444);
or U6790 (N_6790,N_4205,N_922);
nand U6791 (N_6791,N_4509,N_3744);
nand U6792 (N_6792,N_472,N_2552);
nor U6793 (N_6793,N_3518,N_3147);
nor U6794 (N_6794,N_732,N_3732);
or U6795 (N_6795,N_776,N_3331);
nor U6796 (N_6796,N_2589,N_4054);
nand U6797 (N_6797,N_4426,N_252);
nor U6798 (N_6798,N_145,N_491);
nand U6799 (N_6799,N_2366,N_2613);
or U6800 (N_6800,N_933,N_2046);
and U6801 (N_6801,N_2661,N_1870);
nor U6802 (N_6802,N_3404,N_311);
and U6803 (N_6803,N_553,N_2662);
nor U6804 (N_6804,N_344,N_1037);
nand U6805 (N_6805,N_1503,N_25);
nor U6806 (N_6806,N_2932,N_93);
nor U6807 (N_6807,N_1616,N_1022);
nor U6808 (N_6808,N_3978,N_3424);
nand U6809 (N_6809,N_3565,N_4698);
nor U6810 (N_6810,N_2585,N_296);
nand U6811 (N_6811,N_4178,N_1825);
or U6812 (N_6812,N_2320,N_2911);
nand U6813 (N_6813,N_4436,N_4513);
nand U6814 (N_6814,N_3273,N_2514);
or U6815 (N_6815,N_2260,N_2442);
and U6816 (N_6816,N_525,N_1203);
nand U6817 (N_6817,N_2079,N_3296);
nor U6818 (N_6818,N_1977,N_3960);
nand U6819 (N_6819,N_2461,N_692);
or U6820 (N_6820,N_1114,N_2759);
nor U6821 (N_6821,N_1319,N_4339);
or U6822 (N_6822,N_1341,N_3580);
or U6823 (N_6823,N_4147,N_1372);
or U6824 (N_6824,N_1366,N_3092);
nor U6825 (N_6825,N_1307,N_1165);
nor U6826 (N_6826,N_3837,N_958);
and U6827 (N_6827,N_984,N_1907);
and U6828 (N_6828,N_4132,N_1630);
and U6829 (N_6829,N_1742,N_4070);
and U6830 (N_6830,N_376,N_1397);
nand U6831 (N_6831,N_1223,N_4505);
nand U6832 (N_6832,N_4140,N_2034);
or U6833 (N_6833,N_343,N_879);
and U6834 (N_6834,N_4293,N_1549);
and U6835 (N_6835,N_171,N_1904);
nor U6836 (N_6836,N_3863,N_854);
and U6837 (N_6837,N_1088,N_4395);
nand U6838 (N_6838,N_3585,N_1388);
nand U6839 (N_6839,N_3681,N_2153);
nand U6840 (N_6840,N_966,N_1214);
and U6841 (N_6841,N_2005,N_204);
or U6842 (N_6842,N_2788,N_1316);
nor U6843 (N_6843,N_3702,N_1812);
and U6844 (N_6844,N_2506,N_3969);
or U6845 (N_6845,N_2659,N_1128);
and U6846 (N_6846,N_861,N_1751);
and U6847 (N_6847,N_2776,N_1169);
nand U6848 (N_6848,N_4394,N_2770);
or U6849 (N_6849,N_4521,N_3440);
nand U6850 (N_6850,N_113,N_2951);
nand U6851 (N_6851,N_325,N_2282);
and U6852 (N_6852,N_701,N_3759);
and U6853 (N_6853,N_2272,N_2067);
and U6854 (N_6854,N_2353,N_2937);
nor U6855 (N_6855,N_542,N_674);
nor U6856 (N_6856,N_2255,N_3616);
nor U6857 (N_6857,N_3722,N_4811);
and U6858 (N_6858,N_4563,N_1281);
or U6859 (N_6859,N_4907,N_521);
nand U6860 (N_6860,N_1033,N_1112);
and U6861 (N_6861,N_1916,N_790);
xor U6862 (N_6862,N_253,N_3176);
nor U6863 (N_6863,N_2621,N_4201);
xnor U6864 (N_6864,N_1487,N_2605);
or U6865 (N_6865,N_3961,N_2579);
or U6866 (N_6866,N_3211,N_4690);
or U6867 (N_6867,N_1258,N_259);
nor U6868 (N_6868,N_3168,N_2368);
nand U6869 (N_6869,N_2077,N_2938);
nor U6870 (N_6870,N_1143,N_1896);
nor U6871 (N_6871,N_281,N_3502);
nand U6872 (N_6872,N_4997,N_407);
nor U6873 (N_6873,N_2185,N_1664);
nand U6874 (N_6874,N_3015,N_2090);
and U6875 (N_6875,N_4787,N_1448);
and U6876 (N_6876,N_4890,N_2469);
nor U6877 (N_6877,N_3249,N_2226);
nand U6878 (N_6878,N_1384,N_484);
or U6879 (N_6879,N_1290,N_3099);
nor U6880 (N_6880,N_4375,N_735);
nor U6881 (N_6881,N_4832,N_3200);
and U6882 (N_6882,N_1394,N_1682);
and U6883 (N_6883,N_669,N_2477);
nor U6884 (N_6884,N_4064,N_3131);
nand U6885 (N_6885,N_2264,N_3193);
or U6886 (N_6886,N_1594,N_2988);
and U6887 (N_6887,N_4032,N_4580);
nand U6888 (N_6888,N_4532,N_4554);
nand U6889 (N_6889,N_4812,N_4862);
or U6890 (N_6890,N_719,N_4404);
or U6891 (N_6891,N_4995,N_1985);
nand U6892 (N_6892,N_4256,N_2256);
nand U6893 (N_6893,N_2768,N_454);
nor U6894 (N_6894,N_4682,N_3351);
or U6895 (N_6895,N_1928,N_3385);
or U6896 (N_6896,N_2773,N_4318);
or U6897 (N_6897,N_2721,N_3850);
nand U6898 (N_6898,N_255,N_431);
or U6899 (N_6899,N_2999,N_2547);
nor U6900 (N_6900,N_3692,N_2443);
or U6901 (N_6901,N_1716,N_3870);
and U6902 (N_6902,N_3906,N_963);
nand U6903 (N_6903,N_1479,N_1805);
nor U6904 (N_6904,N_2235,N_216);
nand U6905 (N_6905,N_4938,N_2010);
nand U6906 (N_6906,N_3340,N_556);
or U6907 (N_6907,N_896,N_908);
nand U6908 (N_6908,N_3669,N_4462);
and U6909 (N_6909,N_4750,N_1983);
nor U6910 (N_6910,N_4641,N_977);
nand U6911 (N_6911,N_3642,N_4148);
nand U6912 (N_6912,N_408,N_4204);
and U6913 (N_6913,N_595,N_4387);
and U6914 (N_6914,N_3457,N_4667);
or U6915 (N_6915,N_2709,N_3792);
and U6916 (N_6916,N_4021,N_178);
nand U6917 (N_6917,N_2565,N_4199);
nor U6918 (N_6918,N_785,N_2843);
nor U6919 (N_6919,N_2914,N_2068);
and U6920 (N_6920,N_2206,N_1216);
and U6921 (N_6921,N_494,N_3856);
nor U6922 (N_6922,N_3428,N_1208);
nand U6923 (N_6923,N_42,N_3654);
nand U6924 (N_6924,N_965,N_1225);
nor U6925 (N_6925,N_4298,N_3592);
and U6926 (N_6926,N_386,N_1185);
nor U6927 (N_6927,N_2795,N_738);
and U6928 (N_6928,N_363,N_2313);
nor U6929 (N_6929,N_991,N_4537);
and U6930 (N_6930,N_1768,N_1510);
or U6931 (N_6931,N_1234,N_2599);
nand U6932 (N_6932,N_1787,N_2432);
nand U6933 (N_6933,N_3386,N_2279);
and U6934 (N_6934,N_1350,N_3975);
nor U6935 (N_6935,N_47,N_1481);
nor U6936 (N_6936,N_4487,N_4177);
nand U6937 (N_6937,N_4609,N_2141);
and U6938 (N_6938,N_775,N_4729);
and U6939 (N_6939,N_1078,N_750);
nor U6940 (N_6940,N_3685,N_4489);
or U6941 (N_6941,N_2227,N_1415);
nor U6942 (N_6942,N_219,N_202);
or U6943 (N_6943,N_1312,N_2237);
or U6944 (N_6944,N_1638,N_3800);
or U6945 (N_6945,N_4855,N_2489);
xor U6946 (N_6946,N_3676,N_4321);
nand U6947 (N_6947,N_1733,N_2936);
nor U6948 (N_6948,N_4861,N_2378);
and U6949 (N_6949,N_4061,N_4014);
and U6950 (N_6950,N_4338,N_1735);
or U6951 (N_6951,N_1044,N_2790);
nor U6952 (N_6952,N_461,N_3337);
or U6953 (N_6953,N_3106,N_576);
nand U6954 (N_6954,N_3035,N_3400);
nand U6955 (N_6955,N_1762,N_3783);
or U6956 (N_6956,N_2250,N_3811);
nor U6957 (N_6957,N_2856,N_399);
nand U6958 (N_6958,N_4801,N_1120);
or U6959 (N_6959,N_1547,N_643);
and U6960 (N_6960,N_4662,N_4894);
or U6961 (N_6961,N_2979,N_1567);
nand U6962 (N_6962,N_1795,N_4715);
nand U6963 (N_6963,N_650,N_226);
nand U6964 (N_6964,N_2247,N_3281);
nor U6965 (N_6965,N_212,N_641);
or U6966 (N_6966,N_3847,N_1838);
or U6967 (N_6967,N_4456,N_3287);
and U6968 (N_6968,N_4096,N_2060);
and U6969 (N_6969,N_828,N_3916);
and U6970 (N_6970,N_2909,N_3403);
nand U6971 (N_6971,N_4074,N_856);
nand U6972 (N_6972,N_1873,N_537);
nor U6973 (N_6973,N_1663,N_3559);
or U6974 (N_6974,N_279,N_2070);
or U6975 (N_6975,N_1706,N_4407);
and U6976 (N_6976,N_1026,N_2149);
and U6977 (N_6977,N_1291,N_911);
nand U6978 (N_6978,N_3840,N_919);
or U6979 (N_6979,N_3452,N_3857);
nor U6980 (N_6980,N_1493,N_4322);
nand U6981 (N_6981,N_2556,N_1790);
or U6982 (N_6982,N_3038,N_2485);
nor U6983 (N_6983,N_4675,N_1710);
and U6984 (N_6984,N_3020,N_2373);
or U6985 (N_6985,N_2196,N_4186);
nand U6986 (N_6986,N_3480,N_3415);
nand U6987 (N_6987,N_2194,N_3921);
nor U6988 (N_6988,N_2630,N_2854);
and U6989 (N_6989,N_2825,N_3543);
and U6990 (N_6990,N_4746,N_2163);
and U6991 (N_6991,N_1558,N_956);
and U6992 (N_6992,N_10,N_2299);
nor U6993 (N_6993,N_4410,N_369);
or U6994 (N_6994,N_4535,N_1802);
nor U6995 (N_6995,N_4839,N_2199);
nor U6996 (N_6996,N_1364,N_269);
or U6997 (N_6997,N_3266,N_1259);
and U6998 (N_6998,N_2512,N_1488);
nor U6999 (N_6999,N_2177,N_3317);
and U7000 (N_7000,N_527,N_3851);
nand U7001 (N_7001,N_3458,N_3678);
and U7002 (N_7002,N_3635,N_82);
or U7003 (N_7003,N_4867,N_2520);
or U7004 (N_7004,N_700,N_2455);
nand U7005 (N_7005,N_2147,N_2252);
nand U7006 (N_7006,N_244,N_1349);
or U7007 (N_7007,N_1553,N_3713);
or U7008 (N_7008,N_2157,N_4237);
nand U7009 (N_7009,N_4213,N_4071);
nor U7010 (N_7010,N_2602,N_4573);
nand U7011 (N_7011,N_4844,N_2240);
and U7012 (N_7012,N_3084,N_1118);
and U7013 (N_7013,N_3537,N_939);
nor U7014 (N_7014,N_3225,N_4477);
and U7015 (N_7015,N_4708,N_2686);
and U7016 (N_7016,N_3380,N_3886);
and U7017 (N_7017,N_3517,N_4086);
nand U7018 (N_7018,N_3696,N_4190);
nand U7019 (N_7019,N_4511,N_1852);
and U7020 (N_7020,N_3754,N_3270);
nand U7021 (N_7021,N_4921,N_4999);
or U7022 (N_7022,N_663,N_1818);
nand U7023 (N_7023,N_4101,N_2995);
nor U7024 (N_7024,N_3974,N_206);
nor U7025 (N_7025,N_3447,N_3929);
nor U7026 (N_7026,N_3845,N_3758);
or U7027 (N_7027,N_68,N_4326);
and U7028 (N_7028,N_2957,N_3540);
and U7029 (N_7029,N_1096,N_721);
and U7030 (N_7030,N_2168,N_3374);
and U7031 (N_7031,N_2318,N_2689);
nor U7032 (N_7032,N_3372,N_3358);
nand U7033 (N_7033,N_927,N_3453);
nor U7034 (N_7034,N_1996,N_3882);
or U7035 (N_7035,N_1641,N_489);
and U7036 (N_7036,N_1644,N_1688);
nand U7037 (N_7037,N_389,N_2987);
nand U7038 (N_7038,N_3363,N_1604);
nor U7039 (N_7039,N_1831,N_703);
nand U7040 (N_7040,N_2467,N_4747);
and U7041 (N_7041,N_2544,N_3740);
and U7042 (N_7042,N_3573,N_924);
nand U7043 (N_7043,N_4330,N_2597);
and U7044 (N_7044,N_551,N_1150);
nand U7045 (N_7045,N_2117,N_3680);
nand U7046 (N_7046,N_2831,N_1971);
or U7047 (N_7047,N_2963,N_579);
xnor U7048 (N_7048,N_2021,N_2798);
nor U7049 (N_7049,N_3112,N_4872);
nand U7050 (N_7050,N_2309,N_1839);
and U7051 (N_7051,N_4598,N_3165);
or U7052 (N_7052,N_533,N_243);
or U7053 (N_7053,N_3183,N_2566);
or U7054 (N_7054,N_946,N_1891);
nand U7055 (N_7055,N_3907,N_4491);
or U7056 (N_7056,N_3788,N_2685);
or U7057 (N_7057,N_210,N_4275);
nand U7058 (N_7058,N_425,N_816);
nand U7059 (N_7059,N_3602,N_4518);
and U7060 (N_7060,N_601,N_1175);
and U7061 (N_7061,N_1036,N_3218);
nand U7062 (N_7062,N_2411,N_4882);
and U7063 (N_7063,N_3098,N_3128);
or U7064 (N_7064,N_218,N_48);
or U7065 (N_7065,N_4217,N_3327);
or U7066 (N_7066,N_2053,N_992);
nand U7067 (N_7067,N_1538,N_2710);
and U7068 (N_7068,N_2904,N_459);
and U7069 (N_7069,N_3542,N_3928);
nor U7070 (N_7070,N_435,N_4153);
and U7071 (N_7071,N_2849,N_4596);
nand U7072 (N_7072,N_2977,N_599);
nand U7073 (N_7073,N_3809,N_2859);
and U7074 (N_7074,N_3319,N_3127);
nand U7075 (N_7075,N_3687,N_4606);
or U7076 (N_7076,N_658,N_1920);
or U7077 (N_7077,N_3325,N_3609);
and U7078 (N_7078,N_8,N_818);
nor U7079 (N_7079,N_295,N_881);
nor U7080 (N_7080,N_3186,N_4807);
and U7081 (N_7081,N_2134,N_3243);
nor U7082 (N_7082,N_1959,N_4448);
nor U7083 (N_7083,N_2072,N_3392);
or U7084 (N_7084,N_354,N_3943);
nor U7085 (N_7085,N_1634,N_2000);
nand U7086 (N_7086,N_857,N_467);
nor U7087 (N_7087,N_3632,N_505);
nand U7088 (N_7088,N_2012,N_2984);
and U7089 (N_7089,N_4587,N_3701);
nor U7090 (N_7090,N_3455,N_4810);
nand U7091 (N_7091,N_1779,N_3971);
nor U7092 (N_7092,N_157,N_787);
and U7093 (N_7093,N_4073,N_4176);
or U7094 (N_7094,N_1110,N_747);
nor U7095 (N_7095,N_4799,N_1094);
nand U7096 (N_7096,N_797,N_1287);
or U7097 (N_7097,N_256,N_350);
or U7098 (N_7098,N_3626,N_456);
nand U7099 (N_7099,N_1065,N_905);
or U7100 (N_7100,N_4226,N_3778);
nor U7101 (N_7101,N_2741,N_2891);
or U7102 (N_7102,N_2498,N_483);
nor U7103 (N_7103,N_2080,N_2559);
nand U7104 (N_7104,N_4325,N_567);
nor U7105 (N_7105,N_2176,N_169);
or U7106 (N_7106,N_1921,N_2019);
and U7107 (N_7107,N_3528,N_1195);
nand U7108 (N_7108,N_2098,N_2956);
nand U7109 (N_7109,N_813,N_3729);
and U7110 (N_7110,N_4109,N_4956);
nand U7111 (N_7111,N_80,N_1840);
and U7112 (N_7112,N_117,N_3923);
or U7113 (N_7113,N_1899,N_1828);
nand U7114 (N_7114,N_4360,N_677);
and U7115 (N_7115,N_220,N_3066);
or U7116 (N_7116,N_1490,N_2828);
and U7117 (N_7117,N_3429,N_513);
nor U7118 (N_7118,N_4948,N_3067);
nor U7119 (N_7119,N_2775,N_3027);
nor U7120 (N_7120,N_694,N_3593);
and U7121 (N_7121,N_1054,N_1373);
and U7122 (N_7122,N_4591,N_4088);
nand U7123 (N_7123,N_38,N_2302);
or U7124 (N_7124,N_4267,N_167);
nor U7125 (N_7125,N_566,N_2305);
or U7126 (N_7126,N_967,N_3182);
nand U7127 (N_7127,N_4222,N_2837);
and U7128 (N_7128,N_1406,N_1346);
or U7129 (N_7129,N_603,N_2696);
nand U7130 (N_7130,N_3651,N_2845);
or U7131 (N_7131,N_2004,N_479);
and U7132 (N_7132,N_3539,N_4336);
nor U7133 (N_7133,N_1059,N_4996);
nand U7134 (N_7134,N_3762,N_4207);
and U7135 (N_7135,N_827,N_2672);
nor U7136 (N_7136,N_1194,N_3263);
or U7137 (N_7137,N_1090,N_1967);
nand U7138 (N_7138,N_3930,N_891);
nand U7139 (N_7139,N_4869,N_1640);
or U7140 (N_7140,N_1436,N_2745);
nand U7141 (N_7141,N_1222,N_3423);
or U7142 (N_7142,N_4525,N_1238);
nand U7143 (N_7143,N_2052,N_3922);
and U7144 (N_7144,N_3771,N_2407);
nand U7145 (N_7145,N_1163,N_4723);
and U7146 (N_7146,N_4683,N_4572);
nand U7147 (N_7147,N_258,N_4551);
and U7148 (N_7148,N_2627,N_375);
and U7149 (N_7149,N_2450,N_2216);
or U7150 (N_7150,N_1958,N_4688);
nor U7151 (N_7151,N_1905,N_2501);
nor U7152 (N_7152,N_3240,N_4623);
and U7153 (N_7153,N_132,N_4700);
nand U7154 (N_7154,N_4957,N_1062);
nand U7155 (N_7155,N_2031,N_2171);
nand U7156 (N_7156,N_1115,N_1987);
and U7157 (N_7157,N_3146,N_1134);
or U7158 (N_7158,N_697,N_280);
nand U7159 (N_7159,N_2229,N_1402);
nand U7160 (N_7160,N_402,N_3931);
nor U7161 (N_7161,N_3010,N_973);
nor U7162 (N_7162,N_2583,N_3885);
nand U7163 (N_7163,N_885,N_4791);
nor U7164 (N_7164,N_358,N_1586);
and U7165 (N_7165,N_1061,N_4401);
nor U7166 (N_7166,N_901,N_173);
nor U7167 (N_7167,N_778,N_4302);
nand U7168 (N_7168,N_3449,N_524);
nor U7169 (N_7169,N_1018,N_657);
nand U7170 (N_7170,N_4846,N_3034);
or U7171 (N_7171,N_800,N_4817);
or U7172 (N_7172,N_2396,N_3045);
nand U7173 (N_7173,N_794,N_2973);
nor U7174 (N_7174,N_1343,N_340);
or U7175 (N_7175,N_2677,N_4854);
and U7176 (N_7176,N_56,N_1434);
nand U7177 (N_7177,N_4008,N_3202);
nand U7178 (N_7178,N_837,N_1204);
nor U7179 (N_7179,N_3278,N_153);
nand U7180 (N_7180,N_3011,N_107);
and U7181 (N_7181,N_4993,N_434);
nand U7182 (N_7182,N_1121,N_1516);
nand U7183 (N_7183,N_997,N_4282);
nor U7184 (N_7184,N_4597,N_4253);
and U7185 (N_7185,N_1015,N_1552);
or U7186 (N_7186,N_1994,N_2502);
nor U7187 (N_7187,N_1678,N_2231);
or U7188 (N_7188,N_3321,N_4517);
nor U7189 (N_7189,N_2403,N_440);
nor U7190 (N_7190,N_4701,N_3940);
and U7191 (N_7191,N_2483,N_935);
or U7192 (N_7192,N_3836,N_822);
and U7193 (N_7193,N_4331,N_2352);
or U7194 (N_7194,N_3444,N_779);
nand U7195 (N_7195,N_4337,N_2905);
or U7196 (N_7196,N_3675,N_4328);
and U7197 (N_7197,N_4702,N_2001);
or U7198 (N_7198,N_798,N_1857);
nor U7199 (N_7199,N_3420,N_1199);
and U7200 (N_7200,N_1585,N_1427);
and U7201 (N_7201,N_2306,N_1180);
nand U7202 (N_7202,N_945,N_3491);
nand U7203 (N_7203,N_335,N_1801);
or U7204 (N_7204,N_125,N_804);
nand U7205 (N_7205,N_4284,N_4614);
or U7206 (N_7206,N_2303,N_3291);
or U7207 (N_7207,N_4802,N_4157);
and U7208 (N_7208,N_888,N_4742);
or U7209 (N_7209,N_2126,N_765);
or U7210 (N_7210,N_1071,N_321);
nor U7211 (N_7211,N_3607,N_449);
nand U7212 (N_7212,N_3814,N_4494);
or U7213 (N_7213,N_4392,N_170);
or U7214 (N_7214,N_1763,N_3329);
nand U7215 (N_7215,N_635,N_1785);
and U7216 (N_7216,N_1177,N_764);
nand U7217 (N_7217,N_4457,N_2164);
and U7218 (N_7218,N_1894,N_4346);
and U7219 (N_7219,N_2428,N_2691);
or U7220 (N_7220,N_3587,N_1370);
and U7221 (N_7221,N_2290,N_2719);
nor U7222 (N_7222,N_660,N_3286);
or U7223 (N_7223,N_4356,N_2571);
and U7224 (N_7224,N_2160,N_2304);
nor U7225 (N_7225,N_4379,N_1800);
nor U7226 (N_7226,N_328,N_2942);
and U7227 (N_7227,N_1440,N_4528);
nand U7228 (N_7228,N_3421,N_3405);
or U7229 (N_7229,N_1926,N_2241);
nand U7230 (N_7230,N_523,N_3755);
or U7231 (N_7231,N_172,N_4943);
nor U7232 (N_7232,N_4765,N_2611);
and U7233 (N_7233,N_1153,N_4853);
nor U7234 (N_7234,N_2,N_834);
nand U7235 (N_7235,N_2967,N_1660);
nand U7236 (N_7236,N_2099,N_4441);
nand U7237 (N_7237,N_3441,N_230);
nor U7238 (N_7238,N_232,N_4442);
or U7239 (N_7239,N_1231,N_304);
nand U7240 (N_7240,N_4632,N_4718);
or U7241 (N_7241,N_453,N_4555);
nand U7242 (N_7242,N_4399,N_4574);
or U7243 (N_7243,N_5,N_242);
nor U7244 (N_7244,N_3456,N_2869);
or U7245 (N_7245,N_2542,N_3476);
and U7246 (N_7246,N_3697,N_1076);
or U7247 (N_7247,N_4065,N_2336);
and U7248 (N_7248,N_809,N_1745);
and U7249 (N_7249,N_2162,N_2972);
and U7250 (N_7250,N_164,N_1001);
and U7251 (N_7251,N_4250,N_4497);
and U7252 (N_7252,N_588,N_4915);
nand U7253 (N_7253,N_659,N_994);
nor U7254 (N_7254,N_1629,N_1374);
nor U7255 (N_7255,N_699,N_3646);
nor U7256 (N_7256,N_2720,N_3614);
nor U7257 (N_7257,N_2075,N_2369);
nor U7258 (N_7258,N_2156,N_3058);
nand U7259 (N_7259,N_1685,N_4849);
nor U7260 (N_7260,N_4964,N_3933);
nor U7261 (N_7261,N_162,N_16);
nand U7262 (N_7262,N_458,N_3145);
nand U7263 (N_7263,N_2697,N_4209);
nand U7264 (N_7264,N_4719,N_786);
nand U7265 (N_7265,N_1582,N_3309);
or U7266 (N_7266,N_4058,N_970);
nand U7267 (N_7267,N_850,N_4188);
or U7268 (N_7268,N_789,N_4972);
nor U7269 (N_7269,N_2572,N_3848);
nor U7270 (N_7270,N_1233,N_1897);
nand U7271 (N_7271,N_4818,N_1965);
nor U7272 (N_7272,N_3828,N_3178);
nor U7273 (N_7273,N_662,N_4672);
nand U7274 (N_7274,N_4978,N_148);
or U7275 (N_7275,N_899,N_387);
and U7276 (N_7276,N_3947,N_2262);
nor U7277 (N_7277,N_1159,N_3357);
nor U7278 (N_7278,N_3373,N_3001);
nand U7279 (N_7279,N_4821,N_2926);
nand U7280 (N_7280,N_2885,N_3426);
nand U7281 (N_7281,N_2402,N_736);
nor U7282 (N_7282,N_4003,N_1526);
nor U7283 (N_7283,N_2197,N_3384);
nand U7284 (N_7284,N_910,N_3496);
nor U7285 (N_7285,N_3530,N_772);
nor U7286 (N_7286,N_2298,N_2733);
nor U7287 (N_7287,N_4767,N_3584);
xnor U7288 (N_7288,N_1097,N_3264);
or U7289 (N_7289,N_4901,N_3761);
or U7290 (N_7290,N_2086,N_2470);
or U7291 (N_7291,N_3089,N_4304);
and U7292 (N_7292,N_3538,N_4111);
or U7293 (N_7293,N_2549,N_2124);
nand U7294 (N_7294,N_3689,N_4600);
or U7295 (N_7295,N_3970,N_2629);
and U7296 (N_7296,N_1196,N_555);
nor U7297 (N_7297,N_4423,N_4417);
or U7298 (N_7298,N_141,N_1162);
nand U7299 (N_7299,N_2675,N_3861);
nor U7300 (N_7300,N_3948,N_442);
or U7301 (N_7301,N_3074,N_233);
or U7302 (N_7302,N_3715,N_1438);
and U7303 (N_7303,N_3622,N_1003);
nand U7304 (N_7304,N_3594,N_19);
nand U7305 (N_7305,N_680,N_217);
or U7306 (N_7306,N_1376,N_575);
nand U7307 (N_7307,N_959,N_3206);
nand U7308 (N_7308,N_2420,N_2663);
or U7309 (N_7309,N_208,N_2750);
nand U7310 (N_7310,N_4677,N_3499);
and U7311 (N_7311,N_4706,N_4530);
nor U7312 (N_7312,N_593,N_31);
and U7313 (N_7313,N_2154,N_28);
or U7314 (N_7314,N_2499,N_2085);
nor U7315 (N_7315,N_3275,N_4048);
and U7316 (N_7316,N_1570,N_3433);
or U7317 (N_7317,N_791,N_1773);
nand U7318 (N_7318,N_4628,N_1179);
and U7319 (N_7319,N_3915,N_2626);
nand U7320 (N_7320,N_3181,N_3269);
and U7321 (N_7321,N_2139,N_4484);
and U7322 (N_7322,N_3492,N_1524);
nand U7323 (N_7323,N_2342,N_1284);
nand U7324 (N_7324,N_2786,N_4136);
or U7325 (N_7325,N_1074,N_229);
and U7326 (N_7326,N_3332,N_2405);
and U7327 (N_7327,N_4434,N_1940);
or U7328 (N_7328,N_71,N_4939);
nand U7329 (N_7329,N_2288,N_546);
nor U7330 (N_7330,N_615,N_3203);
or U7331 (N_7331,N_4687,N_2809);
and U7332 (N_7332,N_730,N_3610);
and U7333 (N_7333,N_4916,N_370);
or U7334 (N_7334,N_1010,N_4595);
nor U7335 (N_7335,N_2064,N_4648);
or U7336 (N_7336,N_4047,N_4725);
nor U7337 (N_7337,N_3406,N_1342);
nand U7338 (N_7338,N_2358,N_4749);
nand U7339 (N_7339,N_142,N_4355);
nor U7340 (N_7340,N_3599,N_339);
nand U7341 (N_7341,N_3866,N_4160);
or U7342 (N_7342,N_1006,N_3904);
or U7343 (N_7343,N_4320,N_4626);
or U7344 (N_7344,N_4635,N_432);
or U7345 (N_7345,N_3417,N_2093);
and U7346 (N_7346,N_954,N_4332);
and U7347 (N_7347,N_2916,N_4607);
and U7348 (N_7348,N_2797,N_3061);
and U7349 (N_7349,N_582,N_1998);
nor U7350 (N_7350,N_4278,N_3285);
and U7351 (N_7351,N_1007,N_3091);
and U7352 (N_7352,N_2908,N_1158);
and U7353 (N_7353,N_4653,N_3566);
and U7354 (N_7354,N_4660,N_2707);
nor U7355 (N_7355,N_497,N_2439);
and U7356 (N_7356,N_2444,N_289);
nor U7357 (N_7357,N_540,N_3353);
or U7358 (N_7358,N_500,N_4247);
or U7359 (N_7359,N_3712,N_4009);
and U7360 (N_7360,N_3624,N_2893);
nand U7361 (N_7361,N_4631,N_515);
or U7362 (N_7362,N_1226,N_2102);
nand U7363 (N_7363,N_2693,N_565);
and U7364 (N_7364,N_3049,N_3515);
nor U7365 (N_7365,N_3717,N_1527);
or U7366 (N_7366,N_1161,N_3090);
nor U7367 (N_7367,N_3812,N_3520);
nor U7368 (N_7368,N_17,N_613);
and U7369 (N_7369,N_1140,N_3085);
nor U7370 (N_7370,N_4351,N_1867);
or U7371 (N_7371,N_569,N_1997);
and U7372 (N_7372,N_629,N_3825);
nor U7373 (N_7373,N_1639,N_1086);
nor U7374 (N_7374,N_2178,N_149);
nand U7375 (N_7375,N_3927,N_1687);
nor U7376 (N_7376,N_2492,N_866);
nor U7377 (N_7377,N_1027,N_3900);
nor U7378 (N_7378,N_1512,N_3649);
nor U7379 (N_7379,N_2017,N_774);
nand U7380 (N_7380,N_1390,N_2438);
or U7381 (N_7381,N_564,N_3201);
nor U7382 (N_7382,N_1654,N_3171);
and U7383 (N_7383,N_655,N_473);
or U7384 (N_7384,N_2133,N_1633);
or U7385 (N_7385,N_4341,N_215);
and U7386 (N_7386,N_3451,N_2249);
nor U7387 (N_7387,N_159,N_4028);
and U7388 (N_7388,N_1689,N_1404);
nor U7389 (N_7389,N_3554,N_3509);
and U7390 (N_7390,N_123,N_3605);
nand U7391 (N_7391,N_2479,N_1925);
nor U7392 (N_7392,N_423,N_4919);
and U7393 (N_7393,N_936,N_1011);
or U7394 (N_7394,N_3220,N_2722);
nor U7395 (N_7395,N_859,N_678);
and U7396 (N_7396,N_3643,N_3749);
xnor U7397 (N_7397,N_3742,N_3728);
or U7398 (N_7398,N_4772,N_886);
nor U7399 (N_7399,N_3156,N_134);
and U7400 (N_7400,N_2796,N_352);
and U7401 (N_7401,N_4228,N_194);
or U7402 (N_7402,N_1345,N_3986);
and U7403 (N_7403,N_1990,N_3076);
or U7404 (N_7404,N_3674,N_300);
and U7405 (N_7405,N_400,N_3013);
or U7406 (N_7406,N_1769,N_4164);
nand U7407 (N_7407,N_3608,N_606);
nor U7408 (N_7408,N_4686,N_3244);
nor U7409 (N_7409,N_4156,N_3823);
and U7410 (N_7410,N_3621,N_4191);
xnor U7411 (N_7411,N_193,N_2482);
or U7412 (N_7412,N_2929,N_4099);
nand U7413 (N_7413,N_1590,N_3288);
or U7414 (N_7414,N_1172,N_1945);
nand U7415 (N_7415,N_4238,N_1485);
nand U7416 (N_7416,N_122,N_392);
xnor U7417 (N_7417,N_1827,N_44);
or U7418 (N_7418,N_2350,N_57);
and U7419 (N_7419,N_84,N_4840);
or U7420 (N_7420,N_1551,N_884);
xor U7421 (N_7421,N_2531,N_1338);
nand U7422 (N_7422,N_4234,N_2040);
nand U7423 (N_7423,N_155,N_307);
or U7424 (N_7424,N_1189,N_1220);
nand U7425 (N_7425,N_3073,N_2923);
and U7426 (N_7426,N_1500,N_450);
and U7427 (N_7427,N_4393,N_2351);
or U7428 (N_7428,N_2819,N_3418);
and U7429 (N_7429,N_2504,N_1327);
or U7430 (N_7430,N_1257,N_4352);
and U7431 (N_7431,N_3700,N_4624);
or U7432 (N_7432,N_993,N_2705);
or U7433 (N_7433,N_2503,N_4552);
or U7434 (N_7434,N_2577,N_766);
xnor U7435 (N_7435,N_4370,N_4039);
and U7436 (N_7436,N_2861,N_3258);
nor U7437 (N_7437,N_4889,N_144);
nor U7438 (N_7438,N_81,N_4482);
nor U7439 (N_7439,N_1,N_1822);
and U7440 (N_7440,N_3140,N_4949);
nand U7441 (N_7441,N_3756,N_409);
nor U7442 (N_7442,N_3095,N_2315);
or U7443 (N_7443,N_3601,N_3568);
and U7444 (N_7444,N_2982,N_3795);
nand U7445 (N_7445,N_2895,N_2734);
nand U7446 (N_7446,N_4911,N_4559);
or U7447 (N_7447,N_1771,N_1635);
nor U7448 (N_7448,N_2051,N_58);
nand U7449 (N_7449,N_2564,N_621);
nor U7450 (N_7450,N_1123,N_2595);
and U7451 (N_7451,N_2297,N_3497);
nor U7452 (N_7452,N_3615,N_163);
or U7453 (N_7453,N_3059,N_2273);
or U7454 (N_7454,N_2007,N_1734);
or U7455 (N_7455,N_4947,N_308);
and U7456 (N_7456,N_2948,N_4976);
and U7457 (N_7457,N_1922,N_2950);
and U7458 (N_7458,N_873,N_2827);
and U7459 (N_7459,N_1387,N_2848);
or U7460 (N_7460,N_2635,N_1810);
nor U7461 (N_7461,N_1416,N_1557);
and U7462 (N_7462,N_2447,N_4829);
nor U7463 (N_7463,N_2817,N_989);
nand U7464 (N_7464,N_2567,N_4556);
nor U7465 (N_7465,N_2615,N_3371);
nand U7466 (N_7466,N_1138,N_4276);
or U7467 (N_7467,N_1205,N_4926);
nand U7468 (N_7468,N_930,N_1835);
nor U7469 (N_7469,N_3890,N_4674);
nor U7470 (N_7470,N_3153,N_3879);
nor U7471 (N_7471,N_4193,N_2774);
and U7472 (N_7472,N_3490,N_4474);
or U7473 (N_7473,N_2063,N_628);
nor U7474 (N_7474,N_1025,N_2143);
nor U7475 (N_7475,N_3494,N_4757);
and U7476 (N_7476,N_234,N_2002);
nand U7477 (N_7477,N_1938,N_1562);
nor U7478 (N_7478,N_3071,N_396);
nor U7479 (N_7479,N_4440,N_2456);
nand U7480 (N_7480,N_1141,N_3652);
nand U7481 (N_7481,N_1829,N_890);
or U7482 (N_7482,N_1249,N_2054);
or U7483 (N_7483,N_4243,N_2548);
or U7484 (N_7484,N_2344,N_4023);
and U7485 (N_7485,N_2899,N_3653);
nor U7486 (N_7486,N_4933,N_2634);
nor U7487 (N_7487,N_2608,N_3767);
nand U7488 (N_7488,N_3951,N_971);
nand U7489 (N_7489,N_4382,N_469);
and U7490 (N_7490,N_4881,N_4097);
nand U7491 (N_7491,N_1854,N_4049);
nor U7492 (N_7492,N_4165,N_4035);
and U7493 (N_7493,N_1066,N_4834);
and U7494 (N_7494,N_1659,N_1267);
and U7495 (N_7495,N_346,N_4627);
or U7496 (N_7496,N_3251,N_3764);
nand U7497 (N_7497,N_530,N_2437);
or U7498 (N_7498,N_3086,N_2481);
nand U7499 (N_7499,N_3068,N_3077);
and U7500 (N_7500,N_4415,N_1114);
nor U7501 (N_7501,N_3013,N_1540);
nand U7502 (N_7502,N_1282,N_4191);
nor U7503 (N_7503,N_4081,N_1796);
nor U7504 (N_7504,N_1068,N_4262);
or U7505 (N_7505,N_627,N_4377);
nor U7506 (N_7506,N_4717,N_1558);
nor U7507 (N_7507,N_1968,N_3120);
nor U7508 (N_7508,N_3112,N_1117);
nor U7509 (N_7509,N_2551,N_3686);
or U7510 (N_7510,N_3543,N_1975);
nor U7511 (N_7511,N_983,N_2661);
and U7512 (N_7512,N_3543,N_3956);
nand U7513 (N_7513,N_4211,N_288);
nand U7514 (N_7514,N_3445,N_2098);
or U7515 (N_7515,N_2813,N_1170);
nand U7516 (N_7516,N_4246,N_4654);
nor U7517 (N_7517,N_4850,N_930);
xor U7518 (N_7518,N_1999,N_3784);
or U7519 (N_7519,N_1894,N_2857);
nand U7520 (N_7520,N_678,N_3760);
and U7521 (N_7521,N_4997,N_3638);
nand U7522 (N_7522,N_1149,N_1801);
nand U7523 (N_7523,N_513,N_1415);
nor U7524 (N_7524,N_1751,N_3420);
nand U7525 (N_7525,N_3267,N_3107);
and U7526 (N_7526,N_4895,N_1136);
or U7527 (N_7527,N_3742,N_1558);
and U7528 (N_7528,N_4822,N_4047);
or U7529 (N_7529,N_967,N_4560);
or U7530 (N_7530,N_3006,N_1368);
and U7531 (N_7531,N_3196,N_4228);
nor U7532 (N_7532,N_3000,N_3299);
and U7533 (N_7533,N_2108,N_3239);
nand U7534 (N_7534,N_83,N_2256);
and U7535 (N_7535,N_4998,N_705);
or U7536 (N_7536,N_3480,N_1780);
and U7537 (N_7537,N_1554,N_1466);
and U7538 (N_7538,N_1163,N_2353);
and U7539 (N_7539,N_4704,N_362);
or U7540 (N_7540,N_770,N_4603);
nand U7541 (N_7541,N_3961,N_2347);
or U7542 (N_7542,N_914,N_1557);
or U7543 (N_7543,N_3521,N_2640);
nor U7544 (N_7544,N_1374,N_2159);
nor U7545 (N_7545,N_4964,N_4967);
and U7546 (N_7546,N_2890,N_4358);
and U7547 (N_7547,N_2452,N_3867);
or U7548 (N_7548,N_4982,N_4878);
or U7549 (N_7549,N_1518,N_2186);
xor U7550 (N_7550,N_873,N_3864);
and U7551 (N_7551,N_4884,N_3647);
or U7552 (N_7552,N_3264,N_2566);
or U7553 (N_7553,N_1787,N_2305);
and U7554 (N_7554,N_2481,N_4504);
nand U7555 (N_7555,N_2557,N_441);
and U7556 (N_7556,N_4557,N_1273);
or U7557 (N_7557,N_2877,N_897);
or U7558 (N_7558,N_1327,N_2977);
and U7559 (N_7559,N_1333,N_1274);
and U7560 (N_7560,N_2456,N_296);
nor U7561 (N_7561,N_204,N_962);
and U7562 (N_7562,N_4217,N_4830);
and U7563 (N_7563,N_3570,N_1114);
nand U7564 (N_7564,N_2413,N_40);
and U7565 (N_7565,N_2252,N_818);
nor U7566 (N_7566,N_3427,N_2711);
nor U7567 (N_7567,N_2697,N_594);
and U7568 (N_7568,N_4894,N_4531);
nor U7569 (N_7569,N_2351,N_56);
and U7570 (N_7570,N_936,N_1595);
or U7571 (N_7571,N_2883,N_1429);
or U7572 (N_7572,N_3793,N_2673);
nand U7573 (N_7573,N_4020,N_4078);
nand U7574 (N_7574,N_4267,N_3524);
or U7575 (N_7575,N_3115,N_729);
nand U7576 (N_7576,N_3243,N_2545);
and U7577 (N_7577,N_1931,N_3693);
nand U7578 (N_7578,N_3484,N_540);
and U7579 (N_7579,N_4272,N_4104);
nand U7580 (N_7580,N_1145,N_2706);
nand U7581 (N_7581,N_4914,N_4500);
nand U7582 (N_7582,N_567,N_2705);
nor U7583 (N_7583,N_4173,N_3429);
nor U7584 (N_7584,N_2996,N_649);
and U7585 (N_7585,N_3603,N_3894);
and U7586 (N_7586,N_3287,N_1360);
and U7587 (N_7587,N_438,N_4396);
and U7588 (N_7588,N_1066,N_366);
nor U7589 (N_7589,N_522,N_372);
and U7590 (N_7590,N_3506,N_4062);
nand U7591 (N_7591,N_1692,N_1911);
xor U7592 (N_7592,N_3261,N_4886);
nor U7593 (N_7593,N_578,N_1575);
and U7594 (N_7594,N_1797,N_2713);
and U7595 (N_7595,N_4786,N_4620);
and U7596 (N_7596,N_2418,N_4152);
and U7597 (N_7597,N_1794,N_1066);
or U7598 (N_7598,N_3602,N_4953);
nand U7599 (N_7599,N_592,N_521);
and U7600 (N_7600,N_2915,N_4503);
nor U7601 (N_7601,N_4767,N_1050);
and U7602 (N_7602,N_3162,N_1918);
nor U7603 (N_7603,N_4243,N_380);
nand U7604 (N_7604,N_4262,N_1881);
and U7605 (N_7605,N_1189,N_1416);
nor U7606 (N_7606,N_2552,N_4054);
nand U7607 (N_7607,N_2473,N_2663);
nand U7608 (N_7608,N_3825,N_565);
nor U7609 (N_7609,N_3143,N_146);
nor U7610 (N_7610,N_886,N_4262);
or U7611 (N_7611,N_4074,N_2964);
nand U7612 (N_7612,N_4497,N_3537);
and U7613 (N_7613,N_4266,N_4354);
and U7614 (N_7614,N_4530,N_3966);
nor U7615 (N_7615,N_3453,N_4427);
nor U7616 (N_7616,N_3097,N_3763);
nor U7617 (N_7617,N_1804,N_3698);
nand U7618 (N_7618,N_2088,N_3609);
nand U7619 (N_7619,N_4100,N_4961);
nand U7620 (N_7620,N_1943,N_1930);
nor U7621 (N_7621,N_4089,N_2677);
nand U7622 (N_7622,N_419,N_4028);
or U7623 (N_7623,N_2048,N_2107);
nor U7624 (N_7624,N_2382,N_3317);
nor U7625 (N_7625,N_3490,N_2514);
nand U7626 (N_7626,N_3781,N_266);
and U7627 (N_7627,N_2022,N_383);
nor U7628 (N_7628,N_3212,N_1900);
or U7629 (N_7629,N_3191,N_28);
nor U7630 (N_7630,N_2134,N_1013);
or U7631 (N_7631,N_1264,N_2712);
nand U7632 (N_7632,N_4676,N_56);
nand U7633 (N_7633,N_4623,N_1563);
nor U7634 (N_7634,N_4554,N_3169);
or U7635 (N_7635,N_2421,N_4268);
nor U7636 (N_7636,N_4295,N_3843);
nand U7637 (N_7637,N_2337,N_1720);
or U7638 (N_7638,N_3076,N_1946);
nor U7639 (N_7639,N_2762,N_2513);
or U7640 (N_7640,N_910,N_3411);
and U7641 (N_7641,N_988,N_3454);
nor U7642 (N_7642,N_4714,N_4166);
nor U7643 (N_7643,N_909,N_3603);
and U7644 (N_7644,N_4996,N_2224);
or U7645 (N_7645,N_858,N_2935);
nor U7646 (N_7646,N_1167,N_3118);
or U7647 (N_7647,N_1001,N_2937);
and U7648 (N_7648,N_3619,N_4702);
and U7649 (N_7649,N_2533,N_3779);
nor U7650 (N_7650,N_2748,N_746);
or U7651 (N_7651,N_2413,N_2940);
nand U7652 (N_7652,N_4151,N_1890);
nor U7653 (N_7653,N_1825,N_343);
nand U7654 (N_7654,N_324,N_1278);
nor U7655 (N_7655,N_3926,N_427);
or U7656 (N_7656,N_1841,N_2792);
and U7657 (N_7657,N_4858,N_3529);
or U7658 (N_7658,N_306,N_1928);
and U7659 (N_7659,N_298,N_1304);
or U7660 (N_7660,N_411,N_84);
or U7661 (N_7661,N_4062,N_4441);
nand U7662 (N_7662,N_1292,N_205);
and U7663 (N_7663,N_550,N_4615);
nor U7664 (N_7664,N_3490,N_2954);
and U7665 (N_7665,N_2153,N_2004);
nor U7666 (N_7666,N_1851,N_4256);
nor U7667 (N_7667,N_3772,N_3362);
nand U7668 (N_7668,N_1611,N_943);
nor U7669 (N_7669,N_929,N_3948);
nand U7670 (N_7670,N_1650,N_1839);
nand U7671 (N_7671,N_1947,N_2204);
or U7672 (N_7672,N_4325,N_3337);
and U7673 (N_7673,N_1245,N_3087);
or U7674 (N_7674,N_469,N_3139);
nor U7675 (N_7675,N_3704,N_3291);
and U7676 (N_7676,N_2430,N_3300);
nor U7677 (N_7677,N_371,N_3991);
or U7678 (N_7678,N_4996,N_435);
nand U7679 (N_7679,N_821,N_1286);
and U7680 (N_7680,N_224,N_1215);
nor U7681 (N_7681,N_444,N_4949);
nand U7682 (N_7682,N_4292,N_3401);
nor U7683 (N_7683,N_3151,N_3824);
or U7684 (N_7684,N_808,N_804);
or U7685 (N_7685,N_4481,N_4691);
nor U7686 (N_7686,N_2242,N_2673);
or U7687 (N_7687,N_2724,N_4451);
and U7688 (N_7688,N_4398,N_3177);
nor U7689 (N_7689,N_1954,N_1663);
nand U7690 (N_7690,N_4513,N_4433);
and U7691 (N_7691,N_3643,N_2850);
nand U7692 (N_7692,N_2419,N_2354);
xnor U7693 (N_7693,N_426,N_265);
nor U7694 (N_7694,N_1927,N_2139);
and U7695 (N_7695,N_4487,N_597);
nand U7696 (N_7696,N_2642,N_1544);
nor U7697 (N_7697,N_3479,N_1294);
or U7698 (N_7698,N_3676,N_495);
or U7699 (N_7699,N_766,N_1473);
or U7700 (N_7700,N_2492,N_3779);
nand U7701 (N_7701,N_4791,N_1581);
nor U7702 (N_7702,N_642,N_3702);
nor U7703 (N_7703,N_3720,N_2677);
nor U7704 (N_7704,N_2148,N_821);
nor U7705 (N_7705,N_1371,N_3781);
nand U7706 (N_7706,N_3530,N_2367);
nand U7707 (N_7707,N_14,N_702);
nand U7708 (N_7708,N_4280,N_785);
nand U7709 (N_7709,N_1918,N_378);
or U7710 (N_7710,N_499,N_4271);
or U7711 (N_7711,N_4538,N_1987);
and U7712 (N_7712,N_2186,N_713);
and U7713 (N_7713,N_2459,N_4284);
nand U7714 (N_7714,N_4252,N_679);
nand U7715 (N_7715,N_4350,N_2725);
nor U7716 (N_7716,N_4098,N_1909);
nor U7717 (N_7717,N_779,N_2524);
and U7718 (N_7718,N_4183,N_3827);
nor U7719 (N_7719,N_4652,N_677);
and U7720 (N_7720,N_1878,N_3811);
or U7721 (N_7721,N_1638,N_1534);
nor U7722 (N_7722,N_3131,N_1795);
or U7723 (N_7723,N_3459,N_2680);
nor U7724 (N_7724,N_2727,N_1417);
nand U7725 (N_7725,N_2383,N_2846);
and U7726 (N_7726,N_1527,N_2322);
nor U7727 (N_7727,N_606,N_2641);
or U7728 (N_7728,N_2674,N_147);
nand U7729 (N_7729,N_1421,N_172);
nor U7730 (N_7730,N_60,N_873);
and U7731 (N_7731,N_1216,N_2349);
nand U7732 (N_7732,N_3967,N_3164);
nor U7733 (N_7733,N_4533,N_815);
or U7734 (N_7734,N_4887,N_3139);
and U7735 (N_7735,N_1504,N_2713);
and U7736 (N_7736,N_4768,N_2201);
nand U7737 (N_7737,N_4435,N_2251);
and U7738 (N_7738,N_4723,N_1792);
and U7739 (N_7739,N_4443,N_1632);
and U7740 (N_7740,N_176,N_2033);
nor U7741 (N_7741,N_3787,N_1483);
nand U7742 (N_7742,N_4665,N_3467);
nor U7743 (N_7743,N_3445,N_755);
nand U7744 (N_7744,N_4856,N_214);
and U7745 (N_7745,N_3862,N_779);
and U7746 (N_7746,N_2760,N_3379);
nor U7747 (N_7747,N_3032,N_1776);
and U7748 (N_7748,N_3116,N_2968);
or U7749 (N_7749,N_792,N_3915);
nor U7750 (N_7750,N_1797,N_4380);
or U7751 (N_7751,N_1144,N_4651);
nor U7752 (N_7752,N_3843,N_4720);
or U7753 (N_7753,N_1541,N_3609);
nand U7754 (N_7754,N_4308,N_2520);
nor U7755 (N_7755,N_3113,N_2856);
or U7756 (N_7756,N_932,N_1471);
nand U7757 (N_7757,N_414,N_1272);
nor U7758 (N_7758,N_2085,N_1558);
and U7759 (N_7759,N_699,N_1393);
and U7760 (N_7760,N_252,N_1843);
or U7761 (N_7761,N_111,N_2566);
or U7762 (N_7762,N_4131,N_3500);
and U7763 (N_7763,N_1576,N_96);
and U7764 (N_7764,N_2389,N_3191);
or U7765 (N_7765,N_2044,N_3464);
or U7766 (N_7766,N_3158,N_3346);
and U7767 (N_7767,N_3578,N_2443);
nor U7768 (N_7768,N_2974,N_154);
nand U7769 (N_7769,N_3456,N_2052);
or U7770 (N_7770,N_283,N_4636);
or U7771 (N_7771,N_1579,N_879);
nor U7772 (N_7772,N_4583,N_4732);
or U7773 (N_7773,N_4198,N_3686);
and U7774 (N_7774,N_3246,N_790);
and U7775 (N_7775,N_1899,N_3260);
or U7776 (N_7776,N_4891,N_3526);
or U7777 (N_7777,N_1990,N_1188);
or U7778 (N_7778,N_4682,N_2148);
and U7779 (N_7779,N_3166,N_4783);
and U7780 (N_7780,N_3348,N_4962);
or U7781 (N_7781,N_4153,N_2873);
or U7782 (N_7782,N_2595,N_1515);
nand U7783 (N_7783,N_4474,N_1014);
or U7784 (N_7784,N_3925,N_4297);
nor U7785 (N_7785,N_4527,N_3029);
and U7786 (N_7786,N_592,N_2351);
or U7787 (N_7787,N_1145,N_1625);
or U7788 (N_7788,N_4856,N_4071);
nand U7789 (N_7789,N_4402,N_2800);
nor U7790 (N_7790,N_1692,N_981);
nand U7791 (N_7791,N_1317,N_3385);
nand U7792 (N_7792,N_132,N_265);
or U7793 (N_7793,N_4634,N_2852);
and U7794 (N_7794,N_3886,N_3823);
nor U7795 (N_7795,N_3027,N_4396);
and U7796 (N_7796,N_2567,N_741);
nor U7797 (N_7797,N_1645,N_1738);
or U7798 (N_7798,N_1703,N_2355);
nor U7799 (N_7799,N_832,N_1754);
nand U7800 (N_7800,N_2864,N_2669);
or U7801 (N_7801,N_154,N_933);
or U7802 (N_7802,N_2335,N_338);
xnor U7803 (N_7803,N_1655,N_3193);
nand U7804 (N_7804,N_1106,N_4120);
nand U7805 (N_7805,N_3100,N_3428);
and U7806 (N_7806,N_2540,N_1087);
and U7807 (N_7807,N_1244,N_2526);
nor U7808 (N_7808,N_571,N_3823);
nand U7809 (N_7809,N_3527,N_666);
nand U7810 (N_7810,N_883,N_1077);
nand U7811 (N_7811,N_300,N_4241);
nand U7812 (N_7812,N_4101,N_224);
nand U7813 (N_7813,N_3847,N_3845);
nand U7814 (N_7814,N_301,N_4090);
or U7815 (N_7815,N_3554,N_4016);
nor U7816 (N_7816,N_2559,N_3859);
and U7817 (N_7817,N_4244,N_3140);
nor U7818 (N_7818,N_3724,N_2923);
or U7819 (N_7819,N_3222,N_1159);
or U7820 (N_7820,N_1462,N_3230);
and U7821 (N_7821,N_2612,N_4768);
nor U7822 (N_7822,N_1531,N_888);
nor U7823 (N_7823,N_921,N_2382);
or U7824 (N_7824,N_4489,N_1624);
nand U7825 (N_7825,N_1425,N_821);
or U7826 (N_7826,N_1290,N_1110);
or U7827 (N_7827,N_1833,N_2290);
and U7828 (N_7828,N_1158,N_2453);
or U7829 (N_7829,N_4557,N_3107);
or U7830 (N_7830,N_1568,N_4113);
nand U7831 (N_7831,N_1378,N_3565);
nor U7832 (N_7832,N_3660,N_1337);
or U7833 (N_7833,N_1530,N_4017);
nand U7834 (N_7834,N_1485,N_3770);
and U7835 (N_7835,N_336,N_416);
and U7836 (N_7836,N_2015,N_3397);
and U7837 (N_7837,N_328,N_1196);
nor U7838 (N_7838,N_444,N_3830);
or U7839 (N_7839,N_4726,N_2475);
nand U7840 (N_7840,N_332,N_3044);
or U7841 (N_7841,N_3127,N_3641);
and U7842 (N_7842,N_1352,N_2840);
nor U7843 (N_7843,N_2165,N_2405);
and U7844 (N_7844,N_1662,N_2491);
nor U7845 (N_7845,N_2659,N_4016);
or U7846 (N_7846,N_2361,N_2081);
or U7847 (N_7847,N_2902,N_1150);
nand U7848 (N_7848,N_4233,N_2410);
nor U7849 (N_7849,N_3122,N_1886);
and U7850 (N_7850,N_4947,N_4642);
or U7851 (N_7851,N_3705,N_3481);
nor U7852 (N_7852,N_1892,N_1712);
nand U7853 (N_7853,N_1657,N_413);
and U7854 (N_7854,N_3370,N_97);
and U7855 (N_7855,N_4359,N_4209);
xnor U7856 (N_7856,N_1286,N_3456);
and U7857 (N_7857,N_2772,N_2917);
nor U7858 (N_7858,N_475,N_317);
and U7859 (N_7859,N_4661,N_3643);
nor U7860 (N_7860,N_191,N_3570);
nand U7861 (N_7861,N_4172,N_107);
or U7862 (N_7862,N_3745,N_3419);
and U7863 (N_7863,N_1844,N_433);
nand U7864 (N_7864,N_769,N_617);
nor U7865 (N_7865,N_4649,N_4651);
or U7866 (N_7866,N_4794,N_3588);
and U7867 (N_7867,N_810,N_3166);
or U7868 (N_7868,N_1077,N_2625);
or U7869 (N_7869,N_3048,N_2918);
and U7870 (N_7870,N_2231,N_1816);
or U7871 (N_7871,N_4116,N_2765);
or U7872 (N_7872,N_6,N_299);
and U7873 (N_7873,N_4727,N_2661);
or U7874 (N_7874,N_1094,N_1796);
nand U7875 (N_7875,N_1259,N_3594);
and U7876 (N_7876,N_2112,N_1675);
nand U7877 (N_7877,N_4571,N_200);
or U7878 (N_7878,N_3097,N_2271);
and U7879 (N_7879,N_531,N_730);
nor U7880 (N_7880,N_4740,N_494);
xor U7881 (N_7881,N_873,N_2946);
nor U7882 (N_7882,N_67,N_4218);
nand U7883 (N_7883,N_4909,N_2562);
nand U7884 (N_7884,N_4029,N_2923);
nor U7885 (N_7885,N_3641,N_156);
and U7886 (N_7886,N_3809,N_2638);
and U7887 (N_7887,N_1260,N_3523);
or U7888 (N_7888,N_2181,N_960);
nor U7889 (N_7889,N_236,N_1442);
or U7890 (N_7890,N_3187,N_2578);
nor U7891 (N_7891,N_2913,N_3471);
nor U7892 (N_7892,N_3746,N_4450);
and U7893 (N_7893,N_1628,N_1916);
and U7894 (N_7894,N_1645,N_2864);
and U7895 (N_7895,N_92,N_1536);
or U7896 (N_7896,N_680,N_4074);
nand U7897 (N_7897,N_2468,N_1655);
nand U7898 (N_7898,N_4081,N_1221);
or U7899 (N_7899,N_672,N_2737);
nand U7900 (N_7900,N_276,N_1403);
or U7901 (N_7901,N_2855,N_330);
nor U7902 (N_7902,N_1944,N_3664);
nand U7903 (N_7903,N_3912,N_3057);
or U7904 (N_7904,N_3042,N_228);
nand U7905 (N_7905,N_4199,N_2403);
nand U7906 (N_7906,N_4787,N_1244);
or U7907 (N_7907,N_1137,N_4921);
or U7908 (N_7908,N_1220,N_2110);
or U7909 (N_7909,N_3774,N_3184);
or U7910 (N_7910,N_1272,N_1910);
or U7911 (N_7911,N_1798,N_377);
nor U7912 (N_7912,N_476,N_4720);
and U7913 (N_7913,N_1126,N_4917);
and U7914 (N_7914,N_1764,N_1755);
nor U7915 (N_7915,N_4299,N_1104);
nor U7916 (N_7916,N_1828,N_695);
nor U7917 (N_7917,N_2211,N_2879);
nand U7918 (N_7918,N_1622,N_4842);
or U7919 (N_7919,N_4280,N_2867);
nor U7920 (N_7920,N_5,N_2994);
or U7921 (N_7921,N_3878,N_3020);
and U7922 (N_7922,N_364,N_4072);
nand U7923 (N_7923,N_2399,N_2697);
nand U7924 (N_7924,N_3234,N_963);
or U7925 (N_7925,N_4284,N_3426);
nand U7926 (N_7926,N_2591,N_3222);
and U7927 (N_7927,N_3446,N_993);
nor U7928 (N_7928,N_4620,N_748);
or U7929 (N_7929,N_4834,N_1738);
and U7930 (N_7930,N_3218,N_2604);
nand U7931 (N_7931,N_867,N_4105);
and U7932 (N_7932,N_3377,N_51);
nor U7933 (N_7933,N_387,N_2875);
and U7934 (N_7934,N_3834,N_2139);
or U7935 (N_7935,N_3849,N_2794);
nor U7936 (N_7936,N_510,N_1456);
or U7937 (N_7937,N_1048,N_2607);
and U7938 (N_7938,N_3414,N_3005);
and U7939 (N_7939,N_3900,N_2593);
nand U7940 (N_7940,N_1989,N_4903);
or U7941 (N_7941,N_373,N_2694);
nor U7942 (N_7942,N_1207,N_2920);
or U7943 (N_7943,N_2065,N_3866);
and U7944 (N_7944,N_3909,N_2857);
nor U7945 (N_7945,N_964,N_900);
and U7946 (N_7946,N_325,N_4702);
or U7947 (N_7947,N_1892,N_4407);
or U7948 (N_7948,N_779,N_2854);
or U7949 (N_7949,N_3288,N_1622);
or U7950 (N_7950,N_3288,N_609);
and U7951 (N_7951,N_1670,N_2429);
and U7952 (N_7952,N_4878,N_3895);
or U7953 (N_7953,N_347,N_2926);
or U7954 (N_7954,N_1288,N_915);
or U7955 (N_7955,N_4561,N_798);
or U7956 (N_7956,N_3544,N_4263);
or U7957 (N_7957,N_3105,N_4565);
nand U7958 (N_7958,N_2433,N_2695);
and U7959 (N_7959,N_4720,N_430);
nor U7960 (N_7960,N_1234,N_2353);
or U7961 (N_7961,N_1366,N_1383);
nand U7962 (N_7962,N_846,N_3791);
and U7963 (N_7963,N_2945,N_4251);
or U7964 (N_7964,N_978,N_1246);
nand U7965 (N_7965,N_4589,N_1993);
nor U7966 (N_7966,N_1824,N_2757);
nand U7967 (N_7967,N_2390,N_4623);
nor U7968 (N_7968,N_4221,N_3146);
nor U7969 (N_7969,N_1964,N_4665);
or U7970 (N_7970,N_1110,N_2976);
nand U7971 (N_7971,N_4009,N_292);
nor U7972 (N_7972,N_3623,N_4804);
nor U7973 (N_7973,N_1680,N_984);
nor U7974 (N_7974,N_1398,N_531);
or U7975 (N_7975,N_1180,N_1468);
nand U7976 (N_7976,N_3704,N_361);
and U7977 (N_7977,N_138,N_12);
or U7978 (N_7978,N_2485,N_774);
and U7979 (N_7979,N_4727,N_3902);
or U7980 (N_7980,N_4707,N_4280);
nor U7981 (N_7981,N_2581,N_4756);
and U7982 (N_7982,N_3022,N_909);
or U7983 (N_7983,N_2314,N_3789);
and U7984 (N_7984,N_2857,N_1581);
nand U7985 (N_7985,N_1122,N_2092);
nand U7986 (N_7986,N_2221,N_4307);
or U7987 (N_7987,N_3524,N_3462);
or U7988 (N_7988,N_603,N_30);
nand U7989 (N_7989,N_79,N_1946);
and U7990 (N_7990,N_4220,N_2907);
nand U7991 (N_7991,N_3701,N_1169);
nand U7992 (N_7992,N_1394,N_4841);
or U7993 (N_7993,N_310,N_2896);
nand U7994 (N_7994,N_4661,N_3145);
nand U7995 (N_7995,N_1143,N_4289);
nor U7996 (N_7996,N_142,N_1879);
or U7997 (N_7997,N_3584,N_1374);
nand U7998 (N_7998,N_2249,N_963);
and U7999 (N_7999,N_125,N_3099);
nand U8000 (N_8000,N_517,N_2805);
nand U8001 (N_8001,N_3884,N_4944);
nor U8002 (N_8002,N_3244,N_1586);
or U8003 (N_8003,N_3869,N_2516);
or U8004 (N_8004,N_357,N_2350);
and U8005 (N_8005,N_3764,N_3731);
and U8006 (N_8006,N_4673,N_67);
nand U8007 (N_8007,N_2108,N_277);
nand U8008 (N_8008,N_3496,N_3270);
nand U8009 (N_8009,N_4697,N_912);
nor U8010 (N_8010,N_4645,N_4463);
nand U8011 (N_8011,N_2468,N_3063);
nor U8012 (N_8012,N_4907,N_324);
nand U8013 (N_8013,N_753,N_3400);
nand U8014 (N_8014,N_4264,N_3892);
and U8015 (N_8015,N_1425,N_1777);
nor U8016 (N_8016,N_2289,N_3885);
nand U8017 (N_8017,N_2456,N_3922);
and U8018 (N_8018,N_1198,N_1953);
and U8019 (N_8019,N_3103,N_4657);
and U8020 (N_8020,N_1039,N_282);
and U8021 (N_8021,N_2755,N_664);
nand U8022 (N_8022,N_94,N_3556);
nor U8023 (N_8023,N_89,N_4937);
nand U8024 (N_8024,N_1714,N_803);
and U8025 (N_8025,N_3350,N_3113);
or U8026 (N_8026,N_81,N_4841);
and U8027 (N_8027,N_864,N_127);
nand U8028 (N_8028,N_3689,N_3385);
and U8029 (N_8029,N_3191,N_1880);
nor U8030 (N_8030,N_3751,N_707);
nand U8031 (N_8031,N_602,N_66);
nand U8032 (N_8032,N_418,N_4348);
or U8033 (N_8033,N_1926,N_4663);
or U8034 (N_8034,N_707,N_4697);
nand U8035 (N_8035,N_1069,N_2452);
and U8036 (N_8036,N_4647,N_4316);
nor U8037 (N_8037,N_3827,N_4428);
or U8038 (N_8038,N_2065,N_4346);
or U8039 (N_8039,N_3170,N_1381);
or U8040 (N_8040,N_426,N_3507);
or U8041 (N_8041,N_756,N_2223);
nor U8042 (N_8042,N_4975,N_227);
nor U8043 (N_8043,N_4649,N_536);
or U8044 (N_8044,N_809,N_1601);
nand U8045 (N_8045,N_4645,N_1072);
and U8046 (N_8046,N_1124,N_1964);
nand U8047 (N_8047,N_4698,N_4156);
nand U8048 (N_8048,N_2241,N_4354);
and U8049 (N_8049,N_3856,N_4007);
or U8050 (N_8050,N_1329,N_2923);
nor U8051 (N_8051,N_715,N_4945);
and U8052 (N_8052,N_3639,N_3032);
and U8053 (N_8053,N_3851,N_4827);
nand U8054 (N_8054,N_2966,N_1492);
nand U8055 (N_8055,N_2468,N_4150);
nand U8056 (N_8056,N_4640,N_4459);
nand U8057 (N_8057,N_934,N_2781);
or U8058 (N_8058,N_3893,N_1817);
nand U8059 (N_8059,N_597,N_1516);
nor U8060 (N_8060,N_3060,N_1303);
and U8061 (N_8061,N_1874,N_172);
nor U8062 (N_8062,N_818,N_1641);
nor U8063 (N_8063,N_1318,N_2709);
or U8064 (N_8064,N_2241,N_2640);
nor U8065 (N_8065,N_4574,N_1453);
nand U8066 (N_8066,N_3856,N_4952);
nand U8067 (N_8067,N_1887,N_1591);
or U8068 (N_8068,N_660,N_2732);
nor U8069 (N_8069,N_293,N_4719);
nor U8070 (N_8070,N_4302,N_3085);
or U8071 (N_8071,N_2775,N_2680);
or U8072 (N_8072,N_1884,N_4998);
nand U8073 (N_8073,N_1234,N_594);
and U8074 (N_8074,N_4000,N_3606);
nand U8075 (N_8075,N_3743,N_3637);
nand U8076 (N_8076,N_172,N_708);
nor U8077 (N_8077,N_3689,N_3223);
or U8078 (N_8078,N_3730,N_2737);
and U8079 (N_8079,N_4624,N_150);
nor U8080 (N_8080,N_477,N_569);
or U8081 (N_8081,N_4750,N_314);
nand U8082 (N_8082,N_4303,N_2095);
nand U8083 (N_8083,N_2184,N_3970);
nand U8084 (N_8084,N_4797,N_3728);
nor U8085 (N_8085,N_1243,N_3432);
and U8086 (N_8086,N_3676,N_3071);
nand U8087 (N_8087,N_1386,N_3346);
and U8088 (N_8088,N_3455,N_3740);
and U8089 (N_8089,N_2073,N_4202);
or U8090 (N_8090,N_414,N_81);
nand U8091 (N_8091,N_2490,N_2771);
or U8092 (N_8092,N_2919,N_2491);
and U8093 (N_8093,N_4238,N_2507);
nand U8094 (N_8094,N_4542,N_900);
or U8095 (N_8095,N_2863,N_1655);
nor U8096 (N_8096,N_4004,N_840);
nand U8097 (N_8097,N_1530,N_3065);
nor U8098 (N_8098,N_1924,N_188);
or U8099 (N_8099,N_4769,N_3693);
nor U8100 (N_8100,N_1721,N_1413);
or U8101 (N_8101,N_2556,N_1283);
nor U8102 (N_8102,N_936,N_2362);
and U8103 (N_8103,N_411,N_2809);
nand U8104 (N_8104,N_4867,N_3328);
and U8105 (N_8105,N_3105,N_3772);
or U8106 (N_8106,N_263,N_842);
or U8107 (N_8107,N_2452,N_2867);
nor U8108 (N_8108,N_575,N_4910);
or U8109 (N_8109,N_1625,N_3482);
or U8110 (N_8110,N_3797,N_523);
or U8111 (N_8111,N_4173,N_193);
nand U8112 (N_8112,N_3268,N_2546);
nor U8113 (N_8113,N_3218,N_1851);
and U8114 (N_8114,N_1423,N_483);
or U8115 (N_8115,N_3961,N_2988);
nor U8116 (N_8116,N_1443,N_2029);
nand U8117 (N_8117,N_911,N_1071);
or U8118 (N_8118,N_2363,N_2997);
and U8119 (N_8119,N_4061,N_4218);
nand U8120 (N_8120,N_4511,N_3608);
nand U8121 (N_8121,N_4064,N_3362);
nor U8122 (N_8122,N_3181,N_82);
and U8123 (N_8123,N_2959,N_1562);
and U8124 (N_8124,N_871,N_3037);
nand U8125 (N_8125,N_4880,N_1213);
nor U8126 (N_8126,N_3446,N_437);
or U8127 (N_8127,N_4566,N_1320);
or U8128 (N_8128,N_3944,N_3128);
nand U8129 (N_8129,N_1723,N_3450);
and U8130 (N_8130,N_4677,N_243);
nand U8131 (N_8131,N_3763,N_817);
and U8132 (N_8132,N_228,N_4363);
or U8133 (N_8133,N_1579,N_953);
nand U8134 (N_8134,N_3849,N_3698);
or U8135 (N_8135,N_3318,N_4837);
nor U8136 (N_8136,N_4014,N_1492);
or U8137 (N_8137,N_3101,N_302);
nand U8138 (N_8138,N_2336,N_4929);
nand U8139 (N_8139,N_489,N_1878);
or U8140 (N_8140,N_934,N_2229);
and U8141 (N_8141,N_2190,N_1598);
nand U8142 (N_8142,N_2290,N_4865);
and U8143 (N_8143,N_4060,N_1995);
nor U8144 (N_8144,N_3905,N_306);
and U8145 (N_8145,N_1794,N_1434);
and U8146 (N_8146,N_537,N_2222);
nor U8147 (N_8147,N_985,N_847);
nand U8148 (N_8148,N_3561,N_2288);
nand U8149 (N_8149,N_3708,N_1456);
nor U8150 (N_8150,N_1497,N_3740);
or U8151 (N_8151,N_128,N_4676);
nand U8152 (N_8152,N_86,N_4546);
nor U8153 (N_8153,N_2210,N_2163);
nor U8154 (N_8154,N_4011,N_3576);
and U8155 (N_8155,N_823,N_1144);
or U8156 (N_8156,N_940,N_4320);
nand U8157 (N_8157,N_1592,N_789);
or U8158 (N_8158,N_4646,N_3920);
or U8159 (N_8159,N_1243,N_2072);
nand U8160 (N_8160,N_3770,N_4006);
nor U8161 (N_8161,N_315,N_357);
nand U8162 (N_8162,N_1219,N_194);
nand U8163 (N_8163,N_4748,N_182);
or U8164 (N_8164,N_3738,N_998);
and U8165 (N_8165,N_3433,N_72);
or U8166 (N_8166,N_854,N_127);
and U8167 (N_8167,N_3537,N_1257);
nor U8168 (N_8168,N_3646,N_3537);
nor U8169 (N_8169,N_2991,N_1774);
nor U8170 (N_8170,N_290,N_2568);
and U8171 (N_8171,N_4485,N_2967);
nor U8172 (N_8172,N_1174,N_4156);
and U8173 (N_8173,N_4914,N_1708);
and U8174 (N_8174,N_2620,N_2026);
and U8175 (N_8175,N_1885,N_4266);
nand U8176 (N_8176,N_4559,N_1994);
nor U8177 (N_8177,N_2112,N_2065);
or U8178 (N_8178,N_1371,N_682);
and U8179 (N_8179,N_4899,N_1251);
nor U8180 (N_8180,N_4428,N_3202);
nor U8181 (N_8181,N_2565,N_767);
and U8182 (N_8182,N_193,N_4064);
or U8183 (N_8183,N_362,N_4804);
or U8184 (N_8184,N_2961,N_399);
or U8185 (N_8185,N_4579,N_2799);
nor U8186 (N_8186,N_2582,N_888);
nand U8187 (N_8187,N_3931,N_4287);
or U8188 (N_8188,N_3446,N_2871);
nand U8189 (N_8189,N_2824,N_744);
and U8190 (N_8190,N_4479,N_4802);
and U8191 (N_8191,N_1957,N_2239);
or U8192 (N_8192,N_3672,N_4347);
and U8193 (N_8193,N_9,N_2985);
nand U8194 (N_8194,N_3962,N_3445);
nand U8195 (N_8195,N_3231,N_2062);
nor U8196 (N_8196,N_3891,N_1684);
nand U8197 (N_8197,N_3200,N_4422);
nor U8198 (N_8198,N_4078,N_181);
or U8199 (N_8199,N_2936,N_1115);
nand U8200 (N_8200,N_2755,N_450);
nand U8201 (N_8201,N_3355,N_4387);
nor U8202 (N_8202,N_4531,N_2594);
and U8203 (N_8203,N_4324,N_452);
and U8204 (N_8204,N_335,N_4936);
or U8205 (N_8205,N_1512,N_3977);
or U8206 (N_8206,N_2917,N_3720);
nand U8207 (N_8207,N_4018,N_3002);
and U8208 (N_8208,N_4945,N_2510);
nand U8209 (N_8209,N_3802,N_4844);
nor U8210 (N_8210,N_893,N_826);
or U8211 (N_8211,N_2973,N_638);
or U8212 (N_8212,N_2498,N_3137);
and U8213 (N_8213,N_1670,N_4372);
and U8214 (N_8214,N_3993,N_4000);
nor U8215 (N_8215,N_2400,N_902);
nand U8216 (N_8216,N_355,N_1064);
or U8217 (N_8217,N_2831,N_1004);
nor U8218 (N_8218,N_1551,N_3634);
nor U8219 (N_8219,N_1839,N_925);
and U8220 (N_8220,N_3092,N_2992);
nor U8221 (N_8221,N_319,N_3847);
or U8222 (N_8222,N_3610,N_968);
or U8223 (N_8223,N_4087,N_4768);
nor U8224 (N_8224,N_4453,N_1244);
nand U8225 (N_8225,N_4837,N_724);
nand U8226 (N_8226,N_2431,N_4012);
and U8227 (N_8227,N_1932,N_1528);
or U8228 (N_8228,N_3738,N_3766);
nor U8229 (N_8229,N_538,N_2575);
and U8230 (N_8230,N_469,N_2757);
or U8231 (N_8231,N_4818,N_1544);
nor U8232 (N_8232,N_1769,N_1752);
nor U8233 (N_8233,N_1550,N_3610);
nand U8234 (N_8234,N_3121,N_1639);
nor U8235 (N_8235,N_3416,N_4130);
xnor U8236 (N_8236,N_3080,N_1265);
or U8237 (N_8237,N_2904,N_4753);
and U8238 (N_8238,N_569,N_3037);
and U8239 (N_8239,N_1932,N_275);
nand U8240 (N_8240,N_2071,N_2636);
and U8241 (N_8241,N_3194,N_3079);
nor U8242 (N_8242,N_1955,N_1390);
and U8243 (N_8243,N_817,N_2652);
and U8244 (N_8244,N_4804,N_4943);
and U8245 (N_8245,N_3058,N_4942);
or U8246 (N_8246,N_1466,N_1630);
nand U8247 (N_8247,N_3038,N_2439);
nand U8248 (N_8248,N_2061,N_3572);
or U8249 (N_8249,N_4945,N_1486);
nor U8250 (N_8250,N_4930,N_2682);
or U8251 (N_8251,N_4357,N_1548);
nand U8252 (N_8252,N_1720,N_1229);
nand U8253 (N_8253,N_1805,N_2186);
nor U8254 (N_8254,N_3462,N_3909);
nand U8255 (N_8255,N_749,N_936);
or U8256 (N_8256,N_3792,N_2630);
nor U8257 (N_8257,N_2321,N_2625);
and U8258 (N_8258,N_3740,N_4321);
nand U8259 (N_8259,N_1751,N_3155);
nor U8260 (N_8260,N_2261,N_849);
or U8261 (N_8261,N_3119,N_1478);
nor U8262 (N_8262,N_1934,N_3347);
nor U8263 (N_8263,N_524,N_1899);
nand U8264 (N_8264,N_3659,N_3128);
nand U8265 (N_8265,N_2150,N_2994);
nand U8266 (N_8266,N_2789,N_525);
nand U8267 (N_8267,N_2947,N_2436);
and U8268 (N_8268,N_2013,N_970);
nor U8269 (N_8269,N_2643,N_1005);
or U8270 (N_8270,N_2002,N_2121);
and U8271 (N_8271,N_3597,N_1827);
nand U8272 (N_8272,N_2080,N_4443);
nand U8273 (N_8273,N_2827,N_3820);
nor U8274 (N_8274,N_1251,N_207);
or U8275 (N_8275,N_2838,N_2394);
and U8276 (N_8276,N_1351,N_4020);
or U8277 (N_8277,N_2013,N_4168);
or U8278 (N_8278,N_4153,N_4137);
and U8279 (N_8279,N_895,N_2201);
and U8280 (N_8280,N_2351,N_2462);
and U8281 (N_8281,N_4453,N_2402);
nand U8282 (N_8282,N_724,N_2565);
or U8283 (N_8283,N_757,N_3395);
and U8284 (N_8284,N_2760,N_529);
nor U8285 (N_8285,N_4626,N_2853);
nor U8286 (N_8286,N_2397,N_2567);
and U8287 (N_8287,N_3226,N_786);
nand U8288 (N_8288,N_2699,N_588);
nor U8289 (N_8289,N_1463,N_4784);
nand U8290 (N_8290,N_2797,N_3700);
nor U8291 (N_8291,N_4382,N_1441);
xnor U8292 (N_8292,N_2902,N_4126);
nor U8293 (N_8293,N_334,N_3378);
nor U8294 (N_8294,N_792,N_4263);
nor U8295 (N_8295,N_3779,N_1756);
nor U8296 (N_8296,N_2628,N_4525);
nor U8297 (N_8297,N_1212,N_4503);
and U8298 (N_8298,N_2282,N_416);
and U8299 (N_8299,N_4256,N_1899);
nand U8300 (N_8300,N_757,N_158);
and U8301 (N_8301,N_2937,N_424);
nor U8302 (N_8302,N_4354,N_2180);
and U8303 (N_8303,N_4624,N_980);
nand U8304 (N_8304,N_3138,N_1103);
nor U8305 (N_8305,N_1665,N_662);
nor U8306 (N_8306,N_4796,N_2728);
nand U8307 (N_8307,N_3580,N_2902);
nor U8308 (N_8308,N_1610,N_238);
nor U8309 (N_8309,N_2015,N_1097);
nor U8310 (N_8310,N_3939,N_4381);
nor U8311 (N_8311,N_287,N_2545);
nand U8312 (N_8312,N_3339,N_3241);
nand U8313 (N_8313,N_1821,N_4348);
and U8314 (N_8314,N_1751,N_417);
nor U8315 (N_8315,N_3322,N_4900);
or U8316 (N_8316,N_4359,N_3796);
or U8317 (N_8317,N_2928,N_2729);
nor U8318 (N_8318,N_3076,N_1310);
or U8319 (N_8319,N_1310,N_4891);
nand U8320 (N_8320,N_4599,N_4534);
nor U8321 (N_8321,N_431,N_4946);
or U8322 (N_8322,N_1758,N_3489);
nor U8323 (N_8323,N_1583,N_52);
or U8324 (N_8324,N_343,N_825);
and U8325 (N_8325,N_3268,N_4396);
or U8326 (N_8326,N_2021,N_2438);
nor U8327 (N_8327,N_3971,N_3735);
and U8328 (N_8328,N_2923,N_1634);
or U8329 (N_8329,N_3302,N_1277);
nor U8330 (N_8330,N_2072,N_3418);
or U8331 (N_8331,N_1636,N_807);
and U8332 (N_8332,N_2958,N_4784);
nand U8333 (N_8333,N_2668,N_1166);
or U8334 (N_8334,N_2238,N_3503);
and U8335 (N_8335,N_828,N_3831);
nand U8336 (N_8336,N_480,N_4353);
nor U8337 (N_8337,N_2661,N_4522);
nor U8338 (N_8338,N_335,N_775);
nor U8339 (N_8339,N_1528,N_4215);
nor U8340 (N_8340,N_608,N_919);
nor U8341 (N_8341,N_1070,N_3337);
xnor U8342 (N_8342,N_1395,N_739);
or U8343 (N_8343,N_2819,N_4985);
or U8344 (N_8344,N_3085,N_3063);
or U8345 (N_8345,N_2080,N_601);
nor U8346 (N_8346,N_786,N_3720);
nor U8347 (N_8347,N_2645,N_964);
nor U8348 (N_8348,N_4163,N_4730);
nand U8349 (N_8349,N_3194,N_3008);
or U8350 (N_8350,N_322,N_3031);
or U8351 (N_8351,N_4424,N_3977);
nor U8352 (N_8352,N_3381,N_1258);
nor U8353 (N_8353,N_136,N_3644);
nor U8354 (N_8354,N_1248,N_2221);
and U8355 (N_8355,N_3635,N_889);
and U8356 (N_8356,N_2619,N_1666);
and U8357 (N_8357,N_1183,N_169);
nand U8358 (N_8358,N_2744,N_697);
nand U8359 (N_8359,N_4682,N_3709);
and U8360 (N_8360,N_1568,N_2075);
nand U8361 (N_8361,N_3367,N_3867);
nor U8362 (N_8362,N_2675,N_161);
nor U8363 (N_8363,N_1194,N_1174);
nor U8364 (N_8364,N_76,N_4647);
and U8365 (N_8365,N_211,N_4062);
or U8366 (N_8366,N_4852,N_1871);
and U8367 (N_8367,N_2543,N_351);
and U8368 (N_8368,N_2949,N_2052);
nand U8369 (N_8369,N_932,N_3808);
and U8370 (N_8370,N_1962,N_4988);
and U8371 (N_8371,N_3849,N_3502);
nand U8372 (N_8372,N_675,N_3321);
and U8373 (N_8373,N_2133,N_4640);
or U8374 (N_8374,N_1359,N_4290);
nor U8375 (N_8375,N_248,N_4858);
or U8376 (N_8376,N_3768,N_2133);
nand U8377 (N_8377,N_4357,N_3900);
nor U8378 (N_8378,N_847,N_4450);
nor U8379 (N_8379,N_419,N_1698);
nor U8380 (N_8380,N_4366,N_2010);
and U8381 (N_8381,N_1950,N_3000);
and U8382 (N_8382,N_1867,N_4866);
and U8383 (N_8383,N_3391,N_4031);
or U8384 (N_8384,N_4059,N_3179);
nand U8385 (N_8385,N_3160,N_322);
or U8386 (N_8386,N_4746,N_31);
or U8387 (N_8387,N_3749,N_2636);
nand U8388 (N_8388,N_345,N_3110);
or U8389 (N_8389,N_978,N_4638);
nand U8390 (N_8390,N_1193,N_4492);
or U8391 (N_8391,N_3805,N_255);
nand U8392 (N_8392,N_1002,N_2165);
or U8393 (N_8393,N_3902,N_970);
or U8394 (N_8394,N_4170,N_4302);
nand U8395 (N_8395,N_2625,N_856);
nand U8396 (N_8396,N_4367,N_3830);
and U8397 (N_8397,N_4038,N_1300);
or U8398 (N_8398,N_1737,N_81);
and U8399 (N_8399,N_833,N_4619);
nor U8400 (N_8400,N_180,N_2254);
and U8401 (N_8401,N_4438,N_267);
and U8402 (N_8402,N_3149,N_4597);
nor U8403 (N_8403,N_3507,N_1789);
or U8404 (N_8404,N_1991,N_1577);
nor U8405 (N_8405,N_1115,N_1561);
and U8406 (N_8406,N_613,N_2195);
and U8407 (N_8407,N_2222,N_2634);
or U8408 (N_8408,N_369,N_225);
nand U8409 (N_8409,N_2904,N_222);
nor U8410 (N_8410,N_4776,N_1228);
nand U8411 (N_8411,N_4400,N_634);
nor U8412 (N_8412,N_3162,N_2490);
and U8413 (N_8413,N_1468,N_2516);
nand U8414 (N_8414,N_4318,N_1188);
nor U8415 (N_8415,N_2209,N_4592);
nor U8416 (N_8416,N_4880,N_55);
and U8417 (N_8417,N_2602,N_1840);
and U8418 (N_8418,N_2983,N_1969);
or U8419 (N_8419,N_1491,N_281);
and U8420 (N_8420,N_2146,N_4839);
and U8421 (N_8421,N_1176,N_455);
nand U8422 (N_8422,N_3767,N_2893);
nand U8423 (N_8423,N_4421,N_316);
nand U8424 (N_8424,N_4055,N_3827);
nor U8425 (N_8425,N_3270,N_3495);
or U8426 (N_8426,N_3682,N_4408);
and U8427 (N_8427,N_4846,N_3537);
nand U8428 (N_8428,N_2417,N_1431);
nand U8429 (N_8429,N_1902,N_3168);
xnor U8430 (N_8430,N_306,N_623);
or U8431 (N_8431,N_3732,N_760);
nand U8432 (N_8432,N_2581,N_345);
nand U8433 (N_8433,N_2453,N_4931);
and U8434 (N_8434,N_3613,N_3544);
nor U8435 (N_8435,N_2247,N_54);
and U8436 (N_8436,N_769,N_1651);
nand U8437 (N_8437,N_1793,N_4633);
and U8438 (N_8438,N_3925,N_4962);
nor U8439 (N_8439,N_1719,N_2793);
and U8440 (N_8440,N_193,N_3358);
or U8441 (N_8441,N_1973,N_2017);
nor U8442 (N_8442,N_4143,N_29);
and U8443 (N_8443,N_2341,N_1727);
nor U8444 (N_8444,N_3585,N_2937);
nand U8445 (N_8445,N_3711,N_2250);
nand U8446 (N_8446,N_3257,N_2160);
nand U8447 (N_8447,N_2604,N_59);
or U8448 (N_8448,N_2534,N_1177);
nor U8449 (N_8449,N_251,N_2597);
and U8450 (N_8450,N_4497,N_4466);
nand U8451 (N_8451,N_1496,N_2429);
nor U8452 (N_8452,N_3927,N_2494);
nor U8453 (N_8453,N_456,N_1987);
and U8454 (N_8454,N_931,N_4955);
nand U8455 (N_8455,N_3775,N_2652);
or U8456 (N_8456,N_1423,N_150);
nand U8457 (N_8457,N_2918,N_725);
or U8458 (N_8458,N_2050,N_1252);
or U8459 (N_8459,N_3564,N_2780);
or U8460 (N_8460,N_2234,N_4473);
and U8461 (N_8461,N_1946,N_4813);
nor U8462 (N_8462,N_3974,N_3525);
nand U8463 (N_8463,N_3099,N_2016);
and U8464 (N_8464,N_4407,N_1544);
and U8465 (N_8465,N_1714,N_863);
or U8466 (N_8466,N_3603,N_2994);
and U8467 (N_8467,N_2700,N_1883);
nor U8468 (N_8468,N_587,N_3880);
nand U8469 (N_8469,N_1175,N_668);
nand U8470 (N_8470,N_4575,N_4967);
nor U8471 (N_8471,N_3342,N_508);
nand U8472 (N_8472,N_1106,N_4881);
or U8473 (N_8473,N_596,N_4085);
nand U8474 (N_8474,N_345,N_2735);
and U8475 (N_8475,N_4874,N_2154);
and U8476 (N_8476,N_4810,N_2419);
and U8477 (N_8477,N_4025,N_3258);
or U8478 (N_8478,N_4889,N_4838);
and U8479 (N_8479,N_939,N_3459);
or U8480 (N_8480,N_2821,N_2571);
nand U8481 (N_8481,N_4899,N_2490);
nor U8482 (N_8482,N_1282,N_2739);
or U8483 (N_8483,N_789,N_3543);
or U8484 (N_8484,N_3521,N_1378);
nor U8485 (N_8485,N_3855,N_3664);
nor U8486 (N_8486,N_187,N_1458);
nand U8487 (N_8487,N_4378,N_2956);
nor U8488 (N_8488,N_4483,N_4602);
nor U8489 (N_8489,N_2872,N_234);
or U8490 (N_8490,N_3670,N_1643);
xnor U8491 (N_8491,N_4562,N_840);
nor U8492 (N_8492,N_4109,N_4275);
and U8493 (N_8493,N_4035,N_641);
nand U8494 (N_8494,N_3652,N_1098);
or U8495 (N_8495,N_1108,N_4333);
nor U8496 (N_8496,N_2208,N_3225);
or U8497 (N_8497,N_1276,N_2002);
or U8498 (N_8498,N_4713,N_2803);
nand U8499 (N_8499,N_2299,N_4845);
and U8500 (N_8500,N_1951,N_4916);
nor U8501 (N_8501,N_1674,N_1813);
and U8502 (N_8502,N_4592,N_1731);
nand U8503 (N_8503,N_2670,N_3463);
nor U8504 (N_8504,N_1730,N_1111);
or U8505 (N_8505,N_2290,N_1821);
nor U8506 (N_8506,N_4831,N_4109);
nand U8507 (N_8507,N_2170,N_2027);
or U8508 (N_8508,N_4610,N_52);
nand U8509 (N_8509,N_3995,N_2494);
nor U8510 (N_8510,N_4524,N_1547);
nand U8511 (N_8511,N_3605,N_3563);
and U8512 (N_8512,N_2735,N_2596);
nor U8513 (N_8513,N_2170,N_1666);
nand U8514 (N_8514,N_4720,N_3656);
nand U8515 (N_8515,N_115,N_4312);
nor U8516 (N_8516,N_3575,N_1093);
or U8517 (N_8517,N_3376,N_4666);
and U8518 (N_8518,N_4504,N_1156);
and U8519 (N_8519,N_628,N_56);
and U8520 (N_8520,N_850,N_2146);
nand U8521 (N_8521,N_85,N_4985);
nand U8522 (N_8522,N_877,N_647);
nand U8523 (N_8523,N_2952,N_149);
nand U8524 (N_8524,N_629,N_1327);
and U8525 (N_8525,N_3435,N_4709);
nand U8526 (N_8526,N_819,N_337);
and U8527 (N_8527,N_3022,N_191);
or U8528 (N_8528,N_2932,N_3471);
or U8529 (N_8529,N_900,N_4250);
or U8530 (N_8530,N_3233,N_3904);
or U8531 (N_8531,N_4152,N_4225);
nor U8532 (N_8532,N_2877,N_1961);
nor U8533 (N_8533,N_2754,N_359);
nand U8534 (N_8534,N_727,N_2535);
nand U8535 (N_8535,N_3000,N_4430);
nand U8536 (N_8536,N_4289,N_4617);
nand U8537 (N_8537,N_4415,N_4259);
and U8538 (N_8538,N_4206,N_623);
nand U8539 (N_8539,N_2776,N_1281);
nor U8540 (N_8540,N_3798,N_2173);
and U8541 (N_8541,N_756,N_3430);
and U8542 (N_8542,N_174,N_162);
nor U8543 (N_8543,N_1576,N_3154);
or U8544 (N_8544,N_2720,N_4448);
and U8545 (N_8545,N_1881,N_2114);
nor U8546 (N_8546,N_1374,N_4304);
and U8547 (N_8547,N_724,N_2987);
nor U8548 (N_8548,N_843,N_2179);
nand U8549 (N_8549,N_3843,N_2498);
nor U8550 (N_8550,N_3063,N_2947);
nand U8551 (N_8551,N_2832,N_3080);
nor U8552 (N_8552,N_4089,N_2035);
nand U8553 (N_8553,N_3440,N_1925);
and U8554 (N_8554,N_1114,N_1312);
nand U8555 (N_8555,N_3126,N_2712);
or U8556 (N_8556,N_4737,N_1115);
nand U8557 (N_8557,N_37,N_1576);
nand U8558 (N_8558,N_561,N_3459);
and U8559 (N_8559,N_4918,N_4337);
and U8560 (N_8560,N_2447,N_508);
nand U8561 (N_8561,N_4312,N_388);
and U8562 (N_8562,N_2703,N_847);
nand U8563 (N_8563,N_4886,N_564);
and U8564 (N_8564,N_869,N_2911);
nor U8565 (N_8565,N_3346,N_1001);
nand U8566 (N_8566,N_4152,N_1670);
and U8567 (N_8567,N_2743,N_2910);
nand U8568 (N_8568,N_1938,N_1347);
nor U8569 (N_8569,N_2689,N_4711);
or U8570 (N_8570,N_242,N_4680);
nand U8571 (N_8571,N_610,N_2239);
and U8572 (N_8572,N_996,N_4906);
nor U8573 (N_8573,N_1827,N_595);
nand U8574 (N_8574,N_631,N_4634);
or U8575 (N_8575,N_535,N_520);
nand U8576 (N_8576,N_3597,N_3560);
and U8577 (N_8577,N_2616,N_2534);
nor U8578 (N_8578,N_2808,N_1191);
and U8579 (N_8579,N_1590,N_4353);
or U8580 (N_8580,N_3476,N_3581);
nand U8581 (N_8581,N_1695,N_3382);
nand U8582 (N_8582,N_2224,N_2760);
or U8583 (N_8583,N_3874,N_3907);
and U8584 (N_8584,N_74,N_2977);
nand U8585 (N_8585,N_1690,N_1073);
nand U8586 (N_8586,N_2240,N_4868);
nand U8587 (N_8587,N_803,N_4919);
nor U8588 (N_8588,N_1652,N_936);
nor U8589 (N_8589,N_754,N_134);
and U8590 (N_8590,N_757,N_118);
and U8591 (N_8591,N_3881,N_2223);
nand U8592 (N_8592,N_795,N_4264);
and U8593 (N_8593,N_3202,N_708);
or U8594 (N_8594,N_2077,N_2588);
xnor U8595 (N_8595,N_1083,N_1601);
and U8596 (N_8596,N_478,N_4407);
and U8597 (N_8597,N_1980,N_2509);
or U8598 (N_8598,N_3910,N_1895);
nand U8599 (N_8599,N_951,N_2980);
nand U8600 (N_8600,N_3540,N_2254);
nor U8601 (N_8601,N_3863,N_1322);
or U8602 (N_8602,N_4865,N_3691);
or U8603 (N_8603,N_3956,N_18);
or U8604 (N_8604,N_456,N_1839);
nor U8605 (N_8605,N_4023,N_2765);
or U8606 (N_8606,N_2862,N_647);
nor U8607 (N_8607,N_3287,N_2707);
nor U8608 (N_8608,N_1861,N_585);
nor U8609 (N_8609,N_4847,N_3166);
or U8610 (N_8610,N_4903,N_1990);
or U8611 (N_8611,N_93,N_2833);
or U8612 (N_8612,N_3294,N_2369);
and U8613 (N_8613,N_4004,N_1998);
xor U8614 (N_8614,N_3306,N_1910);
or U8615 (N_8615,N_4103,N_4328);
or U8616 (N_8616,N_1854,N_3607);
nand U8617 (N_8617,N_1111,N_259);
or U8618 (N_8618,N_3214,N_2477);
or U8619 (N_8619,N_160,N_4609);
nor U8620 (N_8620,N_3108,N_1743);
and U8621 (N_8621,N_3960,N_3898);
and U8622 (N_8622,N_754,N_2125);
nand U8623 (N_8623,N_3301,N_4616);
and U8624 (N_8624,N_2200,N_1565);
or U8625 (N_8625,N_598,N_2691);
or U8626 (N_8626,N_351,N_2058);
and U8627 (N_8627,N_2141,N_1682);
or U8628 (N_8628,N_4533,N_3720);
and U8629 (N_8629,N_318,N_275);
or U8630 (N_8630,N_2712,N_3837);
and U8631 (N_8631,N_2060,N_2835);
or U8632 (N_8632,N_4799,N_2179);
nor U8633 (N_8633,N_193,N_3930);
and U8634 (N_8634,N_2831,N_2621);
nor U8635 (N_8635,N_2878,N_4372);
nor U8636 (N_8636,N_1790,N_2867);
nand U8637 (N_8637,N_3069,N_1167);
nor U8638 (N_8638,N_1796,N_4329);
nand U8639 (N_8639,N_477,N_1644);
and U8640 (N_8640,N_446,N_2204);
nand U8641 (N_8641,N_811,N_3300);
nand U8642 (N_8642,N_1784,N_79);
nor U8643 (N_8643,N_1720,N_716);
and U8644 (N_8644,N_4959,N_147);
and U8645 (N_8645,N_547,N_2566);
and U8646 (N_8646,N_4232,N_4327);
and U8647 (N_8647,N_1779,N_4643);
and U8648 (N_8648,N_364,N_1853);
nor U8649 (N_8649,N_2374,N_851);
nor U8650 (N_8650,N_4330,N_2634);
nand U8651 (N_8651,N_4384,N_4527);
nor U8652 (N_8652,N_4462,N_4985);
nand U8653 (N_8653,N_189,N_4588);
nor U8654 (N_8654,N_2916,N_2471);
nand U8655 (N_8655,N_3893,N_726);
or U8656 (N_8656,N_763,N_115);
nand U8657 (N_8657,N_537,N_3013);
and U8658 (N_8658,N_1540,N_193);
nand U8659 (N_8659,N_4062,N_3179);
nand U8660 (N_8660,N_601,N_4794);
nor U8661 (N_8661,N_1080,N_3119);
or U8662 (N_8662,N_4308,N_3211);
nand U8663 (N_8663,N_1207,N_4209);
and U8664 (N_8664,N_349,N_2197);
and U8665 (N_8665,N_1487,N_265);
nor U8666 (N_8666,N_3930,N_3755);
and U8667 (N_8667,N_2211,N_691);
and U8668 (N_8668,N_3994,N_1773);
nand U8669 (N_8669,N_4269,N_3332);
nand U8670 (N_8670,N_3216,N_2210);
and U8671 (N_8671,N_3262,N_1986);
nand U8672 (N_8672,N_4831,N_3160);
and U8673 (N_8673,N_1619,N_597);
or U8674 (N_8674,N_521,N_1391);
and U8675 (N_8675,N_273,N_2565);
nor U8676 (N_8676,N_4446,N_2862);
and U8677 (N_8677,N_2953,N_778);
or U8678 (N_8678,N_4420,N_827);
or U8679 (N_8679,N_4663,N_4849);
xnor U8680 (N_8680,N_2200,N_3509);
and U8681 (N_8681,N_2967,N_302);
and U8682 (N_8682,N_1389,N_3654);
and U8683 (N_8683,N_544,N_3803);
or U8684 (N_8684,N_1925,N_4549);
nand U8685 (N_8685,N_1704,N_630);
nor U8686 (N_8686,N_3515,N_4235);
and U8687 (N_8687,N_761,N_4090);
nand U8688 (N_8688,N_1196,N_1471);
and U8689 (N_8689,N_2519,N_2864);
and U8690 (N_8690,N_4973,N_1889);
nor U8691 (N_8691,N_155,N_3046);
nor U8692 (N_8692,N_973,N_1765);
nand U8693 (N_8693,N_789,N_4684);
and U8694 (N_8694,N_4318,N_3625);
or U8695 (N_8695,N_1817,N_836);
nor U8696 (N_8696,N_219,N_2263);
or U8697 (N_8697,N_805,N_3088);
and U8698 (N_8698,N_3492,N_1288);
or U8699 (N_8699,N_4460,N_555);
nand U8700 (N_8700,N_1895,N_4147);
and U8701 (N_8701,N_4096,N_2758);
nand U8702 (N_8702,N_303,N_3265);
and U8703 (N_8703,N_2588,N_3331);
nor U8704 (N_8704,N_4798,N_4157);
or U8705 (N_8705,N_649,N_2777);
nand U8706 (N_8706,N_3680,N_1586);
or U8707 (N_8707,N_4940,N_1169);
nand U8708 (N_8708,N_4342,N_608);
or U8709 (N_8709,N_2314,N_679);
or U8710 (N_8710,N_1177,N_4010);
nor U8711 (N_8711,N_1086,N_4255);
nand U8712 (N_8712,N_1951,N_2535);
nand U8713 (N_8713,N_1750,N_2238);
nand U8714 (N_8714,N_4071,N_2841);
nand U8715 (N_8715,N_2568,N_4921);
nand U8716 (N_8716,N_4944,N_3778);
and U8717 (N_8717,N_1698,N_4033);
nand U8718 (N_8718,N_97,N_197);
and U8719 (N_8719,N_172,N_2757);
and U8720 (N_8720,N_2455,N_2759);
nor U8721 (N_8721,N_4156,N_4427);
nor U8722 (N_8722,N_1383,N_3945);
nand U8723 (N_8723,N_3376,N_3365);
or U8724 (N_8724,N_4288,N_1429);
or U8725 (N_8725,N_2425,N_1511);
and U8726 (N_8726,N_1289,N_473);
nor U8727 (N_8727,N_4821,N_516);
and U8728 (N_8728,N_2532,N_3543);
or U8729 (N_8729,N_3282,N_2312);
or U8730 (N_8730,N_4043,N_2685);
nand U8731 (N_8731,N_3390,N_4337);
and U8732 (N_8732,N_144,N_723);
and U8733 (N_8733,N_3604,N_2583);
and U8734 (N_8734,N_2124,N_1555);
or U8735 (N_8735,N_951,N_770);
nor U8736 (N_8736,N_4721,N_977);
nor U8737 (N_8737,N_4762,N_3738);
and U8738 (N_8738,N_3524,N_1444);
and U8739 (N_8739,N_3965,N_3406);
and U8740 (N_8740,N_1051,N_3204);
nor U8741 (N_8741,N_388,N_1179);
nand U8742 (N_8742,N_4543,N_2108);
nor U8743 (N_8743,N_294,N_1397);
nor U8744 (N_8744,N_3977,N_103);
nor U8745 (N_8745,N_4847,N_607);
or U8746 (N_8746,N_2906,N_4994);
nor U8747 (N_8747,N_3825,N_1314);
nor U8748 (N_8748,N_1299,N_1360);
nand U8749 (N_8749,N_1873,N_613);
nand U8750 (N_8750,N_2907,N_468);
and U8751 (N_8751,N_1098,N_242);
nand U8752 (N_8752,N_677,N_2667);
and U8753 (N_8753,N_561,N_2166);
and U8754 (N_8754,N_4635,N_1797);
nand U8755 (N_8755,N_3099,N_2474);
and U8756 (N_8756,N_2366,N_1884);
nand U8757 (N_8757,N_4872,N_2437);
and U8758 (N_8758,N_3024,N_1056);
nand U8759 (N_8759,N_2616,N_1611);
nand U8760 (N_8760,N_2099,N_264);
nor U8761 (N_8761,N_1652,N_3339);
nor U8762 (N_8762,N_148,N_3536);
nor U8763 (N_8763,N_2708,N_4116);
nand U8764 (N_8764,N_2162,N_2128);
and U8765 (N_8765,N_4612,N_3979);
nand U8766 (N_8766,N_2879,N_96);
nand U8767 (N_8767,N_2141,N_657);
or U8768 (N_8768,N_3627,N_825);
or U8769 (N_8769,N_2129,N_371);
and U8770 (N_8770,N_3017,N_891);
and U8771 (N_8771,N_3974,N_3892);
nand U8772 (N_8772,N_51,N_1147);
and U8773 (N_8773,N_1470,N_714);
and U8774 (N_8774,N_1459,N_2449);
or U8775 (N_8775,N_4609,N_3671);
or U8776 (N_8776,N_3344,N_2717);
nor U8777 (N_8777,N_3679,N_716);
nand U8778 (N_8778,N_1533,N_4991);
and U8779 (N_8779,N_4210,N_2119);
nor U8780 (N_8780,N_3392,N_1267);
nor U8781 (N_8781,N_276,N_2260);
nor U8782 (N_8782,N_4175,N_259);
or U8783 (N_8783,N_2772,N_3844);
or U8784 (N_8784,N_4864,N_1716);
or U8785 (N_8785,N_2936,N_4637);
or U8786 (N_8786,N_483,N_1138);
xor U8787 (N_8787,N_4966,N_4680);
and U8788 (N_8788,N_1530,N_1104);
nor U8789 (N_8789,N_4931,N_3384);
nand U8790 (N_8790,N_2102,N_4989);
nand U8791 (N_8791,N_4766,N_640);
or U8792 (N_8792,N_3641,N_1904);
nand U8793 (N_8793,N_45,N_4080);
or U8794 (N_8794,N_1937,N_520);
and U8795 (N_8795,N_1428,N_1800);
nand U8796 (N_8796,N_2019,N_2654);
nand U8797 (N_8797,N_4740,N_3679);
or U8798 (N_8798,N_694,N_2929);
nand U8799 (N_8799,N_1585,N_4185);
nand U8800 (N_8800,N_3267,N_223);
nand U8801 (N_8801,N_4603,N_1495);
and U8802 (N_8802,N_4317,N_102);
or U8803 (N_8803,N_3912,N_392);
nor U8804 (N_8804,N_1504,N_1848);
nand U8805 (N_8805,N_2308,N_399);
nor U8806 (N_8806,N_3023,N_51);
nand U8807 (N_8807,N_2934,N_2806);
nand U8808 (N_8808,N_2650,N_994);
nand U8809 (N_8809,N_98,N_1430);
and U8810 (N_8810,N_4331,N_2759);
or U8811 (N_8811,N_4152,N_4232);
nor U8812 (N_8812,N_3484,N_3);
and U8813 (N_8813,N_32,N_4002);
nand U8814 (N_8814,N_4287,N_3165);
nor U8815 (N_8815,N_3637,N_1844);
and U8816 (N_8816,N_2231,N_4200);
and U8817 (N_8817,N_934,N_4186);
or U8818 (N_8818,N_1417,N_2091);
or U8819 (N_8819,N_787,N_693);
or U8820 (N_8820,N_2223,N_2982);
nor U8821 (N_8821,N_4940,N_923);
and U8822 (N_8822,N_4464,N_216);
nand U8823 (N_8823,N_2046,N_4969);
nand U8824 (N_8824,N_3749,N_2110);
nand U8825 (N_8825,N_764,N_4936);
or U8826 (N_8826,N_4689,N_2318);
and U8827 (N_8827,N_3881,N_3267);
nor U8828 (N_8828,N_4606,N_3139);
or U8829 (N_8829,N_3192,N_4102);
nand U8830 (N_8830,N_1936,N_3946);
nor U8831 (N_8831,N_4787,N_475);
nand U8832 (N_8832,N_2641,N_1282);
nand U8833 (N_8833,N_2259,N_3728);
and U8834 (N_8834,N_4724,N_3434);
nor U8835 (N_8835,N_544,N_3157);
and U8836 (N_8836,N_4875,N_1405);
and U8837 (N_8837,N_3617,N_4108);
nand U8838 (N_8838,N_2910,N_1500);
nand U8839 (N_8839,N_4303,N_4150);
nor U8840 (N_8840,N_576,N_1062);
nand U8841 (N_8841,N_385,N_4713);
or U8842 (N_8842,N_1954,N_1193);
nor U8843 (N_8843,N_4717,N_1341);
nor U8844 (N_8844,N_3537,N_3851);
and U8845 (N_8845,N_1512,N_1528);
nand U8846 (N_8846,N_3184,N_633);
and U8847 (N_8847,N_3477,N_4849);
and U8848 (N_8848,N_496,N_1917);
and U8849 (N_8849,N_4765,N_3529);
nand U8850 (N_8850,N_4529,N_2851);
and U8851 (N_8851,N_3057,N_1225);
nor U8852 (N_8852,N_2034,N_1699);
or U8853 (N_8853,N_105,N_321);
nand U8854 (N_8854,N_2909,N_344);
nor U8855 (N_8855,N_3213,N_2390);
or U8856 (N_8856,N_2312,N_4317);
nor U8857 (N_8857,N_1270,N_3756);
nand U8858 (N_8858,N_4259,N_2995);
nor U8859 (N_8859,N_1476,N_1585);
nor U8860 (N_8860,N_493,N_3631);
nor U8861 (N_8861,N_514,N_4972);
or U8862 (N_8862,N_4654,N_535);
and U8863 (N_8863,N_886,N_3982);
xnor U8864 (N_8864,N_4424,N_4076);
nor U8865 (N_8865,N_4192,N_4528);
and U8866 (N_8866,N_3011,N_3282);
nor U8867 (N_8867,N_4808,N_2490);
nor U8868 (N_8868,N_1779,N_1658);
nor U8869 (N_8869,N_4418,N_741);
nand U8870 (N_8870,N_2397,N_4451);
nor U8871 (N_8871,N_761,N_360);
nand U8872 (N_8872,N_1945,N_1275);
nand U8873 (N_8873,N_3437,N_950);
or U8874 (N_8874,N_836,N_4835);
xor U8875 (N_8875,N_3540,N_2333);
and U8876 (N_8876,N_4465,N_1825);
nor U8877 (N_8877,N_951,N_1535);
and U8878 (N_8878,N_644,N_3958);
or U8879 (N_8879,N_3895,N_3865);
and U8880 (N_8880,N_4264,N_4437);
xor U8881 (N_8881,N_2519,N_2598);
or U8882 (N_8882,N_2993,N_1666);
xor U8883 (N_8883,N_4820,N_4844);
nor U8884 (N_8884,N_1765,N_3796);
and U8885 (N_8885,N_1684,N_4920);
and U8886 (N_8886,N_2324,N_2821);
and U8887 (N_8887,N_1502,N_1676);
and U8888 (N_8888,N_1417,N_4835);
nor U8889 (N_8889,N_731,N_3087);
nor U8890 (N_8890,N_1040,N_1386);
and U8891 (N_8891,N_3092,N_3477);
nand U8892 (N_8892,N_2746,N_3648);
or U8893 (N_8893,N_3145,N_2529);
or U8894 (N_8894,N_2128,N_3805);
nand U8895 (N_8895,N_2418,N_4068);
or U8896 (N_8896,N_4580,N_4075);
nor U8897 (N_8897,N_698,N_3222);
or U8898 (N_8898,N_4511,N_2382);
nand U8899 (N_8899,N_5,N_1791);
nor U8900 (N_8900,N_4116,N_3846);
nor U8901 (N_8901,N_2468,N_4193);
nand U8902 (N_8902,N_3151,N_277);
or U8903 (N_8903,N_3262,N_4085);
nand U8904 (N_8904,N_383,N_2410);
and U8905 (N_8905,N_3540,N_2751);
nand U8906 (N_8906,N_2711,N_148);
nor U8907 (N_8907,N_858,N_1948);
nand U8908 (N_8908,N_4116,N_4805);
nor U8909 (N_8909,N_4155,N_2943);
nand U8910 (N_8910,N_3126,N_1619);
nor U8911 (N_8911,N_503,N_2933);
and U8912 (N_8912,N_1771,N_2268);
nand U8913 (N_8913,N_2529,N_909);
nor U8914 (N_8914,N_3625,N_3526);
nor U8915 (N_8915,N_4508,N_1463);
nand U8916 (N_8916,N_3662,N_1225);
nand U8917 (N_8917,N_3495,N_1397);
or U8918 (N_8918,N_2264,N_735);
and U8919 (N_8919,N_2066,N_2167);
nor U8920 (N_8920,N_1706,N_4550);
and U8921 (N_8921,N_2768,N_2012);
or U8922 (N_8922,N_3073,N_192);
nand U8923 (N_8923,N_3362,N_3200);
nor U8924 (N_8924,N_192,N_4170);
and U8925 (N_8925,N_1826,N_1521);
or U8926 (N_8926,N_467,N_307);
nor U8927 (N_8927,N_1533,N_4241);
and U8928 (N_8928,N_3014,N_1736);
and U8929 (N_8929,N_2748,N_1322);
and U8930 (N_8930,N_2099,N_4468);
or U8931 (N_8931,N_4605,N_1236);
nor U8932 (N_8932,N_3363,N_2478);
or U8933 (N_8933,N_4682,N_3338);
nand U8934 (N_8934,N_3006,N_2769);
and U8935 (N_8935,N_2977,N_349);
and U8936 (N_8936,N_3892,N_2703);
nand U8937 (N_8937,N_2703,N_3937);
nor U8938 (N_8938,N_11,N_1929);
nand U8939 (N_8939,N_3483,N_4409);
nor U8940 (N_8940,N_3555,N_1870);
nand U8941 (N_8941,N_4298,N_3150);
and U8942 (N_8942,N_3254,N_61);
and U8943 (N_8943,N_2015,N_84);
or U8944 (N_8944,N_1923,N_1794);
nor U8945 (N_8945,N_3644,N_848);
nor U8946 (N_8946,N_3077,N_3678);
or U8947 (N_8947,N_1649,N_4775);
or U8948 (N_8948,N_2024,N_633);
nand U8949 (N_8949,N_4914,N_3326);
or U8950 (N_8950,N_4762,N_1461);
nand U8951 (N_8951,N_4190,N_4502);
nand U8952 (N_8952,N_50,N_419);
and U8953 (N_8953,N_4789,N_1441);
and U8954 (N_8954,N_4185,N_3741);
nand U8955 (N_8955,N_4480,N_1484);
nor U8956 (N_8956,N_4485,N_4964);
nand U8957 (N_8957,N_684,N_1777);
or U8958 (N_8958,N_1614,N_4662);
nand U8959 (N_8959,N_2930,N_774);
and U8960 (N_8960,N_2309,N_4579);
nand U8961 (N_8961,N_2735,N_1557);
and U8962 (N_8962,N_1068,N_3774);
or U8963 (N_8963,N_4996,N_2240);
or U8964 (N_8964,N_4424,N_1940);
or U8965 (N_8965,N_2188,N_4489);
or U8966 (N_8966,N_935,N_2850);
or U8967 (N_8967,N_3434,N_1479);
and U8968 (N_8968,N_775,N_4946);
nand U8969 (N_8969,N_1189,N_1757);
nand U8970 (N_8970,N_2599,N_10);
or U8971 (N_8971,N_3283,N_590);
or U8972 (N_8972,N_1536,N_2344);
nor U8973 (N_8973,N_1101,N_3012);
and U8974 (N_8974,N_598,N_1945);
or U8975 (N_8975,N_4733,N_3574);
nand U8976 (N_8976,N_2758,N_264);
nor U8977 (N_8977,N_4435,N_4726);
and U8978 (N_8978,N_4444,N_1620);
and U8979 (N_8979,N_275,N_4764);
nand U8980 (N_8980,N_160,N_610);
nor U8981 (N_8981,N_245,N_4841);
and U8982 (N_8982,N_513,N_728);
nor U8983 (N_8983,N_3228,N_21);
or U8984 (N_8984,N_3818,N_234);
nand U8985 (N_8985,N_2233,N_3291);
and U8986 (N_8986,N_2938,N_4510);
and U8987 (N_8987,N_1448,N_3830);
or U8988 (N_8988,N_1873,N_4707);
nor U8989 (N_8989,N_3835,N_2132);
nor U8990 (N_8990,N_1784,N_3940);
and U8991 (N_8991,N_4053,N_1895);
nor U8992 (N_8992,N_1377,N_2284);
and U8993 (N_8993,N_2003,N_792);
and U8994 (N_8994,N_1542,N_3183);
nor U8995 (N_8995,N_2098,N_3760);
or U8996 (N_8996,N_3528,N_1088);
nor U8997 (N_8997,N_2975,N_4517);
nor U8998 (N_8998,N_486,N_195);
nand U8999 (N_8999,N_4968,N_2781);
nor U9000 (N_9000,N_1839,N_1610);
nand U9001 (N_9001,N_3820,N_2136);
nor U9002 (N_9002,N_2196,N_1024);
and U9003 (N_9003,N_1035,N_2589);
or U9004 (N_9004,N_875,N_1854);
and U9005 (N_9005,N_3424,N_289);
or U9006 (N_9006,N_4082,N_1890);
and U9007 (N_9007,N_2522,N_4326);
and U9008 (N_9008,N_4829,N_4640);
or U9009 (N_9009,N_3582,N_532);
and U9010 (N_9010,N_1171,N_1609);
or U9011 (N_9011,N_4790,N_3826);
or U9012 (N_9012,N_1709,N_2276);
nand U9013 (N_9013,N_3178,N_2034);
nor U9014 (N_9014,N_4539,N_1185);
or U9015 (N_9015,N_1345,N_53);
nor U9016 (N_9016,N_248,N_380);
and U9017 (N_9017,N_1199,N_663);
and U9018 (N_9018,N_4881,N_2370);
and U9019 (N_9019,N_4659,N_2108);
nand U9020 (N_9020,N_149,N_1131);
and U9021 (N_9021,N_2669,N_3388);
nand U9022 (N_9022,N_3061,N_355);
and U9023 (N_9023,N_3983,N_4840);
xnor U9024 (N_9024,N_4380,N_307);
and U9025 (N_9025,N_669,N_2622);
or U9026 (N_9026,N_829,N_2483);
nor U9027 (N_9027,N_3401,N_4027);
nand U9028 (N_9028,N_2369,N_2483);
and U9029 (N_9029,N_756,N_1453);
nand U9030 (N_9030,N_646,N_1455);
nand U9031 (N_9031,N_1286,N_762);
or U9032 (N_9032,N_961,N_3156);
nand U9033 (N_9033,N_4379,N_4486);
nor U9034 (N_9034,N_1622,N_1207);
nor U9035 (N_9035,N_4535,N_3172);
and U9036 (N_9036,N_2283,N_650);
nor U9037 (N_9037,N_2818,N_4746);
nand U9038 (N_9038,N_715,N_1287);
nand U9039 (N_9039,N_4735,N_1534);
or U9040 (N_9040,N_718,N_1869);
or U9041 (N_9041,N_2710,N_2341);
or U9042 (N_9042,N_1523,N_2697);
nand U9043 (N_9043,N_4081,N_2629);
nand U9044 (N_9044,N_3852,N_1058);
nand U9045 (N_9045,N_4461,N_1724);
and U9046 (N_9046,N_281,N_815);
nand U9047 (N_9047,N_627,N_832);
nand U9048 (N_9048,N_3594,N_539);
nand U9049 (N_9049,N_896,N_111);
and U9050 (N_9050,N_4392,N_1975);
and U9051 (N_9051,N_4491,N_978);
or U9052 (N_9052,N_4314,N_375);
nor U9053 (N_9053,N_3666,N_808);
nand U9054 (N_9054,N_4502,N_134);
and U9055 (N_9055,N_2804,N_4085);
or U9056 (N_9056,N_1407,N_3149);
nor U9057 (N_9057,N_1718,N_1021);
nand U9058 (N_9058,N_4281,N_4044);
and U9059 (N_9059,N_3564,N_2238);
or U9060 (N_9060,N_3604,N_1795);
and U9061 (N_9061,N_1267,N_942);
nor U9062 (N_9062,N_2206,N_3949);
and U9063 (N_9063,N_2128,N_2279);
and U9064 (N_9064,N_537,N_2738);
nor U9065 (N_9065,N_1145,N_2058);
nor U9066 (N_9066,N_3750,N_879);
and U9067 (N_9067,N_2903,N_3938);
nand U9068 (N_9068,N_3190,N_278);
nand U9069 (N_9069,N_2926,N_2645);
and U9070 (N_9070,N_574,N_4484);
or U9071 (N_9071,N_4923,N_4858);
nor U9072 (N_9072,N_3447,N_3632);
nand U9073 (N_9073,N_4241,N_2386);
or U9074 (N_9074,N_3321,N_1696);
nand U9075 (N_9075,N_4735,N_4560);
or U9076 (N_9076,N_2594,N_4080);
and U9077 (N_9077,N_4902,N_4360);
or U9078 (N_9078,N_280,N_1643);
or U9079 (N_9079,N_1497,N_3091);
nor U9080 (N_9080,N_1672,N_3945);
nand U9081 (N_9081,N_916,N_3047);
nand U9082 (N_9082,N_71,N_1729);
and U9083 (N_9083,N_3657,N_275);
and U9084 (N_9084,N_443,N_4410);
nor U9085 (N_9085,N_642,N_3467);
or U9086 (N_9086,N_4257,N_4368);
nand U9087 (N_9087,N_782,N_1039);
nand U9088 (N_9088,N_1090,N_1859);
or U9089 (N_9089,N_4199,N_1753);
nor U9090 (N_9090,N_866,N_3094);
nor U9091 (N_9091,N_4408,N_1667);
nand U9092 (N_9092,N_951,N_1105);
nor U9093 (N_9093,N_1411,N_3328);
and U9094 (N_9094,N_4046,N_701);
nand U9095 (N_9095,N_4141,N_2871);
nor U9096 (N_9096,N_3755,N_1532);
or U9097 (N_9097,N_2398,N_3072);
or U9098 (N_9098,N_4679,N_2363);
and U9099 (N_9099,N_1750,N_2549);
and U9100 (N_9100,N_4810,N_1221);
nand U9101 (N_9101,N_1962,N_2468);
nand U9102 (N_9102,N_4686,N_3612);
nand U9103 (N_9103,N_167,N_4770);
and U9104 (N_9104,N_3815,N_571);
nor U9105 (N_9105,N_2093,N_189);
and U9106 (N_9106,N_2906,N_4849);
or U9107 (N_9107,N_4526,N_230);
nor U9108 (N_9108,N_3458,N_1274);
nand U9109 (N_9109,N_4832,N_4254);
nor U9110 (N_9110,N_4688,N_3193);
nand U9111 (N_9111,N_1783,N_1013);
or U9112 (N_9112,N_3464,N_3471);
nor U9113 (N_9113,N_4449,N_4745);
or U9114 (N_9114,N_1739,N_3114);
nand U9115 (N_9115,N_3665,N_1272);
and U9116 (N_9116,N_4843,N_2541);
nor U9117 (N_9117,N_4854,N_4155);
and U9118 (N_9118,N_2363,N_4150);
nand U9119 (N_9119,N_4164,N_1210);
nor U9120 (N_9120,N_4876,N_4337);
nor U9121 (N_9121,N_4236,N_2997);
or U9122 (N_9122,N_1299,N_1103);
nor U9123 (N_9123,N_2954,N_2142);
nand U9124 (N_9124,N_3056,N_1193);
nand U9125 (N_9125,N_2822,N_58);
and U9126 (N_9126,N_3071,N_2365);
nand U9127 (N_9127,N_2671,N_249);
nor U9128 (N_9128,N_3925,N_870);
xnor U9129 (N_9129,N_349,N_2894);
or U9130 (N_9130,N_1190,N_2399);
or U9131 (N_9131,N_3117,N_3916);
nor U9132 (N_9132,N_4346,N_3733);
or U9133 (N_9133,N_1424,N_3284);
xor U9134 (N_9134,N_3023,N_903);
nand U9135 (N_9135,N_1368,N_3177);
nand U9136 (N_9136,N_4195,N_148);
nor U9137 (N_9137,N_3075,N_3352);
nand U9138 (N_9138,N_838,N_2936);
or U9139 (N_9139,N_2301,N_4088);
or U9140 (N_9140,N_3593,N_2172);
or U9141 (N_9141,N_4485,N_4880);
nand U9142 (N_9142,N_2868,N_2946);
and U9143 (N_9143,N_3640,N_2534);
nand U9144 (N_9144,N_1869,N_4643);
nand U9145 (N_9145,N_2296,N_4656);
nor U9146 (N_9146,N_4522,N_269);
or U9147 (N_9147,N_316,N_3184);
nand U9148 (N_9148,N_973,N_4155);
and U9149 (N_9149,N_3167,N_2014);
or U9150 (N_9150,N_1195,N_991);
nor U9151 (N_9151,N_1211,N_3079);
or U9152 (N_9152,N_3156,N_1922);
nor U9153 (N_9153,N_1101,N_4940);
and U9154 (N_9154,N_1407,N_1938);
or U9155 (N_9155,N_402,N_2641);
or U9156 (N_9156,N_2851,N_3194);
or U9157 (N_9157,N_3491,N_4466);
nand U9158 (N_9158,N_3939,N_4257);
or U9159 (N_9159,N_75,N_2059);
nand U9160 (N_9160,N_4873,N_496);
nor U9161 (N_9161,N_3066,N_3861);
or U9162 (N_9162,N_4677,N_2544);
and U9163 (N_9163,N_180,N_3679);
or U9164 (N_9164,N_4621,N_2659);
nor U9165 (N_9165,N_4981,N_1385);
and U9166 (N_9166,N_3088,N_4912);
and U9167 (N_9167,N_2404,N_4492);
and U9168 (N_9168,N_457,N_4441);
or U9169 (N_9169,N_2526,N_1514);
nor U9170 (N_9170,N_455,N_3621);
or U9171 (N_9171,N_1170,N_2989);
nand U9172 (N_9172,N_4357,N_1960);
or U9173 (N_9173,N_1440,N_4497);
nand U9174 (N_9174,N_4227,N_1509);
or U9175 (N_9175,N_3371,N_212);
or U9176 (N_9176,N_2083,N_3826);
nor U9177 (N_9177,N_1016,N_4535);
and U9178 (N_9178,N_2734,N_4088);
and U9179 (N_9179,N_3756,N_92);
nand U9180 (N_9180,N_1970,N_3878);
nand U9181 (N_9181,N_3167,N_4285);
or U9182 (N_9182,N_4483,N_996);
or U9183 (N_9183,N_1887,N_1246);
or U9184 (N_9184,N_2027,N_4482);
and U9185 (N_9185,N_928,N_1447);
and U9186 (N_9186,N_235,N_3550);
nand U9187 (N_9187,N_3215,N_1575);
or U9188 (N_9188,N_4823,N_573);
or U9189 (N_9189,N_3955,N_1516);
nor U9190 (N_9190,N_480,N_722);
xor U9191 (N_9191,N_4211,N_546);
nand U9192 (N_9192,N_1137,N_4381);
nor U9193 (N_9193,N_4095,N_241);
nand U9194 (N_9194,N_2486,N_1266);
nor U9195 (N_9195,N_3413,N_1101);
nor U9196 (N_9196,N_172,N_4514);
nor U9197 (N_9197,N_2964,N_4866);
nand U9198 (N_9198,N_370,N_2212);
nor U9199 (N_9199,N_4399,N_4051);
and U9200 (N_9200,N_4745,N_1462);
nor U9201 (N_9201,N_2680,N_1492);
nor U9202 (N_9202,N_2243,N_1562);
or U9203 (N_9203,N_3538,N_4623);
nor U9204 (N_9204,N_1537,N_4497);
nand U9205 (N_9205,N_367,N_4736);
nor U9206 (N_9206,N_342,N_2752);
nor U9207 (N_9207,N_2186,N_350);
nand U9208 (N_9208,N_1298,N_622);
nor U9209 (N_9209,N_2791,N_1697);
nand U9210 (N_9210,N_4904,N_1212);
and U9211 (N_9211,N_1575,N_1165);
nor U9212 (N_9212,N_346,N_1040);
or U9213 (N_9213,N_318,N_4305);
and U9214 (N_9214,N_2900,N_224);
nor U9215 (N_9215,N_4300,N_1988);
nor U9216 (N_9216,N_640,N_2104);
and U9217 (N_9217,N_3342,N_3605);
or U9218 (N_9218,N_2946,N_4600);
nand U9219 (N_9219,N_891,N_366);
and U9220 (N_9220,N_4499,N_610);
and U9221 (N_9221,N_4632,N_1115);
nand U9222 (N_9222,N_2340,N_3131);
nor U9223 (N_9223,N_2589,N_635);
or U9224 (N_9224,N_343,N_1927);
nor U9225 (N_9225,N_1870,N_4879);
nand U9226 (N_9226,N_4038,N_1149);
nor U9227 (N_9227,N_3747,N_2804);
nand U9228 (N_9228,N_1559,N_1198);
nor U9229 (N_9229,N_47,N_4252);
nand U9230 (N_9230,N_1447,N_112);
or U9231 (N_9231,N_4376,N_2287);
and U9232 (N_9232,N_3694,N_2873);
nand U9233 (N_9233,N_1471,N_2097);
and U9234 (N_9234,N_3367,N_3372);
nor U9235 (N_9235,N_4007,N_2212);
nor U9236 (N_9236,N_3952,N_2521);
and U9237 (N_9237,N_4707,N_602);
nor U9238 (N_9238,N_2716,N_1354);
and U9239 (N_9239,N_190,N_3312);
nand U9240 (N_9240,N_2990,N_878);
nor U9241 (N_9241,N_2503,N_1533);
nor U9242 (N_9242,N_28,N_3868);
nor U9243 (N_9243,N_4490,N_3725);
and U9244 (N_9244,N_2153,N_4851);
or U9245 (N_9245,N_2767,N_4406);
nand U9246 (N_9246,N_3459,N_2080);
and U9247 (N_9247,N_336,N_1818);
and U9248 (N_9248,N_130,N_567);
nand U9249 (N_9249,N_1783,N_2542);
nand U9250 (N_9250,N_3789,N_3093);
nor U9251 (N_9251,N_2181,N_1012);
nor U9252 (N_9252,N_385,N_20);
nor U9253 (N_9253,N_281,N_523);
and U9254 (N_9254,N_1663,N_3413);
and U9255 (N_9255,N_264,N_2813);
nor U9256 (N_9256,N_952,N_4861);
nor U9257 (N_9257,N_2533,N_4707);
nor U9258 (N_9258,N_2270,N_3438);
and U9259 (N_9259,N_3474,N_1974);
nand U9260 (N_9260,N_365,N_1911);
and U9261 (N_9261,N_56,N_1431);
and U9262 (N_9262,N_4346,N_1227);
nand U9263 (N_9263,N_2835,N_3807);
nor U9264 (N_9264,N_2910,N_2228);
and U9265 (N_9265,N_2733,N_1134);
and U9266 (N_9266,N_482,N_1568);
and U9267 (N_9267,N_4722,N_4048);
nor U9268 (N_9268,N_1791,N_3909);
nor U9269 (N_9269,N_1806,N_2094);
or U9270 (N_9270,N_3168,N_3756);
or U9271 (N_9271,N_1687,N_396);
nand U9272 (N_9272,N_4565,N_14);
and U9273 (N_9273,N_461,N_886);
or U9274 (N_9274,N_2731,N_3125);
nand U9275 (N_9275,N_4187,N_232);
and U9276 (N_9276,N_1888,N_289);
or U9277 (N_9277,N_1074,N_1229);
nand U9278 (N_9278,N_357,N_325);
or U9279 (N_9279,N_2243,N_4379);
and U9280 (N_9280,N_731,N_1085);
nor U9281 (N_9281,N_3727,N_4738);
and U9282 (N_9282,N_4094,N_2445);
and U9283 (N_9283,N_1801,N_4596);
or U9284 (N_9284,N_1994,N_923);
nor U9285 (N_9285,N_1836,N_4960);
and U9286 (N_9286,N_3324,N_781);
or U9287 (N_9287,N_2031,N_4297);
and U9288 (N_9288,N_895,N_2878);
and U9289 (N_9289,N_4319,N_4514);
nor U9290 (N_9290,N_4551,N_187);
and U9291 (N_9291,N_1306,N_244);
nor U9292 (N_9292,N_4443,N_3416);
or U9293 (N_9293,N_1043,N_1585);
and U9294 (N_9294,N_1291,N_2152);
nor U9295 (N_9295,N_3614,N_634);
nor U9296 (N_9296,N_3316,N_1315);
or U9297 (N_9297,N_3499,N_1907);
nor U9298 (N_9298,N_89,N_97);
and U9299 (N_9299,N_810,N_2879);
nand U9300 (N_9300,N_4776,N_447);
or U9301 (N_9301,N_436,N_2843);
or U9302 (N_9302,N_1773,N_1708);
nor U9303 (N_9303,N_2680,N_3549);
nor U9304 (N_9304,N_1582,N_3511);
nand U9305 (N_9305,N_4694,N_3325);
nor U9306 (N_9306,N_4151,N_4662);
nor U9307 (N_9307,N_2575,N_145);
or U9308 (N_9308,N_2023,N_2466);
nor U9309 (N_9309,N_327,N_2987);
or U9310 (N_9310,N_4808,N_150);
and U9311 (N_9311,N_4575,N_4821);
nand U9312 (N_9312,N_4686,N_3291);
and U9313 (N_9313,N_1815,N_4146);
or U9314 (N_9314,N_1225,N_3368);
or U9315 (N_9315,N_3486,N_132);
or U9316 (N_9316,N_4429,N_1661);
nand U9317 (N_9317,N_2537,N_3521);
nand U9318 (N_9318,N_3217,N_1668);
nand U9319 (N_9319,N_3232,N_2916);
nand U9320 (N_9320,N_1923,N_4594);
and U9321 (N_9321,N_2522,N_3403);
nand U9322 (N_9322,N_4050,N_3885);
nor U9323 (N_9323,N_1202,N_4318);
or U9324 (N_9324,N_146,N_4004);
xnor U9325 (N_9325,N_3434,N_1053);
nor U9326 (N_9326,N_1284,N_4601);
xnor U9327 (N_9327,N_2515,N_3325);
and U9328 (N_9328,N_3284,N_780);
xnor U9329 (N_9329,N_4190,N_2720);
nor U9330 (N_9330,N_2128,N_1025);
or U9331 (N_9331,N_1703,N_4742);
nand U9332 (N_9332,N_1737,N_4290);
or U9333 (N_9333,N_2951,N_3326);
nand U9334 (N_9334,N_809,N_4811);
and U9335 (N_9335,N_2453,N_3102);
nand U9336 (N_9336,N_1381,N_4383);
nor U9337 (N_9337,N_1275,N_1704);
nand U9338 (N_9338,N_4051,N_4153);
or U9339 (N_9339,N_421,N_2738);
and U9340 (N_9340,N_4597,N_4981);
nor U9341 (N_9341,N_275,N_821);
or U9342 (N_9342,N_4434,N_2199);
and U9343 (N_9343,N_2211,N_2900);
nor U9344 (N_9344,N_2382,N_1426);
nor U9345 (N_9345,N_796,N_2971);
nor U9346 (N_9346,N_2634,N_2873);
nand U9347 (N_9347,N_2677,N_2389);
and U9348 (N_9348,N_921,N_3072);
nand U9349 (N_9349,N_3360,N_1643);
nand U9350 (N_9350,N_2727,N_874);
nand U9351 (N_9351,N_2868,N_2919);
or U9352 (N_9352,N_4942,N_4229);
and U9353 (N_9353,N_3176,N_1685);
or U9354 (N_9354,N_693,N_4982);
nor U9355 (N_9355,N_554,N_1710);
and U9356 (N_9356,N_3012,N_1054);
nand U9357 (N_9357,N_4924,N_933);
nor U9358 (N_9358,N_1587,N_4232);
or U9359 (N_9359,N_4667,N_3491);
nor U9360 (N_9360,N_4534,N_3114);
xor U9361 (N_9361,N_4559,N_790);
and U9362 (N_9362,N_1894,N_2247);
nor U9363 (N_9363,N_719,N_4670);
or U9364 (N_9364,N_3580,N_716);
nor U9365 (N_9365,N_3808,N_81);
or U9366 (N_9366,N_3390,N_2863);
nor U9367 (N_9367,N_3867,N_1803);
and U9368 (N_9368,N_2977,N_695);
nor U9369 (N_9369,N_4004,N_162);
and U9370 (N_9370,N_2666,N_4933);
nor U9371 (N_9371,N_1246,N_1729);
nor U9372 (N_9372,N_1873,N_2436);
and U9373 (N_9373,N_2460,N_1295);
and U9374 (N_9374,N_1337,N_2301);
or U9375 (N_9375,N_3956,N_2900);
or U9376 (N_9376,N_2646,N_3989);
nor U9377 (N_9377,N_1326,N_4242);
nor U9378 (N_9378,N_590,N_377);
nor U9379 (N_9379,N_4052,N_2526);
nand U9380 (N_9380,N_3240,N_4259);
nand U9381 (N_9381,N_2662,N_1822);
or U9382 (N_9382,N_2364,N_4115);
or U9383 (N_9383,N_4765,N_2221);
nor U9384 (N_9384,N_1249,N_4451);
nor U9385 (N_9385,N_4258,N_4514);
nor U9386 (N_9386,N_1090,N_1519);
nor U9387 (N_9387,N_13,N_64);
or U9388 (N_9388,N_2157,N_377);
and U9389 (N_9389,N_1732,N_1446);
nand U9390 (N_9390,N_3452,N_3435);
and U9391 (N_9391,N_636,N_1632);
and U9392 (N_9392,N_1115,N_3341);
or U9393 (N_9393,N_1962,N_2363);
nand U9394 (N_9394,N_764,N_3699);
or U9395 (N_9395,N_3611,N_268);
nand U9396 (N_9396,N_3518,N_1208);
nand U9397 (N_9397,N_3905,N_45);
or U9398 (N_9398,N_2702,N_1224);
nand U9399 (N_9399,N_1450,N_1103);
or U9400 (N_9400,N_1413,N_2676);
and U9401 (N_9401,N_1814,N_62);
or U9402 (N_9402,N_4546,N_4197);
nand U9403 (N_9403,N_2850,N_3784);
nor U9404 (N_9404,N_4847,N_4902);
nor U9405 (N_9405,N_967,N_4381);
nand U9406 (N_9406,N_1649,N_4802);
and U9407 (N_9407,N_1407,N_2213);
and U9408 (N_9408,N_3186,N_1284);
nand U9409 (N_9409,N_4164,N_1612);
nand U9410 (N_9410,N_1372,N_2790);
nand U9411 (N_9411,N_2386,N_1100);
or U9412 (N_9412,N_1404,N_2214);
nand U9413 (N_9413,N_1895,N_3680);
and U9414 (N_9414,N_4733,N_593);
or U9415 (N_9415,N_730,N_1618);
nor U9416 (N_9416,N_4173,N_2563);
nand U9417 (N_9417,N_3301,N_332);
and U9418 (N_9418,N_2122,N_1225);
or U9419 (N_9419,N_1977,N_4206);
and U9420 (N_9420,N_4481,N_4081);
or U9421 (N_9421,N_2548,N_4371);
nor U9422 (N_9422,N_2096,N_2867);
or U9423 (N_9423,N_4762,N_4583);
nand U9424 (N_9424,N_2027,N_1764);
and U9425 (N_9425,N_462,N_3936);
or U9426 (N_9426,N_2969,N_4014);
nor U9427 (N_9427,N_4352,N_3605);
and U9428 (N_9428,N_4451,N_288);
nor U9429 (N_9429,N_236,N_1426);
nand U9430 (N_9430,N_3721,N_4935);
or U9431 (N_9431,N_700,N_4645);
or U9432 (N_9432,N_4444,N_4611);
nand U9433 (N_9433,N_1629,N_2053);
or U9434 (N_9434,N_2113,N_3819);
and U9435 (N_9435,N_151,N_535);
and U9436 (N_9436,N_3776,N_1774);
and U9437 (N_9437,N_2482,N_3392);
nand U9438 (N_9438,N_2724,N_4916);
and U9439 (N_9439,N_737,N_4604);
nand U9440 (N_9440,N_2673,N_319);
nand U9441 (N_9441,N_324,N_1897);
or U9442 (N_9442,N_3255,N_1386);
or U9443 (N_9443,N_2602,N_487);
nand U9444 (N_9444,N_249,N_4454);
nand U9445 (N_9445,N_4811,N_3090);
or U9446 (N_9446,N_4133,N_3108);
or U9447 (N_9447,N_1612,N_910);
nor U9448 (N_9448,N_3301,N_2455);
or U9449 (N_9449,N_3803,N_3575);
or U9450 (N_9450,N_4392,N_2104);
nor U9451 (N_9451,N_1503,N_3823);
or U9452 (N_9452,N_4149,N_3175);
nor U9453 (N_9453,N_3898,N_4346);
and U9454 (N_9454,N_2303,N_1603);
nand U9455 (N_9455,N_4382,N_1115);
and U9456 (N_9456,N_594,N_4337);
and U9457 (N_9457,N_514,N_1080);
nor U9458 (N_9458,N_4784,N_1795);
and U9459 (N_9459,N_3545,N_2422);
or U9460 (N_9460,N_1861,N_1027);
and U9461 (N_9461,N_2801,N_4954);
or U9462 (N_9462,N_4401,N_1335);
and U9463 (N_9463,N_4087,N_2125);
nand U9464 (N_9464,N_59,N_4624);
and U9465 (N_9465,N_4037,N_1308);
or U9466 (N_9466,N_4898,N_1097);
and U9467 (N_9467,N_2863,N_2802);
nand U9468 (N_9468,N_1571,N_4415);
and U9469 (N_9469,N_3412,N_3587);
nor U9470 (N_9470,N_1627,N_4993);
and U9471 (N_9471,N_602,N_2458);
nand U9472 (N_9472,N_299,N_2794);
nor U9473 (N_9473,N_1057,N_492);
and U9474 (N_9474,N_3799,N_2626);
xor U9475 (N_9475,N_4986,N_2976);
or U9476 (N_9476,N_434,N_3910);
and U9477 (N_9477,N_762,N_1351);
and U9478 (N_9478,N_824,N_2068);
and U9479 (N_9479,N_2767,N_4773);
and U9480 (N_9480,N_2517,N_2551);
nand U9481 (N_9481,N_3359,N_20);
and U9482 (N_9482,N_2822,N_3610);
nand U9483 (N_9483,N_4489,N_4637);
nand U9484 (N_9484,N_1523,N_4484);
xor U9485 (N_9485,N_1680,N_834);
and U9486 (N_9486,N_2399,N_2124);
nor U9487 (N_9487,N_4157,N_1908);
nor U9488 (N_9488,N_2206,N_116);
or U9489 (N_9489,N_3863,N_940);
nor U9490 (N_9490,N_4346,N_628);
and U9491 (N_9491,N_3326,N_1551);
and U9492 (N_9492,N_1011,N_3261);
and U9493 (N_9493,N_2879,N_238);
or U9494 (N_9494,N_4910,N_98);
nand U9495 (N_9495,N_1859,N_1233);
and U9496 (N_9496,N_3632,N_2210);
nand U9497 (N_9497,N_2878,N_1847);
nor U9498 (N_9498,N_1521,N_2878);
and U9499 (N_9499,N_3998,N_4466);
nand U9500 (N_9500,N_4058,N_613);
and U9501 (N_9501,N_2569,N_827);
or U9502 (N_9502,N_4148,N_3306);
and U9503 (N_9503,N_4947,N_3731);
xnor U9504 (N_9504,N_2807,N_2093);
nor U9505 (N_9505,N_2338,N_4973);
and U9506 (N_9506,N_977,N_4655);
and U9507 (N_9507,N_98,N_3995);
nor U9508 (N_9508,N_832,N_734);
nor U9509 (N_9509,N_2860,N_3181);
nor U9510 (N_9510,N_4896,N_4834);
or U9511 (N_9511,N_4285,N_462);
and U9512 (N_9512,N_3395,N_2740);
nor U9513 (N_9513,N_1443,N_1080);
nor U9514 (N_9514,N_3328,N_3577);
nand U9515 (N_9515,N_1963,N_150);
nand U9516 (N_9516,N_1208,N_2131);
and U9517 (N_9517,N_581,N_2904);
nand U9518 (N_9518,N_3592,N_3770);
nand U9519 (N_9519,N_4148,N_3802);
or U9520 (N_9520,N_224,N_3756);
or U9521 (N_9521,N_2752,N_2008);
nand U9522 (N_9522,N_2859,N_2244);
and U9523 (N_9523,N_2969,N_750);
and U9524 (N_9524,N_3137,N_1107);
or U9525 (N_9525,N_3912,N_1764);
or U9526 (N_9526,N_185,N_2981);
and U9527 (N_9527,N_2852,N_1657);
nor U9528 (N_9528,N_2100,N_4620);
nor U9529 (N_9529,N_2489,N_2875);
nor U9530 (N_9530,N_4399,N_2606);
or U9531 (N_9531,N_554,N_3570);
nor U9532 (N_9532,N_3455,N_919);
nand U9533 (N_9533,N_111,N_1132);
or U9534 (N_9534,N_2217,N_722);
and U9535 (N_9535,N_1089,N_643);
and U9536 (N_9536,N_1927,N_2274);
nand U9537 (N_9537,N_844,N_1076);
nand U9538 (N_9538,N_3313,N_3396);
nor U9539 (N_9539,N_4113,N_4510);
and U9540 (N_9540,N_3254,N_3377);
nand U9541 (N_9541,N_3176,N_2114);
and U9542 (N_9542,N_2652,N_4314);
or U9543 (N_9543,N_4564,N_3358);
and U9544 (N_9544,N_2357,N_1354);
or U9545 (N_9545,N_1252,N_3706);
or U9546 (N_9546,N_326,N_1895);
xnor U9547 (N_9547,N_403,N_1524);
or U9548 (N_9548,N_3656,N_1485);
or U9549 (N_9549,N_2810,N_2555);
and U9550 (N_9550,N_3269,N_2701);
and U9551 (N_9551,N_4018,N_3385);
or U9552 (N_9552,N_373,N_4281);
and U9553 (N_9553,N_1718,N_1278);
or U9554 (N_9554,N_280,N_3813);
nand U9555 (N_9555,N_1153,N_4384);
nor U9556 (N_9556,N_2388,N_429);
nand U9557 (N_9557,N_4316,N_1682);
nand U9558 (N_9558,N_4473,N_1024);
and U9559 (N_9559,N_2871,N_4500);
and U9560 (N_9560,N_2912,N_3537);
nand U9561 (N_9561,N_3706,N_16);
nor U9562 (N_9562,N_861,N_2901);
and U9563 (N_9563,N_556,N_1755);
or U9564 (N_9564,N_4249,N_3574);
nand U9565 (N_9565,N_3193,N_925);
or U9566 (N_9566,N_1697,N_1019);
or U9567 (N_9567,N_3879,N_3288);
and U9568 (N_9568,N_2788,N_3113);
and U9569 (N_9569,N_911,N_3764);
nor U9570 (N_9570,N_297,N_4437);
nand U9571 (N_9571,N_301,N_2506);
nor U9572 (N_9572,N_5,N_2743);
nand U9573 (N_9573,N_4501,N_3348);
nand U9574 (N_9574,N_2370,N_251);
nor U9575 (N_9575,N_3977,N_899);
xor U9576 (N_9576,N_1502,N_2891);
nor U9577 (N_9577,N_4433,N_4315);
nor U9578 (N_9578,N_2036,N_1664);
nor U9579 (N_9579,N_4961,N_992);
nand U9580 (N_9580,N_2905,N_3820);
nor U9581 (N_9581,N_4085,N_2490);
nand U9582 (N_9582,N_573,N_2401);
nor U9583 (N_9583,N_356,N_1419);
nor U9584 (N_9584,N_2715,N_3600);
and U9585 (N_9585,N_3415,N_107);
or U9586 (N_9586,N_1521,N_2985);
nor U9587 (N_9587,N_2719,N_3111);
and U9588 (N_9588,N_2482,N_4869);
nor U9589 (N_9589,N_4645,N_2289);
and U9590 (N_9590,N_56,N_217);
and U9591 (N_9591,N_3154,N_3478);
nand U9592 (N_9592,N_1459,N_3362);
or U9593 (N_9593,N_2979,N_2580);
and U9594 (N_9594,N_4624,N_3656);
or U9595 (N_9595,N_724,N_356);
and U9596 (N_9596,N_4733,N_1469);
nor U9597 (N_9597,N_1547,N_3292);
or U9598 (N_9598,N_4545,N_3857);
or U9599 (N_9599,N_509,N_2473);
and U9600 (N_9600,N_2798,N_4279);
or U9601 (N_9601,N_3220,N_4361);
and U9602 (N_9602,N_407,N_1377);
and U9603 (N_9603,N_998,N_1709);
nand U9604 (N_9604,N_3143,N_4401);
and U9605 (N_9605,N_4888,N_3225);
nand U9606 (N_9606,N_4399,N_3779);
or U9607 (N_9607,N_543,N_2775);
and U9608 (N_9608,N_750,N_97);
and U9609 (N_9609,N_4511,N_1779);
nand U9610 (N_9610,N_1462,N_656);
nor U9611 (N_9611,N_4679,N_2595);
nand U9612 (N_9612,N_1346,N_1115);
and U9613 (N_9613,N_1520,N_1130);
and U9614 (N_9614,N_3884,N_2736);
nor U9615 (N_9615,N_4026,N_2079);
or U9616 (N_9616,N_4516,N_747);
nor U9617 (N_9617,N_297,N_3302);
and U9618 (N_9618,N_3673,N_4528);
or U9619 (N_9619,N_4998,N_4731);
nand U9620 (N_9620,N_3243,N_1830);
or U9621 (N_9621,N_778,N_2850);
or U9622 (N_9622,N_4006,N_4327);
and U9623 (N_9623,N_4152,N_2545);
nor U9624 (N_9624,N_4752,N_426);
and U9625 (N_9625,N_583,N_2816);
or U9626 (N_9626,N_558,N_1428);
and U9627 (N_9627,N_78,N_3242);
and U9628 (N_9628,N_3390,N_4788);
nor U9629 (N_9629,N_4465,N_2374);
or U9630 (N_9630,N_230,N_1557);
xor U9631 (N_9631,N_3215,N_1684);
nand U9632 (N_9632,N_2448,N_3132);
nor U9633 (N_9633,N_4435,N_4249);
or U9634 (N_9634,N_2405,N_1107);
nor U9635 (N_9635,N_493,N_3264);
or U9636 (N_9636,N_3829,N_1919);
nor U9637 (N_9637,N_37,N_98);
and U9638 (N_9638,N_889,N_4636);
and U9639 (N_9639,N_4326,N_3256);
and U9640 (N_9640,N_2704,N_1305);
and U9641 (N_9641,N_3215,N_2991);
or U9642 (N_9642,N_4953,N_2774);
or U9643 (N_9643,N_2552,N_2203);
nand U9644 (N_9644,N_4212,N_4395);
nand U9645 (N_9645,N_212,N_3625);
nor U9646 (N_9646,N_2860,N_1561);
nor U9647 (N_9647,N_4432,N_3453);
and U9648 (N_9648,N_2566,N_3274);
or U9649 (N_9649,N_3464,N_2343);
nor U9650 (N_9650,N_4851,N_3349);
and U9651 (N_9651,N_3748,N_1120);
nand U9652 (N_9652,N_4572,N_2375);
nand U9653 (N_9653,N_2667,N_2395);
or U9654 (N_9654,N_985,N_4851);
and U9655 (N_9655,N_1723,N_314);
and U9656 (N_9656,N_4031,N_7);
nand U9657 (N_9657,N_4858,N_3203);
nand U9658 (N_9658,N_2810,N_820);
nor U9659 (N_9659,N_4795,N_2320);
nand U9660 (N_9660,N_610,N_1526);
nand U9661 (N_9661,N_2295,N_1544);
and U9662 (N_9662,N_3052,N_1620);
nand U9663 (N_9663,N_680,N_1436);
and U9664 (N_9664,N_4972,N_416);
and U9665 (N_9665,N_2634,N_635);
and U9666 (N_9666,N_3083,N_4105);
or U9667 (N_9667,N_3204,N_3262);
nor U9668 (N_9668,N_2495,N_3009);
or U9669 (N_9669,N_571,N_4718);
nand U9670 (N_9670,N_1930,N_3317);
or U9671 (N_9671,N_380,N_168);
nand U9672 (N_9672,N_3908,N_3771);
nand U9673 (N_9673,N_4167,N_767);
nand U9674 (N_9674,N_901,N_886);
or U9675 (N_9675,N_1658,N_925);
or U9676 (N_9676,N_2013,N_2320);
nand U9677 (N_9677,N_4461,N_3548);
nor U9678 (N_9678,N_550,N_2520);
and U9679 (N_9679,N_1418,N_3925);
nor U9680 (N_9680,N_289,N_4706);
and U9681 (N_9681,N_479,N_4896);
and U9682 (N_9682,N_80,N_1508);
nand U9683 (N_9683,N_4184,N_4866);
and U9684 (N_9684,N_1732,N_2877);
or U9685 (N_9685,N_1479,N_757);
nor U9686 (N_9686,N_4096,N_1499);
nand U9687 (N_9687,N_3224,N_1939);
nand U9688 (N_9688,N_2945,N_3332);
nor U9689 (N_9689,N_3281,N_4444);
and U9690 (N_9690,N_1372,N_9);
or U9691 (N_9691,N_692,N_560);
and U9692 (N_9692,N_4998,N_1475);
and U9693 (N_9693,N_3685,N_3356);
and U9694 (N_9694,N_393,N_4567);
or U9695 (N_9695,N_3786,N_1221);
nor U9696 (N_9696,N_1310,N_2696);
nand U9697 (N_9697,N_2153,N_2231);
nand U9698 (N_9698,N_907,N_2845);
and U9699 (N_9699,N_2467,N_15);
or U9700 (N_9700,N_4259,N_3004);
and U9701 (N_9701,N_454,N_2634);
or U9702 (N_9702,N_3408,N_1787);
nand U9703 (N_9703,N_4651,N_4404);
xor U9704 (N_9704,N_2045,N_4907);
or U9705 (N_9705,N_917,N_2963);
nand U9706 (N_9706,N_950,N_2398);
or U9707 (N_9707,N_4378,N_3139);
nand U9708 (N_9708,N_758,N_2427);
nand U9709 (N_9709,N_4299,N_1944);
and U9710 (N_9710,N_716,N_2204);
nand U9711 (N_9711,N_4622,N_1579);
or U9712 (N_9712,N_649,N_650);
or U9713 (N_9713,N_4988,N_4787);
and U9714 (N_9714,N_64,N_2390);
or U9715 (N_9715,N_4322,N_4725);
and U9716 (N_9716,N_266,N_2919);
and U9717 (N_9717,N_2125,N_1103);
or U9718 (N_9718,N_2659,N_512);
nor U9719 (N_9719,N_2698,N_2993);
or U9720 (N_9720,N_3883,N_4739);
nor U9721 (N_9721,N_435,N_3460);
nand U9722 (N_9722,N_4773,N_2659);
and U9723 (N_9723,N_203,N_1892);
or U9724 (N_9724,N_2620,N_2884);
or U9725 (N_9725,N_2517,N_4783);
nor U9726 (N_9726,N_4979,N_3886);
or U9727 (N_9727,N_2845,N_2840);
nand U9728 (N_9728,N_1038,N_3702);
nand U9729 (N_9729,N_4797,N_4322);
or U9730 (N_9730,N_734,N_2391);
and U9731 (N_9731,N_3678,N_416);
or U9732 (N_9732,N_2560,N_326);
and U9733 (N_9733,N_2628,N_4688);
or U9734 (N_9734,N_1732,N_3957);
or U9735 (N_9735,N_4317,N_3896);
nand U9736 (N_9736,N_2817,N_2008);
or U9737 (N_9737,N_2714,N_4961);
nand U9738 (N_9738,N_876,N_1639);
or U9739 (N_9739,N_2544,N_3035);
nand U9740 (N_9740,N_1350,N_689);
nand U9741 (N_9741,N_4700,N_1756);
nand U9742 (N_9742,N_4491,N_3342);
nand U9743 (N_9743,N_2816,N_3630);
nor U9744 (N_9744,N_3616,N_2698);
and U9745 (N_9745,N_747,N_4376);
or U9746 (N_9746,N_2394,N_4975);
or U9747 (N_9747,N_2404,N_4404);
nor U9748 (N_9748,N_374,N_4133);
and U9749 (N_9749,N_3556,N_1918);
and U9750 (N_9750,N_876,N_3194);
or U9751 (N_9751,N_688,N_3148);
nand U9752 (N_9752,N_3117,N_720);
nand U9753 (N_9753,N_2634,N_1350);
nor U9754 (N_9754,N_3592,N_4160);
and U9755 (N_9755,N_3335,N_2193);
nor U9756 (N_9756,N_4866,N_291);
xor U9757 (N_9757,N_2079,N_1105);
nand U9758 (N_9758,N_3009,N_2238);
and U9759 (N_9759,N_3605,N_2522);
nor U9760 (N_9760,N_892,N_2276);
nand U9761 (N_9761,N_1710,N_1877);
nor U9762 (N_9762,N_3488,N_54);
and U9763 (N_9763,N_3266,N_413);
or U9764 (N_9764,N_2183,N_1339);
or U9765 (N_9765,N_1498,N_2936);
or U9766 (N_9766,N_2337,N_3960);
nand U9767 (N_9767,N_3846,N_4265);
and U9768 (N_9768,N_1749,N_2910);
or U9769 (N_9769,N_3467,N_2923);
nand U9770 (N_9770,N_900,N_2717);
or U9771 (N_9771,N_4119,N_3791);
nor U9772 (N_9772,N_3150,N_4872);
nor U9773 (N_9773,N_687,N_936);
and U9774 (N_9774,N_1469,N_2603);
or U9775 (N_9775,N_2344,N_1202);
and U9776 (N_9776,N_1759,N_3375);
and U9777 (N_9777,N_4990,N_4792);
nor U9778 (N_9778,N_1590,N_4222);
nand U9779 (N_9779,N_4178,N_2459);
nor U9780 (N_9780,N_2641,N_4647);
or U9781 (N_9781,N_3314,N_358);
or U9782 (N_9782,N_1393,N_1249);
and U9783 (N_9783,N_2440,N_2449);
and U9784 (N_9784,N_4249,N_3203);
nor U9785 (N_9785,N_4849,N_4130);
nor U9786 (N_9786,N_2810,N_1166);
and U9787 (N_9787,N_2436,N_552);
nand U9788 (N_9788,N_1085,N_1608);
nor U9789 (N_9789,N_1179,N_2797);
or U9790 (N_9790,N_594,N_4480);
and U9791 (N_9791,N_534,N_2067);
nor U9792 (N_9792,N_2029,N_2113);
or U9793 (N_9793,N_3063,N_4046);
nor U9794 (N_9794,N_1129,N_1059);
nand U9795 (N_9795,N_3421,N_3486);
nand U9796 (N_9796,N_4014,N_3123);
and U9797 (N_9797,N_4471,N_694);
and U9798 (N_9798,N_2399,N_615);
nand U9799 (N_9799,N_2757,N_1537);
or U9800 (N_9800,N_1381,N_4222);
nand U9801 (N_9801,N_303,N_2781);
nor U9802 (N_9802,N_3695,N_1754);
nor U9803 (N_9803,N_399,N_4766);
nand U9804 (N_9804,N_950,N_4359);
or U9805 (N_9805,N_2827,N_2866);
nor U9806 (N_9806,N_1014,N_676);
or U9807 (N_9807,N_3956,N_4548);
or U9808 (N_9808,N_3563,N_4411);
and U9809 (N_9809,N_4787,N_1046);
or U9810 (N_9810,N_3901,N_319);
nand U9811 (N_9811,N_3091,N_2835);
nand U9812 (N_9812,N_2842,N_3763);
nand U9813 (N_9813,N_3895,N_2230);
nand U9814 (N_9814,N_1494,N_1788);
nand U9815 (N_9815,N_3429,N_983);
nand U9816 (N_9816,N_1046,N_4077);
nor U9817 (N_9817,N_4623,N_159);
or U9818 (N_9818,N_4468,N_1414);
nand U9819 (N_9819,N_2774,N_4843);
nand U9820 (N_9820,N_1418,N_621);
nand U9821 (N_9821,N_3266,N_1420);
or U9822 (N_9822,N_1769,N_200);
nand U9823 (N_9823,N_3044,N_282);
or U9824 (N_9824,N_2477,N_2999);
nor U9825 (N_9825,N_687,N_1568);
nand U9826 (N_9826,N_2233,N_2059);
nor U9827 (N_9827,N_2535,N_2447);
nor U9828 (N_9828,N_1194,N_1112);
nand U9829 (N_9829,N_2871,N_3024);
or U9830 (N_9830,N_1243,N_1910);
nor U9831 (N_9831,N_314,N_3762);
and U9832 (N_9832,N_4851,N_1667);
or U9833 (N_9833,N_2849,N_2579);
nor U9834 (N_9834,N_3025,N_897);
nand U9835 (N_9835,N_1383,N_4378);
and U9836 (N_9836,N_81,N_702);
or U9837 (N_9837,N_4467,N_1752);
nor U9838 (N_9838,N_3608,N_4733);
nor U9839 (N_9839,N_564,N_1407);
or U9840 (N_9840,N_228,N_531);
or U9841 (N_9841,N_1354,N_1977);
and U9842 (N_9842,N_994,N_1397);
nand U9843 (N_9843,N_2859,N_4593);
or U9844 (N_9844,N_4845,N_2365);
nand U9845 (N_9845,N_2076,N_1109);
nor U9846 (N_9846,N_2103,N_1638);
nand U9847 (N_9847,N_741,N_4125);
nor U9848 (N_9848,N_1796,N_1540);
and U9849 (N_9849,N_3951,N_4823);
or U9850 (N_9850,N_4436,N_1287);
or U9851 (N_9851,N_1619,N_1274);
nand U9852 (N_9852,N_3217,N_4408);
nand U9853 (N_9853,N_4926,N_1065);
and U9854 (N_9854,N_2479,N_457);
nand U9855 (N_9855,N_1929,N_1849);
nor U9856 (N_9856,N_995,N_3187);
nand U9857 (N_9857,N_4626,N_4910);
and U9858 (N_9858,N_54,N_1459);
nor U9859 (N_9859,N_4317,N_2800);
nor U9860 (N_9860,N_465,N_4291);
and U9861 (N_9861,N_3157,N_2831);
nand U9862 (N_9862,N_3575,N_3006);
and U9863 (N_9863,N_2145,N_2434);
or U9864 (N_9864,N_1589,N_433);
nand U9865 (N_9865,N_129,N_3804);
nand U9866 (N_9866,N_3620,N_278);
and U9867 (N_9867,N_2066,N_502);
and U9868 (N_9868,N_3203,N_1564);
nor U9869 (N_9869,N_2717,N_3216);
nor U9870 (N_9870,N_4686,N_4613);
or U9871 (N_9871,N_117,N_2557);
or U9872 (N_9872,N_1168,N_107);
or U9873 (N_9873,N_4672,N_4853);
or U9874 (N_9874,N_3677,N_256);
or U9875 (N_9875,N_1408,N_3357);
or U9876 (N_9876,N_183,N_3283);
nand U9877 (N_9877,N_2307,N_3284);
nor U9878 (N_9878,N_30,N_1442);
and U9879 (N_9879,N_4478,N_1452);
or U9880 (N_9880,N_2170,N_4910);
or U9881 (N_9881,N_1061,N_2250);
nor U9882 (N_9882,N_2365,N_4380);
or U9883 (N_9883,N_2985,N_2023);
or U9884 (N_9884,N_1553,N_2977);
nand U9885 (N_9885,N_4968,N_2701);
nand U9886 (N_9886,N_4054,N_2703);
or U9887 (N_9887,N_579,N_1519);
or U9888 (N_9888,N_3879,N_1643);
nor U9889 (N_9889,N_2536,N_8);
and U9890 (N_9890,N_2094,N_0);
nor U9891 (N_9891,N_1132,N_2034);
and U9892 (N_9892,N_3169,N_553);
and U9893 (N_9893,N_4739,N_4326);
or U9894 (N_9894,N_1908,N_1127);
nand U9895 (N_9895,N_3192,N_848);
nor U9896 (N_9896,N_2298,N_1693);
nor U9897 (N_9897,N_3723,N_1222);
nand U9898 (N_9898,N_3589,N_4444);
nand U9899 (N_9899,N_1313,N_63);
nand U9900 (N_9900,N_1340,N_2204);
nor U9901 (N_9901,N_1457,N_2845);
or U9902 (N_9902,N_1283,N_3681);
nand U9903 (N_9903,N_3219,N_2786);
or U9904 (N_9904,N_4322,N_675);
and U9905 (N_9905,N_2736,N_3192);
or U9906 (N_9906,N_1778,N_4138);
nor U9907 (N_9907,N_1181,N_423);
and U9908 (N_9908,N_4797,N_3458);
or U9909 (N_9909,N_4188,N_2886);
nand U9910 (N_9910,N_3478,N_2337);
and U9911 (N_9911,N_4037,N_2719);
or U9912 (N_9912,N_1047,N_3174);
nand U9913 (N_9913,N_3385,N_1586);
and U9914 (N_9914,N_4043,N_1180);
nand U9915 (N_9915,N_1177,N_1426);
nor U9916 (N_9916,N_2245,N_2222);
nor U9917 (N_9917,N_1835,N_3404);
and U9918 (N_9918,N_4414,N_3853);
or U9919 (N_9919,N_750,N_4791);
or U9920 (N_9920,N_2852,N_4313);
nor U9921 (N_9921,N_3392,N_4154);
nor U9922 (N_9922,N_2492,N_1636);
nand U9923 (N_9923,N_3054,N_400);
or U9924 (N_9924,N_3734,N_2535);
nand U9925 (N_9925,N_2662,N_1968);
or U9926 (N_9926,N_3201,N_828);
and U9927 (N_9927,N_2597,N_4734);
nand U9928 (N_9928,N_2148,N_1259);
and U9929 (N_9929,N_4628,N_4551);
and U9930 (N_9930,N_2088,N_899);
and U9931 (N_9931,N_1661,N_1495);
and U9932 (N_9932,N_4700,N_2069);
or U9933 (N_9933,N_1184,N_1851);
nand U9934 (N_9934,N_2443,N_4806);
or U9935 (N_9935,N_3929,N_702);
nand U9936 (N_9936,N_4336,N_3248);
nor U9937 (N_9937,N_4948,N_162);
or U9938 (N_9938,N_50,N_1772);
nor U9939 (N_9939,N_4669,N_2224);
and U9940 (N_9940,N_2829,N_1756);
and U9941 (N_9941,N_3220,N_3071);
or U9942 (N_9942,N_3776,N_1541);
and U9943 (N_9943,N_612,N_1247);
nor U9944 (N_9944,N_1190,N_1086);
and U9945 (N_9945,N_881,N_696);
and U9946 (N_9946,N_2906,N_3576);
and U9947 (N_9947,N_2688,N_4558);
nor U9948 (N_9948,N_2988,N_1492);
and U9949 (N_9949,N_3316,N_3754);
or U9950 (N_9950,N_3083,N_2468);
and U9951 (N_9951,N_3389,N_2560);
nor U9952 (N_9952,N_2351,N_4875);
and U9953 (N_9953,N_148,N_4715);
nor U9954 (N_9954,N_4533,N_2991);
nor U9955 (N_9955,N_2086,N_4567);
or U9956 (N_9956,N_672,N_1309);
or U9957 (N_9957,N_173,N_1299);
nor U9958 (N_9958,N_3708,N_4742);
and U9959 (N_9959,N_1426,N_1079);
or U9960 (N_9960,N_3220,N_954);
nor U9961 (N_9961,N_4672,N_1086);
or U9962 (N_9962,N_3942,N_1369);
nor U9963 (N_9963,N_1706,N_2316);
nor U9964 (N_9964,N_14,N_1114);
and U9965 (N_9965,N_377,N_2275);
nand U9966 (N_9966,N_3802,N_4525);
and U9967 (N_9967,N_1377,N_894);
or U9968 (N_9968,N_3261,N_4469);
or U9969 (N_9969,N_4408,N_2633);
or U9970 (N_9970,N_2559,N_3536);
nand U9971 (N_9971,N_2138,N_3205);
and U9972 (N_9972,N_934,N_2176);
nor U9973 (N_9973,N_2169,N_508);
and U9974 (N_9974,N_4547,N_135);
or U9975 (N_9975,N_3694,N_1773);
nor U9976 (N_9976,N_1312,N_1557);
nand U9977 (N_9977,N_4320,N_565);
and U9978 (N_9978,N_3783,N_3802);
nor U9979 (N_9979,N_2923,N_194);
nor U9980 (N_9980,N_2270,N_4567);
or U9981 (N_9981,N_1516,N_2508);
or U9982 (N_9982,N_2704,N_2564);
and U9983 (N_9983,N_4557,N_4283);
xnor U9984 (N_9984,N_1529,N_1669);
nand U9985 (N_9985,N_4043,N_461);
nand U9986 (N_9986,N_3277,N_29);
nor U9987 (N_9987,N_4076,N_1687);
nor U9988 (N_9988,N_4177,N_2575);
and U9989 (N_9989,N_1437,N_884);
nand U9990 (N_9990,N_25,N_976);
and U9991 (N_9991,N_503,N_3448);
nand U9992 (N_9992,N_4874,N_4473);
nand U9993 (N_9993,N_3255,N_14);
or U9994 (N_9994,N_2262,N_2958);
or U9995 (N_9995,N_2172,N_3542);
or U9996 (N_9996,N_942,N_2721);
and U9997 (N_9997,N_3967,N_4559);
nor U9998 (N_9998,N_2717,N_3256);
nand U9999 (N_9999,N_2508,N_1052);
or U10000 (N_10000,N_6680,N_5309);
or U10001 (N_10001,N_7172,N_8912);
nor U10002 (N_10002,N_9190,N_8980);
nor U10003 (N_10003,N_5353,N_9006);
nor U10004 (N_10004,N_6271,N_8513);
nand U10005 (N_10005,N_7980,N_8807);
nor U10006 (N_10006,N_9521,N_8114);
nand U10007 (N_10007,N_8578,N_8519);
and U10008 (N_10008,N_7804,N_5613);
or U10009 (N_10009,N_6784,N_7679);
and U10010 (N_10010,N_5902,N_6583);
nor U10011 (N_10011,N_9005,N_6515);
nor U10012 (N_10012,N_8023,N_9402);
or U10013 (N_10013,N_5458,N_6207);
nor U10014 (N_10014,N_5924,N_7547);
xnor U10015 (N_10015,N_8010,N_5444);
or U10016 (N_10016,N_6701,N_5857);
and U10017 (N_10017,N_7373,N_6971);
or U10018 (N_10018,N_9291,N_7341);
nand U10019 (N_10019,N_9479,N_5650);
or U10020 (N_10020,N_8693,N_9246);
and U10021 (N_10021,N_9518,N_7195);
or U10022 (N_10022,N_8176,N_8420);
or U10023 (N_10023,N_9222,N_6428);
nor U10024 (N_10024,N_7220,N_5408);
nand U10025 (N_10025,N_8848,N_9644);
and U10026 (N_10026,N_9310,N_8045);
and U10027 (N_10027,N_7561,N_6614);
or U10028 (N_10028,N_7386,N_7984);
or U10029 (N_10029,N_7592,N_9220);
nor U10030 (N_10030,N_7815,N_7872);
xor U10031 (N_10031,N_8988,N_9829);
or U10032 (N_10032,N_5971,N_5319);
nor U10033 (N_10033,N_5139,N_7329);
or U10034 (N_10034,N_6400,N_5637);
nor U10035 (N_10035,N_5615,N_6972);
or U10036 (N_10036,N_7800,N_6490);
and U10037 (N_10037,N_8650,N_8028);
or U10038 (N_10038,N_5571,N_8813);
or U10039 (N_10039,N_6613,N_8091);
and U10040 (N_10040,N_7994,N_8704);
nor U10041 (N_10041,N_5017,N_9027);
and U10042 (N_10042,N_6588,N_5546);
or U10043 (N_10043,N_5523,N_5069);
nand U10044 (N_10044,N_5829,N_8049);
or U10045 (N_10045,N_9195,N_6112);
or U10046 (N_10046,N_5832,N_9556);
nor U10047 (N_10047,N_9315,N_6966);
or U10048 (N_10048,N_9877,N_7781);
or U10049 (N_10049,N_6562,N_6949);
and U10050 (N_10050,N_7265,N_6069);
or U10051 (N_10051,N_9363,N_7462);
and U10052 (N_10052,N_8722,N_7808);
or U10053 (N_10053,N_6557,N_9467);
nand U10054 (N_10054,N_7623,N_5126);
nand U10055 (N_10055,N_6355,N_8262);
nor U10056 (N_10056,N_6965,N_8130);
nand U10057 (N_10057,N_5743,N_9164);
or U10058 (N_10058,N_8349,N_9238);
and U10059 (N_10059,N_9562,N_7945);
and U10060 (N_10060,N_6290,N_9489);
nor U10061 (N_10061,N_7532,N_7059);
or U10062 (N_10062,N_6103,N_8145);
and U10063 (N_10063,N_7423,N_7505);
xnor U10064 (N_10064,N_6461,N_6028);
and U10065 (N_10065,N_9243,N_5778);
or U10066 (N_10066,N_8802,N_8962);
nor U10067 (N_10067,N_9503,N_5675);
nor U10068 (N_10068,N_7251,N_6171);
or U10069 (N_10069,N_5860,N_6174);
nand U10070 (N_10070,N_9616,N_7779);
and U10071 (N_10071,N_6546,N_9380);
nand U10072 (N_10072,N_6994,N_8356);
or U10073 (N_10073,N_7605,N_8221);
nand U10074 (N_10074,N_6002,N_6566);
nand U10075 (N_10075,N_8670,N_9797);
nand U10076 (N_10076,N_7965,N_7014);
nand U10077 (N_10077,N_8332,N_7807);
and U10078 (N_10078,N_5898,N_8089);
and U10079 (N_10079,N_7231,N_7347);
nor U10080 (N_10080,N_6829,N_6740);
and U10081 (N_10081,N_6399,N_9858);
xnor U10082 (N_10082,N_5967,N_8697);
nor U10083 (N_10083,N_8526,N_7687);
and U10084 (N_10084,N_7876,N_6853);
nor U10085 (N_10085,N_6860,N_7069);
nor U10086 (N_10086,N_8799,N_7752);
and U10087 (N_10087,N_8762,N_7333);
and U10088 (N_10088,N_5887,N_8217);
or U10089 (N_10089,N_6045,N_5979);
or U10090 (N_10090,N_9882,N_5375);
nand U10091 (N_10091,N_6033,N_7999);
nand U10092 (N_10092,N_6749,N_6686);
and U10093 (N_10093,N_8795,N_8779);
and U10094 (N_10094,N_6439,N_7413);
nand U10095 (N_10095,N_7543,N_6020);
or U10096 (N_10096,N_7828,N_9016);
nor U10097 (N_10097,N_9376,N_7092);
nor U10098 (N_10098,N_7756,N_9676);
xnor U10099 (N_10099,N_9669,N_5081);
nor U10100 (N_10100,N_6536,N_9811);
nor U10101 (N_10101,N_7272,N_6106);
nand U10102 (N_10102,N_6509,N_6167);
and U10103 (N_10103,N_8470,N_6459);
nor U10104 (N_10104,N_7785,N_9911);
nor U10105 (N_10105,N_9345,N_9841);
nand U10106 (N_10106,N_8075,N_9459);
and U10107 (N_10107,N_5918,N_6506);
or U10108 (N_10108,N_7664,N_7396);
xor U10109 (N_10109,N_9768,N_8445);
nor U10110 (N_10110,N_5032,N_6135);
nand U10111 (N_10111,N_6595,N_6093);
nand U10112 (N_10112,N_9043,N_5271);
and U10113 (N_10113,N_5657,N_8921);
nor U10114 (N_10114,N_5443,N_9427);
nand U10115 (N_10115,N_8721,N_6162);
and U10116 (N_10116,N_7825,N_5321);
and U10117 (N_10117,N_7482,N_8982);
and U10118 (N_10118,N_6296,N_6009);
nor U10119 (N_10119,N_8327,N_5781);
nor U10120 (N_10120,N_7254,N_9286);
or U10121 (N_10121,N_5256,N_5817);
and U10122 (N_10122,N_6465,N_9646);
nor U10123 (N_10123,N_5322,N_8767);
nand U10124 (N_10124,N_8462,N_9872);
or U10125 (N_10125,N_7439,N_7502);
or U10126 (N_10126,N_5407,N_7349);
nor U10127 (N_10127,N_5312,N_9683);
or U10128 (N_10128,N_5378,N_5555);
and U10129 (N_10129,N_6672,N_9274);
or U10130 (N_10130,N_9405,N_6646);
and U10131 (N_10131,N_7319,N_6426);
and U10132 (N_10132,N_5972,N_9808);
or U10133 (N_10133,N_7004,N_7564);
nand U10134 (N_10134,N_5945,N_9952);
nand U10135 (N_10135,N_5264,N_5027);
or U10136 (N_10136,N_9927,N_7754);
nor U10137 (N_10137,N_8699,N_8020);
or U10138 (N_10138,N_7746,N_8371);
or U10139 (N_10139,N_7435,N_6429);
or U10140 (N_10140,N_5262,N_5384);
nor U10141 (N_10141,N_8885,N_6633);
and U10142 (N_10142,N_6513,N_6573);
or U10143 (N_10143,N_5628,N_9301);
and U10144 (N_10144,N_9444,N_8173);
nand U10145 (N_10145,N_5270,N_6435);
nand U10146 (N_10146,N_9697,N_8021);
and U10147 (N_10147,N_7761,N_9745);
nand U10148 (N_10148,N_7879,N_8644);
and U10149 (N_10149,N_9650,N_6607);
or U10150 (N_10150,N_8206,N_7971);
and U10151 (N_10151,N_6144,N_9598);
and U10152 (N_10152,N_6669,N_9638);
or U10153 (N_10153,N_7880,N_9211);
or U10154 (N_10154,N_6525,N_6410);
nor U10155 (N_10155,N_7714,N_7839);
nor U10156 (N_10156,N_8934,N_8450);
and U10157 (N_10157,N_8861,N_5012);
nand U10158 (N_10158,N_5298,N_6064);
nor U10159 (N_10159,N_6365,N_7657);
or U10160 (N_10160,N_8435,N_6305);
or U10161 (N_10161,N_5981,N_6063);
or U10162 (N_10162,N_8576,N_8160);
nand U10163 (N_10163,N_8769,N_8047);
or U10164 (N_10164,N_7010,N_9543);
and U10165 (N_10165,N_5869,N_9523);
nor U10166 (N_10166,N_9559,N_6974);
and U10167 (N_10167,N_5581,N_7404);
nand U10168 (N_10168,N_6511,N_7812);
nor U10169 (N_10169,N_6990,N_7689);
nand U10170 (N_10170,N_5314,N_6988);
nor U10171 (N_10171,N_5789,N_7813);
and U10172 (N_10172,N_7136,N_9773);
or U10173 (N_10173,N_8283,N_8613);
nor U10174 (N_10174,N_6074,N_5761);
nor U10175 (N_10175,N_8355,N_9497);
nor U10176 (N_10176,N_9892,N_8225);
nand U10177 (N_10177,N_9799,N_9864);
or U10178 (N_10178,N_5693,N_6978);
nand U10179 (N_10179,N_9434,N_6370);
and U10180 (N_10180,N_5899,N_7098);
and U10181 (N_10181,N_9487,N_7155);
nand U10182 (N_10182,N_6755,N_6474);
and U10183 (N_10183,N_7629,N_7832);
nor U10184 (N_10184,N_5151,N_9194);
nand U10185 (N_10185,N_7449,N_5195);
nand U10186 (N_10186,N_7944,N_8341);
nor U10187 (N_10187,N_6434,N_6295);
nor U10188 (N_10188,N_5226,N_9072);
nor U10189 (N_10189,N_6552,N_6361);
or U10190 (N_10190,N_5411,N_9404);
and U10191 (N_10191,N_8598,N_6024);
nor U10192 (N_10192,N_6512,N_9140);
and U10193 (N_10193,N_6099,N_7757);
or U10194 (N_10194,N_8106,N_9789);
nor U10195 (N_10195,N_7628,N_9965);
nor U10196 (N_10196,N_6313,N_7217);
nand U10197 (N_10197,N_5459,N_9601);
nand U10198 (N_10198,N_7453,N_9553);
and U10199 (N_10199,N_7022,N_5327);
and U10200 (N_10200,N_7093,N_6431);
nand U10201 (N_10201,N_7916,N_8960);
nand U10202 (N_10202,N_7701,N_9844);
nor U10203 (N_10203,N_7708,N_8455);
and U10204 (N_10204,N_5293,N_9493);
nand U10205 (N_10205,N_7488,N_7478);
and U10206 (N_10206,N_8387,N_7044);
and U10207 (N_10207,N_5995,N_5835);
nand U10208 (N_10208,N_9649,N_8678);
nand U10209 (N_10209,N_5954,N_6161);
and U10210 (N_10210,N_7572,N_8858);
nor U10211 (N_10211,N_6156,N_7335);
or U10212 (N_10212,N_7034,N_5791);
or U10213 (N_10213,N_5597,N_9230);
and U10214 (N_10214,N_6412,N_6420);
or U10215 (N_10215,N_9256,N_6270);
and U10216 (N_10216,N_8417,N_9641);
nor U10217 (N_10217,N_6222,N_9464);
nor U10218 (N_10218,N_7148,N_7552);
nand U10219 (N_10219,N_6341,N_7540);
nand U10220 (N_10220,N_8241,N_8961);
nand U10221 (N_10221,N_7131,N_7745);
and U10222 (N_10222,N_8497,N_8579);
nor U10223 (N_10223,N_5846,N_6141);
nor U10224 (N_10224,N_8529,N_8756);
nor U10225 (N_10225,N_6705,N_5429);
nand U10226 (N_10226,N_9428,N_5395);
and U10227 (N_10227,N_7151,N_5082);
nand U10228 (N_10228,N_8755,N_6991);
and U10229 (N_10229,N_5131,N_9623);
xor U10230 (N_10230,N_7917,N_6837);
and U10231 (N_10231,N_9533,N_9259);
nand U10232 (N_10232,N_7042,N_6952);
nor U10233 (N_10233,N_5323,N_6143);
and U10234 (N_10234,N_6882,N_5457);
xor U10235 (N_10235,N_8062,N_9851);
xor U10236 (N_10236,N_9852,N_8549);
and U10237 (N_10237,N_5341,N_9171);
nand U10238 (N_10238,N_5720,N_6761);
nor U10239 (N_10239,N_8304,N_8302);
or U10240 (N_10240,N_6812,N_9378);
nor U10241 (N_10241,N_8466,N_6010);
and U10242 (N_10242,N_9353,N_6856);
or U10243 (N_10243,N_9282,N_7168);
and U10244 (N_10244,N_6262,N_6387);
nand U10245 (N_10245,N_6501,N_9316);
nor U10246 (N_10246,N_7614,N_8607);
nor U10247 (N_10247,N_7226,N_7078);
nand U10248 (N_10248,N_8984,N_9704);
nand U10249 (N_10249,N_7602,N_6481);
or U10250 (N_10250,N_5683,N_5706);
or U10251 (N_10251,N_6356,N_5472);
nand U10252 (N_10252,N_5794,N_5496);
nor U10253 (N_10253,N_6780,N_8212);
and U10254 (N_10254,N_8015,N_7989);
nor U10255 (N_10255,N_5705,N_7245);
nor U10256 (N_10256,N_5570,N_7143);
nor U10257 (N_10257,N_7273,N_7270);
nor U10258 (N_10258,N_5197,N_7891);
or U10259 (N_10259,N_7608,N_9415);
and U10260 (N_10260,N_6084,N_6922);
or U10261 (N_10261,N_9906,N_7018);
nor U10262 (N_10262,N_9702,N_8600);
or U10263 (N_10263,N_9197,N_6319);
and U10264 (N_10264,N_7787,N_8299);
nand U10265 (N_10265,N_9040,N_8259);
and U10266 (N_10266,N_9870,N_6497);
and U10267 (N_10267,N_9981,N_9805);
nand U10268 (N_10268,N_7823,N_6608);
and U10269 (N_10269,N_5799,N_7416);
nand U10270 (N_10270,N_5281,N_5431);
and U10271 (N_10271,N_5773,N_7621);
nor U10272 (N_10272,N_8643,N_7598);
nand U10273 (N_10273,N_8680,N_9552);
nor U10274 (N_10274,N_5545,N_5218);
nand U10275 (N_10275,N_5834,N_6152);
nor U10276 (N_10276,N_9807,N_9099);
and U10277 (N_10277,N_8994,N_9122);
xnor U10278 (N_10278,N_7674,N_7189);
nor U10279 (N_10279,N_5342,N_6699);
or U10280 (N_10280,N_5109,N_5054);
nor U10281 (N_10281,N_9654,N_5527);
or U10282 (N_10282,N_6508,N_9269);
and U10283 (N_10283,N_6021,N_6560);
and U10284 (N_10284,N_7101,N_9751);
nor U10285 (N_10285,N_5931,N_7321);
nand U10286 (N_10286,N_8750,N_9983);
nand U10287 (N_10287,N_7672,N_8659);
nand U10288 (N_10288,N_7869,N_6752);
nand U10289 (N_10289,N_5075,N_9401);
nand U10290 (N_10290,N_8027,N_8257);
and U10291 (N_10291,N_5369,N_9454);
nand U10292 (N_10292,N_8174,N_5494);
and U10293 (N_10293,N_7244,N_5940);
nand U10294 (N_10294,N_7974,N_8528);
nand U10295 (N_10295,N_7569,N_9723);
nand U10296 (N_10296,N_9390,N_7109);
nor U10297 (N_10297,N_9081,N_6968);
nor U10298 (N_10298,N_5664,N_8451);
and U10299 (N_10299,N_9823,N_6598);
nor U10300 (N_10300,N_9835,N_6083);
or U10301 (N_10301,N_8475,N_9391);
nand U10302 (N_10302,N_9795,N_7499);
nor U10303 (N_10303,N_5007,N_6214);
nand U10304 (N_10304,N_6671,N_6217);
and U10305 (N_10305,N_7514,N_5631);
or U10306 (N_10306,N_7577,N_5721);
and U10307 (N_10307,N_7571,N_5041);
nand U10308 (N_10308,N_9311,N_9137);
nor U10309 (N_10309,N_5452,N_7328);
or U10310 (N_10310,N_9226,N_6424);
or U10311 (N_10311,N_8682,N_8737);
and U10312 (N_10312,N_6788,N_9962);
nand U10313 (N_10313,N_5826,N_5461);
nor U10314 (N_10314,N_5752,N_7356);
nand U10315 (N_10315,N_8998,N_7410);
and U10316 (N_10316,N_9421,N_7052);
nor U10317 (N_10317,N_9532,N_9959);
nor U10318 (N_10318,N_5176,N_9707);
nor U10319 (N_10319,N_8036,N_5175);
nor U10320 (N_10320,N_8515,N_9340);
or U10321 (N_10321,N_8692,N_7904);
or U10322 (N_10322,N_9991,N_8830);
and U10323 (N_10323,N_8163,N_5101);
nor U10324 (N_10324,N_9347,N_6272);
nand U10325 (N_10325,N_8637,N_7892);
nand U10326 (N_10326,N_7312,N_8496);
nor U10327 (N_10327,N_9091,N_8282);
and U10328 (N_10328,N_8149,N_7035);
or U10329 (N_10329,N_9619,N_5646);
nand U10330 (N_10330,N_5167,N_7461);
nor U10331 (N_10331,N_5793,N_8395);
or U10332 (N_10332,N_5166,N_8557);
nand U10333 (N_10333,N_6845,N_8281);
nor U10334 (N_10334,N_9058,N_7649);
or U10335 (N_10335,N_7447,N_8296);
nand U10336 (N_10336,N_5883,N_6872);
nand U10337 (N_10337,N_8118,N_9414);
or U10338 (N_10338,N_9208,N_7243);
nand U10339 (N_10339,N_7730,N_8862);
and U10340 (N_10340,N_9411,N_9847);
nand U10341 (N_10341,N_7282,N_9648);
and U10342 (N_10342,N_9449,N_8425);
nand U10343 (N_10343,N_8922,N_9228);
nand U10344 (N_10344,N_8477,N_6884);
or U10345 (N_10345,N_9838,N_8624);
and U10346 (N_10346,N_7990,N_7769);
nor U10347 (N_10347,N_5292,N_7307);
and U10348 (N_10348,N_9191,N_9097);
and U10349 (N_10349,N_8179,N_7051);
or U10350 (N_10350,N_9344,N_5718);
and U10351 (N_10351,N_5679,N_7591);
nor U10352 (N_10352,N_6995,N_6219);
nor U10353 (N_10353,N_8571,N_6797);
nand U10354 (N_10354,N_8347,N_8824);
or U10355 (N_10355,N_6941,N_9389);
and U10356 (N_10356,N_7337,N_6537);
nand U10357 (N_10357,N_6364,N_7635);
nor U10358 (N_10358,N_7970,N_9678);
nor U10359 (N_10359,N_8316,N_6638);
and U10360 (N_10360,N_8155,N_9519);
and U10361 (N_10361,N_5172,N_6401);
or U10362 (N_10362,N_6180,N_7234);
and U10363 (N_10363,N_7088,N_9033);
nor U10364 (N_10364,N_5225,N_8788);
and U10365 (N_10365,N_9276,N_7859);
nor U10366 (N_10366,N_8431,N_5333);
nor U10367 (N_10367,N_9323,N_8765);
and U10368 (N_10368,N_9944,N_8538);
or U10369 (N_10369,N_8187,N_7384);
nor U10370 (N_10370,N_9100,N_7019);
nand U10371 (N_10371,N_7652,N_6594);
nand U10372 (N_10372,N_9537,N_7176);
nor U10373 (N_10373,N_9742,N_8636);
or U10374 (N_10374,N_9388,N_7766);
nor U10375 (N_10375,N_6229,N_8523);
or U10376 (N_10376,N_6215,N_8907);
nand U10377 (N_10377,N_5142,N_6070);
nand U10378 (N_10378,N_5158,N_9878);
nor U10379 (N_10379,N_5379,N_7773);
and U10380 (N_10380,N_8266,N_5838);
or U10381 (N_10381,N_5801,N_5800);
and U10382 (N_10382,N_8246,N_5662);
or U10383 (N_10383,N_7320,N_6432);
or U10384 (N_10384,N_6667,N_7430);
and U10385 (N_10385,N_5823,N_9869);
xor U10386 (N_10386,N_6902,N_6979);
nand U10387 (N_10387,N_6846,N_9744);
nand U10388 (N_10388,N_6231,N_7500);
nand U10389 (N_10389,N_8310,N_5623);
nand U10390 (N_10390,N_5874,N_9573);
or U10391 (N_10391,N_9051,N_8090);
or U10392 (N_10392,N_9365,N_7894);
nand U10393 (N_10393,N_6661,N_9236);
and U10394 (N_10394,N_6159,N_5134);
and U10395 (N_10395,N_5783,N_5612);
nor U10396 (N_10396,N_5638,N_6418);
or U10397 (N_10397,N_8318,N_8152);
nor U10398 (N_10398,N_8928,N_5576);
and U10399 (N_10399,N_9903,N_5973);
nand U10400 (N_10400,N_8336,N_9472);
and U10401 (N_10401,N_6036,N_5482);
xnor U10402 (N_10402,N_5161,N_8370);
nand U10403 (N_10403,N_6380,N_5814);
nor U10404 (N_10404,N_5518,N_7620);
nor U10405 (N_10405,N_5403,N_6774);
nor U10406 (N_10406,N_9514,N_6538);
nor U10407 (N_10407,N_5450,N_5816);
nand U10408 (N_10408,N_5876,N_7278);
and U10409 (N_10409,N_8000,N_7290);
nand U10410 (N_10410,N_9158,N_8610);
nor U10411 (N_10411,N_5330,N_8007);
nor U10412 (N_10412,N_7986,N_5311);
nand U10413 (N_10413,N_8868,N_6737);
nand U10414 (N_10414,N_7369,N_8674);
nand U10415 (N_10415,N_5553,N_6331);
nor U10416 (N_10416,N_5599,N_6635);
and U10417 (N_10417,N_9127,N_9978);
or U10418 (N_10418,N_7931,N_7852);
nor U10419 (N_10419,N_5632,N_6351);
nor U10420 (N_10420,N_6657,N_5279);
xnor U10421 (N_10421,N_6201,N_7331);
nand U10422 (N_10422,N_6066,N_6321);
nor U10423 (N_10423,N_9067,N_8398);
nand U10424 (N_10424,N_8662,N_7090);
nand U10425 (N_10425,N_8512,N_9827);
and U10426 (N_10426,N_8843,N_8639);
and U10427 (N_10427,N_7512,N_8162);
and U10428 (N_10428,N_6395,N_8172);
nor U10429 (N_10429,N_5456,N_8017);
and U10430 (N_10430,N_5676,N_5241);
nor U10431 (N_10431,N_6483,N_8111);
or U10432 (N_10432,N_9485,N_6281);
or U10433 (N_10433,N_9242,N_7846);
nand U10434 (N_10434,N_6188,N_9592);
xor U10435 (N_10435,N_9071,N_8540);
xnor U10436 (N_10436,N_6891,N_5583);
nand U10437 (N_10437,N_5483,N_8158);
and U10438 (N_10438,N_9342,N_5602);
nor U10439 (N_10439,N_9379,N_5211);
or U10440 (N_10440,N_9156,N_7829);
nor U10441 (N_10441,N_5890,N_7031);
nand U10442 (N_10442,N_8066,N_6170);
nand U10443 (N_10443,N_9212,N_7201);
nor U10444 (N_10444,N_9483,N_5357);
nand U10445 (N_10445,N_5021,N_6254);
or U10446 (N_10446,N_8072,N_9326);
xnor U10447 (N_10447,N_5196,N_5877);
or U10448 (N_10448,N_5694,N_6430);
or U10449 (N_10449,N_6176,N_7465);
nand U10450 (N_10450,N_9661,N_9828);
nor U10451 (N_10451,N_9002,N_8731);
and U10452 (N_10452,N_6119,N_5627);
nand U10453 (N_10453,N_8043,N_6417);
and U10454 (N_10454,N_8418,N_5879);
nor U10455 (N_10455,N_9115,N_8734);
nor U10456 (N_10456,N_9409,N_9207);
and U10457 (N_10457,N_5564,N_9132);
nand U10458 (N_10458,N_8973,N_7676);
or U10459 (N_10459,N_5004,N_8819);
and U10460 (N_10460,N_7023,N_6589);
and U10461 (N_10461,N_9810,N_5715);
and U10462 (N_10462,N_7097,N_7655);
and U10463 (N_10463,N_5941,N_9684);
and U10464 (N_10464,N_6586,N_7075);
nor U10465 (N_10465,N_8073,N_9939);
nand U10466 (N_10466,N_8129,N_8055);
or U10467 (N_10467,N_7383,N_6098);
or U10468 (N_10468,N_9187,N_5290);
nand U10469 (N_10469,N_6443,N_8666);
xnor U10470 (N_10470,N_8429,N_9787);
nor U10471 (N_10471,N_5219,N_5684);
or U10472 (N_10472,N_7299,N_7276);
and U10473 (N_10473,N_9447,N_7469);
and U10474 (N_10474,N_5010,N_5036);
or U10475 (N_10475,N_9740,N_5061);
nand U10476 (N_10476,N_8238,N_8766);
or U10477 (N_10477,N_5359,N_9473);
and U10478 (N_10478,N_6944,N_8042);
and U10479 (N_10479,N_9725,N_5747);
nor U10480 (N_10480,N_6390,N_9551);
nand U10481 (N_10481,N_8743,N_9695);
xnor U10482 (N_10482,N_6023,N_8159);
nand U10483 (N_10483,N_9897,N_5208);
nand U10484 (N_10484,N_7072,N_6245);
or U10485 (N_10485,N_6678,N_6377);
and U10486 (N_10486,N_9266,N_6291);
nor U10487 (N_10487,N_6190,N_8291);
and U10488 (N_10488,N_9701,N_7164);
and U10489 (N_10489,N_7402,N_8877);
or U10490 (N_10490,N_8913,N_5795);
nor U10491 (N_10491,N_9957,N_7388);
nor U10492 (N_10492,N_6772,N_7861);
nand U10493 (N_10493,N_8323,N_5233);
or U10494 (N_10494,N_9622,N_7048);
nor U10495 (N_10495,N_5065,N_9224);
nor U10496 (N_10496,N_6751,N_5467);
or U10497 (N_10497,N_6849,N_6158);
or U10498 (N_10498,N_7011,N_9331);
nor U10499 (N_10499,N_7821,N_5317);
nand U10500 (N_10500,N_6275,N_9923);
nor U10501 (N_10501,N_7029,N_6352);
nor U10502 (N_10502,N_9934,N_7115);
nand U10503 (N_10503,N_8991,N_5119);
or U10504 (N_10504,N_9609,N_5957);
or U10505 (N_10505,N_6411,N_5454);
nand U10506 (N_10506,N_9337,N_8559);
or U10507 (N_10507,N_6577,N_5144);
or U10508 (N_10508,N_9031,N_5983);
nor U10509 (N_10509,N_8153,N_7930);
and U10510 (N_10510,N_7146,N_8237);
or U10511 (N_10511,N_5837,N_5727);
and U10512 (N_10512,N_8248,N_8943);
and U10513 (N_10513,N_6817,N_7125);
nor U10514 (N_10514,N_8683,N_7929);
or U10515 (N_10515,N_9038,N_8113);
nand U10516 (N_10516,N_8353,N_5647);
and U10517 (N_10517,N_7067,N_7489);
nor U10518 (N_10518,N_6842,N_9515);
nand U10519 (N_10519,N_9902,N_7137);
or U10520 (N_10520,N_8761,N_9721);
and U10521 (N_10521,N_7988,N_8537);
and U10522 (N_10522,N_5308,N_8286);
nand U10523 (N_10523,N_5230,N_9364);
nor U10524 (N_10524,N_6526,N_9223);
or U10525 (N_10525,N_6796,N_8718);
xor U10526 (N_10526,N_8889,N_6204);
nor U10527 (N_10527,N_6114,N_7911);
nand U10528 (N_10528,N_8808,N_7332);
and U10529 (N_10529,N_7106,N_8741);
or U10530 (N_10530,N_8927,N_9152);
nor U10531 (N_10531,N_9969,N_9214);
nand U10532 (N_10532,N_7665,N_9203);
or U10533 (N_10533,N_6468,N_7236);
nor U10534 (N_10534,N_8975,N_9972);
and U10535 (N_10535,N_8604,N_6942);
nand U10536 (N_10536,N_8224,N_8953);
and U10537 (N_10537,N_6839,N_9069);
and U10538 (N_10538,N_8071,N_7824);
or U10539 (N_10539,N_9184,N_9946);
nor U10540 (N_10540,N_9780,N_9798);
and U10541 (N_10541,N_8508,N_8285);
nand U10542 (N_10542,N_7962,N_9408);
nor U10543 (N_10543,N_5989,N_7429);
and U10544 (N_10544,N_9997,N_9284);
nor U10545 (N_10545,N_8527,N_7012);
and U10546 (N_10546,N_9831,N_5325);
or U10547 (N_10547,N_9620,N_6149);
nand U10548 (N_10548,N_8256,N_5073);
or U10549 (N_10549,N_5751,N_9087);
and U10550 (N_10550,N_6575,N_9296);
or U10551 (N_10551,N_8204,N_9816);
nand U10552 (N_10552,N_7741,N_5579);
and U10553 (N_10553,N_7798,N_8013);
nor U10554 (N_10554,N_6444,N_5617);
nor U10555 (N_10555,N_5239,N_5433);
and U10556 (N_10556,N_6962,N_5222);
nor U10557 (N_10557,N_8178,N_5260);
nand U10558 (N_10558,N_6825,N_5779);
or U10559 (N_10559,N_7545,N_8433);
nand U10560 (N_10560,N_9568,N_8189);
and U10561 (N_10561,N_9840,N_9445);
nor U10562 (N_10562,N_6031,N_6603);
xnor U10563 (N_10563,N_8702,N_8742);
nor U10564 (N_10564,N_7438,N_8358);
nand U10565 (N_10565,N_9430,N_6854);
nor U10566 (N_10566,N_5034,N_5499);
or U10567 (N_10567,N_6904,N_7968);
nand U10568 (N_10568,N_8979,N_9192);
and U10569 (N_10569,N_8612,N_7267);
nand U10570 (N_10570,N_6736,N_6600);
or U10571 (N_10571,N_6239,N_7100);
nor U10572 (N_10572,N_5393,N_8916);
or U10573 (N_10573,N_5360,N_9018);
or U10574 (N_10574,N_7576,N_7718);
and U10575 (N_10575,N_5700,N_6264);
or U10576 (N_10576,N_8937,N_9586);
and U10577 (N_10577,N_7463,N_7995);
nand U10578 (N_10578,N_6591,N_9716);
and U10579 (N_10579,N_9700,N_9280);
nor U10580 (N_10580,N_8486,N_9837);
and U10581 (N_10581,N_6155,N_9637);
nand U10582 (N_10582,N_9992,N_8040);
nor U10583 (N_10583,N_5993,N_6998);
and U10584 (N_10584,N_9956,N_7574);
and U10585 (N_10585,N_5689,N_7673);
and U10586 (N_10586,N_7353,N_8880);
nand U10587 (N_10587,N_8708,N_7419);
nand U10588 (N_10588,N_8570,N_8597);
nor U10589 (N_10589,N_6259,N_7311);
nor U10590 (N_10590,N_5120,N_9261);
nand U10591 (N_10591,N_5115,N_9596);
and U10592 (N_10592,N_8524,N_6720);
or U10593 (N_10593,N_9086,N_5337);
nor U10594 (N_10594,N_8102,N_7152);
nand U10595 (N_10595,N_7492,N_7959);
or U10596 (N_10596,N_6791,N_8148);
nor U10597 (N_10597,N_9866,N_7996);
or U10598 (N_10598,N_8838,N_9362);
or U10599 (N_10599,N_7856,N_5667);
nand U10600 (N_10600,N_8003,N_7428);
nand U10601 (N_10601,N_5478,N_8669);
and U10602 (N_10602,N_6383,N_7870);
nor U10603 (N_10603,N_7844,N_7070);
and U10604 (N_10604,N_6189,N_6534);
nor U10605 (N_10605,N_8936,N_5100);
nand U10606 (N_10606,N_7433,N_5183);
and U10607 (N_10607,N_5616,N_5373);
nand U10608 (N_10608,N_6531,N_8331);
and U10609 (N_10609,N_6110,N_8501);
or U10610 (N_10610,N_8029,N_6654);
or U10611 (N_10611,N_6168,N_5666);
nand U10612 (N_10612,N_6880,N_7578);
and U10613 (N_10613,N_5372,N_6987);
and U10614 (N_10614,N_6407,N_5808);
nor U10615 (N_10615,N_7440,N_9491);
nand U10616 (N_10616,N_9566,N_6581);
and U10617 (N_10617,N_8125,N_8048);
nand U10618 (N_10618,N_5093,N_8273);
or U10619 (N_10619,N_8931,N_6357);
or U10620 (N_10620,N_5383,N_9988);
nor U10621 (N_10621,N_7056,N_8183);
or U10622 (N_10622,N_9607,N_6206);
and U10623 (N_10623,N_8190,N_7796);
or U10624 (N_10624,N_5284,N_6993);
or U10625 (N_10625,N_6615,N_6279);
and U10626 (N_10626,N_8705,N_8696);
and U10627 (N_10627,N_5641,N_5930);
nand U10628 (N_10628,N_5177,N_9836);
xnor U10629 (N_10629,N_5505,N_6623);
nor U10630 (N_10630,N_6997,N_7113);
nand U10631 (N_10631,N_8458,N_5251);
nor U10632 (N_10632,N_6930,N_7156);
or U10633 (N_10633,N_6675,N_5301);
and U10634 (N_10634,N_9001,N_5604);
and U10635 (N_10635,N_5740,N_9312);
nor U10636 (N_10636,N_9576,N_8312);
nor U10637 (N_10637,N_5697,N_8456);
and U10638 (N_10638,N_5668,N_9657);
nor U10639 (N_10639,N_8530,N_7921);
nor U10640 (N_10640,N_7768,N_5358);
or U10641 (N_10641,N_6234,N_7531);
nor U10642 (N_10642,N_7625,N_8098);
nand U10643 (N_10643,N_5191,N_9169);
nand U10644 (N_10644,N_5228,N_8424);
nor U10645 (N_10645,N_8628,N_9332);
nor U10646 (N_10646,N_9689,N_5964);
nand U10647 (N_10647,N_8865,N_6961);
and U10648 (N_10648,N_8646,N_8097);
and U10649 (N_10649,N_7275,N_8058);
nor U10650 (N_10650,N_8606,N_7841);
or U10651 (N_10651,N_7262,N_7456);
nor U10652 (N_10652,N_9617,N_7127);
nor U10653 (N_10653,N_5210,N_5338);
nor U10654 (N_10654,N_6488,N_8191);
xnor U10655 (N_10655,N_5315,N_7058);
or U10656 (N_10656,N_8236,N_7391);
nor U10657 (N_10657,N_5076,N_6460);
nand U10658 (N_10658,N_9564,N_6054);
nand U10659 (N_10659,N_7316,N_8284);
and U10660 (N_10660,N_9613,N_5371);
or U10661 (N_10661,N_8630,N_5405);
or U10662 (N_10662,N_5394,N_5299);
nor U10663 (N_10663,N_6486,N_9542);
nor U10664 (N_10664,N_6203,N_5376);
nand U10665 (N_10665,N_6674,N_8511);
or U10666 (N_10666,N_8834,N_7471);
nand U10667 (N_10667,N_5749,N_7498);
and U10668 (N_10668,N_8359,N_6900);
or U10669 (N_10669,N_8464,N_6802);
or U10670 (N_10670,N_7733,N_9372);
nand U10671 (N_10671,N_8132,N_6869);
and U10672 (N_10672,N_7960,N_8038);
nor U10673 (N_10673,N_5148,N_7399);
or U10674 (N_10674,N_8277,N_6126);
and U10675 (N_10675,N_7858,N_8269);
nor U10676 (N_10676,N_6362,N_5422);
and U10677 (N_10677,N_8253,N_8245);
nor U10678 (N_10678,N_7723,N_8728);
or U10679 (N_10679,N_5188,N_8825);
and U10680 (N_10680,N_5305,N_9413);
or U10681 (N_10681,N_5095,N_9511);
and U10682 (N_10682,N_9778,N_7782);
and U10683 (N_10683,N_6721,N_6912);
or U10684 (N_10684,N_5432,N_9662);
nand U10685 (N_10685,N_6283,N_6004);
or U10686 (N_10686,N_7436,N_7837);
and U10687 (N_10687,N_6266,N_6068);
and U10688 (N_10688,N_6636,N_6220);
and U10689 (N_10689,N_9821,N_9260);
nand U10690 (N_10690,N_7468,N_9412);
and U10691 (N_10691,N_5901,N_8992);
nand U10692 (N_10692,N_6298,N_7554);
or U10693 (N_10693,N_7950,N_8346);
and U10694 (N_10694,N_5605,N_7103);
or U10695 (N_10695,N_7784,N_9426);
or U10696 (N_10696,N_6241,N_7910);
nor U10697 (N_10697,N_5243,N_8184);
or U10698 (N_10698,N_6344,N_9126);
or U10699 (N_10699,N_8660,N_8276);
and U10700 (N_10700,N_5479,N_9582);
or U10701 (N_10701,N_6933,N_6403);
nand U10702 (N_10702,N_5220,N_5080);
and U10703 (N_10703,N_6195,N_7076);
and U10704 (N_10704,N_8499,N_9201);
nor U10705 (N_10705,N_8397,N_7585);
nor U10706 (N_10706,N_7414,N_7795);
and U10707 (N_10707,N_7339,N_8366);
nand U10708 (N_10708,N_5114,N_7711);
or U10709 (N_10709,N_8590,N_8653);
xnor U10710 (N_10710,N_7642,N_5502);
nor U10711 (N_10711,N_6824,N_6263);
nand U10712 (N_10712,N_5286,N_9106);
nor U10713 (N_10713,N_6905,N_6419);
or U10714 (N_10714,N_9726,N_8782);
nor U10715 (N_10715,N_9814,N_6406);
nand U10716 (N_10716,N_8033,N_8344);
or U10717 (N_10717,N_5488,N_9951);
nand U10718 (N_10718,N_5610,N_9182);
nor U10719 (N_10719,N_7174,N_7024);
nand U10720 (N_10720,N_9819,N_6656);
and U10721 (N_10721,N_8385,N_5880);
nor U10722 (N_10722,N_6601,N_8959);
and U10723 (N_10723,N_7933,N_5624);
nor U10724 (N_10724,N_5003,N_8471);
or U10725 (N_10725,N_8260,N_5848);
or U10726 (N_10726,N_6771,N_6467);
or U10727 (N_10727,N_7160,N_6696);
nor U10728 (N_10728,N_9397,N_8999);
nand U10729 (N_10729,N_7640,N_8541);
nor U10730 (N_10730,N_8474,N_5551);
nor U10731 (N_10731,N_7032,N_6379);
nand U10732 (N_10732,N_7343,N_9728);
nand U10733 (N_10733,N_9004,N_8778);
nor U10734 (N_10734,N_8375,N_9933);
nor U10735 (N_10735,N_6823,N_8093);
and U10736 (N_10736,N_8226,N_5345);
nand U10737 (N_10737,N_5618,N_6857);
or U10738 (N_10738,N_7728,N_9580);
or U10739 (N_10739,N_9967,N_7760);
xor U10740 (N_10740,N_9237,N_8319);
and U10741 (N_10741,N_5854,N_8820);
nor U10742 (N_10742,N_5122,N_5364);
nor U10743 (N_10743,N_9679,N_7406);
or U10744 (N_10744,N_6910,N_7291);
nand U10745 (N_10745,N_5821,N_5803);
and U10746 (N_10746,N_9065,N_5269);
nand U10747 (N_10747,N_5905,N_9949);
nand U10748 (N_10748,N_8100,N_5170);
nor U10749 (N_10749,N_6814,N_8514);
nor U10750 (N_10750,N_7318,N_5283);
nand U10751 (N_10751,N_7184,N_5904);
nand U10752 (N_10752,N_7896,N_5370);
nor U10753 (N_10753,N_6145,N_9677);
nand U10754 (N_10754,N_6062,N_6367);
and U10755 (N_10755,N_9984,N_7736);
nor U10756 (N_10756,N_9890,N_8723);
nor U10757 (N_10757,N_5047,N_6813);
or U10758 (N_10758,N_9541,N_8064);
and U10759 (N_10759,N_9231,N_5129);
and U10760 (N_10760,N_9931,N_5077);
nor U10761 (N_10761,N_5784,N_8574);
nor U10762 (N_10762,N_5366,N_6378);
and U10763 (N_10763,N_7751,N_6007);
and U10764 (N_10764,N_5728,N_9652);
nand U10765 (N_10765,N_8550,N_6042);
nor U10766 (N_10766,N_6628,N_6855);
and U10767 (N_10767,N_7348,N_5229);
or U10768 (N_10768,N_7181,N_7405);
and U10769 (N_10769,N_7675,N_7977);
nand U10770 (N_10770,N_9368,N_7250);
nand U10771 (N_10771,N_9288,N_9561);
nor U10772 (N_10772,N_8725,N_7963);
nor U10773 (N_10773,N_7102,N_5713);
or U10774 (N_10774,N_8196,N_6369);
nand U10775 (N_10775,N_8006,N_8459);
or U10776 (N_10776,N_8416,N_9011);
nor U10777 (N_10777,N_8175,N_8208);
nand U10778 (N_10778,N_7119,N_9971);
nor U10779 (N_10779,N_8635,N_5634);
nor U10780 (N_10780,N_6479,N_8584);
nand U10781 (N_10781,N_5707,N_5636);
nor U10782 (N_10782,N_9741,N_9037);
and U10783 (N_10783,N_5741,N_8383);
nand U10784 (N_10784,N_8985,N_6640);
nand U10785 (N_10785,N_6147,N_7490);
and U10786 (N_10786,N_7246,N_8144);
nand U10787 (N_10787,N_9336,N_8531);
and U10788 (N_10788,N_5040,N_7344);
and U10789 (N_10789,N_9193,N_7095);
nor U10790 (N_10790,N_8580,N_8230);
or U10791 (N_10791,N_9452,N_6695);
xor U10792 (N_10792,N_5424,N_8789);
nand U10793 (N_10793,N_7134,N_9642);
or U10794 (N_10794,N_8641,N_5258);
or U10795 (N_10795,N_5221,N_5831);
and U10796 (N_10796,N_9830,N_6746);
nor U10797 (N_10797,N_7533,N_7460);
xnor U10798 (N_10798,N_7871,N_7283);
xnor U10799 (N_10799,N_6647,N_6127);
nor U10800 (N_10800,N_8078,N_7289);
nand U10801 (N_10801,N_8135,N_8167);
and U10802 (N_10802,N_7124,N_6394);
nand U10803 (N_10803,N_8303,N_6087);
or U10804 (N_10804,N_9756,N_5030);
nor U10805 (N_10805,N_8354,N_8768);
xor U10806 (N_10806,N_6967,N_6252);
and U10807 (N_10807,N_9356,N_7706);
or U10808 (N_10808,N_6392,N_7802);
nor U10809 (N_10809,N_7130,N_8083);
and U10810 (N_10810,N_7229,N_5427);
nand U10811 (N_10811,N_5714,N_6197);
and U10812 (N_10812,N_7953,N_5691);
and U10813 (N_10813,N_5756,N_9073);
or U10814 (N_10814,N_7755,N_9501);
nand U10815 (N_10815,N_8522,N_9149);
nor U10816 (N_10816,N_6287,N_9254);
and U10817 (N_10817,N_5089,N_8556);
xnor U10818 (N_10818,N_8770,N_9539);
nor U10819 (N_10819,N_8258,N_8904);
nand U10820 (N_10820,N_8809,N_6945);
nor U10821 (N_10821,N_5192,N_5549);
or U10822 (N_10822,N_9887,N_6484);
or U10823 (N_10823,N_9633,N_9857);
or U10824 (N_10824,N_5285,N_7759);
nand U10825 (N_10825,N_8565,N_5897);
nand U10826 (N_10826,N_5884,N_9535);
or U10827 (N_10827,N_5303,N_5023);
nand U10828 (N_10828,N_9163,N_5173);
or U10829 (N_10829,N_8009,N_8428);
nor U10830 (N_10830,N_8532,N_8810);
or U10831 (N_10831,N_8521,N_5155);
nor U10832 (N_10832,N_6117,N_5417);
nand U10833 (N_10833,N_9024,N_7973);
nand U10834 (N_10834,N_5392,N_8415);
nand U10835 (N_10835,N_5547,N_6694);
and U10836 (N_10836,N_8828,N_6704);
nor U10837 (N_10837,N_9109,N_5839);
nor U10838 (N_10838,N_8430,N_6086);
or U10839 (N_10839,N_9039,N_9893);
and U10840 (N_10840,N_7816,N_8272);
xnor U10841 (N_10841,N_5094,N_7688);
nand U10842 (N_10842,N_5926,N_5765);
and U10843 (N_10843,N_5060,N_6323);
nor U10844 (N_10844,N_6801,N_7426);
and U10845 (N_10845,N_6150,N_9287);
and U10846 (N_10846,N_7789,N_9225);
and U10847 (N_10847,N_9277,N_8494);
nor U10848 (N_10848,N_9423,N_7323);
and U10849 (N_10849,N_9177,N_8667);
nor U10850 (N_10850,N_9818,N_7288);
nor U10851 (N_10851,N_6702,N_5377);
nor U10852 (N_10852,N_9019,N_8544);
nand U10853 (N_10853,N_9666,N_5858);
and U10854 (N_10854,N_5187,N_9796);
nor U10855 (N_10855,N_8181,N_8891);
nand U10856 (N_10856,N_7099,N_7707);
nor U10857 (N_10857,N_5949,N_8517);
and U10858 (N_10858,N_9842,N_5015);
or U10859 (N_10859,N_6946,N_6652);
nand U10860 (N_10860,N_6533,N_8625);
or U10861 (N_10861,N_7351,N_8067);
and U10862 (N_10862,N_5244,N_9791);
and U10863 (N_10863,N_7644,N_8806);
and U10864 (N_10864,N_7515,N_5272);
or U10865 (N_10865,N_8432,N_5385);
and U10866 (N_10866,N_8855,N_8896);
nand U10867 (N_10867,N_8616,N_8804);
or U10868 (N_10868,N_5753,N_7864);
and U10869 (N_10869,N_5595,N_8698);
and U10870 (N_10870,N_8651,N_5820);
nor U10871 (N_10871,N_8974,N_5398);
nor U10872 (N_10872,N_8603,N_7987);
or U10873 (N_10873,N_7432,N_9021);
or U10874 (N_10874,N_8568,N_9585);
nand U10875 (N_10875,N_8817,N_5157);
or U10876 (N_10876,N_6157,N_9753);
or U10877 (N_10877,N_8647,N_6725);
or U10878 (N_10878,N_6210,N_9671);
nor U10879 (N_10879,N_9198,N_6832);
or U10880 (N_10880,N_7497,N_9131);
nand U10881 (N_10881,N_7803,N_8773);
and U10882 (N_10882,N_7269,N_9699);
nor U10883 (N_10883,N_6726,N_5859);
and U10884 (N_10884,N_9252,N_8965);
and U10885 (N_10885,N_7293,N_9730);
and U10886 (N_10886,N_9891,N_8157);
and U10887 (N_10887,N_7593,N_6447);
nor U10888 (N_10888,N_6992,N_7918);
nor U10889 (N_10889,N_7992,N_5160);
nand U10890 (N_10890,N_9658,N_6804);
nor U10891 (N_10891,N_9327,N_5535);
and U10892 (N_10892,N_8661,N_9801);
nand U10893 (N_10893,N_5343,N_8878);
and U10894 (N_10894,N_8293,N_8631);
and U10895 (N_10895,N_7317,N_9690);
and U10896 (N_10896,N_6113,N_9507);
nor U10897 (N_10897,N_6999,N_6182);
and U10898 (N_10898,N_5106,N_8957);
or U10899 (N_10899,N_5209,N_7313);
nand U10900 (N_10900,N_6469,N_5111);
and U10901 (N_10901,N_8869,N_5538);
nor U10902 (N_10902,N_8169,N_6255);
and U10903 (N_10903,N_5236,N_7354);
nand U10904 (N_10904,N_7441,N_8730);
or U10905 (N_10905,N_6019,N_7065);
xor U10906 (N_10906,N_5600,N_8059);
nand U10907 (N_10907,N_9711,N_6037);
nor U10908 (N_10908,N_9628,N_7470);
or U10909 (N_10909,N_5438,N_9527);
nor U10910 (N_10910,N_6897,N_7955);
or U10911 (N_10911,N_5639,N_7636);
nor U10912 (N_10912,N_8300,N_5214);
and U10913 (N_10913,N_8648,N_5204);
or U10914 (N_10914,N_9680,N_5585);
or U10915 (N_10915,N_8287,N_8271);
or U10916 (N_10916,N_8933,N_6013);
or U10917 (N_10917,N_8909,N_7848);
nor U10918 (N_10918,N_7527,N_8234);
nand U10919 (N_10919,N_5696,N_8037);
or U10920 (N_10920,N_7908,N_6133);
and U10921 (N_10921,N_5868,N_7626);
or U10922 (N_10922,N_9724,N_5936);
and U10923 (N_10923,N_8542,N_9111);
nand U10924 (N_10924,N_6913,N_9781);
nor U10925 (N_10925,N_7163,N_5153);
nor U10926 (N_10926,N_5217,N_9834);
and U10927 (N_10927,N_8056,N_6690);
and U10928 (N_10928,N_7612,N_9525);
nand U10929 (N_10929,N_8746,N_8449);
nor U10930 (N_10930,N_9270,N_9880);
nor U10931 (N_10931,N_6359,N_9929);
and U10932 (N_10932,N_6914,N_7411);
nand U10933 (N_10933,N_8195,N_5288);
and U10934 (N_10934,N_7266,N_8853);
and U10935 (N_10935,N_8239,N_6888);
and U10936 (N_10936,N_8314,N_6895);
or U10937 (N_10937,N_9350,N_6984);
xor U10938 (N_10938,N_6519,N_8533);
nor U10939 (N_10939,N_5557,N_5038);
or U10940 (N_10940,N_6915,N_5988);
nor U10941 (N_10941,N_9257,N_5997);
and U10942 (N_10942,N_5382,N_6520);
and U10943 (N_10943,N_5917,N_8011);
or U10944 (N_10944,N_7669,N_7511);
nor U10945 (N_10945,N_9121,N_8490);
and U10946 (N_10946,N_5762,N_9070);
nand U10947 (N_10947,N_7216,N_9440);
and U10948 (N_10948,N_9715,N_7685);
nand U10949 (N_10949,N_5086,N_6485);
nor U10950 (N_10950,N_9921,N_5416);
nor U10951 (N_10951,N_6228,N_9456);
or U10952 (N_10952,N_8796,N_8847);
and U10953 (N_10953,N_9839,N_7671);
nand U10954 (N_10954,N_5181,N_7057);
or U10955 (N_10955,N_8852,N_5909);
nor U10956 (N_10956,N_7595,N_8495);
and U10957 (N_10957,N_9324,N_6368);
or U10958 (N_10958,N_8235,N_9524);
nor U10959 (N_10959,N_6811,N_6717);
xor U10960 (N_10960,N_6303,N_8857);
or U10961 (N_10961,N_8822,N_6757);
and U10962 (N_10962,N_9794,N_7927);
nand U10963 (N_10963,N_6790,N_6570);
xnor U10964 (N_10964,N_7020,N_9060);
nand U10965 (N_10965,N_9549,N_9595);
or U10966 (N_10966,N_6136,N_6440);
nand U10967 (N_10967,N_7425,N_9846);
nor U10968 (N_10968,N_8087,N_5661);
and U10969 (N_10969,N_5648,N_6848);
and U10970 (N_10970,N_5815,N_9982);
nor U10971 (N_10971,N_7737,N_6541);
or U10972 (N_10972,N_6558,N_9119);
nand U10973 (N_10973,N_6620,N_7161);
nor U10974 (N_10974,N_9629,N_8774);
or U10975 (N_10975,N_9142,N_6427);
nor U10976 (N_10976,N_8841,N_5528);
nor U10977 (N_10977,N_5586,N_7912);
or U10978 (N_10978,N_8161,N_8860);
or U10979 (N_10979,N_7303,N_5695);
nor U10980 (N_10980,N_5733,N_5116);
and U10981 (N_10981,N_5959,N_9333);
or U10982 (N_10982,N_8076,N_9153);
or U10983 (N_10983,N_5532,N_6216);
nor U10984 (N_10984,N_7338,N_6218);
nand U10985 (N_10985,N_7535,N_6125);
nor U10986 (N_10986,N_7091,N_8448);
or U10987 (N_10987,N_7631,N_8695);
and U10988 (N_10988,N_8888,N_7372);
nor U10989 (N_10989,N_6561,N_5146);
or U10990 (N_10990,N_6609,N_7696);
nand U10991 (N_10991,N_5764,N_6768);
and U10992 (N_10992,N_6192,N_5529);
and U10993 (N_10993,N_8836,N_8031);
or U10994 (N_10994,N_8338,N_9985);
and U10995 (N_10995,N_9213,N_9775);
and U10996 (N_10996,N_8726,N_6346);
or U10997 (N_10997,N_8070,N_6307);
nand U10998 (N_10998,N_9935,N_6448);
and U10999 (N_10999,N_6970,N_7393);
nor U11000 (N_11000,N_6051,N_8468);
nand U11001 (N_11001,N_5651,N_6890);
and U11002 (N_11002,N_5991,N_8454);
nand U11003 (N_11003,N_6350,N_7104);
nand U11004 (N_11004,N_6936,N_5223);
nand U11005 (N_11005,N_8617,N_9516);
and U11006 (N_11006,N_6977,N_6003);
or U11007 (N_11007,N_9014,N_6666);
nor U11008 (N_11008,N_6396,N_9560);
and U11009 (N_11009,N_6008,N_7528);
nand U11010 (N_11010,N_7510,N_8082);
xor U11011 (N_11011,N_9612,N_6080);
nor U11012 (N_11012,N_9748,N_5026);
and U11013 (N_11013,N_5594,N_5464);
or U11014 (N_11014,N_8566,N_9078);
or U11015 (N_11015,N_9167,N_9554);
nor U11016 (N_11016,N_9322,N_6238);
or U11017 (N_11017,N_6748,N_6901);
nor U11018 (N_11018,N_7363,N_7094);
nor U11019 (N_11019,N_5351,N_7210);
nand U11020 (N_11020,N_7053,N_5575);
and U11021 (N_11021,N_6826,N_5052);
nor U11022 (N_11022,N_7898,N_5087);
and U11023 (N_11023,N_8360,N_7681);
nand U11024 (N_11024,N_5952,N_8452);
xor U11025 (N_11025,N_9278,N_8703);
nand U11026 (N_11026,N_9719,N_9602);
or U11027 (N_11027,N_9107,N_9804);
nor U11028 (N_11028,N_5182,N_9186);
and U11029 (N_11029,N_7073,N_6115);
nor U11030 (N_11030,N_9367,N_5827);
nor U11031 (N_11031,N_5231,N_6599);
nand U11032 (N_11032,N_8546,N_6756);
and U11033 (N_11033,N_6276,N_5572);
nor U11034 (N_11034,N_5103,N_5324);
and U11035 (N_11035,N_8754,N_8663);
and U11036 (N_11036,N_7740,N_5865);
nor U11037 (N_11037,N_6956,N_9597);
nand U11038 (N_11038,N_5414,N_8792);
or U11039 (N_11039,N_7982,N_8390);
nand U11040 (N_11040,N_6937,N_6921);
nand U11041 (N_11041,N_7190,N_7597);
and U11042 (N_11042,N_7464,N_8791);
or U11043 (N_11043,N_9166,N_9868);
or U11044 (N_11044,N_5259,N_6665);
and U11045 (N_11045,N_5071,N_7778);
or U11046 (N_11046,N_8164,N_8599);
or U11047 (N_11047,N_7427,N_5310);
or U11048 (N_11048,N_5152,N_8052);
nand U11049 (N_11049,N_7187,N_7764);
nor U11050 (N_11050,N_5966,N_8294);
or U11051 (N_11051,N_8301,N_6191);
and U11052 (N_11052,N_6026,N_8199);
or U11053 (N_11053,N_5044,N_5133);
and U11054 (N_11054,N_6315,N_9651);
nand U11055 (N_11055,N_6374,N_7114);
and U11056 (N_11056,N_5025,N_7583);
and U11057 (N_11057,N_5185,N_7909);
nand U11058 (N_11058,N_7882,N_6522);
nand U11059 (N_11059,N_7412,N_8315);
or U11060 (N_11060,N_8560,N_7225);
or U11061 (N_11061,N_7797,N_9922);
or U11062 (N_11062,N_8827,N_6810);
nand U11063 (N_11063,N_6934,N_6981);
and U11064 (N_11064,N_5609,N_9904);
nor U11065 (N_11065,N_9540,N_7506);
and U11066 (N_11066,N_9438,N_7638);
and U11067 (N_11067,N_7817,N_9659);
nor U11068 (N_11068,N_5190,N_8480);
nand U11069 (N_11069,N_8681,N_9486);
and U11070 (N_11070,N_9484,N_6327);
nand U11071 (N_11071,N_8688,N_8409);
nand U11072 (N_11072,N_6879,N_5486);
nor U11073 (N_11073,N_9495,N_6451);
and U11074 (N_11074,N_7036,N_5818);
and U11075 (N_11075,N_5888,N_6932);
nand U11076 (N_11076,N_9199,N_9268);
nand U11077 (N_11077,N_5712,N_8060);
and U11078 (N_11078,N_8112,N_7009);
nand U11079 (N_11079,N_7523,N_7637);
or U11080 (N_11080,N_6187,N_7336);
or U11081 (N_11081,N_9029,N_6556);
or U11082 (N_11082,N_9663,N_8487);
nand U11083 (N_11083,N_8290,N_6258);
nor U11084 (N_11084,N_9581,N_6408);
nor U11085 (N_11085,N_8041,N_5982);
or U11086 (N_11086,N_9615,N_6571);
or U11087 (N_11087,N_7483,N_5560);
nand U11088 (N_11088,N_8733,N_7334);
or U11089 (N_11089,N_6107,N_5083);
nand U11090 (N_11090,N_6122,N_5881);
and U11091 (N_11091,N_8744,N_6294);
and U11092 (N_11092,N_9545,N_5058);
nor U11093 (N_11093,N_5203,N_9863);
nand U11094 (N_11094,N_5462,N_7271);
nand U11095 (N_11095,N_9656,N_5234);
and U11096 (N_11096,N_7952,N_8214);
nand U11097 (N_11097,N_6874,N_5029);
nand U11098 (N_11098,N_8611,N_9233);
or U11099 (N_11099,N_9028,N_8443);
nand U11100 (N_11100,N_6587,N_7487);
and U11101 (N_11101,N_7698,N_8330);
or U11102 (N_11102,N_8990,N_6627);
or U11103 (N_11103,N_6975,N_8168);
xnor U11104 (N_11104,N_7889,N_7767);
nand U11105 (N_11105,N_6183,N_9920);
or U11106 (N_11106,N_8032,N_9134);
and U11107 (N_11107,N_7557,N_8849);
or U11108 (N_11108,N_6293,N_9133);
or U11109 (N_11109,N_7221,N_9432);
and U11110 (N_11110,N_7814,N_6551);
nor U11111 (N_11111,N_7292,N_6078);
or U11112 (N_11112,N_5802,N_7667);
nor U11113 (N_11113,N_6689,N_7919);
nand U11114 (N_11114,N_6101,N_8993);
nor U11115 (N_11115,N_5536,N_8121);
nor U11116 (N_11116,N_6760,N_6631);
and U11117 (N_11117,N_8202,N_6532);
and U11118 (N_11118,N_6416,N_9387);
nor U11119 (N_11119,N_8516,N_5489);
or U11120 (N_11120,N_7525,N_8005);
or U11121 (N_11121,N_5977,N_5336);
nand U11122 (N_11122,N_9318,N_9154);
nand U11123 (N_11123,N_6651,N_6951);
and U11124 (N_11124,N_5716,N_9571);
or U11125 (N_11125,N_9334,N_6859);
and U11126 (N_11126,N_8555,N_6040);
or U11127 (N_11127,N_8902,N_8213);
or U11128 (N_11128,N_7579,N_7401);
and U11129 (N_11129,N_7899,N_6807);
and U11130 (N_11130,N_5550,N_7936);
or U11131 (N_11131,N_6763,N_8709);
nor U11132 (N_11132,N_7129,N_7025);
nor U11133 (N_11133,N_6316,N_7260);
nor U11134 (N_11134,N_5329,N_9961);
or U11135 (N_11135,N_8137,N_9548);
and U11136 (N_11136,N_6065,N_5929);
nand U11137 (N_11137,N_9000,N_5804);
and U11138 (N_11138,N_9047,N_5117);
nand U11139 (N_11139,N_6503,N_9603);
nor U11140 (N_11140,N_5566,N_7107);
or U11141 (N_11141,N_6624,N_6693);
nor U11142 (N_11142,N_8712,N_8897);
nand U11143 (N_11143,N_9088,N_9307);
nor U11144 (N_11144,N_5198,N_7656);
and U11145 (N_11145,N_5630,N_9800);
nor U11146 (N_11146,N_8101,N_6634);
nor U11147 (N_11147,N_6898,N_7326);
nand U11148 (N_11148,N_5893,N_8305);
or U11149 (N_11149,N_7179,N_7403);
or U11150 (N_11150,N_6765,N_8012);
and U11151 (N_11151,N_8536,N_9995);
nor U11152 (N_11152,N_6494,N_6172);
nand U11153 (N_11153,N_8585,N_6286);
nand U11154 (N_11154,N_5542,N_9061);
nor U11155 (N_11155,N_8180,N_8334);
nand U11156 (N_11156,N_5178,N_8664);
nand U11157 (N_11157,N_6871,N_6916);
or U11158 (N_11158,N_9386,N_7310);
or U11159 (N_11159,N_9928,N_6477);
or U11160 (N_11160,N_8919,N_8562);
and U11161 (N_11161,N_7049,N_6148);
and U11162 (N_11162,N_5790,N_7893);
nand U11163 (N_11163,N_8764,N_5480);
or U11164 (N_11164,N_8945,N_6896);
and U11165 (N_11165,N_5517,N_9103);
or U11166 (N_11166,N_8918,N_7788);
nand U11167 (N_11167,N_9853,N_8077);
and U11168 (N_11168,N_8263,N_8222);
nor U11169 (N_11169,N_7061,N_6200);
nand U11170 (N_11170,N_5614,N_5097);
and U11171 (N_11171,N_8182,N_9565);
or U11172 (N_11172,N_9859,N_7584);
nand U11173 (N_11173,N_7417,N_8095);
nor U11174 (N_11174,N_7758,N_7040);
nand U11175 (N_11175,N_5923,N_5278);
and U11176 (N_11176,N_8434,N_5130);
nand U11177 (N_11177,N_6405,N_8220);
and U11178 (N_11178,N_7359,N_8298);
or U11179 (N_11179,N_8786,N_7526);
or U11180 (N_11180,N_7915,N_5912);
nand U11181 (N_11181,N_8640,N_7793);
nand U11182 (N_11182,N_8127,N_6339);
and U11183 (N_11183,N_8881,N_8714);
nand U11184 (N_11184,N_7619,N_5339);
or U11185 (N_11185,N_7081,N_7770);
nand U11186 (N_11186,N_7833,N_9575);
and U11187 (N_11187,N_6502,N_6082);
nand U11188 (N_11188,N_9092,N_5635);
and U11189 (N_11189,N_8684,N_6822);
nor U11190 (N_11190,N_7158,N_6249);
or U11191 (N_11191,N_9588,N_6246);
and U11192 (N_11192,N_6337,N_5938);
nand U11193 (N_11193,N_5849,N_9743);
and U11194 (N_11194,N_5387,N_6292);
or U11195 (N_11195,N_6985,N_6163);
nor U11196 (N_11196,N_6375,N_5235);
and U11197 (N_11197,N_5558,N_8335);
nor U11198 (N_11198,N_9508,N_7609);
nor U11199 (N_11199,N_9113,N_6044);
nand U11200 (N_11200,N_8019,N_8261);
and U11201 (N_11201,N_5987,N_9752);
nand U11202 (N_11202,N_8198,N_8627);
or U11203 (N_11203,N_6782,N_8348);
and U11204 (N_11204,N_6622,N_8794);
or U11205 (N_11205,N_5806,N_6043);
or U11206 (N_11206,N_5734,N_7153);
or U11207 (N_11207,N_6317,N_8069);
and U11208 (N_11208,N_9055,N_5735);
and U11209 (N_11209,N_7791,N_9351);
nand U11210 (N_11210,N_7783,N_8053);
nand U11211 (N_11211,N_7550,N_6179);
and U11212 (N_11212,N_9477,N_5460);
or U11213 (N_11213,N_9494,N_7294);
and U11214 (N_11214,N_6075,N_7519);
and U11215 (N_11215,N_8402,N_5856);
or U11216 (N_11216,N_7838,N_9849);
nor U11217 (N_11217,N_9974,N_6658);
and U11218 (N_11218,N_9970,N_6833);
nor U11219 (N_11219,N_5674,N_9417);
and U11220 (N_11220,N_8201,N_5522);
and U11221 (N_11221,N_7700,N_5937);
and U11222 (N_11222,N_7923,N_8812);
nor U11223 (N_11223,N_6918,N_7682);
nand U11224 (N_11224,N_5328,N_5171);
nor U11225 (N_11225,N_9884,N_5589);
nand U11226 (N_11226,N_7805,N_7182);
nand U11227 (N_11227,N_7135,N_8352);
and U11228 (N_11228,N_9692,N_9820);
or U11229 (N_11229,N_9079,N_8747);
and U11230 (N_11230,N_9765,N_9631);
nand U11231 (N_11231,N_7287,N_6109);
nor U11232 (N_11232,N_5976,N_7806);
or U11233 (N_11233,N_7692,N_9189);
or U11234 (N_11234,N_9915,N_8964);
nor U11235 (N_11235,N_9439,N_9357);
nand U11236 (N_11236,N_5777,N_8309);
or U11237 (N_11237,N_5035,N_8905);
or U11238 (N_11238,N_9112,N_8479);
nand U11239 (N_11239,N_8115,N_6924);
and U11240 (N_11240,N_7001,N_9883);
or U11241 (N_11241,N_6733,N_8870);
and U11242 (N_11242,N_9150,N_9146);
nor U11243 (N_11243,N_5138,N_9833);
and U11244 (N_11244,N_6781,N_7559);
nor U11245 (N_11245,N_9817,N_9299);
nand U11246 (N_11246,N_5099,N_7627);
nor U11247 (N_11247,N_7041,N_6572);
or U11248 (N_11248,N_9241,N_9172);
and U11249 (N_11249,N_7503,N_9110);
nor U11250 (N_11250,N_9098,N_7748);
nand U11251 (N_11251,N_6779,N_7939);
and U11252 (N_11252,N_8966,N_9610);
nand U11253 (N_11253,N_9462,N_9788);
or U11254 (N_11254,N_9674,N_6310);
nor U11255 (N_11255,N_5867,N_7240);
nor U11256 (N_11256,N_8969,N_8340);
nor U11257 (N_11257,N_8126,N_5500);
and U11258 (N_11258,N_5267,N_9672);
and U11259 (N_11259,N_5852,N_7546);
nand U11260 (N_11260,N_5824,N_8882);
and U11261 (N_11261,N_8103,N_6059);
nor U11262 (N_11262,N_7725,N_6793);
or U11263 (N_11263,N_5763,N_5962);
nor U11264 (N_11264,N_6529,N_9298);
and U11265 (N_11265,N_9774,N_5147);
and U11266 (N_11266,N_7166,N_7836);
and U11267 (N_11267,N_6057,N_7196);
xor U11268 (N_11268,N_5677,N_9950);
or U11269 (N_11269,N_5390,N_8609);
and U11270 (N_11270,N_9076,N_9366);
nor U11271 (N_11271,N_6311,N_9036);
and U11272 (N_11272,N_8194,N_5302);
nor U11273 (N_11273,N_5248,N_6792);
nor U11274 (N_11274,N_5782,N_8798);
nor U11275 (N_11275,N_7903,N_5435);
nand U11276 (N_11276,N_7529,N_6224);
or U11277 (N_11277,N_6268,N_6175);
nor U11278 (N_11278,N_5746,N_5018);
and U11279 (N_11279,N_7617,N_6478);
and U11280 (N_11280,N_9856,N_5754);
nor U11281 (N_11281,N_7575,N_8377);
and U11282 (N_11282,N_9032,N_9080);
and U11283 (N_11283,N_9966,N_6492);
and U11284 (N_11284,N_8065,N_7117);
and U11285 (N_11285,N_8485,N_5644);
nor U11286 (N_11286,N_7678,N_6353);
and U11287 (N_11287,N_9210,N_6284);
and U11288 (N_11288,N_5340,N_6329);
and U11289 (N_11289,N_5999,N_6450);
nand U11290 (N_11290,N_5974,N_7877);
or U11291 (N_11291,N_8057,N_7938);
nand U11292 (N_11292,N_8337,N_7914);
and U11293 (N_11293,N_8626,N_9206);
nor U11294 (N_11294,N_9900,N_8586);
or U11295 (N_11295,N_5678,N_8233);
or U11296 (N_11296,N_7937,N_9007);
nor U11297 (N_11297,N_6251,N_5625);
nand U11298 (N_11298,N_6322,N_7030);
xnor U11299 (N_11299,N_8329,N_7253);
nand U11300 (N_11300,N_7518,N_5449);
or U11301 (N_11301,N_6750,N_7476);
nand U11302 (N_11302,N_7096,N_6683);
nor U11303 (N_11303,N_8803,N_8551);
nor U11304 (N_11304,N_5541,N_7205);
nand U11305 (N_11305,N_6619,N_5591);
nor U11306 (N_11306,N_9986,N_7398);
nand U11307 (N_11307,N_6630,N_9375);
nand U11308 (N_11308,N_8324,N_6139);
nor U11309 (N_11309,N_7886,N_9955);
nand U11310 (N_11310,N_6280,N_8655);
or U11311 (N_11311,N_8989,N_9424);
and U11312 (N_11312,N_6366,N_8423);
xnor U11313 (N_11313,N_5442,N_6332);
nor U11314 (N_11314,N_6336,N_7183);
nor U11315 (N_11315,N_8249,N_8080);
nand U11316 (N_11316,N_7633,N_9117);
nand U11317 (N_11317,N_7888,N_5510);
nor U11318 (N_11318,N_8971,N_5184);
nor U11319 (N_11319,N_7780,N_7501);
or U11320 (N_11320,N_6643,N_6097);
and U11321 (N_11321,N_7255,N_7203);
nor U11322 (N_11322,N_8815,N_8935);
nor U11323 (N_11323,N_9673,N_5516);
nand U11324 (N_11324,N_9123,N_8138);
and U11325 (N_11325,N_6053,N_9977);
nand U11326 (N_11326,N_5396,N_7738);
nand U11327 (N_11327,N_7604,N_6085);
and U11328 (N_11328,N_5698,N_9352);
or U11329 (N_11329,N_8592,N_8141);
or U11330 (N_11330,N_5335,N_8510);
and U11331 (N_11331,N_7558,N_9498);
nor U11332 (N_11332,N_6677,N_6659);
and U11333 (N_11333,N_7381,N_8757);
nand U11334 (N_11334,N_5587,N_7279);
or U11335 (N_11335,N_5915,N_8414);
nor U11336 (N_11336,N_6038,N_5475);
and U11337 (N_11337,N_5049,N_6134);
and U11338 (N_11338,N_5404,N_7415);
nand U11339 (N_11339,N_6285,N_8805);
or U11340 (N_11340,N_7123,N_7504);
nor U11341 (N_11341,N_6402,N_5354);
and U11342 (N_11342,N_7455,N_9496);
nor U11343 (N_11343,N_9578,N_6542);
and U11344 (N_11344,N_7901,N_7188);
nand U11345 (N_11345,N_9157,N_7949);
nand U11346 (N_11346,N_7697,N_9873);
nor U11347 (N_11347,N_9587,N_6385);
xor U11348 (N_11348,N_9151,N_9895);
nor U11349 (N_11349,N_8192,N_5836);
or U11350 (N_11350,N_7454,N_6843);
or U11351 (N_11351,N_6470,N_7235);
nand U11352 (N_11352,N_8926,N_5067);
and U11353 (N_11353,N_6703,N_8970);
nor U11354 (N_11354,N_5548,N_5833);
nor U11355 (N_11355,N_5508,N_8972);
or U11356 (N_11356,N_8380,N_5202);
nand U11357 (N_11357,N_7277,N_5078);
or U11358 (N_11358,N_6046,N_7305);
or U11359 (N_11359,N_8133,N_6923);
and U11360 (N_11360,N_6670,N_7368);
nand U11361 (N_11361,N_5554,N_7570);
nand U11362 (N_11362,N_7724,N_7066);
and U11363 (N_11363,N_6095,N_9634);
and U11364 (N_11364,N_8123,N_8170);
nor U11365 (N_11365,N_5519,N_7387);
nor U11366 (N_11366,N_5626,N_9625);
nand U11367 (N_11367,N_5745,N_7530);
nor U11368 (N_11368,N_8108,N_8400);
nand U11369 (N_11369,N_9247,N_8950);
nor U11370 (N_11370,N_6160,N_8632);
or U11371 (N_11371,N_7304,N_6852);
and U11372 (N_11372,N_5611,N_5289);
nand U11373 (N_11373,N_5348,N_9400);
or U11374 (N_11374,N_7855,N_6863);
and U11375 (N_11375,N_6173,N_9441);
or U11376 (N_11376,N_7618,N_9764);
or U11377 (N_11377,N_7539,N_9290);
nor U11378 (N_11378,N_7998,N_8706);
xnor U11379 (N_11379,N_8364,N_8952);
nand U11380 (N_11380,N_9547,N_7956);
and U11381 (N_11381,N_6071,N_8787);
or U11382 (N_11382,N_9176,N_6709);
or U11383 (N_11383,N_6504,N_5622);
nand U11384 (N_11384,N_8379,N_5005);
or U11385 (N_11385,N_6642,N_5163);
or U11386 (N_11386,N_9135,N_6735);
or U11387 (N_11387,N_8854,N_9295);
nand U11388 (N_11388,N_8025,N_5788);
nor U11389 (N_11389,N_8117,N_6983);
and U11390 (N_11390,N_5984,N_6827);
or U11391 (N_11391,N_9567,N_8844);
and U11392 (N_11392,N_5840,N_7315);
or U11393 (N_11393,N_9437,N_6495);
nor U11394 (N_11394,N_6475,N_9855);
or U11395 (N_11395,N_7645,N_5506);
and U11396 (N_11396,N_5079,N_5796);
and U11397 (N_11397,N_6330,N_6809);
nand U11398 (N_11398,N_5162,N_6260);
nand U11399 (N_11399,N_9136,N_8240);
or U11400 (N_11400,N_7357,N_8292);
and U11401 (N_11401,N_9396,N_5574);
xor U11402 (N_11402,N_7831,N_7509);
nor U11403 (N_11403,N_7145,N_8621);
or U11404 (N_11404,N_5711,N_6524);
or U11405 (N_11405,N_7084,N_7776);
and U11406 (N_11406,N_8577,N_5096);
and U11407 (N_11407,N_5563,N_8422);
nand U11408 (N_11408,N_5772,N_6867);
nand U11409 (N_11409,N_7684,N_6948);
or U11410 (N_11410,N_5423,N_9319);
or U11411 (N_11411,N_9647,N_6498);
xnor U11412 (N_11412,N_6012,N_5980);
nand U11413 (N_11413,N_7224,N_9750);
and U11414 (N_11414,N_5135,N_9293);
nand U11415 (N_11415,N_9371,N_8545);
nand U11416 (N_11416,N_7481,N_7774);
nor U11417 (N_11417,N_8906,N_7457);
or U11418 (N_11418,N_5994,N_6545);
and U11419 (N_11419,N_6454,N_5332);
nand U11420 (N_11420,N_5640,N_8658);
nor U11421 (N_11421,N_9235,N_5491);
or U11422 (N_11422,N_7925,N_9052);
nor U11423 (N_11423,N_8061,N_5530);
nand U11424 (N_11424,N_9875,N_7375);
and U11425 (N_11425,N_9733,N_6304);
nand U11426 (N_11426,N_5819,N_5750);
nand U11427 (N_11427,N_5507,N_7739);
nor U11428 (N_11428,N_8136,N_7544);
nand U11429 (N_11429,N_7133,N_5866);
and U11430 (N_11430,N_9786,N_7434);
nand U11431 (N_11431,N_6345,N_9694);
or U11432 (N_11432,N_9862,N_5388);
nand U11433 (N_11433,N_8720,N_9431);
nand U11434 (N_11434,N_6372,N_5780);
nand U11435 (N_11435,N_6724,N_8867);
and U11436 (N_11436,N_8978,N_5537);
nor U11437 (N_11437,N_5056,N_8758);
or U11438 (N_11438,N_9160,N_6058);
nand U11439 (N_11439,N_9914,N_6637);
nand U11440 (N_11440,N_7458,N_9691);
or U11441 (N_11441,N_9359,N_8122);
or U11442 (N_11442,N_7442,N_6653);
or U11443 (N_11443,N_6089,N_7284);
nand U11444 (N_11444,N_9709,N_7258);
nor U11445 (N_11445,N_7370,N_8506);
nand U11446 (N_11446,N_6673,N_7749);
and U11447 (N_11447,N_6253,N_9041);
and U11448 (N_11448,N_6776,N_9305);
or U11449 (N_11449,N_5511,N_5608);
and U11450 (N_11450,N_5642,N_8629);
nor U11451 (N_11451,N_5421,N_9714);
and U11452 (N_11452,N_7340,N_9913);
nand U11453 (N_11453,N_5501,N_6184);
nand U11454 (N_11454,N_6090,N_6205);
or U11455 (N_11455,N_7920,N_6496);
or U11456 (N_11456,N_7801,N_5520);
nand U11457 (N_11457,N_7180,N_5985);
nor U11458 (N_11458,N_7377,N_5265);
or U11459 (N_11459,N_7144,N_8735);
or U11460 (N_11460,N_5512,N_9930);
nor U11461 (N_11461,N_9267,N_5732);
and U11462 (N_11462,N_5921,N_6820);
and U11463 (N_11463,N_8923,N_7281);
and U11464 (N_11464,N_6092,N_7650);
nor U11465 (N_11465,N_9960,N_5582);
or U11466 (N_11466,N_6865,N_8835);
nor U11467 (N_11467,N_9888,N_9450);
and U11468 (N_11468,N_5737,N_8254);
nor U11469 (N_11469,N_5864,N_9802);
nand U11470 (N_11470,N_8963,N_5169);
or U11471 (N_11471,N_8649,N_6516);
nand U11472 (N_11472,N_6816,N_8255);
or U11473 (N_11473,N_5844,N_6129);
or U11474 (N_11474,N_9300,N_6491);
nor U11475 (N_11475,N_5194,N_9180);
xor U11476 (N_11476,N_9958,N_8775);
nand U11477 (N_11477,N_6349,N_8079);
or U11478 (N_11478,N_8339,N_9599);
nor U11479 (N_11479,N_5944,N_6715);
nand U11480 (N_11480,N_6535,N_6527);
or U11481 (N_11481,N_5692,N_6001);
and U11482 (N_11482,N_7424,N_6957);
or U11483 (N_11483,N_8399,N_8267);
nand U11484 (N_11484,N_9746,N_8925);
nor U11485 (N_11485,N_6668,N_8378);
or U11486 (N_11486,N_9793,N_7854);
or U11487 (N_11487,N_9406,N_6660);
nand U11488 (N_11488,N_8563,N_6719);
nor U11489 (N_11489,N_7560,N_6861);
nand U11490 (N_11490,N_8200,N_6716);
nor U11491 (N_11491,N_7966,N_6959);
and U11492 (N_11492,N_8996,N_6456);
or U11493 (N_11493,N_6334,N_6199);
and U11494 (N_11494,N_9499,N_5046);
nand U11495 (N_11495,N_7420,N_9763);
or U11496 (N_11496,N_6306,N_7573);
and U11497 (N_11497,N_7346,N_6213);
and U11498 (N_11498,N_7116,N_9916);
or U11499 (N_11499,N_5766,N_7395);
or U11500 (N_11500,N_9500,N_7228);
or U11501 (N_11501,N_5468,N_7895);
or U11502 (N_11502,N_5380,N_8910);
and U11503 (N_11503,N_9941,N_7691);
nor U11504 (N_11504,N_9717,N_5043);
or U11505 (N_11505,N_6664,N_8831);
and U11506 (N_11506,N_8369,N_7845);
nor U11507 (N_11507,N_6553,N_7060);
nor U11508 (N_11508,N_8552,N_5822);
and U11509 (N_11509,N_9147,N_5397);
or U11510 (N_11510,N_5960,N_5006);
nand U11511 (N_11511,N_5107,N_7632);
nand U11512 (N_11512,N_9458,N_7551);
or U11513 (N_11513,N_7900,N_5347);
or U11514 (N_11514,N_9546,N_9407);
or U11515 (N_11515,N_7843,N_6342);
or U11516 (N_11516,N_9626,N_5598);
nand U11517 (N_11517,N_5247,N_7295);
or U11518 (N_11518,N_6423,N_6834);
nand U11519 (N_11519,N_5619,N_5128);
or U11520 (N_11520,N_5212,N_6954);
nand U11521 (N_11521,N_6835,N_5873);
nor U11522 (N_11522,N_6976,N_6645);
and U11523 (N_11523,N_5419,N_5020);
nor U11524 (N_11524,N_9608,N_5703);
or U11525 (N_11525,N_5870,N_9665);
nor U11526 (N_11526,N_7257,N_7274);
or U11527 (N_11527,N_9976,N_9947);
nor U11528 (N_11528,N_9303,N_7199);
and U11529 (N_11529,N_5320,N_5525);
nand U11530 (N_11530,N_5748,N_6118);
or U11531 (N_11531,N_7407,N_6518);
nor U11532 (N_11532,N_8150,N_5453);
nand U11533 (N_11533,N_9188,N_6393);
nand U11534 (N_11534,N_6409,N_9755);
and U11535 (N_11535,N_5365,N_7450);
and U11536 (N_11536,N_8686,N_5055);
nor U11537 (N_11537,N_7712,N_8361);
or U11538 (N_11538,N_7361,N_9465);
and U11539 (N_11539,N_5900,N_6493);
nor U11540 (N_11540,N_6471,N_7000);
nand U11541 (N_11541,N_7555,N_6014);
nor U11542 (N_11542,N_9482,N_6938);
or U11543 (N_11543,N_6088,N_6441);
nor U11544 (N_11544,N_9258,N_6232);
nor U11545 (N_11545,N_7491,N_9244);
nor U11546 (N_11546,N_9251,N_5282);
xor U11547 (N_11547,N_8981,N_6499);
and U11548 (N_11548,N_8393,N_7418);
nand U11549 (N_11549,N_8492,N_5811);
or U11550 (N_11550,N_8685,N_6326);
and U11551 (N_11551,N_5719,N_7979);
or U11552 (N_11552,N_9583,N_8995);
and U11553 (N_11553,N_7941,N_7197);
nor U11554 (N_11554,N_8759,N_9643);
nor U11555 (N_11555,N_7599,N_8001);
and U11556 (N_11556,N_8177,N_9529);
or U11557 (N_11557,N_9185,N_6862);
nor U11558 (N_11558,N_7750,N_5969);
or U11559 (N_11559,N_7358,N_8223);
and U11560 (N_11560,N_7364,N_9218);
nand U11561 (N_11561,N_9729,N_6789);
nor U11562 (N_11562,N_9738,N_7849);
nor U11563 (N_11563,N_6413,N_7241);
nor U11564 (N_11564,N_5786,N_9713);
nor U11565 (N_11565,N_7634,N_7043);
and U11566 (N_11566,N_6335,N_8924);
and U11567 (N_11567,N_8593,N_8587);
and U11568 (N_11568,N_7790,N_7508);
and U11569 (N_11569,N_9049,N_6382);
or U11570 (N_11570,N_9360,N_8583);
or U11571 (N_11571,N_5402,N_7200);
nand U11572 (N_11572,N_8151,N_6463);
or U11573 (N_11573,N_6505,N_6011);
nand U11574 (N_11574,N_9639,N_5048);
xnor U11575 (N_11575,N_5996,N_5316);
nand U11576 (N_11576,N_9685,N_8050);
nand U11577 (N_11577,N_6104,N_7443);
nor U11578 (N_11578,N_8317,N_7686);
or U11579 (N_11579,N_7452,N_8142);
and U11580 (N_11580,N_9881,N_9614);
nor U11581 (N_11581,N_8748,N_5875);
nand U11582 (N_11582,N_5409,N_8951);
nand U11583 (N_11583,N_7641,N_9074);
nor U11584 (N_11584,N_8345,N_5297);
nand U11585 (N_11585,N_8426,N_6102);
and U11586 (N_11586,N_7459,N_9422);
or U11587 (N_11587,N_5643,N_7873);
nand U11588 (N_11588,N_9645,N_8463);
nand U11589 (N_11589,N_6655,N_6688);
nand U11590 (N_11590,N_7495,N_8401);
nand U11591 (N_11591,N_5349,N_6881);
and U11592 (N_11592,N_5596,N_5361);
nor U11593 (N_11593,N_5584,N_9050);
and U11594 (N_11594,N_9905,N_8736);
nand U11595 (N_11595,N_6743,N_9053);
nand U11596 (N_11596,N_9563,N_7486);
or U11597 (N_11597,N_8654,N_6578);
or U11598 (N_11598,N_5771,N_6940);
and U11599 (N_11599,N_7568,N_6707);
nor U11600 (N_11600,N_5413,N_6828);
and U11601 (N_11601,N_9655,N_9082);
nand U11602 (N_11602,N_6018,N_7567);
or U11603 (N_11603,N_9263,N_8968);
nand U11604 (N_11604,N_8763,N_9766);
or U11605 (N_11605,N_6549,N_8460);
nand U11606 (N_11606,N_6729,N_5885);
xnor U11607 (N_11607,N_8481,N_8413);
nand U11608 (N_11608,N_9273,N_5280);
nand U11609 (N_11609,N_5240,N_9698);
or U11610 (N_11610,N_9272,N_8105);
nand U11611 (N_11611,N_6265,N_8591);
nand U11612 (N_11612,N_6584,N_5729);
or U11613 (N_11613,N_7983,N_7222);
or U11614 (N_11614,N_9118,N_6567);
and U11615 (N_11615,N_7670,N_5473);
nand U11616 (N_11616,N_6489,N_9924);
and U11617 (N_11617,N_5350,N_7957);
nor U11618 (N_11618,N_7021,N_8419);
or U11619 (N_11619,N_9104,N_5118);
or U11620 (N_11620,N_9083,N_8143);
nor U11621 (N_11621,N_6886,N_5592);
nand U11622 (N_11622,N_5889,N_9370);
and U11623 (N_11623,N_8700,N_8491);
or U11624 (N_11624,N_6878,N_6539);
and U11625 (N_11625,N_9784,N_9304);
or U11626 (N_11626,N_5513,N_5274);
or U11627 (N_11627,N_9433,N_9936);
nor U11628 (N_11628,N_6691,N_8209);
and U11629 (N_11629,N_9129,N_7651);
nand U11630 (N_11630,N_9325,N_5701);
and U11631 (N_11631,N_6178,N_6015);
or U11632 (N_11632,N_8436,N_6146);
nor U11633 (N_11633,N_9373,N_5346);
nor U11634 (N_11634,N_7951,N_6876);
nor U11635 (N_11635,N_6373,N_8251);
or U11636 (N_11636,N_8478,N_7743);
nor U11637 (N_11637,N_7851,N_8892);
nand U11638 (N_11638,N_5504,N_7695);
nand U11639 (N_11639,N_7715,N_7475);
nor U11640 (N_11640,N_5051,N_8740);
nor U11641 (N_11641,N_5352,N_5767);
and U11642 (N_11642,N_5965,N_8751);
nand U11643 (N_11643,N_8034,N_8582);
nand U11644 (N_11644,N_5368,N_7374);
nand U11645 (N_11645,N_9179,N_7622);
xor U11646 (N_11646,N_7147,N_9635);
nor U11647 (N_11647,N_9410,N_7132);
and U11648 (N_11648,N_5205,N_5001);
xor U11649 (N_11649,N_6596,N_7392);
nor U11650 (N_11650,N_5687,N_6894);
nor U11651 (N_11651,N_7389,N_6138);
or U11652 (N_11652,N_9317,N_8328);
nand U11653 (N_11653,N_6108,N_6754);
nor U11654 (N_11654,N_5213,N_8833);
nor U11655 (N_11655,N_9806,N_5381);
nor U11656 (N_11656,N_5068,N_6094);
and U11657 (N_11657,N_6982,N_9062);
nor U11658 (N_11658,N_9670,N_6783);
nand U11659 (N_11659,N_7588,N_7702);
and U11660 (N_11660,N_5759,N_8793);
or U11661 (N_11661,N_9918,N_6154);
or U11662 (N_11662,N_5064,N_9161);
nand U11663 (N_11663,N_7365,N_5232);
nand U11664 (N_11664,N_7238,N_8940);
nand U11665 (N_11665,N_8322,N_6464);
or U11666 (N_11666,N_8596,N_8846);
nor U11667 (N_11667,N_6617,N_7142);
nand U11668 (N_11668,N_9461,N_8026);
nor U11669 (N_11669,N_9017,N_8717);
nand U11670 (N_11670,N_5455,N_5412);
and U11671 (N_11671,N_8752,N_8265);
nand U11672 (N_11672,N_9096,N_7594);
nand U11673 (N_11673,N_6208,N_8171);
and U11674 (N_11674,N_5871,N_5355);
nor U11675 (N_11675,N_8800,N_7826);
nor U11676 (N_11676,N_7536,N_5934);
or U11677 (N_11677,N_8535,N_7327);
or U11678 (N_11678,N_7630,N_9809);
or U11679 (N_11679,N_6986,N_7606);
nand U11680 (N_11680,N_5261,N_7958);
or U11681 (N_11681,N_9480,N_5304);
and U11682 (N_11682,N_5809,N_6892);
or U11683 (N_11683,N_9398,N_8215);
nor U11684 (N_11684,N_9403,N_5418);
and U11685 (N_11685,N_6079,N_5658);
and U11686 (N_11686,N_9116,N_6730);
nand U11687 (N_11687,N_5084,N_8453);
or U11688 (N_11688,N_8575,N_6632);
xnor U11689 (N_11689,N_5313,N_5273);
nor U11690 (N_11690,N_9528,N_7350);
nor U11691 (N_11691,N_6067,N_5725);
and U11692 (N_11692,N_6775,N_6787);
nor U11693 (N_11693,N_7693,N_5903);
or U11694 (N_11694,N_6706,N_9510);
nand U11695 (N_11695,N_7362,N_6679);
nand U11696 (N_11696,N_8938,N_6230);
nor U11697 (N_11697,N_8096,N_8367);
and U11698 (N_11698,N_5156,N_5659);
or U11699 (N_11699,N_8362,N_8140);
or U11700 (N_11700,N_6318,N_8895);
or U11701 (N_11701,N_8376,N_9054);
or U11702 (N_11702,N_8941,N_5224);
nor U11703 (N_11703,N_5164,N_8351);
and U11704 (N_11704,N_5249,N_5503);
nand U11705 (N_11705,N_5237,N_5655);
nor U11706 (N_11706,N_8381,N_9066);
or U11707 (N_11707,N_9471,N_7699);
or U11708 (N_11708,N_8110,N_7074);
or U11709 (N_11709,N_9349,N_9718);
and U11710 (N_11710,N_9899,N_6593);
and U11711 (N_11711,N_9355,N_9346);
nor U11712 (N_11712,N_7522,N_9989);
nand U11713 (N_11713,N_5470,N_5108);
nand U11714 (N_11714,N_7639,N_5252);
nand U11715 (N_11715,N_7496,N_8932);
nand U11716 (N_11716,N_8915,N_5374);
or U11717 (N_11717,N_8502,N_8929);
nor U11718 (N_11718,N_9329,N_6047);
and U11719 (N_11719,N_6433,N_6734);
or U11720 (N_11720,N_8389,N_6685);
and U11721 (N_11721,N_5062,N_7466);
nand U11722 (N_11722,N_7493,N_9681);
nor U11723 (N_11723,N_6030,N_9776);
nand U11724 (N_11724,N_7280,N_7378);
nor U11725 (N_11725,N_9954,N_8116);
and U11726 (N_11726,N_8872,N_6885);
or U11727 (N_11727,N_5463,N_5490);
nor U11728 (N_11728,N_5033,N_7159);
nor U11729 (N_11729,N_9557,N_5420);
nand U11730 (N_11730,N_9399,N_8874);
nor U11731 (N_11731,N_9867,N_8675);
or U11732 (N_11732,N_9686,N_5448);
and U11733 (N_11733,N_7232,N_7819);
and U11734 (N_11734,N_6973,N_7380);
and U11735 (N_11735,N_8403,N_7451);
nor U11736 (N_11736,N_6221,N_7792);
nand U11737 (N_11737,N_6909,N_7324);
nand U11738 (N_11738,N_9502,N_9030);
and U11739 (N_11739,N_9942,N_7772);
and U11740 (N_11740,N_6883,N_5024);
or U11741 (N_11741,N_6376,N_9570);
and U11742 (N_11742,N_7268,N_8920);
nor U11743 (N_11743,N_9285,N_7534);
and U11744 (N_11744,N_9003,N_7513);
and U11745 (N_11745,N_9973,N_9077);
and U11746 (N_11746,N_8210,N_9760);
nor U11747 (N_11747,N_5649,N_9783);
or U11748 (N_11748,N_8588,N_7926);
nand U11749 (N_11749,N_7878,N_5645);
nor U11750 (N_11750,N_6032,N_9442);
nor U11751 (N_11751,N_6543,N_5389);
nor U11752 (N_11752,N_7818,N_9341);
and U11753 (N_11753,N_7516,N_9250);
nand U11754 (N_11754,N_9538,N_8785);
nor U11755 (N_11755,N_5892,N_8391);
nor U11756 (N_11756,N_5415,N_9505);
or U11757 (N_11757,N_9885,N_8619);
nor U11758 (N_11758,N_9987,N_8307);
nor U11759 (N_11759,N_8392,N_8890);
or U11760 (N_11760,N_6140,N_6767);
nor U11761 (N_11761,N_8908,N_7446);
and U11762 (N_11762,N_5787,N_7177);
and U11763 (N_11763,N_6844,N_9506);
and U11764 (N_11764,N_9705,N_8716);
nor U11765 (N_11765,N_7863,N_9604);
and U11766 (N_11766,N_5812,N_7193);
nor U11767 (N_11767,N_9975,N_5140);
nor U11768 (N_11768,N_9175,N_9045);
or U11769 (N_11769,N_7538,N_8866);
nor U11770 (N_11770,N_6676,N_9513);
and U11771 (N_11771,N_9898,N_5474);
nor U11772 (N_11772,N_7705,N_6917);
and U11773 (N_11773,N_8205,N_9063);
nor U11774 (N_11774,N_6996,N_8749);
nor U11775 (N_11775,N_8851,N_9343);
and U11776 (N_11776,N_9937,N_9221);
nor U11777 (N_11777,N_6963,N_5724);
or U11778 (N_11778,N_7747,N_5975);
nor U11779 (N_11779,N_8898,N_6482);
or U11780 (N_11780,N_5031,N_7654);
or U11781 (N_11781,N_9239,N_6773);
and U11782 (N_11782,N_9183,N_9630);
nor U11783 (N_11783,N_9860,N_9874);
or U11784 (N_11784,N_8701,N_5088);
xor U11785 (N_11785,N_6592,N_5037);
or U11786 (N_11786,N_8388,N_6723);
and U11787 (N_11787,N_6648,N_5895);
nand U11788 (N_11788,N_6242,N_6457);
and U11789 (N_11789,N_8539,N_8665);
nor U11790 (N_11790,N_5845,N_9013);
xnor U11791 (N_11791,N_7400,N_8671);
and U11792 (N_11792,N_5861,N_8407);
nand U11793 (N_11793,N_9703,N_7355);
xnor U11794 (N_11794,N_6000,N_9504);
nand U11795 (N_11795,N_7479,N_5813);
and U11796 (N_11796,N_9229,N_6142);
nand U11797 (N_11797,N_5465,N_9105);
and U11798 (N_11798,N_6061,N_8467);
nand U11799 (N_11799,N_5606,N_8342);
or U11800 (N_11800,N_8673,N_9308);
nand U11801 (N_11801,N_9420,N_8930);
xor U11802 (N_11802,N_5603,N_9907);
or U11803 (N_11803,N_9302,N_5123);
or U11804 (N_11804,N_5059,N_7118);
nand U11805 (N_11805,N_5206,N_5104);
and U11806 (N_11806,N_9688,N_9383);
and U11807 (N_11807,N_7771,N_9785);
nor U11808 (N_11808,N_8350,N_7121);
nand U11809 (N_11809,N_6186,N_8569);
and U11810 (N_11810,N_6227,N_6731);
or U11811 (N_11811,N_8365,N_6629);
and U11812 (N_11812,N_7985,N_5717);
and U11813 (N_11813,N_6742,N_8288);
nor U11814 (N_11814,N_6663,N_6908);
and U11815 (N_11815,N_7122,N_5947);
or U11816 (N_11816,N_9008,N_9354);
xnor U11817 (N_11817,N_8421,N_6564);
and U11818 (N_11818,N_9125,N_6785);
nand U11819 (N_11819,N_6579,N_8441);
nand U11820 (N_11820,N_5768,N_6302);
nor U11821 (N_11821,N_8022,N_8997);
nand U11822 (N_11822,N_7120,N_9022);
nand U11823 (N_11823,N_5723,N_8197);
nor U11824 (N_11824,N_7002,N_6299);
and U11825 (N_11825,N_7860,N_8051);
and U11826 (N_11826,N_9777,N_8203);
nand U11827 (N_11827,N_9034,N_8457);
and U11828 (N_11828,N_8900,N_5102);
nor U11829 (N_11829,N_6181,N_8227);
or U11830 (N_11830,N_5531,N_8645);
nor U11831 (N_11831,N_8207,N_9606);
nor U11832 (N_11832,N_6687,N_7259);
and U11833 (N_11833,N_9632,N_9227);
nand U11834 (N_11834,N_5653,N_8967);
nand U11835 (N_11835,N_5855,N_9476);
nand U11836 (N_11836,N_7261,N_5710);
nor U11837 (N_11837,N_7542,N_5367);
nor U11838 (N_11838,N_8382,N_6712);
and U11839 (N_11839,N_7212,N_6466);
and U11840 (N_11840,N_9832,N_8185);
or U11841 (N_11841,N_5344,N_6931);
and U11842 (N_11842,N_6831,N_8247);
and U11843 (N_11843,N_8879,N_5113);
nand U11844 (N_11844,N_7192,N_9374);
or U11845 (N_11845,N_5074,N_5428);
nand U11846 (N_11846,N_7223,N_8901);
and U11847 (N_11847,N_5776,N_9457);
or U11848 (N_11848,N_9139,N_5939);
and U11849 (N_11849,N_6875,N_8534);
nor U11850 (N_11850,N_8250,N_5663);
nor U11851 (N_11851,N_7379,N_9443);
nor U11852 (N_11852,N_6514,N_5008);
and U11853 (N_11853,N_8104,N_5186);
xnor U11854 (N_11854,N_8086,N_6989);
nand U11855 (N_11855,N_5590,N_7431);
nand U11856 (N_11856,N_6120,N_8745);
or U11857 (N_11857,N_6764,N_7517);
nor U11858 (N_11858,N_5476,N_6212);
nand U11859 (N_11859,N_9048,N_8165);
or U11860 (N_11860,N_5708,N_8193);
or U11861 (N_11861,N_7264,N_7016);
nor U11862 (N_11862,N_7008,N_9708);
nand U11863 (N_11863,N_8279,N_5922);
or U11864 (N_11864,N_9338,N_8947);
xor U11865 (N_11865,N_7421,N_6698);
nand U11866 (N_11866,N_9124,N_6282);
and U11867 (N_11867,N_9762,N_7422);
nand U11868 (N_11868,N_8894,N_9668);
or U11869 (N_11869,N_6415,N_8955);
and U11870 (N_11870,N_7170,N_5057);
nand U11871 (N_11871,N_7954,N_5179);
nand U11872 (N_11872,N_7082,N_7607);
or U11873 (N_11873,N_7734,N_6209);
nor U11874 (N_11874,N_6035,N_8325);
nand U11875 (N_11875,N_8218,N_8771);
or U11876 (N_11876,N_5709,N_6641);
or U11877 (N_11877,N_9392,N_7840);
and U11878 (N_11878,N_9757,N_7071);
nor U11879 (N_11879,N_5493,N_6903);
nand U11880 (N_11880,N_9255,N_5149);
nand U11881 (N_11881,N_5066,N_7709);
nand U11882 (N_11882,N_6404,N_9416);
nand U11883 (N_11883,N_9178,N_9675);
and U11884 (N_11884,N_7068,N_8219);
and U11885 (N_11885,N_8875,N_8707);
nand U11886 (N_11886,N_5593,N_8605);
nor U11887 (N_11887,N_7661,N_9240);
or U11888 (N_11888,N_6626,N_8760);
nor U11889 (N_11889,N_7230,N_9057);
and U11890 (N_11890,N_7409,N_8690);
nor U11891 (N_11891,N_6682,N_9143);
nor U11892 (N_11892,N_5543,N_7263);
nor U11893 (N_11893,N_9020,N_8739);
and U11894 (N_11894,N_9579,N_5828);
nand U11895 (N_11895,N_6256,N_9385);
nor U11896 (N_11896,N_5673,N_8472);
and U11897 (N_11897,N_9732,N_9056);
or U11898 (N_11898,N_6758,N_9998);
and U11899 (N_11899,N_6517,N_6240);
nor U11900 (N_11900,N_5797,N_7050);
and U11901 (N_11901,N_9824,N_8719);
or U11902 (N_11902,N_8404,N_9384);
nor U11903 (N_11903,N_6700,N_8139);
nor U11904 (N_11904,N_7590,N_5399);
or U11905 (N_11905,N_5002,N_6360);
nor U11906 (N_11906,N_7704,N_9734);
nand U11907 (N_11907,N_9660,N_6132);
and U11908 (N_11908,N_6388,N_8438);
nor U11909 (N_11909,N_7360,N_7437);
nand U11910 (N_11910,N_6325,N_6582);
and U11911 (N_11911,N_7064,N_7352);
and U11912 (N_11912,N_7382,N_8850);
and U11913 (N_11913,N_6277,N_9204);
nor U11914 (N_11914,N_7077,N_9314);
and U11915 (N_11915,N_8504,N_7653);
and U11916 (N_11916,N_8732,N_9009);
or U11917 (N_11917,N_9682,N_6953);
or U11918 (N_11918,N_8829,N_9478);
nand U11919 (N_11919,N_6458,N_6274);
nor U11920 (N_11920,N_7961,N_9593);
and U11921 (N_11921,N_9271,N_9084);
and U11922 (N_11922,N_7033,N_6778);
or U11923 (N_11923,N_9979,N_7596);
or U11924 (N_11924,N_8772,N_6523);
nor U11925 (N_11925,N_9120,N_5843);
nand U11926 (N_11926,N_6662,N_6193);
and U11927 (N_11927,N_5953,N_9429);
nand U11928 (N_11928,N_5019,N_9141);
or U11929 (N_11929,N_5400,N_7298);
nand U11930 (N_11930,N_9640,N_6738);
nor U11931 (N_11931,N_8444,N_6052);
and U11932 (N_11932,N_7850,N_9114);
and U11933 (N_11933,N_6612,N_8498);
nor U11934 (N_11934,N_5287,N_9917);
and U11935 (N_11935,N_7948,N_8797);
and U11936 (N_11936,N_9591,N_9306);
or U11937 (N_11937,N_6198,N_6223);
and U11938 (N_11938,N_9782,N_7905);
nand U11939 (N_11939,N_8814,N_6237);
nor U11940 (N_11940,N_9023,N_9470);
nor U11941 (N_11941,N_8547,N_9618);
nor U11942 (N_11942,N_7325,N_8622);
nor U11943 (N_11943,N_8311,N_7237);
nand U11944 (N_11944,N_6055,N_8525);
or U11945 (N_11945,N_6226,N_5189);
and U11946 (N_11946,N_5275,N_9926);
or U11947 (N_11947,N_7038,N_5670);
nor U11948 (N_11948,N_7658,N_6870);
xor U11949 (N_11949,N_9948,N_6121);
nor U11950 (N_11950,N_9990,N_6500);
or U11951 (N_11951,N_7006,N_5466);
xnor U11952 (N_11952,N_7366,N_9772);
nor U11953 (N_11953,N_8887,N_5484);
and U11954 (N_11954,N_5894,N_9159);
and U11955 (N_11955,N_6510,N_7112);
or U11956 (N_11956,N_7643,N_7603);
nor U11957 (N_11957,N_6384,N_6769);
nand U11958 (N_11958,N_5956,N_8948);
or U11959 (N_11959,N_7028,N_7875);
and U11960 (N_11960,N_6169,N_6550);
or U11961 (N_11961,N_6371,N_5539);
or U11962 (N_11962,N_5842,N_7735);
nor U11963 (N_11963,N_9245,N_6819);
nand U11964 (N_11964,N_6267,N_9908);
and U11965 (N_11965,N_7397,N_5872);
nor U11966 (N_11966,N_8119,N_6196);
or U11967 (N_11967,N_5331,N_8864);
nor U11968 (N_11968,N_9993,N_6250);
nand U11969 (N_11969,N_5447,N_9825);
nand U11970 (N_11970,N_8949,N_8306);
and U11971 (N_11971,N_6697,N_9321);
or U11972 (N_11972,N_6006,N_8956);
nor U11973 (N_11973,N_9530,N_5810);
nor U11974 (N_11974,N_8146,N_5268);
or U11975 (N_11975,N_5200,N_8394);
or U11976 (N_11976,N_9253,N_9200);
or U11977 (N_11977,N_8476,N_9876);
or U11978 (N_11978,N_7171,N_7140);
and U11979 (N_11979,N_8543,N_5446);
nand U11980 (N_11980,N_5942,N_5127);
or U11981 (N_11981,N_8886,N_8614);
and U11982 (N_11982,N_5391,N_5306);
nor U11983 (N_11983,N_9064,N_8594);
or U11984 (N_11984,N_9463,N_9348);
nand U11985 (N_11985,N_5216,N_8859);
or U11986 (N_11986,N_7141,N_5757);
or U11987 (N_11987,N_8081,N_8821);
and U11988 (N_11988,N_8372,N_6943);
nor U11989 (N_11989,N_5654,N_7003);
xnor U11990 (N_11990,N_6202,N_5481);
and U11991 (N_11991,N_7978,N_9735);
and U11992 (N_11992,N_5742,N_7128);
nor U11993 (N_11993,N_6288,N_9812);
or U11994 (N_11994,N_7902,N_6611);
and U11995 (N_11995,N_8408,N_9693);
nor U11996 (N_11996,N_6563,N_8274);
nand U11997 (N_11997,N_5830,N_9909);
or U11998 (N_11998,N_9667,N_8147);
or U11999 (N_11999,N_9474,N_9865);
or U12000 (N_12000,N_9455,N_8437);
or U12001 (N_12001,N_8977,N_7330);
or U12002 (N_12002,N_9155,N_5968);
nand U12003 (N_12003,N_7302,N_5702);
and U12004 (N_12004,N_7867,N_5928);
xor U12005 (N_12005,N_6919,N_9968);
or U12006 (N_12006,N_6436,N_7940);
nand U12007 (N_12007,N_5731,N_7178);
nor U12008 (N_12008,N_8046,N_9555);
and U12009 (N_12009,N_6166,N_7296);
nand U12010 (N_12010,N_5022,N_5681);
nor U12011 (N_12011,N_6105,N_7762);
nand U12012 (N_12012,N_7677,N_9181);
nand U12013 (N_12013,N_5970,N_6363);
or U12014 (N_12014,N_8509,N_5669);
and U12015 (N_12015,N_7204,N_8488);
nand U12016 (N_12016,N_8679,N_8816);
or U12017 (N_12017,N_6935,N_7371);
nor U12018 (N_12018,N_9803,N_8088);
nor U12019 (N_12019,N_7732,N_6713);
nand U12020 (N_12020,N_7085,N_9094);
and U12021 (N_12021,N_7089,N_6320);
and U12022 (N_12022,N_7976,N_8252);
nor U12023 (N_12023,N_6681,N_9727);
and U12024 (N_12024,N_7549,N_9624);
or U12025 (N_12025,N_9025,N_9234);
or U12026 (N_12026,N_8672,N_9335);
or U12027 (N_12027,N_7165,N_6480);
nand U12028 (N_12028,N_5690,N_6455);
nand U12029 (N_12029,N_6925,N_7309);
or U12030 (N_12030,N_6950,N_5521);
nand U12031 (N_12031,N_6818,N_5250);
or U12032 (N_12032,N_5565,N_7729);
nand U12033 (N_12033,N_8558,N_8446);
nor U12034 (N_12034,N_7485,N_6927);
nand U12035 (N_12035,N_7581,N_9358);
or U12036 (N_12036,N_7286,N_6745);
and U12037 (N_12037,N_6056,N_9101);
nand U12038 (N_12038,N_5853,N_9712);
or U12039 (N_12039,N_8676,N_6096);
and U12040 (N_12040,N_8268,N_9309);
xor U12041 (N_12041,N_7810,N_8092);
nor U12042 (N_12042,N_8710,N_6544);
or U12043 (N_12043,N_8729,N_5878);
and U12044 (N_12044,N_9910,N_6438);
nor U12045 (N_12045,N_5629,N_8166);
nor U12046 (N_12046,N_8482,N_6236);
and U12047 (N_12047,N_7830,N_6815);
and U12048 (N_12048,N_5736,N_7794);
nor U12049 (N_12049,N_8618,N_8410);
and U12050 (N_12050,N_7208,N_9894);
nor U12051 (N_12051,N_7138,N_8518);
or U12052 (N_12052,N_7297,N_8987);
or U12053 (N_12053,N_7477,N_5573);
and U12054 (N_12054,N_8447,N_7753);
and U12055 (N_12055,N_5016,N_7742);
nand U12056 (N_12056,N_6739,N_6487);
or U12057 (N_12057,N_8243,N_6130);
nor U12058 (N_12058,N_9722,N_7907);
or U12059 (N_12059,N_6597,N_6414);
or U12060 (N_12060,N_7663,N_9754);
nand U12061 (N_12061,N_6151,N_5792);
and U12062 (N_12062,N_6072,N_7680);
or U12063 (N_12063,N_6714,N_8035);
nor U12064 (N_12064,N_9759,N_8713);
or U12065 (N_12065,N_8295,N_8244);
and U12066 (N_12066,N_6939,N_5199);
or U12067 (N_12067,N_5946,N_7827);
nand U12068 (N_12068,N_9418,N_9531);
nor U12069 (N_12069,N_8018,N_7507);
nor U12070 (N_12070,N_5925,N_7887);
or U12071 (N_12071,N_9747,N_8211);
nor U12072 (N_12072,N_8561,N_8489);
or U12073 (N_12073,N_5561,N_9394);
nand U12074 (N_12074,N_7394,N_5207);
and U12075 (N_12075,N_8694,N_7820);
nor U12076 (N_12076,N_8589,N_9605);
or U12077 (N_12077,N_9085,N_7086);
or U12078 (N_12078,N_5578,N_7946);
nand U12079 (N_12079,N_7935,N_9522);
and U12080 (N_12080,N_8320,N_8689);
nand U12081 (N_12081,N_8687,N_7967);
or U12082 (N_12082,N_8131,N_8691);
and U12083 (N_12083,N_6111,N_9980);
and U12084 (N_12084,N_6308,N_6604);
nand U12085 (N_12085,N_7716,N_6442);
nand U12086 (N_12086,N_6808,N_7610);
and U12087 (N_12087,N_7198,N_9145);
and U12088 (N_12088,N_6777,N_7211);
nand U12089 (N_12089,N_9779,N_7613);
and U12090 (N_12090,N_9919,N_9215);
nand U12091 (N_12091,N_6049,N_9999);
nand U12092 (N_12092,N_7997,N_5110);
or U12093 (N_12093,N_5577,N_6766);
or U12094 (N_12094,N_5028,N_8278);
nor U12095 (N_12095,N_7703,N_6421);
nor U12096 (N_12096,N_9436,N_6081);
nand U12097 (N_12097,N_7883,N_9209);
nand U12098 (N_12098,N_5436,N_5950);
or U12099 (N_12099,N_8124,N_5471);
nand U12100 (N_12100,N_6398,N_6446);
or U12101 (N_12101,N_8564,N_6233);
nand U12102 (N_12102,N_5441,N_6786);
nand U12103 (N_12103,N_9996,N_9148);
nand U12104 (N_12104,N_5524,N_9611);
nand U12105 (N_12105,N_8186,N_5296);
and U12106 (N_12106,N_5680,N_9196);
nor U12107 (N_12107,N_8842,N_5000);
and U12108 (N_12108,N_5318,N_9767);
or U12109 (N_12109,N_8711,N_5927);
or U12110 (N_12110,N_8840,N_6747);
nand U12111 (N_12111,N_5526,N_5891);
or U12112 (N_12112,N_6555,N_7026);
or U12113 (N_12113,N_8633,N_8883);
and U12114 (N_12114,N_7308,N_9216);
nand U12115 (N_12115,N_6741,N_5245);
and U12116 (N_12116,N_6873,N_7342);
nor U12117 (N_12117,N_5291,N_6124);
and U12118 (N_12118,N_9492,N_8884);
and U12119 (N_12119,N_6960,N_5726);
and U12120 (N_12120,N_9945,N_6269);
nor U12121 (N_12121,N_7981,N_6569);
nor U12122 (N_12122,N_7731,N_6565);
or U12123 (N_12123,N_6840,N_5174);
nand U12124 (N_12124,N_5907,N_6955);
nor U12125 (N_12125,N_5862,N_8823);
nand U12126 (N_12126,N_8781,N_9102);
nor U12127 (N_12127,N_9095,N_6868);
and U12128 (N_12128,N_5863,N_5699);
nand U12129 (N_12129,N_9964,N_9138);
or U12130 (N_12130,N_8572,N_8373);
nand U12131 (N_12131,N_5277,N_8954);
or U12132 (N_12132,N_8917,N_8411);
or U12133 (N_12133,N_7157,N_7242);
or U12134 (N_12134,N_8784,N_6605);
nor U12135 (N_12135,N_7175,N_5567);
nor U12136 (N_12136,N_9173,N_6348);
nand U12137 (N_12137,N_5682,N_7922);
nor U12138 (N_12138,N_9369,N_9550);
or U12139 (N_12139,N_7108,N_6027);
or U12140 (N_12140,N_9520,N_5722);
nand U12141 (N_12141,N_6257,N_9813);
nor U12142 (N_12142,N_6273,N_9281);
or U12143 (N_12143,N_6858,N_9170);
nor U12144 (N_12144,N_7717,N_7932);
or U12145 (N_12145,N_6590,N_5948);
nor U12146 (N_12146,N_7080,N_7777);
nand U12147 (N_12147,N_9512,N_8343);
and U12148 (N_12148,N_7111,N_6568);
and U12149 (N_12149,N_7890,N_7775);
and U12150 (N_12150,N_6795,N_6453);
nand U12151 (N_12151,N_8134,N_7047);
nand U12152 (N_12152,N_6386,N_8074);
or U12153 (N_12153,N_6076,N_6381);
nor U12154 (N_12154,N_7046,N_9328);
nor U12155 (N_12155,N_5807,N_7580);
or U12156 (N_12156,N_6354,N_9621);
or U12157 (N_12157,N_7390,N_8642);
nand U12158 (N_12158,N_5014,N_5607);
nand U12159 (N_12159,N_8396,N_8876);
and U12160 (N_12160,N_8873,N_7713);
and U12161 (N_12161,N_8275,N_7367);
nand U12162 (N_12162,N_6016,N_9294);
or U12163 (N_12163,N_6528,N_5990);
nor U12164 (N_12164,N_8548,N_6314);
and U12165 (N_12165,N_7185,N_7494);
nand U12166 (N_12166,N_5932,N_9963);
and U12167 (N_12167,N_9446,N_7248);
nor U12168 (N_12168,N_6100,N_9165);
or U12169 (N_12169,N_6616,N_7964);
nand U12170 (N_12170,N_7991,N_6799);
nor U12171 (N_12171,N_9737,N_6830);
and U12172 (N_12172,N_7521,N_7874);
or U12173 (N_12173,N_5150,N_6899);
nand U12174 (N_12174,N_6472,N_6644);
nand U12175 (N_12175,N_8634,N_7799);
and U12176 (N_12176,N_8229,N_8326);
nand U12177 (N_12177,N_9879,N_8406);
nand U12178 (N_12178,N_5951,N_8863);
and U12179 (N_12179,N_5620,N_7345);
nand U12180 (N_12180,N_5955,N_6309);
nand U12181 (N_12181,N_8983,N_6711);
and U12182 (N_12182,N_7194,N_5410);
nor U12183 (N_12183,N_8242,N_8986);
and U12184 (N_12184,N_5091,N_9636);
and U12185 (N_12185,N_6621,N_5307);
and U12186 (N_12186,N_8668,N_6911);
nand U12187 (N_12187,N_9584,N_6650);
or U12188 (N_12188,N_5514,N_8944);
nor U12189 (N_12189,N_9249,N_7993);
or U12190 (N_12190,N_9706,N_6449);
and U12191 (N_12191,N_5730,N_7247);
or U12192 (N_12192,N_8520,N_6618);
nand U12193 (N_12193,N_5253,N_7660);
or U12194 (N_12194,N_6907,N_8567);
nand U12195 (N_12195,N_5326,N_5770);
and U12196 (N_12196,N_8818,N_8044);
nor U12197 (N_12197,N_8008,N_9901);
and U12198 (N_12198,N_7444,N_5254);
nor U12199 (N_12199,N_8030,N_8500);
or U12200 (N_12200,N_6445,N_9108);
nor U12201 (N_12201,N_7615,N_8608);
or U12202 (N_12202,N_6328,N_9696);
or U12203 (N_12203,N_9925,N_6177);
and U12204 (N_12204,N_7087,N_8623);
and U12205 (N_12205,N_6610,N_6244);
nand U12206 (N_12206,N_9219,N_8652);
and U12207 (N_12207,N_8313,N_5978);
nand U12208 (N_12208,N_8107,N_8677);
and U12209 (N_12209,N_5910,N_7624);
nand U12210 (N_12210,N_6029,N_7524);
nand U12211 (N_12211,N_5652,N_7169);
or U12212 (N_12212,N_5497,N_5660);
or U12213 (N_12213,N_6060,N_7206);
nor U12214 (N_12214,N_8503,N_7472);
and U12215 (N_12215,N_7537,N_6821);
nor U12216 (N_12216,N_5193,N_8493);
and U12217 (N_12217,N_7928,N_7027);
or U12218 (N_12218,N_6800,N_6847);
nor U12219 (N_12219,N_7239,N_9279);
and U12220 (N_12220,N_5363,N_6841);
nor U12221 (N_12221,N_9536,N_8573);
nor U12222 (N_12222,N_7601,N_7202);
nor U12223 (N_12223,N_9854,N_9769);
and U12224 (N_12224,N_5515,N_6866);
nor U12225 (N_12225,N_9297,N_6017);
and U12226 (N_12226,N_7207,N_7079);
and U12227 (N_12227,N_5445,N_9275);
nand U12228 (N_12228,N_6422,N_8638);
nor U12229 (N_12229,N_8553,N_9361);
and U12230 (N_12230,N_8412,N_7063);
or U12231 (N_12231,N_6343,N_5266);
and U12232 (N_12232,N_9770,N_7306);
and U12233 (N_12233,N_7972,N_9589);
nor U12234 (N_12234,N_8469,N_5136);
or U12235 (N_12235,N_6708,N_5665);
and U12236 (N_12236,N_7690,N_9822);
and U12237 (N_12237,N_5009,N_9481);
nor U12238 (N_12238,N_8002,N_5090);
or U12239 (N_12239,N_6836,N_6131);
nor U12240 (N_12240,N_6425,N_5498);
nor U12241 (N_12241,N_5053,N_8014);
nand U12242 (N_12242,N_9162,N_9090);
nor U12243 (N_12243,N_7083,N_6877);
nand U12244 (N_12244,N_5125,N_9938);
nor U12245 (N_12245,N_5334,N_5227);
nor U12246 (N_12246,N_8903,N_9792);
nand U12247 (N_12247,N_9509,N_9264);
or U12248 (N_12248,N_8465,N_9075);
nand U12249 (N_12249,N_5143,N_8231);
and U12250 (N_12250,N_5744,N_6926);
nor U12251 (N_12251,N_7587,N_9590);
xor U12252 (N_12252,N_5013,N_7150);
nor U12253 (N_12253,N_7710,N_9889);
nand U12254 (N_12254,N_7045,N_8270);
nand U12255 (N_12255,N_7301,N_5760);
nand U12256 (N_12256,N_6289,N_5401);
nand U12257 (N_12257,N_6389,N_5552);
nor U12258 (N_12258,N_6798,N_8016);
or U12259 (N_12259,N_7285,N_5798);
nor U12260 (N_12260,N_8656,N_9953);
and U12261 (N_12261,N_9664,N_9932);
or U12262 (N_12262,N_6297,N_5092);
or U12263 (N_12263,N_7233,N_7556);
or U12264 (N_12264,N_8321,N_5685);
nand U12265 (N_12265,N_7582,N_5825);
and U12266 (N_12266,N_6887,N_9289);
or U12267 (N_12267,N_5246,N_7186);
nand U12268 (N_12268,N_7139,N_6211);
nand U12269 (N_12269,N_8811,N_9419);
or U12270 (N_12270,N_5738,N_7744);
nor U12271 (N_12271,N_6759,N_7647);
or U12272 (N_12272,N_9569,N_8738);
or U12273 (N_12273,N_5533,N_7473);
or U12274 (N_12274,N_5958,N_5704);
nand U12275 (N_12275,N_6580,N_7942);
nor U12276 (N_12276,N_9627,N_5257);
and U12277 (N_12277,N_7480,N_9012);
and U12278 (N_12278,N_5906,N_9339);
or U12279 (N_12279,N_8363,N_6928);
nand U12280 (N_12280,N_6684,N_5919);
and U12281 (N_12281,N_6278,N_8386);
or U12282 (N_12282,N_6235,N_7376);
nor U12283 (N_12283,N_6347,N_9435);
and U12284 (N_12284,N_9313,N_9577);
and U12285 (N_12285,N_6039,N_8473);
nand U12286 (N_12286,N_6540,N_5159);
and U12287 (N_12287,N_8801,N_7822);
and U12288 (N_12288,N_5633,N_5920);
or U12289 (N_12289,N_8461,N_9736);
or U12290 (N_12290,N_9896,N_7834);
nor U12291 (N_12291,N_8484,N_5755);
and U12292 (N_12292,N_8427,N_5851);
nor U12293 (N_12293,N_9861,N_9130);
nand U12294 (N_12294,N_9174,N_9382);
nand U12295 (N_12295,N_7149,N_6649);
nand U12296 (N_12296,N_7666,N_5534);
and U12297 (N_12297,N_6728,N_8976);
and U12298 (N_12298,N_6128,N_7969);
nand U12299 (N_12299,N_7975,N_7722);
nor U12300 (N_12300,N_5242,N_9600);
or U12301 (N_12301,N_6243,N_8004);
nor U12302 (N_12302,N_7548,N_5406);
nor U12303 (N_12303,N_9425,N_9248);
nand U12304 (N_12304,N_5451,N_7566);
nor U12305 (N_12305,N_8958,N_6718);
nand U12306 (N_12306,N_6732,N_7007);
nor U12307 (N_12307,N_9393,N_7191);
nand U12308 (N_12308,N_8554,N_6077);
nand U12309 (N_12309,N_7565,N_5998);
nand U12310 (N_12310,N_5132,N_9044);
nor U12311 (N_12311,N_7209,N_7847);
and U12312 (N_12312,N_9653,N_6548);
nand U12313 (N_12313,N_8120,N_8505);
and U12314 (N_12314,N_8094,N_6397);
nand U12315 (N_12315,N_9330,N_9451);
and U12316 (N_12316,N_7314,N_5992);
or U12317 (N_12317,N_5154,N_7943);
or U12318 (N_12318,N_8911,N_9292);
nand U12319 (N_12319,N_6803,N_8845);
nand U12320 (N_12320,N_7720,N_5882);
nand U12321 (N_12321,N_7694,N_6929);
and U12322 (N_12322,N_9710,N_5943);
or U12323 (N_12323,N_5300,N_6005);
nand U12324 (N_12324,N_6602,N_6194);
nor U12325 (N_12325,N_7173,N_7611);
nand U12326 (N_12326,N_7484,N_6123);
or U12327 (N_12327,N_5294,N_5386);
nor U12328 (N_12328,N_9466,N_9848);
and U12329 (N_12329,N_6358,N_7616);
nand U12330 (N_12330,N_6805,N_5039);
nand U12331 (N_12331,N_5672,N_8188);
nand U12332 (N_12332,N_9010,N_6091);
and U12333 (N_12333,N_7467,N_5961);
or U12334 (N_12334,N_6452,N_7037);
or U12335 (N_12335,N_8099,N_8232);
or U12336 (N_12336,N_6165,N_8856);
and U12337 (N_12337,N_5908,N_6073);
or U12338 (N_12338,N_6554,N_7857);
nor U12339 (N_12339,N_6300,N_9015);
nor U12340 (N_12340,N_6794,N_5933);
and U12341 (N_12341,N_7809,N_6920);
or U12342 (N_12342,N_7252,N_9128);
and U12343 (N_12343,N_6185,N_8601);
and U12344 (N_12344,N_7013,N_5050);
nor U12345 (N_12345,N_9453,N_7448);
nand U12346 (N_12346,N_8657,N_6041);
xnor U12347 (N_12347,N_8128,N_5671);
or U12348 (N_12348,N_7385,N_6947);
nand U12349 (N_12349,N_8374,N_9168);
nand U12350 (N_12350,N_7866,N_9544);
nand U12351 (N_12351,N_5098,N_6025);
nand U12352 (N_12352,N_7727,N_7105);
and U12353 (N_12353,N_6889,N_7553);
and U12354 (N_12354,N_9490,N_5011);
nand U12355 (N_12355,N_8297,N_8357);
nor U12356 (N_12356,N_9042,N_5105);
and U12357 (N_12357,N_8156,N_7881);
and U12358 (N_12358,N_8333,N_5063);
or U12359 (N_12359,N_5569,N_9687);
and U12360 (N_12360,N_7589,N_7162);
and U12361 (N_12361,N_8753,N_5914);
nand U12362 (N_12362,N_5255,N_6980);
nand U12363 (N_12363,N_5137,N_9749);
and U12364 (N_12364,N_5739,N_7213);
nor U12365 (N_12365,N_5559,N_9534);
and U12366 (N_12366,N_7055,N_9886);
nor U12367 (N_12367,N_5070,N_6838);
or U12368 (N_12368,N_7054,N_7219);
nor U12369 (N_12369,N_6521,N_6116);
nor U12370 (N_12370,N_8727,N_5356);
nor U12371 (N_12371,N_6906,N_7445);
nor U12372 (N_12372,N_5896,N_8839);
nand U12373 (N_12373,N_9731,N_7110);
and U12374 (N_12374,N_7842,N_6473);
nor U12375 (N_12375,N_8595,N_8783);
nand U12376 (N_12376,N_6576,N_7563);
nor U12377 (N_12377,N_9469,N_5509);
nand U12378 (N_12378,N_6964,N_9943);
or U12379 (N_12379,N_6744,N_8615);
or U12380 (N_12380,N_9144,N_7721);
nor U12381 (N_12381,N_8581,N_9994);
and U12382 (N_12382,N_6333,N_7541);
nor U12383 (N_12383,N_5124,N_8780);
nor U12384 (N_12384,N_6710,N_6247);
nor U12385 (N_12385,N_6301,N_6137);
and U12386 (N_12386,N_9572,N_8405);
and U12387 (N_12387,N_5556,N_9739);
and U12388 (N_12388,N_7586,N_9790);
nor U12389 (N_12389,N_7154,N_5913);
or U12390 (N_12390,N_9912,N_7906);
nor U12391 (N_12391,N_5215,N_8777);
or U12392 (N_12392,N_8216,N_8440);
nor U12393 (N_12393,N_8109,N_9815);
and U12394 (N_12394,N_9558,N_6851);
or U12395 (N_12395,N_5425,N_5430);
and U12396 (N_12396,N_5588,N_5911);
or U12397 (N_12397,N_7726,N_5295);
nor U12398 (N_12398,N_7600,N_5437);
and U12399 (N_12399,N_7885,N_5434);
nor U12400 (N_12400,N_6248,N_7227);
or U12401 (N_12401,N_9035,N_6048);
nand U12402 (N_12402,N_9845,N_5686);
nand U12403 (N_12403,N_5238,N_7786);
or U12404 (N_12404,N_7005,N_5935);
or U12405 (N_12405,N_7668,N_5439);
and U12406 (N_12406,N_6547,N_5850);
nand U12407 (N_12407,N_8289,N_5145);
and U12408 (N_12408,N_5758,N_6391);
or U12409 (N_12409,N_7835,N_7215);
xor U12410 (N_12410,N_6606,N_8893);
and U12411 (N_12411,N_9232,N_6559);
nor U12412 (N_12412,N_5769,N_5045);
nor U12413 (N_12413,N_9262,N_6340);
nor U12414 (N_12414,N_9202,N_5485);
or U12415 (N_12415,N_9850,N_7646);
nand U12416 (N_12416,N_8837,N_9217);
and U12417 (N_12417,N_7015,N_9488);
nor U12418 (N_12418,N_8715,N_5165);
and U12419 (N_12419,N_5544,N_6462);
nor U12420 (N_12420,N_8039,N_8384);
xnor U12421 (N_12421,N_8871,N_7256);
nand U12422 (N_12422,N_9517,N_5487);
nand U12423 (N_12423,N_8899,N_6476);
nor U12424 (N_12424,N_8068,N_5580);
nor U12425 (N_12425,N_8085,N_7853);
nor U12426 (N_12426,N_9843,N_9761);
and U12427 (N_12427,N_7865,N_5141);
or U12428 (N_12428,N_7167,N_9068);
and U12429 (N_12429,N_6727,N_9320);
and U12430 (N_12430,N_6164,N_5785);
nor U12431 (N_12431,N_8507,N_7811);
and U12432 (N_12432,N_9448,N_6050);
and U12433 (N_12433,N_5085,N_7947);
nand U12434 (N_12434,N_9871,N_7934);
nand U12435 (N_12435,N_6722,N_8442);
nand U12436 (N_12436,N_8483,N_6153);
and U12437 (N_12437,N_7408,N_7913);
or U12438 (N_12438,N_7249,N_8063);
or U12439 (N_12439,N_9093,N_7017);
and U12440 (N_12440,N_5168,N_6770);
and U12441 (N_12441,N_9594,N_8308);
nor U12442 (N_12442,N_9468,N_7868);
nor U12443 (N_12443,N_5656,N_7062);
nand U12444 (N_12444,N_5263,N_5886);
nand U12445 (N_12445,N_5601,N_6034);
nor U12446 (N_12446,N_8939,N_7474);
nand U12447 (N_12447,N_6639,N_9574);
nand U12448 (N_12448,N_7039,N_6312);
nand U12449 (N_12449,N_8826,N_8914);
nand U12450 (N_12450,N_5847,N_6574);
or U12451 (N_12451,N_8776,N_5540);
nand U12452 (N_12452,N_5963,N_8264);
or U12453 (N_12453,N_5042,N_5688);
or U12454 (N_12454,N_8439,N_9475);
nor U12455 (N_12455,N_6762,N_6225);
or U12456 (N_12456,N_5492,N_9720);
or U12457 (N_12457,N_6864,N_5469);
and U12458 (N_12458,N_8228,N_6437);
or U12459 (N_12459,N_5495,N_6806);
nand U12460 (N_12460,N_8084,N_5201);
or U12461 (N_12461,N_7897,N_5621);
or U12462 (N_12462,N_7884,N_7763);
nor U12463 (N_12463,N_6338,N_5276);
nor U12464 (N_12464,N_7218,N_8154);
nand U12465 (N_12465,N_7648,N_6585);
and U12466 (N_12466,N_7126,N_9526);
and U12467 (N_12467,N_5568,N_7662);
nor U12468 (N_12468,N_8368,N_5362);
or U12469 (N_12469,N_5562,N_6969);
nor U12470 (N_12470,N_9758,N_7659);
nor U12471 (N_12471,N_9377,N_6530);
or U12472 (N_12472,N_8280,N_5440);
or U12473 (N_12473,N_9265,N_9771);
nand U12474 (N_12474,N_9046,N_8790);
or U12475 (N_12475,N_9205,N_6261);
nor U12476 (N_12476,N_5775,N_8946);
xor U12477 (N_12477,N_8942,N_5477);
nor U12478 (N_12478,N_5121,N_5986);
nor U12479 (N_12479,N_5774,N_8724);
nor U12480 (N_12480,N_8054,N_8832);
nor U12481 (N_12481,N_9026,N_5805);
and U12482 (N_12482,N_6022,N_7862);
or U12483 (N_12483,N_6893,N_5841);
nor U12484 (N_12484,N_6324,N_7520);
and U12485 (N_12485,N_6692,N_6507);
nor U12486 (N_12486,N_7300,N_7683);
or U12487 (N_12487,N_8620,N_9940);
and U12488 (N_12488,N_9283,N_7322);
xor U12489 (N_12489,N_9826,N_5916);
nand U12490 (N_12490,N_7214,N_7562);
and U12491 (N_12491,N_9089,N_6850);
nand U12492 (N_12492,N_5426,N_6753);
nor U12493 (N_12493,N_9460,N_8602);
and U12494 (N_12494,N_7719,N_7765);
or U12495 (N_12495,N_6958,N_5112);
xor U12496 (N_12496,N_9059,N_5072);
nor U12497 (N_12497,N_5180,N_9395);
nand U12498 (N_12498,N_8024,N_6625);
or U12499 (N_12499,N_9381,N_7924);
nor U12500 (N_12500,N_5229,N_5058);
and U12501 (N_12501,N_6900,N_8773);
nand U12502 (N_12502,N_5733,N_6980);
nand U12503 (N_12503,N_7857,N_9643);
nand U12504 (N_12504,N_9620,N_6980);
or U12505 (N_12505,N_5393,N_5368);
nor U12506 (N_12506,N_7223,N_7529);
or U12507 (N_12507,N_9940,N_9304);
nor U12508 (N_12508,N_7728,N_5931);
and U12509 (N_12509,N_5462,N_8341);
nand U12510 (N_12510,N_6436,N_9782);
nor U12511 (N_12511,N_5169,N_8565);
nand U12512 (N_12512,N_7691,N_7175);
nor U12513 (N_12513,N_6192,N_8238);
nor U12514 (N_12514,N_9575,N_8919);
and U12515 (N_12515,N_6920,N_8473);
nor U12516 (N_12516,N_8518,N_8249);
or U12517 (N_12517,N_6855,N_6047);
nor U12518 (N_12518,N_9273,N_5590);
nor U12519 (N_12519,N_9642,N_8119);
and U12520 (N_12520,N_9174,N_8391);
or U12521 (N_12521,N_8819,N_5293);
nor U12522 (N_12522,N_6145,N_9912);
or U12523 (N_12523,N_8301,N_5658);
nor U12524 (N_12524,N_5618,N_8365);
nor U12525 (N_12525,N_5527,N_5565);
and U12526 (N_12526,N_8178,N_8191);
and U12527 (N_12527,N_7219,N_9578);
and U12528 (N_12528,N_6138,N_6079);
nor U12529 (N_12529,N_8243,N_8436);
nand U12530 (N_12530,N_9022,N_7131);
nand U12531 (N_12531,N_6344,N_9464);
or U12532 (N_12532,N_6259,N_5692);
or U12533 (N_12533,N_9995,N_5871);
nand U12534 (N_12534,N_7273,N_9667);
and U12535 (N_12535,N_6042,N_8279);
nand U12536 (N_12536,N_9227,N_8831);
nor U12537 (N_12537,N_5882,N_7567);
nand U12538 (N_12538,N_7258,N_6935);
nor U12539 (N_12539,N_5635,N_9054);
nor U12540 (N_12540,N_7412,N_9801);
nor U12541 (N_12541,N_5225,N_9860);
and U12542 (N_12542,N_9445,N_9943);
nand U12543 (N_12543,N_5489,N_5677);
and U12544 (N_12544,N_7723,N_9114);
and U12545 (N_12545,N_8127,N_5430);
nor U12546 (N_12546,N_8331,N_9783);
nand U12547 (N_12547,N_8408,N_5488);
nor U12548 (N_12548,N_5806,N_7467);
nand U12549 (N_12549,N_5895,N_9648);
nor U12550 (N_12550,N_8850,N_6710);
and U12551 (N_12551,N_6701,N_6806);
nand U12552 (N_12552,N_5386,N_5342);
or U12553 (N_12553,N_9358,N_8981);
nor U12554 (N_12554,N_8520,N_7618);
or U12555 (N_12555,N_8149,N_5861);
or U12556 (N_12556,N_5379,N_7417);
and U12557 (N_12557,N_9128,N_5586);
nand U12558 (N_12558,N_7570,N_5035);
nand U12559 (N_12559,N_7583,N_9927);
or U12560 (N_12560,N_9998,N_9819);
and U12561 (N_12561,N_8657,N_6319);
nor U12562 (N_12562,N_6719,N_7619);
or U12563 (N_12563,N_9944,N_5732);
nand U12564 (N_12564,N_6260,N_6697);
or U12565 (N_12565,N_9198,N_9223);
or U12566 (N_12566,N_6017,N_7911);
and U12567 (N_12567,N_8553,N_9636);
and U12568 (N_12568,N_9684,N_7619);
or U12569 (N_12569,N_9075,N_6555);
or U12570 (N_12570,N_6104,N_5577);
or U12571 (N_12571,N_8602,N_9821);
nor U12572 (N_12572,N_9243,N_8203);
nor U12573 (N_12573,N_9317,N_8008);
and U12574 (N_12574,N_9786,N_8231);
or U12575 (N_12575,N_7112,N_8179);
or U12576 (N_12576,N_9416,N_7814);
nor U12577 (N_12577,N_5543,N_6644);
or U12578 (N_12578,N_7225,N_6170);
and U12579 (N_12579,N_8747,N_7674);
or U12580 (N_12580,N_5648,N_8517);
and U12581 (N_12581,N_6476,N_6534);
nor U12582 (N_12582,N_5187,N_7395);
and U12583 (N_12583,N_6636,N_8442);
or U12584 (N_12584,N_5346,N_8347);
nand U12585 (N_12585,N_7970,N_6318);
and U12586 (N_12586,N_6861,N_5555);
nor U12587 (N_12587,N_8855,N_7791);
nor U12588 (N_12588,N_6762,N_6005);
nand U12589 (N_12589,N_7453,N_8008);
and U12590 (N_12590,N_5978,N_5513);
and U12591 (N_12591,N_7032,N_5721);
nor U12592 (N_12592,N_8744,N_8933);
nor U12593 (N_12593,N_9229,N_5951);
and U12594 (N_12594,N_6532,N_6943);
and U12595 (N_12595,N_6214,N_7507);
nor U12596 (N_12596,N_6565,N_8080);
or U12597 (N_12597,N_6997,N_5523);
nand U12598 (N_12598,N_7400,N_5201);
and U12599 (N_12599,N_7687,N_8276);
nor U12600 (N_12600,N_9857,N_5276);
nor U12601 (N_12601,N_5479,N_9637);
nand U12602 (N_12602,N_5788,N_6856);
and U12603 (N_12603,N_8279,N_9052);
nand U12604 (N_12604,N_7788,N_5216);
and U12605 (N_12605,N_5015,N_9652);
or U12606 (N_12606,N_9733,N_6169);
nor U12607 (N_12607,N_7866,N_6924);
nor U12608 (N_12608,N_5510,N_5635);
xnor U12609 (N_12609,N_8149,N_7882);
nor U12610 (N_12610,N_9119,N_5737);
and U12611 (N_12611,N_8666,N_5946);
nor U12612 (N_12612,N_7562,N_6353);
or U12613 (N_12613,N_7169,N_9289);
nand U12614 (N_12614,N_5008,N_9805);
nor U12615 (N_12615,N_6754,N_7007);
nor U12616 (N_12616,N_6846,N_5166);
or U12617 (N_12617,N_8044,N_6862);
nor U12618 (N_12618,N_9887,N_6883);
and U12619 (N_12619,N_8525,N_5945);
nor U12620 (N_12620,N_5400,N_8093);
nor U12621 (N_12621,N_5556,N_7212);
nand U12622 (N_12622,N_8265,N_6309);
nand U12623 (N_12623,N_8705,N_6128);
nor U12624 (N_12624,N_9733,N_7268);
or U12625 (N_12625,N_6539,N_7463);
and U12626 (N_12626,N_7042,N_8812);
nor U12627 (N_12627,N_8022,N_7060);
nor U12628 (N_12628,N_6395,N_6406);
nor U12629 (N_12629,N_9604,N_9942);
nand U12630 (N_12630,N_6769,N_6613);
nor U12631 (N_12631,N_7557,N_7512);
or U12632 (N_12632,N_9130,N_6499);
nor U12633 (N_12633,N_5927,N_8655);
or U12634 (N_12634,N_5612,N_8150);
nor U12635 (N_12635,N_6810,N_5892);
or U12636 (N_12636,N_6297,N_8227);
nand U12637 (N_12637,N_9108,N_8741);
and U12638 (N_12638,N_7672,N_6166);
nor U12639 (N_12639,N_9490,N_7116);
nand U12640 (N_12640,N_5916,N_7485);
nand U12641 (N_12641,N_8347,N_5122);
and U12642 (N_12642,N_7224,N_7209);
nand U12643 (N_12643,N_7689,N_5878);
nand U12644 (N_12644,N_9383,N_5784);
nor U12645 (N_12645,N_6933,N_8287);
and U12646 (N_12646,N_5729,N_6957);
or U12647 (N_12647,N_6448,N_7598);
or U12648 (N_12648,N_7680,N_9379);
nand U12649 (N_12649,N_7127,N_5088);
and U12650 (N_12650,N_5087,N_5288);
nand U12651 (N_12651,N_9377,N_7199);
nand U12652 (N_12652,N_5542,N_5327);
nand U12653 (N_12653,N_5931,N_7598);
nand U12654 (N_12654,N_6588,N_9123);
or U12655 (N_12655,N_5711,N_6320);
nor U12656 (N_12656,N_6859,N_6327);
xor U12657 (N_12657,N_5830,N_8204);
nor U12658 (N_12658,N_5877,N_5071);
nand U12659 (N_12659,N_9753,N_8155);
nand U12660 (N_12660,N_8173,N_9860);
or U12661 (N_12661,N_9279,N_7820);
or U12662 (N_12662,N_7927,N_5715);
nand U12663 (N_12663,N_5899,N_8722);
or U12664 (N_12664,N_8180,N_9377);
or U12665 (N_12665,N_5262,N_9772);
nand U12666 (N_12666,N_8881,N_9434);
and U12667 (N_12667,N_5001,N_5643);
and U12668 (N_12668,N_6926,N_6749);
or U12669 (N_12669,N_9131,N_9355);
and U12670 (N_12670,N_9133,N_5514);
and U12671 (N_12671,N_6550,N_6784);
nor U12672 (N_12672,N_7641,N_7389);
and U12673 (N_12673,N_9417,N_9096);
and U12674 (N_12674,N_6672,N_7850);
and U12675 (N_12675,N_5866,N_6156);
or U12676 (N_12676,N_5912,N_9715);
or U12677 (N_12677,N_7326,N_6466);
nor U12678 (N_12678,N_7159,N_5002);
or U12679 (N_12679,N_6279,N_8446);
nor U12680 (N_12680,N_8061,N_5595);
or U12681 (N_12681,N_6173,N_6531);
nand U12682 (N_12682,N_7539,N_8443);
nand U12683 (N_12683,N_6448,N_8108);
nand U12684 (N_12684,N_7534,N_6240);
nand U12685 (N_12685,N_6762,N_8244);
and U12686 (N_12686,N_7997,N_7044);
nand U12687 (N_12687,N_9069,N_5745);
nor U12688 (N_12688,N_9024,N_5676);
or U12689 (N_12689,N_7935,N_6382);
or U12690 (N_12690,N_8655,N_8377);
or U12691 (N_12691,N_8667,N_6011);
nor U12692 (N_12692,N_5701,N_7633);
and U12693 (N_12693,N_9503,N_6903);
xnor U12694 (N_12694,N_5209,N_7256);
and U12695 (N_12695,N_6259,N_8996);
nand U12696 (N_12696,N_6649,N_8241);
nand U12697 (N_12697,N_6368,N_5340);
or U12698 (N_12698,N_7555,N_8270);
or U12699 (N_12699,N_8694,N_9535);
nand U12700 (N_12700,N_8378,N_8870);
nor U12701 (N_12701,N_5065,N_6713);
or U12702 (N_12702,N_8270,N_6609);
or U12703 (N_12703,N_7893,N_7220);
nor U12704 (N_12704,N_9122,N_7642);
nor U12705 (N_12705,N_5882,N_8182);
or U12706 (N_12706,N_5920,N_9071);
or U12707 (N_12707,N_5046,N_8722);
nand U12708 (N_12708,N_6188,N_6544);
nand U12709 (N_12709,N_8790,N_5030);
xor U12710 (N_12710,N_8299,N_6302);
nand U12711 (N_12711,N_7375,N_7987);
nand U12712 (N_12712,N_7542,N_8237);
and U12713 (N_12713,N_5458,N_8419);
nand U12714 (N_12714,N_8465,N_8353);
nand U12715 (N_12715,N_7694,N_7108);
and U12716 (N_12716,N_8796,N_7352);
or U12717 (N_12717,N_7954,N_7212);
nor U12718 (N_12718,N_7499,N_8711);
or U12719 (N_12719,N_8456,N_5542);
and U12720 (N_12720,N_5448,N_6126);
nand U12721 (N_12721,N_6957,N_8553);
and U12722 (N_12722,N_7696,N_7081);
and U12723 (N_12723,N_9049,N_8943);
nand U12724 (N_12724,N_6571,N_8524);
nand U12725 (N_12725,N_8838,N_9662);
nand U12726 (N_12726,N_5499,N_7550);
or U12727 (N_12727,N_8801,N_8985);
or U12728 (N_12728,N_9071,N_7810);
and U12729 (N_12729,N_6731,N_6497);
nand U12730 (N_12730,N_7062,N_6278);
and U12731 (N_12731,N_6197,N_9470);
nand U12732 (N_12732,N_5025,N_6197);
nor U12733 (N_12733,N_7928,N_7971);
and U12734 (N_12734,N_9680,N_7428);
or U12735 (N_12735,N_9549,N_9512);
nor U12736 (N_12736,N_5734,N_8150);
and U12737 (N_12737,N_7154,N_5705);
or U12738 (N_12738,N_9811,N_8985);
nand U12739 (N_12739,N_7265,N_5905);
or U12740 (N_12740,N_7516,N_5874);
nand U12741 (N_12741,N_9029,N_6915);
nor U12742 (N_12742,N_6463,N_7585);
nand U12743 (N_12743,N_9968,N_9720);
nor U12744 (N_12744,N_6990,N_7903);
or U12745 (N_12745,N_5362,N_7462);
or U12746 (N_12746,N_7426,N_6261);
nand U12747 (N_12747,N_7262,N_8967);
and U12748 (N_12748,N_9432,N_7623);
and U12749 (N_12749,N_8665,N_6854);
and U12750 (N_12750,N_7947,N_8119);
and U12751 (N_12751,N_7065,N_9324);
nor U12752 (N_12752,N_8430,N_6769);
nor U12753 (N_12753,N_5601,N_5566);
nor U12754 (N_12754,N_8588,N_7411);
nand U12755 (N_12755,N_5902,N_9826);
and U12756 (N_12756,N_7541,N_9864);
xnor U12757 (N_12757,N_6038,N_8951);
or U12758 (N_12758,N_8418,N_7413);
or U12759 (N_12759,N_6686,N_7359);
or U12760 (N_12760,N_7115,N_8374);
or U12761 (N_12761,N_8047,N_9624);
or U12762 (N_12762,N_8484,N_8723);
nor U12763 (N_12763,N_6534,N_5955);
or U12764 (N_12764,N_8793,N_8719);
and U12765 (N_12765,N_8389,N_5037);
nor U12766 (N_12766,N_6161,N_7542);
and U12767 (N_12767,N_6949,N_8623);
or U12768 (N_12768,N_5216,N_7253);
and U12769 (N_12769,N_6056,N_9621);
nand U12770 (N_12770,N_7582,N_7041);
and U12771 (N_12771,N_8376,N_6347);
nand U12772 (N_12772,N_6494,N_7737);
or U12773 (N_12773,N_9737,N_5176);
and U12774 (N_12774,N_6636,N_6482);
and U12775 (N_12775,N_6559,N_5437);
and U12776 (N_12776,N_6994,N_8817);
nand U12777 (N_12777,N_5919,N_7883);
nor U12778 (N_12778,N_5472,N_6167);
nand U12779 (N_12779,N_7746,N_6371);
nand U12780 (N_12780,N_7207,N_6514);
or U12781 (N_12781,N_7303,N_5619);
and U12782 (N_12782,N_8871,N_7709);
and U12783 (N_12783,N_7134,N_7638);
nor U12784 (N_12784,N_8522,N_8866);
and U12785 (N_12785,N_9493,N_5246);
and U12786 (N_12786,N_9704,N_7821);
nor U12787 (N_12787,N_8551,N_8152);
xnor U12788 (N_12788,N_7149,N_5135);
nand U12789 (N_12789,N_7077,N_8217);
and U12790 (N_12790,N_5204,N_7307);
and U12791 (N_12791,N_8904,N_5065);
nor U12792 (N_12792,N_7041,N_8548);
and U12793 (N_12793,N_9688,N_5559);
and U12794 (N_12794,N_9819,N_5083);
xor U12795 (N_12795,N_5597,N_7092);
nor U12796 (N_12796,N_7484,N_8471);
or U12797 (N_12797,N_6500,N_6339);
nand U12798 (N_12798,N_9492,N_5153);
nor U12799 (N_12799,N_6494,N_5994);
nor U12800 (N_12800,N_5435,N_6368);
or U12801 (N_12801,N_6681,N_8012);
nor U12802 (N_12802,N_8949,N_6193);
nand U12803 (N_12803,N_8583,N_8722);
or U12804 (N_12804,N_5036,N_7657);
and U12805 (N_12805,N_8373,N_5203);
and U12806 (N_12806,N_5298,N_9903);
xnor U12807 (N_12807,N_8690,N_9267);
or U12808 (N_12808,N_8787,N_8401);
or U12809 (N_12809,N_6217,N_9333);
or U12810 (N_12810,N_7841,N_8171);
nand U12811 (N_12811,N_6306,N_5450);
nand U12812 (N_12812,N_5824,N_5079);
nor U12813 (N_12813,N_9703,N_6655);
nor U12814 (N_12814,N_8525,N_5613);
nor U12815 (N_12815,N_9916,N_5599);
nor U12816 (N_12816,N_8694,N_6244);
nand U12817 (N_12817,N_5013,N_7345);
and U12818 (N_12818,N_6942,N_5038);
and U12819 (N_12819,N_8940,N_5990);
nand U12820 (N_12820,N_5733,N_9163);
nor U12821 (N_12821,N_5276,N_7119);
or U12822 (N_12822,N_6986,N_6522);
or U12823 (N_12823,N_9056,N_8388);
nor U12824 (N_12824,N_9061,N_5261);
or U12825 (N_12825,N_9560,N_7781);
nand U12826 (N_12826,N_5807,N_8739);
nor U12827 (N_12827,N_9764,N_8823);
nand U12828 (N_12828,N_9248,N_6181);
or U12829 (N_12829,N_6011,N_5028);
or U12830 (N_12830,N_6292,N_8155);
nor U12831 (N_12831,N_6103,N_8100);
or U12832 (N_12832,N_6277,N_6378);
nor U12833 (N_12833,N_6113,N_9094);
nand U12834 (N_12834,N_9444,N_6040);
and U12835 (N_12835,N_7504,N_8490);
nand U12836 (N_12836,N_9014,N_7472);
nor U12837 (N_12837,N_8691,N_8927);
and U12838 (N_12838,N_8676,N_5503);
and U12839 (N_12839,N_8321,N_8660);
and U12840 (N_12840,N_7382,N_6724);
nor U12841 (N_12841,N_6985,N_6962);
and U12842 (N_12842,N_5578,N_5665);
and U12843 (N_12843,N_7714,N_9999);
nor U12844 (N_12844,N_6407,N_5104);
or U12845 (N_12845,N_8992,N_9110);
nor U12846 (N_12846,N_5119,N_8482);
nor U12847 (N_12847,N_7640,N_6446);
and U12848 (N_12848,N_8210,N_5150);
or U12849 (N_12849,N_8464,N_7339);
xor U12850 (N_12850,N_7532,N_6635);
and U12851 (N_12851,N_8146,N_6833);
and U12852 (N_12852,N_5539,N_6996);
nand U12853 (N_12853,N_6458,N_5952);
nand U12854 (N_12854,N_8710,N_7189);
nand U12855 (N_12855,N_6712,N_7973);
nor U12856 (N_12856,N_7848,N_5425);
or U12857 (N_12857,N_6215,N_7451);
and U12858 (N_12858,N_5569,N_8217);
nor U12859 (N_12859,N_8440,N_5810);
nand U12860 (N_12860,N_5212,N_8029);
and U12861 (N_12861,N_6188,N_5643);
nor U12862 (N_12862,N_5089,N_7809);
or U12863 (N_12863,N_7302,N_8267);
and U12864 (N_12864,N_9214,N_5997);
nor U12865 (N_12865,N_5163,N_9519);
and U12866 (N_12866,N_5812,N_7720);
and U12867 (N_12867,N_5386,N_8263);
nor U12868 (N_12868,N_7400,N_8746);
and U12869 (N_12869,N_6070,N_6842);
and U12870 (N_12870,N_6374,N_5602);
or U12871 (N_12871,N_8142,N_5854);
or U12872 (N_12872,N_5224,N_5815);
and U12873 (N_12873,N_6480,N_9908);
nor U12874 (N_12874,N_6839,N_9606);
nand U12875 (N_12875,N_8223,N_5233);
nor U12876 (N_12876,N_7903,N_8500);
or U12877 (N_12877,N_7440,N_5640);
or U12878 (N_12878,N_8571,N_7079);
nand U12879 (N_12879,N_6320,N_8126);
and U12880 (N_12880,N_7604,N_5306);
and U12881 (N_12881,N_9865,N_5493);
nand U12882 (N_12882,N_6469,N_6941);
nand U12883 (N_12883,N_7251,N_5028);
and U12884 (N_12884,N_9739,N_9110);
and U12885 (N_12885,N_8040,N_8802);
nand U12886 (N_12886,N_5054,N_9267);
and U12887 (N_12887,N_7460,N_5623);
or U12888 (N_12888,N_7131,N_9299);
nor U12889 (N_12889,N_5260,N_6960);
nor U12890 (N_12890,N_6977,N_7427);
or U12891 (N_12891,N_8540,N_5836);
and U12892 (N_12892,N_9143,N_8535);
or U12893 (N_12893,N_7230,N_8480);
and U12894 (N_12894,N_8654,N_8144);
nor U12895 (N_12895,N_9116,N_8962);
nand U12896 (N_12896,N_7856,N_6145);
and U12897 (N_12897,N_7242,N_9427);
nand U12898 (N_12898,N_7996,N_5837);
nand U12899 (N_12899,N_5665,N_6014);
nor U12900 (N_12900,N_9288,N_8828);
nand U12901 (N_12901,N_9320,N_8454);
nor U12902 (N_12902,N_6079,N_7290);
nand U12903 (N_12903,N_9672,N_8456);
nand U12904 (N_12904,N_6232,N_5666);
nand U12905 (N_12905,N_5776,N_6831);
and U12906 (N_12906,N_9738,N_7482);
nor U12907 (N_12907,N_7129,N_7143);
and U12908 (N_12908,N_9909,N_5874);
or U12909 (N_12909,N_6536,N_5648);
nor U12910 (N_12910,N_5715,N_9011);
nor U12911 (N_12911,N_8262,N_6809);
nor U12912 (N_12912,N_7552,N_7053);
or U12913 (N_12913,N_8183,N_7267);
or U12914 (N_12914,N_7798,N_7148);
nand U12915 (N_12915,N_6815,N_9707);
nor U12916 (N_12916,N_5044,N_7330);
and U12917 (N_12917,N_7102,N_9616);
and U12918 (N_12918,N_7741,N_5424);
and U12919 (N_12919,N_7851,N_6093);
nor U12920 (N_12920,N_6328,N_8399);
and U12921 (N_12921,N_5907,N_6404);
nand U12922 (N_12922,N_8038,N_8438);
and U12923 (N_12923,N_6065,N_9477);
and U12924 (N_12924,N_8020,N_6566);
nand U12925 (N_12925,N_7439,N_8326);
nor U12926 (N_12926,N_5901,N_5829);
nor U12927 (N_12927,N_7019,N_5536);
nor U12928 (N_12928,N_5397,N_7066);
and U12929 (N_12929,N_7713,N_9901);
nor U12930 (N_12930,N_9097,N_8776);
or U12931 (N_12931,N_6204,N_9647);
nor U12932 (N_12932,N_7829,N_8396);
nand U12933 (N_12933,N_7702,N_6081);
or U12934 (N_12934,N_6599,N_8221);
nor U12935 (N_12935,N_7982,N_6369);
and U12936 (N_12936,N_7944,N_7353);
and U12937 (N_12937,N_9173,N_9179);
xnor U12938 (N_12938,N_8725,N_9186);
nor U12939 (N_12939,N_5618,N_6761);
nor U12940 (N_12940,N_6971,N_8562);
or U12941 (N_12941,N_9229,N_6755);
and U12942 (N_12942,N_8437,N_5907);
nand U12943 (N_12943,N_7473,N_5434);
and U12944 (N_12944,N_7931,N_6763);
nand U12945 (N_12945,N_7890,N_5735);
or U12946 (N_12946,N_9082,N_9171);
nor U12947 (N_12947,N_7968,N_8611);
nor U12948 (N_12948,N_7983,N_5229);
or U12949 (N_12949,N_7641,N_7395);
and U12950 (N_12950,N_9838,N_8831);
and U12951 (N_12951,N_7678,N_5334);
nor U12952 (N_12952,N_7171,N_6427);
nor U12953 (N_12953,N_9759,N_7277);
nand U12954 (N_12954,N_5030,N_7287);
nor U12955 (N_12955,N_7975,N_5306);
nor U12956 (N_12956,N_7947,N_5983);
nand U12957 (N_12957,N_8781,N_8979);
or U12958 (N_12958,N_9178,N_9315);
nand U12959 (N_12959,N_7565,N_7017);
and U12960 (N_12960,N_7468,N_9018);
or U12961 (N_12961,N_7087,N_5274);
and U12962 (N_12962,N_7206,N_5964);
nor U12963 (N_12963,N_8737,N_6230);
and U12964 (N_12964,N_8013,N_7506);
or U12965 (N_12965,N_7886,N_8899);
nand U12966 (N_12966,N_8423,N_7184);
nand U12967 (N_12967,N_8686,N_9776);
and U12968 (N_12968,N_7727,N_8018);
and U12969 (N_12969,N_9071,N_5760);
or U12970 (N_12970,N_5364,N_6312);
nor U12971 (N_12971,N_6878,N_5309);
or U12972 (N_12972,N_5184,N_5265);
and U12973 (N_12973,N_9697,N_6466);
or U12974 (N_12974,N_6030,N_9964);
or U12975 (N_12975,N_5064,N_9222);
nand U12976 (N_12976,N_6258,N_6086);
and U12977 (N_12977,N_6048,N_9819);
nand U12978 (N_12978,N_8984,N_7380);
or U12979 (N_12979,N_9917,N_6376);
or U12980 (N_12980,N_6426,N_7359);
nand U12981 (N_12981,N_7075,N_8720);
and U12982 (N_12982,N_6257,N_6383);
nand U12983 (N_12983,N_5711,N_7083);
nor U12984 (N_12984,N_5128,N_8578);
and U12985 (N_12985,N_6190,N_7377);
nor U12986 (N_12986,N_8882,N_9906);
nand U12987 (N_12987,N_5090,N_6619);
nor U12988 (N_12988,N_7269,N_6204);
nor U12989 (N_12989,N_8975,N_9001);
nor U12990 (N_12990,N_7665,N_8225);
and U12991 (N_12991,N_6344,N_7723);
nand U12992 (N_12992,N_8741,N_9402);
or U12993 (N_12993,N_8064,N_6167);
nand U12994 (N_12994,N_8575,N_6748);
nand U12995 (N_12995,N_5576,N_5769);
or U12996 (N_12996,N_6947,N_6793);
nand U12997 (N_12997,N_9367,N_6473);
or U12998 (N_12998,N_7086,N_8451);
and U12999 (N_12999,N_8161,N_7657);
and U13000 (N_13000,N_7127,N_7413);
nand U13001 (N_13001,N_6263,N_6527);
nor U13002 (N_13002,N_9141,N_7708);
and U13003 (N_13003,N_5678,N_5111);
and U13004 (N_13004,N_5788,N_8182);
nand U13005 (N_13005,N_5025,N_6730);
or U13006 (N_13006,N_6923,N_9986);
nand U13007 (N_13007,N_9886,N_5196);
nor U13008 (N_13008,N_6721,N_6870);
nand U13009 (N_13009,N_8040,N_9019);
and U13010 (N_13010,N_8685,N_7436);
and U13011 (N_13011,N_8730,N_5354);
nor U13012 (N_13012,N_5828,N_7569);
nand U13013 (N_13013,N_6540,N_9698);
and U13014 (N_13014,N_5619,N_6350);
nand U13015 (N_13015,N_7858,N_6895);
nor U13016 (N_13016,N_6129,N_9329);
and U13017 (N_13017,N_5419,N_5102);
and U13018 (N_13018,N_8299,N_8592);
or U13019 (N_13019,N_7268,N_5505);
or U13020 (N_13020,N_5604,N_6392);
xnor U13021 (N_13021,N_8179,N_7796);
nand U13022 (N_13022,N_5813,N_7760);
and U13023 (N_13023,N_6256,N_7774);
nor U13024 (N_13024,N_5853,N_5633);
nor U13025 (N_13025,N_9466,N_6680);
nor U13026 (N_13026,N_9593,N_9983);
nor U13027 (N_13027,N_9423,N_9312);
and U13028 (N_13028,N_5104,N_6198);
nor U13029 (N_13029,N_7749,N_9370);
nor U13030 (N_13030,N_8276,N_7337);
nand U13031 (N_13031,N_5642,N_6377);
and U13032 (N_13032,N_7659,N_6212);
nor U13033 (N_13033,N_7074,N_5654);
and U13034 (N_13034,N_7773,N_5787);
or U13035 (N_13035,N_5490,N_9239);
nor U13036 (N_13036,N_9121,N_7872);
and U13037 (N_13037,N_6447,N_8308);
nor U13038 (N_13038,N_7936,N_9169);
and U13039 (N_13039,N_6343,N_7828);
nor U13040 (N_13040,N_8722,N_9766);
nor U13041 (N_13041,N_7935,N_6197);
or U13042 (N_13042,N_5467,N_9088);
nand U13043 (N_13043,N_7048,N_8386);
nor U13044 (N_13044,N_6090,N_6571);
nor U13045 (N_13045,N_7767,N_6906);
or U13046 (N_13046,N_9327,N_5338);
or U13047 (N_13047,N_9813,N_9575);
or U13048 (N_13048,N_5968,N_6115);
nand U13049 (N_13049,N_7439,N_8161);
nor U13050 (N_13050,N_5141,N_9218);
or U13051 (N_13051,N_6451,N_5935);
and U13052 (N_13052,N_6990,N_9834);
nor U13053 (N_13053,N_7400,N_5600);
nor U13054 (N_13054,N_5220,N_8022);
and U13055 (N_13055,N_9299,N_9394);
and U13056 (N_13056,N_6843,N_6376);
and U13057 (N_13057,N_6993,N_9702);
or U13058 (N_13058,N_8261,N_6551);
and U13059 (N_13059,N_5687,N_8392);
nand U13060 (N_13060,N_8648,N_9330);
nor U13061 (N_13061,N_8834,N_6981);
nor U13062 (N_13062,N_9961,N_8113);
nand U13063 (N_13063,N_9160,N_7956);
nand U13064 (N_13064,N_7630,N_9975);
and U13065 (N_13065,N_6334,N_6220);
and U13066 (N_13066,N_7885,N_5502);
nand U13067 (N_13067,N_9727,N_6629);
nor U13068 (N_13068,N_8827,N_7471);
nand U13069 (N_13069,N_7267,N_5949);
nor U13070 (N_13070,N_9581,N_7533);
nand U13071 (N_13071,N_8433,N_9321);
or U13072 (N_13072,N_6643,N_7238);
and U13073 (N_13073,N_5562,N_8928);
and U13074 (N_13074,N_9868,N_8449);
nand U13075 (N_13075,N_7011,N_9838);
or U13076 (N_13076,N_8437,N_5963);
nor U13077 (N_13077,N_8442,N_5191);
nand U13078 (N_13078,N_6112,N_6344);
or U13079 (N_13079,N_6511,N_5988);
and U13080 (N_13080,N_5218,N_5387);
and U13081 (N_13081,N_9088,N_5758);
nor U13082 (N_13082,N_8442,N_6232);
or U13083 (N_13083,N_7479,N_8720);
nor U13084 (N_13084,N_5104,N_9278);
or U13085 (N_13085,N_8489,N_9067);
or U13086 (N_13086,N_5585,N_9467);
xor U13087 (N_13087,N_6594,N_6876);
and U13088 (N_13088,N_9565,N_6251);
nor U13089 (N_13089,N_6936,N_6305);
and U13090 (N_13090,N_8688,N_9612);
nor U13091 (N_13091,N_9158,N_8878);
or U13092 (N_13092,N_7148,N_6946);
and U13093 (N_13093,N_9912,N_5874);
nand U13094 (N_13094,N_7041,N_8460);
nand U13095 (N_13095,N_8301,N_6058);
and U13096 (N_13096,N_9442,N_6314);
nor U13097 (N_13097,N_9899,N_7360);
or U13098 (N_13098,N_7928,N_8898);
nand U13099 (N_13099,N_5920,N_7321);
or U13100 (N_13100,N_8511,N_8273);
nand U13101 (N_13101,N_9452,N_9008);
nor U13102 (N_13102,N_7859,N_6705);
nor U13103 (N_13103,N_7742,N_7691);
nor U13104 (N_13104,N_5113,N_5134);
or U13105 (N_13105,N_7262,N_5011);
or U13106 (N_13106,N_7411,N_7528);
nor U13107 (N_13107,N_6435,N_8038);
or U13108 (N_13108,N_9577,N_9801);
nor U13109 (N_13109,N_5483,N_6592);
nor U13110 (N_13110,N_9045,N_9281);
or U13111 (N_13111,N_5566,N_7591);
and U13112 (N_13112,N_9786,N_9324);
nor U13113 (N_13113,N_8452,N_5101);
nand U13114 (N_13114,N_7294,N_5251);
nand U13115 (N_13115,N_7456,N_9195);
and U13116 (N_13116,N_9993,N_5161);
nor U13117 (N_13117,N_5203,N_6009);
nor U13118 (N_13118,N_7694,N_6178);
or U13119 (N_13119,N_9965,N_9897);
or U13120 (N_13120,N_9126,N_9525);
nor U13121 (N_13121,N_6997,N_6274);
and U13122 (N_13122,N_5984,N_9142);
nand U13123 (N_13123,N_7640,N_8560);
nand U13124 (N_13124,N_9655,N_6715);
or U13125 (N_13125,N_8610,N_6430);
nor U13126 (N_13126,N_7143,N_8508);
nand U13127 (N_13127,N_5946,N_7370);
or U13128 (N_13128,N_7993,N_9021);
or U13129 (N_13129,N_8059,N_6500);
and U13130 (N_13130,N_9852,N_8366);
or U13131 (N_13131,N_8315,N_5288);
nand U13132 (N_13132,N_7331,N_6355);
or U13133 (N_13133,N_5153,N_7202);
nand U13134 (N_13134,N_5291,N_7096);
or U13135 (N_13135,N_7869,N_5109);
nand U13136 (N_13136,N_9483,N_5386);
nor U13137 (N_13137,N_7611,N_5528);
or U13138 (N_13138,N_8793,N_6085);
and U13139 (N_13139,N_8055,N_7912);
nand U13140 (N_13140,N_7775,N_7514);
nor U13141 (N_13141,N_9379,N_5065);
and U13142 (N_13142,N_9772,N_6532);
or U13143 (N_13143,N_6223,N_5159);
nor U13144 (N_13144,N_5512,N_8054);
nand U13145 (N_13145,N_6895,N_5374);
nand U13146 (N_13146,N_6790,N_8036);
xor U13147 (N_13147,N_6571,N_9619);
nand U13148 (N_13148,N_5164,N_5572);
or U13149 (N_13149,N_6311,N_9021);
nand U13150 (N_13150,N_7804,N_9074);
nor U13151 (N_13151,N_5607,N_7266);
nor U13152 (N_13152,N_5143,N_5675);
nor U13153 (N_13153,N_6378,N_6323);
nor U13154 (N_13154,N_9046,N_9411);
and U13155 (N_13155,N_5975,N_7894);
nand U13156 (N_13156,N_9231,N_9578);
or U13157 (N_13157,N_9779,N_5167);
nand U13158 (N_13158,N_9627,N_9533);
nand U13159 (N_13159,N_8445,N_6937);
nor U13160 (N_13160,N_6167,N_5515);
or U13161 (N_13161,N_8140,N_9823);
nand U13162 (N_13162,N_5667,N_6072);
or U13163 (N_13163,N_7804,N_5761);
and U13164 (N_13164,N_7278,N_8659);
or U13165 (N_13165,N_7886,N_8788);
and U13166 (N_13166,N_8497,N_6487);
and U13167 (N_13167,N_8592,N_6621);
nor U13168 (N_13168,N_7452,N_5038);
or U13169 (N_13169,N_9156,N_9606);
and U13170 (N_13170,N_7190,N_9517);
nor U13171 (N_13171,N_9570,N_9816);
nand U13172 (N_13172,N_7220,N_9134);
nand U13173 (N_13173,N_5999,N_5608);
nand U13174 (N_13174,N_5364,N_7748);
nor U13175 (N_13175,N_6049,N_8783);
or U13176 (N_13176,N_6456,N_5513);
and U13177 (N_13177,N_7112,N_7981);
and U13178 (N_13178,N_7013,N_6908);
nor U13179 (N_13179,N_5894,N_9874);
nor U13180 (N_13180,N_6497,N_6605);
nand U13181 (N_13181,N_5185,N_5654);
and U13182 (N_13182,N_9474,N_7010);
or U13183 (N_13183,N_7620,N_6808);
nor U13184 (N_13184,N_8693,N_5592);
nor U13185 (N_13185,N_6968,N_8664);
or U13186 (N_13186,N_8612,N_9669);
and U13187 (N_13187,N_5563,N_7064);
nand U13188 (N_13188,N_6530,N_5696);
nand U13189 (N_13189,N_5839,N_7161);
or U13190 (N_13190,N_7340,N_9763);
or U13191 (N_13191,N_9980,N_8032);
or U13192 (N_13192,N_8505,N_8651);
nor U13193 (N_13193,N_8160,N_5259);
and U13194 (N_13194,N_5342,N_5405);
nand U13195 (N_13195,N_9895,N_9651);
or U13196 (N_13196,N_5189,N_6740);
nand U13197 (N_13197,N_5359,N_9602);
nor U13198 (N_13198,N_6283,N_9479);
and U13199 (N_13199,N_6089,N_6816);
or U13200 (N_13200,N_8168,N_5275);
or U13201 (N_13201,N_5990,N_7600);
and U13202 (N_13202,N_8353,N_5685);
and U13203 (N_13203,N_9359,N_6161);
nor U13204 (N_13204,N_9490,N_7969);
and U13205 (N_13205,N_6619,N_8450);
or U13206 (N_13206,N_5840,N_8745);
and U13207 (N_13207,N_6145,N_8170);
nand U13208 (N_13208,N_7871,N_9279);
or U13209 (N_13209,N_9298,N_6984);
nand U13210 (N_13210,N_6313,N_5965);
and U13211 (N_13211,N_5943,N_8588);
nor U13212 (N_13212,N_6701,N_8803);
nand U13213 (N_13213,N_9463,N_9767);
or U13214 (N_13214,N_8230,N_7667);
nand U13215 (N_13215,N_6331,N_5043);
or U13216 (N_13216,N_7860,N_5122);
and U13217 (N_13217,N_5097,N_9185);
nor U13218 (N_13218,N_9959,N_5909);
nor U13219 (N_13219,N_7760,N_6044);
and U13220 (N_13220,N_7347,N_8584);
or U13221 (N_13221,N_6098,N_6116);
nand U13222 (N_13222,N_5893,N_8495);
or U13223 (N_13223,N_8067,N_7549);
or U13224 (N_13224,N_6400,N_8736);
nor U13225 (N_13225,N_5722,N_8003);
nor U13226 (N_13226,N_7492,N_9657);
and U13227 (N_13227,N_9185,N_5414);
nand U13228 (N_13228,N_6359,N_9693);
nor U13229 (N_13229,N_9078,N_5564);
or U13230 (N_13230,N_6913,N_7281);
and U13231 (N_13231,N_9742,N_8317);
or U13232 (N_13232,N_7039,N_6844);
or U13233 (N_13233,N_7252,N_6962);
nor U13234 (N_13234,N_8520,N_8556);
nand U13235 (N_13235,N_6561,N_5662);
and U13236 (N_13236,N_5518,N_9455);
nand U13237 (N_13237,N_9032,N_7166);
nor U13238 (N_13238,N_6500,N_9653);
and U13239 (N_13239,N_7578,N_8067);
and U13240 (N_13240,N_7570,N_9500);
nand U13241 (N_13241,N_9438,N_6758);
nor U13242 (N_13242,N_6296,N_8506);
or U13243 (N_13243,N_9923,N_7034);
nor U13244 (N_13244,N_7587,N_7605);
nand U13245 (N_13245,N_9813,N_8973);
nor U13246 (N_13246,N_5852,N_5862);
nor U13247 (N_13247,N_5578,N_6027);
nand U13248 (N_13248,N_5361,N_7675);
nand U13249 (N_13249,N_8308,N_7616);
nor U13250 (N_13250,N_8212,N_5399);
nor U13251 (N_13251,N_8348,N_6237);
and U13252 (N_13252,N_5203,N_6210);
nor U13253 (N_13253,N_9407,N_9041);
and U13254 (N_13254,N_6157,N_5671);
nor U13255 (N_13255,N_8167,N_8825);
nand U13256 (N_13256,N_9679,N_8325);
or U13257 (N_13257,N_8473,N_6626);
nand U13258 (N_13258,N_7628,N_6021);
and U13259 (N_13259,N_8827,N_8202);
nor U13260 (N_13260,N_5979,N_8928);
nand U13261 (N_13261,N_6374,N_7089);
xnor U13262 (N_13262,N_9937,N_8749);
and U13263 (N_13263,N_5784,N_5542);
and U13264 (N_13264,N_8630,N_8539);
or U13265 (N_13265,N_7555,N_9561);
nand U13266 (N_13266,N_8592,N_6599);
nor U13267 (N_13267,N_6503,N_6844);
and U13268 (N_13268,N_9241,N_6972);
nor U13269 (N_13269,N_7060,N_9849);
nor U13270 (N_13270,N_6965,N_5249);
or U13271 (N_13271,N_5920,N_6034);
nor U13272 (N_13272,N_7721,N_7693);
nand U13273 (N_13273,N_8723,N_8993);
nor U13274 (N_13274,N_7497,N_8083);
or U13275 (N_13275,N_5051,N_6653);
nand U13276 (N_13276,N_5284,N_8269);
nand U13277 (N_13277,N_7636,N_6809);
nor U13278 (N_13278,N_5381,N_5799);
xnor U13279 (N_13279,N_9284,N_9565);
and U13280 (N_13280,N_8256,N_6479);
nand U13281 (N_13281,N_8219,N_8004);
or U13282 (N_13282,N_9486,N_8425);
and U13283 (N_13283,N_5743,N_9943);
nor U13284 (N_13284,N_8019,N_7731);
nor U13285 (N_13285,N_9745,N_6693);
nor U13286 (N_13286,N_8354,N_5640);
or U13287 (N_13287,N_8224,N_5258);
nor U13288 (N_13288,N_7185,N_5748);
nand U13289 (N_13289,N_8741,N_7840);
nor U13290 (N_13290,N_6648,N_8562);
nor U13291 (N_13291,N_9811,N_6802);
nor U13292 (N_13292,N_8684,N_6733);
nor U13293 (N_13293,N_5303,N_5456);
nand U13294 (N_13294,N_5777,N_6216);
and U13295 (N_13295,N_9010,N_5954);
and U13296 (N_13296,N_8916,N_9597);
nor U13297 (N_13297,N_6516,N_7930);
and U13298 (N_13298,N_9287,N_9854);
or U13299 (N_13299,N_8011,N_6865);
nor U13300 (N_13300,N_5074,N_6804);
and U13301 (N_13301,N_8605,N_8204);
and U13302 (N_13302,N_6688,N_9232);
or U13303 (N_13303,N_7858,N_9577);
and U13304 (N_13304,N_8284,N_7063);
nand U13305 (N_13305,N_6706,N_8624);
nand U13306 (N_13306,N_9289,N_6814);
nor U13307 (N_13307,N_6122,N_9541);
nand U13308 (N_13308,N_7491,N_8740);
and U13309 (N_13309,N_5474,N_9074);
or U13310 (N_13310,N_5748,N_7509);
and U13311 (N_13311,N_8886,N_7045);
and U13312 (N_13312,N_5345,N_5524);
and U13313 (N_13313,N_5474,N_8743);
or U13314 (N_13314,N_6353,N_7498);
and U13315 (N_13315,N_8750,N_5301);
xnor U13316 (N_13316,N_9189,N_5110);
or U13317 (N_13317,N_7150,N_6768);
or U13318 (N_13318,N_6515,N_5439);
nand U13319 (N_13319,N_7357,N_8284);
nand U13320 (N_13320,N_5133,N_5893);
or U13321 (N_13321,N_6332,N_7807);
or U13322 (N_13322,N_6945,N_7560);
nor U13323 (N_13323,N_9127,N_9069);
nor U13324 (N_13324,N_9832,N_9011);
and U13325 (N_13325,N_6782,N_9951);
and U13326 (N_13326,N_7556,N_8560);
nand U13327 (N_13327,N_8327,N_5510);
and U13328 (N_13328,N_6779,N_5287);
and U13329 (N_13329,N_6386,N_9640);
nand U13330 (N_13330,N_5372,N_6561);
nand U13331 (N_13331,N_8967,N_6876);
nand U13332 (N_13332,N_9719,N_9772);
and U13333 (N_13333,N_7986,N_8906);
nor U13334 (N_13334,N_7155,N_5708);
nor U13335 (N_13335,N_7400,N_7362);
nor U13336 (N_13336,N_7649,N_7960);
and U13337 (N_13337,N_5628,N_9389);
and U13338 (N_13338,N_6541,N_8475);
and U13339 (N_13339,N_9073,N_5777);
and U13340 (N_13340,N_7390,N_7020);
or U13341 (N_13341,N_8551,N_8346);
nand U13342 (N_13342,N_5479,N_5549);
nand U13343 (N_13343,N_6524,N_8609);
and U13344 (N_13344,N_9965,N_6142);
and U13345 (N_13345,N_8338,N_8997);
nor U13346 (N_13346,N_9463,N_9469);
nand U13347 (N_13347,N_9928,N_8083);
and U13348 (N_13348,N_6576,N_7541);
and U13349 (N_13349,N_9668,N_8930);
and U13350 (N_13350,N_7883,N_5032);
nand U13351 (N_13351,N_9816,N_5417);
nor U13352 (N_13352,N_7182,N_7283);
nor U13353 (N_13353,N_6813,N_5941);
and U13354 (N_13354,N_5908,N_8338);
nor U13355 (N_13355,N_5940,N_9480);
nand U13356 (N_13356,N_6793,N_8615);
and U13357 (N_13357,N_6805,N_5229);
or U13358 (N_13358,N_9007,N_8253);
or U13359 (N_13359,N_8182,N_9693);
nor U13360 (N_13360,N_6956,N_6424);
nand U13361 (N_13361,N_6678,N_6113);
or U13362 (N_13362,N_5767,N_6123);
nand U13363 (N_13363,N_6616,N_9779);
nor U13364 (N_13364,N_5737,N_5981);
and U13365 (N_13365,N_8050,N_7510);
nor U13366 (N_13366,N_5659,N_6055);
or U13367 (N_13367,N_8845,N_7992);
nand U13368 (N_13368,N_8572,N_5533);
nor U13369 (N_13369,N_5836,N_6586);
nand U13370 (N_13370,N_5506,N_5575);
and U13371 (N_13371,N_5166,N_7944);
nand U13372 (N_13372,N_6861,N_8657);
or U13373 (N_13373,N_5589,N_9493);
nor U13374 (N_13374,N_9263,N_6415);
nor U13375 (N_13375,N_9906,N_6423);
and U13376 (N_13376,N_5724,N_6400);
nand U13377 (N_13377,N_6080,N_6749);
or U13378 (N_13378,N_9563,N_7387);
nand U13379 (N_13379,N_8050,N_6522);
nand U13380 (N_13380,N_7013,N_6318);
and U13381 (N_13381,N_5407,N_9206);
nand U13382 (N_13382,N_7360,N_8306);
nor U13383 (N_13383,N_8616,N_5378);
nor U13384 (N_13384,N_9520,N_7487);
or U13385 (N_13385,N_5573,N_7577);
nand U13386 (N_13386,N_8479,N_5042);
or U13387 (N_13387,N_8464,N_8706);
nor U13388 (N_13388,N_7605,N_9786);
nand U13389 (N_13389,N_5295,N_7764);
nor U13390 (N_13390,N_5189,N_8529);
and U13391 (N_13391,N_9456,N_5681);
or U13392 (N_13392,N_5593,N_8145);
or U13393 (N_13393,N_7061,N_9487);
and U13394 (N_13394,N_9258,N_5364);
or U13395 (N_13395,N_9483,N_8569);
nand U13396 (N_13396,N_8948,N_8515);
nor U13397 (N_13397,N_6164,N_6970);
or U13398 (N_13398,N_8476,N_7810);
and U13399 (N_13399,N_7055,N_8977);
nand U13400 (N_13400,N_9465,N_8969);
or U13401 (N_13401,N_9700,N_9803);
nor U13402 (N_13402,N_5531,N_5042);
and U13403 (N_13403,N_9065,N_9813);
nand U13404 (N_13404,N_8805,N_7414);
and U13405 (N_13405,N_7672,N_6809);
xor U13406 (N_13406,N_8497,N_5846);
nand U13407 (N_13407,N_7661,N_7489);
and U13408 (N_13408,N_6930,N_6073);
nand U13409 (N_13409,N_6043,N_9898);
and U13410 (N_13410,N_9565,N_9450);
or U13411 (N_13411,N_8754,N_9592);
or U13412 (N_13412,N_9740,N_8919);
nor U13413 (N_13413,N_7006,N_9016);
nor U13414 (N_13414,N_8841,N_7317);
nor U13415 (N_13415,N_6435,N_9343);
and U13416 (N_13416,N_6314,N_8014);
nor U13417 (N_13417,N_7844,N_7602);
nor U13418 (N_13418,N_6351,N_8657);
or U13419 (N_13419,N_7097,N_7705);
nand U13420 (N_13420,N_7644,N_5437);
and U13421 (N_13421,N_6199,N_7517);
nand U13422 (N_13422,N_7513,N_6608);
and U13423 (N_13423,N_8914,N_7086);
or U13424 (N_13424,N_8522,N_9535);
and U13425 (N_13425,N_5391,N_7693);
nand U13426 (N_13426,N_6852,N_6714);
nand U13427 (N_13427,N_8120,N_7216);
nand U13428 (N_13428,N_7906,N_7210);
nand U13429 (N_13429,N_9909,N_8133);
xor U13430 (N_13430,N_9174,N_5062);
nor U13431 (N_13431,N_7583,N_8666);
and U13432 (N_13432,N_9535,N_7831);
and U13433 (N_13433,N_8733,N_8295);
nand U13434 (N_13434,N_9035,N_8069);
nor U13435 (N_13435,N_5456,N_5381);
xnor U13436 (N_13436,N_5178,N_6750);
or U13437 (N_13437,N_9388,N_7651);
or U13438 (N_13438,N_9847,N_5535);
and U13439 (N_13439,N_9217,N_7077);
nand U13440 (N_13440,N_7494,N_5815);
nor U13441 (N_13441,N_5084,N_5286);
or U13442 (N_13442,N_9871,N_5524);
nand U13443 (N_13443,N_9025,N_8707);
and U13444 (N_13444,N_6146,N_5395);
xor U13445 (N_13445,N_8949,N_5158);
nor U13446 (N_13446,N_7979,N_6593);
or U13447 (N_13447,N_6952,N_8069);
nand U13448 (N_13448,N_7441,N_6270);
nand U13449 (N_13449,N_5101,N_7699);
nand U13450 (N_13450,N_8969,N_8012);
nor U13451 (N_13451,N_5504,N_8779);
and U13452 (N_13452,N_8494,N_9206);
nand U13453 (N_13453,N_9104,N_5201);
or U13454 (N_13454,N_9725,N_9400);
or U13455 (N_13455,N_6759,N_6439);
nor U13456 (N_13456,N_6811,N_7409);
or U13457 (N_13457,N_6373,N_6917);
or U13458 (N_13458,N_9663,N_6829);
or U13459 (N_13459,N_6742,N_7989);
nand U13460 (N_13460,N_8623,N_5028);
and U13461 (N_13461,N_8147,N_5816);
and U13462 (N_13462,N_8843,N_6955);
or U13463 (N_13463,N_9655,N_5002);
and U13464 (N_13464,N_6775,N_5402);
nand U13465 (N_13465,N_6075,N_9881);
nand U13466 (N_13466,N_9188,N_5350);
or U13467 (N_13467,N_7713,N_9694);
or U13468 (N_13468,N_8983,N_9043);
nor U13469 (N_13469,N_9232,N_6298);
or U13470 (N_13470,N_7047,N_6081);
or U13471 (N_13471,N_7804,N_7669);
or U13472 (N_13472,N_6223,N_8363);
nor U13473 (N_13473,N_9750,N_7393);
or U13474 (N_13474,N_9810,N_6855);
or U13475 (N_13475,N_6875,N_9630);
or U13476 (N_13476,N_7660,N_7674);
and U13477 (N_13477,N_7446,N_6942);
nor U13478 (N_13478,N_8679,N_6252);
and U13479 (N_13479,N_8097,N_6438);
or U13480 (N_13480,N_8882,N_8477);
and U13481 (N_13481,N_5680,N_9549);
and U13482 (N_13482,N_6564,N_5588);
or U13483 (N_13483,N_6062,N_9584);
nand U13484 (N_13484,N_8081,N_5480);
nor U13485 (N_13485,N_7977,N_9926);
nand U13486 (N_13486,N_6557,N_6491);
or U13487 (N_13487,N_9160,N_9118);
and U13488 (N_13488,N_5694,N_7570);
or U13489 (N_13489,N_9833,N_7159);
nand U13490 (N_13490,N_6057,N_7625);
or U13491 (N_13491,N_5895,N_6935);
or U13492 (N_13492,N_8934,N_6660);
or U13493 (N_13493,N_5271,N_7409);
nor U13494 (N_13494,N_8061,N_5810);
or U13495 (N_13495,N_9082,N_9185);
nand U13496 (N_13496,N_7778,N_7797);
and U13497 (N_13497,N_7401,N_7375);
nor U13498 (N_13498,N_8876,N_8965);
nor U13499 (N_13499,N_6200,N_6294);
nor U13500 (N_13500,N_6605,N_9251);
nor U13501 (N_13501,N_8937,N_8156);
nor U13502 (N_13502,N_8942,N_5544);
and U13503 (N_13503,N_9363,N_5126);
and U13504 (N_13504,N_7438,N_9469);
xor U13505 (N_13505,N_5955,N_7185);
or U13506 (N_13506,N_9424,N_7442);
nor U13507 (N_13507,N_6553,N_5542);
nand U13508 (N_13508,N_5998,N_8788);
nand U13509 (N_13509,N_8186,N_7163);
nor U13510 (N_13510,N_8043,N_5084);
and U13511 (N_13511,N_9402,N_7246);
and U13512 (N_13512,N_5707,N_8522);
and U13513 (N_13513,N_6710,N_5493);
and U13514 (N_13514,N_6278,N_6295);
nand U13515 (N_13515,N_9575,N_5117);
nor U13516 (N_13516,N_9279,N_8453);
nor U13517 (N_13517,N_6267,N_6714);
nor U13518 (N_13518,N_6546,N_9757);
or U13519 (N_13519,N_9657,N_5723);
or U13520 (N_13520,N_7800,N_5921);
nand U13521 (N_13521,N_8718,N_7531);
or U13522 (N_13522,N_7840,N_5523);
nand U13523 (N_13523,N_8343,N_8905);
and U13524 (N_13524,N_9808,N_7687);
nor U13525 (N_13525,N_8982,N_6415);
or U13526 (N_13526,N_9599,N_9392);
or U13527 (N_13527,N_8885,N_9729);
nor U13528 (N_13528,N_6156,N_9684);
nor U13529 (N_13529,N_5042,N_6599);
or U13530 (N_13530,N_5117,N_6314);
nor U13531 (N_13531,N_9094,N_7440);
and U13532 (N_13532,N_9645,N_5814);
and U13533 (N_13533,N_6793,N_9088);
and U13534 (N_13534,N_7175,N_8013);
nor U13535 (N_13535,N_7554,N_9568);
and U13536 (N_13536,N_9118,N_7672);
nand U13537 (N_13537,N_5548,N_6570);
and U13538 (N_13538,N_9069,N_5948);
nand U13539 (N_13539,N_8446,N_8963);
nand U13540 (N_13540,N_7551,N_5278);
and U13541 (N_13541,N_8038,N_9653);
or U13542 (N_13542,N_7328,N_7633);
or U13543 (N_13543,N_7020,N_5142);
and U13544 (N_13544,N_7044,N_6615);
nand U13545 (N_13545,N_9462,N_7553);
and U13546 (N_13546,N_6264,N_8977);
or U13547 (N_13547,N_7332,N_9697);
nor U13548 (N_13548,N_7411,N_8542);
nand U13549 (N_13549,N_8888,N_5121);
or U13550 (N_13550,N_8924,N_8384);
or U13551 (N_13551,N_5158,N_7195);
or U13552 (N_13552,N_5316,N_8270);
or U13553 (N_13553,N_8030,N_6415);
or U13554 (N_13554,N_5175,N_5684);
nor U13555 (N_13555,N_5442,N_7613);
nor U13556 (N_13556,N_9056,N_6137);
and U13557 (N_13557,N_7694,N_8655);
and U13558 (N_13558,N_7115,N_8851);
and U13559 (N_13559,N_6497,N_9884);
and U13560 (N_13560,N_8308,N_8649);
nand U13561 (N_13561,N_9033,N_9265);
xor U13562 (N_13562,N_8594,N_7158);
nor U13563 (N_13563,N_9487,N_8853);
nand U13564 (N_13564,N_8483,N_7308);
or U13565 (N_13565,N_6158,N_5159);
nand U13566 (N_13566,N_8953,N_8483);
nor U13567 (N_13567,N_9691,N_6933);
nand U13568 (N_13568,N_9210,N_6841);
or U13569 (N_13569,N_6952,N_8015);
nor U13570 (N_13570,N_9132,N_5394);
nand U13571 (N_13571,N_6029,N_8528);
nand U13572 (N_13572,N_6620,N_8521);
and U13573 (N_13573,N_7171,N_6842);
nor U13574 (N_13574,N_6238,N_5055);
nor U13575 (N_13575,N_7366,N_6573);
nand U13576 (N_13576,N_8889,N_6587);
or U13577 (N_13577,N_8999,N_5349);
or U13578 (N_13578,N_8575,N_9763);
and U13579 (N_13579,N_7856,N_6717);
and U13580 (N_13580,N_6875,N_8794);
xnor U13581 (N_13581,N_6798,N_5041);
and U13582 (N_13582,N_9426,N_5680);
nor U13583 (N_13583,N_6733,N_9427);
nand U13584 (N_13584,N_8192,N_5446);
nand U13585 (N_13585,N_6438,N_7276);
nand U13586 (N_13586,N_9604,N_6489);
nand U13587 (N_13587,N_8072,N_8143);
nand U13588 (N_13588,N_8906,N_7797);
or U13589 (N_13589,N_8853,N_8221);
nand U13590 (N_13590,N_6455,N_6811);
and U13591 (N_13591,N_8072,N_5756);
nor U13592 (N_13592,N_5013,N_5368);
or U13593 (N_13593,N_8994,N_5775);
nand U13594 (N_13594,N_9934,N_8152);
nand U13595 (N_13595,N_5617,N_5046);
nand U13596 (N_13596,N_8134,N_9491);
nand U13597 (N_13597,N_7659,N_8380);
or U13598 (N_13598,N_9091,N_9462);
or U13599 (N_13599,N_9252,N_7310);
nand U13600 (N_13600,N_8390,N_8695);
nor U13601 (N_13601,N_7456,N_7005);
and U13602 (N_13602,N_5578,N_9112);
nor U13603 (N_13603,N_5720,N_5469);
nor U13604 (N_13604,N_5310,N_7964);
and U13605 (N_13605,N_5832,N_7110);
nor U13606 (N_13606,N_7302,N_6153);
and U13607 (N_13607,N_5235,N_8956);
nand U13608 (N_13608,N_8040,N_8949);
nor U13609 (N_13609,N_7315,N_6179);
or U13610 (N_13610,N_6548,N_8796);
nor U13611 (N_13611,N_6893,N_8669);
nand U13612 (N_13612,N_8326,N_5421);
nand U13613 (N_13613,N_8313,N_7012);
and U13614 (N_13614,N_6862,N_8227);
nand U13615 (N_13615,N_6040,N_5545);
nor U13616 (N_13616,N_5132,N_8015);
nor U13617 (N_13617,N_7212,N_7957);
nor U13618 (N_13618,N_7048,N_5963);
nand U13619 (N_13619,N_5318,N_5658);
or U13620 (N_13620,N_5683,N_9466);
nor U13621 (N_13621,N_8565,N_5806);
nor U13622 (N_13622,N_9235,N_7652);
and U13623 (N_13623,N_7330,N_9984);
nand U13624 (N_13624,N_6063,N_9584);
nand U13625 (N_13625,N_5171,N_9575);
xnor U13626 (N_13626,N_7358,N_8987);
or U13627 (N_13627,N_9236,N_5518);
nand U13628 (N_13628,N_6956,N_8464);
nor U13629 (N_13629,N_8795,N_7421);
or U13630 (N_13630,N_7789,N_7580);
and U13631 (N_13631,N_5033,N_7468);
or U13632 (N_13632,N_8902,N_8317);
and U13633 (N_13633,N_8269,N_5397);
and U13634 (N_13634,N_5003,N_8439);
and U13635 (N_13635,N_7671,N_9530);
and U13636 (N_13636,N_6340,N_5209);
and U13637 (N_13637,N_6542,N_7008);
or U13638 (N_13638,N_8042,N_6508);
and U13639 (N_13639,N_9727,N_9132);
nand U13640 (N_13640,N_9846,N_9466);
and U13641 (N_13641,N_7417,N_8486);
nand U13642 (N_13642,N_8316,N_9705);
and U13643 (N_13643,N_6665,N_5499);
nor U13644 (N_13644,N_7653,N_5336);
or U13645 (N_13645,N_7498,N_9896);
nor U13646 (N_13646,N_6542,N_6622);
and U13647 (N_13647,N_9020,N_9526);
and U13648 (N_13648,N_9937,N_7662);
and U13649 (N_13649,N_5590,N_6961);
and U13650 (N_13650,N_5223,N_5844);
and U13651 (N_13651,N_9476,N_9938);
nand U13652 (N_13652,N_7550,N_7524);
nor U13653 (N_13653,N_9420,N_8960);
nand U13654 (N_13654,N_8517,N_9046);
nand U13655 (N_13655,N_7866,N_8292);
or U13656 (N_13656,N_7702,N_6200);
or U13657 (N_13657,N_7304,N_9237);
or U13658 (N_13658,N_8116,N_7037);
nor U13659 (N_13659,N_7884,N_6864);
nor U13660 (N_13660,N_7120,N_7782);
nor U13661 (N_13661,N_8362,N_8981);
nor U13662 (N_13662,N_9737,N_6408);
nor U13663 (N_13663,N_9348,N_9160);
or U13664 (N_13664,N_9173,N_7744);
nor U13665 (N_13665,N_5646,N_6688);
or U13666 (N_13666,N_8351,N_9364);
or U13667 (N_13667,N_6406,N_8275);
or U13668 (N_13668,N_6473,N_5437);
nor U13669 (N_13669,N_7272,N_7300);
nor U13670 (N_13670,N_9160,N_5933);
or U13671 (N_13671,N_6452,N_7506);
or U13672 (N_13672,N_9096,N_6792);
nand U13673 (N_13673,N_8059,N_5066);
or U13674 (N_13674,N_9309,N_5966);
and U13675 (N_13675,N_6389,N_9321);
nor U13676 (N_13676,N_5490,N_5804);
and U13677 (N_13677,N_5482,N_9148);
and U13678 (N_13678,N_9724,N_5722);
nor U13679 (N_13679,N_5877,N_5364);
or U13680 (N_13680,N_5152,N_6669);
nor U13681 (N_13681,N_7023,N_5200);
or U13682 (N_13682,N_5135,N_6896);
nor U13683 (N_13683,N_5176,N_7353);
and U13684 (N_13684,N_6982,N_6657);
nor U13685 (N_13685,N_6009,N_5230);
nand U13686 (N_13686,N_9289,N_6112);
nand U13687 (N_13687,N_8327,N_5957);
and U13688 (N_13688,N_8689,N_6869);
or U13689 (N_13689,N_5607,N_6726);
and U13690 (N_13690,N_9777,N_6833);
nor U13691 (N_13691,N_8270,N_8813);
nor U13692 (N_13692,N_9701,N_9803);
and U13693 (N_13693,N_8611,N_6194);
nor U13694 (N_13694,N_5866,N_7427);
or U13695 (N_13695,N_7744,N_6707);
nor U13696 (N_13696,N_9216,N_8504);
nor U13697 (N_13697,N_9653,N_7503);
or U13698 (N_13698,N_7513,N_8211);
or U13699 (N_13699,N_7486,N_9262);
and U13700 (N_13700,N_6862,N_5959);
or U13701 (N_13701,N_9424,N_5731);
nand U13702 (N_13702,N_9115,N_7076);
nand U13703 (N_13703,N_8933,N_5362);
nor U13704 (N_13704,N_5595,N_9528);
and U13705 (N_13705,N_8020,N_5649);
or U13706 (N_13706,N_9632,N_7431);
and U13707 (N_13707,N_8944,N_5782);
nand U13708 (N_13708,N_7708,N_5523);
and U13709 (N_13709,N_7355,N_9434);
or U13710 (N_13710,N_8391,N_9396);
or U13711 (N_13711,N_8379,N_9687);
nor U13712 (N_13712,N_6160,N_8177);
or U13713 (N_13713,N_5172,N_9131);
nand U13714 (N_13714,N_5797,N_6746);
or U13715 (N_13715,N_6713,N_8543);
and U13716 (N_13716,N_7565,N_6883);
nor U13717 (N_13717,N_6782,N_7856);
and U13718 (N_13718,N_6383,N_5716);
or U13719 (N_13719,N_8063,N_7264);
nor U13720 (N_13720,N_7576,N_9291);
nand U13721 (N_13721,N_9356,N_6745);
or U13722 (N_13722,N_7163,N_7268);
and U13723 (N_13723,N_9402,N_7148);
and U13724 (N_13724,N_8135,N_5206);
and U13725 (N_13725,N_5201,N_8529);
or U13726 (N_13726,N_7492,N_9971);
nand U13727 (N_13727,N_6243,N_9783);
and U13728 (N_13728,N_9759,N_6878);
nor U13729 (N_13729,N_9112,N_7818);
and U13730 (N_13730,N_5844,N_9631);
nor U13731 (N_13731,N_7977,N_9243);
nand U13732 (N_13732,N_5980,N_6015);
xnor U13733 (N_13733,N_5440,N_6875);
nor U13734 (N_13734,N_6288,N_9224);
nand U13735 (N_13735,N_8404,N_6842);
xor U13736 (N_13736,N_6564,N_5229);
nand U13737 (N_13737,N_9345,N_6361);
nand U13738 (N_13738,N_5654,N_8215);
and U13739 (N_13739,N_5637,N_6742);
and U13740 (N_13740,N_6399,N_8964);
or U13741 (N_13741,N_7477,N_8656);
nand U13742 (N_13742,N_5694,N_9384);
and U13743 (N_13743,N_9600,N_5607);
nor U13744 (N_13744,N_5102,N_8166);
nor U13745 (N_13745,N_7374,N_7932);
or U13746 (N_13746,N_5302,N_9441);
or U13747 (N_13747,N_8492,N_8535);
nand U13748 (N_13748,N_7631,N_7770);
and U13749 (N_13749,N_5857,N_9001);
and U13750 (N_13750,N_5839,N_9366);
and U13751 (N_13751,N_5634,N_8932);
or U13752 (N_13752,N_9689,N_8550);
nand U13753 (N_13753,N_6571,N_5152);
nor U13754 (N_13754,N_7456,N_7855);
nor U13755 (N_13755,N_8118,N_8588);
nand U13756 (N_13756,N_6155,N_9015);
or U13757 (N_13757,N_8156,N_7584);
or U13758 (N_13758,N_8735,N_5107);
nor U13759 (N_13759,N_9651,N_9993);
or U13760 (N_13760,N_6090,N_8637);
nand U13761 (N_13761,N_8955,N_8052);
nor U13762 (N_13762,N_6320,N_6120);
or U13763 (N_13763,N_5627,N_9756);
or U13764 (N_13764,N_5843,N_7688);
nand U13765 (N_13765,N_7549,N_7237);
nor U13766 (N_13766,N_9876,N_6275);
and U13767 (N_13767,N_9190,N_5775);
nor U13768 (N_13768,N_7665,N_9872);
and U13769 (N_13769,N_8916,N_7916);
nor U13770 (N_13770,N_6193,N_9131);
nand U13771 (N_13771,N_9257,N_5650);
nand U13772 (N_13772,N_6154,N_9948);
nor U13773 (N_13773,N_6470,N_5995);
or U13774 (N_13774,N_7587,N_6697);
nand U13775 (N_13775,N_9417,N_7063);
and U13776 (N_13776,N_9001,N_8355);
and U13777 (N_13777,N_8298,N_8023);
or U13778 (N_13778,N_7722,N_8374);
and U13779 (N_13779,N_9431,N_9667);
and U13780 (N_13780,N_6594,N_5004);
and U13781 (N_13781,N_9520,N_9880);
nor U13782 (N_13782,N_8880,N_6026);
nand U13783 (N_13783,N_6239,N_9881);
nand U13784 (N_13784,N_7729,N_9368);
nand U13785 (N_13785,N_6064,N_7944);
or U13786 (N_13786,N_6750,N_9519);
nand U13787 (N_13787,N_7793,N_5944);
and U13788 (N_13788,N_6194,N_7194);
and U13789 (N_13789,N_5906,N_9053);
or U13790 (N_13790,N_5266,N_8764);
nor U13791 (N_13791,N_8143,N_9233);
or U13792 (N_13792,N_9347,N_6612);
nand U13793 (N_13793,N_7705,N_8652);
nand U13794 (N_13794,N_8903,N_8070);
or U13795 (N_13795,N_9631,N_7521);
xor U13796 (N_13796,N_5513,N_8207);
nor U13797 (N_13797,N_7379,N_6897);
nand U13798 (N_13798,N_8203,N_7107);
and U13799 (N_13799,N_8100,N_6528);
nor U13800 (N_13800,N_9260,N_7018);
or U13801 (N_13801,N_7150,N_5386);
nor U13802 (N_13802,N_7244,N_5289);
or U13803 (N_13803,N_7079,N_9949);
or U13804 (N_13804,N_6833,N_9577);
or U13805 (N_13805,N_5921,N_8526);
nor U13806 (N_13806,N_8507,N_8578);
and U13807 (N_13807,N_7102,N_5491);
or U13808 (N_13808,N_6465,N_8053);
or U13809 (N_13809,N_6111,N_5192);
nand U13810 (N_13810,N_6910,N_6159);
nand U13811 (N_13811,N_5329,N_5528);
and U13812 (N_13812,N_8282,N_6039);
or U13813 (N_13813,N_6657,N_6781);
and U13814 (N_13814,N_8391,N_9791);
nor U13815 (N_13815,N_6361,N_6717);
nor U13816 (N_13816,N_9346,N_6089);
or U13817 (N_13817,N_5142,N_8822);
and U13818 (N_13818,N_6493,N_8743);
or U13819 (N_13819,N_6673,N_5885);
or U13820 (N_13820,N_8535,N_6400);
and U13821 (N_13821,N_5009,N_7868);
and U13822 (N_13822,N_8015,N_6093);
or U13823 (N_13823,N_5985,N_6916);
nor U13824 (N_13824,N_5020,N_9390);
nor U13825 (N_13825,N_5616,N_5085);
nand U13826 (N_13826,N_7640,N_5787);
and U13827 (N_13827,N_8656,N_8956);
nor U13828 (N_13828,N_7345,N_7737);
or U13829 (N_13829,N_9461,N_6020);
nand U13830 (N_13830,N_6424,N_5619);
nor U13831 (N_13831,N_8177,N_6558);
nor U13832 (N_13832,N_8300,N_9558);
nand U13833 (N_13833,N_7877,N_6050);
nand U13834 (N_13834,N_7050,N_7782);
or U13835 (N_13835,N_9535,N_7947);
nor U13836 (N_13836,N_6291,N_7615);
and U13837 (N_13837,N_7665,N_6758);
nor U13838 (N_13838,N_8588,N_9964);
xnor U13839 (N_13839,N_7319,N_8739);
and U13840 (N_13840,N_9736,N_6243);
and U13841 (N_13841,N_9478,N_5356);
or U13842 (N_13842,N_5853,N_8081);
nor U13843 (N_13843,N_5822,N_5728);
and U13844 (N_13844,N_8954,N_6151);
or U13845 (N_13845,N_6501,N_8388);
nor U13846 (N_13846,N_6696,N_9995);
nor U13847 (N_13847,N_5278,N_9600);
nand U13848 (N_13848,N_9066,N_9334);
nor U13849 (N_13849,N_9323,N_7950);
or U13850 (N_13850,N_5626,N_6165);
nor U13851 (N_13851,N_6627,N_8477);
nand U13852 (N_13852,N_7243,N_8826);
or U13853 (N_13853,N_9271,N_7904);
and U13854 (N_13854,N_6970,N_9280);
or U13855 (N_13855,N_7195,N_9440);
nand U13856 (N_13856,N_8520,N_6377);
nor U13857 (N_13857,N_8924,N_5002);
and U13858 (N_13858,N_7286,N_9137);
or U13859 (N_13859,N_9564,N_7005);
or U13860 (N_13860,N_7178,N_5023);
and U13861 (N_13861,N_6471,N_8254);
and U13862 (N_13862,N_6494,N_6039);
or U13863 (N_13863,N_9147,N_5036);
and U13864 (N_13864,N_6617,N_7016);
and U13865 (N_13865,N_8105,N_7536);
and U13866 (N_13866,N_9360,N_6243);
nor U13867 (N_13867,N_7864,N_8278);
or U13868 (N_13868,N_8045,N_5121);
or U13869 (N_13869,N_8868,N_7234);
or U13870 (N_13870,N_9628,N_8203);
nand U13871 (N_13871,N_7364,N_9960);
nor U13872 (N_13872,N_9510,N_6226);
nor U13873 (N_13873,N_6302,N_8577);
nor U13874 (N_13874,N_8977,N_6365);
nor U13875 (N_13875,N_7177,N_8452);
nand U13876 (N_13876,N_7591,N_9001);
and U13877 (N_13877,N_6144,N_8874);
and U13878 (N_13878,N_9316,N_7466);
or U13879 (N_13879,N_6031,N_9100);
nor U13880 (N_13880,N_8364,N_6757);
nor U13881 (N_13881,N_6097,N_9707);
and U13882 (N_13882,N_9431,N_9424);
and U13883 (N_13883,N_6117,N_9970);
and U13884 (N_13884,N_5775,N_7436);
nand U13885 (N_13885,N_8061,N_9331);
and U13886 (N_13886,N_8283,N_7179);
nand U13887 (N_13887,N_5220,N_6517);
nor U13888 (N_13888,N_5959,N_6663);
or U13889 (N_13889,N_9499,N_5545);
nor U13890 (N_13890,N_7951,N_9779);
or U13891 (N_13891,N_6052,N_9316);
and U13892 (N_13892,N_7464,N_5041);
nor U13893 (N_13893,N_9456,N_9165);
and U13894 (N_13894,N_5262,N_5208);
or U13895 (N_13895,N_8284,N_9505);
or U13896 (N_13896,N_7171,N_5108);
and U13897 (N_13897,N_6609,N_9190);
and U13898 (N_13898,N_8849,N_7562);
nor U13899 (N_13899,N_8000,N_5579);
nand U13900 (N_13900,N_7597,N_5522);
or U13901 (N_13901,N_8897,N_8340);
nand U13902 (N_13902,N_6777,N_9866);
nand U13903 (N_13903,N_9458,N_7570);
nor U13904 (N_13904,N_9482,N_7617);
or U13905 (N_13905,N_9272,N_8703);
and U13906 (N_13906,N_6516,N_7826);
nand U13907 (N_13907,N_5047,N_7647);
nand U13908 (N_13908,N_5687,N_5376);
and U13909 (N_13909,N_8453,N_6138);
xor U13910 (N_13910,N_9566,N_9286);
nor U13911 (N_13911,N_5671,N_9652);
nor U13912 (N_13912,N_8104,N_9810);
and U13913 (N_13913,N_6250,N_7288);
and U13914 (N_13914,N_5992,N_9730);
or U13915 (N_13915,N_9799,N_7416);
or U13916 (N_13916,N_7854,N_6935);
nand U13917 (N_13917,N_6757,N_5883);
nor U13918 (N_13918,N_8483,N_5828);
nor U13919 (N_13919,N_7174,N_8973);
nor U13920 (N_13920,N_5439,N_6082);
nand U13921 (N_13921,N_6367,N_6391);
or U13922 (N_13922,N_8587,N_6427);
nor U13923 (N_13923,N_9276,N_6465);
and U13924 (N_13924,N_5377,N_8861);
nand U13925 (N_13925,N_9749,N_9285);
and U13926 (N_13926,N_9859,N_7647);
nor U13927 (N_13927,N_9994,N_6610);
nor U13928 (N_13928,N_8437,N_9535);
xnor U13929 (N_13929,N_8724,N_6905);
nand U13930 (N_13930,N_8682,N_5945);
nand U13931 (N_13931,N_9342,N_5605);
and U13932 (N_13932,N_5736,N_9643);
or U13933 (N_13933,N_8593,N_5838);
nor U13934 (N_13934,N_9026,N_6669);
and U13935 (N_13935,N_8387,N_8355);
nand U13936 (N_13936,N_7797,N_9213);
and U13937 (N_13937,N_6962,N_7371);
nand U13938 (N_13938,N_9683,N_6232);
nor U13939 (N_13939,N_7429,N_8998);
nor U13940 (N_13940,N_6248,N_6934);
or U13941 (N_13941,N_5764,N_5442);
and U13942 (N_13942,N_8459,N_5386);
nand U13943 (N_13943,N_5885,N_7383);
nor U13944 (N_13944,N_8946,N_6066);
nor U13945 (N_13945,N_5710,N_9884);
nor U13946 (N_13946,N_5005,N_5511);
nor U13947 (N_13947,N_8871,N_5546);
and U13948 (N_13948,N_6924,N_9640);
nand U13949 (N_13949,N_6492,N_5251);
nand U13950 (N_13950,N_9708,N_8040);
or U13951 (N_13951,N_6536,N_6287);
xor U13952 (N_13952,N_7193,N_5303);
nand U13953 (N_13953,N_7724,N_8168);
or U13954 (N_13954,N_9382,N_6680);
and U13955 (N_13955,N_8925,N_7990);
nor U13956 (N_13956,N_6019,N_9882);
or U13957 (N_13957,N_5103,N_7942);
and U13958 (N_13958,N_9022,N_6017);
nand U13959 (N_13959,N_6954,N_7765);
nand U13960 (N_13960,N_6539,N_7053);
and U13961 (N_13961,N_5794,N_8754);
nor U13962 (N_13962,N_9719,N_9312);
nand U13963 (N_13963,N_7423,N_6831);
nor U13964 (N_13964,N_6024,N_7241);
nor U13965 (N_13965,N_9710,N_9611);
nand U13966 (N_13966,N_9647,N_9201);
and U13967 (N_13967,N_7910,N_8998);
or U13968 (N_13968,N_5657,N_7020);
nor U13969 (N_13969,N_7821,N_9554);
and U13970 (N_13970,N_9781,N_7655);
xor U13971 (N_13971,N_9482,N_6915);
and U13972 (N_13972,N_5298,N_9411);
and U13973 (N_13973,N_7437,N_7714);
nand U13974 (N_13974,N_9060,N_9999);
nand U13975 (N_13975,N_5702,N_9649);
nor U13976 (N_13976,N_7279,N_5792);
or U13977 (N_13977,N_7243,N_7208);
nand U13978 (N_13978,N_5946,N_5969);
and U13979 (N_13979,N_7845,N_6683);
and U13980 (N_13980,N_7031,N_7883);
and U13981 (N_13981,N_7598,N_7811);
nor U13982 (N_13982,N_7462,N_6391);
and U13983 (N_13983,N_8434,N_5105);
and U13984 (N_13984,N_6845,N_5066);
nor U13985 (N_13985,N_5938,N_9681);
nand U13986 (N_13986,N_8322,N_9019);
nor U13987 (N_13987,N_7060,N_8256);
or U13988 (N_13988,N_8466,N_8284);
nor U13989 (N_13989,N_7846,N_9015);
nor U13990 (N_13990,N_7505,N_8953);
and U13991 (N_13991,N_9829,N_8482);
nor U13992 (N_13992,N_8384,N_6798);
and U13993 (N_13993,N_5283,N_5258);
and U13994 (N_13994,N_9961,N_5517);
and U13995 (N_13995,N_8465,N_6012);
nand U13996 (N_13996,N_8177,N_7948);
nand U13997 (N_13997,N_5588,N_8271);
and U13998 (N_13998,N_9524,N_6040);
nand U13999 (N_13999,N_9082,N_7209);
and U14000 (N_14000,N_5787,N_6499);
nand U14001 (N_14001,N_7988,N_9466);
and U14002 (N_14002,N_5592,N_9549);
nor U14003 (N_14003,N_5935,N_7721);
nor U14004 (N_14004,N_9251,N_6416);
nor U14005 (N_14005,N_6467,N_8142);
nand U14006 (N_14006,N_7955,N_8983);
nor U14007 (N_14007,N_8691,N_7809);
or U14008 (N_14008,N_6173,N_7322);
nand U14009 (N_14009,N_8801,N_8311);
and U14010 (N_14010,N_7750,N_8477);
and U14011 (N_14011,N_8635,N_5460);
nand U14012 (N_14012,N_5342,N_5693);
xor U14013 (N_14013,N_7804,N_9836);
or U14014 (N_14014,N_5386,N_8763);
nor U14015 (N_14015,N_9284,N_8165);
nor U14016 (N_14016,N_9545,N_5475);
nand U14017 (N_14017,N_7167,N_8849);
nand U14018 (N_14018,N_6258,N_5608);
or U14019 (N_14019,N_5376,N_9193);
nand U14020 (N_14020,N_8416,N_7482);
and U14021 (N_14021,N_6406,N_7481);
nand U14022 (N_14022,N_8522,N_6514);
or U14023 (N_14023,N_7537,N_8323);
and U14024 (N_14024,N_6947,N_8706);
or U14025 (N_14025,N_8084,N_7995);
or U14026 (N_14026,N_9562,N_7288);
nand U14027 (N_14027,N_8120,N_9702);
nand U14028 (N_14028,N_6090,N_9330);
and U14029 (N_14029,N_8658,N_8191);
or U14030 (N_14030,N_8191,N_9996);
and U14031 (N_14031,N_8017,N_9854);
nor U14032 (N_14032,N_5014,N_7160);
nand U14033 (N_14033,N_9801,N_5469);
or U14034 (N_14034,N_5887,N_7358);
or U14035 (N_14035,N_8226,N_5658);
nor U14036 (N_14036,N_9790,N_8146);
and U14037 (N_14037,N_7634,N_6017);
nor U14038 (N_14038,N_9999,N_7338);
nor U14039 (N_14039,N_6518,N_8180);
nor U14040 (N_14040,N_7757,N_8985);
nor U14041 (N_14041,N_5951,N_7679);
nor U14042 (N_14042,N_9678,N_8557);
nand U14043 (N_14043,N_6229,N_5472);
nor U14044 (N_14044,N_6064,N_6683);
or U14045 (N_14045,N_5971,N_8088);
nor U14046 (N_14046,N_8550,N_8974);
nand U14047 (N_14047,N_9727,N_8194);
nand U14048 (N_14048,N_7998,N_6320);
or U14049 (N_14049,N_9235,N_7719);
nor U14050 (N_14050,N_8624,N_5607);
nand U14051 (N_14051,N_7150,N_9155);
nand U14052 (N_14052,N_7282,N_7428);
nor U14053 (N_14053,N_7458,N_7942);
or U14054 (N_14054,N_7424,N_8624);
nand U14055 (N_14055,N_5478,N_9844);
nand U14056 (N_14056,N_6616,N_5348);
nor U14057 (N_14057,N_8618,N_7146);
and U14058 (N_14058,N_9089,N_6434);
nand U14059 (N_14059,N_6751,N_9472);
or U14060 (N_14060,N_7795,N_7508);
or U14061 (N_14061,N_9104,N_7909);
and U14062 (N_14062,N_9080,N_7460);
nor U14063 (N_14063,N_9672,N_7645);
or U14064 (N_14064,N_9094,N_7441);
or U14065 (N_14065,N_8441,N_8278);
nand U14066 (N_14066,N_9673,N_5141);
or U14067 (N_14067,N_6711,N_5925);
nor U14068 (N_14068,N_8112,N_8141);
nor U14069 (N_14069,N_6386,N_9683);
and U14070 (N_14070,N_8046,N_5406);
nand U14071 (N_14071,N_7321,N_5944);
nand U14072 (N_14072,N_5810,N_5739);
or U14073 (N_14073,N_7479,N_7889);
nand U14074 (N_14074,N_8954,N_8160);
and U14075 (N_14075,N_9441,N_9148);
nor U14076 (N_14076,N_7800,N_7971);
nor U14077 (N_14077,N_9182,N_8658);
and U14078 (N_14078,N_5624,N_5628);
and U14079 (N_14079,N_7570,N_5962);
nand U14080 (N_14080,N_5511,N_7264);
or U14081 (N_14081,N_8265,N_7725);
and U14082 (N_14082,N_7165,N_9127);
nor U14083 (N_14083,N_7043,N_6529);
or U14084 (N_14084,N_8935,N_5755);
nor U14085 (N_14085,N_7139,N_8641);
or U14086 (N_14086,N_5849,N_7014);
nor U14087 (N_14087,N_5828,N_8258);
nand U14088 (N_14088,N_9716,N_6927);
nor U14089 (N_14089,N_5301,N_7630);
or U14090 (N_14090,N_6455,N_5601);
nor U14091 (N_14091,N_8202,N_5382);
and U14092 (N_14092,N_7596,N_9088);
nand U14093 (N_14093,N_7045,N_5573);
and U14094 (N_14094,N_6427,N_7806);
nand U14095 (N_14095,N_8611,N_9761);
and U14096 (N_14096,N_6667,N_8342);
or U14097 (N_14097,N_8083,N_9455);
or U14098 (N_14098,N_6393,N_8979);
nand U14099 (N_14099,N_7793,N_6694);
nor U14100 (N_14100,N_5337,N_8946);
or U14101 (N_14101,N_8690,N_5446);
nor U14102 (N_14102,N_6066,N_8126);
nand U14103 (N_14103,N_6604,N_6878);
or U14104 (N_14104,N_8793,N_9654);
nor U14105 (N_14105,N_6681,N_9541);
and U14106 (N_14106,N_7743,N_7792);
nand U14107 (N_14107,N_9207,N_9530);
and U14108 (N_14108,N_7207,N_6141);
nor U14109 (N_14109,N_7804,N_7535);
nor U14110 (N_14110,N_7153,N_9950);
or U14111 (N_14111,N_7652,N_7234);
or U14112 (N_14112,N_5479,N_8098);
nand U14113 (N_14113,N_8138,N_5754);
or U14114 (N_14114,N_8499,N_6392);
and U14115 (N_14115,N_6588,N_9925);
nor U14116 (N_14116,N_5884,N_9479);
and U14117 (N_14117,N_6360,N_6735);
or U14118 (N_14118,N_5084,N_6467);
nand U14119 (N_14119,N_9352,N_9647);
and U14120 (N_14120,N_8174,N_5353);
and U14121 (N_14121,N_5683,N_8210);
or U14122 (N_14122,N_5891,N_6874);
or U14123 (N_14123,N_9291,N_8866);
nor U14124 (N_14124,N_7828,N_7501);
nand U14125 (N_14125,N_8658,N_5354);
nor U14126 (N_14126,N_8553,N_9547);
and U14127 (N_14127,N_8045,N_8347);
or U14128 (N_14128,N_5152,N_9916);
or U14129 (N_14129,N_8792,N_8102);
and U14130 (N_14130,N_6253,N_9051);
xor U14131 (N_14131,N_6581,N_8270);
nand U14132 (N_14132,N_5389,N_7349);
nand U14133 (N_14133,N_8789,N_7486);
nor U14134 (N_14134,N_5832,N_6517);
or U14135 (N_14135,N_8400,N_5295);
and U14136 (N_14136,N_6264,N_5067);
and U14137 (N_14137,N_7940,N_7396);
nor U14138 (N_14138,N_6053,N_8871);
nand U14139 (N_14139,N_9250,N_9013);
and U14140 (N_14140,N_9480,N_5410);
nand U14141 (N_14141,N_5611,N_5566);
or U14142 (N_14142,N_6825,N_6876);
nor U14143 (N_14143,N_5766,N_7830);
xor U14144 (N_14144,N_7130,N_9163);
or U14145 (N_14145,N_6251,N_6992);
nand U14146 (N_14146,N_9475,N_8788);
nand U14147 (N_14147,N_9733,N_5939);
nand U14148 (N_14148,N_8245,N_9066);
nand U14149 (N_14149,N_5026,N_6063);
and U14150 (N_14150,N_8762,N_7679);
xor U14151 (N_14151,N_5580,N_6109);
nor U14152 (N_14152,N_9208,N_5432);
nand U14153 (N_14153,N_9734,N_7980);
nor U14154 (N_14154,N_9717,N_9634);
and U14155 (N_14155,N_9534,N_5071);
or U14156 (N_14156,N_5074,N_9258);
or U14157 (N_14157,N_9513,N_8937);
nand U14158 (N_14158,N_7314,N_8891);
or U14159 (N_14159,N_7033,N_6363);
or U14160 (N_14160,N_7419,N_8058);
nor U14161 (N_14161,N_6472,N_5485);
or U14162 (N_14162,N_5463,N_6806);
and U14163 (N_14163,N_9460,N_7383);
nor U14164 (N_14164,N_9224,N_8869);
and U14165 (N_14165,N_8577,N_7658);
or U14166 (N_14166,N_6757,N_8813);
or U14167 (N_14167,N_7381,N_7047);
nor U14168 (N_14168,N_6715,N_5403);
nand U14169 (N_14169,N_5278,N_8307);
nand U14170 (N_14170,N_6230,N_6359);
nand U14171 (N_14171,N_5219,N_6448);
nor U14172 (N_14172,N_8166,N_5964);
nor U14173 (N_14173,N_7383,N_7916);
nand U14174 (N_14174,N_5273,N_6720);
and U14175 (N_14175,N_9168,N_5993);
and U14176 (N_14176,N_8798,N_8204);
nor U14177 (N_14177,N_8572,N_6377);
and U14178 (N_14178,N_5570,N_9046);
and U14179 (N_14179,N_6752,N_5113);
nor U14180 (N_14180,N_6009,N_6814);
nand U14181 (N_14181,N_5839,N_5077);
nand U14182 (N_14182,N_9113,N_8578);
or U14183 (N_14183,N_5882,N_6760);
nor U14184 (N_14184,N_5950,N_7339);
nand U14185 (N_14185,N_6296,N_6971);
nor U14186 (N_14186,N_5447,N_7302);
nand U14187 (N_14187,N_7826,N_9543);
and U14188 (N_14188,N_9731,N_7361);
or U14189 (N_14189,N_9389,N_9450);
or U14190 (N_14190,N_5360,N_9701);
and U14191 (N_14191,N_7570,N_8944);
or U14192 (N_14192,N_8969,N_6829);
or U14193 (N_14193,N_5515,N_7170);
and U14194 (N_14194,N_5437,N_7313);
or U14195 (N_14195,N_5782,N_6002);
nand U14196 (N_14196,N_6432,N_9738);
and U14197 (N_14197,N_5602,N_6503);
nor U14198 (N_14198,N_5909,N_6957);
or U14199 (N_14199,N_6242,N_6926);
or U14200 (N_14200,N_9386,N_6076);
or U14201 (N_14201,N_6453,N_9255);
nor U14202 (N_14202,N_6870,N_9561);
xnor U14203 (N_14203,N_8786,N_5006);
or U14204 (N_14204,N_6807,N_9943);
or U14205 (N_14205,N_6729,N_5227);
nand U14206 (N_14206,N_6594,N_9643);
nor U14207 (N_14207,N_5203,N_8253);
nand U14208 (N_14208,N_5509,N_7127);
or U14209 (N_14209,N_9570,N_5730);
or U14210 (N_14210,N_7164,N_7621);
and U14211 (N_14211,N_5209,N_6702);
and U14212 (N_14212,N_9932,N_9158);
nor U14213 (N_14213,N_8043,N_7862);
nor U14214 (N_14214,N_6583,N_7145);
and U14215 (N_14215,N_8441,N_9429);
nand U14216 (N_14216,N_6041,N_9009);
and U14217 (N_14217,N_5635,N_5035);
nand U14218 (N_14218,N_5215,N_8365);
nand U14219 (N_14219,N_9709,N_9490);
and U14220 (N_14220,N_5154,N_6706);
xor U14221 (N_14221,N_8622,N_6998);
nand U14222 (N_14222,N_8245,N_6614);
nor U14223 (N_14223,N_8059,N_6243);
nor U14224 (N_14224,N_6118,N_5854);
or U14225 (N_14225,N_7646,N_9655);
nor U14226 (N_14226,N_9625,N_9767);
nor U14227 (N_14227,N_6037,N_5959);
and U14228 (N_14228,N_9929,N_5309);
or U14229 (N_14229,N_7592,N_6992);
and U14230 (N_14230,N_7402,N_9153);
nand U14231 (N_14231,N_8105,N_6796);
nand U14232 (N_14232,N_9349,N_6831);
and U14233 (N_14233,N_7482,N_8918);
nor U14234 (N_14234,N_9028,N_5661);
and U14235 (N_14235,N_7632,N_9642);
nand U14236 (N_14236,N_5654,N_7088);
nor U14237 (N_14237,N_6431,N_7915);
or U14238 (N_14238,N_9793,N_8192);
and U14239 (N_14239,N_7285,N_9205);
or U14240 (N_14240,N_7718,N_8107);
nor U14241 (N_14241,N_8089,N_9534);
or U14242 (N_14242,N_7920,N_9770);
and U14243 (N_14243,N_6019,N_9565);
and U14244 (N_14244,N_5240,N_9297);
nand U14245 (N_14245,N_5200,N_7500);
and U14246 (N_14246,N_9529,N_6176);
or U14247 (N_14247,N_7142,N_5831);
and U14248 (N_14248,N_8155,N_5220);
or U14249 (N_14249,N_8898,N_8591);
and U14250 (N_14250,N_8131,N_7963);
or U14251 (N_14251,N_5219,N_6800);
and U14252 (N_14252,N_5067,N_9396);
nand U14253 (N_14253,N_5905,N_9472);
nand U14254 (N_14254,N_9242,N_5754);
nand U14255 (N_14255,N_7548,N_9147);
or U14256 (N_14256,N_6054,N_6474);
and U14257 (N_14257,N_9978,N_9574);
or U14258 (N_14258,N_5248,N_5027);
nor U14259 (N_14259,N_5281,N_5415);
nor U14260 (N_14260,N_6416,N_9864);
or U14261 (N_14261,N_8119,N_7701);
and U14262 (N_14262,N_9730,N_5772);
nor U14263 (N_14263,N_9534,N_7484);
and U14264 (N_14264,N_7350,N_5717);
nor U14265 (N_14265,N_6584,N_6637);
nor U14266 (N_14266,N_6424,N_5513);
nor U14267 (N_14267,N_8278,N_5497);
xor U14268 (N_14268,N_5968,N_8512);
or U14269 (N_14269,N_6421,N_6427);
nand U14270 (N_14270,N_8249,N_6719);
and U14271 (N_14271,N_6826,N_6786);
nand U14272 (N_14272,N_7689,N_8244);
nand U14273 (N_14273,N_5432,N_6334);
or U14274 (N_14274,N_8252,N_7639);
nand U14275 (N_14275,N_5653,N_5351);
or U14276 (N_14276,N_7721,N_5547);
and U14277 (N_14277,N_5458,N_7304);
xor U14278 (N_14278,N_9885,N_9241);
and U14279 (N_14279,N_9263,N_5598);
or U14280 (N_14280,N_7011,N_9353);
and U14281 (N_14281,N_9450,N_5720);
and U14282 (N_14282,N_5449,N_6327);
or U14283 (N_14283,N_6776,N_9843);
and U14284 (N_14284,N_5378,N_7334);
and U14285 (N_14285,N_8659,N_6587);
nand U14286 (N_14286,N_8552,N_5051);
nand U14287 (N_14287,N_6984,N_5794);
nor U14288 (N_14288,N_9102,N_7985);
and U14289 (N_14289,N_9680,N_9422);
and U14290 (N_14290,N_8511,N_8768);
and U14291 (N_14291,N_7997,N_5172);
and U14292 (N_14292,N_5815,N_7839);
nor U14293 (N_14293,N_6442,N_7902);
and U14294 (N_14294,N_7324,N_7820);
xor U14295 (N_14295,N_9083,N_7812);
nor U14296 (N_14296,N_7079,N_6521);
nand U14297 (N_14297,N_5958,N_6461);
and U14298 (N_14298,N_9944,N_8758);
and U14299 (N_14299,N_9959,N_8770);
or U14300 (N_14300,N_7846,N_5832);
and U14301 (N_14301,N_5840,N_7351);
or U14302 (N_14302,N_9524,N_5495);
or U14303 (N_14303,N_6123,N_5855);
or U14304 (N_14304,N_8859,N_8074);
or U14305 (N_14305,N_9495,N_5635);
nor U14306 (N_14306,N_9173,N_5076);
nand U14307 (N_14307,N_6473,N_6485);
or U14308 (N_14308,N_7928,N_9122);
nor U14309 (N_14309,N_6718,N_9163);
nor U14310 (N_14310,N_5042,N_5992);
or U14311 (N_14311,N_7246,N_9161);
or U14312 (N_14312,N_6463,N_6107);
and U14313 (N_14313,N_7668,N_5486);
and U14314 (N_14314,N_9615,N_8549);
nand U14315 (N_14315,N_5174,N_5996);
nand U14316 (N_14316,N_7103,N_7675);
and U14317 (N_14317,N_8125,N_8660);
or U14318 (N_14318,N_6308,N_8986);
nand U14319 (N_14319,N_9881,N_9233);
nor U14320 (N_14320,N_6074,N_5545);
or U14321 (N_14321,N_7613,N_8553);
and U14322 (N_14322,N_5488,N_9194);
nand U14323 (N_14323,N_9810,N_8576);
nand U14324 (N_14324,N_7493,N_9726);
nor U14325 (N_14325,N_8333,N_6713);
and U14326 (N_14326,N_6522,N_8964);
nand U14327 (N_14327,N_7045,N_7473);
nand U14328 (N_14328,N_7009,N_5581);
nand U14329 (N_14329,N_7946,N_8788);
nand U14330 (N_14330,N_8541,N_8149);
nor U14331 (N_14331,N_6729,N_8421);
nand U14332 (N_14332,N_8277,N_7350);
nor U14333 (N_14333,N_8238,N_6731);
or U14334 (N_14334,N_5226,N_5238);
or U14335 (N_14335,N_5246,N_8179);
or U14336 (N_14336,N_7586,N_9735);
nand U14337 (N_14337,N_9302,N_6192);
or U14338 (N_14338,N_9375,N_8289);
nand U14339 (N_14339,N_7891,N_8740);
nor U14340 (N_14340,N_8209,N_9322);
nor U14341 (N_14341,N_8640,N_5520);
and U14342 (N_14342,N_6078,N_5462);
nor U14343 (N_14343,N_5301,N_9556);
and U14344 (N_14344,N_7137,N_9291);
nor U14345 (N_14345,N_6730,N_5427);
and U14346 (N_14346,N_9147,N_6012);
nor U14347 (N_14347,N_5524,N_5259);
and U14348 (N_14348,N_5343,N_6939);
or U14349 (N_14349,N_9022,N_9721);
nand U14350 (N_14350,N_6287,N_5352);
or U14351 (N_14351,N_5872,N_8923);
or U14352 (N_14352,N_5492,N_8405);
or U14353 (N_14353,N_7130,N_9691);
nor U14354 (N_14354,N_8039,N_6841);
nor U14355 (N_14355,N_8121,N_9938);
and U14356 (N_14356,N_7180,N_6764);
and U14357 (N_14357,N_5570,N_9492);
nor U14358 (N_14358,N_9586,N_6299);
and U14359 (N_14359,N_6288,N_7171);
and U14360 (N_14360,N_9119,N_5855);
or U14361 (N_14361,N_8948,N_5912);
nand U14362 (N_14362,N_8919,N_8577);
or U14363 (N_14363,N_9599,N_9701);
nor U14364 (N_14364,N_9425,N_7558);
and U14365 (N_14365,N_9722,N_9658);
nand U14366 (N_14366,N_8664,N_9975);
and U14367 (N_14367,N_7921,N_8615);
nand U14368 (N_14368,N_7163,N_7787);
or U14369 (N_14369,N_8309,N_7957);
nand U14370 (N_14370,N_8996,N_9809);
or U14371 (N_14371,N_5123,N_6504);
nand U14372 (N_14372,N_9937,N_5383);
nand U14373 (N_14373,N_9742,N_5064);
or U14374 (N_14374,N_9005,N_5907);
nor U14375 (N_14375,N_5706,N_5749);
or U14376 (N_14376,N_9933,N_5068);
xnor U14377 (N_14377,N_7137,N_9123);
nor U14378 (N_14378,N_5008,N_8659);
nor U14379 (N_14379,N_8784,N_8792);
nor U14380 (N_14380,N_6146,N_8491);
nand U14381 (N_14381,N_6993,N_5209);
nand U14382 (N_14382,N_9697,N_5674);
or U14383 (N_14383,N_9720,N_8723);
nand U14384 (N_14384,N_6979,N_7235);
and U14385 (N_14385,N_9494,N_8899);
and U14386 (N_14386,N_9935,N_5628);
and U14387 (N_14387,N_8687,N_7323);
and U14388 (N_14388,N_7503,N_7721);
nand U14389 (N_14389,N_5066,N_8702);
and U14390 (N_14390,N_6377,N_5213);
or U14391 (N_14391,N_5079,N_8821);
nand U14392 (N_14392,N_7648,N_6134);
and U14393 (N_14393,N_5583,N_5076);
nand U14394 (N_14394,N_9546,N_7588);
nand U14395 (N_14395,N_9311,N_7482);
nand U14396 (N_14396,N_6995,N_7358);
or U14397 (N_14397,N_5825,N_5692);
or U14398 (N_14398,N_9797,N_9366);
nand U14399 (N_14399,N_6956,N_9055);
nor U14400 (N_14400,N_8758,N_8944);
or U14401 (N_14401,N_9141,N_5103);
nor U14402 (N_14402,N_7830,N_7478);
nand U14403 (N_14403,N_6558,N_9771);
and U14404 (N_14404,N_5927,N_8629);
nor U14405 (N_14405,N_9175,N_8329);
nand U14406 (N_14406,N_5035,N_5636);
or U14407 (N_14407,N_9785,N_5387);
nor U14408 (N_14408,N_5492,N_8193);
nand U14409 (N_14409,N_6014,N_7689);
nand U14410 (N_14410,N_8682,N_5750);
nor U14411 (N_14411,N_5587,N_6246);
and U14412 (N_14412,N_8774,N_9153);
nor U14413 (N_14413,N_9886,N_5953);
nand U14414 (N_14414,N_8063,N_7927);
and U14415 (N_14415,N_5006,N_9496);
and U14416 (N_14416,N_5487,N_9752);
nor U14417 (N_14417,N_7441,N_6334);
and U14418 (N_14418,N_8171,N_6384);
and U14419 (N_14419,N_6289,N_8339);
and U14420 (N_14420,N_9043,N_6196);
nor U14421 (N_14421,N_5420,N_7914);
nand U14422 (N_14422,N_6067,N_9500);
nand U14423 (N_14423,N_5864,N_5981);
nor U14424 (N_14424,N_5467,N_7875);
nor U14425 (N_14425,N_6762,N_6943);
or U14426 (N_14426,N_6288,N_8063);
or U14427 (N_14427,N_7534,N_6874);
nand U14428 (N_14428,N_7604,N_8100);
and U14429 (N_14429,N_5891,N_7071);
nor U14430 (N_14430,N_6243,N_8345);
nand U14431 (N_14431,N_7012,N_7963);
nand U14432 (N_14432,N_8313,N_8074);
nand U14433 (N_14433,N_8694,N_8443);
or U14434 (N_14434,N_6851,N_9982);
and U14435 (N_14435,N_6330,N_9421);
or U14436 (N_14436,N_6335,N_6576);
and U14437 (N_14437,N_8288,N_9311);
and U14438 (N_14438,N_5252,N_8394);
and U14439 (N_14439,N_7758,N_7115);
or U14440 (N_14440,N_5318,N_8375);
nor U14441 (N_14441,N_8030,N_7527);
nor U14442 (N_14442,N_6946,N_8066);
nor U14443 (N_14443,N_5322,N_8762);
nand U14444 (N_14444,N_5352,N_6378);
nor U14445 (N_14445,N_7131,N_7613);
or U14446 (N_14446,N_9763,N_9244);
or U14447 (N_14447,N_7088,N_8521);
or U14448 (N_14448,N_7845,N_7105);
nand U14449 (N_14449,N_5526,N_7050);
or U14450 (N_14450,N_7693,N_7918);
or U14451 (N_14451,N_9508,N_6365);
nand U14452 (N_14452,N_9398,N_9509);
nor U14453 (N_14453,N_6099,N_8572);
and U14454 (N_14454,N_8527,N_7216);
nor U14455 (N_14455,N_5961,N_5468);
and U14456 (N_14456,N_6406,N_6216);
nor U14457 (N_14457,N_6387,N_9077);
nor U14458 (N_14458,N_8787,N_9942);
or U14459 (N_14459,N_5739,N_6146);
nand U14460 (N_14460,N_6227,N_8610);
or U14461 (N_14461,N_9593,N_8021);
nand U14462 (N_14462,N_8890,N_6117);
nand U14463 (N_14463,N_5365,N_5850);
nor U14464 (N_14464,N_8117,N_8162);
and U14465 (N_14465,N_8726,N_6298);
nor U14466 (N_14466,N_9068,N_8040);
or U14467 (N_14467,N_5843,N_6545);
or U14468 (N_14468,N_8769,N_5591);
nor U14469 (N_14469,N_6885,N_6888);
nand U14470 (N_14470,N_7639,N_5390);
and U14471 (N_14471,N_5785,N_6252);
and U14472 (N_14472,N_9047,N_7805);
xor U14473 (N_14473,N_7274,N_6329);
or U14474 (N_14474,N_7644,N_8606);
nand U14475 (N_14475,N_6115,N_7254);
nand U14476 (N_14476,N_9761,N_8487);
xor U14477 (N_14477,N_8632,N_7217);
or U14478 (N_14478,N_7799,N_8394);
and U14479 (N_14479,N_7709,N_6959);
nand U14480 (N_14480,N_8342,N_7694);
nand U14481 (N_14481,N_6265,N_7771);
or U14482 (N_14482,N_8319,N_5710);
nor U14483 (N_14483,N_7307,N_8992);
or U14484 (N_14484,N_9974,N_7300);
or U14485 (N_14485,N_6059,N_6194);
or U14486 (N_14486,N_6046,N_5667);
nor U14487 (N_14487,N_6799,N_5673);
nor U14488 (N_14488,N_8404,N_9170);
nand U14489 (N_14489,N_7385,N_7649);
or U14490 (N_14490,N_9884,N_9427);
nor U14491 (N_14491,N_6291,N_7100);
and U14492 (N_14492,N_8736,N_7325);
or U14493 (N_14493,N_6255,N_6431);
or U14494 (N_14494,N_9747,N_9442);
nand U14495 (N_14495,N_8413,N_7122);
or U14496 (N_14496,N_8844,N_6126);
nor U14497 (N_14497,N_8584,N_7586);
and U14498 (N_14498,N_6568,N_6981);
nand U14499 (N_14499,N_5491,N_7558);
and U14500 (N_14500,N_9137,N_5491);
nand U14501 (N_14501,N_8397,N_7842);
and U14502 (N_14502,N_9516,N_7442);
or U14503 (N_14503,N_7656,N_5473);
and U14504 (N_14504,N_9694,N_8342);
nand U14505 (N_14505,N_5598,N_5029);
nor U14506 (N_14506,N_7267,N_9857);
or U14507 (N_14507,N_5389,N_5272);
or U14508 (N_14508,N_6417,N_6128);
nor U14509 (N_14509,N_5816,N_5594);
and U14510 (N_14510,N_6463,N_7347);
nor U14511 (N_14511,N_9547,N_9155);
and U14512 (N_14512,N_7472,N_8149);
and U14513 (N_14513,N_6038,N_6163);
and U14514 (N_14514,N_6574,N_7374);
nor U14515 (N_14515,N_6223,N_6066);
and U14516 (N_14516,N_9913,N_5828);
nor U14517 (N_14517,N_5862,N_8991);
nor U14518 (N_14518,N_7616,N_9276);
nand U14519 (N_14519,N_7587,N_7789);
or U14520 (N_14520,N_6011,N_6749);
nand U14521 (N_14521,N_7870,N_7081);
nor U14522 (N_14522,N_5463,N_8954);
nand U14523 (N_14523,N_9098,N_5296);
nor U14524 (N_14524,N_5927,N_6862);
and U14525 (N_14525,N_8865,N_5454);
nand U14526 (N_14526,N_7984,N_6261);
and U14527 (N_14527,N_6896,N_6096);
nor U14528 (N_14528,N_7801,N_7053);
and U14529 (N_14529,N_8416,N_6160);
and U14530 (N_14530,N_7172,N_8567);
xnor U14531 (N_14531,N_5155,N_6697);
or U14532 (N_14532,N_5234,N_9427);
and U14533 (N_14533,N_7411,N_6126);
nand U14534 (N_14534,N_6146,N_6347);
and U14535 (N_14535,N_9795,N_9807);
or U14536 (N_14536,N_8715,N_5022);
and U14537 (N_14537,N_8394,N_8847);
or U14538 (N_14538,N_5907,N_9696);
and U14539 (N_14539,N_5659,N_5980);
and U14540 (N_14540,N_9467,N_7083);
nor U14541 (N_14541,N_7964,N_5646);
or U14542 (N_14542,N_6443,N_6088);
nor U14543 (N_14543,N_7898,N_8830);
nor U14544 (N_14544,N_6573,N_5947);
or U14545 (N_14545,N_5747,N_9900);
or U14546 (N_14546,N_7639,N_9639);
or U14547 (N_14547,N_5335,N_8853);
or U14548 (N_14548,N_5285,N_9841);
nand U14549 (N_14549,N_9200,N_6215);
nor U14550 (N_14550,N_5254,N_7641);
nor U14551 (N_14551,N_5450,N_9676);
or U14552 (N_14552,N_5708,N_5994);
nor U14553 (N_14553,N_5208,N_6792);
nand U14554 (N_14554,N_7793,N_7080);
or U14555 (N_14555,N_7970,N_9352);
or U14556 (N_14556,N_7100,N_5803);
nand U14557 (N_14557,N_9171,N_8411);
xor U14558 (N_14558,N_9475,N_7785);
or U14559 (N_14559,N_5150,N_7157);
and U14560 (N_14560,N_5981,N_5885);
nor U14561 (N_14561,N_6813,N_5675);
nor U14562 (N_14562,N_9786,N_5250);
nor U14563 (N_14563,N_5796,N_7387);
or U14564 (N_14564,N_6507,N_9006);
and U14565 (N_14565,N_9202,N_5126);
nor U14566 (N_14566,N_6331,N_6496);
nor U14567 (N_14567,N_8582,N_6447);
nand U14568 (N_14568,N_7001,N_7902);
or U14569 (N_14569,N_6322,N_6366);
nand U14570 (N_14570,N_5308,N_8031);
nand U14571 (N_14571,N_5217,N_5104);
nand U14572 (N_14572,N_7053,N_8797);
or U14573 (N_14573,N_6604,N_7737);
or U14574 (N_14574,N_6352,N_6162);
nor U14575 (N_14575,N_6658,N_5228);
nand U14576 (N_14576,N_9782,N_8691);
and U14577 (N_14577,N_8414,N_8355);
nor U14578 (N_14578,N_7888,N_8937);
nand U14579 (N_14579,N_7413,N_5836);
nor U14580 (N_14580,N_8952,N_8971);
nor U14581 (N_14581,N_8552,N_7531);
and U14582 (N_14582,N_6811,N_7669);
nor U14583 (N_14583,N_6286,N_7310);
or U14584 (N_14584,N_8827,N_7451);
and U14585 (N_14585,N_7585,N_6606);
or U14586 (N_14586,N_6881,N_6962);
and U14587 (N_14587,N_9605,N_9497);
nand U14588 (N_14588,N_6852,N_5021);
or U14589 (N_14589,N_5628,N_9889);
and U14590 (N_14590,N_8427,N_5388);
and U14591 (N_14591,N_6466,N_5090);
nand U14592 (N_14592,N_6421,N_5632);
nor U14593 (N_14593,N_7858,N_7515);
nor U14594 (N_14594,N_5019,N_6210);
and U14595 (N_14595,N_9185,N_9292);
nand U14596 (N_14596,N_6698,N_6867);
nand U14597 (N_14597,N_6012,N_5753);
or U14598 (N_14598,N_8936,N_7453);
nor U14599 (N_14599,N_7504,N_9845);
nand U14600 (N_14600,N_5878,N_9655);
nor U14601 (N_14601,N_9321,N_7797);
or U14602 (N_14602,N_6699,N_6633);
nor U14603 (N_14603,N_5251,N_9335);
nor U14604 (N_14604,N_6499,N_8289);
or U14605 (N_14605,N_8917,N_7701);
or U14606 (N_14606,N_5081,N_8762);
and U14607 (N_14607,N_9266,N_9767);
and U14608 (N_14608,N_5715,N_8085);
nor U14609 (N_14609,N_9621,N_9374);
and U14610 (N_14610,N_7146,N_7045);
nor U14611 (N_14611,N_5742,N_8301);
and U14612 (N_14612,N_9604,N_5068);
xor U14613 (N_14613,N_8435,N_5005);
or U14614 (N_14614,N_8641,N_5572);
or U14615 (N_14615,N_7797,N_6768);
and U14616 (N_14616,N_7979,N_7851);
nor U14617 (N_14617,N_7949,N_8633);
and U14618 (N_14618,N_5675,N_9878);
nor U14619 (N_14619,N_8806,N_9396);
nor U14620 (N_14620,N_8606,N_9907);
nor U14621 (N_14621,N_9017,N_6338);
or U14622 (N_14622,N_6221,N_5330);
or U14623 (N_14623,N_9283,N_9771);
and U14624 (N_14624,N_8616,N_5565);
nand U14625 (N_14625,N_5126,N_7848);
or U14626 (N_14626,N_5606,N_9671);
nor U14627 (N_14627,N_6189,N_5237);
and U14628 (N_14628,N_8845,N_7891);
nor U14629 (N_14629,N_5766,N_6686);
and U14630 (N_14630,N_9295,N_6323);
nand U14631 (N_14631,N_6575,N_9126);
or U14632 (N_14632,N_5437,N_8564);
or U14633 (N_14633,N_6682,N_8983);
nor U14634 (N_14634,N_8939,N_7479);
and U14635 (N_14635,N_6460,N_5884);
nand U14636 (N_14636,N_9566,N_7204);
nor U14637 (N_14637,N_9714,N_5982);
or U14638 (N_14638,N_7520,N_7449);
and U14639 (N_14639,N_9904,N_8198);
nand U14640 (N_14640,N_8233,N_6334);
and U14641 (N_14641,N_5621,N_8313);
and U14642 (N_14642,N_6799,N_8402);
nand U14643 (N_14643,N_5790,N_9799);
and U14644 (N_14644,N_6870,N_6840);
nor U14645 (N_14645,N_9679,N_7016);
or U14646 (N_14646,N_9048,N_9606);
nor U14647 (N_14647,N_6972,N_5246);
nand U14648 (N_14648,N_6527,N_9566);
and U14649 (N_14649,N_9521,N_9687);
nand U14650 (N_14650,N_5172,N_7339);
nor U14651 (N_14651,N_8674,N_5823);
nor U14652 (N_14652,N_9038,N_5894);
nor U14653 (N_14653,N_5424,N_6285);
or U14654 (N_14654,N_8158,N_9279);
nand U14655 (N_14655,N_9869,N_8051);
and U14656 (N_14656,N_7046,N_6771);
and U14657 (N_14657,N_9682,N_7543);
nor U14658 (N_14658,N_6165,N_7809);
or U14659 (N_14659,N_9098,N_8085);
nand U14660 (N_14660,N_8296,N_9270);
and U14661 (N_14661,N_9654,N_7497);
nand U14662 (N_14662,N_6180,N_9252);
nand U14663 (N_14663,N_9403,N_8992);
nand U14664 (N_14664,N_6977,N_8851);
or U14665 (N_14665,N_9584,N_6646);
nand U14666 (N_14666,N_7942,N_5828);
nand U14667 (N_14667,N_8956,N_7537);
nor U14668 (N_14668,N_9476,N_7162);
nor U14669 (N_14669,N_6667,N_6596);
nand U14670 (N_14670,N_5021,N_9617);
and U14671 (N_14671,N_8385,N_7298);
or U14672 (N_14672,N_7712,N_6164);
and U14673 (N_14673,N_7999,N_5896);
or U14674 (N_14674,N_9339,N_9876);
nand U14675 (N_14675,N_8527,N_9284);
nor U14676 (N_14676,N_6473,N_5356);
or U14677 (N_14677,N_5923,N_6343);
or U14678 (N_14678,N_8635,N_8519);
and U14679 (N_14679,N_5919,N_5862);
nor U14680 (N_14680,N_5487,N_5638);
or U14681 (N_14681,N_7537,N_7442);
and U14682 (N_14682,N_5340,N_7531);
nor U14683 (N_14683,N_6054,N_7997);
nor U14684 (N_14684,N_7254,N_5473);
or U14685 (N_14685,N_7090,N_6109);
nor U14686 (N_14686,N_6098,N_8064);
or U14687 (N_14687,N_9829,N_7665);
and U14688 (N_14688,N_5261,N_7343);
nor U14689 (N_14689,N_6261,N_8743);
or U14690 (N_14690,N_7974,N_5739);
nor U14691 (N_14691,N_8625,N_5440);
nor U14692 (N_14692,N_9297,N_8369);
or U14693 (N_14693,N_5139,N_9091);
and U14694 (N_14694,N_9435,N_9636);
or U14695 (N_14695,N_9045,N_8276);
nor U14696 (N_14696,N_6801,N_8356);
or U14697 (N_14697,N_7940,N_7017);
or U14698 (N_14698,N_6353,N_8507);
or U14699 (N_14699,N_8542,N_8690);
and U14700 (N_14700,N_8989,N_6831);
and U14701 (N_14701,N_5279,N_7222);
or U14702 (N_14702,N_7255,N_9977);
or U14703 (N_14703,N_6707,N_8126);
or U14704 (N_14704,N_5249,N_9667);
or U14705 (N_14705,N_9418,N_9670);
or U14706 (N_14706,N_9564,N_7685);
and U14707 (N_14707,N_8931,N_6619);
and U14708 (N_14708,N_5758,N_5872);
or U14709 (N_14709,N_7299,N_9238);
nor U14710 (N_14710,N_6647,N_6165);
nand U14711 (N_14711,N_8143,N_7788);
and U14712 (N_14712,N_7412,N_6736);
nand U14713 (N_14713,N_9872,N_9134);
nor U14714 (N_14714,N_8034,N_9329);
or U14715 (N_14715,N_8158,N_8258);
nor U14716 (N_14716,N_5635,N_6149);
nand U14717 (N_14717,N_8268,N_8625);
nor U14718 (N_14718,N_9717,N_7972);
and U14719 (N_14719,N_7761,N_5174);
nand U14720 (N_14720,N_8395,N_8216);
or U14721 (N_14721,N_8682,N_5844);
nor U14722 (N_14722,N_7875,N_9004);
and U14723 (N_14723,N_6203,N_6508);
nand U14724 (N_14724,N_7403,N_7099);
nor U14725 (N_14725,N_5522,N_8146);
nand U14726 (N_14726,N_5565,N_6329);
xor U14727 (N_14727,N_9091,N_7217);
nor U14728 (N_14728,N_7986,N_6853);
and U14729 (N_14729,N_6703,N_6983);
nand U14730 (N_14730,N_9878,N_9860);
or U14731 (N_14731,N_5149,N_8943);
nand U14732 (N_14732,N_6629,N_9923);
nor U14733 (N_14733,N_9604,N_9340);
nand U14734 (N_14734,N_8395,N_5246);
nand U14735 (N_14735,N_7108,N_8989);
and U14736 (N_14736,N_8297,N_8977);
nor U14737 (N_14737,N_9963,N_9179);
nand U14738 (N_14738,N_8607,N_7388);
or U14739 (N_14739,N_7165,N_9986);
or U14740 (N_14740,N_9517,N_6714);
xnor U14741 (N_14741,N_8636,N_6719);
nand U14742 (N_14742,N_8648,N_6114);
or U14743 (N_14743,N_9913,N_6102);
or U14744 (N_14744,N_9571,N_6721);
and U14745 (N_14745,N_6000,N_7243);
nor U14746 (N_14746,N_6023,N_8752);
and U14747 (N_14747,N_8669,N_8117);
and U14748 (N_14748,N_9011,N_7184);
or U14749 (N_14749,N_5729,N_9709);
or U14750 (N_14750,N_6877,N_5925);
nor U14751 (N_14751,N_9420,N_5274);
nand U14752 (N_14752,N_6537,N_6406);
and U14753 (N_14753,N_6365,N_9448);
and U14754 (N_14754,N_8830,N_9418);
nand U14755 (N_14755,N_7351,N_9378);
or U14756 (N_14756,N_8051,N_7056);
and U14757 (N_14757,N_9043,N_9361);
nor U14758 (N_14758,N_5590,N_5727);
nand U14759 (N_14759,N_8993,N_9993);
nand U14760 (N_14760,N_8800,N_9303);
and U14761 (N_14761,N_9410,N_9267);
nor U14762 (N_14762,N_5804,N_7259);
and U14763 (N_14763,N_9129,N_8574);
nor U14764 (N_14764,N_8691,N_6558);
nor U14765 (N_14765,N_9180,N_5122);
nor U14766 (N_14766,N_8293,N_7468);
or U14767 (N_14767,N_7402,N_5689);
nor U14768 (N_14768,N_9805,N_9371);
nor U14769 (N_14769,N_5405,N_5980);
or U14770 (N_14770,N_9293,N_6101);
nand U14771 (N_14771,N_8253,N_8339);
nor U14772 (N_14772,N_8977,N_8855);
nor U14773 (N_14773,N_8756,N_8296);
or U14774 (N_14774,N_7741,N_9517);
or U14775 (N_14775,N_5724,N_9722);
and U14776 (N_14776,N_7042,N_8722);
nor U14777 (N_14777,N_9243,N_6420);
nor U14778 (N_14778,N_7978,N_9420);
or U14779 (N_14779,N_6653,N_6140);
nor U14780 (N_14780,N_9616,N_6086);
or U14781 (N_14781,N_9816,N_5390);
nand U14782 (N_14782,N_8743,N_5937);
and U14783 (N_14783,N_8929,N_7110);
or U14784 (N_14784,N_8330,N_9454);
nor U14785 (N_14785,N_7837,N_8967);
nand U14786 (N_14786,N_9480,N_7709);
or U14787 (N_14787,N_6607,N_7438);
or U14788 (N_14788,N_7911,N_8551);
nand U14789 (N_14789,N_6305,N_9504);
or U14790 (N_14790,N_8243,N_8121);
and U14791 (N_14791,N_5732,N_6901);
and U14792 (N_14792,N_9425,N_7440);
nand U14793 (N_14793,N_8738,N_9909);
and U14794 (N_14794,N_7804,N_7824);
nand U14795 (N_14795,N_8522,N_7296);
nand U14796 (N_14796,N_9187,N_7386);
nor U14797 (N_14797,N_8025,N_5634);
and U14798 (N_14798,N_5778,N_7727);
nor U14799 (N_14799,N_9692,N_6174);
and U14800 (N_14800,N_6967,N_6698);
and U14801 (N_14801,N_7362,N_5865);
or U14802 (N_14802,N_8885,N_6286);
nand U14803 (N_14803,N_5498,N_8921);
and U14804 (N_14804,N_7619,N_8175);
nor U14805 (N_14805,N_5224,N_8772);
nand U14806 (N_14806,N_5742,N_9331);
nor U14807 (N_14807,N_9799,N_5572);
and U14808 (N_14808,N_6939,N_8413);
nor U14809 (N_14809,N_6519,N_5853);
or U14810 (N_14810,N_7086,N_7035);
nand U14811 (N_14811,N_8557,N_7829);
and U14812 (N_14812,N_6361,N_7004);
nand U14813 (N_14813,N_9288,N_5645);
nor U14814 (N_14814,N_9005,N_7955);
nor U14815 (N_14815,N_5229,N_9444);
nand U14816 (N_14816,N_8906,N_7850);
nor U14817 (N_14817,N_8387,N_8821);
or U14818 (N_14818,N_6556,N_8401);
or U14819 (N_14819,N_8613,N_8063);
and U14820 (N_14820,N_5637,N_6941);
nand U14821 (N_14821,N_8678,N_6113);
nor U14822 (N_14822,N_8067,N_8510);
nand U14823 (N_14823,N_8860,N_8250);
and U14824 (N_14824,N_7400,N_6697);
and U14825 (N_14825,N_6419,N_6366);
nand U14826 (N_14826,N_6001,N_5291);
nand U14827 (N_14827,N_6355,N_9153);
or U14828 (N_14828,N_6803,N_6267);
and U14829 (N_14829,N_6135,N_7670);
or U14830 (N_14830,N_9700,N_7030);
nand U14831 (N_14831,N_5680,N_6426);
and U14832 (N_14832,N_5074,N_6316);
and U14833 (N_14833,N_6949,N_6341);
nor U14834 (N_14834,N_9101,N_8432);
or U14835 (N_14835,N_8036,N_9060);
or U14836 (N_14836,N_7530,N_6036);
nand U14837 (N_14837,N_9012,N_6577);
or U14838 (N_14838,N_5118,N_5562);
and U14839 (N_14839,N_8942,N_5248);
nand U14840 (N_14840,N_9879,N_6159);
nor U14841 (N_14841,N_8522,N_8195);
or U14842 (N_14842,N_5042,N_9310);
or U14843 (N_14843,N_7929,N_7347);
or U14844 (N_14844,N_9983,N_6324);
nor U14845 (N_14845,N_7249,N_5237);
nor U14846 (N_14846,N_6690,N_8658);
nor U14847 (N_14847,N_6252,N_6557);
or U14848 (N_14848,N_8963,N_7352);
nor U14849 (N_14849,N_6430,N_6098);
or U14850 (N_14850,N_8331,N_9705);
nor U14851 (N_14851,N_8548,N_5097);
nor U14852 (N_14852,N_7675,N_5494);
nor U14853 (N_14853,N_8782,N_7202);
nand U14854 (N_14854,N_5446,N_5554);
nor U14855 (N_14855,N_9733,N_5970);
or U14856 (N_14856,N_8949,N_5010);
nor U14857 (N_14857,N_9974,N_5782);
or U14858 (N_14858,N_6191,N_6181);
and U14859 (N_14859,N_8122,N_6544);
nor U14860 (N_14860,N_9469,N_8388);
nand U14861 (N_14861,N_9896,N_7380);
nand U14862 (N_14862,N_8351,N_9174);
nor U14863 (N_14863,N_6239,N_8705);
nor U14864 (N_14864,N_6468,N_6512);
or U14865 (N_14865,N_7672,N_8130);
nand U14866 (N_14866,N_8029,N_8375);
nand U14867 (N_14867,N_9027,N_6130);
nand U14868 (N_14868,N_8949,N_8116);
and U14869 (N_14869,N_8012,N_9125);
nand U14870 (N_14870,N_8106,N_9772);
nand U14871 (N_14871,N_8244,N_6690);
xor U14872 (N_14872,N_8603,N_9660);
and U14873 (N_14873,N_5182,N_6534);
and U14874 (N_14874,N_7261,N_5117);
nor U14875 (N_14875,N_8428,N_7758);
nand U14876 (N_14876,N_7818,N_6026);
or U14877 (N_14877,N_8979,N_5334);
nand U14878 (N_14878,N_7791,N_7265);
nand U14879 (N_14879,N_8178,N_8904);
and U14880 (N_14880,N_6168,N_8951);
nand U14881 (N_14881,N_5046,N_9730);
nor U14882 (N_14882,N_6742,N_9872);
nand U14883 (N_14883,N_6688,N_5504);
nor U14884 (N_14884,N_6363,N_7762);
nor U14885 (N_14885,N_6697,N_9602);
and U14886 (N_14886,N_9452,N_5384);
nor U14887 (N_14887,N_8536,N_9248);
and U14888 (N_14888,N_6081,N_8671);
and U14889 (N_14889,N_9961,N_6473);
nor U14890 (N_14890,N_5880,N_9645);
nand U14891 (N_14891,N_5104,N_6134);
nand U14892 (N_14892,N_8222,N_9885);
nor U14893 (N_14893,N_7489,N_5068);
nand U14894 (N_14894,N_8281,N_7427);
nand U14895 (N_14895,N_8132,N_6037);
nor U14896 (N_14896,N_7756,N_7844);
or U14897 (N_14897,N_7631,N_9862);
nand U14898 (N_14898,N_6919,N_6015);
nand U14899 (N_14899,N_8811,N_8796);
nand U14900 (N_14900,N_8541,N_6051);
nand U14901 (N_14901,N_9474,N_6734);
nand U14902 (N_14902,N_6196,N_7293);
nor U14903 (N_14903,N_8676,N_9266);
nand U14904 (N_14904,N_8112,N_5668);
and U14905 (N_14905,N_8692,N_8588);
or U14906 (N_14906,N_5448,N_6352);
nor U14907 (N_14907,N_6291,N_7949);
or U14908 (N_14908,N_6896,N_5866);
or U14909 (N_14909,N_9933,N_8653);
and U14910 (N_14910,N_7001,N_5261);
nor U14911 (N_14911,N_7812,N_5797);
and U14912 (N_14912,N_8422,N_8372);
nor U14913 (N_14913,N_5716,N_8013);
nor U14914 (N_14914,N_9253,N_6385);
nor U14915 (N_14915,N_8032,N_7025);
nand U14916 (N_14916,N_8649,N_6426);
and U14917 (N_14917,N_6622,N_8050);
nor U14918 (N_14918,N_8539,N_5128);
nand U14919 (N_14919,N_9261,N_6218);
or U14920 (N_14920,N_5867,N_6474);
nand U14921 (N_14921,N_8508,N_5102);
nand U14922 (N_14922,N_7040,N_7454);
and U14923 (N_14923,N_7930,N_7462);
or U14924 (N_14924,N_8742,N_6768);
nor U14925 (N_14925,N_5905,N_6067);
nand U14926 (N_14926,N_7698,N_8902);
nor U14927 (N_14927,N_6601,N_7125);
nor U14928 (N_14928,N_5035,N_9638);
or U14929 (N_14929,N_7907,N_6942);
nand U14930 (N_14930,N_5407,N_9420);
and U14931 (N_14931,N_8846,N_9259);
nor U14932 (N_14932,N_8823,N_7808);
nand U14933 (N_14933,N_8806,N_8990);
nor U14934 (N_14934,N_5949,N_5023);
or U14935 (N_14935,N_5284,N_6128);
nand U14936 (N_14936,N_5330,N_8683);
or U14937 (N_14937,N_6237,N_8141);
or U14938 (N_14938,N_7131,N_8679);
nor U14939 (N_14939,N_8653,N_7988);
and U14940 (N_14940,N_7046,N_9379);
nor U14941 (N_14941,N_9901,N_8361);
nand U14942 (N_14942,N_7116,N_7798);
or U14943 (N_14943,N_7884,N_7846);
nor U14944 (N_14944,N_8326,N_7693);
nand U14945 (N_14945,N_7974,N_9707);
or U14946 (N_14946,N_5334,N_8711);
nor U14947 (N_14947,N_8022,N_8594);
nand U14948 (N_14948,N_9276,N_6967);
nand U14949 (N_14949,N_9922,N_5738);
nor U14950 (N_14950,N_6483,N_8858);
nor U14951 (N_14951,N_7550,N_7014);
nand U14952 (N_14952,N_7690,N_8939);
nand U14953 (N_14953,N_9229,N_5703);
nand U14954 (N_14954,N_7918,N_5929);
nor U14955 (N_14955,N_6940,N_9812);
nor U14956 (N_14956,N_6671,N_8401);
or U14957 (N_14957,N_7670,N_6746);
nand U14958 (N_14958,N_6148,N_8027);
and U14959 (N_14959,N_7168,N_9111);
nand U14960 (N_14960,N_9742,N_9850);
nor U14961 (N_14961,N_6565,N_8040);
nand U14962 (N_14962,N_5458,N_9785);
nor U14963 (N_14963,N_6374,N_7975);
nor U14964 (N_14964,N_5646,N_6112);
nor U14965 (N_14965,N_6603,N_6906);
or U14966 (N_14966,N_8150,N_6196);
nor U14967 (N_14967,N_6904,N_9168);
or U14968 (N_14968,N_5319,N_8137);
and U14969 (N_14969,N_8540,N_8488);
and U14970 (N_14970,N_7457,N_6765);
or U14971 (N_14971,N_7694,N_9604);
and U14972 (N_14972,N_9218,N_9464);
nand U14973 (N_14973,N_8814,N_9129);
and U14974 (N_14974,N_8222,N_6820);
and U14975 (N_14975,N_7579,N_7931);
and U14976 (N_14976,N_8866,N_6233);
and U14977 (N_14977,N_9305,N_6829);
nand U14978 (N_14978,N_5066,N_7704);
nand U14979 (N_14979,N_6304,N_5675);
nor U14980 (N_14980,N_6739,N_5406);
nor U14981 (N_14981,N_5682,N_9940);
or U14982 (N_14982,N_5054,N_6156);
nor U14983 (N_14983,N_5268,N_7968);
nand U14984 (N_14984,N_9862,N_5222);
nor U14985 (N_14985,N_9540,N_7083);
or U14986 (N_14986,N_5968,N_8141);
nor U14987 (N_14987,N_5383,N_9487);
or U14988 (N_14988,N_8514,N_9923);
nor U14989 (N_14989,N_9645,N_9245);
or U14990 (N_14990,N_5264,N_8690);
or U14991 (N_14991,N_9172,N_7131);
and U14992 (N_14992,N_7123,N_7660);
nand U14993 (N_14993,N_6545,N_7135);
or U14994 (N_14994,N_6415,N_5201);
or U14995 (N_14995,N_8103,N_6392);
xnor U14996 (N_14996,N_7731,N_8792);
nor U14997 (N_14997,N_9398,N_6260);
nand U14998 (N_14998,N_5638,N_8493);
nand U14999 (N_14999,N_6879,N_8551);
or UO_0 (O_0,N_11287,N_10650);
nand UO_1 (O_1,N_11171,N_12642);
nand UO_2 (O_2,N_11490,N_13996);
nor UO_3 (O_3,N_12607,N_11911);
nor UO_4 (O_4,N_10173,N_13054);
and UO_5 (O_5,N_12059,N_12131);
nor UO_6 (O_6,N_11099,N_13953);
and UO_7 (O_7,N_11964,N_12898);
or UO_8 (O_8,N_12198,N_12687);
or UO_9 (O_9,N_14229,N_11571);
and UO_10 (O_10,N_13278,N_12044);
nand UO_11 (O_11,N_14463,N_10192);
nor UO_12 (O_12,N_10344,N_11149);
or UO_13 (O_13,N_10047,N_14163);
and UO_14 (O_14,N_11644,N_10203);
nand UO_15 (O_15,N_12956,N_10868);
nor UO_16 (O_16,N_10652,N_13734);
nor UO_17 (O_17,N_13992,N_14625);
and UO_18 (O_18,N_11971,N_11085);
and UO_19 (O_19,N_10582,N_14742);
nor UO_20 (O_20,N_12285,N_10918);
nor UO_21 (O_21,N_10766,N_12776);
and UO_22 (O_22,N_12424,N_10338);
nand UO_23 (O_23,N_12186,N_11892);
nand UO_24 (O_24,N_10842,N_14503);
or UO_25 (O_25,N_11973,N_13473);
nand UO_26 (O_26,N_10887,N_13338);
and UO_27 (O_27,N_11422,N_13907);
nor UO_28 (O_28,N_14725,N_11703);
nand UO_29 (O_29,N_12858,N_11044);
or UO_30 (O_30,N_14111,N_11706);
nor UO_31 (O_31,N_10520,N_12705);
nor UO_32 (O_32,N_13335,N_14487);
nor UO_33 (O_33,N_10911,N_12148);
xor UO_34 (O_34,N_11327,N_12461);
nand UO_35 (O_35,N_14181,N_10053);
and UO_36 (O_36,N_11531,N_10783);
nor UO_37 (O_37,N_10011,N_12241);
or UO_38 (O_38,N_12344,N_14902);
nor UO_39 (O_39,N_10807,N_13920);
nand UO_40 (O_40,N_10443,N_12791);
or UO_41 (O_41,N_10504,N_14031);
and UO_42 (O_42,N_13990,N_12287);
or UO_43 (O_43,N_11557,N_14046);
or UO_44 (O_44,N_13056,N_12158);
nor UO_45 (O_45,N_12874,N_13080);
or UO_46 (O_46,N_11834,N_10681);
nor UO_47 (O_47,N_10050,N_13847);
or UO_48 (O_48,N_14235,N_13012);
nor UO_49 (O_49,N_13523,N_11204);
or UO_50 (O_50,N_13120,N_14314);
or UO_51 (O_51,N_10406,N_12740);
and UO_52 (O_52,N_13937,N_10511);
or UO_53 (O_53,N_11712,N_12704);
nand UO_54 (O_54,N_13709,N_10424);
or UO_55 (O_55,N_12384,N_11846);
xnor UO_56 (O_56,N_13194,N_10316);
and UO_57 (O_57,N_12267,N_11297);
nand UO_58 (O_58,N_10874,N_11966);
nor UO_59 (O_59,N_11745,N_14696);
and UO_60 (O_60,N_12895,N_12093);
nand UO_61 (O_61,N_10724,N_11372);
nor UO_62 (O_62,N_10866,N_14521);
and UO_63 (O_63,N_14849,N_12981);
or UO_64 (O_64,N_10353,N_13133);
and UO_65 (O_65,N_13929,N_11123);
or UO_66 (O_66,N_14177,N_10917);
or UO_67 (O_67,N_14873,N_14891);
nor UO_68 (O_68,N_12659,N_14093);
nor UO_69 (O_69,N_14722,N_13893);
and UO_70 (O_70,N_12584,N_14472);
and UO_71 (O_71,N_10749,N_14476);
and UO_72 (O_72,N_11690,N_14126);
nor UO_73 (O_73,N_11033,N_11214);
nand UO_74 (O_74,N_11254,N_13565);
xnor UO_75 (O_75,N_12069,N_14278);
nand UO_76 (O_76,N_10287,N_12410);
nor UO_77 (O_77,N_12798,N_11489);
and UO_78 (O_78,N_10544,N_11616);
nor UO_79 (O_79,N_13817,N_10666);
nand UO_80 (O_80,N_10243,N_14395);
and UO_81 (O_81,N_13468,N_12645);
and UO_82 (O_82,N_12989,N_14005);
nor UO_83 (O_83,N_14867,N_12819);
nor UO_84 (O_84,N_12019,N_13557);
and UO_85 (O_85,N_11007,N_10389);
nor UO_86 (O_86,N_10375,N_10909);
nor UO_87 (O_87,N_13906,N_12516);
nor UO_88 (O_88,N_13434,N_14875);
and UO_89 (O_89,N_11987,N_13222);
nand UO_90 (O_90,N_12374,N_11244);
nor UO_91 (O_91,N_10997,N_14378);
and UO_92 (O_92,N_11350,N_10041);
nand UO_93 (O_93,N_11707,N_10065);
or UO_94 (O_94,N_12153,N_13266);
or UO_95 (O_95,N_12234,N_12112);
nand UO_96 (O_96,N_11437,N_14876);
and UO_97 (O_97,N_12110,N_13437);
nor UO_98 (O_98,N_13701,N_10174);
and UO_99 (O_99,N_11855,N_14890);
and UO_100 (O_100,N_10518,N_13615);
nand UO_101 (O_101,N_11116,N_12692);
nor UO_102 (O_102,N_11902,N_10605);
nor UO_103 (O_103,N_13533,N_11511);
and UO_104 (O_104,N_12454,N_11808);
nand UO_105 (O_105,N_14652,N_14604);
nor UO_106 (O_106,N_13454,N_13551);
or UO_107 (O_107,N_10221,N_12312);
nand UO_108 (O_108,N_11818,N_11110);
and UO_109 (O_109,N_10527,N_14069);
and UO_110 (O_110,N_10610,N_11551);
or UO_111 (O_111,N_10684,N_13935);
and UO_112 (O_112,N_10165,N_12191);
nand UO_113 (O_113,N_14247,N_11603);
and UO_114 (O_114,N_14335,N_14736);
or UO_115 (O_115,N_11972,N_14948);
nand UO_116 (O_116,N_12724,N_12385);
nor UO_117 (O_117,N_13349,N_12929);
nand UO_118 (O_118,N_11330,N_12465);
or UO_119 (O_119,N_10811,N_13573);
or UO_120 (O_120,N_13553,N_11383);
nand UO_121 (O_121,N_14915,N_14687);
or UO_122 (O_122,N_14405,N_14071);
and UO_123 (O_123,N_14889,N_12006);
nand UO_124 (O_124,N_13544,N_13815);
nor UO_125 (O_125,N_13518,N_10356);
nor UO_126 (O_126,N_11505,N_14998);
nand UO_127 (O_127,N_14318,N_10642);
nand UO_128 (O_128,N_11715,N_10071);
nor UO_129 (O_129,N_14353,N_12202);
or UO_130 (O_130,N_11311,N_13035);
and UO_131 (O_131,N_10458,N_13084);
nand UO_132 (O_132,N_10034,N_12435);
or UO_133 (O_133,N_10562,N_12652);
nand UO_134 (O_134,N_11938,N_12715);
nor UO_135 (O_135,N_12595,N_11431);
or UO_136 (O_136,N_12327,N_11402);
nor UO_137 (O_137,N_13968,N_11692);
and UO_138 (O_138,N_13407,N_12236);
or UO_139 (O_139,N_12095,N_12007);
or UO_140 (O_140,N_10004,N_12275);
nor UO_141 (O_141,N_11373,N_13641);
and UO_142 (O_142,N_13424,N_12184);
nand UO_143 (O_143,N_10485,N_11433);
nor UO_144 (O_144,N_10301,N_14106);
nand UO_145 (O_145,N_13303,N_14439);
nor UO_146 (O_146,N_11849,N_11087);
and UO_147 (O_147,N_10095,N_10154);
nand UO_148 (O_148,N_13810,N_12086);
and UO_149 (O_149,N_10627,N_11702);
nand UO_150 (O_150,N_14061,N_11436);
nand UO_151 (O_151,N_11182,N_13017);
or UO_152 (O_152,N_14465,N_10029);
or UO_153 (O_153,N_14404,N_14790);
nor UO_154 (O_154,N_14598,N_12179);
or UO_155 (O_155,N_10619,N_14938);
or UO_156 (O_156,N_12180,N_14081);
or UO_157 (O_157,N_12683,N_14008);
nand UO_158 (O_158,N_11251,N_13825);
or UO_159 (O_159,N_13046,N_11158);
nand UO_160 (O_160,N_10200,N_13831);
nor UO_161 (O_161,N_14004,N_13258);
nand UO_162 (O_162,N_10100,N_11376);
xor UO_163 (O_163,N_11861,N_10415);
nand UO_164 (O_164,N_14735,N_13886);
nand UO_165 (O_165,N_12310,N_10594);
nand UO_166 (O_166,N_14509,N_10473);
nand UO_167 (O_167,N_10372,N_10856);
and UO_168 (O_168,N_13100,N_13652);
and UO_169 (O_169,N_13461,N_11624);
or UO_170 (O_170,N_13376,N_11065);
nand UO_171 (O_171,N_14574,N_10283);
and UO_172 (O_172,N_10324,N_12885);
and UO_173 (O_173,N_12482,N_10555);
nor UO_174 (O_174,N_13070,N_10757);
or UO_175 (O_175,N_13067,N_13366);
nor UO_176 (O_176,N_12458,N_13803);
nand UO_177 (O_177,N_13691,N_11732);
nand UO_178 (O_178,N_10347,N_12300);
and UO_179 (O_179,N_13238,N_10576);
xnor UO_180 (O_180,N_11225,N_14198);
and UO_181 (O_181,N_13945,N_12398);
nor UO_182 (O_182,N_10869,N_11890);
and UO_183 (O_183,N_10699,N_11819);
nor UO_184 (O_184,N_11396,N_11628);
and UO_185 (O_185,N_10566,N_12864);
or UO_186 (O_186,N_13524,N_13208);
and UO_187 (O_187,N_12205,N_14881);
or UO_188 (O_188,N_12262,N_12831);
and UO_189 (O_189,N_11039,N_11443);
and UO_190 (O_190,N_10878,N_12544);
nor UO_191 (O_191,N_13268,N_10785);
or UO_192 (O_192,N_10569,N_12916);
nor UO_193 (O_193,N_11111,N_14223);
nor UO_194 (O_194,N_14820,N_14263);
nand UO_195 (O_195,N_12115,N_12338);
nor UO_196 (O_196,N_14689,N_14775);
nor UO_197 (O_197,N_12391,N_12486);
nand UO_198 (O_198,N_10252,N_12045);
nor UO_199 (O_199,N_13542,N_14603);
and UO_200 (O_200,N_13209,N_14110);
nand UO_201 (O_201,N_14317,N_14549);
and UO_202 (O_202,N_12272,N_14923);
and UO_203 (O_203,N_10275,N_12032);
nand UO_204 (O_204,N_10147,N_10908);
nand UO_205 (O_205,N_10967,N_11174);
nor UO_206 (O_206,N_10841,N_11594);
nor UO_207 (O_207,N_11992,N_10467);
or UO_208 (O_208,N_10670,N_12558);
or UO_209 (O_209,N_14442,N_11030);
nand UO_210 (O_210,N_12547,N_13939);
or UO_211 (O_211,N_11345,N_13055);
and UO_212 (O_212,N_12809,N_11854);
and UO_213 (O_213,N_11169,N_11078);
or UO_214 (O_214,N_13746,N_11960);
and UO_215 (O_215,N_13900,N_14692);
nand UO_216 (O_216,N_14070,N_14878);
and UO_217 (O_217,N_14011,N_10806);
nand UO_218 (O_218,N_12713,N_14690);
nand UO_219 (O_219,N_12256,N_10452);
and UO_220 (O_220,N_10169,N_12484);
and UO_221 (O_221,N_13173,N_13879);
or UO_222 (O_222,N_13739,N_12756);
and UO_223 (O_223,N_14467,N_11893);
nand UO_224 (O_224,N_14863,N_14744);
or UO_225 (O_225,N_12507,N_11500);
nor UO_226 (O_226,N_13058,N_10059);
nand UO_227 (O_227,N_12274,N_12985);
or UO_228 (O_228,N_13282,N_10108);
and UO_229 (O_229,N_10431,N_10257);
nand UO_230 (O_230,N_12644,N_14806);
nor UO_231 (O_231,N_12416,N_13806);
nand UO_232 (O_232,N_13769,N_14363);
or UO_233 (O_233,N_10278,N_13586);
or UO_234 (O_234,N_13675,N_14786);
or UO_235 (O_235,N_13203,N_12536);
nand UO_236 (O_236,N_11572,N_12141);
or UO_237 (O_237,N_11922,N_10012);
xor UO_238 (O_238,N_12915,N_13978);
xnor UO_239 (O_239,N_11979,N_14771);
nor UO_240 (O_240,N_14075,N_14436);
or UO_241 (O_241,N_10982,N_10947);
nand UO_242 (O_242,N_10737,N_13529);
and UO_243 (O_243,N_10360,N_10560);
and UO_244 (O_244,N_13711,N_10337);
or UO_245 (O_245,N_12297,N_10744);
nor UO_246 (O_246,N_10726,N_14906);
or UO_247 (O_247,N_12075,N_13995);
or UO_248 (O_248,N_13587,N_12015);
nand UO_249 (O_249,N_14033,N_11999);
nand UO_250 (O_250,N_10098,N_14481);
nor UO_251 (O_251,N_14695,N_10710);
and UO_252 (O_252,N_14566,N_13983);
and UO_253 (O_253,N_12639,N_13311);
nand UO_254 (O_254,N_12364,N_10671);
and UO_255 (O_255,N_10027,N_10043);
or UO_256 (O_256,N_11850,N_14458);
and UO_257 (O_257,N_13220,N_14675);
nand UO_258 (O_258,N_10035,N_11006);
nor UO_259 (O_259,N_13211,N_11894);
and UO_260 (O_260,N_13325,N_13917);
or UO_261 (O_261,N_11982,N_13805);
and UO_262 (O_262,N_11454,N_14864);
or UO_263 (O_263,N_11659,N_14698);
or UO_264 (O_264,N_14200,N_13576);
and UO_265 (O_265,N_12942,N_11643);
and UO_266 (O_266,N_10274,N_11568);
nand UO_267 (O_267,N_10591,N_14387);
nand UO_268 (O_268,N_11695,N_10224);
nand UO_269 (O_269,N_10077,N_13853);
or UO_270 (O_270,N_10408,N_12406);
nand UO_271 (O_271,N_12650,N_13766);
nand UO_272 (O_272,N_10531,N_11167);
nand UO_273 (O_273,N_14469,N_11828);
or UO_274 (O_274,N_11951,N_13247);
xnor UO_275 (O_275,N_13490,N_12829);
nand UO_276 (O_276,N_13638,N_14269);
nand UO_277 (O_277,N_11374,N_10730);
nor UO_278 (O_278,N_12210,N_11259);
or UO_279 (O_279,N_12701,N_10371);
and UO_280 (O_280,N_13854,N_12280);
nor UO_281 (O_281,N_12330,N_10793);
and UO_282 (O_282,N_12031,N_12407);
nand UO_283 (O_283,N_14173,N_12881);
nand UO_284 (O_284,N_10510,N_14019);
nand UO_285 (O_285,N_13657,N_13154);
nand UO_286 (O_286,N_14136,N_13840);
nor UO_287 (O_287,N_12096,N_10404);
and UO_288 (O_288,N_13808,N_13137);
or UO_289 (O_289,N_12358,N_11115);
or UO_290 (O_290,N_12042,N_14840);
or UO_291 (O_291,N_11426,N_12087);
nor UO_292 (O_292,N_13037,N_13126);
nand UO_293 (O_293,N_11965,N_10623);
nand UO_294 (O_294,N_14874,N_11170);
nor UO_295 (O_295,N_10139,N_12303);
and UO_296 (O_296,N_11636,N_14280);
nor UO_297 (O_297,N_14538,N_10378);
nor UO_298 (O_298,N_13453,N_11637);
nand UO_299 (O_299,N_12356,N_12654);
or UO_300 (O_300,N_12538,N_13663);
nor UO_301 (O_301,N_11660,N_10326);
xnor UO_302 (O_302,N_12611,N_11059);
and UO_303 (O_303,N_14795,N_10926);
and UO_304 (O_304,N_12412,N_13728);
or UO_305 (O_305,N_13412,N_11632);
nand UO_306 (O_306,N_12508,N_10630);
nand UO_307 (O_307,N_11755,N_10864);
nand UO_308 (O_308,N_14723,N_11506);
or UO_309 (O_309,N_10541,N_12602);
nor UO_310 (O_310,N_10172,N_11219);
nor UO_311 (O_311,N_12306,N_13799);
nand UO_312 (O_312,N_10548,N_12389);
nor UO_313 (O_313,N_12387,N_12512);
and UO_314 (O_314,N_13789,N_14780);
nor UO_315 (O_315,N_10872,N_10604);
nand UO_316 (O_316,N_12835,N_13399);
nand UO_317 (O_317,N_14374,N_11309);
or UO_318 (O_318,N_10660,N_11203);
nor UO_319 (O_319,N_14792,N_11790);
and UO_320 (O_320,N_11701,N_10054);
and UO_321 (O_321,N_14379,N_11963);
nor UO_322 (O_322,N_14016,N_13098);
and UO_323 (O_323,N_12166,N_11625);
nand UO_324 (O_324,N_14298,N_10417);
nor UO_325 (O_325,N_13949,N_11710);
nor UO_326 (O_326,N_14933,N_13109);
and UO_327 (O_327,N_11906,N_11190);
nand UO_328 (O_328,N_12397,N_13578);
and UO_329 (O_329,N_11887,N_14715);
and UO_330 (O_330,N_12647,N_10786);
nand UO_331 (O_331,N_13672,N_14919);
nand UO_332 (O_332,N_12729,N_13870);
nand UO_333 (O_333,N_13319,N_14921);
or UO_334 (O_334,N_12730,N_11598);
nor UO_335 (O_335,N_12711,N_12760);
nand UO_336 (O_336,N_10564,N_12905);
nor UO_337 (O_337,N_10542,N_11763);
nand UO_338 (O_338,N_11026,N_14709);
nor UO_339 (O_339,N_12553,N_14900);
nor UO_340 (O_340,N_14757,N_13823);
or UO_341 (O_341,N_13302,N_11492);
or UO_342 (O_342,N_10055,N_10537);
or UO_343 (O_343,N_12244,N_11985);
or UO_344 (O_344,N_12057,N_14804);
and UO_345 (O_345,N_14410,N_13448);
and UO_346 (O_346,N_13654,N_11853);
or UO_347 (O_347,N_10130,N_14309);
nor UO_348 (O_348,N_11546,N_14697);
and UO_349 (O_349,N_12493,N_12009);
nand UO_350 (O_350,N_12626,N_11407);
and UO_351 (O_351,N_10157,N_11576);
or UO_352 (O_352,N_10668,N_10899);
and UO_353 (O_353,N_11184,N_13300);
nor UO_354 (O_354,N_14785,N_11786);
and UO_355 (O_355,N_11682,N_12106);
and UO_356 (O_356,N_14428,N_11406);
or UO_357 (O_357,N_13198,N_13132);
nor UO_358 (O_358,N_12071,N_10675);
or UO_359 (O_359,N_13610,N_14265);
and UO_360 (O_360,N_12296,N_10302);
nand UO_361 (O_361,N_13758,N_10507);
or UO_362 (O_362,N_10683,N_13487);
nand UO_363 (O_363,N_10954,N_14770);
and UO_364 (O_364,N_12780,N_10184);
and UO_365 (O_365,N_11294,N_12594);
or UO_366 (O_366,N_13871,N_11118);
nand UO_367 (O_367,N_14519,N_14951);
and UO_368 (O_368,N_11410,N_11959);
and UO_369 (O_369,N_10898,N_11769);
nor UO_370 (O_370,N_10770,N_14327);
xnor UO_371 (O_371,N_12961,N_12927);
nor UO_372 (O_372,N_12257,N_12997);
or UO_373 (O_373,N_13496,N_11548);
or UO_374 (O_374,N_11375,N_10391);
and UO_375 (O_375,N_11439,N_11575);
or UO_376 (O_376,N_12965,N_14164);
xnor UO_377 (O_377,N_11235,N_11897);
nand UO_378 (O_378,N_10804,N_13633);
nand UO_379 (O_379,N_14289,N_14520);
and UO_380 (O_380,N_14291,N_14669);
nand UO_381 (O_381,N_13406,N_13076);
or UO_382 (O_382,N_11322,N_14120);
or UO_383 (O_383,N_11106,N_14040);
and UO_384 (O_384,N_10885,N_11621);
and UO_385 (O_385,N_10019,N_10538);
and UO_386 (O_386,N_11720,N_10386);
nor UO_387 (O_387,N_14774,N_12359);
nand UO_388 (O_388,N_12233,N_10112);
and UO_389 (O_389,N_11619,N_12868);
and UO_390 (O_390,N_10118,N_14674);
and UO_391 (O_391,N_12919,N_10494);
nor UO_392 (O_392,N_14232,N_10107);
nand UO_393 (O_393,N_12608,N_11403);
nor UO_394 (O_394,N_13296,N_14172);
nand UO_395 (O_395,N_10902,N_11343);
or UO_396 (O_396,N_13536,N_10575);
nor UO_397 (O_397,N_12987,N_11234);
and UO_398 (O_398,N_10953,N_13494);
nor UO_399 (O_399,N_11891,N_10478);
nor UO_400 (O_400,N_10444,N_13892);
or UO_401 (O_401,N_11515,N_13230);
nand UO_402 (O_402,N_12268,N_11095);
nand UO_403 (O_403,N_14313,N_12160);
nor UO_404 (O_404,N_10709,N_13057);
nor UO_405 (O_405,N_13234,N_14992);
and UO_406 (O_406,N_14745,N_13770);
nand UO_407 (O_407,N_10940,N_10113);
or UO_408 (O_408,N_10592,N_14788);
or UO_409 (O_409,N_10426,N_12423);
nand UO_410 (O_410,N_13271,N_12081);
nor UO_411 (O_411,N_13495,N_13326);
and UO_412 (O_412,N_11997,N_14386);
nor UO_413 (O_413,N_10839,N_11495);
and UO_414 (O_414,N_11599,N_11336);
nor UO_415 (O_415,N_13219,N_12053);
nor UO_416 (O_416,N_11884,N_10574);
or UO_417 (O_417,N_11043,N_12549);
nand UO_418 (O_418,N_12795,N_11306);
nand UO_419 (O_419,N_14734,N_14304);
nand UO_420 (O_420,N_12865,N_11542);
or UO_421 (O_421,N_14225,N_14322);
or UO_422 (O_422,N_12746,N_11928);
or UO_423 (O_423,N_10472,N_12646);
nand UO_424 (O_424,N_13567,N_11880);
nor UO_425 (O_425,N_10127,N_12316);
nand UO_426 (O_426,N_13186,N_10907);
or UO_427 (O_427,N_13753,N_11121);
or UO_428 (O_428,N_11829,N_10428);
nor UO_429 (O_429,N_14577,N_12853);
and UO_430 (O_430,N_10125,N_13855);
and UO_431 (O_431,N_10232,N_11477);
nand UO_432 (O_432,N_14294,N_10912);
or UO_433 (O_433,N_14147,N_12278);
nor UO_434 (O_434,N_14018,N_14001);
or UO_435 (O_435,N_10821,N_14594);
nand UO_436 (O_436,N_13379,N_12900);
or UO_437 (O_437,N_10006,N_13446);
or UO_438 (O_438,N_12621,N_11215);
or UO_439 (O_439,N_10495,N_13779);
or UO_440 (O_440,N_11937,N_11385);
nor UO_441 (O_441,N_10105,N_12737);
nand UO_442 (O_442,N_12008,N_13738);
and UO_443 (O_443,N_13862,N_10245);
nor UO_444 (O_444,N_10291,N_11771);
nor UO_445 (O_445,N_12415,N_13092);
nand UO_446 (O_446,N_13874,N_12792);
and UO_447 (O_447,N_11040,N_10355);
or UO_448 (O_448,N_10400,N_12666);
or UO_449 (O_449,N_14370,N_14989);
and UO_450 (O_450,N_12567,N_10010);
nor UO_451 (O_451,N_13526,N_12311);
or UO_452 (O_452,N_14391,N_13780);
or UO_453 (O_453,N_14582,N_11393);
nor UO_454 (O_454,N_10844,N_13532);
nor UO_455 (O_455,N_13015,N_11113);
nand UO_456 (O_456,N_12675,N_14726);
or UO_457 (O_457,N_13605,N_10568);
nand UO_458 (O_458,N_12703,N_12640);
nand UO_459 (O_459,N_13032,N_14375);
nor UO_460 (O_460,N_12313,N_11936);
or UO_461 (O_461,N_11986,N_11479);
nand UO_462 (O_462,N_14344,N_13510);
nor UO_463 (O_463,N_14552,N_12432);
or UO_464 (O_464,N_12943,N_11315);
nor UO_465 (O_465,N_11057,N_14234);
nand UO_466 (O_466,N_11995,N_11222);
nor UO_467 (O_467,N_14022,N_12510);
nand UO_468 (O_468,N_12249,N_11905);
nand UO_469 (O_469,N_11451,N_14202);
xnor UO_470 (O_470,N_12206,N_14107);
nor UO_471 (O_471,N_14168,N_10694);
nor UO_472 (O_472,N_13818,N_11248);
nor UO_473 (O_473,N_13981,N_13118);
and UO_474 (O_474,N_10137,N_14239);
nor UO_475 (O_475,N_11940,N_13351);
nand UO_476 (O_476,N_13373,N_14080);
and UO_477 (O_477,N_14909,N_10539);
or UO_478 (O_478,N_12734,N_13139);
or UO_479 (O_479,N_10817,N_13398);
or UO_480 (O_480,N_12863,N_13069);
or UO_481 (O_481,N_13890,N_11411);
nand UO_482 (O_482,N_12719,N_14418);
or UO_483 (O_483,N_11283,N_10973);
nand UO_484 (O_484,N_11915,N_11080);
and UO_485 (O_485,N_10076,N_13506);
nand UO_486 (O_486,N_13287,N_14051);
nand UO_487 (O_487,N_11475,N_10923);
and UO_488 (O_488,N_11899,N_11726);
nor UO_489 (O_489,N_11930,N_10655);
nor UO_490 (O_490,N_14079,N_13571);
xor UO_491 (O_491,N_14017,N_13635);
or UO_492 (O_492,N_12419,N_11014);
nand UO_493 (O_493,N_13647,N_12260);
xor UO_494 (O_494,N_11989,N_10719);
and UO_495 (O_495,N_12321,N_10771);
or UO_496 (O_496,N_11669,N_13471);
nor UO_497 (O_497,N_14869,N_14701);
and UO_498 (O_498,N_14296,N_10981);
nand UO_499 (O_499,N_10731,N_10455);
and UO_500 (O_500,N_10074,N_14224);
or UO_501 (O_501,N_10760,N_13721);
nor UO_502 (O_502,N_11307,N_11811);
and UO_503 (O_503,N_14994,N_14209);
nand UO_504 (O_504,N_13987,N_11245);
nor UO_505 (O_505,N_13798,N_13408);
or UO_506 (O_506,N_14609,N_12147);
and UO_507 (O_507,N_11626,N_13707);
nand UO_508 (O_508,N_14116,N_11381);
nor UO_509 (O_509,N_13600,N_11198);
nor UO_510 (O_510,N_12661,N_12264);
nor UO_511 (O_511,N_12967,N_12789);
nand UO_512 (O_512,N_12177,N_11998);
or UO_513 (O_513,N_13090,N_11466);
and UO_514 (O_514,N_13322,N_11662);
nand UO_515 (O_515,N_14233,N_12337);
nor UO_516 (O_516,N_14750,N_12823);
or UO_517 (O_517,N_10342,N_14255);
nand UO_518 (O_518,N_12699,N_14610);
or UO_519 (O_519,N_11197,N_10672);
nand UO_520 (O_520,N_12347,N_14781);
nand UO_521 (O_521,N_12755,N_12794);
and UO_522 (O_522,N_12518,N_10622);
or UO_523 (O_523,N_13748,N_12766);
nor UO_524 (O_524,N_13514,N_13024);
nor UO_525 (O_525,N_10476,N_11614);
nand UO_526 (O_526,N_11883,N_10182);
and UO_527 (O_527,N_10625,N_13370);
nor UO_528 (O_528,N_13259,N_13135);
nand UO_529 (O_529,N_10383,N_12085);
or UO_530 (O_530,N_11879,N_12571);
or UO_531 (O_531,N_12324,N_10734);
and UO_532 (O_532,N_12686,N_14028);
nor UO_533 (O_533,N_13041,N_11770);
nand UO_534 (O_534,N_14602,N_13484);
nand UO_535 (O_535,N_14419,N_14429);
or UO_536 (O_536,N_11832,N_13757);
nand UO_537 (O_537,N_13264,N_14199);
nor UO_538 (O_538,N_13918,N_12909);
nor UO_539 (O_539,N_12497,N_14749);
or UO_540 (O_540,N_13517,N_14708);
nor UO_541 (O_541,N_14451,N_10937);
and UO_542 (O_542,N_14455,N_11996);
nor UO_543 (O_543,N_10003,N_13465);
or UO_544 (O_544,N_13188,N_11063);
and UO_545 (O_545,N_12903,N_11278);
and UO_546 (O_546,N_11131,N_14166);
nand UO_547 (O_547,N_11804,N_10965);
nand UO_548 (O_548,N_11903,N_10618);
nor UO_549 (O_549,N_10206,N_12842);
xnor UO_550 (O_550,N_12718,N_10831);
nor UO_551 (O_551,N_13839,N_12372);
xnor UO_552 (O_552,N_12893,N_12299);
nand UO_553 (O_553,N_13025,N_12560);
nand UO_554 (O_554,N_14980,N_12124);
nor UO_555 (O_555,N_11794,N_14035);
nand UO_556 (O_556,N_11356,N_14393);
nand UO_557 (O_557,N_13679,N_11714);
or UO_558 (O_558,N_10658,N_11036);
nand UO_559 (O_559,N_14895,N_14337);
or UO_560 (O_560,N_13458,N_12872);
nor UO_561 (O_561,N_13556,N_10094);
or UO_562 (O_562,N_14479,N_11363);
nand UO_563 (O_563,N_11200,N_12117);
and UO_564 (O_564,N_12688,N_11268);
or UO_565 (O_565,N_10809,N_12400);
nor UO_566 (O_566,N_12976,N_14787);
or UO_567 (O_567,N_11606,N_11053);
and UO_568 (O_568,N_12098,N_14189);
or UO_569 (O_569,N_14539,N_10269);
nor UO_570 (O_570,N_11767,N_12641);
or UO_571 (O_571,N_13275,N_14212);
or UO_572 (O_572,N_14431,N_14024);
or UO_573 (O_573,N_10889,N_12557);
nor UO_574 (O_574,N_10886,N_13700);
nor UO_575 (O_575,N_14970,N_11502);
or UO_576 (O_576,N_11942,N_12790);
and UO_577 (O_577,N_14532,N_13733);
nand UO_578 (O_578,N_13527,N_11210);
and UO_579 (O_579,N_12759,N_10608);
or UO_580 (O_580,N_13944,N_14956);
and UO_581 (O_581,N_12240,N_12660);
or UO_582 (O_582,N_12357,N_11666);
and UO_583 (O_583,N_12726,N_13593);
and UO_584 (O_584,N_13696,N_10716);
or UO_585 (O_585,N_10585,N_13613);
or UO_586 (O_586,N_14856,N_12801);
nand UO_587 (O_587,N_10171,N_10438);
nor UO_588 (O_588,N_10140,N_13106);
nor UO_589 (O_589,N_10850,N_14416);
nor UO_590 (O_590,N_10432,N_13119);
or UO_591 (O_591,N_14753,N_13380);
nand UO_592 (O_592,N_12103,N_11077);
nor UO_593 (O_593,N_12332,N_12152);
nor UO_594 (O_594,N_14184,N_12975);
or UO_595 (O_595,N_10867,N_10497);
and UO_596 (O_596,N_10776,N_11954);
or UO_597 (O_597,N_14169,N_10161);
or UO_598 (O_598,N_10180,N_10546);
nor UO_599 (O_599,N_14800,N_10999);
nor UO_600 (O_600,N_13156,N_12906);
and UO_601 (O_601,N_11471,N_14302);
nand UO_602 (O_602,N_13229,N_12761);
nor UO_603 (O_603,N_13143,N_13440);
nor UO_604 (O_604,N_12343,N_11062);
nor UO_605 (O_605,N_10039,N_11877);
nor UO_606 (O_606,N_12388,N_12922);
nor UO_607 (O_607,N_14424,N_14557);
or UO_608 (O_608,N_11747,N_14086);
nor UO_609 (O_609,N_11323,N_12473);
and UO_610 (O_610,N_12521,N_11369);
or UO_611 (O_611,N_10032,N_14991);
or UO_612 (O_612,N_11773,N_14884);
nor UO_613 (O_613,N_11634,N_14480);
nand UO_614 (O_614,N_14510,N_14121);
nor UO_615 (O_615,N_14243,N_11961);
nand UO_616 (O_616,N_10995,N_14118);
and UO_617 (O_617,N_13947,N_10549);
and UO_618 (O_618,N_13888,N_11852);
nand UO_619 (O_619,N_13813,N_14185);
nand UO_620 (O_620,N_12481,N_10052);
nor UO_621 (O_621,N_12744,N_10922);
and UO_622 (O_622,N_14947,N_10031);
or UO_623 (O_623,N_12248,N_13082);
nor UO_624 (O_624,N_10341,N_13620);
nand UO_625 (O_625,N_11047,N_13217);
nand UO_626 (O_626,N_12774,N_11814);
or UO_627 (O_627,N_13970,N_12392);
and UO_628 (O_628,N_13348,N_14127);
nor UO_629 (O_629,N_14897,N_12505);
and UO_630 (O_630,N_12772,N_13612);
and UO_631 (O_631,N_11579,N_12702);
nand UO_632 (O_632,N_12000,N_13105);
or UO_633 (O_633,N_11013,N_10398);
or UO_634 (O_634,N_14426,N_14829);
and UO_635 (O_635,N_14534,N_13162);
nor UO_636 (O_636,N_14411,N_12690);
and UO_637 (O_637,N_14073,N_14142);
and UO_638 (O_638,N_13552,N_14963);
nand UO_639 (O_639,N_10246,N_14694);
or UO_640 (O_640,N_14050,N_11812);
and UO_641 (O_641,N_14977,N_14935);
or UO_642 (O_642,N_10732,N_11484);
nand UO_643 (O_643,N_14733,N_14684);
xnor UO_644 (O_644,N_14516,N_10414);
nand UO_645 (O_645,N_12928,N_11019);
nand UO_646 (O_646,N_11545,N_14067);
or UO_647 (O_647,N_12573,N_13796);
or UO_648 (O_648,N_10832,N_10499);
and UO_649 (O_649,N_12228,N_10122);
or UO_650 (O_650,N_10097,N_10138);
or UO_651 (O_651,N_13669,N_10002);
nor UO_652 (O_652,N_10939,N_12810);
or UO_653 (O_653,N_10932,N_10293);
nand UO_654 (O_654,N_11453,N_13117);
nor UO_655 (O_655,N_14072,N_10930);
nand UO_656 (O_656,N_10530,N_11321);
or UO_657 (O_657,N_14145,N_11912);
nand UO_658 (O_658,N_11263,N_14330);
nand UO_659 (O_659,N_12504,N_14858);
nand UO_660 (O_660,N_13531,N_13984);
and UO_661 (O_661,N_12052,N_13511);
or UO_662 (O_662,N_14474,N_12813);
nand UO_663 (O_663,N_14010,N_11816);
nand UO_664 (O_664,N_11610,N_12532);
or UO_665 (O_665,N_12208,N_14522);
nand UO_666 (O_666,N_14454,N_14460);
nand UO_667 (O_667,N_14210,N_10420);
nand UO_668 (O_668,N_13622,N_14440);
nand UO_669 (O_669,N_10026,N_13497);
and UO_670 (O_670,N_12488,N_11886);
nand UO_671 (O_671,N_12932,N_13788);
nand UO_672 (O_672,N_13625,N_10397);
nand UO_673 (O_673,N_13443,N_13395);
nor UO_674 (O_674,N_11236,N_10208);
nor UO_675 (O_675,N_11536,N_14037);
and UO_676 (O_676,N_10411,N_12684);
and UO_677 (O_677,N_13729,N_13963);
nor UO_678 (O_678,N_14942,N_13213);
nor UO_679 (O_679,N_14656,N_10128);
and UO_680 (O_680,N_11205,N_13327);
nor UO_681 (O_681,N_11822,N_10265);
and UO_682 (O_682,N_14270,N_13224);
nand UO_683 (O_683,N_14585,N_11027);
and UO_684 (O_684,N_13243,N_10522);
or UO_685 (O_685,N_10309,N_14953);
nor UO_686 (O_686,N_10974,N_14838);
nor UO_687 (O_687,N_13199,N_12574);
and UO_688 (O_688,N_11866,N_13979);
or UO_689 (O_689,N_14568,N_12517);
nand UO_690 (O_690,N_13626,N_11896);
and UO_691 (O_691,N_12682,N_13171);
or UO_692 (O_692,N_10020,N_11050);
or UO_693 (O_693,N_14588,N_14506);
and UO_694 (O_694,N_10942,N_13110);
nor UO_695 (O_695,N_11127,N_10480);
and UO_696 (O_696,N_14308,N_14155);
or UO_697 (O_697,N_10351,N_14959);
nor UO_698 (O_698,N_13914,N_10217);
nand UO_699 (O_699,N_14920,N_10056);
and UO_700 (O_700,N_10405,N_13762);
xnor UO_701 (O_701,N_14082,N_10178);
nand UO_702 (O_702,N_10516,N_14347);
nand UO_703 (O_703,N_10779,N_12739);
nor UO_704 (O_704,N_14596,N_13819);
or UO_705 (O_705,N_13123,N_10290);
nor UO_706 (O_706,N_12869,N_12991);
and UO_707 (O_707,N_12632,N_12531);
nor UO_708 (O_708,N_12149,N_12192);
or UO_709 (O_709,N_14290,N_13280);
and UO_710 (O_710,N_10213,N_12748);
nand UO_711 (O_711,N_10363,N_10000);
or UO_712 (O_712,N_13637,N_10815);
nor UO_713 (O_713,N_10863,N_11105);
and UO_714 (O_714,N_14180,N_13640);
or UO_715 (O_715,N_13385,N_10563);
or UO_716 (O_716,N_11175,N_10288);
and UO_717 (O_717,N_10033,N_10960);
nor UO_718 (O_718,N_13013,N_11835);
nand UO_719 (O_719,N_11071,N_12172);
nand UO_720 (O_720,N_12616,N_11139);
nor UO_721 (O_721,N_12509,N_11765);
and UO_722 (O_722,N_14409,N_11290);
nand UO_723 (O_723,N_14352,N_12068);
and UO_724 (O_724,N_11382,N_13659);
and UO_725 (O_725,N_12527,N_10451);
or UO_726 (O_726,N_13200,N_10600);
and UO_727 (O_727,N_13097,N_12250);
nor UO_728 (O_728,N_12167,N_12873);
or UO_729 (O_729,N_11386,N_12021);
or UO_730 (O_730,N_14592,N_12762);
or UO_731 (O_731,N_11314,N_10349);
nor UO_732 (O_732,N_14427,N_11012);
nor UO_733 (O_733,N_10750,N_10014);
or UO_734 (O_734,N_14276,N_12421);
and UO_735 (O_735,N_14724,N_11932);
xor UO_736 (O_736,N_12457,N_14731);
and UO_737 (O_737,N_11750,N_14946);
and UO_738 (O_738,N_12277,N_11830);
and UO_739 (O_739,N_14357,N_13867);
and UO_740 (O_740,N_12217,N_13252);
nor UO_741 (O_741,N_12940,N_12373);
and UO_742 (O_742,N_13122,N_12139);
nand UO_743 (O_743,N_14922,N_14975);
nand UO_744 (O_744,N_10153,N_14595);
or UO_745 (O_745,N_12055,N_12771);
nand UO_746 (O_746,N_13040,N_12393);
nand UO_747 (O_747,N_13396,N_12623);
nand UO_748 (O_748,N_14730,N_14167);
or UO_749 (O_749,N_12060,N_11871);
nand UO_750 (O_750,N_14174,N_14396);
nor UO_751 (O_751,N_11258,N_12575);
or UO_752 (O_752,N_10847,N_10460);
and UO_753 (O_753,N_11267,N_12200);
or UO_754 (O_754,N_10456,N_14221);
nor UO_755 (O_755,N_11857,N_12295);
nand UO_756 (O_756,N_14649,N_14836);
nand UO_757 (O_757,N_11586,N_11813);
nand UO_758 (O_758,N_12951,N_12029);
nand UO_759 (O_759,N_12751,N_10667);
or UO_760 (O_760,N_14537,N_11344);
and UO_761 (O_761,N_13631,N_10711);
or UO_762 (O_762,N_11756,N_13590);
or UO_763 (O_763,N_12450,N_11859);
or UO_764 (O_764,N_13315,N_10319);
and UO_765 (O_765,N_10895,N_10023);
and UO_766 (O_766,N_12665,N_12342);
and UO_767 (O_767,N_13923,N_13756);
nand UO_768 (O_768,N_14249,N_10114);
and UO_769 (O_769,N_14809,N_12769);
nor UO_770 (O_770,N_13190,N_12620);
nor UO_771 (O_771,N_12298,N_14706);
nor UO_772 (O_772,N_14102,N_10272);
and UO_773 (O_773,N_13397,N_11483);
and UO_774 (O_774,N_14277,N_13539);
nand UO_775 (O_775,N_14648,N_11563);
nand UO_776 (O_776,N_11218,N_10254);
or UO_777 (O_777,N_11281,N_13836);
nand UO_778 (O_778,N_10462,N_14345);
nand UO_779 (O_779,N_10838,N_10693);
nand UO_780 (O_780,N_11524,N_12434);
or UO_781 (O_781,N_13812,N_11277);
nand UO_782 (O_782,N_13059,N_13841);
or UO_783 (O_783,N_13394,N_10828);
and UO_784 (O_784,N_12805,N_12840);
and UO_785 (O_785,N_10703,N_10823);
nand UO_786 (O_786,N_14619,N_10259);
and UO_787 (O_787,N_12768,N_10166);
nand UO_788 (O_788,N_12464,N_13583);
and UO_789 (O_789,N_13639,N_13585);
nor UO_790 (O_790,N_13865,N_12673);
nor UO_791 (O_791,N_11398,N_11025);
xnor UO_792 (O_792,N_11134,N_10084);
nor UO_793 (O_793,N_14464,N_11247);
or UO_794 (O_794,N_11566,N_11649);
or UO_795 (O_795,N_10567,N_10904);
or UO_796 (O_796,N_11318,N_11847);
and UO_797 (O_797,N_10743,N_12972);
and UO_798 (O_798,N_11117,N_12209);
and UO_799 (O_799,N_13581,N_10300);
nor UO_800 (O_800,N_10990,N_10168);
and UO_801 (O_801,N_11180,N_12290);
nor UO_802 (O_802,N_10673,N_13782);
nand UO_803 (O_803,N_10214,N_10461);
nand UO_804 (O_804,N_11749,N_10827);
and UO_805 (O_805,N_10964,N_14718);
nor UO_806 (O_806,N_14489,N_14853);
or UO_807 (O_807,N_14197,N_13601);
nand UO_808 (O_808,N_14192,N_11103);
or UO_809 (O_809,N_11679,N_12100);
nor UO_810 (O_810,N_13042,N_14219);
nand UO_811 (O_811,N_12259,N_11055);
and UO_812 (O_812,N_14518,N_10805);
nor UO_813 (O_813,N_12720,N_14432);
or UO_814 (O_814,N_12614,N_14311);
nor UO_815 (O_815,N_14285,N_11494);
nand UO_816 (O_816,N_13298,N_13103);
nand UO_817 (O_817,N_13433,N_13671);
and UO_818 (O_818,N_11587,N_14916);
or UO_819 (O_819,N_10088,N_12777);
nor UO_820 (O_820,N_14917,N_13462);
and UO_821 (O_821,N_14195,N_11667);
nor UO_822 (O_822,N_10134,N_14282);
nor UO_823 (O_823,N_14758,N_12700);
nand UO_824 (O_824,N_12235,N_12197);
or UO_825 (O_825,N_14835,N_10044);
nor UO_826 (O_826,N_12401,N_14186);
or UO_827 (O_827,N_13483,N_13334);
or UO_828 (O_828,N_14178,N_12716);
or UO_829 (O_829,N_14272,N_10145);
or UO_830 (O_830,N_14196,N_10685);
or UO_831 (O_831,N_14362,N_11137);
and UO_832 (O_832,N_12109,N_11445);
nand UO_833 (O_833,N_14562,N_13007);
and UO_834 (O_834,N_13389,N_10812);
nand UO_835 (O_835,N_13952,N_14839);
nand UO_836 (O_836,N_12561,N_11337);
and UO_837 (O_837,N_14634,N_11564);
nor UO_838 (O_838,N_12899,N_10106);
nor UO_839 (O_839,N_10970,N_12663);
and UO_840 (O_840,N_12078,N_14320);
or UO_841 (O_841,N_10800,N_13916);
nor UO_842 (O_842,N_10789,N_13617);
and UO_843 (O_843,N_10661,N_10956);
or UO_844 (O_844,N_13724,N_11460);
or UO_845 (O_845,N_12496,N_11387);
or UO_846 (O_846,N_14501,N_11419);
and UO_847 (O_847,N_12123,N_14646);
nor UO_848 (O_848,N_10170,N_12866);
nor UO_849 (O_849,N_13233,N_12157);
and UO_850 (O_850,N_10938,N_14662);
or UO_851 (O_851,N_10755,N_12983);
and UO_852 (O_852,N_12566,N_13852);
and UO_853 (O_853,N_13052,N_12292);
nand UO_854 (O_854,N_10808,N_11743);
nor UO_855 (O_855,N_14230,N_10880);
nor UO_856 (O_856,N_14350,N_14324);
nor UO_857 (O_857,N_10773,N_10949);
nor UO_858 (O_858,N_13664,N_12994);
nor UO_859 (O_859,N_13689,N_12023);
and UO_860 (O_860,N_11538,N_11708);
nor UO_861 (O_861,N_14083,N_10598);
nor UO_862 (O_862,N_10296,N_12212);
nand UO_863 (O_863,N_11320,N_13921);
and UO_864 (O_864,N_13540,N_12440);
or UO_865 (O_865,N_10270,N_13744);
nand UO_866 (O_866,N_13442,N_11391);
nand UO_867 (O_867,N_12500,N_11780);
nand UO_868 (O_868,N_10109,N_10915);
and UO_869 (O_869,N_14997,N_13314);
and UO_870 (O_870,N_12129,N_11962);
nand UO_871 (O_871,N_11474,N_12698);
nand UO_872 (O_872,N_14482,N_13816);
nor UO_873 (O_873,N_14264,N_10336);
nor UO_874 (O_874,N_12145,N_13342);
nand UO_875 (O_875,N_10679,N_12920);
nand UO_876 (O_876,N_10536,N_12048);
or UO_877 (O_877,N_12947,N_11487);
nand UO_878 (O_878,N_11104,N_13400);
nor UO_879 (O_879,N_14905,N_10104);
nand UO_880 (O_880,N_13492,N_13047);
nand UO_881 (O_881,N_12930,N_14297);
nor UO_882 (O_882,N_14644,N_10677);
nor UO_883 (O_883,N_14310,N_11230);
and UO_884 (O_884,N_11839,N_11086);
or UO_885 (O_885,N_12807,N_10558);
or UO_886 (O_886,N_14825,N_10240);
and UO_887 (O_887,N_13289,N_12012);
or UO_888 (O_888,N_12913,N_10725);
nand UO_889 (O_889,N_11430,N_12847);
nor UO_890 (O_890,N_11530,N_14663);
nand UO_891 (O_891,N_13313,N_12979);
nor UO_892 (O_892,N_11152,N_13566);
nand UO_893 (O_893,N_12383,N_10352);
nor UO_894 (O_894,N_12442,N_14329);
or UO_895 (O_895,N_12476,N_11827);
nand UO_896 (O_896,N_11862,N_14700);
nand UO_897 (O_897,N_12818,N_10374);
and UO_898 (O_898,N_14660,N_12775);
and UO_899 (O_899,N_13305,N_10928);
nor UO_900 (O_900,N_13464,N_14719);
nand UO_901 (O_901,N_12604,N_10062);
nand UO_902 (O_902,N_11464,N_12062);
or UO_903 (O_903,N_14258,N_12127);
nand UO_904 (O_904,N_11878,N_10754);
nand UO_905 (O_905,N_12822,N_13114);
and UO_906 (O_906,N_14632,N_11319);
xor UO_907 (O_907,N_12914,N_14996);
and UO_908 (O_908,N_11596,N_12271);
or UO_909 (O_909,N_11178,N_13245);
nor UO_910 (O_910,N_10787,N_10952);
and UO_911 (O_911,N_14571,N_12588);
nand UO_912 (O_912,N_10230,N_14767);
or UO_913 (O_913,N_12072,N_12207);
and UO_914 (O_914,N_10407,N_12832);
nand UO_915 (O_915,N_11064,N_10440);
or UO_916 (O_916,N_13759,N_13096);
xor UO_917 (O_917,N_10482,N_14376);
nand UO_918 (O_918,N_12570,N_11528);
nand UO_919 (O_919,N_10816,N_11274);
and UO_920 (O_920,N_11168,N_14242);
nand UO_921 (O_921,N_12013,N_14654);
nand UO_922 (O_922,N_11128,N_12779);
or UO_923 (O_923,N_11629,N_13002);
and UO_924 (O_924,N_12018,N_12061);
or UO_925 (O_925,N_13832,N_12901);
and UO_926 (O_926,N_11604,N_13958);
and UO_927 (O_927,N_10236,N_13814);
or UO_928 (O_928,N_13882,N_11355);
nor UO_929 (O_929,N_10881,N_11736);
nand UO_930 (O_930,N_11573,N_14146);
nand UO_931 (O_931,N_11716,N_10129);
nor UO_932 (O_932,N_13094,N_14215);
and UO_933 (O_933,N_10489,N_12778);
or UO_934 (O_934,N_10080,N_13153);
nand UO_935 (O_935,N_12314,N_14012);
nor UO_936 (O_936,N_11286,N_13235);
or UO_937 (O_937,N_14545,N_10736);
xor UO_938 (O_938,N_12293,N_13265);
and UO_939 (O_939,N_12396,N_14211);
and UO_940 (O_940,N_13894,N_12199);
and UO_941 (O_941,N_10164,N_13681);
and UO_942 (O_942,N_10729,N_14176);
nand UO_943 (O_943,N_12710,N_11527);
or UO_944 (O_944,N_10393,N_11029);
and UO_945 (O_945,N_14226,N_10361);
nand UO_946 (O_946,N_14974,N_14090);
or UO_947 (O_947,N_10723,N_11740);
nand UO_948 (O_948,N_14556,N_14385);
nand UO_949 (O_949,N_14672,N_10231);
nor UO_950 (O_950,N_11298,N_14096);
and UO_951 (O_951,N_10235,N_12382);
and UO_952 (O_952,N_13065,N_11157);
or UO_953 (O_953,N_11498,N_10903);
nand UO_954 (O_954,N_11024,N_11221);
nand UO_955 (O_955,N_14950,N_14325);
nand UO_956 (O_956,N_14097,N_14605);
nand UO_957 (O_957,N_12352,N_14153);
nor UO_958 (O_958,N_12902,N_10640);
and UO_959 (O_959,N_10545,N_13697);
nor UO_960 (O_960,N_10297,N_14101);
or UO_961 (O_961,N_12263,N_13964);
nand UO_962 (O_962,N_12067,N_14000);
nor UO_963 (O_963,N_13662,N_13113);
and UO_964 (O_964,N_13295,N_13183);
nand UO_965 (O_965,N_11917,N_11676);
and UO_966 (O_966,N_14740,N_12437);
or UO_967 (O_967,N_10514,N_11733);
nand UO_968 (O_968,N_10306,N_14587);
and UO_969 (O_969,N_13802,N_13644);
nand UO_970 (O_970,N_12882,N_13754);
nor UO_971 (O_971,N_12525,N_10523);
or UO_972 (O_972,N_12732,N_10506);
nor UO_973 (O_973,N_11627,N_13582);
nand UO_974 (O_974,N_11378,N_14315);
and UO_975 (O_975,N_13904,N_10984);
nor UO_976 (O_976,N_11358,N_13131);
nand UO_977 (O_977,N_10078,N_12728);
nor UO_978 (O_978,N_13850,N_14020);
nand UO_979 (O_979,N_12656,N_14990);
or UO_980 (O_980,N_14686,N_10840);
and UO_981 (O_981,N_14316,N_14885);
and UO_982 (O_982,N_14848,N_13323);
nor UO_983 (O_983,N_14551,N_13673);
nor UO_984 (O_984,N_12957,N_13698);
nand UO_985 (O_985,N_13164,N_13241);
nor UO_986 (O_986,N_10951,N_11447);
nand UO_987 (O_987,N_11974,N_14681);
nand UO_988 (O_988,N_14527,N_14914);
or UO_989 (O_989,N_10888,N_10820);
or UO_990 (O_990,N_11181,N_10330);
and UO_991 (O_991,N_12403,N_13343);
xor UO_992 (O_992,N_14967,N_12676);
and UO_993 (O_993,N_14438,N_12017);
nand UO_994 (O_994,N_14085,N_14629);
and UO_995 (O_995,N_14236,N_14336);
nand UO_996 (O_996,N_12568,N_13185);
nand UO_997 (O_997,N_10612,N_14668);
and UO_998 (O_998,N_13755,N_14003);
and UO_999 (O_999,N_14470,N_10141);
nor UO_1000 (O_1000,N_10791,N_11823);
or UO_1001 (O_1001,N_11580,N_10205);
or UO_1002 (O_1002,N_11070,N_12662);
and UO_1003 (O_1003,N_14851,N_11162);
nor UO_1004 (O_1004,N_13476,N_13432);
nor UO_1005 (O_1005,N_12670,N_13857);
or UO_1006 (O_1006,N_14621,N_13668);
nand UO_1007 (O_1007,N_11956,N_13128);
nor UO_1008 (O_1008,N_10322,N_13774);
or UO_1009 (O_1009,N_10412,N_10163);
and UO_1010 (O_1010,N_14499,N_12378);
and UO_1011 (O_1011,N_10016,N_11609);
nor UO_1012 (O_1012,N_12788,N_13651);
nand UO_1013 (O_1013,N_10085,N_12224);
or UO_1014 (O_1014,N_14268,N_10535);
and UO_1015 (O_1015,N_11155,N_11179);
or UO_1016 (O_1016,N_13856,N_13261);
nand UO_1017 (O_1017,N_11876,N_14928);
nor UO_1018 (O_1018,N_10633,N_12037);
nand UO_1019 (O_1019,N_12741,N_14371);
nand UO_1020 (O_1020,N_13438,N_11389);
and UO_1021 (O_1021,N_10962,N_14100);
nand UO_1022 (O_1022,N_11943,N_13833);
nor UO_1023 (O_1023,N_10588,N_11612);
nand UO_1024 (O_1024,N_12305,N_11192);
nand UO_1025 (O_1025,N_12757,N_13201);
and UO_1026 (O_1026,N_10654,N_10307);
and UO_1027 (O_1027,N_11789,N_11655);
nand UO_1028 (O_1028,N_11907,N_13390);
and UO_1029 (O_1029,N_12011,N_14620);
or UO_1030 (O_1030,N_13416,N_11653);
and UO_1031 (O_1031,N_12108,N_11008);
or UO_1032 (O_1032,N_14569,N_10553);
or UO_1033 (O_1033,N_10466,N_14679);
or UO_1034 (O_1034,N_10312,N_14053);
and UO_1035 (O_1035,N_11457,N_11473);
or UO_1036 (O_1036,N_10759,N_12697);
and UO_1037 (O_1037,N_11895,N_12120);
and UO_1038 (O_1038,N_10571,N_14300);
nor UO_1039 (O_1039,N_11058,N_14613);
nor UO_1040 (O_1040,N_11870,N_14267);
nand UO_1041 (O_1041,N_12721,N_11910);
and UO_1042 (O_1042,N_11449,N_13500);
and UO_1043 (O_1043,N_10613,N_11224);
nand UO_1044 (O_1044,N_13598,N_14025);
or UO_1045 (O_1045,N_12024,N_13924);
and UO_1046 (O_1046,N_14333,N_10454);
and UO_1047 (O_1047,N_10150,N_13623);
and UO_1048 (O_1048,N_13512,N_12695);
and UO_1049 (O_1049,N_13027,N_14377);
nor UO_1050 (O_1050,N_14036,N_12269);
nand UO_1051 (O_1051,N_12001,N_11978);
nor UO_1052 (O_1052,N_14407,N_13554);
nor UO_1053 (O_1053,N_13676,N_11015);
or UO_1054 (O_1054,N_13149,N_13959);
and UO_1055 (O_1055,N_14845,N_10653);
or UO_1056 (O_1056,N_13071,N_12170);
nor UO_1057 (O_1057,N_12143,N_10069);
or UO_1058 (O_1058,N_10958,N_10359);
or UO_1059 (O_1059,N_13928,N_14653);
nor UO_1060 (O_1060,N_12386,N_14485);
or UO_1061 (O_1061,N_11567,N_10705);
or UO_1062 (O_1062,N_14794,N_10849);
and UO_1063 (O_1063,N_12459,N_13402);
nand UO_1064 (O_1064,N_13546,N_14607);
and UO_1065 (O_1065,N_11774,N_12307);
nor UO_1066 (O_1066,N_12917,N_10993);
nand UO_1067 (O_1067,N_13791,N_10194);
or UO_1068 (O_1068,N_14303,N_11686);
or UO_1069 (O_1069,N_11216,N_14449);
nor UO_1070 (O_1070,N_14507,N_10198);
or UO_1071 (O_1071,N_14608,N_10561);
xnor UO_1072 (O_1072,N_12137,N_10496);
or UO_1073 (O_1073,N_10580,N_14842);
and UO_1074 (O_1074,N_10445,N_13479);
nor UO_1075 (O_1075,N_10261,N_14565);
nand UO_1076 (O_1076,N_14252,N_13555);
or UO_1077 (O_1077,N_10758,N_11421);
or UO_1078 (O_1078,N_13018,N_10038);
and UO_1079 (O_1079,N_11346,N_13478);
nor UO_1080 (O_1080,N_11122,N_14883);
nand UO_1081 (O_1081,N_12064,N_11207);
and UO_1082 (O_1082,N_13475,N_10468);
xnor UO_1083 (O_1083,N_11658,N_14643);
nand UO_1084 (O_1084,N_12146,N_12322);
or UO_1085 (O_1085,N_12555,N_14213);
nand UO_1086 (O_1086,N_13001,N_13868);
nand UO_1087 (O_1087,N_13975,N_10350);
nor UO_1088 (O_1088,N_11289,N_12627);
nand UO_1089 (O_1089,N_13685,N_14122);
and UO_1090 (O_1090,N_10124,N_12879);
and UO_1091 (O_1091,N_13538,N_11721);
nand UO_1092 (O_1092,N_14535,N_14616);
nor UO_1093 (O_1093,N_13530,N_14816);
or UO_1094 (O_1094,N_14623,N_10339);
and UO_1095 (O_1095,N_14941,N_13621);
and UO_1096 (O_1096,N_10643,N_12034);
nand UO_1097 (O_1097,N_13477,N_13049);
and UO_1098 (O_1098,N_10572,N_10794);
and UO_1099 (O_1099,N_11388,N_12094);
nor UO_1100 (O_1100,N_11969,N_12283);
nand UO_1101 (O_1101,N_12040,N_12409);
or UO_1102 (O_1102,N_10365,N_12513);
nor UO_1103 (O_1103,N_10073,N_12725);
nor UO_1104 (O_1104,N_10429,N_11704);
nor UO_1105 (O_1105,N_13466,N_11303);
or UO_1106 (O_1106,N_13087,N_13360);
nor UO_1107 (O_1107,N_12097,N_14584);
nand UO_1108 (O_1108,N_12178,N_13033);
nor UO_1109 (O_1109,N_10943,N_14819);
xor UO_1110 (O_1110,N_14484,N_10271);
and UO_1111 (O_1111,N_13628,N_10228);
or UO_1112 (O_1112,N_13048,N_13752);
nand UO_1113 (O_1113,N_14727,N_12955);
or UO_1114 (O_1114,N_14677,N_14583);
nand UO_1115 (O_1115,N_13706,N_13973);
and UO_1116 (O_1116,N_12624,N_12787);
or UO_1117 (O_1117,N_14940,N_13004);
nand UO_1118 (O_1118,N_12326,N_14425);
and UO_1119 (O_1119,N_11858,N_13430);
nor UO_1120 (O_1120,N_11824,N_13932);
nand UO_1121 (O_1121,N_11766,N_14417);
and UO_1122 (O_1122,N_10829,N_13277);
nor UO_1123 (O_1123,N_13111,N_11994);
nor UO_1124 (O_1124,N_11408,N_13152);
and UO_1125 (O_1125,N_12446,N_12159);
or UO_1126 (O_1126,N_14398,N_13125);
nor UO_1127 (O_1127,N_10072,N_10738);
or UO_1128 (O_1128,N_14319,N_10512);
or UO_1129 (O_1129,N_11272,N_12781);
or UO_1130 (O_1130,N_12520,N_13439);
nand UO_1131 (O_1131,N_10893,N_13257);
or UO_1132 (O_1132,N_12089,N_11472);
and UO_1133 (O_1133,N_13444,N_14704);
and UO_1134 (O_1134,N_11725,N_12033);
nand UO_1135 (O_1135,N_14821,N_14743);
or UO_1136 (O_1136,N_11642,N_11772);
and UO_1137 (O_1137,N_12693,N_10332);
or UO_1138 (O_1138,N_14389,N_10860);
and UO_1139 (O_1139,N_10748,N_13457);
or UO_1140 (O_1140,N_13827,N_10256);
nor UO_1141 (O_1141,N_12861,N_13260);
or UO_1142 (O_1142,N_11958,N_14918);
and UO_1143 (O_1143,N_10959,N_11295);
nand UO_1144 (O_1144,N_13270,N_11413);
nand UO_1145 (O_1145,N_10061,N_10282);
or UO_1146 (O_1146,N_10457,N_14765);
nor UO_1147 (O_1147,N_11261,N_12582);
or UO_1148 (O_1148,N_12291,N_14231);
nor UO_1149 (O_1149,N_12121,N_10621);
nand UO_1150 (O_1150,N_11864,N_12242);
and UO_1151 (O_1151,N_10310,N_12664);
or UO_1152 (O_1152,N_13000,N_13104);
or UO_1153 (O_1153,N_12050,N_10123);
and UO_1154 (O_1154,N_14659,N_10394);
or UO_1155 (O_1155,N_11232,N_13388);
and UO_1156 (O_1156,N_12986,N_11631);
or UO_1157 (O_1157,N_10481,N_11685);
and UO_1158 (O_1158,N_12231,N_10160);
nand UO_1159 (O_1159,N_11731,N_12543);
nand UO_1160 (O_1160,N_11488,N_11147);
nand UO_1161 (O_1161,N_12354,N_12056);
and UO_1162 (O_1162,N_13926,N_14307);
and UO_1163 (O_1163,N_11705,N_13371);
or UO_1164 (O_1164,N_14321,N_13568);
nand UO_1165 (O_1165,N_13761,N_11865);
nand UO_1166 (O_1166,N_10985,N_10722);
nand UO_1167 (O_1167,N_10782,N_10632);
or UO_1168 (O_1168,N_10687,N_12294);
or UO_1169 (O_1169,N_14043,N_12118);
and UO_1170 (O_1170,N_13344,N_10111);
or UO_1171 (O_1171,N_14355,N_12470);
and UO_1172 (O_1172,N_14034,N_12921);
and UO_1173 (O_1173,N_11980,N_14913);
and UO_1174 (O_1174,N_10935,N_12880);
nor UO_1175 (O_1175,N_11243,N_12657);
or UO_1176 (O_1176,N_10427,N_11291);
nand UO_1177 (O_1177,N_11739,N_10500);
nand UO_1178 (O_1178,N_12467,N_14760);
and UO_1179 (O_1179,N_10855,N_14162);
nand UO_1180 (O_1180,N_14443,N_10799);
or UO_1181 (O_1181,N_13560,N_12468);
nand UO_1182 (O_1182,N_11074,N_11920);
nor UO_1183 (O_1183,N_10284,N_12002);
and UO_1184 (O_1184,N_11432,N_12163);
nand UO_1185 (O_1185,N_10784,N_10136);
nand UO_1186 (O_1186,N_13369,N_12841);
nor UO_1187 (O_1187,N_10646,N_14713);
nor UO_1188 (O_1188,N_12562,N_10484);
nand UO_1189 (O_1189,N_11955,N_12845);
nor UO_1190 (O_1190,N_14206,N_13362);
and UO_1191 (O_1191,N_13771,N_11083);
or UO_1192 (O_1192,N_11729,N_12452);
nor UO_1193 (O_1193,N_13205,N_11461);
and UO_1194 (O_1194,N_11130,N_13745);
and UO_1195 (O_1195,N_14631,N_11518);
nor UO_1196 (O_1196,N_11496,N_11693);
nor UO_1197 (O_1197,N_13045,N_11435);
nor UO_1198 (O_1198,N_12878,N_13961);
or UO_1199 (O_1199,N_13881,N_11073);
nand UO_1200 (O_1200,N_13246,N_14988);
and UO_1201 (O_1201,N_11266,N_12954);
and UO_1202 (O_1202,N_10091,N_13521);
nand UO_1203 (O_1203,N_11977,N_14240);
nor UO_1204 (O_1204,N_12038,N_14589);
nor UO_1205 (O_1205,N_13860,N_13182);
and UO_1206 (O_1206,N_14088,N_11561);
nor UO_1207 (O_1207,N_10624,N_12941);
nor UO_1208 (O_1208,N_12239,N_13297);
and UO_1209 (O_1209,N_12950,N_12035);
or UO_1210 (O_1210,N_11144,N_12599);
or UO_1211 (O_1211,N_13988,N_11384);
or UO_1212 (O_1212,N_14452,N_13562);
and UO_1213 (O_1213,N_13594,N_10083);
and UO_1214 (O_1214,N_14486,N_12828);
xor UO_1215 (O_1215,N_10924,N_11761);
or UO_1216 (O_1216,N_14260,N_11482);
or UO_1217 (O_1217,N_13842,N_12414);
nand UO_1218 (O_1218,N_11428,N_11957);
and UO_1219 (O_1219,N_12155,N_11177);
nor UO_1220 (O_1220,N_11577,N_14888);
and UO_1221 (O_1221,N_12447,N_11371);
or UO_1222 (O_1222,N_11760,N_12417);
and UO_1223 (O_1223,N_14156,N_14128);
or UO_1224 (O_1224,N_12816,N_13800);
and UO_1225 (O_1225,N_12394,N_13714);
nand UO_1226 (O_1226,N_13274,N_13737);
and UO_1227 (O_1227,N_10251,N_12216);
nand UO_1228 (O_1228,N_14323,N_13140);
nor UO_1229 (O_1229,N_11793,N_14497);
or UO_1230 (O_1230,N_13804,N_10871);
and UO_1231 (O_1231,N_13597,N_13324);
and UO_1232 (O_1232,N_11788,N_14769);
or UO_1233 (O_1233,N_14105,N_10788);
or UO_1234 (O_1234,N_11723,N_13677);
or UO_1235 (O_1235,N_11673,N_12931);
nand UO_1236 (O_1236,N_12827,N_11051);
or UO_1237 (O_1237,N_12369,N_10207);
nor UO_1238 (O_1238,N_14982,N_13820);
xor UO_1239 (O_1239,N_13897,N_13193);
and UO_1240 (O_1240,N_13749,N_14717);
or UO_1241 (O_1241,N_10552,N_13172);
or UO_1242 (O_1242,N_12605,N_11507);
and UO_1243 (O_1243,N_11552,N_12912);
nor UO_1244 (O_1244,N_14638,N_14218);
nor UO_1245 (O_1245,N_14216,N_13014);
and UO_1246 (O_1246,N_10543,N_11145);
nor UO_1247 (O_1247,N_14295,N_14117);
and UO_1248 (O_1248,N_11349,N_14673);
nand UO_1249 (O_1249,N_14453,N_13124);
or UO_1250 (O_1250,N_13053,N_14339);
or UO_1251 (O_1251,N_13130,N_13482);
nand UO_1252 (O_1252,N_11161,N_13044);
nand UO_1253 (O_1253,N_11328,N_13005);
nor UO_1254 (O_1254,N_12886,N_10464);
and UO_1255 (O_1255,N_14658,N_12243);
or UO_1256 (O_1256,N_14908,N_10186);
or UO_1257 (O_1257,N_10697,N_13835);
nand UO_1258 (O_1258,N_14861,N_13913);
and UO_1259 (O_1259,N_11752,N_14478);
nor UO_1260 (O_1260,N_11285,N_10557);
and UO_1261 (O_1261,N_14799,N_12622);
nor UO_1262 (O_1262,N_12348,N_10209);
and UO_1263 (O_1263,N_10846,N_13239);
or UO_1264 (O_1264,N_12548,N_12563);
nand UO_1265 (O_1265,N_10638,N_12556);
and UO_1266 (O_1266,N_11227,N_12526);
and UO_1267 (O_1267,N_10067,N_14635);
or UO_1268 (O_1268,N_11656,N_11570);
and UO_1269 (O_1269,N_13826,N_14705);
or UO_1270 (O_1270,N_14870,N_10657);
and UO_1271 (O_1271,N_13572,N_14394);
or UO_1272 (O_1272,N_12529,N_12377);
or UO_1273 (O_1273,N_13872,N_10248);
nor UO_1274 (O_1274,N_13848,N_10701);
or UO_1275 (O_1275,N_14373,N_12107);
and UO_1276 (O_1276,N_12130,N_10950);
nor UO_1277 (O_1277,N_14707,N_11032);
nand UO_1278 (O_1278,N_13575,N_14812);
nor UO_1279 (O_1279,N_10116,N_10304);
and UO_1280 (O_1280,N_12685,N_13498);
xor UO_1281 (O_1281,N_11252,N_10626);
nand UO_1282 (O_1282,N_10762,N_10641);
nor UO_1283 (O_1283,N_11746,N_14779);
or UO_1284 (O_1284,N_12974,N_12195);
nand UO_1285 (O_1285,N_12851,N_11717);
nand UO_1286 (O_1286,N_11639,N_11079);
or UO_1287 (O_1287,N_10321,N_14871);
nand UO_1288 (O_1288,N_13039,N_11154);
nor UO_1289 (O_1289,N_12279,N_11623);
or UO_1290 (O_1290,N_11129,N_13741);
nand UO_1291 (O_1291,N_12964,N_12892);
nor UO_1292 (O_1292,N_10151,N_11067);
or UO_1293 (O_1293,N_14039,N_10948);
nor UO_1294 (O_1294,N_13649,N_12923);
nor UO_1295 (O_1295,N_11519,N_10739);
nand UO_1296 (O_1296,N_13822,N_11727);
xnor UO_1297 (O_1297,N_12533,N_14114);
and UO_1298 (O_1298,N_13267,N_14747);
and UO_1299 (O_1299,N_10008,N_13773);
and UO_1300 (O_1300,N_10662,N_14862);
nand UO_1301 (O_1301,N_11362,N_11925);
nor UO_1302 (O_1302,N_10848,N_10781);
nor UO_1303 (O_1303,N_10796,N_11734);
or UO_1304 (O_1304,N_10439,N_11529);
nor UO_1305 (O_1305,N_11292,N_13168);
and UO_1306 (O_1306,N_11377,N_13157);
nand UO_1307 (O_1307,N_12185,N_14756);
or UO_1308 (O_1308,N_11276,N_13778);
or UO_1309 (O_1309,N_11400,N_14170);
nand UO_1310 (O_1310,N_10810,N_13723);
and UO_1311 (O_1311,N_10547,N_11217);
and UO_1312 (O_1312,N_12784,N_14133);
nand UO_1313 (O_1313,N_14531,N_12288);
nand UO_1314 (O_1314,N_14009,N_13898);
and UO_1315 (O_1315,N_14581,N_11312);
nand UO_1316 (O_1316,N_11533,N_13602);
xnor UO_1317 (O_1317,N_13450,N_12475);
nand UO_1318 (O_1318,N_11581,N_12846);
xnor UO_1319 (O_1319,N_12430,N_12077);
and UO_1320 (O_1320,N_11650,N_13683);
and UO_1321 (O_1321,N_11613,N_13927);
and UO_1322 (O_1322,N_12222,N_12990);
or UO_1323 (O_1323,N_10521,N_11754);
and UO_1324 (O_1324,N_12350,N_12193);
and UO_1325 (O_1325,N_11331,N_13361);
or UO_1326 (O_1326,N_12204,N_14752);
nand UO_1327 (O_1327,N_12884,N_14254);
nor UO_1328 (O_1328,N_11476,N_13355);
and UO_1329 (O_1329,N_13516,N_14135);
nand UO_1330 (O_1330,N_12843,N_13228);
or UO_1331 (O_1331,N_12753,N_14833);
and UO_1332 (O_1332,N_11091,N_10131);
or UO_1333 (O_1333,N_10196,N_11753);
nand UO_1334 (O_1334,N_13910,N_11602);
nand UO_1335 (O_1335,N_12877,N_12937);
or UO_1336 (O_1336,N_13347,N_13829);
and UO_1337 (O_1337,N_14032,N_14965);
nor UO_1338 (O_1338,N_12681,N_10247);
or UO_1339 (O_1339,N_11270,N_11904);
and UO_1340 (O_1340,N_11353,N_10916);
nand UO_1341 (O_1341,N_14647,N_12070);
nor UO_1342 (O_1342,N_11762,N_13786);
or UO_1343 (O_1343,N_11456,N_14746);
or UO_1344 (O_1344,N_14346,N_13488);
or UO_1345 (O_1345,N_10144,N_10616);
and UO_1346 (O_1346,N_11405,N_11901);
nand UO_1347 (O_1347,N_10733,N_10589);
nand UO_1348 (O_1348,N_14714,N_12883);
nor UO_1349 (O_1349,N_12783,N_13710);
and UO_1350 (O_1350,N_14492,N_13936);
nand UO_1351 (O_1351,N_10434,N_14358);
and UO_1352 (O_1352,N_10223,N_13455);
and UO_1353 (O_1353,N_12945,N_13470);
or UO_1354 (O_1354,N_14341,N_10927);
or UO_1355 (O_1355,N_12586,N_10584);
or UO_1356 (O_1356,N_14554,N_11100);
and UO_1357 (O_1357,N_11820,N_10148);
nor UO_1358 (O_1358,N_11921,N_10854);
nand UO_1359 (O_1359,N_11368,N_11840);
or UO_1360 (O_1360,N_11444,N_13212);
or UO_1361 (O_1361,N_12363,N_12854);
xnor UO_1362 (O_1362,N_11256,N_14065);
or UO_1363 (O_1363,N_10477,N_10315);
or UO_1364 (O_1364,N_10853,N_14412);
nand UO_1365 (O_1365,N_13145,N_14929);
nor UO_1366 (O_1366,N_11555,N_13382);
nand UO_1367 (O_1367,N_14563,N_14886);
nor UO_1368 (O_1368,N_13147,N_11301);
nor UO_1369 (O_1369,N_14952,N_14547);
nor UO_1370 (O_1370,N_13020,N_12105);
nand UO_1371 (O_1371,N_13328,N_10752);
nand UO_1372 (O_1372,N_14685,N_10919);
nand UO_1373 (O_1373,N_12438,N_13160);
or UO_1374 (O_1374,N_11638,N_11458);
and UO_1375 (O_1375,N_12365,N_13410);
nor UO_1376 (O_1376,N_13011,N_13074);
nor UO_1377 (O_1377,N_14667,N_14402);
or UO_1378 (O_1378,N_13207,N_11516);
nand UO_1379 (O_1379,N_12043,N_13767);
nor UO_1380 (O_1380,N_10237,N_10609);
nand UO_1381 (O_1381,N_10826,N_12653);
and UO_1382 (O_1382,N_12583,N_14266);
nor UO_1383 (O_1383,N_13618,N_12456);
or UO_1384 (O_1384,N_12333,N_11090);
nand UO_1385 (O_1385,N_13064,N_10447);
or UO_1386 (O_1386,N_12449,N_11869);
nor UO_1387 (O_1387,N_10691,N_12995);
nor UO_1388 (O_1388,N_10900,N_13121);
nor UO_1389 (O_1389,N_14400,N_10051);
nor UO_1390 (O_1390,N_14661,N_11582);
xor UO_1391 (O_1391,N_13101,N_11335);
or UO_1392 (O_1392,N_13449,N_14782);
nor UO_1393 (O_1393,N_13787,N_10983);
nor UO_1394 (O_1394,N_13905,N_12266);
nor UO_1395 (O_1395,N_13550,N_13742);
nor UO_1396 (O_1396,N_14514,N_11931);
nor UO_1397 (O_1397,N_10682,N_13223);
nor UO_1398 (O_1398,N_10595,N_12857);
nand UO_1399 (O_1399,N_12936,N_12834);
and UO_1400 (O_1400,N_10435,N_11775);
nand UO_1401 (O_1401,N_13129,N_10593);
nor UO_1402 (O_1402,N_10897,N_11440);
nand UO_1403 (O_1403,N_11253,N_11919);
nor UO_1404 (O_1404,N_12973,N_13345);
or UO_1405 (O_1405,N_10329,N_13811);
nand UO_1406 (O_1406,N_12782,N_13656);
nand UO_1407 (O_1407,N_14802,N_13997);
or UO_1408 (O_1408,N_14413,N_13584);
or UO_1409 (O_1409,N_12926,N_13807);
and UO_1410 (O_1410,N_10822,N_12420);
nor UO_1411 (O_1411,N_10712,N_13447);
nand UO_1412 (O_1412,N_10233,N_12289);
or UO_1413 (O_1413,N_11593,N_13419);
or UO_1414 (O_1414,N_11452,N_11000);
nor UO_1415 (O_1415,N_11084,N_11522);
or UO_1416 (O_1416,N_12380,N_13547);
and UO_1417 (O_1417,N_13878,N_13248);
and UO_1418 (O_1418,N_10423,N_11641);
and UO_1419 (O_1419,N_13304,N_13184);
and UO_1420 (O_1420,N_13616,N_10441);
or UO_1421 (O_1421,N_13943,N_12390);
nor UO_1422 (O_1422,N_11427,N_11993);
nand UO_1423 (O_1423,N_13515,N_13951);
and UO_1424 (O_1424,N_13686,N_13352);
and UO_1425 (O_1425,N_12276,N_11279);
or UO_1426 (O_1426,N_14068,N_13629);
nor UO_1427 (O_1427,N_12619,N_11429);
and UO_1428 (O_1428,N_10747,N_14691);
nand UO_1429 (O_1429,N_12963,N_13933);
nor UO_1430 (O_1430,N_14637,N_12738);
and UO_1431 (O_1431,N_13772,N_14435);
nor UO_1432 (O_1432,N_14191,N_13255);
nand UO_1433 (O_1433,N_14540,N_10459);
nor UO_1434 (O_1434,N_10745,N_10966);
and UO_1435 (O_1435,N_10222,N_13980);
nor UO_1436 (O_1436,N_10583,N_11462);
and UO_1437 (O_1437,N_14529,N_11068);
nand UO_1438 (O_1438,N_12477,N_10115);
and UO_1439 (O_1439,N_13368,N_13386);
or UO_1440 (O_1440,N_13993,N_12889);
nand UO_1441 (O_1441,N_14972,N_13115);
nor UO_1442 (O_1442,N_11114,N_14515);
or UO_1443 (O_1443,N_11185,N_10798);
nand UO_1444 (O_1444,N_12041,N_11724);
xnor UO_1445 (O_1445,N_13112,N_14815);
xnor UO_1446 (O_1446,N_11049,N_11946);
nor UO_1447 (O_1447,N_13329,N_13722);
nand UO_1448 (O_1448,N_10778,N_13364);
nor UO_1449 (O_1449,N_10505,N_11299);
nor UO_1450 (O_1450,N_11781,N_10873);
nor UO_1451 (O_1451,N_12897,N_10273);
nor UO_1452 (O_1452,N_11467,N_12515);
nand UO_1453 (O_1453,N_13330,N_10132);
nor UO_1454 (O_1454,N_12826,N_13971);
nor UO_1455 (O_1455,N_12519,N_12635);
and UO_1456 (O_1456,N_11945,N_12539);
nand UO_1457 (O_1457,N_11648,N_13611);
or UO_1458 (O_1458,N_14597,N_13429);
or UO_1459 (O_1459,N_14633,N_12402);
and UO_1460 (O_1460,N_12833,N_11783);
and UO_1461 (O_1461,N_12027,N_10187);
or UO_1462 (O_1462,N_14627,N_10298);
or UO_1463 (O_1463,N_11260,N_10891);
and UO_1464 (O_1464,N_12552,N_13276);
and UO_1465 (O_1465,N_12674,N_10617);
xor UO_1466 (O_1466,N_12168,N_13073);
and UO_1467 (O_1467,N_14561,N_14098);
nand UO_1468 (O_1468,N_10093,N_12088);
or UO_1469 (O_1469,N_12960,N_12850);
and UO_1470 (O_1470,N_12054,N_12678);
nand UO_1471 (O_1471,N_13655,N_14526);
or UO_1472 (O_1472,N_14201,N_12514);
and UO_1473 (O_1473,N_10167,N_11271);
nand UO_1474 (O_1474,N_13286,N_12980);
nor UO_1475 (O_1475,N_11718,N_10215);
and UO_1476 (O_1476,N_13946,N_10513);
or UO_1477 (O_1477,N_14351,N_12194);
or UO_1478 (O_1478,N_12581,N_11611);
and UO_1479 (O_1479,N_10579,N_10975);
and UO_1480 (O_1480,N_12733,N_10483);
nor UO_1481 (O_1481,N_12366,N_12752);
and UO_1482 (O_1482,N_10721,N_11872);
nand UO_1483 (O_1483,N_14502,N_13891);
nor UO_1484 (O_1484,N_12443,N_14284);
nand UO_1485 (O_1485,N_14553,N_14459);
nor UO_1486 (O_1486,N_11370,N_11617);
nand UO_1487 (O_1487,N_11630,N_13451);
nor UO_1488 (O_1488,N_11934,N_11241);
nand UO_1489 (O_1489,N_13941,N_10488);
nor UO_1490 (O_1490,N_14651,N_10714);
and UO_1491 (O_1491,N_11565,N_11226);
or UO_1492 (O_1492,N_10570,N_10046);
nand UO_1493 (O_1493,N_13083,N_12319);
nand UO_1494 (O_1494,N_12128,N_14256);
nor UO_1495 (O_1495,N_11338,N_13008);
and UO_1496 (O_1496,N_10769,N_10216);
nor UO_1497 (O_1497,N_14832,N_10387);
nand UO_1498 (O_1498,N_12796,N_12466);
nor UO_1499 (O_1499,N_14729,N_10774);
and UO_1500 (O_1500,N_13291,N_10663);
nor UO_1501 (O_1501,N_13785,N_14060);
and UO_1502 (O_1502,N_12600,N_12910);
and UO_1503 (O_1503,N_14796,N_10082);
nor UO_1504 (O_1504,N_13505,N_11537);
nor UO_1505 (O_1505,N_14762,N_12966);
and UO_1506 (O_1506,N_14793,N_11867);
xnor UO_1507 (O_1507,N_10577,N_11037);
nor UO_1508 (O_1508,N_14193,N_11670);
xnor UO_1509 (O_1509,N_12183,N_13763);
or UO_1510 (O_1510,N_10152,N_10720);
nand UO_1511 (O_1511,N_14015,N_10858);
and UO_1512 (O_1512,N_10385,N_10280);
nor UO_1513 (O_1513,N_10204,N_12325);
nor UO_1514 (O_1514,N_14456,N_10479);
or UO_1515 (O_1515,N_10707,N_11601);
nand UO_1516 (O_1516,N_14814,N_14807);
or UO_1517 (O_1517,N_13292,N_14559);
xor UO_1518 (O_1518,N_12301,N_14751);
and UO_1519 (O_1519,N_11696,N_14130);
nor UO_1520 (O_1520,N_13619,N_12478);
nor UO_1521 (O_1521,N_10833,N_12534);
and UO_1522 (O_1522,N_13010,N_14368);
and UO_1523 (O_1523,N_14910,N_14650);
nor UO_1524 (O_1524,N_10756,N_12472);
or UO_1525 (O_1525,N_11153,N_14968);
xor UO_1526 (O_1526,N_11924,N_11694);
nor UO_1527 (O_1527,N_10851,N_10244);
and UO_1528 (O_1528,N_10637,N_13155);
or UO_1529 (O_1529,N_10601,N_11671);
nor UO_1530 (O_1530,N_10493,N_14898);
or UO_1531 (O_1531,N_12371,N_13596);
nand UO_1532 (O_1532,N_10279,N_11635);
and UO_1533 (O_1533,N_11881,N_13441);
or UO_1534 (O_1534,N_14615,N_11481);
nor UO_1535 (O_1535,N_13502,N_12859);
or UO_1536 (O_1536,N_10991,N_13404);
or UO_1537 (O_1537,N_13513,N_12958);
nor UO_1538 (O_1538,N_14384,N_14683);
nand UO_1539 (O_1539,N_13415,N_10340);
or UO_1540 (O_1540,N_10884,N_13365);
nand UO_1541 (O_1541,N_10433,N_14528);
or UO_1542 (O_1542,N_10704,N_13950);
or UO_1543 (O_1543,N_13249,N_10212);
nor UO_1544 (O_1544,N_14158,N_12804);
nor UO_1545 (O_1545,N_10690,N_11166);
and UO_1546 (O_1546,N_12173,N_13436);
or UO_1547 (O_1547,N_14274,N_11578);
and UO_1548 (O_1548,N_11737,N_12188);
nand UO_1549 (O_1549,N_14179,N_14361);
or UO_1550 (O_1550,N_13072,N_14505);
or UO_1551 (O_1551,N_12637,N_10241);
and UO_1552 (O_1552,N_10910,N_10611);
nand UO_1553 (O_1553,N_13086,N_10834);
and UO_1554 (O_1554,N_13317,N_12651);
nor UO_1555 (O_1555,N_10994,N_13930);
and UO_1556 (O_1556,N_14572,N_13684);
nand UO_1557 (O_1557,N_12317,N_13174);
and UO_1558 (O_1558,N_10692,N_14803);
or UO_1559 (O_1559,N_14617,N_12648);
nand UO_1560 (O_1560,N_10977,N_11841);
or UO_1561 (O_1561,N_11360,N_10961);
nand UO_1562 (O_1562,N_10802,N_14437);
and UO_1563 (O_1563,N_11361,N_14064);
nor UO_1564 (O_1564,N_14525,N_11842);
nor UO_1565 (O_1565,N_10629,N_13095);
and UO_1566 (O_1566,N_14058,N_13050);
nand UO_1567 (O_1567,N_14152,N_13889);
and UO_1568 (O_1568,N_10007,N_14171);
or UO_1569 (O_1569,N_14332,N_14732);
or UO_1570 (O_1570,N_14214,N_13577);
nand UO_1571 (O_1571,N_14969,N_11416);
nor UO_1572 (O_1572,N_12460,N_12302);
nand UO_1573 (O_1573,N_13776,N_11194);
nand UO_1574 (O_1574,N_14712,N_14491);
nor UO_1575 (O_1575,N_10362,N_10765);
nand UO_1576 (O_1576,N_13864,N_13085);
and UO_1577 (O_1577,N_13491,N_13634);
or UO_1578 (O_1578,N_10185,N_13384);
and UO_1579 (O_1579,N_10914,N_12176);
nor UO_1580 (O_1580,N_13977,N_12451);
nand UO_1581 (O_1581,N_10238,N_13632);
and UO_1582 (O_1582,N_11159,N_10183);
nor UO_1583 (O_1583,N_12999,N_11273);
or UO_1584 (O_1584,N_13163,N_13972);
or UO_1585 (O_1585,N_12142,N_13545);
nor UO_1586 (O_1586,N_14738,N_13504);
or UO_1587 (O_1587,N_13099,N_10048);
or UO_1588 (O_1588,N_11141,N_11941);
and UO_1589 (O_1589,N_11101,N_12911);
nand UO_1590 (O_1590,N_13341,N_13332);
and UO_1591 (O_1591,N_13066,N_13895);
or UO_1592 (O_1592,N_11591,N_10490);
nor UO_1593 (O_1593,N_11438,N_14281);
and UO_1594 (O_1594,N_11888,N_14430);
nand UO_1595 (O_1595,N_10980,N_14279);
nor UO_1596 (O_1596,N_14768,N_10377);
and UO_1597 (O_1597,N_13426,N_14899);
nand UO_1598 (O_1598,N_12837,N_14995);
or UO_1599 (O_1599,N_13743,N_13670);
nand UO_1600 (O_1600,N_14618,N_11677);
nand UO_1601 (O_1601,N_13940,N_12213);
nor UO_1602 (O_1602,N_11615,N_14161);
nor UO_1603 (O_1603,N_13991,N_10715);
nor UO_1604 (O_1604,N_10814,N_13392);
and UO_1605 (O_1605,N_14693,N_13021);
nand UO_1606 (O_1606,N_10474,N_11404);
or UO_1607 (O_1607,N_12968,N_10049);
or UO_1608 (O_1608,N_11202,N_12214);
and UO_1609 (O_1609,N_11652,N_13161);
xnor UO_1610 (O_1610,N_10502,N_13285);
and UO_1611 (O_1611,N_12785,N_13068);
nor UO_1612 (O_1612,N_14461,N_12345);
and UO_1613 (O_1613,N_11056,N_10181);
or UO_1614 (O_1614,N_11035,N_12439);
or UO_1615 (O_1615,N_14737,N_11909);
and UO_1616 (O_1616,N_14149,N_12308);
nor UO_1617 (O_1617,N_14077,N_10865);
nor UO_1618 (O_1618,N_13401,N_10825);
nand UO_1619 (O_1619,N_13902,N_14104);
nand UO_1620 (O_1620,N_14857,N_14238);
and UO_1621 (O_1621,N_14640,N_11782);
nand UO_1622 (O_1622,N_13537,N_13151);
nand UO_1623 (O_1623,N_14273,N_14007);
nand UO_1624 (O_1624,N_14131,N_13225);
xor UO_1625 (O_1625,N_10410,N_12587);
nor UO_1626 (O_1626,N_10419,N_10193);
or UO_1627 (O_1627,N_13176,N_11399);
or UO_1628 (O_1628,N_10751,N_13310);
xor UO_1629 (O_1629,N_10018,N_13859);
nand UO_1630 (O_1630,N_12723,N_12134);
and UO_1631 (O_1631,N_13214,N_11709);
nor UO_1632 (O_1632,N_11640,N_12925);
nor UO_1633 (O_1633,N_11282,N_10921);
or UO_1634 (O_1634,N_14334,N_11072);
nor UO_1635 (O_1635,N_12540,N_11365);
and UO_1636 (O_1636,N_14047,N_14894);
or UO_1637 (O_1637,N_13354,N_14445);
or UO_1638 (O_1638,N_13781,N_10266);
nor UO_1639 (O_1639,N_13197,N_14882);
nor UO_1640 (O_1640,N_14828,N_14383);
nand UO_1641 (O_1641,N_13414,N_12535);
nand UO_1642 (O_1642,N_10603,N_11046);
nand UO_1643 (O_1643,N_10957,N_12254);
or UO_1644 (O_1644,N_13727,N_10813);
nor UO_1645 (O_1645,N_13712,N_10845);
and UO_1646 (O_1646,N_10242,N_13281);
nor UO_1647 (O_1647,N_14784,N_10819);
nor UO_1648 (O_1648,N_11390,N_11589);
nor UO_1649 (O_1649,N_14112,N_10713);
nand UO_1650 (O_1650,N_13851,N_10602);
or UO_1651 (O_1651,N_14084,N_12282);
and UO_1652 (O_1652,N_14847,N_12463);
nand UO_1653 (O_1653,N_11003,N_14063);
or UO_1654 (O_1654,N_14390,N_12049);
nor UO_1655 (O_1655,N_12341,N_11738);
and UO_1656 (O_1656,N_14029,N_11534);
and UO_1657 (O_1657,N_12576,N_11764);
and UO_1658 (O_1658,N_13858,N_10202);
nor UO_1659 (O_1659,N_11485,N_10976);
nand UO_1660 (O_1660,N_12712,N_10969);
nor UO_1661 (O_1661,N_11004,N_13043);
or UO_1662 (O_1662,N_10317,N_12786);
nand UO_1663 (O_1663,N_12113,N_14388);
nand UO_1664 (O_1664,N_13801,N_11209);
or UO_1665 (O_1665,N_14123,N_12978);
nand UO_1666 (O_1666,N_12150,N_12836);
nor UO_1667 (O_1667,N_10075,N_12551);
or UO_1668 (O_1668,N_11787,N_13372);
nand UO_1669 (O_1669,N_13783,N_13717);
and UO_1670 (O_1670,N_12655,N_14879);
nor UO_1671 (O_1671,N_13422,N_14340);
nor UO_1672 (O_1672,N_11231,N_13989);
or UO_1673 (O_1673,N_12238,N_11675);
nor UO_1674 (O_1674,N_13784,N_10790);
nor UO_1675 (O_1675,N_12618,N_12598);
nor UO_1676 (O_1676,N_13148,N_12154);
and UO_1677 (O_1677,N_10179,N_10998);
and UO_1678 (O_1678,N_11304,N_11140);
nand UO_1679 (O_1679,N_11719,N_13607);
or UO_1680 (O_1680,N_10381,N_12694);
nand UO_1681 (O_1681,N_14066,N_13648);
nor UO_1682 (O_1682,N_13986,N_10581);
and UO_1683 (O_1683,N_11394,N_11800);
nor UO_1684 (O_1684,N_14380,N_10767);
nand UO_1685 (O_1685,N_12005,N_13658);
nand UO_1686 (O_1686,N_11220,N_11333);
nand UO_1687 (O_1687,N_11935,N_13934);
nand UO_1688 (O_1688,N_10664,N_12119);
or UO_1689 (O_1689,N_13948,N_10486);
nand UO_1690 (O_1690,N_11556,N_12140);
nand UO_1691 (O_1691,N_14030,N_13378);
nand UO_1692 (O_1692,N_13253,N_11052);
nor UO_1693 (O_1693,N_10267,N_10348);
nor UO_1694 (O_1694,N_10346,N_10596);
and UO_1695 (O_1695,N_13469,N_10413);
and UO_1696 (O_1696,N_12411,N_14493);
nand UO_1697 (O_1697,N_12754,N_11698);
nor UO_1698 (O_1698,N_12844,N_10992);
or UO_1699 (O_1699,N_14299,N_10901);
and UO_1700 (O_1700,N_14132,N_14958);
nand UO_1701 (O_1701,N_12073,N_12413);
nand UO_1702 (O_1702,N_11674,N_10001);
nand UO_1703 (O_1703,N_11510,N_10892);
or UO_1704 (O_1704,N_11186,N_14343);
nor UO_1705 (O_1705,N_13699,N_13192);
nor UO_1706 (O_1706,N_12181,N_13403);
and UO_1707 (O_1707,N_12542,N_10859);
nand UO_1708 (O_1708,N_13606,N_10620);
nor UO_1709 (O_1709,N_14887,N_11663);
or UO_1710 (O_1710,N_11142,N_14244);
nand UO_1711 (O_1711,N_10528,N_14183);
or UO_1712 (O_1712,N_11826,N_14699);
and UO_1713 (O_1713,N_14513,N_10430);
nand UO_1714 (O_1714,N_10735,N_12628);
or UO_1715 (O_1715,N_14253,N_11844);
and UO_1716 (O_1716,N_14739,N_12151);
nand UO_1717 (O_1717,N_14636,N_14624);
nor UO_1718 (O_1718,N_14590,N_13391);
nor UO_1719 (O_1719,N_11588,N_14945);
or UO_1720 (O_1720,N_14062,N_13159);
or UO_1721 (O_1721,N_14092,N_13167);
and UO_1722 (O_1722,N_14408,N_13138);
nor UO_1723 (O_1723,N_12714,N_14907);
and UO_1724 (O_1724,N_13144,N_14846);
and UO_1725 (O_1725,N_12144,N_14544);
nor UO_1726 (O_1726,N_13608,N_13880);
and UO_1727 (O_1727,N_11163,N_10665);
and UO_1728 (O_1728,N_10955,N_13166);
or UO_1729 (O_1729,N_13792,N_10063);
and UO_1730 (O_1730,N_12745,N_10022);
or UO_1731 (O_1731,N_10742,N_12735);
or UO_1732 (O_1732,N_13875,N_10934);
nand UO_1733 (O_1733,N_11201,N_13393);
or UO_1734 (O_1734,N_11863,N_11228);
nand UO_1735 (O_1735,N_12546,N_13705);
and UO_1736 (O_1736,N_12506,N_10698);
and UO_1737 (O_1737,N_12962,N_14844);
nand UO_1738 (O_1738,N_10159,N_11339);
and UO_1739 (O_1739,N_10689,N_14944);
nor UO_1740 (O_1740,N_11544,N_14773);
and UO_1741 (O_1741,N_14359,N_13294);
nand UO_1742 (O_1742,N_11305,N_14262);
nor UO_1743 (O_1743,N_11357,N_10896);
and UO_1744 (O_1744,N_12503,N_10741);
and UO_1745 (O_1745,N_13312,N_14150);
nand UO_1746 (O_1746,N_12474,N_11126);
nor UO_1747 (O_1747,N_12211,N_10648);
nor UO_1748 (O_1748,N_13318,N_13178);
nor UO_1749 (O_1749,N_13719,N_12219);
nand UO_1750 (O_1750,N_12585,N_14057);
nand UO_1751 (O_1751,N_14558,N_10373);
nor UO_1752 (O_1752,N_14129,N_10659);
nor UO_1753 (O_1753,N_13028,N_12083);
and UO_1754 (O_1754,N_12174,N_11017);
nand UO_1755 (O_1755,N_14523,N_10963);
nand UO_1756 (O_1756,N_12189,N_14817);
nor UO_1757 (O_1757,N_10718,N_10327);
nand UO_1758 (O_1758,N_11423,N_11334);
nor UO_1759 (O_1759,N_12803,N_10875);
nor UO_1760 (O_1760,N_13283,N_10931);
nand UO_1761 (O_1761,N_11680,N_14850);
nand UO_1762 (O_1762,N_10913,N_13290);
nor UO_1763 (O_1763,N_12890,N_11837);
and UO_1764 (O_1764,N_11562,N_11352);
and UO_1765 (O_1765,N_14328,N_11469);
or UO_1766 (O_1766,N_14931,N_14369);
or UO_1767 (O_1767,N_12252,N_13030);
or UO_1768 (O_1768,N_11136,N_13427);
nand UO_1769 (O_1769,N_12852,N_11983);
nor UO_1770 (O_1770,N_12672,N_12934);
or UO_1771 (O_1771,N_10614,N_11414);
nor UO_1772 (O_1772,N_10906,N_11288);
nor UO_1773 (O_1773,N_13687,N_11183);
nand UO_1774 (O_1774,N_10066,N_10155);
nor UO_1775 (O_1775,N_10402,N_13760);
nor UO_1776 (O_1776,N_13377,N_11164);
nand UO_1777 (O_1777,N_14517,N_14593);
or UO_1778 (O_1778,N_10471,N_11525);
or UO_1779 (O_1779,N_11075,N_13036);
and UO_1780 (O_1780,N_14250,N_10156);
or UO_1781 (O_1781,N_10883,N_13216);
nand UO_1782 (O_1782,N_11441,N_13665);
and UO_1783 (O_1783,N_10396,N_13708);
or UO_1784 (O_1784,N_12076,N_12904);
and UO_1785 (O_1785,N_13974,N_12084);
nor UO_1786 (O_1786,N_10775,N_12633);
nor UO_1787 (O_1787,N_12631,N_12797);
or UO_1788 (O_1788,N_11326,N_10870);
nand UO_1789 (O_1789,N_12743,N_13206);
nor UO_1790 (O_1790,N_11459,N_14141);
and UO_1791 (O_1791,N_11975,N_14755);
nand UO_1792 (O_1792,N_10971,N_11246);
or UO_1793 (O_1793,N_11412,N_11465);
or UO_1794 (O_1794,N_12079,N_12601);
nor UO_1795 (O_1795,N_12727,N_12590);
nor UO_1796 (O_1796,N_12164,N_13509);
xor UO_1797 (O_1797,N_11953,N_13288);
nor UO_1798 (O_1798,N_12428,N_14716);
or UO_1799 (O_1799,N_12770,N_14026);
or UO_1800 (O_1800,N_11815,N_11908);
and UO_1801 (O_1801,N_10768,N_13485);
nand UO_1802 (O_1802,N_13081,N_13254);
nand UO_1803 (O_1803,N_14048,N_12090);
and UO_1804 (O_1804,N_10772,N_11223);
and UO_1805 (O_1805,N_12237,N_10281);
nor UO_1806 (O_1806,N_10119,N_11094);
or UO_1807 (O_1807,N_12988,N_10392);
nor UO_1808 (O_1808,N_12758,N_14680);
and UO_1809 (O_1809,N_12530,N_11803);
nor UO_1810 (O_1810,N_13346,N_10081);
and UO_1811 (O_1811,N_11501,N_10469);
nand UO_1812 (O_1812,N_11583,N_10368);
or UO_1813 (O_1813,N_13579,N_13061);
and UO_1814 (O_1814,N_14573,N_13725);
or UO_1815 (O_1815,N_10727,N_10177);
or UO_1816 (O_1816,N_10606,N_10669);
nor UO_1817 (O_1817,N_11981,N_14957);
or UO_1818 (O_1818,N_13418,N_10313);
or UO_1819 (O_1819,N_13751,N_12817);
and UO_1820 (O_1820,N_12613,N_10058);
nand UO_1821 (O_1821,N_13912,N_14904);
nand UO_1822 (O_1822,N_13493,N_10803);
or UO_1823 (O_1823,N_14099,N_14579);
and UO_1824 (O_1824,N_11595,N_12247);
nand UO_1825 (O_1825,N_11284,N_11532);
nor UO_1826 (O_1826,N_13911,N_10343);
nand UO_1827 (O_1827,N_11240,N_13210);
and UO_1828 (O_1828,N_14720,N_11463);
and UO_1829 (O_1829,N_14665,N_13630);
xnor UO_1830 (O_1830,N_12436,N_13522);
or UO_1831 (O_1831,N_11176,N_14113);
nor UO_1832 (O_1832,N_14641,N_10040);
and UO_1833 (O_1833,N_10277,N_14422);
or UO_1834 (O_1834,N_14468,N_13703);
nand UO_1835 (O_1835,N_13204,N_12593);
or UO_1836 (O_1836,N_13824,N_11758);
nand UO_1837 (O_1837,N_13321,N_11681);
and UO_1838 (O_1838,N_12643,N_14049);
and UO_1839 (O_1839,N_14087,N_11584);
nand UO_1840 (O_1840,N_10103,N_14892);
and UO_1841 (O_1841,N_10835,N_12036);
nor UO_1842 (O_1842,N_12609,N_11317);
nor UO_1843 (O_1843,N_14536,N_11213);
nand UO_1844 (O_1844,N_10070,N_11434);
or UO_1845 (O_1845,N_13543,N_10335);
nand UO_1846 (O_1846,N_11810,N_14115);
and UO_1847 (O_1847,N_11031,N_11265);
or UO_1848 (O_1848,N_13191,N_10126);
nand UO_1849 (O_1849,N_10524,N_14810);
and UO_1850 (O_1850,N_14283,N_10318);
nor UO_1851 (O_1851,N_10005,N_11926);
and UO_1852 (O_1852,N_12329,N_14471);
and UO_1853 (O_1853,N_12938,N_12349);
xor UO_1854 (O_1854,N_10987,N_11875);
or UO_1855 (O_1855,N_11119,N_10096);
nand UO_1856 (O_1856,N_13232,N_13107);
and UO_1857 (O_1857,N_14841,N_12225);
nor UO_1858 (O_1858,N_14926,N_10421);
or UO_1859 (O_1859,N_12136,N_11016);
nor UO_1860 (O_1860,N_11513,N_10289);
nor UO_1861 (O_1861,N_12537,N_13181);
nor UO_1862 (O_1862,N_12848,N_11900);
nand UO_1863 (O_1863,N_13667,N_12335);
and UO_1864 (O_1864,N_13102,N_10920);
nor UO_1865 (O_1865,N_10929,N_13609);
or UO_1866 (O_1866,N_10090,N_13425);
or UO_1867 (O_1867,N_10226,N_14896);
or UO_1868 (O_1868,N_13718,N_12830);
and UO_1869 (O_1869,N_12649,N_13413);
and UO_1870 (O_1870,N_12039,N_14288);
or UO_1871 (O_1871,N_14976,N_14877);
nand UO_1872 (O_1872,N_13340,N_14175);
or UO_1873 (O_1873,N_12939,N_14041);
and UO_1874 (O_1874,N_10706,N_14504);
and UO_1875 (O_1875,N_13019,N_14397);
or UO_1876 (O_1876,N_11269,N_11873);
nand UO_1877 (O_1877,N_12870,N_12404);
nor UO_1878 (O_1878,N_12578,N_14203);
nand UO_1879 (O_1879,N_14140,N_14639);
nand UO_1880 (O_1880,N_10674,N_14801);
nand UO_1881 (O_1881,N_10945,N_13589);
or UO_1882 (O_1882,N_14855,N_13387);
nand UO_1883 (O_1883,N_13704,N_10416);
and UO_1884 (O_1884,N_12849,N_10508);
or UO_1885 (O_1885,N_13421,N_11664);
nor UO_1886 (O_1886,N_12462,N_12499);
and UO_1887 (O_1887,N_10370,N_12498);
nand UO_1888 (O_1888,N_14764,N_12490);
nand UO_1889 (O_1889,N_12887,N_14600);
nand UO_1890 (O_1890,N_14286,N_11499);
or UO_1891 (O_1891,N_13740,N_13507);
nor UO_1892 (O_1892,N_11021,N_11504);
or UO_1893 (O_1893,N_10143,N_10746);
or UO_1894 (O_1894,N_13357,N_14360);
nand UO_1895 (O_1895,N_14999,N_14567);
and UO_1896 (O_1896,N_14054,N_10409);
and UO_1897 (O_1897,N_13519,N_10376);
nor UO_1898 (O_1898,N_11927,N_14257);
nand UO_1899 (O_1899,N_13603,N_13463);
nand UO_1900 (O_1900,N_13251,N_11002);
nand UO_1901 (O_1901,N_14448,N_14606);
nor UO_1902 (O_1902,N_13006,N_14006);
nand UO_1903 (O_1903,N_14546,N_12815);
nor UO_1904 (O_1904,N_10028,N_14766);
nor UO_1905 (O_1905,N_13736,N_10379);
nor UO_1906 (O_1906,N_13508,N_11665);
and UO_1907 (O_1907,N_14678,N_11212);
nor UO_1908 (O_1908,N_11711,N_11211);
nor UO_1909 (O_1909,N_14789,N_11296);
or UO_1910 (O_1910,N_10644,N_11018);
nor UO_1911 (O_1911,N_12422,N_10989);
and UO_1912 (O_1912,N_13960,N_11093);
nor UO_1913 (O_1913,N_13127,N_13227);
or UO_1914 (O_1914,N_14961,N_14834);
and UO_1915 (O_1915,N_12709,N_12948);
and UO_1916 (O_1916,N_13480,N_14144);
or UO_1917 (O_1917,N_14301,N_13187);
or UO_1918 (O_1918,N_13861,N_12875);
nor UO_1919 (O_1919,N_11316,N_11107);
nand UO_1920 (O_1920,N_12610,N_11409);
nand UO_1921 (O_1921,N_11300,N_10515);
and UO_1922 (O_1922,N_13692,N_14622);
nand UO_1923 (O_1923,N_13409,N_10425);
or UO_1924 (O_1924,N_13591,N_13876);
nand UO_1925 (O_1925,N_13242,N_12221);
and UO_1926 (O_1926,N_14511,N_11947);
or UO_1927 (O_1927,N_13284,N_14960);
or UO_1928 (O_1928,N_11645,N_11041);
xnor UO_1929 (O_1929,N_10219,N_14125);
nor UO_1930 (O_1930,N_11672,N_14993);
or UO_1931 (O_1931,N_10384,N_10021);
or UO_1932 (O_1932,N_14423,N_12577);
and UO_1933 (O_1933,N_10498,N_10060);
and UO_1934 (O_1934,N_13794,N_12495);
nor UO_1935 (O_1935,N_14165,N_12441);
and UO_1936 (O_1936,N_11280,N_12867);
nand UO_1937 (O_1937,N_13472,N_10503);
or UO_1938 (O_1938,N_13489,N_11856);
nor UO_1939 (O_1939,N_10024,N_13956);
nor UO_1940 (O_1940,N_12918,N_11590);
and UO_1941 (O_1941,N_13023,N_11950);
xnor UO_1942 (O_1942,N_10121,N_13026);
nor UO_1943 (O_1943,N_12638,N_11395);
or UO_1944 (O_1944,N_10388,N_12126);
nor UO_1945 (O_1945,N_11851,N_12907);
and UO_1946 (O_1946,N_11678,N_10299);
and UO_1947 (O_1947,N_11802,N_12589);
and UO_1948 (O_1948,N_14305,N_11549);
nor UO_1949 (O_1949,N_14365,N_12229);
and UO_1950 (O_1950,N_12360,N_13244);
and UO_1951 (O_1951,N_10728,N_12634);
nand UO_1952 (O_1952,N_12227,N_11868);
nand UO_1953 (O_1953,N_14880,N_13674);
and UO_1954 (O_1954,N_10292,N_14524);
and UO_1955 (O_1955,N_14936,N_13957);
nand UO_1956 (O_1956,N_13293,N_13534);
nand UO_1957 (O_1957,N_13925,N_10199);
or UO_1958 (O_1958,N_11354,N_10551);
or UO_1959 (O_1959,N_10578,N_10597);
and UO_1960 (O_1960,N_11668,N_14494);
nor UO_1961 (O_1961,N_14103,N_12004);
nand UO_1962 (O_1962,N_14354,N_12891);
nand UO_1963 (O_1963,N_13680,N_11417);
or UO_1964 (O_1964,N_12340,N_11125);
nor UO_1965 (O_1965,N_10068,N_11784);
nand UO_1966 (O_1966,N_12706,N_13240);
nor UO_1967 (O_1967,N_10635,N_13645);
nor UO_1968 (O_1968,N_10442,N_12101);
and UO_1969 (O_1969,N_13999,N_10220);
or UO_1970 (O_1970,N_10357,N_12479);
or UO_1971 (O_1971,N_12182,N_12218);
nor UO_1972 (O_1972,N_13666,N_12799);
and UO_1973 (O_1973,N_13967,N_13306);
nand UO_1974 (O_1974,N_11415,N_11257);
and UO_1975 (O_1975,N_11558,N_10079);
nand UO_1976 (O_1976,N_11509,N_13777);
nor UO_1977 (O_1977,N_12559,N_13170);
nand UO_1978 (O_1978,N_14666,N_14763);
nand UO_1979 (O_1979,N_12946,N_11098);
or UO_1980 (O_1980,N_10323,N_12471);
or UO_1981 (O_1981,N_14204,N_13075);
nand UO_1982 (O_1982,N_11124,N_14293);
nand UO_1983 (O_1983,N_12564,N_12082);
or UO_1984 (O_1984,N_14356,N_14776);
or UO_1985 (O_1985,N_10680,N_11831);
or UO_1986 (O_1986,N_13525,N_12051);
nand UO_1987 (O_1987,N_12617,N_11776);
and UO_1988 (O_1988,N_13694,N_11700);
and UO_1989 (O_1989,N_14194,N_11898);
nor UO_1990 (O_1990,N_14710,N_14777);
and UO_1991 (O_1991,N_10882,N_11605);
and UO_1992 (O_1992,N_14962,N_12825);
and UO_1993 (O_1993,N_11699,N_14488);
nand UO_1994 (O_1994,N_12232,N_12824);
and UO_1995 (O_1995,N_12708,N_10852);
nand UO_1996 (O_1996,N_13016,N_12812);
or UO_1997 (O_1997,N_13838,N_12323);
and UO_1998 (O_1998,N_12984,N_14925);
nand UO_1999 (O_1999,N_11191,N_11801);
endmodule