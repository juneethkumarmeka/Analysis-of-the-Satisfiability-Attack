module basic_500_3000_500_60_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_3,In_262);
nand U1 (N_1,In_97,In_404);
nor U2 (N_2,In_487,In_355);
or U3 (N_3,In_127,In_309);
or U4 (N_4,In_111,In_55);
and U5 (N_5,In_420,In_198);
and U6 (N_6,In_192,In_363);
or U7 (N_7,In_256,In_146);
nand U8 (N_8,In_277,In_341);
nor U9 (N_9,In_78,In_423);
nor U10 (N_10,In_128,In_467);
nand U11 (N_11,In_223,In_63);
and U12 (N_12,In_5,In_435);
and U13 (N_13,In_279,In_83);
and U14 (N_14,In_181,In_163);
nor U15 (N_15,In_483,In_178);
nor U16 (N_16,In_330,In_312);
and U17 (N_17,In_189,In_336);
nand U18 (N_18,In_106,In_314);
and U19 (N_19,In_327,In_145);
and U20 (N_20,In_286,In_75);
or U21 (N_21,In_61,In_313);
and U22 (N_22,In_46,In_406);
nor U23 (N_23,In_160,In_74);
nand U24 (N_24,In_477,In_369);
nor U25 (N_25,In_11,In_233);
nand U26 (N_26,In_284,In_271);
and U27 (N_27,In_441,In_134);
nor U28 (N_28,In_246,In_212);
nand U29 (N_29,In_305,In_356);
and U30 (N_30,In_138,In_428);
or U31 (N_31,In_370,In_278);
nor U32 (N_32,In_207,In_342);
nor U33 (N_33,In_195,In_110);
or U34 (N_34,In_155,In_352);
nand U35 (N_35,In_85,In_333);
nand U36 (N_36,In_65,In_325);
nand U37 (N_37,In_417,In_166);
and U38 (N_38,In_339,In_232);
nor U39 (N_39,In_269,In_402);
and U40 (N_40,In_209,In_48);
or U41 (N_41,In_40,In_267);
and U42 (N_42,In_432,In_371);
nand U43 (N_43,In_30,In_259);
nor U44 (N_44,In_20,In_457);
and U45 (N_45,In_306,In_250);
nand U46 (N_46,In_288,In_228);
and U47 (N_47,In_485,In_359);
nor U48 (N_48,In_401,In_105);
nor U49 (N_49,In_357,In_37);
or U50 (N_50,In_492,In_185);
nor U51 (N_51,In_98,In_95);
and U52 (N_52,In_307,In_320);
nor U53 (N_53,In_253,In_177);
nor U54 (N_54,In_414,In_431);
or U55 (N_55,In_495,In_135);
and U56 (N_56,In_291,In_454);
or U57 (N_57,In_67,In_488);
nand U58 (N_58,In_174,In_244);
xnor U59 (N_59,In_179,In_116);
nor U60 (N_60,In_335,In_26);
nor U61 (N_61,In_173,In_270);
nand U62 (N_62,In_167,N_3);
nand U63 (N_63,In_409,In_458);
or U64 (N_64,N_29,In_257);
or U65 (N_65,In_281,In_461);
nor U66 (N_66,In_41,In_443);
nand U67 (N_67,In_234,In_439);
or U68 (N_68,In_28,In_310);
and U69 (N_69,In_260,In_392);
or U70 (N_70,In_222,In_115);
or U71 (N_71,In_216,In_290);
and U72 (N_72,In_482,In_27);
or U73 (N_73,In_8,In_129);
or U74 (N_74,In_470,In_114);
nor U75 (N_75,In_358,In_491);
and U76 (N_76,In_112,In_194);
and U77 (N_77,In_6,In_452);
nand U78 (N_78,In_31,In_49);
nor U79 (N_79,N_32,In_263);
and U80 (N_80,In_239,In_360);
nand U81 (N_81,In_175,In_54);
and U82 (N_82,In_449,In_318);
nand U83 (N_83,In_438,In_351);
and U84 (N_84,In_468,In_39);
or U85 (N_85,N_18,In_453);
or U86 (N_86,In_153,In_165);
nor U87 (N_87,In_101,In_411);
or U88 (N_88,In_201,In_272);
or U89 (N_89,In_32,In_252);
or U90 (N_90,In_92,In_44);
and U91 (N_91,In_400,In_368);
nor U92 (N_92,In_455,In_413);
nand U93 (N_93,In_324,N_45);
nand U94 (N_94,N_43,In_231);
or U95 (N_95,In_407,In_149);
nand U96 (N_96,In_204,In_186);
nor U97 (N_97,In_247,In_385);
or U98 (N_98,In_136,In_133);
nand U99 (N_99,In_376,In_476);
or U100 (N_100,In_274,In_123);
or U101 (N_101,N_26,N_95);
nand U102 (N_102,N_67,In_462);
and U103 (N_103,In_171,In_447);
and U104 (N_104,In_268,In_121);
and U105 (N_105,In_465,In_226);
nand U106 (N_106,N_19,In_103);
nor U107 (N_107,In_182,In_399);
and U108 (N_108,In_132,In_162);
or U109 (N_109,In_70,N_76);
and U110 (N_110,In_19,In_345);
nand U111 (N_111,In_264,In_317);
nand U112 (N_112,In_499,In_445);
nand U113 (N_113,In_300,In_169);
nand U114 (N_114,In_130,In_120);
nand U115 (N_115,In_122,In_489);
and U116 (N_116,In_161,In_113);
nor U117 (N_117,N_44,N_55);
or U118 (N_118,In_148,In_29);
nor U119 (N_119,In_394,In_297);
nor U120 (N_120,In_493,In_79);
nand U121 (N_121,In_390,In_321);
nand U122 (N_122,In_346,In_47);
and U123 (N_123,In_299,In_202);
nor U124 (N_124,In_24,In_415);
or U125 (N_125,In_353,N_51);
or U126 (N_126,In_152,In_380);
nor U127 (N_127,In_191,In_304);
and U128 (N_128,N_53,N_71);
or U129 (N_129,N_72,In_450);
nand U130 (N_130,In_475,In_227);
or U131 (N_131,In_142,N_92);
nor U132 (N_132,In_375,N_86);
or U133 (N_133,In_301,In_190);
nand U134 (N_134,In_89,In_34);
nor U135 (N_135,In_294,In_296);
nand U136 (N_136,In_430,In_416);
xor U137 (N_137,In_285,In_347);
nor U138 (N_138,N_30,In_104);
nor U139 (N_139,In_200,N_68);
nand U140 (N_140,N_4,In_303);
and U141 (N_141,In_94,N_13);
nor U142 (N_142,In_283,N_69);
nor U143 (N_143,In_168,In_205);
nor U144 (N_144,In_344,In_157);
and U145 (N_145,In_282,In_211);
nor U146 (N_146,N_84,N_75);
nand U147 (N_147,In_151,In_56);
xnor U148 (N_148,In_275,In_422);
nand U149 (N_149,In_0,In_10);
or U150 (N_150,In_124,N_106);
nand U151 (N_151,N_46,N_52);
and U152 (N_152,In_315,In_102);
or U153 (N_153,In_57,N_128);
and U154 (N_154,In_52,N_1);
nor U155 (N_155,In_436,N_91);
nor U156 (N_156,N_120,N_80);
and U157 (N_157,In_463,N_73);
nor U158 (N_158,In_326,In_498);
or U159 (N_159,In_287,In_15);
or U160 (N_160,In_273,In_364);
and U161 (N_161,N_117,N_70);
and U162 (N_162,N_11,N_42);
xnor U163 (N_163,In_484,In_91);
nand U164 (N_164,N_7,N_24);
nand U165 (N_165,In_18,N_14);
nor U166 (N_166,N_2,In_295);
nor U167 (N_167,N_125,In_350);
nand U168 (N_168,In_480,In_90);
nor U169 (N_169,In_473,In_419);
or U170 (N_170,In_38,In_140);
or U171 (N_171,In_472,In_14);
and U172 (N_172,N_50,In_280);
or U173 (N_173,In_348,In_71);
nand U174 (N_174,N_134,In_214);
nor U175 (N_175,In_184,In_68);
nand U176 (N_176,N_116,N_109);
and U177 (N_177,In_446,In_340);
nand U178 (N_178,N_88,In_183);
or U179 (N_179,In_494,In_265);
nor U180 (N_180,In_4,N_60);
and U181 (N_181,In_354,In_448);
and U182 (N_182,N_145,In_60);
nor U183 (N_183,N_81,In_316);
and U184 (N_184,In_62,In_383);
nand U185 (N_185,In_210,In_403);
and U186 (N_186,In_84,In_224);
and U187 (N_187,N_123,N_110);
nor U188 (N_188,In_197,In_33);
and U189 (N_189,N_40,In_16);
or U190 (N_190,N_48,In_125);
or U191 (N_191,In_96,In_193);
or U192 (N_192,N_122,N_101);
nand U193 (N_193,N_115,N_58);
and U194 (N_194,In_1,In_119);
nor U195 (N_195,In_319,N_99);
nand U196 (N_196,In_377,In_382);
and U197 (N_197,In_444,In_218);
nor U198 (N_198,N_9,In_100);
and U199 (N_199,N_49,In_408);
nand U200 (N_200,In_241,In_66);
or U201 (N_201,In_64,In_393);
or U202 (N_202,N_118,N_28);
nand U203 (N_203,In_388,In_378);
nor U204 (N_204,In_53,In_405);
and U205 (N_205,N_138,In_7);
nor U206 (N_206,In_176,N_126);
nand U207 (N_207,N_196,N_178);
and U208 (N_208,In_158,In_237);
and U209 (N_209,N_121,In_93);
and U210 (N_210,In_249,In_386);
or U211 (N_211,N_12,In_410);
or U212 (N_212,N_63,In_42);
nor U213 (N_213,In_73,In_429);
nor U214 (N_214,N_17,N_157);
nand U215 (N_215,In_217,N_169);
nor U216 (N_216,N_93,In_235);
and U217 (N_217,In_397,N_187);
nor U218 (N_218,N_127,In_236);
and U219 (N_219,N_31,N_141);
nand U220 (N_220,N_82,N_78);
nor U221 (N_221,In_332,N_172);
and U222 (N_222,In_238,In_418);
and U223 (N_223,N_142,In_187);
nand U224 (N_224,In_206,In_289);
and U225 (N_225,In_343,N_94);
nand U226 (N_226,N_158,In_372);
nor U227 (N_227,N_148,N_0);
or U228 (N_228,N_171,In_466);
or U229 (N_229,N_27,N_140);
and U230 (N_230,In_384,N_168);
or U231 (N_231,N_165,In_391);
and U232 (N_232,N_192,N_112);
nand U233 (N_233,N_90,N_35);
nand U234 (N_234,In_107,N_186);
and U235 (N_235,In_334,In_424);
nand U236 (N_236,N_124,In_150);
nor U237 (N_237,N_6,N_83);
and U238 (N_238,N_195,N_89);
nand U239 (N_239,N_22,In_254);
and U240 (N_240,In_86,In_59);
and U241 (N_241,N_54,In_311);
or U242 (N_242,In_242,In_219);
and U243 (N_243,N_143,N_132);
nand U244 (N_244,In_373,In_76);
and U245 (N_245,In_456,N_175);
and U246 (N_246,N_25,In_398);
or U247 (N_247,In_365,N_34);
nor U248 (N_248,N_21,In_328);
nor U249 (N_249,In_395,N_155);
or U250 (N_250,N_36,N_216);
nand U251 (N_251,N_194,N_162);
nand U252 (N_252,N_247,N_41);
and U253 (N_253,In_460,In_88);
and U254 (N_254,N_136,In_17);
nor U255 (N_255,N_160,N_104);
and U256 (N_256,N_199,N_166);
nand U257 (N_257,N_150,In_87);
and U258 (N_258,In_143,N_62);
and U259 (N_259,N_225,In_387);
nand U260 (N_260,N_176,N_198);
nand U261 (N_261,N_193,N_77);
nand U262 (N_262,In_433,N_65);
nand U263 (N_263,N_102,N_203);
nand U264 (N_264,In_170,In_118);
and U265 (N_265,N_87,N_179);
or U266 (N_266,In_12,In_337);
and U267 (N_267,N_10,N_249);
xor U268 (N_268,In_258,In_230);
and U269 (N_269,In_126,In_381);
nand U270 (N_270,N_200,N_243);
and U271 (N_271,In_137,In_50);
nand U272 (N_272,N_227,N_222);
and U273 (N_273,N_137,N_208);
or U274 (N_274,N_246,N_244);
nor U275 (N_275,N_129,N_131);
nand U276 (N_276,N_201,N_156);
nand U277 (N_277,In_9,In_481);
or U278 (N_278,N_97,N_100);
nor U279 (N_279,N_241,N_139);
nor U280 (N_280,In_486,N_66);
or U281 (N_281,N_173,N_191);
or U282 (N_282,In_362,In_425);
and U283 (N_283,In_25,N_107);
nand U284 (N_284,N_189,In_229);
nor U285 (N_285,N_239,N_61);
and U286 (N_286,In_266,N_33);
nand U287 (N_287,In_23,N_237);
nand U288 (N_288,N_238,In_220);
and U289 (N_289,In_43,In_13);
nor U290 (N_290,N_230,N_228);
and U291 (N_291,In_199,N_232);
nor U292 (N_292,N_153,N_236);
or U293 (N_293,In_338,In_164);
nor U294 (N_294,N_108,N_130);
and U295 (N_295,In_180,N_159);
or U296 (N_296,In_82,In_440);
and U297 (N_297,In_35,N_229);
nand U298 (N_298,In_225,N_174);
or U299 (N_299,N_38,In_80);
or U300 (N_300,N_16,In_427);
and U301 (N_301,N_161,In_261);
or U302 (N_302,In_479,In_331);
or U303 (N_303,N_164,In_255);
nor U304 (N_304,N_245,N_184);
and U305 (N_305,N_218,N_177);
nand U306 (N_306,N_255,In_117);
or U307 (N_307,N_215,In_276);
or U308 (N_308,N_272,N_220);
and U309 (N_309,In_240,N_96);
and U310 (N_310,N_273,N_202);
nor U311 (N_311,N_226,N_250);
or U312 (N_312,N_251,In_77);
or U313 (N_313,N_268,N_113);
nor U314 (N_314,In_434,N_296);
nor U315 (N_315,N_224,N_151);
nand U316 (N_316,In_292,In_469);
or U317 (N_317,N_213,N_205);
and U318 (N_318,In_474,N_144);
nor U319 (N_319,In_322,In_221);
nand U320 (N_320,N_154,In_497);
and U321 (N_321,N_149,N_15);
nor U322 (N_322,N_254,N_188);
nor U323 (N_323,In_2,N_182);
nand U324 (N_324,N_264,N_287);
or U325 (N_325,In_159,N_275);
and U326 (N_326,In_437,N_231);
nor U327 (N_327,In_144,N_214);
nand U328 (N_328,N_103,In_22);
and U329 (N_329,In_251,N_85);
and U330 (N_330,In_293,N_133);
or U331 (N_331,N_210,N_293);
and U332 (N_332,In_426,N_185);
nor U333 (N_333,N_211,N_292);
nor U334 (N_334,N_280,In_196);
and U335 (N_335,In_109,N_56);
nor U336 (N_336,In_349,N_283);
nand U337 (N_337,In_367,In_298);
nand U338 (N_338,N_180,N_290);
nand U339 (N_339,N_266,N_274);
nor U340 (N_340,N_265,N_285);
nor U341 (N_341,In_139,N_288);
nand U342 (N_342,In_478,In_459);
nand U343 (N_343,N_114,N_147);
nand U344 (N_344,N_276,N_267);
nor U345 (N_345,In_396,In_45);
or U346 (N_346,N_98,In_374);
and U347 (N_347,N_5,N_260);
nand U348 (N_348,In_208,N_253);
nor U349 (N_349,N_286,N_242);
nor U350 (N_350,N_248,N_306);
and U351 (N_351,N_20,N_324);
nor U352 (N_352,N_233,N_281);
nor U353 (N_353,N_291,N_321);
and U354 (N_354,N_340,N_146);
nand U355 (N_355,N_278,N_39);
and U356 (N_356,N_105,In_323);
nand U357 (N_357,N_269,N_341);
or U358 (N_358,N_47,In_108);
and U359 (N_359,N_261,N_263);
or U360 (N_360,N_335,N_345);
nand U361 (N_361,N_344,N_343);
nor U362 (N_362,In_442,N_135);
nor U363 (N_363,N_257,N_308);
nor U364 (N_364,N_119,N_311);
nor U365 (N_365,N_183,In_471);
and U366 (N_366,In_329,N_302);
or U367 (N_367,In_141,N_303);
nand U368 (N_368,In_21,N_339);
and U369 (N_369,N_314,N_282);
nor U370 (N_370,N_299,In_361);
nor U371 (N_371,N_307,N_317);
nor U372 (N_372,N_197,N_346);
nand U373 (N_373,N_295,In_215);
and U374 (N_374,N_338,In_245);
or U375 (N_375,N_337,N_315);
nor U376 (N_376,N_334,In_51);
or U377 (N_377,N_331,N_310);
nor U378 (N_378,N_320,N_223);
and U379 (N_379,N_23,N_207);
nor U380 (N_380,N_209,N_259);
or U381 (N_381,In_451,N_206);
nor U382 (N_382,In_72,N_219);
nor U383 (N_383,N_79,N_326);
and U384 (N_384,In_36,In_213);
nor U385 (N_385,N_111,N_298);
and U386 (N_386,N_204,N_37);
nand U387 (N_387,In_203,N_74);
and U388 (N_388,N_212,In_156);
nor U389 (N_389,N_349,N_297);
nor U390 (N_390,In_366,N_336);
or U391 (N_391,In_248,N_167);
nand U392 (N_392,N_234,In_188);
and U393 (N_393,N_270,N_342);
and U394 (N_394,N_284,N_258);
nand U395 (N_395,In_147,N_348);
nor U396 (N_396,N_312,N_294);
or U397 (N_397,N_289,N_240);
nor U398 (N_398,N_163,N_152);
nand U399 (N_399,In_379,N_318);
nand U400 (N_400,N_170,N_333);
nor U401 (N_401,N_356,In_302);
and U402 (N_402,N_300,N_370);
or U403 (N_403,N_316,N_362);
nand U404 (N_404,N_377,N_279);
or U405 (N_405,N_369,N_390);
or U406 (N_406,N_359,In_99);
and U407 (N_407,N_366,N_373);
xnor U408 (N_408,N_397,N_386);
nor U409 (N_409,N_313,N_59);
or U410 (N_410,In_154,N_360);
nor U411 (N_411,N_389,N_271);
xnor U412 (N_412,N_319,N_325);
or U413 (N_413,N_304,N_64);
nor U414 (N_414,N_384,N_375);
nor U415 (N_415,In_412,N_395);
or U416 (N_416,In_490,N_367);
nand U417 (N_417,N_378,In_131);
or U418 (N_418,N_329,N_394);
or U419 (N_419,N_217,N_382);
or U420 (N_420,N_305,N_374);
nand U421 (N_421,N_392,In_464);
or U422 (N_422,N_357,N_381);
and U423 (N_423,N_388,N_301);
nor U424 (N_424,N_277,N_350);
nand U425 (N_425,N_376,N_332);
xnor U426 (N_426,In_172,N_355);
nor U427 (N_427,N_235,N_398);
and U428 (N_428,N_309,N_354);
nor U429 (N_429,N_383,N_353);
and U430 (N_430,In_308,N_190);
nand U431 (N_431,N_387,N_352);
nor U432 (N_432,N_347,N_252);
nand U433 (N_433,N_330,In_496);
nor U434 (N_434,N_379,N_351);
nor U435 (N_435,N_256,N_380);
nand U436 (N_436,N_372,N_363);
nand U437 (N_437,N_327,N_364);
and U438 (N_438,N_8,In_421);
and U439 (N_439,N_393,N_322);
nor U440 (N_440,N_328,N_391);
or U441 (N_441,In_243,In_81);
and U442 (N_442,N_323,N_358);
or U443 (N_443,N_371,N_385);
and U444 (N_444,N_262,N_365);
or U445 (N_445,N_221,N_399);
and U446 (N_446,In_58,N_361);
nand U447 (N_447,N_181,N_57);
and U448 (N_448,In_389,N_396);
and U449 (N_449,N_368,In_69);
and U450 (N_450,N_416,N_415);
and U451 (N_451,N_422,N_408);
nand U452 (N_452,N_443,N_405);
nand U453 (N_453,N_428,N_435);
or U454 (N_454,N_427,N_404);
or U455 (N_455,N_418,N_436);
and U456 (N_456,N_411,N_413);
and U457 (N_457,N_433,N_432);
nand U458 (N_458,N_421,N_417);
and U459 (N_459,N_441,N_447);
or U460 (N_460,N_446,N_424);
nand U461 (N_461,N_400,N_409);
and U462 (N_462,N_414,N_407);
nand U463 (N_463,N_445,N_449);
nand U464 (N_464,N_406,N_403);
nor U465 (N_465,N_430,N_439);
or U466 (N_466,N_444,N_431);
nand U467 (N_467,N_410,N_412);
or U468 (N_468,N_438,N_420);
and U469 (N_469,N_434,N_401);
and U470 (N_470,N_425,N_437);
or U471 (N_471,N_423,N_419);
nand U472 (N_472,N_429,N_440);
nand U473 (N_473,N_426,N_448);
and U474 (N_474,N_442,N_402);
and U475 (N_475,N_440,N_421);
nand U476 (N_476,N_441,N_425);
or U477 (N_477,N_438,N_437);
nor U478 (N_478,N_418,N_439);
nand U479 (N_479,N_422,N_440);
nand U480 (N_480,N_445,N_427);
or U481 (N_481,N_448,N_412);
and U482 (N_482,N_433,N_414);
nand U483 (N_483,N_437,N_419);
or U484 (N_484,N_434,N_444);
nand U485 (N_485,N_433,N_420);
nor U486 (N_486,N_433,N_429);
nand U487 (N_487,N_431,N_403);
nor U488 (N_488,N_445,N_428);
nor U489 (N_489,N_414,N_434);
nand U490 (N_490,N_443,N_420);
nor U491 (N_491,N_427,N_431);
nand U492 (N_492,N_424,N_436);
nand U493 (N_493,N_439,N_407);
or U494 (N_494,N_427,N_423);
and U495 (N_495,N_419,N_447);
nand U496 (N_496,N_401,N_408);
or U497 (N_497,N_449,N_408);
and U498 (N_498,N_422,N_401);
nand U499 (N_499,N_426,N_410);
and U500 (N_500,N_456,N_491);
or U501 (N_501,N_474,N_462);
or U502 (N_502,N_473,N_483);
xor U503 (N_503,N_488,N_486);
nor U504 (N_504,N_471,N_452);
or U505 (N_505,N_489,N_459);
and U506 (N_506,N_485,N_450);
nand U507 (N_507,N_484,N_451);
nor U508 (N_508,N_479,N_463);
and U509 (N_509,N_464,N_467);
and U510 (N_510,N_470,N_475);
nor U511 (N_511,N_477,N_466);
nand U512 (N_512,N_487,N_480);
nor U513 (N_513,N_494,N_469);
nand U514 (N_514,N_497,N_455);
nand U515 (N_515,N_492,N_457);
and U516 (N_516,N_499,N_493);
nand U517 (N_517,N_476,N_481);
nand U518 (N_518,N_453,N_478);
nand U519 (N_519,N_498,N_482);
nor U520 (N_520,N_490,N_460);
or U521 (N_521,N_458,N_461);
or U522 (N_522,N_468,N_495);
and U523 (N_523,N_496,N_472);
nand U524 (N_524,N_465,N_454);
and U525 (N_525,N_481,N_454);
or U526 (N_526,N_469,N_479);
nand U527 (N_527,N_482,N_462);
nor U528 (N_528,N_468,N_462);
nor U529 (N_529,N_455,N_461);
or U530 (N_530,N_466,N_496);
nand U531 (N_531,N_482,N_457);
and U532 (N_532,N_451,N_472);
or U533 (N_533,N_467,N_466);
and U534 (N_534,N_463,N_453);
or U535 (N_535,N_450,N_467);
xnor U536 (N_536,N_467,N_465);
or U537 (N_537,N_487,N_472);
nand U538 (N_538,N_487,N_479);
or U539 (N_539,N_486,N_459);
and U540 (N_540,N_475,N_462);
xor U541 (N_541,N_459,N_476);
or U542 (N_542,N_458,N_493);
and U543 (N_543,N_473,N_481);
nand U544 (N_544,N_488,N_490);
and U545 (N_545,N_472,N_475);
or U546 (N_546,N_465,N_474);
and U547 (N_547,N_450,N_470);
and U548 (N_548,N_482,N_492);
and U549 (N_549,N_458,N_454);
or U550 (N_550,N_521,N_503);
and U551 (N_551,N_516,N_530);
xor U552 (N_552,N_515,N_547);
or U553 (N_553,N_548,N_532);
and U554 (N_554,N_512,N_538);
or U555 (N_555,N_540,N_534);
nand U556 (N_556,N_533,N_504);
nand U557 (N_557,N_546,N_519);
nor U558 (N_558,N_549,N_500);
nand U559 (N_559,N_523,N_502);
nor U560 (N_560,N_545,N_535);
nand U561 (N_561,N_536,N_529);
nor U562 (N_562,N_541,N_539);
or U563 (N_563,N_513,N_542);
nand U564 (N_564,N_518,N_544);
or U565 (N_565,N_505,N_506);
or U566 (N_566,N_509,N_537);
and U567 (N_567,N_525,N_508);
nor U568 (N_568,N_520,N_507);
nand U569 (N_569,N_522,N_526);
and U570 (N_570,N_527,N_528);
or U571 (N_571,N_514,N_543);
nor U572 (N_572,N_524,N_517);
or U573 (N_573,N_511,N_501);
and U574 (N_574,N_531,N_510);
nor U575 (N_575,N_521,N_517);
nand U576 (N_576,N_538,N_543);
nand U577 (N_577,N_535,N_532);
or U578 (N_578,N_544,N_504);
nand U579 (N_579,N_531,N_543);
or U580 (N_580,N_532,N_539);
or U581 (N_581,N_507,N_547);
and U582 (N_582,N_545,N_502);
nor U583 (N_583,N_546,N_503);
or U584 (N_584,N_512,N_518);
nor U585 (N_585,N_535,N_503);
nand U586 (N_586,N_529,N_548);
or U587 (N_587,N_549,N_509);
and U588 (N_588,N_546,N_547);
nor U589 (N_589,N_502,N_532);
and U590 (N_590,N_540,N_519);
nor U591 (N_591,N_535,N_527);
or U592 (N_592,N_531,N_525);
and U593 (N_593,N_549,N_520);
or U594 (N_594,N_513,N_532);
nand U595 (N_595,N_518,N_549);
nor U596 (N_596,N_523,N_513);
nand U597 (N_597,N_530,N_513);
and U598 (N_598,N_532,N_509);
or U599 (N_599,N_504,N_509);
nand U600 (N_600,N_551,N_556);
nor U601 (N_601,N_552,N_581);
and U602 (N_602,N_567,N_591);
or U603 (N_603,N_573,N_599);
or U604 (N_604,N_590,N_575);
and U605 (N_605,N_589,N_561);
nand U606 (N_606,N_558,N_566);
and U607 (N_607,N_582,N_596);
and U608 (N_608,N_571,N_586);
or U609 (N_609,N_559,N_587);
or U610 (N_610,N_563,N_580);
and U611 (N_611,N_583,N_553);
nor U612 (N_612,N_593,N_562);
nor U613 (N_613,N_570,N_594);
or U614 (N_614,N_598,N_585);
nor U615 (N_615,N_557,N_577);
and U616 (N_616,N_555,N_579);
nand U617 (N_617,N_560,N_550);
or U618 (N_618,N_588,N_597);
nor U619 (N_619,N_592,N_554);
or U620 (N_620,N_595,N_564);
and U621 (N_621,N_568,N_572);
and U622 (N_622,N_584,N_574);
and U623 (N_623,N_569,N_576);
or U624 (N_624,N_578,N_565);
nand U625 (N_625,N_574,N_589);
and U626 (N_626,N_552,N_599);
nor U627 (N_627,N_556,N_594);
or U628 (N_628,N_586,N_577);
nor U629 (N_629,N_554,N_569);
or U630 (N_630,N_566,N_550);
or U631 (N_631,N_551,N_589);
and U632 (N_632,N_557,N_595);
nand U633 (N_633,N_558,N_583);
or U634 (N_634,N_561,N_587);
and U635 (N_635,N_574,N_579);
nand U636 (N_636,N_565,N_584);
or U637 (N_637,N_586,N_596);
or U638 (N_638,N_569,N_597);
nor U639 (N_639,N_580,N_590);
nor U640 (N_640,N_576,N_594);
nor U641 (N_641,N_566,N_563);
nor U642 (N_642,N_595,N_571);
or U643 (N_643,N_560,N_588);
and U644 (N_644,N_578,N_562);
or U645 (N_645,N_582,N_576);
nand U646 (N_646,N_593,N_561);
or U647 (N_647,N_567,N_584);
and U648 (N_648,N_567,N_576);
or U649 (N_649,N_594,N_554);
or U650 (N_650,N_642,N_628);
and U651 (N_651,N_609,N_629);
nor U652 (N_652,N_639,N_631);
nor U653 (N_653,N_638,N_610);
nor U654 (N_654,N_603,N_643);
and U655 (N_655,N_623,N_635);
or U656 (N_656,N_611,N_640);
and U657 (N_657,N_617,N_620);
and U658 (N_658,N_600,N_602);
nand U659 (N_659,N_606,N_637);
or U660 (N_660,N_626,N_613);
nand U661 (N_661,N_648,N_614);
and U662 (N_662,N_627,N_646);
and U663 (N_663,N_621,N_649);
xnor U664 (N_664,N_608,N_644);
nor U665 (N_665,N_607,N_605);
or U666 (N_666,N_630,N_625);
and U667 (N_667,N_622,N_647);
and U668 (N_668,N_619,N_618);
or U669 (N_669,N_615,N_636);
or U670 (N_670,N_604,N_601);
nor U671 (N_671,N_624,N_616);
nand U672 (N_672,N_612,N_632);
or U673 (N_673,N_634,N_641);
and U674 (N_674,N_645,N_633);
nor U675 (N_675,N_616,N_627);
nand U676 (N_676,N_628,N_619);
and U677 (N_677,N_640,N_635);
and U678 (N_678,N_622,N_617);
or U679 (N_679,N_639,N_649);
and U680 (N_680,N_607,N_641);
and U681 (N_681,N_610,N_611);
and U682 (N_682,N_637,N_622);
nor U683 (N_683,N_617,N_605);
and U684 (N_684,N_645,N_606);
or U685 (N_685,N_605,N_640);
or U686 (N_686,N_641,N_616);
nor U687 (N_687,N_610,N_635);
nand U688 (N_688,N_643,N_604);
and U689 (N_689,N_629,N_634);
or U690 (N_690,N_603,N_629);
nand U691 (N_691,N_641,N_638);
or U692 (N_692,N_614,N_618);
nor U693 (N_693,N_646,N_638);
nor U694 (N_694,N_637,N_615);
and U695 (N_695,N_608,N_614);
nor U696 (N_696,N_646,N_622);
nand U697 (N_697,N_607,N_632);
or U698 (N_698,N_613,N_612);
nand U699 (N_699,N_609,N_634);
or U700 (N_700,N_679,N_659);
nand U701 (N_701,N_682,N_657);
or U702 (N_702,N_690,N_697);
or U703 (N_703,N_694,N_663);
or U704 (N_704,N_685,N_674);
nor U705 (N_705,N_669,N_660);
or U706 (N_706,N_658,N_664);
nand U707 (N_707,N_673,N_654);
nor U708 (N_708,N_650,N_689);
and U709 (N_709,N_666,N_684);
or U710 (N_710,N_683,N_653);
nor U711 (N_711,N_667,N_670);
nor U712 (N_712,N_681,N_698);
nor U713 (N_713,N_668,N_661);
and U714 (N_714,N_652,N_678);
nand U715 (N_715,N_656,N_671);
nor U716 (N_716,N_677,N_695);
nor U717 (N_717,N_672,N_662);
and U718 (N_718,N_691,N_686);
or U719 (N_719,N_665,N_688);
or U720 (N_720,N_680,N_699);
nand U721 (N_721,N_692,N_676);
xor U722 (N_722,N_651,N_655);
nor U723 (N_723,N_693,N_696);
nand U724 (N_724,N_675,N_687);
nand U725 (N_725,N_678,N_671);
nand U726 (N_726,N_698,N_650);
nor U727 (N_727,N_684,N_693);
nand U728 (N_728,N_699,N_677);
nand U729 (N_729,N_693,N_650);
nand U730 (N_730,N_661,N_677);
and U731 (N_731,N_681,N_664);
or U732 (N_732,N_667,N_696);
nor U733 (N_733,N_673,N_697);
or U734 (N_734,N_654,N_666);
or U735 (N_735,N_681,N_658);
and U736 (N_736,N_688,N_664);
and U737 (N_737,N_655,N_695);
nor U738 (N_738,N_682,N_690);
and U739 (N_739,N_668,N_672);
nor U740 (N_740,N_664,N_652);
nor U741 (N_741,N_672,N_691);
and U742 (N_742,N_681,N_663);
or U743 (N_743,N_655,N_693);
or U744 (N_744,N_654,N_698);
and U745 (N_745,N_668,N_699);
or U746 (N_746,N_660,N_699);
nor U747 (N_747,N_653,N_684);
nor U748 (N_748,N_697,N_689);
nand U749 (N_749,N_683,N_689);
nor U750 (N_750,N_742,N_730);
nor U751 (N_751,N_703,N_709);
or U752 (N_752,N_743,N_727);
nor U753 (N_753,N_724,N_735);
nor U754 (N_754,N_741,N_719);
nand U755 (N_755,N_748,N_701);
nor U756 (N_756,N_712,N_732);
and U757 (N_757,N_737,N_720);
nand U758 (N_758,N_749,N_723);
or U759 (N_759,N_713,N_718);
or U760 (N_760,N_729,N_739);
nand U761 (N_761,N_710,N_731);
nand U762 (N_762,N_711,N_704);
or U763 (N_763,N_706,N_716);
nor U764 (N_764,N_733,N_705);
nor U765 (N_765,N_702,N_707);
or U766 (N_766,N_700,N_728);
and U767 (N_767,N_746,N_745);
or U768 (N_768,N_725,N_736);
and U769 (N_769,N_721,N_726);
or U770 (N_770,N_717,N_734);
nor U771 (N_771,N_738,N_722);
nor U772 (N_772,N_740,N_708);
nand U773 (N_773,N_744,N_747);
nand U774 (N_774,N_715,N_714);
nand U775 (N_775,N_733,N_704);
nand U776 (N_776,N_732,N_720);
or U777 (N_777,N_716,N_705);
nor U778 (N_778,N_728,N_748);
nor U779 (N_779,N_710,N_707);
and U780 (N_780,N_738,N_729);
nand U781 (N_781,N_738,N_736);
and U782 (N_782,N_712,N_731);
nand U783 (N_783,N_715,N_702);
or U784 (N_784,N_744,N_727);
nor U785 (N_785,N_734,N_702);
nor U786 (N_786,N_723,N_705);
nand U787 (N_787,N_740,N_713);
and U788 (N_788,N_723,N_711);
and U789 (N_789,N_749,N_719);
xnor U790 (N_790,N_723,N_737);
nor U791 (N_791,N_742,N_711);
and U792 (N_792,N_735,N_733);
nor U793 (N_793,N_706,N_719);
or U794 (N_794,N_737,N_702);
xnor U795 (N_795,N_735,N_729);
or U796 (N_796,N_735,N_734);
and U797 (N_797,N_743,N_720);
and U798 (N_798,N_704,N_709);
and U799 (N_799,N_731,N_715);
or U800 (N_800,N_784,N_773);
or U801 (N_801,N_762,N_761);
and U802 (N_802,N_777,N_754);
nor U803 (N_803,N_766,N_751);
or U804 (N_804,N_771,N_764);
or U805 (N_805,N_787,N_752);
and U806 (N_806,N_763,N_753);
nor U807 (N_807,N_798,N_790);
nand U808 (N_808,N_796,N_760);
nand U809 (N_809,N_788,N_759);
nor U810 (N_810,N_786,N_769);
nor U811 (N_811,N_757,N_770);
and U812 (N_812,N_780,N_795);
nand U813 (N_813,N_775,N_774);
or U814 (N_814,N_793,N_768);
and U815 (N_815,N_791,N_781);
and U816 (N_816,N_778,N_767);
or U817 (N_817,N_750,N_799);
or U818 (N_818,N_765,N_758);
nor U819 (N_819,N_782,N_789);
and U820 (N_820,N_772,N_792);
nor U821 (N_821,N_797,N_755);
and U822 (N_822,N_779,N_776);
nor U823 (N_823,N_756,N_783);
and U824 (N_824,N_794,N_785);
and U825 (N_825,N_774,N_777);
and U826 (N_826,N_799,N_790);
or U827 (N_827,N_780,N_752);
nand U828 (N_828,N_796,N_799);
or U829 (N_829,N_792,N_774);
and U830 (N_830,N_777,N_789);
nand U831 (N_831,N_752,N_789);
or U832 (N_832,N_783,N_754);
or U833 (N_833,N_790,N_754);
and U834 (N_834,N_789,N_794);
or U835 (N_835,N_770,N_779);
nor U836 (N_836,N_762,N_793);
nor U837 (N_837,N_750,N_753);
nand U838 (N_838,N_750,N_779);
nand U839 (N_839,N_767,N_762);
nor U840 (N_840,N_758,N_761);
and U841 (N_841,N_785,N_798);
nor U842 (N_842,N_768,N_773);
nand U843 (N_843,N_791,N_762);
and U844 (N_844,N_779,N_796);
nand U845 (N_845,N_790,N_765);
or U846 (N_846,N_774,N_750);
or U847 (N_847,N_798,N_756);
nor U848 (N_848,N_753,N_793);
nor U849 (N_849,N_750,N_775);
and U850 (N_850,N_815,N_843);
nor U851 (N_851,N_822,N_825);
nor U852 (N_852,N_820,N_838);
nand U853 (N_853,N_845,N_821);
nand U854 (N_854,N_806,N_816);
and U855 (N_855,N_846,N_830);
and U856 (N_856,N_805,N_802);
nand U857 (N_857,N_827,N_812);
and U858 (N_858,N_814,N_823);
nand U859 (N_859,N_847,N_834);
nor U860 (N_860,N_835,N_844);
or U861 (N_861,N_809,N_841);
or U862 (N_862,N_819,N_828);
nor U863 (N_863,N_817,N_833);
xor U864 (N_864,N_829,N_832);
nand U865 (N_865,N_840,N_803);
nand U866 (N_866,N_849,N_842);
or U867 (N_867,N_810,N_808);
nand U868 (N_868,N_848,N_807);
and U869 (N_869,N_839,N_800);
nor U870 (N_870,N_813,N_811);
nor U871 (N_871,N_824,N_818);
and U872 (N_872,N_804,N_831);
nor U873 (N_873,N_801,N_826);
nor U874 (N_874,N_836,N_837);
and U875 (N_875,N_841,N_813);
nor U876 (N_876,N_830,N_820);
nor U877 (N_877,N_830,N_814);
and U878 (N_878,N_834,N_801);
nand U879 (N_879,N_848,N_846);
nand U880 (N_880,N_808,N_802);
nand U881 (N_881,N_817,N_803);
or U882 (N_882,N_805,N_823);
and U883 (N_883,N_831,N_823);
xor U884 (N_884,N_805,N_812);
or U885 (N_885,N_814,N_833);
nor U886 (N_886,N_809,N_840);
or U887 (N_887,N_801,N_815);
nor U888 (N_888,N_845,N_840);
nand U889 (N_889,N_810,N_835);
and U890 (N_890,N_835,N_842);
nand U891 (N_891,N_802,N_842);
and U892 (N_892,N_846,N_824);
nor U893 (N_893,N_806,N_835);
nor U894 (N_894,N_807,N_834);
nand U895 (N_895,N_845,N_831);
or U896 (N_896,N_825,N_836);
nand U897 (N_897,N_826,N_834);
nand U898 (N_898,N_816,N_800);
nand U899 (N_899,N_827,N_836);
nor U900 (N_900,N_858,N_889);
or U901 (N_901,N_899,N_859);
nand U902 (N_902,N_853,N_878);
and U903 (N_903,N_856,N_888);
and U904 (N_904,N_864,N_883);
nand U905 (N_905,N_880,N_896);
or U906 (N_906,N_894,N_857);
nand U907 (N_907,N_854,N_869);
or U908 (N_908,N_873,N_885);
or U909 (N_909,N_862,N_897);
or U910 (N_910,N_852,N_861);
nor U911 (N_911,N_850,N_868);
or U912 (N_912,N_874,N_890);
nor U913 (N_913,N_893,N_876);
or U914 (N_914,N_886,N_863);
nor U915 (N_915,N_877,N_875);
and U916 (N_916,N_866,N_882);
and U917 (N_917,N_851,N_871);
or U918 (N_918,N_867,N_865);
and U919 (N_919,N_872,N_887);
nand U920 (N_920,N_881,N_891);
nor U921 (N_921,N_879,N_892);
nand U922 (N_922,N_895,N_884);
or U923 (N_923,N_855,N_860);
and U924 (N_924,N_898,N_870);
or U925 (N_925,N_875,N_873);
nand U926 (N_926,N_898,N_881);
and U927 (N_927,N_888,N_892);
and U928 (N_928,N_883,N_897);
nor U929 (N_929,N_869,N_850);
or U930 (N_930,N_885,N_868);
nor U931 (N_931,N_888,N_863);
nor U932 (N_932,N_890,N_870);
nor U933 (N_933,N_857,N_870);
nor U934 (N_934,N_867,N_892);
or U935 (N_935,N_866,N_884);
nor U936 (N_936,N_879,N_867);
and U937 (N_937,N_862,N_866);
and U938 (N_938,N_880,N_856);
nand U939 (N_939,N_895,N_871);
and U940 (N_940,N_856,N_851);
or U941 (N_941,N_886,N_872);
nor U942 (N_942,N_889,N_855);
nor U943 (N_943,N_876,N_862);
nand U944 (N_944,N_898,N_877);
nand U945 (N_945,N_852,N_874);
nand U946 (N_946,N_883,N_865);
or U947 (N_947,N_870,N_855);
xor U948 (N_948,N_878,N_873);
or U949 (N_949,N_874,N_897);
or U950 (N_950,N_906,N_914);
nor U951 (N_951,N_947,N_937);
or U952 (N_952,N_917,N_948);
and U953 (N_953,N_929,N_938);
nand U954 (N_954,N_936,N_905);
and U955 (N_955,N_904,N_918);
nand U956 (N_956,N_933,N_923);
nor U957 (N_957,N_927,N_940);
or U958 (N_958,N_907,N_949);
or U959 (N_959,N_900,N_915);
or U960 (N_960,N_925,N_943);
nor U961 (N_961,N_916,N_922);
nor U962 (N_962,N_912,N_930);
nor U963 (N_963,N_913,N_931);
and U964 (N_964,N_908,N_911);
or U965 (N_965,N_902,N_910);
or U966 (N_966,N_920,N_901);
nor U967 (N_967,N_939,N_921);
and U968 (N_968,N_926,N_909);
nand U969 (N_969,N_934,N_903);
and U970 (N_970,N_945,N_941);
or U971 (N_971,N_935,N_946);
nor U972 (N_972,N_924,N_942);
nor U973 (N_973,N_944,N_919);
and U974 (N_974,N_928,N_932);
nor U975 (N_975,N_917,N_907);
nand U976 (N_976,N_908,N_913);
and U977 (N_977,N_900,N_922);
nor U978 (N_978,N_927,N_942);
nand U979 (N_979,N_945,N_936);
and U980 (N_980,N_910,N_949);
nand U981 (N_981,N_931,N_928);
and U982 (N_982,N_910,N_938);
nor U983 (N_983,N_945,N_906);
and U984 (N_984,N_925,N_929);
or U985 (N_985,N_941,N_906);
nand U986 (N_986,N_938,N_907);
nand U987 (N_987,N_927,N_909);
and U988 (N_988,N_920,N_908);
and U989 (N_989,N_941,N_910);
and U990 (N_990,N_928,N_912);
or U991 (N_991,N_932,N_924);
and U992 (N_992,N_924,N_943);
nand U993 (N_993,N_928,N_937);
nand U994 (N_994,N_946,N_908);
or U995 (N_995,N_924,N_919);
xor U996 (N_996,N_949,N_921);
xnor U997 (N_997,N_906,N_909);
or U998 (N_998,N_900,N_946);
or U999 (N_999,N_931,N_915);
or U1000 (N_1000,N_988,N_990);
nand U1001 (N_1001,N_964,N_957);
xor U1002 (N_1002,N_984,N_986);
and U1003 (N_1003,N_989,N_963);
nand U1004 (N_1004,N_959,N_956);
or U1005 (N_1005,N_974,N_967);
nor U1006 (N_1006,N_998,N_965);
nor U1007 (N_1007,N_979,N_977);
nand U1008 (N_1008,N_985,N_970);
and U1009 (N_1009,N_958,N_973);
and U1010 (N_1010,N_991,N_975);
or U1011 (N_1011,N_968,N_987);
and U1012 (N_1012,N_999,N_952);
and U1013 (N_1013,N_971,N_962);
nand U1014 (N_1014,N_966,N_954);
nand U1015 (N_1015,N_955,N_981);
nand U1016 (N_1016,N_982,N_992);
nor U1017 (N_1017,N_951,N_972);
nand U1018 (N_1018,N_961,N_983);
nand U1019 (N_1019,N_976,N_993);
or U1020 (N_1020,N_950,N_994);
and U1021 (N_1021,N_978,N_995);
or U1022 (N_1022,N_960,N_996);
nor U1023 (N_1023,N_997,N_969);
nor U1024 (N_1024,N_953,N_980);
nand U1025 (N_1025,N_967,N_990);
nor U1026 (N_1026,N_958,N_990);
and U1027 (N_1027,N_988,N_957);
nand U1028 (N_1028,N_953,N_983);
nor U1029 (N_1029,N_962,N_992);
or U1030 (N_1030,N_959,N_963);
or U1031 (N_1031,N_991,N_974);
nor U1032 (N_1032,N_984,N_985);
nor U1033 (N_1033,N_994,N_998);
nand U1034 (N_1034,N_987,N_988);
or U1035 (N_1035,N_989,N_988);
and U1036 (N_1036,N_957,N_950);
and U1037 (N_1037,N_970,N_998);
nand U1038 (N_1038,N_983,N_992);
nor U1039 (N_1039,N_987,N_976);
xnor U1040 (N_1040,N_979,N_992);
nor U1041 (N_1041,N_964,N_972);
or U1042 (N_1042,N_999,N_964);
and U1043 (N_1043,N_988,N_952);
nor U1044 (N_1044,N_985,N_973);
nor U1045 (N_1045,N_955,N_973);
nand U1046 (N_1046,N_974,N_955);
and U1047 (N_1047,N_951,N_997);
and U1048 (N_1048,N_973,N_981);
or U1049 (N_1049,N_989,N_986);
and U1050 (N_1050,N_1015,N_1025);
nor U1051 (N_1051,N_1048,N_1024);
and U1052 (N_1052,N_1021,N_1022);
and U1053 (N_1053,N_1010,N_1029);
nand U1054 (N_1054,N_1035,N_1003);
and U1055 (N_1055,N_1020,N_1028);
nand U1056 (N_1056,N_1018,N_1039);
nor U1057 (N_1057,N_1001,N_1049);
or U1058 (N_1058,N_1002,N_1006);
and U1059 (N_1059,N_1043,N_1016);
and U1060 (N_1060,N_1026,N_1044);
nor U1061 (N_1061,N_1037,N_1013);
nor U1062 (N_1062,N_1040,N_1005);
nand U1063 (N_1063,N_1007,N_1027);
and U1064 (N_1064,N_1000,N_1012);
and U1065 (N_1065,N_1047,N_1046);
and U1066 (N_1066,N_1038,N_1036);
or U1067 (N_1067,N_1042,N_1023);
nand U1068 (N_1068,N_1014,N_1033);
nor U1069 (N_1069,N_1030,N_1031);
nand U1070 (N_1070,N_1041,N_1008);
and U1071 (N_1071,N_1009,N_1019);
nand U1072 (N_1072,N_1034,N_1045);
and U1073 (N_1073,N_1032,N_1004);
and U1074 (N_1074,N_1011,N_1017);
nor U1075 (N_1075,N_1014,N_1005);
and U1076 (N_1076,N_1017,N_1039);
nand U1077 (N_1077,N_1003,N_1010);
nor U1078 (N_1078,N_1023,N_1006);
or U1079 (N_1079,N_1005,N_1000);
nand U1080 (N_1080,N_1007,N_1010);
nand U1081 (N_1081,N_1010,N_1042);
or U1082 (N_1082,N_1015,N_1024);
nand U1083 (N_1083,N_1039,N_1025);
nor U1084 (N_1084,N_1016,N_1039);
nor U1085 (N_1085,N_1026,N_1024);
nand U1086 (N_1086,N_1000,N_1046);
and U1087 (N_1087,N_1012,N_1011);
and U1088 (N_1088,N_1020,N_1047);
nor U1089 (N_1089,N_1002,N_1010);
nor U1090 (N_1090,N_1013,N_1040);
nand U1091 (N_1091,N_1028,N_1045);
nand U1092 (N_1092,N_1003,N_1021);
or U1093 (N_1093,N_1039,N_1043);
nor U1094 (N_1094,N_1010,N_1043);
and U1095 (N_1095,N_1013,N_1045);
and U1096 (N_1096,N_1008,N_1020);
or U1097 (N_1097,N_1040,N_1032);
nor U1098 (N_1098,N_1040,N_1044);
or U1099 (N_1099,N_1044,N_1027);
nor U1100 (N_1100,N_1086,N_1075);
or U1101 (N_1101,N_1052,N_1054);
nand U1102 (N_1102,N_1062,N_1092);
or U1103 (N_1103,N_1067,N_1071);
and U1104 (N_1104,N_1091,N_1056);
or U1105 (N_1105,N_1082,N_1080);
or U1106 (N_1106,N_1063,N_1065);
xnor U1107 (N_1107,N_1051,N_1098);
nand U1108 (N_1108,N_1087,N_1070);
or U1109 (N_1109,N_1069,N_1068);
nor U1110 (N_1110,N_1057,N_1058);
or U1111 (N_1111,N_1061,N_1055);
or U1112 (N_1112,N_1078,N_1060);
nor U1113 (N_1113,N_1084,N_1094);
nor U1114 (N_1114,N_1081,N_1083);
and U1115 (N_1115,N_1066,N_1072);
and U1116 (N_1116,N_1095,N_1090);
nand U1117 (N_1117,N_1096,N_1059);
nor U1118 (N_1118,N_1073,N_1079);
and U1119 (N_1119,N_1077,N_1085);
nand U1120 (N_1120,N_1097,N_1076);
or U1121 (N_1121,N_1053,N_1089);
nor U1122 (N_1122,N_1093,N_1099);
and U1123 (N_1123,N_1088,N_1064);
nand U1124 (N_1124,N_1050,N_1074);
nand U1125 (N_1125,N_1057,N_1052);
and U1126 (N_1126,N_1068,N_1098);
or U1127 (N_1127,N_1052,N_1090);
nor U1128 (N_1128,N_1098,N_1074);
or U1129 (N_1129,N_1097,N_1068);
and U1130 (N_1130,N_1095,N_1070);
and U1131 (N_1131,N_1090,N_1050);
and U1132 (N_1132,N_1067,N_1054);
and U1133 (N_1133,N_1066,N_1083);
and U1134 (N_1134,N_1066,N_1050);
nand U1135 (N_1135,N_1097,N_1061);
nor U1136 (N_1136,N_1051,N_1055);
nor U1137 (N_1137,N_1056,N_1096);
nor U1138 (N_1138,N_1091,N_1093);
nand U1139 (N_1139,N_1050,N_1095);
and U1140 (N_1140,N_1075,N_1066);
nand U1141 (N_1141,N_1067,N_1062);
or U1142 (N_1142,N_1087,N_1088);
or U1143 (N_1143,N_1062,N_1099);
or U1144 (N_1144,N_1070,N_1098);
or U1145 (N_1145,N_1083,N_1091);
or U1146 (N_1146,N_1085,N_1096);
xor U1147 (N_1147,N_1084,N_1074);
nand U1148 (N_1148,N_1084,N_1072);
or U1149 (N_1149,N_1072,N_1094);
and U1150 (N_1150,N_1129,N_1105);
nand U1151 (N_1151,N_1111,N_1106);
nand U1152 (N_1152,N_1133,N_1145);
or U1153 (N_1153,N_1148,N_1144);
and U1154 (N_1154,N_1127,N_1119);
or U1155 (N_1155,N_1121,N_1120);
or U1156 (N_1156,N_1116,N_1122);
nand U1157 (N_1157,N_1143,N_1114);
and U1158 (N_1158,N_1126,N_1100);
and U1159 (N_1159,N_1123,N_1146);
nand U1160 (N_1160,N_1142,N_1103);
nand U1161 (N_1161,N_1130,N_1113);
or U1162 (N_1162,N_1118,N_1147);
or U1163 (N_1163,N_1128,N_1140);
and U1164 (N_1164,N_1102,N_1135);
or U1165 (N_1165,N_1104,N_1125);
nor U1166 (N_1166,N_1134,N_1136);
nand U1167 (N_1167,N_1112,N_1108);
and U1168 (N_1168,N_1137,N_1149);
nor U1169 (N_1169,N_1141,N_1132);
or U1170 (N_1170,N_1138,N_1109);
or U1171 (N_1171,N_1115,N_1107);
nor U1172 (N_1172,N_1101,N_1139);
nor U1173 (N_1173,N_1110,N_1124);
nand U1174 (N_1174,N_1117,N_1131);
or U1175 (N_1175,N_1134,N_1141);
nand U1176 (N_1176,N_1125,N_1143);
nor U1177 (N_1177,N_1103,N_1114);
or U1178 (N_1178,N_1127,N_1137);
nor U1179 (N_1179,N_1128,N_1145);
and U1180 (N_1180,N_1111,N_1146);
and U1181 (N_1181,N_1100,N_1145);
nand U1182 (N_1182,N_1144,N_1120);
nand U1183 (N_1183,N_1144,N_1147);
nand U1184 (N_1184,N_1124,N_1130);
nand U1185 (N_1185,N_1140,N_1109);
nor U1186 (N_1186,N_1121,N_1149);
nand U1187 (N_1187,N_1146,N_1136);
nand U1188 (N_1188,N_1145,N_1131);
nand U1189 (N_1189,N_1111,N_1128);
nor U1190 (N_1190,N_1130,N_1134);
nand U1191 (N_1191,N_1118,N_1135);
nor U1192 (N_1192,N_1103,N_1143);
or U1193 (N_1193,N_1112,N_1138);
and U1194 (N_1194,N_1140,N_1142);
or U1195 (N_1195,N_1143,N_1111);
or U1196 (N_1196,N_1107,N_1100);
nand U1197 (N_1197,N_1149,N_1113);
nand U1198 (N_1198,N_1114,N_1122);
nand U1199 (N_1199,N_1131,N_1136);
or U1200 (N_1200,N_1185,N_1196);
nand U1201 (N_1201,N_1152,N_1162);
and U1202 (N_1202,N_1169,N_1157);
nor U1203 (N_1203,N_1164,N_1182);
and U1204 (N_1204,N_1153,N_1188);
and U1205 (N_1205,N_1179,N_1150);
nand U1206 (N_1206,N_1161,N_1194);
nand U1207 (N_1207,N_1176,N_1174);
nor U1208 (N_1208,N_1186,N_1191);
xnor U1209 (N_1209,N_1158,N_1197);
or U1210 (N_1210,N_1178,N_1171);
nand U1211 (N_1211,N_1154,N_1172);
or U1212 (N_1212,N_1167,N_1184);
nand U1213 (N_1213,N_1151,N_1180);
or U1214 (N_1214,N_1155,N_1166);
nand U1215 (N_1215,N_1159,N_1160);
or U1216 (N_1216,N_1156,N_1181);
and U1217 (N_1217,N_1189,N_1190);
nand U1218 (N_1218,N_1199,N_1193);
nor U1219 (N_1219,N_1183,N_1173);
nand U1220 (N_1220,N_1177,N_1168);
and U1221 (N_1221,N_1165,N_1192);
or U1222 (N_1222,N_1187,N_1198);
or U1223 (N_1223,N_1170,N_1195);
nor U1224 (N_1224,N_1163,N_1175);
nand U1225 (N_1225,N_1159,N_1179);
xor U1226 (N_1226,N_1165,N_1182);
or U1227 (N_1227,N_1156,N_1173);
nand U1228 (N_1228,N_1185,N_1178);
and U1229 (N_1229,N_1180,N_1198);
or U1230 (N_1230,N_1182,N_1168);
and U1231 (N_1231,N_1191,N_1172);
nor U1232 (N_1232,N_1190,N_1159);
or U1233 (N_1233,N_1195,N_1190);
nand U1234 (N_1234,N_1198,N_1194);
nand U1235 (N_1235,N_1195,N_1153);
nor U1236 (N_1236,N_1150,N_1190);
nor U1237 (N_1237,N_1166,N_1163);
and U1238 (N_1238,N_1192,N_1155);
or U1239 (N_1239,N_1199,N_1173);
nor U1240 (N_1240,N_1151,N_1153);
or U1241 (N_1241,N_1181,N_1199);
or U1242 (N_1242,N_1182,N_1151);
nor U1243 (N_1243,N_1159,N_1175);
or U1244 (N_1244,N_1162,N_1177);
or U1245 (N_1245,N_1160,N_1157);
nand U1246 (N_1246,N_1164,N_1197);
nand U1247 (N_1247,N_1172,N_1165);
nand U1248 (N_1248,N_1162,N_1161);
nor U1249 (N_1249,N_1177,N_1164);
nand U1250 (N_1250,N_1233,N_1248);
or U1251 (N_1251,N_1217,N_1214);
or U1252 (N_1252,N_1230,N_1204);
and U1253 (N_1253,N_1234,N_1211);
and U1254 (N_1254,N_1235,N_1240);
and U1255 (N_1255,N_1249,N_1244);
and U1256 (N_1256,N_1247,N_1208);
or U1257 (N_1257,N_1232,N_1219);
nand U1258 (N_1258,N_1205,N_1216);
xor U1259 (N_1259,N_1207,N_1202);
or U1260 (N_1260,N_1209,N_1226);
nand U1261 (N_1261,N_1243,N_1223);
nor U1262 (N_1262,N_1245,N_1222);
and U1263 (N_1263,N_1237,N_1227);
nand U1264 (N_1264,N_1242,N_1224);
and U1265 (N_1265,N_1238,N_1220);
or U1266 (N_1266,N_1228,N_1221);
or U1267 (N_1267,N_1201,N_1229);
nor U1268 (N_1268,N_1206,N_1225);
and U1269 (N_1269,N_1239,N_1215);
and U1270 (N_1270,N_1210,N_1218);
nand U1271 (N_1271,N_1241,N_1203);
or U1272 (N_1272,N_1200,N_1213);
or U1273 (N_1273,N_1236,N_1231);
nor U1274 (N_1274,N_1246,N_1212);
or U1275 (N_1275,N_1246,N_1217);
or U1276 (N_1276,N_1232,N_1248);
nand U1277 (N_1277,N_1237,N_1210);
and U1278 (N_1278,N_1210,N_1214);
nor U1279 (N_1279,N_1227,N_1244);
or U1280 (N_1280,N_1231,N_1225);
nand U1281 (N_1281,N_1240,N_1247);
or U1282 (N_1282,N_1218,N_1237);
nor U1283 (N_1283,N_1245,N_1238);
nand U1284 (N_1284,N_1245,N_1215);
and U1285 (N_1285,N_1231,N_1229);
or U1286 (N_1286,N_1240,N_1220);
or U1287 (N_1287,N_1245,N_1237);
and U1288 (N_1288,N_1232,N_1223);
nand U1289 (N_1289,N_1239,N_1230);
nand U1290 (N_1290,N_1209,N_1243);
nand U1291 (N_1291,N_1235,N_1248);
and U1292 (N_1292,N_1211,N_1212);
and U1293 (N_1293,N_1229,N_1247);
nor U1294 (N_1294,N_1200,N_1230);
or U1295 (N_1295,N_1224,N_1221);
nand U1296 (N_1296,N_1216,N_1238);
and U1297 (N_1297,N_1214,N_1241);
nand U1298 (N_1298,N_1212,N_1201);
nor U1299 (N_1299,N_1235,N_1232);
nand U1300 (N_1300,N_1285,N_1293);
nand U1301 (N_1301,N_1299,N_1251);
nand U1302 (N_1302,N_1264,N_1257);
nor U1303 (N_1303,N_1271,N_1291);
nor U1304 (N_1304,N_1282,N_1269);
and U1305 (N_1305,N_1272,N_1277);
nor U1306 (N_1306,N_1295,N_1276);
nand U1307 (N_1307,N_1294,N_1266);
or U1308 (N_1308,N_1259,N_1260);
nand U1309 (N_1309,N_1270,N_1278);
or U1310 (N_1310,N_1280,N_1275);
nand U1311 (N_1311,N_1298,N_1267);
or U1312 (N_1312,N_1292,N_1273);
and U1313 (N_1313,N_1265,N_1252);
nor U1314 (N_1314,N_1279,N_1262);
nor U1315 (N_1315,N_1261,N_1290);
nor U1316 (N_1316,N_1268,N_1254);
or U1317 (N_1317,N_1256,N_1263);
and U1318 (N_1318,N_1283,N_1281);
nor U1319 (N_1319,N_1255,N_1288);
nand U1320 (N_1320,N_1289,N_1286);
nor U1321 (N_1321,N_1274,N_1253);
nand U1322 (N_1322,N_1250,N_1258);
and U1323 (N_1323,N_1297,N_1287);
nor U1324 (N_1324,N_1284,N_1296);
nor U1325 (N_1325,N_1282,N_1265);
or U1326 (N_1326,N_1277,N_1298);
and U1327 (N_1327,N_1289,N_1270);
nand U1328 (N_1328,N_1283,N_1258);
or U1329 (N_1329,N_1272,N_1254);
and U1330 (N_1330,N_1266,N_1291);
xnor U1331 (N_1331,N_1289,N_1276);
and U1332 (N_1332,N_1253,N_1252);
and U1333 (N_1333,N_1264,N_1299);
or U1334 (N_1334,N_1278,N_1299);
and U1335 (N_1335,N_1288,N_1280);
and U1336 (N_1336,N_1283,N_1279);
and U1337 (N_1337,N_1265,N_1285);
and U1338 (N_1338,N_1280,N_1256);
and U1339 (N_1339,N_1263,N_1251);
nand U1340 (N_1340,N_1263,N_1270);
nor U1341 (N_1341,N_1260,N_1265);
nand U1342 (N_1342,N_1261,N_1286);
or U1343 (N_1343,N_1298,N_1258);
nand U1344 (N_1344,N_1286,N_1267);
nand U1345 (N_1345,N_1262,N_1277);
nand U1346 (N_1346,N_1252,N_1279);
nand U1347 (N_1347,N_1298,N_1260);
or U1348 (N_1348,N_1296,N_1279);
or U1349 (N_1349,N_1279,N_1275);
nor U1350 (N_1350,N_1349,N_1310);
nor U1351 (N_1351,N_1308,N_1335);
nor U1352 (N_1352,N_1322,N_1309);
and U1353 (N_1353,N_1342,N_1338);
nor U1354 (N_1354,N_1307,N_1313);
xnor U1355 (N_1355,N_1301,N_1325);
nand U1356 (N_1356,N_1332,N_1334);
nor U1357 (N_1357,N_1343,N_1318);
or U1358 (N_1358,N_1321,N_1336);
nand U1359 (N_1359,N_1320,N_1319);
nand U1360 (N_1360,N_1348,N_1303);
and U1361 (N_1361,N_1327,N_1306);
or U1362 (N_1362,N_1315,N_1302);
nor U1363 (N_1363,N_1333,N_1314);
or U1364 (N_1364,N_1331,N_1304);
or U1365 (N_1365,N_1323,N_1316);
nor U1366 (N_1366,N_1326,N_1345);
nand U1367 (N_1367,N_1347,N_1312);
and U1368 (N_1368,N_1330,N_1328);
nor U1369 (N_1369,N_1329,N_1344);
xor U1370 (N_1370,N_1346,N_1341);
or U1371 (N_1371,N_1337,N_1339);
or U1372 (N_1372,N_1317,N_1340);
nor U1373 (N_1373,N_1305,N_1311);
nand U1374 (N_1374,N_1300,N_1324);
or U1375 (N_1375,N_1326,N_1304);
and U1376 (N_1376,N_1326,N_1314);
nor U1377 (N_1377,N_1308,N_1331);
and U1378 (N_1378,N_1343,N_1306);
nor U1379 (N_1379,N_1327,N_1337);
or U1380 (N_1380,N_1306,N_1328);
nand U1381 (N_1381,N_1339,N_1326);
and U1382 (N_1382,N_1341,N_1342);
or U1383 (N_1383,N_1316,N_1336);
nand U1384 (N_1384,N_1333,N_1301);
and U1385 (N_1385,N_1321,N_1338);
xor U1386 (N_1386,N_1317,N_1318);
and U1387 (N_1387,N_1304,N_1311);
or U1388 (N_1388,N_1348,N_1302);
or U1389 (N_1389,N_1317,N_1319);
and U1390 (N_1390,N_1314,N_1312);
nor U1391 (N_1391,N_1326,N_1324);
or U1392 (N_1392,N_1340,N_1337);
nand U1393 (N_1393,N_1316,N_1338);
nor U1394 (N_1394,N_1330,N_1304);
nor U1395 (N_1395,N_1337,N_1338);
nand U1396 (N_1396,N_1323,N_1337);
nand U1397 (N_1397,N_1303,N_1304);
and U1398 (N_1398,N_1327,N_1333);
and U1399 (N_1399,N_1311,N_1333);
nor U1400 (N_1400,N_1373,N_1376);
nor U1401 (N_1401,N_1367,N_1390);
nand U1402 (N_1402,N_1387,N_1398);
nor U1403 (N_1403,N_1375,N_1385);
and U1404 (N_1404,N_1353,N_1379);
nor U1405 (N_1405,N_1358,N_1388);
nand U1406 (N_1406,N_1364,N_1363);
nand U1407 (N_1407,N_1391,N_1356);
nand U1408 (N_1408,N_1351,N_1378);
nand U1409 (N_1409,N_1381,N_1359);
and U1410 (N_1410,N_1350,N_1377);
or U1411 (N_1411,N_1395,N_1372);
or U1412 (N_1412,N_1368,N_1361);
nand U1413 (N_1413,N_1374,N_1386);
or U1414 (N_1414,N_1383,N_1389);
nand U1415 (N_1415,N_1384,N_1392);
nor U1416 (N_1416,N_1393,N_1366);
nand U1417 (N_1417,N_1380,N_1354);
and U1418 (N_1418,N_1357,N_1370);
nand U1419 (N_1419,N_1355,N_1399);
and U1420 (N_1420,N_1382,N_1360);
nand U1421 (N_1421,N_1396,N_1369);
or U1422 (N_1422,N_1371,N_1352);
or U1423 (N_1423,N_1362,N_1397);
and U1424 (N_1424,N_1394,N_1365);
and U1425 (N_1425,N_1366,N_1389);
nor U1426 (N_1426,N_1392,N_1364);
or U1427 (N_1427,N_1354,N_1375);
nor U1428 (N_1428,N_1396,N_1373);
and U1429 (N_1429,N_1366,N_1364);
and U1430 (N_1430,N_1370,N_1383);
and U1431 (N_1431,N_1369,N_1357);
nand U1432 (N_1432,N_1375,N_1396);
and U1433 (N_1433,N_1379,N_1355);
nor U1434 (N_1434,N_1397,N_1354);
and U1435 (N_1435,N_1355,N_1378);
nor U1436 (N_1436,N_1364,N_1379);
or U1437 (N_1437,N_1392,N_1367);
nor U1438 (N_1438,N_1371,N_1386);
nor U1439 (N_1439,N_1350,N_1385);
nor U1440 (N_1440,N_1381,N_1391);
and U1441 (N_1441,N_1362,N_1363);
nand U1442 (N_1442,N_1396,N_1383);
and U1443 (N_1443,N_1364,N_1372);
and U1444 (N_1444,N_1360,N_1361);
or U1445 (N_1445,N_1392,N_1385);
or U1446 (N_1446,N_1373,N_1393);
nand U1447 (N_1447,N_1354,N_1396);
and U1448 (N_1448,N_1372,N_1369);
nand U1449 (N_1449,N_1357,N_1362);
nor U1450 (N_1450,N_1422,N_1449);
and U1451 (N_1451,N_1436,N_1438);
or U1452 (N_1452,N_1434,N_1401);
nand U1453 (N_1453,N_1410,N_1447);
nor U1454 (N_1454,N_1417,N_1423);
or U1455 (N_1455,N_1427,N_1412);
nor U1456 (N_1456,N_1441,N_1424);
nand U1457 (N_1457,N_1408,N_1419);
or U1458 (N_1458,N_1407,N_1435);
nand U1459 (N_1459,N_1414,N_1444);
nand U1460 (N_1460,N_1405,N_1411);
and U1461 (N_1461,N_1409,N_1426);
nor U1462 (N_1462,N_1430,N_1442);
nand U1463 (N_1463,N_1448,N_1432);
and U1464 (N_1464,N_1406,N_1431);
and U1465 (N_1465,N_1429,N_1416);
nand U1466 (N_1466,N_1446,N_1437);
and U1467 (N_1467,N_1400,N_1413);
or U1468 (N_1468,N_1428,N_1445);
nor U1469 (N_1469,N_1402,N_1425);
nand U1470 (N_1470,N_1433,N_1403);
nor U1471 (N_1471,N_1439,N_1420);
nand U1472 (N_1472,N_1418,N_1443);
nor U1473 (N_1473,N_1440,N_1404);
or U1474 (N_1474,N_1421,N_1415);
or U1475 (N_1475,N_1405,N_1449);
nor U1476 (N_1476,N_1405,N_1427);
nand U1477 (N_1477,N_1405,N_1413);
and U1478 (N_1478,N_1449,N_1410);
or U1479 (N_1479,N_1437,N_1425);
or U1480 (N_1480,N_1430,N_1410);
nor U1481 (N_1481,N_1415,N_1411);
nor U1482 (N_1482,N_1414,N_1439);
and U1483 (N_1483,N_1401,N_1405);
nor U1484 (N_1484,N_1437,N_1415);
and U1485 (N_1485,N_1422,N_1413);
or U1486 (N_1486,N_1431,N_1447);
nor U1487 (N_1487,N_1424,N_1410);
nand U1488 (N_1488,N_1410,N_1437);
nor U1489 (N_1489,N_1439,N_1426);
or U1490 (N_1490,N_1415,N_1414);
nand U1491 (N_1491,N_1447,N_1401);
or U1492 (N_1492,N_1434,N_1446);
nor U1493 (N_1493,N_1425,N_1415);
or U1494 (N_1494,N_1412,N_1447);
nand U1495 (N_1495,N_1413,N_1447);
nor U1496 (N_1496,N_1436,N_1400);
or U1497 (N_1497,N_1441,N_1402);
nand U1498 (N_1498,N_1404,N_1422);
nand U1499 (N_1499,N_1415,N_1417);
and U1500 (N_1500,N_1499,N_1498);
or U1501 (N_1501,N_1490,N_1492);
nand U1502 (N_1502,N_1484,N_1486);
and U1503 (N_1503,N_1464,N_1485);
or U1504 (N_1504,N_1489,N_1470);
nand U1505 (N_1505,N_1471,N_1475);
or U1506 (N_1506,N_1497,N_1481);
nand U1507 (N_1507,N_1460,N_1474);
nand U1508 (N_1508,N_1494,N_1451);
or U1509 (N_1509,N_1461,N_1467);
or U1510 (N_1510,N_1473,N_1472);
nor U1511 (N_1511,N_1465,N_1479);
nor U1512 (N_1512,N_1478,N_1482);
or U1513 (N_1513,N_1456,N_1458);
nor U1514 (N_1514,N_1457,N_1476);
or U1515 (N_1515,N_1462,N_1468);
nor U1516 (N_1516,N_1466,N_1483);
nor U1517 (N_1517,N_1455,N_1459);
and U1518 (N_1518,N_1495,N_1496);
and U1519 (N_1519,N_1488,N_1453);
or U1520 (N_1520,N_1450,N_1493);
nor U1521 (N_1521,N_1463,N_1454);
or U1522 (N_1522,N_1487,N_1469);
and U1523 (N_1523,N_1477,N_1452);
nand U1524 (N_1524,N_1491,N_1480);
nor U1525 (N_1525,N_1451,N_1484);
or U1526 (N_1526,N_1454,N_1480);
and U1527 (N_1527,N_1474,N_1457);
nor U1528 (N_1528,N_1486,N_1499);
or U1529 (N_1529,N_1471,N_1489);
nor U1530 (N_1530,N_1455,N_1456);
or U1531 (N_1531,N_1461,N_1488);
or U1532 (N_1532,N_1458,N_1489);
nand U1533 (N_1533,N_1490,N_1495);
or U1534 (N_1534,N_1475,N_1490);
or U1535 (N_1535,N_1475,N_1488);
and U1536 (N_1536,N_1497,N_1468);
nor U1537 (N_1537,N_1464,N_1492);
nand U1538 (N_1538,N_1450,N_1459);
and U1539 (N_1539,N_1490,N_1496);
nor U1540 (N_1540,N_1470,N_1450);
or U1541 (N_1541,N_1491,N_1476);
and U1542 (N_1542,N_1465,N_1492);
and U1543 (N_1543,N_1456,N_1486);
nand U1544 (N_1544,N_1494,N_1464);
nand U1545 (N_1545,N_1488,N_1468);
and U1546 (N_1546,N_1453,N_1459);
or U1547 (N_1547,N_1451,N_1486);
or U1548 (N_1548,N_1451,N_1463);
nand U1549 (N_1549,N_1475,N_1464);
nor U1550 (N_1550,N_1533,N_1523);
or U1551 (N_1551,N_1526,N_1543);
or U1552 (N_1552,N_1507,N_1501);
or U1553 (N_1553,N_1528,N_1500);
nand U1554 (N_1554,N_1545,N_1506);
and U1555 (N_1555,N_1535,N_1549);
nor U1556 (N_1556,N_1504,N_1532);
and U1557 (N_1557,N_1538,N_1503);
or U1558 (N_1558,N_1524,N_1505);
nor U1559 (N_1559,N_1512,N_1539);
or U1560 (N_1560,N_1540,N_1531);
or U1561 (N_1561,N_1521,N_1511);
or U1562 (N_1562,N_1547,N_1517);
and U1563 (N_1563,N_1548,N_1519);
nor U1564 (N_1564,N_1536,N_1520);
or U1565 (N_1565,N_1529,N_1546);
nand U1566 (N_1566,N_1541,N_1530);
and U1567 (N_1567,N_1522,N_1515);
nor U1568 (N_1568,N_1525,N_1513);
and U1569 (N_1569,N_1510,N_1514);
and U1570 (N_1570,N_1544,N_1508);
or U1571 (N_1571,N_1502,N_1509);
or U1572 (N_1572,N_1537,N_1516);
or U1573 (N_1573,N_1518,N_1542);
nor U1574 (N_1574,N_1534,N_1527);
nor U1575 (N_1575,N_1547,N_1533);
or U1576 (N_1576,N_1518,N_1508);
nand U1577 (N_1577,N_1542,N_1532);
nor U1578 (N_1578,N_1524,N_1529);
or U1579 (N_1579,N_1529,N_1531);
nor U1580 (N_1580,N_1507,N_1539);
nand U1581 (N_1581,N_1544,N_1515);
xnor U1582 (N_1582,N_1504,N_1508);
nor U1583 (N_1583,N_1523,N_1549);
and U1584 (N_1584,N_1503,N_1546);
nor U1585 (N_1585,N_1520,N_1502);
and U1586 (N_1586,N_1541,N_1503);
nor U1587 (N_1587,N_1524,N_1526);
nand U1588 (N_1588,N_1529,N_1528);
or U1589 (N_1589,N_1545,N_1532);
and U1590 (N_1590,N_1513,N_1522);
or U1591 (N_1591,N_1538,N_1501);
and U1592 (N_1592,N_1504,N_1517);
nor U1593 (N_1593,N_1511,N_1531);
and U1594 (N_1594,N_1524,N_1540);
nand U1595 (N_1595,N_1520,N_1549);
and U1596 (N_1596,N_1548,N_1516);
or U1597 (N_1597,N_1524,N_1528);
or U1598 (N_1598,N_1538,N_1547);
nor U1599 (N_1599,N_1504,N_1513);
nor U1600 (N_1600,N_1588,N_1562);
or U1601 (N_1601,N_1585,N_1576);
nand U1602 (N_1602,N_1582,N_1583);
and U1603 (N_1603,N_1569,N_1592);
nor U1604 (N_1604,N_1570,N_1553);
and U1605 (N_1605,N_1554,N_1577);
nor U1606 (N_1606,N_1552,N_1568);
and U1607 (N_1607,N_1561,N_1597);
and U1608 (N_1608,N_1580,N_1559);
and U1609 (N_1609,N_1573,N_1575);
nand U1610 (N_1610,N_1590,N_1578);
or U1611 (N_1611,N_1550,N_1584);
or U1612 (N_1612,N_1579,N_1564);
nand U1613 (N_1613,N_1567,N_1596);
nand U1614 (N_1614,N_1586,N_1574);
and U1615 (N_1615,N_1581,N_1556);
and U1616 (N_1616,N_1566,N_1555);
nand U1617 (N_1617,N_1551,N_1560);
or U1618 (N_1618,N_1593,N_1558);
or U1619 (N_1619,N_1565,N_1589);
nor U1620 (N_1620,N_1594,N_1599);
nor U1621 (N_1621,N_1571,N_1557);
or U1622 (N_1622,N_1595,N_1587);
nand U1623 (N_1623,N_1591,N_1572);
nor U1624 (N_1624,N_1598,N_1563);
and U1625 (N_1625,N_1599,N_1597);
nor U1626 (N_1626,N_1567,N_1593);
nor U1627 (N_1627,N_1572,N_1586);
and U1628 (N_1628,N_1591,N_1551);
nand U1629 (N_1629,N_1579,N_1560);
or U1630 (N_1630,N_1594,N_1590);
and U1631 (N_1631,N_1550,N_1598);
and U1632 (N_1632,N_1579,N_1567);
or U1633 (N_1633,N_1579,N_1583);
nor U1634 (N_1634,N_1563,N_1565);
and U1635 (N_1635,N_1585,N_1555);
nor U1636 (N_1636,N_1597,N_1594);
and U1637 (N_1637,N_1596,N_1588);
and U1638 (N_1638,N_1574,N_1570);
and U1639 (N_1639,N_1565,N_1577);
and U1640 (N_1640,N_1563,N_1580);
nand U1641 (N_1641,N_1578,N_1581);
nor U1642 (N_1642,N_1579,N_1557);
nand U1643 (N_1643,N_1586,N_1578);
nand U1644 (N_1644,N_1565,N_1559);
and U1645 (N_1645,N_1551,N_1598);
or U1646 (N_1646,N_1558,N_1595);
and U1647 (N_1647,N_1582,N_1567);
and U1648 (N_1648,N_1569,N_1561);
and U1649 (N_1649,N_1584,N_1561);
nor U1650 (N_1650,N_1633,N_1608);
or U1651 (N_1651,N_1641,N_1640);
and U1652 (N_1652,N_1616,N_1626);
or U1653 (N_1653,N_1622,N_1603);
or U1654 (N_1654,N_1630,N_1602);
or U1655 (N_1655,N_1607,N_1604);
or U1656 (N_1656,N_1637,N_1613);
nand U1657 (N_1657,N_1623,N_1644);
and U1658 (N_1658,N_1621,N_1612);
nor U1659 (N_1659,N_1624,N_1632);
or U1660 (N_1660,N_1625,N_1600);
or U1661 (N_1661,N_1649,N_1614);
nor U1662 (N_1662,N_1636,N_1618);
nor U1663 (N_1663,N_1642,N_1634);
nand U1664 (N_1664,N_1646,N_1615);
or U1665 (N_1665,N_1645,N_1610);
or U1666 (N_1666,N_1635,N_1647);
nor U1667 (N_1667,N_1648,N_1611);
or U1668 (N_1668,N_1643,N_1638);
nand U1669 (N_1669,N_1627,N_1628);
or U1670 (N_1670,N_1606,N_1605);
nor U1671 (N_1671,N_1629,N_1620);
nand U1672 (N_1672,N_1601,N_1631);
nand U1673 (N_1673,N_1639,N_1609);
nor U1674 (N_1674,N_1619,N_1617);
nand U1675 (N_1675,N_1633,N_1613);
or U1676 (N_1676,N_1621,N_1634);
and U1677 (N_1677,N_1632,N_1627);
nand U1678 (N_1678,N_1636,N_1644);
nand U1679 (N_1679,N_1605,N_1633);
nor U1680 (N_1680,N_1619,N_1637);
and U1681 (N_1681,N_1601,N_1633);
nor U1682 (N_1682,N_1634,N_1631);
nor U1683 (N_1683,N_1634,N_1627);
or U1684 (N_1684,N_1618,N_1627);
nor U1685 (N_1685,N_1616,N_1640);
nor U1686 (N_1686,N_1616,N_1647);
nor U1687 (N_1687,N_1628,N_1613);
and U1688 (N_1688,N_1638,N_1601);
and U1689 (N_1689,N_1640,N_1622);
nor U1690 (N_1690,N_1638,N_1625);
nor U1691 (N_1691,N_1606,N_1602);
and U1692 (N_1692,N_1638,N_1627);
nand U1693 (N_1693,N_1620,N_1613);
nor U1694 (N_1694,N_1632,N_1621);
or U1695 (N_1695,N_1636,N_1632);
and U1696 (N_1696,N_1630,N_1603);
nor U1697 (N_1697,N_1624,N_1639);
and U1698 (N_1698,N_1603,N_1609);
and U1699 (N_1699,N_1641,N_1634);
nand U1700 (N_1700,N_1662,N_1669);
nand U1701 (N_1701,N_1654,N_1691);
nand U1702 (N_1702,N_1693,N_1695);
and U1703 (N_1703,N_1684,N_1661);
and U1704 (N_1704,N_1671,N_1651);
nor U1705 (N_1705,N_1689,N_1698);
or U1706 (N_1706,N_1663,N_1688);
xnor U1707 (N_1707,N_1673,N_1699);
or U1708 (N_1708,N_1692,N_1694);
and U1709 (N_1709,N_1680,N_1679);
nand U1710 (N_1710,N_1667,N_1660);
nand U1711 (N_1711,N_1677,N_1681);
or U1712 (N_1712,N_1656,N_1653);
and U1713 (N_1713,N_1670,N_1672);
and U1714 (N_1714,N_1685,N_1686);
nand U1715 (N_1715,N_1665,N_1650);
or U1716 (N_1716,N_1682,N_1683);
or U1717 (N_1717,N_1657,N_1696);
nand U1718 (N_1718,N_1674,N_1659);
and U1719 (N_1719,N_1658,N_1668);
or U1720 (N_1720,N_1655,N_1666);
nor U1721 (N_1721,N_1687,N_1652);
nand U1722 (N_1722,N_1690,N_1664);
nand U1723 (N_1723,N_1678,N_1697);
nand U1724 (N_1724,N_1676,N_1675);
and U1725 (N_1725,N_1695,N_1666);
and U1726 (N_1726,N_1693,N_1654);
nor U1727 (N_1727,N_1678,N_1682);
and U1728 (N_1728,N_1699,N_1652);
and U1729 (N_1729,N_1666,N_1699);
nand U1730 (N_1730,N_1684,N_1652);
nand U1731 (N_1731,N_1688,N_1657);
nor U1732 (N_1732,N_1655,N_1681);
or U1733 (N_1733,N_1658,N_1662);
nor U1734 (N_1734,N_1690,N_1654);
nand U1735 (N_1735,N_1652,N_1679);
nand U1736 (N_1736,N_1699,N_1671);
or U1737 (N_1737,N_1655,N_1661);
nor U1738 (N_1738,N_1665,N_1664);
nor U1739 (N_1739,N_1691,N_1683);
nor U1740 (N_1740,N_1666,N_1665);
or U1741 (N_1741,N_1668,N_1698);
nor U1742 (N_1742,N_1657,N_1699);
nand U1743 (N_1743,N_1660,N_1650);
or U1744 (N_1744,N_1650,N_1669);
and U1745 (N_1745,N_1673,N_1670);
nor U1746 (N_1746,N_1689,N_1655);
nand U1747 (N_1747,N_1697,N_1684);
or U1748 (N_1748,N_1658,N_1691);
nor U1749 (N_1749,N_1697,N_1673);
nand U1750 (N_1750,N_1718,N_1737);
nor U1751 (N_1751,N_1713,N_1714);
or U1752 (N_1752,N_1743,N_1740);
and U1753 (N_1753,N_1730,N_1742);
and U1754 (N_1754,N_1736,N_1745);
nor U1755 (N_1755,N_1701,N_1712);
or U1756 (N_1756,N_1729,N_1725);
and U1757 (N_1757,N_1711,N_1722);
or U1758 (N_1758,N_1710,N_1744);
nor U1759 (N_1759,N_1706,N_1702);
and U1760 (N_1760,N_1731,N_1735);
or U1761 (N_1761,N_1732,N_1707);
nor U1762 (N_1762,N_1709,N_1720);
nor U1763 (N_1763,N_1717,N_1739);
and U1764 (N_1764,N_1719,N_1708);
and U1765 (N_1765,N_1746,N_1738);
or U1766 (N_1766,N_1726,N_1715);
or U1767 (N_1767,N_1741,N_1749);
and U1768 (N_1768,N_1716,N_1703);
or U1769 (N_1769,N_1721,N_1704);
or U1770 (N_1770,N_1727,N_1748);
and U1771 (N_1771,N_1724,N_1700);
and U1772 (N_1772,N_1723,N_1728);
nor U1773 (N_1773,N_1733,N_1747);
and U1774 (N_1774,N_1705,N_1734);
and U1775 (N_1775,N_1712,N_1731);
or U1776 (N_1776,N_1746,N_1724);
nand U1777 (N_1777,N_1712,N_1729);
nor U1778 (N_1778,N_1747,N_1704);
nand U1779 (N_1779,N_1705,N_1740);
nand U1780 (N_1780,N_1723,N_1722);
nor U1781 (N_1781,N_1718,N_1708);
nor U1782 (N_1782,N_1738,N_1708);
and U1783 (N_1783,N_1714,N_1735);
nand U1784 (N_1784,N_1712,N_1743);
or U1785 (N_1785,N_1723,N_1709);
or U1786 (N_1786,N_1738,N_1711);
nor U1787 (N_1787,N_1723,N_1718);
or U1788 (N_1788,N_1745,N_1715);
nand U1789 (N_1789,N_1722,N_1714);
or U1790 (N_1790,N_1746,N_1734);
xor U1791 (N_1791,N_1739,N_1724);
or U1792 (N_1792,N_1717,N_1705);
nor U1793 (N_1793,N_1725,N_1735);
or U1794 (N_1794,N_1711,N_1705);
nand U1795 (N_1795,N_1725,N_1709);
nor U1796 (N_1796,N_1723,N_1734);
nor U1797 (N_1797,N_1740,N_1720);
or U1798 (N_1798,N_1703,N_1710);
or U1799 (N_1799,N_1700,N_1718);
and U1800 (N_1800,N_1779,N_1766);
and U1801 (N_1801,N_1782,N_1758);
and U1802 (N_1802,N_1795,N_1762);
nor U1803 (N_1803,N_1776,N_1773);
xor U1804 (N_1804,N_1793,N_1757);
nor U1805 (N_1805,N_1786,N_1792);
and U1806 (N_1806,N_1780,N_1790);
nor U1807 (N_1807,N_1772,N_1775);
nand U1808 (N_1808,N_1783,N_1774);
and U1809 (N_1809,N_1785,N_1759);
or U1810 (N_1810,N_1768,N_1797);
nor U1811 (N_1811,N_1755,N_1799);
or U1812 (N_1812,N_1770,N_1751);
nor U1813 (N_1813,N_1760,N_1769);
nor U1814 (N_1814,N_1771,N_1752);
or U1815 (N_1815,N_1791,N_1794);
nor U1816 (N_1816,N_1789,N_1787);
or U1817 (N_1817,N_1763,N_1788);
or U1818 (N_1818,N_1756,N_1778);
nor U1819 (N_1819,N_1767,N_1798);
nor U1820 (N_1820,N_1764,N_1753);
or U1821 (N_1821,N_1765,N_1784);
or U1822 (N_1822,N_1777,N_1750);
nand U1823 (N_1823,N_1796,N_1781);
and U1824 (N_1824,N_1761,N_1754);
and U1825 (N_1825,N_1764,N_1785);
or U1826 (N_1826,N_1768,N_1759);
and U1827 (N_1827,N_1756,N_1751);
nor U1828 (N_1828,N_1796,N_1777);
nand U1829 (N_1829,N_1792,N_1773);
nor U1830 (N_1830,N_1794,N_1760);
nand U1831 (N_1831,N_1778,N_1760);
or U1832 (N_1832,N_1781,N_1782);
and U1833 (N_1833,N_1783,N_1771);
or U1834 (N_1834,N_1782,N_1773);
nor U1835 (N_1835,N_1771,N_1770);
and U1836 (N_1836,N_1767,N_1756);
nor U1837 (N_1837,N_1791,N_1779);
nand U1838 (N_1838,N_1795,N_1780);
and U1839 (N_1839,N_1790,N_1767);
nand U1840 (N_1840,N_1759,N_1787);
nor U1841 (N_1841,N_1776,N_1752);
nand U1842 (N_1842,N_1760,N_1795);
nand U1843 (N_1843,N_1785,N_1750);
nor U1844 (N_1844,N_1777,N_1778);
nor U1845 (N_1845,N_1791,N_1799);
and U1846 (N_1846,N_1766,N_1780);
and U1847 (N_1847,N_1793,N_1764);
nor U1848 (N_1848,N_1778,N_1795);
nor U1849 (N_1849,N_1766,N_1768);
nor U1850 (N_1850,N_1822,N_1827);
or U1851 (N_1851,N_1813,N_1846);
nor U1852 (N_1852,N_1800,N_1801);
nor U1853 (N_1853,N_1831,N_1804);
and U1854 (N_1854,N_1835,N_1820);
and U1855 (N_1855,N_1817,N_1834);
and U1856 (N_1856,N_1821,N_1805);
or U1857 (N_1857,N_1803,N_1837);
nor U1858 (N_1858,N_1814,N_1802);
nor U1859 (N_1859,N_1828,N_1807);
or U1860 (N_1860,N_1839,N_1824);
or U1861 (N_1861,N_1806,N_1840);
or U1862 (N_1862,N_1836,N_1842);
nor U1863 (N_1863,N_1808,N_1843);
nor U1864 (N_1864,N_1847,N_1810);
or U1865 (N_1865,N_1816,N_1845);
or U1866 (N_1866,N_1811,N_1826);
nor U1867 (N_1867,N_1841,N_1832);
and U1868 (N_1868,N_1849,N_1809);
or U1869 (N_1869,N_1812,N_1829);
and U1870 (N_1870,N_1830,N_1844);
and U1871 (N_1871,N_1818,N_1819);
nand U1872 (N_1872,N_1825,N_1815);
or U1873 (N_1873,N_1833,N_1838);
and U1874 (N_1874,N_1848,N_1823);
or U1875 (N_1875,N_1830,N_1804);
or U1876 (N_1876,N_1838,N_1828);
nor U1877 (N_1877,N_1819,N_1833);
nor U1878 (N_1878,N_1808,N_1832);
and U1879 (N_1879,N_1815,N_1826);
nand U1880 (N_1880,N_1809,N_1822);
nand U1881 (N_1881,N_1841,N_1848);
or U1882 (N_1882,N_1801,N_1849);
nand U1883 (N_1883,N_1822,N_1842);
nor U1884 (N_1884,N_1841,N_1843);
or U1885 (N_1885,N_1816,N_1800);
nand U1886 (N_1886,N_1845,N_1842);
or U1887 (N_1887,N_1821,N_1811);
or U1888 (N_1888,N_1833,N_1845);
nand U1889 (N_1889,N_1805,N_1803);
nand U1890 (N_1890,N_1821,N_1842);
and U1891 (N_1891,N_1847,N_1823);
or U1892 (N_1892,N_1830,N_1825);
nand U1893 (N_1893,N_1833,N_1800);
nor U1894 (N_1894,N_1814,N_1805);
and U1895 (N_1895,N_1808,N_1802);
or U1896 (N_1896,N_1809,N_1801);
nand U1897 (N_1897,N_1847,N_1814);
nand U1898 (N_1898,N_1831,N_1815);
and U1899 (N_1899,N_1825,N_1848);
or U1900 (N_1900,N_1865,N_1858);
nand U1901 (N_1901,N_1859,N_1890);
and U1902 (N_1902,N_1851,N_1878);
and U1903 (N_1903,N_1887,N_1892);
nor U1904 (N_1904,N_1864,N_1894);
and U1905 (N_1905,N_1885,N_1852);
nand U1906 (N_1906,N_1896,N_1895);
or U1907 (N_1907,N_1872,N_1875);
nand U1908 (N_1908,N_1862,N_1899);
or U1909 (N_1909,N_1877,N_1889);
nor U1910 (N_1910,N_1869,N_1870);
nand U1911 (N_1911,N_1854,N_1874);
or U1912 (N_1912,N_1886,N_1857);
nor U1913 (N_1913,N_1871,N_1850);
or U1914 (N_1914,N_1898,N_1855);
and U1915 (N_1915,N_1882,N_1873);
nor U1916 (N_1916,N_1891,N_1860);
or U1917 (N_1917,N_1868,N_1893);
nor U1918 (N_1918,N_1879,N_1856);
or U1919 (N_1919,N_1880,N_1863);
and U1920 (N_1920,N_1883,N_1881);
and U1921 (N_1921,N_1867,N_1853);
or U1922 (N_1922,N_1884,N_1897);
and U1923 (N_1923,N_1876,N_1866);
nor U1924 (N_1924,N_1861,N_1888);
and U1925 (N_1925,N_1894,N_1898);
nand U1926 (N_1926,N_1875,N_1879);
and U1927 (N_1927,N_1858,N_1856);
or U1928 (N_1928,N_1891,N_1854);
nand U1929 (N_1929,N_1897,N_1858);
or U1930 (N_1930,N_1880,N_1865);
nor U1931 (N_1931,N_1856,N_1881);
and U1932 (N_1932,N_1866,N_1893);
or U1933 (N_1933,N_1892,N_1878);
or U1934 (N_1934,N_1887,N_1888);
and U1935 (N_1935,N_1869,N_1857);
nand U1936 (N_1936,N_1889,N_1892);
or U1937 (N_1937,N_1866,N_1883);
nor U1938 (N_1938,N_1879,N_1862);
nand U1939 (N_1939,N_1855,N_1885);
nand U1940 (N_1940,N_1858,N_1877);
or U1941 (N_1941,N_1888,N_1860);
and U1942 (N_1942,N_1867,N_1898);
or U1943 (N_1943,N_1870,N_1876);
or U1944 (N_1944,N_1856,N_1867);
nor U1945 (N_1945,N_1893,N_1885);
nand U1946 (N_1946,N_1891,N_1857);
or U1947 (N_1947,N_1878,N_1886);
and U1948 (N_1948,N_1882,N_1859);
or U1949 (N_1949,N_1853,N_1882);
and U1950 (N_1950,N_1904,N_1902);
and U1951 (N_1951,N_1907,N_1936);
or U1952 (N_1952,N_1934,N_1924);
nor U1953 (N_1953,N_1921,N_1938);
or U1954 (N_1954,N_1911,N_1943);
and U1955 (N_1955,N_1917,N_1946);
or U1956 (N_1956,N_1926,N_1906);
and U1957 (N_1957,N_1920,N_1912);
and U1958 (N_1958,N_1923,N_1941);
nor U1959 (N_1959,N_1909,N_1929);
nor U1960 (N_1960,N_1915,N_1949);
nand U1961 (N_1961,N_1939,N_1948);
or U1962 (N_1962,N_1900,N_1908);
or U1963 (N_1963,N_1910,N_1942);
and U1964 (N_1964,N_1914,N_1922);
nand U1965 (N_1965,N_1940,N_1916);
and U1966 (N_1966,N_1931,N_1930);
nand U1967 (N_1967,N_1927,N_1905);
nor U1968 (N_1968,N_1932,N_1933);
and U1969 (N_1969,N_1903,N_1947);
and U1970 (N_1970,N_1944,N_1918);
nand U1971 (N_1971,N_1928,N_1937);
nor U1972 (N_1972,N_1919,N_1901);
nor U1973 (N_1973,N_1925,N_1945);
and U1974 (N_1974,N_1913,N_1935);
or U1975 (N_1975,N_1915,N_1919);
and U1976 (N_1976,N_1927,N_1944);
and U1977 (N_1977,N_1931,N_1901);
or U1978 (N_1978,N_1910,N_1936);
nor U1979 (N_1979,N_1917,N_1949);
nand U1980 (N_1980,N_1931,N_1916);
nor U1981 (N_1981,N_1939,N_1930);
and U1982 (N_1982,N_1939,N_1924);
nor U1983 (N_1983,N_1907,N_1900);
nor U1984 (N_1984,N_1949,N_1919);
or U1985 (N_1985,N_1915,N_1935);
nor U1986 (N_1986,N_1906,N_1907);
and U1987 (N_1987,N_1910,N_1903);
nand U1988 (N_1988,N_1931,N_1915);
and U1989 (N_1989,N_1924,N_1937);
or U1990 (N_1990,N_1901,N_1907);
or U1991 (N_1991,N_1918,N_1909);
nand U1992 (N_1992,N_1938,N_1931);
and U1993 (N_1993,N_1901,N_1941);
nor U1994 (N_1994,N_1912,N_1930);
and U1995 (N_1995,N_1913,N_1904);
nor U1996 (N_1996,N_1902,N_1935);
and U1997 (N_1997,N_1935,N_1942);
nand U1998 (N_1998,N_1943,N_1933);
nor U1999 (N_1999,N_1913,N_1934);
and U2000 (N_2000,N_1957,N_1958);
or U2001 (N_2001,N_1962,N_1982);
nand U2002 (N_2002,N_1968,N_1984);
and U2003 (N_2003,N_1983,N_1971);
or U2004 (N_2004,N_1975,N_1990);
nand U2005 (N_2005,N_1980,N_1954);
nor U2006 (N_2006,N_1974,N_1963);
and U2007 (N_2007,N_1977,N_1956);
nand U2008 (N_2008,N_1989,N_1964);
and U2009 (N_2009,N_1969,N_1951);
or U2010 (N_2010,N_1991,N_1961);
nand U2011 (N_2011,N_1978,N_1960);
or U2012 (N_2012,N_1999,N_1966);
or U2013 (N_2013,N_1970,N_1988);
or U2014 (N_2014,N_1997,N_1995);
or U2015 (N_2015,N_1996,N_1953);
and U2016 (N_2016,N_1998,N_1965);
nor U2017 (N_2017,N_1950,N_1986);
xnor U2018 (N_2018,N_1985,N_1993);
nor U2019 (N_2019,N_1981,N_1952);
nor U2020 (N_2020,N_1967,N_1987);
nor U2021 (N_2021,N_1973,N_1955);
and U2022 (N_2022,N_1972,N_1994);
and U2023 (N_2023,N_1959,N_1992);
nand U2024 (N_2024,N_1976,N_1979);
nand U2025 (N_2025,N_1997,N_1981);
nor U2026 (N_2026,N_1979,N_1987);
nand U2027 (N_2027,N_1992,N_1983);
or U2028 (N_2028,N_1954,N_1997);
and U2029 (N_2029,N_1985,N_1979);
nand U2030 (N_2030,N_1954,N_1999);
nand U2031 (N_2031,N_1993,N_1975);
nor U2032 (N_2032,N_1977,N_1974);
and U2033 (N_2033,N_1950,N_1974);
or U2034 (N_2034,N_1958,N_1968);
and U2035 (N_2035,N_1972,N_1986);
nor U2036 (N_2036,N_1977,N_1959);
and U2037 (N_2037,N_1986,N_1975);
nor U2038 (N_2038,N_1976,N_1950);
and U2039 (N_2039,N_1975,N_1970);
and U2040 (N_2040,N_1959,N_1966);
and U2041 (N_2041,N_1997,N_1975);
and U2042 (N_2042,N_1957,N_1952);
or U2043 (N_2043,N_1997,N_1968);
or U2044 (N_2044,N_1976,N_1965);
nor U2045 (N_2045,N_1991,N_1969);
nor U2046 (N_2046,N_1995,N_1966);
or U2047 (N_2047,N_1997,N_1984);
nand U2048 (N_2048,N_1974,N_1962);
nor U2049 (N_2049,N_1956,N_1964);
or U2050 (N_2050,N_2041,N_2000);
or U2051 (N_2051,N_2012,N_2010);
nand U2052 (N_2052,N_2006,N_2009);
or U2053 (N_2053,N_2035,N_2007);
nor U2054 (N_2054,N_2034,N_2026);
nor U2055 (N_2055,N_2028,N_2033);
or U2056 (N_2056,N_2037,N_2022);
nor U2057 (N_2057,N_2049,N_2021);
or U2058 (N_2058,N_2029,N_2004);
nand U2059 (N_2059,N_2001,N_2045);
nand U2060 (N_2060,N_2044,N_2040);
or U2061 (N_2061,N_2002,N_2024);
nand U2062 (N_2062,N_2047,N_2019);
and U2063 (N_2063,N_2043,N_2003);
nand U2064 (N_2064,N_2008,N_2031);
nor U2065 (N_2065,N_2039,N_2014);
and U2066 (N_2066,N_2032,N_2027);
or U2067 (N_2067,N_2042,N_2020);
or U2068 (N_2068,N_2011,N_2036);
and U2069 (N_2069,N_2018,N_2016);
or U2070 (N_2070,N_2023,N_2046);
nor U2071 (N_2071,N_2015,N_2017);
or U2072 (N_2072,N_2005,N_2030);
and U2073 (N_2073,N_2048,N_2025);
nor U2074 (N_2074,N_2038,N_2013);
nand U2075 (N_2075,N_2020,N_2028);
or U2076 (N_2076,N_2037,N_2040);
nor U2077 (N_2077,N_2041,N_2031);
xnor U2078 (N_2078,N_2015,N_2022);
or U2079 (N_2079,N_2008,N_2035);
nor U2080 (N_2080,N_2028,N_2038);
nand U2081 (N_2081,N_2039,N_2004);
and U2082 (N_2082,N_2029,N_2006);
nor U2083 (N_2083,N_2021,N_2037);
or U2084 (N_2084,N_2017,N_2030);
nand U2085 (N_2085,N_2020,N_2033);
nand U2086 (N_2086,N_2018,N_2010);
or U2087 (N_2087,N_2043,N_2038);
and U2088 (N_2088,N_2009,N_2048);
and U2089 (N_2089,N_2040,N_2018);
or U2090 (N_2090,N_2016,N_2002);
nor U2091 (N_2091,N_2025,N_2045);
nand U2092 (N_2092,N_2036,N_2021);
and U2093 (N_2093,N_2016,N_2011);
and U2094 (N_2094,N_2007,N_2039);
and U2095 (N_2095,N_2047,N_2032);
or U2096 (N_2096,N_2038,N_2044);
or U2097 (N_2097,N_2021,N_2032);
or U2098 (N_2098,N_2021,N_2048);
nand U2099 (N_2099,N_2048,N_2002);
nand U2100 (N_2100,N_2050,N_2062);
and U2101 (N_2101,N_2075,N_2090);
nand U2102 (N_2102,N_2058,N_2077);
or U2103 (N_2103,N_2051,N_2060);
nand U2104 (N_2104,N_2063,N_2068);
nand U2105 (N_2105,N_2089,N_2069);
and U2106 (N_2106,N_2091,N_2057);
nor U2107 (N_2107,N_2064,N_2098);
and U2108 (N_2108,N_2096,N_2081);
or U2109 (N_2109,N_2087,N_2088);
nand U2110 (N_2110,N_2082,N_2066);
xor U2111 (N_2111,N_2099,N_2052);
xnor U2112 (N_2112,N_2095,N_2076);
nand U2113 (N_2113,N_2080,N_2059);
nand U2114 (N_2114,N_2097,N_2084);
nand U2115 (N_2115,N_2086,N_2071);
nor U2116 (N_2116,N_2093,N_2067);
nand U2117 (N_2117,N_2054,N_2083);
nor U2118 (N_2118,N_2073,N_2074);
or U2119 (N_2119,N_2094,N_2061);
nand U2120 (N_2120,N_2070,N_2065);
nand U2121 (N_2121,N_2079,N_2055);
nor U2122 (N_2122,N_2078,N_2092);
xor U2123 (N_2123,N_2053,N_2072);
nand U2124 (N_2124,N_2056,N_2085);
and U2125 (N_2125,N_2062,N_2057);
nand U2126 (N_2126,N_2089,N_2063);
and U2127 (N_2127,N_2077,N_2065);
and U2128 (N_2128,N_2060,N_2097);
and U2129 (N_2129,N_2087,N_2068);
nor U2130 (N_2130,N_2075,N_2089);
nand U2131 (N_2131,N_2061,N_2083);
and U2132 (N_2132,N_2082,N_2061);
nand U2133 (N_2133,N_2062,N_2068);
nand U2134 (N_2134,N_2087,N_2078);
or U2135 (N_2135,N_2075,N_2073);
or U2136 (N_2136,N_2084,N_2063);
or U2137 (N_2137,N_2085,N_2050);
nor U2138 (N_2138,N_2083,N_2078);
nor U2139 (N_2139,N_2070,N_2061);
nand U2140 (N_2140,N_2092,N_2076);
nor U2141 (N_2141,N_2054,N_2066);
and U2142 (N_2142,N_2073,N_2097);
and U2143 (N_2143,N_2054,N_2095);
or U2144 (N_2144,N_2069,N_2052);
or U2145 (N_2145,N_2053,N_2063);
or U2146 (N_2146,N_2083,N_2073);
and U2147 (N_2147,N_2057,N_2097);
nor U2148 (N_2148,N_2064,N_2054);
and U2149 (N_2149,N_2087,N_2059);
nor U2150 (N_2150,N_2112,N_2132);
nor U2151 (N_2151,N_2137,N_2130);
or U2152 (N_2152,N_2149,N_2147);
nand U2153 (N_2153,N_2138,N_2107);
nor U2154 (N_2154,N_2106,N_2136);
or U2155 (N_2155,N_2146,N_2100);
and U2156 (N_2156,N_2109,N_2110);
or U2157 (N_2157,N_2108,N_2122);
nand U2158 (N_2158,N_2115,N_2140);
and U2159 (N_2159,N_2144,N_2133);
or U2160 (N_2160,N_2104,N_2103);
nand U2161 (N_2161,N_2128,N_2117);
nand U2162 (N_2162,N_2142,N_2143);
and U2163 (N_2163,N_2102,N_2118);
nand U2164 (N_2164,N_2116,N_2105);
nor U2165 (N_2165,N_2121,N_2114);
or U2166 (N_2166,N_2135,N_2141);
and U2167 (N_2167,N_2119,N_2139);
or U2168 (N_2168,N_2101,N_2131);
nand U2169 (N_2169,N_2127,N_2125);
nand U2170 (N_2170,N_2148,N_2120);
and U2171 (N_2171,N_2111,N_2113);
or U2172 (N_2172,N_2134,N_2129);
and U2173 (N_2173,N_2123,N_2126);
and U2174 (N_2174,N_2145,N_2124);
and U2175 (N_2175,N_2107,N_2145);
or U2176 (N_2176,N_2148,N_2149);
or U2177 (N_2177,N_2125,N_2111);
nor U2178 (N_2178,N_2107,N_2109);
nand U2179 (N_2179,N_2146,N_2132);
nand U2180 (N_2180,N_2116,N_2126);
nor U2181 (N_2181,N_2113,N_2148);
nand U2182 (N_2182,N_2145,N_2148);
nand U2183 (N_2183,N_2140,N_2107);
nor U2184 (N_2184,N_2139,N_2130);
nand U2185 (N_2185,N_2116,N_2102);
and U2186 (N_2186,N_2142,N_2104);
nand U2187 (N_2187,N_2134,N_2143);
nand U2188 (N_2188,N_2140,N_2144);
nand U2189 (N_2189,N_2121,N_2127);
or U2190 (N_2190,N_2100,N_2103);
or U2191 (N_2191,N_2129,N_2138);
and U2192 (N_2192,N_2115,N_2148);
nor U2193 (N_2193,N_2111,N_2148);
and U2194 (N_2194,N_2101,N_2130);
or U2195 (N_2195,N_2130,N_2110);
nor U2196 (N_2196,N_2115,N_2143);
and U2197 (N_2197,N_2104,N_2136);
or U2198 (N_2198,N_2115,N_2104);
and U2199 (N_2199,N_2104,N_2133);
or U2200 (N_2200,N_2186,N_2174);
nand U2201 (N_2201,N_2187,N_2163);
nor U2202 (N_2202,N_2188,N_2177);
nor U2203 (N_2203,N_2165,N_2166);
nor U2204 (N_2204,N_2189,N_2170);
or U2205 (N_2205,N_2158,N_2154);
nor U2206 (N_2206,N_2175,N_2195);
nand U2207 (N_2207,N_2167,N_2198);
or U2208 (N_2208,N_2161,N_2179);
nand U2209 (N_2209,N_2183,N_2176);
nand U2210 (N_2210,N_2178,N_2199);
nand U2211 (N_2211,N_2185,N_2157);
nor U2212 (N_2212,N_2172,N_2182);
and U2213 (N_2213,N_2173,N_2156);
nand U2214 (N_2214,N_2151,N_2168);
or U2215 (N_2215,N_2193,N_2191);
nor U2216 (N_2216,N_2194,N_2153);
nand U2217 (N_2217,N_2169,N_2197);
nand U2218 (N_2218,N_2180,N_2164);
nor U2219 (N_2219,N_2159,N_2160);
nor U2220 (N_2220,N_2155,N_2152);
nor U2221 (N_2221,N_2162,N_2196);
and U2222 (N_2222,N_2150,N_2181);
and U2223 (N_2223,N_2171,N_2184);
nor U2224 (N_2224,N_2190,N_2192);
nor U2225 (N_2225,N_2188,N_2180);
or U2226 (N_2226,N_2156,N_2160);
and U2227 (N_2227,N_2157,N_2159);
or U2228 (N_2228,N_2181,N_2183);
nand U2229 (N_2229,N_2165,N_2174);
or U2230 (N_2230,N_2199,N_2185);
and U2231 (N_2231,N_2198,N_2191);
nand U2232 (N_2232,N_2162,N_2161);
and U2233 (N_2233,N_2153,N_2199);
nor U2234 (N_2234,N_2163,N_2167);
nor U2235 (N_2235,N_2176,N_2195);
nor U2236 (N_2236,N_2184,N_2173);
and U2237 (N_2237,N_2156,N_2179);
and U2238 (N_2238,N_2195,N_2190);
and U2239 (N_2239,N_2197,N_2155);
and U2240 (N_2240,N_2192,N_2180);
nand U2241 (N_2241,N_2188,N_2185);
nand U2242 (N_2242,N_2190,N_2179);
or U2243 (N_2243,N_2191,N_2177);
or U2244 (N_2244,N_2158,N_2195);
nor U2245 (N_2245,N_2158,N_2150);
and U2246 (N_2246,N_2163,N_2162);
and U2247 (N_2247,N_2156,N_2187);
nand U2248 (N_2248,N_2198,N_2195);
or U2249 (N_2249,N_2177,N_2152);
or U2250 (N_2250,N_2235,N_2227);
or U2251 (N_2251,N_2225,N_2222);
and U2252 (N_2252,N_2206,N_2211);
nor U2253 (N_2253,N_2220,N_2240);
nand U2254 (N_2254,N_2233,N_2215);
or U2255 (N_2255,N_2228,N_2230);
or U2256 (N_2256,N_2223,N_2224);
nand U2257 (N_2257,N_2203,N_2214);
and U2258 (N_2258,N_2202,N_2232);
or U2259 (N_2259,N_2248,N_2221);
nor U2260 (N_2260,N_2213,N_2207);
nand U2261 (N_2261,N_2205,N_2236);
nor U2262 (N_2262,N_2216,N_2229);
and U2263 (N_2263,N_2242,N_2239);
nor U2264 (N_2264,N_2204,N_2245);
nor U2265 (N_2265,N_2247,N_2243);
nand U2266 (N_2266,N_2238,N_2208);
and U2267 (N_2267,N_2231,N_2218);
nand U2268 (N_2268,N_2241,N_2217);
and U2269 (N_2269,N_2201,N_2237);
and U2270 (N_2270,N_2249,N_2210);
and U2271 (N_2271,N_2209,N_2244);
and U2272 (N_2272,N_2219,N_2234);
nand U2273 (N_2273,N_2200,N_2246);
or U2274 (N_2274,N_2212,N_2226);
xnor U2275 (N_2275,N_2200,N_2227);
or U2276 (N_2276,N_2217,N_2223);
nand U2277 (N_2277,N_2222,N_2206);
and U2278 (N_2278,N_2239,N_2248);
or U2279 (N_2279,N_2201,N_2231);
nor U2280 (N_2280,N_2244,N_2215);
nor U2281 (N_2281,N_2230,N_2217);
or U2282 (N_2282,N_2236,N_2209);
or U2283 (N_2283,N_2248,N_2240);
nand U2284 (N_2284,N_2248,N_2206);
nor U2285 (N_2285,N_2231,N_2213);
or U2286 (N_2286,N_2226,N_2203);
and U2287 (N_2287,N_2231,N_2245);
and U2288 (N_2288,N_2217,N_2209);
or U2289 (N_2289,N_2223,N_2230);
and U2290 (N_2290,N_2215,N_2238);
nand U2291 (N_2291,N_2215,N_2236);
and U2292 (N_2292,N_2218,N_2236);
nand U2293 (N_2293,N_2220,N_2246);
nor U2294 (N_2294,N_2204,N_2217);
nor U2295 (N_2295,N_2246,N_2239);
and U2296 (N_2296,N_2245,N_2232);
nor U2297 (N_2297,N_2232,N_2247);
nor U2298 (N_2298,N_2210,N_2225);
nand U2299 (N_2299,N_2210,N_2214);
or U2300 (N_2300,N_2269,N_2298);
or U2301 (N_2301,N_2282,N_2283);
nor U2302 (N_2302,N_2265,N_2262);
nand U2303 (N_2303,N_2254,N_2299);
and U2304 (N_2304,N_2253,N_2250);
and U2305 (N_2305,N_2257,N_2267);
and U2306 (N_2306,N_2297,N_2272);
or U2307 (N_2307,N_2278,N_2271);
nand U2308 (N_2308,N_2285,N_2255);
nor U2309 (N_2309,N_2270,N_2289);
or U2310 (N_2310,N_2286,N_2264);
nor U2311 (N_2311,N_2263,N_2284);
or U2312 (N_2312,N_2251,N_2275);
nand U2313 (N_2313,N_2274,N_2258);
nor U2314 (N_2314,N_2252,N_2273);
or U2315 (N_2315,N_2287,N_2292);
and U2316 (N_2316,N_2290,N_2296);
and U2317 (N_2317,N_2266,N_2256);
nor U2318 (N_2318,N_2291,N_2288);
and U2319 (N_2319,N_2260,N_2295);
nand U2320 (N_2320,N_2279,N_2276);
nor U2321 (N_2321,N_2280,N_2277);
nand U2322 (N_2322,N_2293,N_2261);
or U2323 (N_2323,N_2294,N_2259);
nand U2324 (N_2324,N_2281,N_2268);
nor U2325 (N_2325,N_2299,N_2286);
or U2326 (N_2326,N_2252,N_2266);
or U2327 (N_2327,N_2294,N_2251);
or U2328 (N_2328,N_2289,N_2279);
nand U2329 (N_2329,N_2274,N_2286);
nor U2330 (N_2330,N_2268,N_2278);
nor U2331 (N_2331,N_2277,N_2257);
nand U2332 (N_2332,N_2276,N_2298);
or U2333 (N_2333,N_2254,N_2271);
nor U2334 (N_2334,N_2256,N_2286);
and U2335 (N_2335,N_2298,N_2274);
or U2336 (N_2336,N_2264,N_2291);
and U2337 (N_2337,N_2278,N_2250);
nand U2338 (N_2338,N_2252,N_2290);
or U2339 (N_2339,N_2256,N_2265);
or U2340 (N_2340,N_2263,N_2295);
nand U2341 (N_2341,N_2259,N_2269);
or U2342 (N_2342,N_2263,N_2277);
nor U2343 (N_2343,N_2299,N_2298);
nor U2344 (N_2344,N_2288,N_2258);
or U2345 (N_2345,N_2297,N_2256);
nor U2346 (N_2346,N_2261,N_2251);
or U2347 (N_2347,N_2287,N_2273);
nor U2348 (N_2348,N_2289,N_2253);
or U2349 (N_2349,N_2258,N_2295);
or U2350 (N_2350,N_2304,N_2332);
or U2351 (N_2351,N_2303,N_2347);
nand U2352 (N_2352,N_2334,N_2325);
and U2353 (N_2353,N_2321,N_2339);
xor U2354 (N_2354,N_2344,N_2320);
and U2355 (N_2355,N_2335,N_2315);
nor U2356 (N_2356,N_2341,N_2337);
nand U2357 (N_2357,N_2301,N_2331);
and U2358 (N_2358,N_2338,N_2333);
or U2359 (N_2359,N_2349,N_2328);
or U2360 (N_2360,N_2340,N_2318);
nand U2361 (N_2361,N_2345,N_2330);
nand U2362 (N_2362,N_2317,N_2309);
or U2363 (N_2363,N_2324,N_2306);
and U2364 (N_2364,N_2302,N_2346);
and U2365 (N_2365,N_2329,N_2336);
and U2366 (N_2366,N_2308,N_2348);
nor U2367 (N_2367,N_2343,N_2305);
nand U2368 (N_2368,N_2310,N_2312);
nand U2369 (N_2369,N_2322,N_2327);
nor U2370 (N_2370,N_2342,N_2326);
or U2371 (N_2371,N_2314,N_2313);
nor U2372 (N_2372,N_2311,N_2300);
nor U2373 (N_2373,N_2319,N_2307);
nor U2374 (N_2374,N_2316,N_2323);
nand U2375 (N_2375,N_2334,N_2313);
nand U2376 (N_2376,N_2330,N_2315);
nand U2377 (N_2377,N_2344,N_2315);
or U2378 (N_2378,N_2328,N_2333);
nor U2379 (N_2379,N_2305,N_2323);
or U2380 (N_2380,N_2347,N_2333);
or U2381 (N_2381,N_2341,N_2344);
and U2382 (N_2382,N_2313,N_2339);
nor U2383 (N_2383,N_2307,N_2330);
nor U2384 (N_2384,N_2306,N_2331);
and U2385 (N_2385,N_2346,N_2318);
nand U2386 (N_2386,N_2317,N_2331);
nand U2387 (N_2387,N_2306,N_2348);
or U2388 (N_2388,N_2329,N_2322);
nor U2389 (N_2389,N_2317,N_2333);
or U2390 (N_2390,N_2344,N_2327);
nor U2391 (N_2391,N_2307,N_2322);
or U2392 (N_2392,N_2338,N_2314);
nor U2393 (N_2393,N_2325,N_2328);
and U2394 (N_2394,N_2344,N_2336);
nand U2395 (N_2395,N_2318,N_2331);
or U2396 (N_2396,N_2303,N_2332);
nand U2397 (N_2397,N_2318,N_2333);
or U2398 (N_2398,N_2320,N_2302);
nand U2399 (N_2399,N_2330,N_2302);
nand U2400 (N_2400,N_2365,N_2361);
nor U2401 (N_2401,N_2387,N_2373);
and U2402 (N_2402,N_2381,N_2383);
nor U2403 (N_2403,N_2385,N_2374);
or U2404 (N_2404,N_2363,N_2353);
nor U2405 (N_2405,N_2356,N_2388);
or U2406 (N_2406,N_2358,N_2372);
nor U2407 (N_2407,N_2375,N_2362);
nand U2408 (N_2408,N_2352,N_2396);
nor U2409 (N_2409,N_2370,N_2380);
nand U2410 (N_2410,N_2364,N_2377);
nand U2411 (N_2411,N_2367,N_2354);
or U2412 (N_2412,N_2368,N_2389);
and U2413 (N_2413,N_2359,N_2394);
or U2414 (N_2414,N_2393,N_2376);
and U2415 (N_2415,N_2355,N_2369);
or U2416 (N_2416,N_2398,N_2382);
nor U2417 (N_2417,N_2371,N_2357);
or U2418 (N_2418,N_2391,N_2392);
nor U2419 (N_2419,N_2386,N_2395);
or U2420 (N_2420,N_2350,N_2379);
and U2421 (N_2421,N_2378,N_2384);
nor U2422 (N_2422,N_2390,N_2351);
nor U2423 (N_2423,N_2360,N_2366);
or U2424 (N_2424,N_2399,N_2397);
and U2425 (N_2425,N_2376,N_2382);
or U2426 (N_2426,N_2360,N_2382);
or U2427 (N_2427,N_2388,N_2372);
and U2428 (N_2428,N_2393,N_2370);
and U2429 (N_2429,N_2351,N_2396);
or U2430 (N_2430,N_2388,N_2384);
nor U2431 (N_2431,N_2361,N_2371);
and U2432 (N_2432,N_2384,N_2376);
and U2433 (N_2433,N_2350,N_2389);
nor U2434 (N_2434,N_2357,N_2385);
or U2435 (N_2435,N_2357,N_2381);
nand U2436 (N_2436,N_2354,N_2382);
nand U2437 (N_2437,N_2397,N_2352);
and U2438 (N_2438,N_2372,N_2374);
nor U2439 (N_2439,N_2352,N_2391);
nand U2440 (N_2440,N_2370,N_2354);
xnor U2441 (N_2441,N_2378,N_2373);
and U2442 (N_2442,N_2399,N_2372);
nand U2443 (N_2443,N_2353,N_2364);
and U2444 (N_2444,N_2372,N_2387);
nand U2445 (N_2445,N_2356,N_2374);
nor U2446 (N_2446,N_2375,N_2365);
nand U2447 (N_2447,N_2382,N_2358);
or U2448 (N_2448,N_2378,N_2381);
or U2449 (N_2449,N_2384,N_2361);
or U2450 (N_2450,N_2429,N_2405);
nand U2451 (N_2451,N_2421,N_2440);
nand U2452 (N_2452,N_2412,N_2441);
nand U2453 (N_2453,N_2432,N_2420);
nor U2454 (N_2454,N_2430,N_2417);
nand U2455 (N_2455,N_2431,N_2414);
xor U2456 (N_2456,N_2434,N_2428);
and U2457 (N_2457,N_2425,N_2449);
nand U2458 (N_2458,N_2415,N_2446);
nor U2459 (N_2459,N_2401,N_2433);
or U2460 (N_2460,N_2413,N_2422);
or U2461 (N_2461,N_2407,N_2436);
and U2462 (N_2462,N_2409,N_2411);
nand U2463 (N_2463,N_2444,N_2418);
or U2464 (N_2464,N_2437,N_2408);
nand U2465 (N_2465,N_2406,N_2419);
and U2466 (N_2466,N_2402,N_2435);
and U2467 (N_2467,N_2424,N_2438);
and U2468 (N_2468,N_2400,N_2445);
nand U2469 (N_2469,N_2443,N_2423);
nor U2470 (N_2470,N_2447,N_2442);
and U2471 (N_2471,N_2404,N_2416);
nand U2472 (N_2472,N_2426,N_2439);
nor U2473 (N_2473,N_2427,N_2448);
nor U2474 (N_2474,N_2410,N_2403);
and U2475 (N_2475,N_2428,N_2445);
and U2476 (N_2476,N_2403,N_2416);
or U2477 (N_2477,N_2416,N_2413);
nor U2478 (N_2478,N_2403,N_2425);
and U2479 (N_2479,N_2403,N_2414);
nand U2480 (N_2480,N_2434,N_2441);
xnor U2481 (N_2481,N_2441,N_2449);
nand U2482 (N_2482,N_2400,N_2430);
or U2483 (N_2483,N_2413,N_2425);
nand U2484 (N_2484,N_2416,N_2432);
nor U2485 (N_2485,N_2428,N_2442);
and U2486 (N_2486,N_2441,N_2432);
nor U2487 (N_2487,N_2441,N_2424);
nor U2488 (N_2488,N_2421,N_2436);
nand U2489 (N_2489,N_2437,N_2443);
nor U2490 (N_2490,N_2433,N_2419);
or U2491 (N_2491,N_2434,N_2419);
nor U2492 (N_2492,N_2432,N_2446);
or U2493 (N_2493,N_2433,N_2402);
nand U2494 (N_2494,N_2427,N_2420);
or U2495 (N_2495,N_2428,N_2409);
nand U2496 (N_2496,N_2401,N_2406);
or U2497 (N_2497,N_2445,N_2412);
and U2498 (N_2498,N_2444,N_2407);
and U2499 (N_2499,N_2436,N_2403);
nor U2500 (N_2500,N_2465,N_2476);
and U2501 (N_2501,N_2454,N_2462);
and U2502 (N_2502,N_2488,N_2487);
xnor U2503 (N_2503,N_2499,N_2482);
and U2504 (N_2504,N_2459,N_2485);
or U2505 (N_2505,N_2495,N_2481);
nand U2506 (N_2506,N_2490,N_2468);
or U2507 (N_2507,N_2475,N_2450);
or U2508 (N_2508,N_2463,N_2492);
nand U2509 (N_2509,N_2469,N_2496);
and U2510 (N_2510,N_2464,N_2451);
or U2511 (N_2511,N_2458,N_2478);
nand U2512 (N_2512,N_2461,N_2474);
nand U2513 (N_2513,N_2486,N_2489);
nor U2514 (N_2514,N_2473,N_2494);
or U2515 (N_2515,N_2466,N_2484);
nor U2516 (N_2516,N_2470,N_2467);
or U2517 (N_2517,N_2456,N_2483);
nand U2518 (N_2518,N_2452,N_2460);
nand U2519 (N_2519,N_2472,N_2455);
and U2520 (N_2520,N_2491,N_2493);
nor U2521 (N_2521,N_2479,N_2471);
or U2522 (N_2522,N_2498,N_2457);
or U2523 (N_2523,N_2497,N_2453);
or U2524 (N_2524,N_2480,N_2477);
nor U2525 (N_2525,N_2498,N_2456);
and U2526 (N_2526,N_2477,N_2493);
nand U2527 (N_2527,N_2454,N_2489);
and U2528 (N_2528,N_2450,N_2473);
nor U2529 (N_2529,N_2456,N_2457);
nand U2530 (N_2530,N_2473,N_2455);
or U2531 (N_2531,N_2470,N_2481);
nand U2532 (N_2532,N_2494,N_2471);
or U2533 (N_2533,N_2489,N_2456);
nand U2534 (N_2534,N_2459,N_2482);
nand U2535 (N_2535,N_2483,N_2465);
nor U2536 (N_2536,N_2458,N_2470);
nor U2537 (N_2537,N_2477,N_2461);
nor U2538 (N_2538,N_2498,N_2481);
nand U2539 (N_2539,N_2458,N_2456);
or U2540 (N_2540,N_2461,N_2475);
nand U2541 (N_2541,N_2456,N_2474);
nand U2542 (N_2542,N_2475,N_2456);
nor U2543 (N_2543,N_2462,N_2483);
nand U2544 (N_2544,N_2491,N_2459);
nor U2545 (N_2545,N_2485,N_2455);
or U2546 (N_2546,N_2492,N_2487);
and U2547 (N_2547,N_2475,N_2481);
or U2548 (N_2548,N_2470,N_2492);
or U2549 (N_2549,N_2496,N_2483);
nor U2550 (N_2550,N_2501,N_2523);
nand U2551 (N_2551,N_2509,N_2536);
and U2552 (N_2552,N_2522,N_2532);
nand U2553 (N_2553,N_2525,N_2519);
or U2554 (N_2554,N_2511,N_2535);
nor U2555 (N_2555,N_2520,N_2518);
nor U2556 (N_2556,N_2543,N_2524);
and U2557 (N_2557,N_2546,N_2503);
nor U2558 (N_2558,N_2547,N_2537);
nand U2559 (N_2559,N_2500,N_2530);
nand U2560 (N_2560,N_2506,N_2528);
nor U2561 (N_2561,N_2534,N_2548);
or U2562 (N_2562,N_2505,N_2533);
or U2563 (N_2563,N_2542,N_2521);
and U2564 (N_2564,N_2517,N_2529);
or U2565 (N_2565,N_2527,N_2526);
nor U2566 (N_2566,N_2508,N_2502);
and U2567 (N_2567,N_2538,N_2514);
and U2568 (N_2568,N_2504,N_2549);
nor U2569 (N_2569,N_2545,N_2510);
nor U2570 (N_2570,N_2541,N_2540);
or U2571 (N_2571,N_2507,N_2512);
nor U2572 (N_2572,N_2544,N_2513);
and U2573 (N_2573,N_2531,N_2516);
nor U2574 (N_2574,N_2515,N_2539);
and U2575 (N_2575,N_2548,N_2527);
nand U2576 (N_2576,N_2544,N_2521);
nand U2577 (N_2577,N_2506,N_2539);
and U2578 (N_2578,N_2549,N_2518);
and U2579 (N_2579,N_2500,N_2519);
nor U2580 (N_2580,N_2544,N_2549);
or U2581 (N_2581,N_2519,N_2516);
nor U2582 (N_2582,N_2503,N_2518);
nor U2583 (N_2583,N_2540,N_2516);
nand U2584 (N_2584,N_2516,N_2509);
nand U2585 (N_2585,N_2529,N_2538);
nor U2586 (N_2586,N_2548,N_2509);
and U2587 (N_2587,N_2527,N_2528);
nand U2588 (N_2588,N_2528,N_2512);
and U2589 (N_2589,N_2501,N_2533);
nor U2590 (N_2590,N_2525,N_2522);
nand U2591 (N_2591,N_2522,N_2523);
and U2592 (N_2592,N_2516,N_2501);
nor U2593 (N_2593,N_2512,N_2539);
and U2594 (N_2594,N_2517,N_2510);
nor U2595 (N_2595,N_2536,N_2548);
nand U2596 (N_2596,N_2516,N_2542);
or U2597 (N_2597,N_2507,N_2546);
or U2598 (N_2598,N_2547,N_2531);
and U2599 (N_2599,N_2521,N_2545);
xor U2600 (N_2600,N_2593,N_2579);
nand U2601 (N_2601,N_2597,N_2594);
and U2602 (N_2602,N_2569,N_2564);
nand U2603 (N_2603,N_2589,N_2558);
nand U2604 (N_2604,N_2570,N_2559);
and U2605 (N_2605,N_2552,N_2557);
and U2606 (N_2606,N_2562,N_2568);
or U2607 (N_2607,N_2554,N_2595);
nand U2608 (N_2608,N_2577,N_2588);
nand U2609 (N_2609,N_2598,N_2571);
nor U2610 (N_2610,N_2580,N_2585);
and U2611 (N_2611,N_2563,N_2582);
nand U2612 (N_2612,N_2560,N_2565);
nor U2613 (N_2613,N_2586,N_2581);
nor U2614 (N_2614,N_2584,N_2578);
or U2615 (N_2615,N_2576,N_2555);
or U2616 (N_2616,N_2573,N_2561);
nand U2617 (N_2617,N_2574,N_2587);
or U2618 (N_2618,N_2566,N_2575);
and U2619 (N_2619,N_2556,N_2583);
and U2620 (N_2620,N_2592,N_2553);
nand U2621 (N_2621,N_2550,N_2590);
or U2622 (N_2622,N_2572,N_2567);
nor U2623 (N_2623,N_2596,N_2599);
nand U2624 (N_2624,N_2591,N_2551);
and U2625 (N_2625,N_2558,N_2596);
xor U2626 (N_2626,N_2585,N_2570);
nand U2627 (N_2627,N_2579,N_2582);
nand U2628 (N_2628,N_2567,N_2562);
and U2629 (N_2629,N_2552,N_2592);
and U2630 (N_2630,N_2576,N_2574);
and U2631 (N_2631,N_2593,N_2569);
nand U2632 (N_2632,N_2591,N_2560);
and U2633 (N_2633,N_2551,N_2552);
xor U2634 (N_2634,N_2552,N_2560);
nor U2635 (N_2635,N_2550,N_2554);
and U2636 (N_2636,N_2566,N_2597);
nor U2637 (N_2637,N_2556,N_2555);
or U2638 (N_2638,N_2585,N_2599);
or U2639 (N_2639,N_2553,N_2583);
or U2640 (N_2640,N_2580,N_2598);
and U2641 (N_2641,N_2579,N_2576);
nor U2642 (N_2642,N_2575,N_2569);
and U2643 (N_2643,N_2559,N_2573);
and U2644 (N_2644,N_2569,N_2578);
nand U2645 (N_2645,N_2556,N_2590);
or U2646 (N_2646,N_2598,N_2590);
nand U2647 (N_2647,N_2554,N_2574);
nor U2648 (N_2648,N_2551,N_2594);
and U2649 (N_2649,N_2565,N_2580);
nand U2650 (N_2650,N_2609,N_2600);
and U2651 (N_2651,N_2604,N_2615);
nand U2652 (N_2652,N_2605,N_2635);
and U2653 (N_2653,N_2643,N_2630);
nor U2654 (N_2654,N_2602,N_2649);
or U2655 (N_2655,N_2647,N_2614);
nor U2656 (N_2656,N_2634,N_2619);
or U2657 (N_2657,N_2636,N_2644);
nand U2658 (N_2658,N_2613,N_2633);
nand U2659 (N_2659,N_2637,N_2646);
and U2660 (N_2660,N_2639,N_2628);
or U2661 (N_2661,N_2612,N_2622);
nand U2662 (N_2662,N_2608,N_2641);
and U2663 (N_2663,N_2632,N_2645);
and U2664 (N_2664,N_2626,N_2611);
and U2665 (N_2665,N_2610,N_2603);
or U2666 (N_2666,N_2648,N_2618);
nand U2667 (N_2667,N_2640,N_2617);
and U2668 (N_2668,N_2623,N_2620);
nand U2669 (N_2669,N_2625,N_2642);
or U2670 (N_2670,N_2606,N_2624);
or U2671 (N_2671,N_2627,N_2616);
or U2672 (N_2672,N_2601,N_2607);
nand U2673 (N_2673,N_2629,N_2621);
nor U2674 (N_2674,N_2638,N_2631);
and U2675 (N_2675,N_2636,N_2647);
or U2676 (N_2676,N_2647,N_2617);
nor U2677 (N_2677,N_2626,N_2630);
and U2678 (N_2678,N_2645,N_2639);
and U2679 (N_2679,N_2636,N_2646);
nand U2680 (N_2680,N_2627,N_2646);
or U2681 (N_2681,N_2604,N_2610);
and U2682 (N_2682,N_2642,N_2632);
or U2683 (N_2683,N_2626,N_2602);
and U2684 (N_2684,N_2648,N_2624);
nor U2685 (N_2685,N_2606,N_2620);
and U2686 (N_2686,N_2612,N_2647);
nand U2687 (N_2687,N_2616,N_2633);
or U2688 (N_2688,N_2638,N_2615);
nor U2689 (N_2689,N_2606,N_2621);
and U2690 (N_2690,N_2605,N_2634);
nand U2691 (N_2691,N_2648,N_2605);
nand U2692 (N_2692,N_2649,N_2604);
nor U2693 (N_2693,N_2633,N_2604);
nand U2694 (N_2694,N_2645,N_2637);
and U2695 (N_2695,N_2626,N_2629);
and U2696 (N_2696,N_2638,N_2611);
xnor U2697 (N_2697,N_2645,N_2600);
nand U2698 (N_2698,N_2631,N_2627);
nand U2699 (N_2699,N_2618,N_2638);
nand U2700 (N_2700,N_2657,N_2689);
or U2701 (N_2701,N_2664,N_2679);
nand U2702 (N_2702,N_2677,N_2676);
or U2703 (N_2703,N_2672,N_2653);
xor U2704 (N_2704,N_2687,N_2684);
nand U2705 (N_2705,N_2675,N_2655);
nor U2706 (N_2706,N_2696,N_2682);
and U2707 (N_2707,N_2681,N_2692);
or U2708 (N_2708,N_2660,N_2650);
nand U2709 (N_2709,N_2698,N_2685);
or U2710 (N_2710,N_2688,N_2659);
or U2711 (N_2711,N_2686,N_2662);
and U2712 (N_2712,N_2683,N_2697);
nor U2713 (N_2713,N_2652,N_2693);
nand U2714 (N_2714,N_2674,N_2658);
and U2715 (N_2715,N_2690,N_2670);
nand U2716 (N_2716,N_2666,N_2678);
nor U2717 (N_2717,N_2695,N_2654);
nor U2718 (N_2718,N_2691,N_2671);
nand U2719 (N_2719,N_2680,N_2667);
and U2720 (N_2720,N_2694,N_2651);
nand U2721 (N_2721,N_2699,N_2661);
nand U2722 (N_2722,N_2669,N_2663);
and U2723 (N_2723,N_2668,N_2673);
nor U2724 (N_2724,N_2656,N_2665);
and U2725 (N_2725,N_2674,N_2693);
and U2726 (N_2726,N_2677,N_2670);
nand U2727 (N_2727,N_2662,N_2655);
nand U2728 (N_2728,N_2657,N_2683);
or U2729 (N_2729,N_2663,N_2667);
or U2730 (N_2730,N_2669,N_2699);
nor U2731 (N_2731,N_2697,N_2656);
or U2732 (N_2732,N_2698,N_2689);
or U2733 (N_2733,N_2663,N_2695);
nor U2734 (N_2734,N_2693,N_2659);
nor U2735 (N_2735,N_2677,N_2684);
nor U2736 (N_2736,N_2695,N_2677);
and U2737 (N_2737,N_2692,N_2684);
and U2738 (N_2738,N_2681,N_2695);
and U2739 (N_2739,N_2675,N_2670);
and U2740 (N_2740,N_2675,N_2666);
or U2741 (N_2741,N_2697,N_2660);
and U2742 (N_2742,N_2656,N_2684);
nor U2743 (N_2743,N_2688,N_2679);
nor U2744 (N_2744,N_2671,N_2652);
nor U2745 (N_2745,N_2667,N_2696);
nor U2746 (N_2746,N_2661,N_2697);
and U2747 (N_2747,N_2694,N_2675);
or U2748 (N_2748,N_2672,N_2652);
or U2749 (N_2749,N_2678,N_2659);
and U2750 (N_2750,N_2703,N_2741);
nand U2751 (N_2751,N_2734,N_2720);
xnor U2752 (N_2752,N_2729,N_2706);
and U2753 (N_2753,N_2708,N_2736);
nor U2754 (N_2754,N_2731,N_2727);
nor U2755 (N_2755,N_2710,N_2714);
or U2756 (N_2756,N_2748,N_2738);
or U2757 (N_2757,N_2745,N_2721);
and U2758 (N_2758,N_2730,N_2735);
and U2759 (N_2759,N_2713,N_2707);
or U2760 (N_2760,N_2733,N_2716);
and U2761 (N_2761,N_2723,N_2728);
nand U2762 (N_2762,N_2722,N_2700);
nand U2763 (N_2763,N_2717,N_2712);
or U2764 (N_2764,N_2726,N_2718);
or U2765 (N_2765,N_2743,N_2732);
or U2766 (N_2766,N_2739,N_2724);
or U2767 (N_2767,N_2709,N_2746);
nor U2768 (N_2768,N_2704,N_2747);
and U2769 (N_2769,N_2705,N_2740);
and U2770 (N_2770,N_2725,N_2719);
or U2771 (N_2771,N_2744,N_2702);
or U2772 (N_2772,N_2711,N_2737);
and U2773 (N_2773,N_2715,N_2742);
nand U2774 (N_2774,N_2749,N_2701);
nand U2775 (N_2775,N_2716,N_2702);
and U2776 (N_2776,N_2735,N_2709);
nor U2777 (N_2777,N_2737,N_2726);
and U2778 (N_2778,N_2749,N_2702);
nand U2779 (N_2779,N_2726,N_2733);
and U2780 (N_2780,N_2700,N_2724);
nand U2781 (N_2781,N_2727,N_2701);
nor U2782 (N_2782,N_2708,N_2733);
or U2783 (N_2783,N_2731,N_2723);
nor U2784 (N_2784,N_2704,N_2736);
and U2785 (N_2785,N_2740,N_2731);
or U2786 (N_2786,N_2701,N_2741);
and U2787 (N_2787,N_2720,N_2745);
and U2788 (N_2788,N_2709,N_2729);
or U2789 (N_2789,N_2744,N_2720);
or U2790 (N_2790,N_2726,N_2740);
xnor U2791 (N_2791,N_2723,N_2727);
nand U2792 (N_2792,N_2746,N_2708);
or U2793 (N_2793,N_2731,N_2745);
nand U2794 (N_2794,N_2736,N_2712);
or U2795 (N_2795,N_2703,N_2713);
and U2796 (N_2796,N_2734,N_2709);
nor U2797 (N_2797,N_2743,N_2747);
and U2798 (N_2798,N_2749,N_2709);
and U2799 (N_2799,N_2737,N_2715);
nor U2800 (N_2800,N_2769,N_2790);
nor U2801 (N_2801,N_2770,N_2750);
nor U2802 (N_2802,N_2752,N_2762);
or U2803 (N_2803,N_2771,N_2765);
or U2804 (N_2804,N_2754,N_2766);
nand U2805 (N_2805,N_2764,N_2753);
or U2806 (N_2806,N_2779,N_2773);
nand U2807 (N_2807,N_2776,N_2777);
nand U2808 (N_2808,N_2792,N_2775);
or U2809 (N_2809,N_2751,N_2799);
or U2810 (N_2810,N_2786,N_2796);
or U2811 (N_2811,N_2759,N_2760);
nand U2812 (N_2812,N_2778,N_2798);
nand U2813 (N_2813,N_2772,N_2787);
nand U2814 (N_2814,N_2758,N_2774);
and U2815 (N_2815,N_2755,N_2763);
nand U2816 (N_2816,N_2794,N_2783);
nor U2817 (N_2817,N_2780,N_2797);
and U2818 (N_2818,N_2757,N_2756);
and U2819 (N_2819,N_2793,N_2781);
nand U2820 (N_2820,N_2768,N_2767);
or U2821 (N_2821,N_2782,N_2788);
nor U2822 (N_2822,N_2795,N_2789);
and U2823 (N_2823,N_2791,N_2785);
nand U2824 (N_2824,N_2761,N_2784);
nand U2825 (N_2825,N_2767,N_2775);
nand U2826 (N_2826,N_2752,N_2780);
nor U2827 (N_2827,N_2770,N_2753);
and U2828 (N_2828,N_2762,N_2794);
and U2829 (N_2829,N_2792,N_2769);
nor U2830 (N_2830,N_2788,N_2754);
nand U2831 (N_2831,N_2762,N_2782);
or U2832 (N_2832,N_2795,N_2751);
or U2833 (N_2833,N_2795,N_2775);
nand U2834 (N_2834,N_2778,N_2768);
or U2835 (N_2835,N_2759,N_2764);
nand U2836 (N_2836,N_2786,N_2755);
nor U2837 (N_2837,N_2755,N_2772);
or U2838 (N_2838,N_2750,N_2791);
and U2839 (N_2839,N_2769,N_2797);
nand U2840 (N_2840,N_2797,N_2777);
nand U2841 (N_2841,N_2766,N_2794);
or U2842 (N_2842,N_2770,N_2756);
nand U2843 (N_2843,N_2756,N_2785);
and U2844 (N_2844,N_2765,N_2795);
nor U2845 (N_2845,N_2785,N_2794);
and U2846 (N_2846,N_2798,N_2751);
or U2847 (N_2847,N_2796,N_2767);
nor U2848 (N_2848,N_2767,N_2794);
nor U2849 (N_2849,N_2768,N_2794);
or U2850 (N_2850,N_2820,N_2842);
or U2851 (N_2851,N_2827,N_2810);
nand U2852 (N_2852,N_2829,N_2807);
nand U2853 (N_2853,N_2818,N_2805);
or U2854 (N_2854,N_2812,N_2802);
nand U2855 (N_2855,N_2825,N_2838);
or U2856 (N_2856,N_2817,N_2830);
or U2857 (N_2857,N_2822,N_2813);
and U2858 (N_2858,N_2844,N_2801);
and U2859 (N_2859,N_2828,N_2848);
and U2860 (N_2860,N_2809,N_2841);
or U2861 (N_2861,N_2806,N_2824);
nor U2862 (N_2862,N_2849,N_2840);
nor U2863 (N_2863,N_2815,N_2836);
xor U2864 (N_2864,N_2816,N_2803);
or U2865 (N_2865,N_2833,N_2845);
nand U2866 (N_2866,N_2821,N_2831);
or U2867 (N_2867,N_2837,N_2800);
and U2868 (N_2868,N_2832,N_2804);
nor U2869 (N_2869,N_2819,N_2847);
or U2870 (N_2870,N_2846,N_2843);
and U2871 (N_2871,N_2814,N_2834);
and U2872 (N_2872,N_2823,N_2826);
and U2873 (N_2873,N_2808,N_2835);
or U2874 (N_2874,N_2839,N_2811);
nor U2875 (N_2875,N_2811,N_2814);
or U2876 (N_2876,N_2806,N_2819);
nand U2877 (N_2877,N_2821,N_2817);
nor U2878 (N_2878,N_2847,N_2810);
or U2879 (N_2879,N_2829,N_2849);
or U2880 (N_2880,N_2826,N_2833);
or U2881 (N_2881,N_2835,N_2822);
nor U2882 (N_2882,N_2838,N_2816);
nor U2883 (N_2883,N_2808,N_2836);
nand U2884 (N_2884,N_2821,N_2845);
nand U2885 (N_2885,N_2806,N_2838);
xnor U2886 (N_2886,N_2836,N_2821);
nand U2887 (N_2887,N_2842,N_2812);
or U2888 (N_2888,N_2833,N_2810);
or U2889 (N_2889,N_2801,N_2834);
and U2890 (N_2890,N_2820,N_2825);
nor U2891 (N_2891,N_2843,N_2820);
and U2892 (N_2892,N_2829,N_2819);
nand U2893 (N_2893,N_2815,N_2830);
or U2894 (N_2894,N_2849,N_2841);
nor U2895 (N_2895,N_2805,N_2825);
or U2896 (N_2896,N_2820,N_2816);
nor U2897 (N_2897,N_2822,N_2818);
nor U2898 (N_2898,N_2842,N_2810);
nand U2899 (N_2899,N_2803,N_2810);
nand U2900 (N_2900,N_2865,N_2877);
or U2901 (N_2901,N_2874,N_2886);
or U2902 (N_2902,N_2898,N_2899);
or U2903 (N_2903,N_2871,N_2882);
and U2904 (N_2904,N_2859,N_2864);
and U2905 (N_2905,N_2893,N_2889);
and U2906 (N_2906,N_2860,N_2876);
nor U2907 (N_2907,N_2851,N_2861);
and U2908 (N_2908,N_2894,N_2867);
or U2909 (N_2909,N_2883,N_2853);
and U2910 (N_2910,N_2855,N_2890);
xnor U2911 (N_2911,N_2858,N_2862);
and U2912 (N_2912,N_2879,N_2887);
nand U2913 (N_2913,N_2896,N_2880);
nand U2914 (N_2914,N_2888,N_2856);
and U2915 (N_2915,N_2866,N_2863);
and U2916 (N_2916,N_2884,N_2878);
or U2917 (N_2917,N_2873,N_2854);
and U2918 (N_2918,N_2895,N_2891);
and U2919 (N_2919,N_2892,N_2850);
nand U2920 (N_2920,N_2869,N_2881);
nand U2921 (N_2921,N_2875,N_2852);
or U2922 (N_2922,N_2885,N_2857);
or U2923 (N_2923,N_2897,N_2868);
and U2924 (N_2924,N_2872,N_2870);
nand U2925 (N_2925,N_2855,N_2894);
and U2926 (N_2926,N_2867,N_2851);
or U2927 (N_2927,N_2861,N_2852);
nand U2928 (N_2928,N_2850,N_2853);
and U2929 (N_2929,N_2898,N_2854);
nor U2930 (N_2930,N_2857,N_2863);
nor U2931 (N_2931,N_2856,N_2861);
nand U2932 (N_2932,N_2884,N_2876);
nor U2933 (N_2933,N_2876,N_2874);
or U2934 (N_2934,N_2892,N_2887);
nand U2935 (N_2935,N_2894,N_2889);
or U2936 (N_2936,N_2875,N_2876);
or U2937 (N_2937,N_2895,N_2854);
and U2938 (N_2938,N_2871,N_2872);
nor U2939 (N_2939,N_2879,N_2860);
nand U2940 (N_2940,N_2889,N_2886);
and U2941 (N_2941,N_2898,N_2888);
nor U2942 (N_2942,N_2869,N_2889);
and U2943 (N_2943,N_2874,N_2852);
or U2944 (N_2944,N_2883,N_2880);
or U2945 (N_2945,N_2858,N_2878);
and U2946 (N_2946,N_2897,N_2886);
or U2947 (N_2947,N_2886,N_2856);
nand U2948 (N_2948,N_2864,N_2858);
xnor U2949 (N_2949,N_2850,N_2857);
or U2950 (N_2950,N_2945,N_2930);
nand U2951 (N_2951,N_2914,N_2943);
nand U2952 (N_2952,N_2909,N_2907);
nand U2953 (N_2953,N_2913,N_2924);
nand U2954 (N_2954,N_2927,N_2906);
nor U2955 (N_2955,N_2942,N_2901);
or U2956 (N_2956,N_2946,N_2949);
and U2957 (N_2957,N_2917,N_2918);
nand U2958 (N_2958,N_2934,N_2902);
and U2959 (N_2959,N_2926,N_2903);
nand U2960 (N_2960,N_2928,N_2939);
or U2961 (N_2961,N_2908,N_2941);
and U2962 (N_2962,N_2947,N_2938);
and U2963 (N_2963,N_2919,N_2915);
and U2964 (N_2964,N_2910,N_2944);
nor U2965 (N_2965,N_2933,N_2937);
nor U2966 (N_2966,N_2935,N_2904);
or U2967 (N_2967,N_2905,N_2922);
and U2968 (N_2968,N_2925,N_2911);
nor U2969 (N_2969,N_2936,N_2900);
and U2970 (N_2970,N_2921,N_2912);
or U2971 (N_2971,N_2932,N_2940);
nand U2972 (N_2972,N_2931,N_2929);
nor U2973 (N_2973,N_2920,N_2948);
and U2974 (N_2974,N_2916,N_2923);
nor U2975 (N_2975,N_2948,N_2933);
and U2976 (N_2976,N_2933,N_2925);
or U2977 (N_2977,N_2932,N_2927);
nand U2978 (N_2978,N_2946,N_2919);
nand U2979 (N_2979,N_2944,N_2936);
or U2980 (N_2980,N_2921,N_2948);
or U2981 (N_2981,N_2939,N_2922);
nor U2982 (N_2982,N_2909,N_2943);
or U2983 (N_2983,N_2929,N_2918);
and U2984 (N_2984,N_2910,N_2902);
nand U2985 (N_2985,N_2917,N_2901);
nor U2986 (N_2986,N_2939,N_2906);
nor U2987 (N_2987,N_2923,N_2947);
or U2988 (N_2988,N_2943,N_2947);
nand U2989 (N_2989,N_2926,N_2917);
nand U2990 (N_2990,N_2905,N_2948);
nor U2991 (N_2991,N_2906,N_2924);
or U2992 (N_2992,N_2947,N_2913);
and U2993 (N_2993,N_2915,N_2912);
nand U2994 (N_2994,N_2934,N_2915);
nor U2995 (N_2995,N_2904,N_2929);
and U2996 (N_2996,N_2923,N_2933);
nor U2997 (N_2997,N_2934,N_2903);
and U2998 (N_2998,N_2905,N_2919);
and U2999 (N_2999,N_2929,N_2944);
and UO_0 (O_0,N_2992,N_2989);
xnor UO_1 (O_1,N_2966,N_2963);
and UO_2 (O_2,N_2968,N_2976);
and UO_3 (O_3,N_2978,N_2956);
nand UO_4 (O_4,N_2981,N_2955);
nand UO_5 (O_5,N_2972,N_2991);
nor UO_6 (O_6,N_2983,N_2971);
and UO_7 (O_7,N_2977,N_2998);
nor UO_8 (O_8,N_2994,N_2984);
nor UO_9 (O_9,N_2999,N_2962);
and UO_10 (O_10,N_2973,N_2979);
and UO_11 (O_11,N_2960,N_2959);
or UO_12 (O_12,N_2974,N_2975);
and UO_13 (O_13,N_2950,N_2980);
and UO_14 (O_14,N_2985,N_2995);
xor UO_15 (O_15,N_2964,N_2969);
nand UO_16 (O_16,N_2951,N_2970);
and UO_17 (O_17,N_2958,N_2952);
or UO_18 (O_18,N_2953,N_2986);
or UO_19 (O_19,N_2954,N_2967);
nand UO_20 (O_20,N_2987,N_2997);
or UO_21 (O_21,N_2996,N_2961);
nand UO_22 (O_22,N_2990,N_2957);
nor UO_23 (O_23,N_2965,N_2988);
or UO_24 (O_24,N_2993,N_2982);
nand UO_25 (O_25,N_2968,N_2983);
nor UO_26 (O_26,N_2987,N_2991);
and UO_27 (O_27,N_2998,N_2997);
nor UO_28 (O_28,N_2957,N_2961);
nor UO_29 (O_29,N_2978,N_2952);
and UO_30 (O_30,N_2987,N_2967);
nor UO_31 (O_31,N_2969,N_2999);
nor UO_32 (O_32,N_2968,N_2991);
and UO_33 (O_33,N_2964,N_2983);
or UO_34 (O_34,N_2996,N_2990);
and UO_35 (O_35,N_2966,N_2950);
and UO_36 (O_36,N_2997,N_2958);
or UO_37 (O_37,N_2981,N_2976);
nor UO_38 (O_38,N_2986,N_2950);
and UO_39 (O_39,N_2961,N_2990);
or UO_40 (O_40,N_2974,N_2960);
and UO_41 (O_41,N_2957,N_2967);
and UO_42 (O_42,N_2961,N_2975);
and UO_43 (O_43,N_2999,N_2981);
or UO_44 (O_44,N_2971,N_2980);
or UO_45 (O_45,N_2978,N_2967);
nor UO_46 (O_46,N_2971,N_2968);
nand UO_47 (O_47,N_2994,N_2965);
and UO_48 (O_48,N_2992,N_2953);
and UO_49 (O_49,N_2976,N_2983);
nand UO_50 (O_50,N_2950,N_2970);
and UO_51 (O_51,N_2983,N_2996);
and UO_52 (O_52,N_2998,N_2951);
and UO_53 (O_53,N_2992,N_2979);
or UO_54 (O_54,N_2985,N_2972);
nor UO_55 (O_55,N_2979,N_2991);
or UO_56 (O_56,N_2961,N_2954);
and UO_57 (O_57,N_2989,N_2964);
and UO_58 (O_58,N_2974,N_2995);
or UO_59 (O_59,N_2981,N_2968);
and UO_60 (O_60,N_2983,N_2979);
nor UO_61 (O_61,N_2982,N_2952);
nand UO_62 (O_62,N_2960,N_2977);
nand UO_63 (O_63,N_2961,N_2974);
or UO_64 (O_64,N_2986,N_2993);
and UO_65 (O_65,N_2992,N_2955);
nor UO_66 (O_66,N_2987,N_2955);
nand UO_67 (O_67,N_2997,N_2976);
nand UO_68 (O_68,N_2994,N_2991);
and UO_69 (O_69,N_2977,N_2974);
and UO_70 (O_70,N_2987,N_2965);
nor UO_71 (O_71,N_2952,N_2994);
and UO_72 (O_72,N_2964,N_2968);
and UO_73 (O_73,N_2986,N_2961);
nand UO_74 (O_74,N_2974,N_2966);
nor UO_75 (O_75,N_2952,N_2996);
or UO_76 (O_76,N_2963,N_2954);
or UO_77 (O_77,N_2977,N_2965);
nor UO_78 (O_78,N_2982,N_2961);
and UO_79 (O_79,N_2961,N_2994);
nor UO_80 (O_80,N_2997,N_2985);
nand UO_81 (O_81,N_2991,N_2975);
nand UO_82 (O_82,N_2992,N_2968);
or UO_83 (O_83,N_2963,N_2985);
nand UO_84 (O_84,N_2996,N_2978);
nor UO_85 (O_85,N_2965,N_2953);
or UO_86 (O_86,N_2967,N_2956);
or UO_87 (O_87,N_2979,N_2960);
and UO_88 (O_88,N_2960,N_2956);
or UO_89 (O_89,N_2982,N_2973);
nand UO_90 (O_90,N_2958,N_2986);
and UO_91 (O_91,N_2971,N_2963);
nand UO_92 (O_92,N_2977,N_2966);
or UO_93 (O_93,N_2971,N_2981);
nand UO_94 (O_94,N_2994,N_2985);
or UO_95 (O_95,N_2997,N_2951);
or UO_96 (O_96,N_2994,N_2993);
or UO_97 (O_97,N_2975,N_2967);
nor UO_98 (O_98,N_2954,N_2998);
and UO_99 (O_99,N_2971,N_2986);
nand UO_100 (O_100,N_2983,N_2973);
and UO_101 (O_101,N_2956,N_2977);
nand UO_102 (O_102,N_2999,N_2963);
nor UO_103 (O_103,N_2997,N_2999);
and UO_104 (O_104,N_2995,N_2996);
or UO_105 (O_105,N_2985,N_2975);
nand UO_106 (O_106,N_2973,N_2960);
and UO_107 (O_107,N_2976,N_2979);
or UO_108 (O_108,N_2962,N_2965);
or UO_109 (O_109,N_2954,N_2984);
nor UO_110 (O_110,N_2984,N_2988);
nor UO_111 (O_111,N_2976,N_2960);
nor UO_112 (O_112,N_2984,N_2993);
nor UO_113 (O_113,N_2951,N_2982);
and UO_114 (O_114,N_2995,N_2954);
and UO_115 (O_115,N_2982,N_2995);
or UO_116 (O_116,N_2988,N_2957);
or UO_117 (O_117,N_2983,N_2966);
nand UO_118 (O_118,N_2984,N_2974);
nor UO_119 (O_119,N_2956,N_2955);
and UO_120 (O_120,N_2992,N_2960);
nand UO_121 (O_121,N_2963,N_2980);
nor UO_122 (O_122,N_2985,N_2959);
nand UO_123 (O_123,N_2967,N_2970);
nand UO_124 (O_124,N_2953,N_2984);
xnor UO_125 (O_125,N_2973,N_2980);
and UO_126 (O_126,N_2989,N_2954);
nor UO_127 (O_127,N_2954,N_2994);
nand UO_128 (O_128,N_2970,N_2961);
or UO_129 (O_129,N_2959,N_2997);
or UO_130 (O_130,N_2998,N_2953);
or UO_131 (O_131,N_2999,N_2965);
or UO_132 (O_132,N_2983,N_2978);
and UO_133 (O_133,N_2974,N_2993);
and UO_134 (O_134,N_2964,N_2974);
nor UO_135 (O_135,N_2967,N_2998);
nor UO_136 (O_136,N_2965,N_2978);
nor UO_137 (O_137,N_2973,N_2958);
or UO_138 (O_138,N_2958,N_2960);
or UO_139 (O_139,N_2955,N_2972);
nor UO_140 (O_140,N_2957,N_2969);
or UO_141 (O_141,N_2969,N_2987);
nor UO_142 (O_142,N_2997,N_2977);
and UO_143 (O_143,N_2979,N_2978);
nand UO_144 (O_144,N_2997,N_2950);
or UO_145 (O_145,N_2971,N_2960);
nand UO_146 (O_146,N_2952,N_2999);
nand UO_147 (O_147,N_2977,N_2996);
or UO_148 (O_148,N_2968,N_2998);
xnor UO_149 (O_149,N_2956,N_2983);
nand UO_150 (O_150,N_2992,N_2978);
nor UO_151 (O_151,N_2987,N_2951);
and UO_152 (O_152,N_2968,N_2954);
or UO_153 (O_153,N_2970,N_2957);
nand UO_154 (O_154,N_2959,N_2957);
nand UO_155 (O_155,N_2953,N_2979);
nand UO_156 (O_156,N_2969,N_2955);
and UO_157 (O_157,N_2987,N_2960);
nand UO_158 (O_158,N_2960,N_2969);
and UO_159 (O_159,N_2975,N_2969);
or UO_160 (O_160,N_2986,N_2960);
nor UO_161 (O_161,N_2982,N_2955);
nand UO_162 (O_162,N_2962,N_2960);
or UO_163 (O_163,N_2967,N_2982);
or UO_164 (O_164,N_2955,N_2976);
nor UO_165 (O_165,N_2955,N_2993);
or UO_166 (O_166,N_2966,N_2960);
and UO_167 (O_167,N_2967,N_2984);
and UO_168 (O_168,N_2953,N_2980);
nand UO_169 (O_169,N_2997,N_2983);
or UO_170 (O_170,N_2992,N_2997);
nor UO_171 (O_171,N_2991,N_2983);
or UO_172 (O_172,N_2982,N_2984);
or UO_173 (O_173,N_2999,N_2972);
or UO_174 (O_174,N_2963,N_2961);
nor UO_175 (O_175,N_2966,N_2982);
or UO_176 (O_176,N_2993,N_2963);
and UO_177 (O_177,N_2997,N_2956);
nor UO_178 (O_178,N_2994,N_2981);
and UO_179 (O_179,N_2979,N_2965);
or UO_180 (O_180,N_2968,N_2985);
nor UO_181 (O_181,N_2980,N_2990);
and UO_182 (O_182,N_2999,N_2966);
nand UO_183 (O_183,N_2961,N_2955);
and UO_184 (O_184,N_2990,N_2981);
nor UO_185 (O_185,N_2971,N_2982);
nand UO_186 (O_186,N_2986,N_2963);
nand UO_187 (O_187,N_2953,N_2985);
or UO_188 (O_188,N_2958,N_2985);
and UO_189 (O_189,N_2953,N_2951);
or UO_190 (O_190,N_2972,N_2967);
or UO_191 (O_191,N_2975,N_2986);
nor UO_192 (O_192,N_2983,N_2988);
nand UO_193 (O_193,N_2959,N_2995);
and UO_194 (O_194,N_2988,N_2954);
or UO_195 (O_195,N_2977,N_2951);
nor UO_196 (O_196,N_2958,N_2982);
nor UO_197 (O_197,N_2979,N_2996);
nor UO_198 (O_198,N_2958,N_2983);
and UO_199 (O_199,N_2993,N_2979);
nand UO_200 (O_200,N_2963,N_2982);
and UO_201 (O_201,N_2953,N_2963);
nand UO_202 (O_202,N_2990,N_2999);
nor UO_203 (O_203,N_2993,N_2991);
nand UO_204 (O_204,N_2996,N_2987);
or UO_205 (O_205,N_2966,N_2975);
and UO_206 (O_206,N_2996,N_2958);
and UO_207 (O_207,N_2992,N_2987);
and UO_208 (O_208,N_2975,N_2978);
or UO_209 (O_209,N_2951,N_2980);
nor UO_210 (O_210,N_2960,N_2994);
and UO_211 (O_211,N_2961,N_2980);
or UO_212 (O_212,N_2957,N_2977);
nand UO_213 (O_213,N_2996,N_2998);
and UO_214 (O_214,N_2954,N_2992);
or UO_215 (O_215,N_2971,N_2989);
and UO_216 (O_216,N_2975,N_2956);
and UO_217 (O_217,N_2973,N_2956);
nand UO_218 (O_218,N_2961,N_2968);
nand UO_219 (O_219,N_2969,N_2992);
nor UO_220 (O_220,N_2981,N_2974);
and UO_221 (O_221,N_2986,N_2982);
or UO_222 (O_222,N_2999,N_2977);
xnor UO_223 (O_223,N_2975,N_2998);
and UO_224 (O_224,N_2999,N_2992);
nor UO_225 (O_225,N_2971,N_2965);
xor UO_226 (O_226,N_2984,N_2992);
nor UO_227 (O_227,N_2982,N_2998);
nand UO_228 (O_228,N_2988,N_2955);
nor UO_229 (O_229,N_2960,N_2996);
or UO_230 (O_230,N_2963,N_2950);
and UO_231 (O_231,N_2956,N_2969);
or UO_232 (O_232,N_2974,N_2952);
and UO_233 (O_233,N_2996,N_2968);
nor UO_234 (O_234,N_2979,N_2950);
nor UO_235 (O_235,N_2989,N_2993);
nor UO_236 (O_236,N_2989,N_2977);
or UO_237 (O_237,N_2976,N_2980);
nand UO_238 (O_238,N_2977,N_2992);
or UO_239 (O_239,N_2980,N_2991);
and UO_240 (O_240,N_2985,N_2954);
and UO_241 (O_241,N_2979,N_2995);
or UO_242 (O_242,N_2994,N_2964);
and UO_243 (O_243,N_2963,N_2956);
nand UO_244 (O_244,N_2989,N_2999);
nand UO_245 (O_245,N_2972,N_2964);
or UO_246 (O_246,N_2986,N_2985);
or UO_247 (O_247,N_2973,N_2974);
nand UO_248 (O_248,N_2965,N_2969);
and UO_249 (O_249,N_2970,N_2965);
nor UO_250 (O_250,N_2963,N_2979);
nor UO_251 (O_251,N_2955,N_2985);
and UO_252 (O_252,N_2954,N_2991);
nor UO_253 (O_253,N_2973,N_2954);
and UO_254 (O_254,N_2987,N_2961);
or UO_255 (O_255,N_2966,N_2976);
nand UO_256 (O_256,N_2958,N_2971);
and UO_257 (O_257,N_2962,N_2961);
or UO_258 (O_258,N_2985,N_2970);
or UO_259 (O_259,N_2966,N_2970);
nand UO_260 (O_260,N_2992,N_2951);
or UO_261 (O_261,N_2964,N_2978);
and UO_262 (O_262,N_2954,N_2976);
or UO_263 (O_263,N_2982,N_2990);
or UO_264 (O_264,N_2979,N_2987);
or UO_265 (O_265,N_2963,N_2972);
nand UO_266 (O_266,N_2964,N_2971);
and UO_267 (O_267,N_2973,N_2972);
or UO_268 (O_268,N_2992,N_2991);
nor UO_269 (O_269,N_2971,N_2984);
and UO_270 (O_270,N_2986,N_2966);
and UO_271 (O_271,N_2981,N_2980);
or UO_272 (O_272,N_2954,N_2970);
nand UO_273 (O_273,N_2970,N_2963);
nand UO_274 (O_274,N_2958,N_2979);
and UO_275 (O_275,N_2984,N_2997);
nand UO_276 (O_276,N_2966,N_2981);
or UO_277 (O_277,N_2974,N_2968);
and UO_278 (O_278,N_2970,N_2969);
nor UO_279 (O_279,N_2981,N_2988);
nor UO_280 (O_280,N_2986,N_2994);
nor UO_281 (O_281,N_2984,N_2972);
or UO_282 (O_282,N_2972,N_2983);
and UO_283 (O_283,N_2964,N_2979);
or UO_284 (O_284,N_2950,N_2959);
or UO_285 (O_285,N_2998,N_2986);
and UO_286 (O_286,N_2976,N_2967);
and UO_287 (O_287,N_2994,N_2982);
nand UO_288 (O_288,N_2996,N_2966);
and UO_289 (O_289,N_2953,N_2954);
or UO_290 (O_290,N_2956,N_2964);
nand UO_291 (O_291,N_2990,N_2994);
and UO_292 (O_292,N_2953,N_2969);
nand UO_293 (O_293,N_2992,N_2957);
or UO_294 (O_294,N_2989,N_2994);
nor UO_295 (O_295,N_2976,N_2984);
nand UO_296 (O_296,N_2952,N_2984);
nand UO_297 (O_297,N_2976,N_2978);
nor UO_298 (O_298,N_2995,N_2991);
nor UO_299 (O_299,N_2995,N_2970);
and UO_300 (O_300,N_2986,N_2976);
nand UO_301 (O_301,N_2958,N_2965);
nor UO_302 (O_302,N_2989,N_2986);
or UO_303 (O_303,N_2997,N_2960);
and UO_304 (O_304,N_2984,N_2985);
nand UO_305 (O_305,N_2992,N_2982);
and UO_306 (O_306,N_2952,N_2964);
or UO_307 (O_307,N_2964,N_2963);
nand UO_308 (O_308,N_2994,N_2963);
and UO_309 (O_309,N_2981,N_2951);
nand UO_310 (O_310,N_2950,N_2967);
nand UO_311 (O_311,N_2964,N_2990);
and UO_312 (O_312,N_2994,N_2999);
nor UO_313 (O_313,N_2986,N_2957);
and UO_314 (O_314,N_2996,N_2957);
or UO_315 (O_315,N_2976,N_2996);
and UO_316 (O_316,N_2984,N_2978);
or UO_317 (O_317,N_2965,N_2968);
and UO_318 (O_318,N_2963,N_2957);
nand UO_319 (O_319,N_2982,N_2972);
and UO_320 (O_320,N_2961,N_2964);
nor UO_321 (O_321,N_2970,N_2955);
nor UO_322 (O_322,N_2955,N_2967);
nand UO_323 (O_323,N_2970,N_2974);
nand UO_324 (O_324,N_2998,N_2965);
or UO_325 (O_325,N_2995,N_2958);
or UO_326 (O_326,N_2975,N_2968);
and UO_327 (O_327,N_2970,N_2958);
and UO_328 (O_328,N_2994,N_2996);
nand UO_329 (O_329,N_2979,N_2972);
nand UO_330 (O_330,N_2984,N_2989);
or UO_331 (O_331,N_2989,N_2953);
nand UO_332 (O_332,N_2990,N_2951);
or UO_333 (O_333,N_2959,N_2994);
nor UO_334 (O_334,N_2993,N_2957);
nor UO_335 (O_335,N_2989,N_2969);
nor UO_336 (O_336,N_2952,N_2953);
nand UO_337 (O_337,N_2974,N_2953);
and UO_338 (O_338,N_2959,N_2996);
nand UO_339 (O_339,N_2995,N_2952);
nor UO_340 (O_340,N_2980,N_2977);
or UO_341 (O_341,N_2953,N_2959);
nand UO_342 (O_342,N_2996,N_2962);
or UO_343 (O_343,N_2981,N_2991);
xnor UO_344 (O_344,N_2966,N_2964);
nand UO_345 (O_345,N_2964,N_2954);
nand UO_346 (O_346,N_2981,N_2978);
nor UO_347 (O_347,N_2994,N_2976);
or UO_348 (O_348,N_2978,N_2989);
nor UO_349 (O_349,N_2960,N_2967);
nor UO_350 (O_350,N_2991,N_2953);
nand UO_351 (O_351,N_2998,N_2958);
and UO_352 (O_352,N_2976,N_2975);
and UO_353 (O_353,N_2993,N_2952);
nor UO_354 (O_354,N_2960,N_2982);
nor UO_355 (O_355,N_2960,N_2970);
or UO_356 (O_356,N_2956,N_2998);
nor UO_357 (O_357,N_2979,N_2999);
or UO_358 (O_358,N_2991,N_2989);
or UO_359 (O_359,N_2988,N_2974);
or UO_360 (O_360,N_2978,N_2950);
or UO_361 (O_361,N_2992,N_2958);
and UO_362 (O_362,N_2983,N_2967);
nand UO_363 (O_363,N_2957,N_2995);
nand UO_364 (O_364,N_2964,N_2998);
nor UO_365 (O_365,N_2979,N_2952);
xor UO_366 (O_366,N_2966,N_2951);
and UO_367 (O_367,N_2971,N_2975);
nor UO_368 (O_368,N_2956,N_2979);
xor UO_369 (O_369,N_2955,N_2971);
nor UO_370 (O_370,N_2995,N_2998);
nand UO_371 (O_371,N_2953,N_2966);
or UO_372 (O_372,N_2978,N_2968);
or UO_373 (O_373,N_2995,N_2987);
and UO_374 (O_374,N_2971,N_2954);
nor UO_375 (O_375,N_2984,N_2983);
or UO_376 (O_376,N_2990,N_2956);
or UO_377 (O_377,N_2988,N_2967);
and UO_378 (O_378,N_2964,N_2957);
nor UO_379 (O_379,N_2969,N_2994);
nor UO_380 (O_380,N_2965,N_2956);
or UO_381 (O_381,N_2986,N_2983);
and UO_382 (O_382,N_2981,N_2984);
and UO_383 (O_383,N_2960,N_2975);
and UO_384 (O_384,N_2990,N_2995);
or UO_385 (O_385,N_2977,N_2994);
nor UO_386 (O_386,N_2970,N_2998);
nand UO_387 (O_387,N_2958,N_2993);
and UO_388 (O_388,N_2990,N_2963);
or UO_389 (O_389,N_2974,N_2990);
and UO_390 (O_390,N_2973,N_2985);
or UO_391 (O_391,N_2981,N_2964);
or UO_392 (O_392,N_2977,N_2982);
nand UO_393 (O_393,N_2987,N_2950);
or UO_394 (O_394,N_2988,N_2972);
and UO_395 (O_395,N_2985,N_2952);
nand UO_396 (O_396,N_2961,N_2953);
or UO_397 (O_397,N_2975,N_2977);
and UO_398 (O_398,N_2955,N_2978);
nor UO_399 (O_399,N_2961,N_2973);
or UO_400 (O_400,N_2973,N_2953);
and UO_401 (O_401,N_2971,N_2976);
or UO_402 (O_402,N_2959,N_2965);
nor UO_403 (O_403,N_2961,N_2952);
nor UO_404 (O_404,N_2980,N_2978);
nor UO_405 (O_405,N_2974,N_2950);
or UO_406 (O_406,N_2994,N_2951);
and UO_407 (O_407,N_2984,N_2957);
or UO_408 (O_408,N_2982,N_2956);
nor UO_409 (O_409,N_2971,N_2951);
nor UO_410 (O_410,N_2994,N_2987);
and UO_411 (O_411,N_2967,N_2964);
nand UO_412 (O_412,N_2963,N_2984);
and UO_413 (O_413,N_2981,N_2970);
nand UO_414 (O_414,N_2968,N_2967);
nand UO_415 (O_415,N_2959,N_2992);
or UO_416 (O_416,N_2991,N_2970);
or UO_417 (O_417,N_2955,N_2965);
nor UO_418 (O_418,N_2975,N_2955);
or UO_419 (O_419,N_2995,N_2950);
or UO_420 (O_420,N_2960,N_2957);
nor UO_421 (O_421,N_2988,N_2971);
xor UO_422 (O_422,N_2988,N_2968);
and UO_423 (O_423,N_2957,N_2985);
nor UO_424 (O_424,N_2999,N_2996);
and UO_425 (O_425,N_2965,N_2976);
nand UO_426 (O_426,N_2959,N_2973);
or UO_427 (O_427,N_2967,N_2997);
nor UO_428 (O_428,N_2983,N_2961);
nand UO_429 (O_429,N_2978,N_2969);
or UO_430 (O_430,N_2955,N_2952);
nor UO_431 (O_431,N_2993,N_2996);
or UO_432 (O_432,N_2989,N_2979);
nand UO_433 (O_433,N_2970,N_2973);
or UO_434 (O_434,N_2982,N_2985);
nor UO_435 (O_435,N_2993,N_2983);
or UO_436 (O_436,N_2981,N_2958);
nor UO_437 (O_437,N_2971,N_2959);
or UO_438 (O_438,N_2950,N_2999);
nor UO_439 (O_439,N_2975,N_2952);
and UO_440 (O_440,N_2981,N_2992);
nand UO_441 (O_441,N_2990,N_2976);
and UO_442 (O_442,N_2951,N_2964);
nand UO_443 (O_443,N_2984,N_2987);
and UO_444 (O_444,N_2970,N_2980);
and UO_445 (O_445,N_2964,N_2988);
nor UO_446 (O_446,N_2998,N_2992);
nor UO_447 (O_447,N_2976,N_2964);
nand UO_448 (O_448,N_2987,N_2953);
or UO_449 (O_449,N_2952,N_2969);
nand UO_450 (O_450,N_2997,N_2953);
nor UO_451 (O_451,N_2957,N_2991);
nand UO_452 (O_452,N_2970,N_2983);
and UO_453 (O_453,N_2996,N_2972);
and UO_454 (O_454,N_2968,N_2959);
or UO_455 (O_455,N_2951,N_2979);
and UO_456 (O_456,N_2968,N_2995);
nor UO_457 (O_457,N_2954,N_2969);
and UO_458 (O_458,N_2963,N_2952);
nor UO_459 (O_459,N_2950,N_2981);
and UO_460 (O_460,N_2980,N_2998);
and UO_461 (O_461,N_2962,N_2988);
and UO_462 (O_462,N_2995,N_2969);
nor UO_463 (O_463,N_2965,N_2991);
nor UO_464 (O_464,N_2999,N_2956);
or UO_465 (O_465,N_2991,N_2951);
or UO_466 (O_466,N_2984,N_2956);
or UO_467 (O_467,N_2974,N_2955);
and UO_468 (O_468,N_2960,N_2993);
nand UO_469 (O_469,N_2985,N_2951);
nand UO_470 (O_470,N_2961,N_2992);
nand UO_471 (O_471,N_2994,N_2971);
or UO_472 (O_472,N_2957,N_2968);
or UO_473 (O_473,N_2973,N_2997);
and UO_474 (O_474,N_2976,N_2993);
nand UO_475 (O_475,N_2973,N_2992);
nor UO_476 (O_476,N_2972,N_2965);
or UO_477 (O_477,N_2955,N_2963);
and UO_478 (O_478,N_2963,N_2975);
nor UO_479 (O_479,N_2950,N_2953);
or UO_480 (O_480,N_2992,N_2974);
and UO_481 (O_481,N_2993,N_2962);
or UO_482 (O_482,N_2953,N_2972);
nand UO_483 (O_483,N_2988,N_2975);
or UO_484 (O_484,N_2960,N_2953);
and UO_485 (O_485,N_2970,N_2992);
or UO_486 (O_486,N_2991,N_2982);
or UO_487 (O_487,N_2959,N_2974);
nand UO_488 (O_488,N_2982,N_2999);
and UO_489 (O_489,N_2984,N_2980);
nand UO_490 (O_490,N_2990,N_2966);
or UO_491 (O_491,N_2989,N_2951);
and UO_492 (O_492,N_2999,N_2955);
or UO_493 (O_493,N_2997,N_2952);
or UO_494 (O_494,N_2973,N_2978);
nand UO_495 (O_495,N_2952,N_2962);
or UO_496 (O_496,N_2950,N_2969);
nand UO_497 (O_497,N_2973,N_2991);
or UO_498 (O_498,N_2975,N_2950);
nor UO_499 (O_499,N_2990,N_2971);
endmodule