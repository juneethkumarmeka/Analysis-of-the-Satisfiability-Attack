module basic_500_3000_500_50_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_306,In_102);
and U1 (N_1,In_307,In_473);
nand U2 (N_2,In_110,In_50);
nand U3 (N_3,In_321,In_212);
and U4 (N_4,In_340,In_484);
nor U5 (N_5,In_79,In_187);
or U6 (N_6,In_23,In_449);
and U7 (N_7,In_425,In_401);
nand U8 (N_8,In_165,In_278);
nor U9 (N_9,In_0,In_331);
and U10 (N_10,In_488,In_422);
or U11 (N_11,In_379,In_477);
nor U12 (N_12,In_43,In_471);
nand U13 (N_13,In_40,In_179);
nor U14 (N_14,In_494,In_103);
and U15 (N_15,In_497,In_465);
nor U16 (N_16,In_383,In_216);
nand U17 (N_17,In_341,In_227);
nor U18 (N_18,In_268,In_89);
nand U19 (N_19,In_262,In_34);
and U20 (N_20,In_226,In_352);
or U21 (N_21,In_232,In_83);
nor U22 (N_22,In_408,In_153);
nor U23 (N_23,In_418,In_255);
xor U24 (N_24,In_325,In_33);
or U25 (N_25,In_239,In_158);
nor U26 (N_26,In_339,In_120);
nor U27 (N_27,In_293,In_481);
and U28 (N_28,In_238,In_27);
or U29 (N_29,In_134,In_97);
and U30 (N_30,In_67,In_295);
nor U31 (N_31,In_461,In_439);
nor U32 (N_32,In_42,In_288);
and U33 (N_33,In_12,In_485);
and U34 (N_34,In_166,In_195);
and U35 (N_35,In_417,In_223);
nand U36 (N_36,In_265,In_73);
nand U37 (N_37,In_427,In_394);
or U38 (N_38,In_132,In_380);
nand U39 (N_39,In_184,In_263);
and U40 (N_40,In_200,In_244);
or U41 (N_41,In_354,In_470);
and U42 (N_42,In_302,In_324);
nor U43 (N_43,In_400,In_177);
xor U44 (N_44,In_234,In_186);
nand U45 (N_45,In_114,In_129);
or U46 (N_46,In_267,In_334);
nand U47 (N_47,In_447,In_251);
xnor U48 (N_48,In_61,In_317);
nand U49 (N_49,In_164,In_289);
nand U50 (N_50,In_453,In_6);
or U51 (N_51,In_296,In_361);
nor U52 (N_52,In_130,In_327);
nand U53 (N_53,In_346,In_249);
and U54 (N_54,In_190,In_229);
nor U55 (N_55,In_264,In_183);
or U56 (N_56,In_148,In_230);
nor U57 (N_57,In_491,In_57);
and U58 (N_58,In_330,In_241);
and U59 (N_59,In_141,In_377);
and U60 (N_60,In_256,In_31);
xor U61 (N_61,In_309,N_47);
nor U62 (N_62,In_434,In_133);
nand U63 (N_63,In_395,In_496);
or U64 (N_64,In_185,In_430);
nand U65 (N_65,In_273,In_174);
and U66 (N_66,In_448,N_44);
nand U67 (N_67,In_207,N_29);
xor U68 (N_68,In_71,In_328);
nor U69 (N_69,In_431,N_41);
nand U70 (N_70,In_369,In_192);
nand U71 (N_71,In_441,In_21);
nand U72 (N_72,In_113,In_245);
and U73 (N_73,In_146,In_45);
nand U74 (N_74,In_66,In_467);
and U75 (N_75,N_12,In_86);
nor U76 (N_76,In_364,In_105);
nor U77 (N_77,N_38,In_299);
and U78 (N_78,In_405,In_283);
and U79 (N_79,In_335,In_167);
nand U80 (N_80,In_106,In_32);
or U81 (N_81,In_301,In_26);
nor U82 (N_82,In_493,In_396);
nor U83 (N_83,In_135,In_161);
nand U84 (N_84,In_197,In_490);
nand U85 (N_85,In_478,In_108);
and U86 (N_86,In_47,In_281);
or U87 (N_87,In_193,N_49);
or U88 (N_88,In_305,In_53);
nand U89 (N_89,In_87,In_218);
and U90 (N_90,In_68,In_19);
nor U91 (N_91,N_28,In_14);
xnor U92 (N_92,In_440,In_5);
nand U93 (N_93,In_215,In_147);
and U94 (N_94,In_127,In_84);
nor U95 (N_95,In_49,In_419);
nor U96 (N_96,N_31,In_411);
nor U97 (N_97,N_56,In_140);
and U98 (N_98,In_112,In_390);
and U99 (N_99,In_287,N_54);
nand U100 (N_100,In_250,In_93);
and U101 (N_101,N_42,In_252);
nand U102 (N_102,In_107,N_36);
or U103 (N_103,In_428,In_367);
or U104 (N_104,In_266,In_65);
nor U105 (N_105,In_257,In_214);
and U106 (N_106,In_237,In_72);
nor U107 (N_107,In_286,In_414);
or U108 (N_108,In_259,In_372);
nand U109 (N_109,N_45,In_150);
nand U110 (N_110,In_55,In_423);
nor U111 (N_111,In_151,In_169);
nand U112 (N_112,In_450,N_24);
nor U113 (N_113,In_409,In_88);
or U114 (N_114,In_499,N_43);
and U115 (N_115,In_385,In_7);
nor U116 (N_116,In_378,In_208);
and U117 (N_117,N_33,In_445);
and U118 (N_118,In_204,In_253);
and U119 (N_119,In_209,In_355);
nand U120 (N_120,N_14,In_111);
and U121 (N_121,In_180,N_117);
nand U122 (N_122,N_87,In_122);
and U123 (N_123,In_375,In_78);
or U124 (N_124,N_15,In_155);
nand U125 (N_125,In_225,N_19);
or U126 (N_126,In_90,In_446);
nand U127 (N_127,In_480,In_443);
or U128 (N_128,N_16,N_1);
or U129 (N_129,In_402,N_77);
nand U130 (N_130,In_95,In_60);
and U131 (N_131,In_243,N_35);
nor U132 (N_132,N_32,In_432);
xnor U133 (N_133,In_152,In_13);
or U134 (N_134,In_397,In_76);
or U135 (N_135,N_7,In_85);
nor U136 (N_136,In_316,In_344);
nor U137 (N_137,In_189,In_362);
and U138 (N_138,In_349,In_9);
or U139 (N_139,In_292,In_435);
nor U140 (N_140,N_64,In_254);
or U141 (N_141,In_406,N_40);
and U142 (N_142,In_220,N_106);
nor U143 (N_143,In_366,In_476);
nand U144 (N_144,In_463,In_224);
nand U145 (N_145,In_365,In_81);
nand U146 (N_146,In_125,N_17);
and U147 (N_147,In_258,In_469);
nor U148 (N_148,N_109,In_415);
and U149 (N_149,In_269,N_60);
and U150 (N_150,In_137,In_194);
and U151 (N_151,In_157,In_462);
nor U152 (N_152,N_70,In_168);
or U153 (N_153,N_66,N_51);
nand U154 (N_154,In_222,N_62);
and U155 (N_155,In_454,N_108);
and U156 (N_156,In_11,N_2);
nor U157 (N_157,In_382,In_171);
xnor U158 (N_158,In_69,In_486);
xor U159 (N_159,N_5,In_8);
nor U160 (N_160,In_139,In_51);
xor U161 (N_161,In_178,In_343);
xor U162 (N_162,N_34,N_23);
nor U163 (N_163,In_272,N_90);
or U164 (N_164,In_119,In_18);
nand U165 (N_165,N_104,In_350);
or U166 (N_166,In_15,N_67);
nand U167 (N_167,In_2,In_199);
xor U168 (N_168,In_271,N_37);
and U169 (N_169,N_75,In_358);
nor U170 (N_170,In_466,N_85);
nand U171 (N_171,In_333,N_8);
and U172 (N_172,In_30,In_424);
nor U173 (N_173,In_464,In_381);
nor U174 (N_174,In_348,In_360);
or U175 (N_175,In_429,N_101);
and U176 (N_176,In_233,In_294);
nand U177 (N_177,N_11,In_246);
nor U178 (N_178,N_39,N_92);
nand U179 (N_179,In_22,In_48);
nand U180 (N_180,N_107,N_149);
or U181 (N_181,In_116,N_63);
nand U182 (N_182,In_458,In_74);
nor U183 (N_183,N_20,In_353);
nor U184 (N_184,N_155,In_159);
or U185 (N_185,N_154,In_181);
nand U186 (N_186,In_332,In_487);
nor U187 (N_187,N_158,In_459);
nand U188 (N_188,N_94,N_84);
nor U189 (N_189,In_38,In_96);
xnor U190 (N_190,In_456,In_303);
or U191 (N_191,In_176,In_421);
and U192 (N_192,In_94,In_160);
and U193 (N_193,In_436,In_475);
or U194 (N_194,In_202,N_150);
or U195 (N_195,In_16,In_247);
or U196 (N_196,N_141,In_373);
nand U197 (N_197,N_55,In_211);
nor U198 (N_198,In_115,In_138);
nor U199 (N_199,N_91,In_392);
nor U200 (N_200,In_280,In_489);
and U201 (N_201,In_70,In_210);
nand U202 (N_202,In_175,N_112);
or U203 (N_203,N_152,In_426);
nor U204 (N_204,In_314,N_153);
nor U205 (N_205,In_279,In_117);
and U206 (N_206,In_20,In_104);
or U207 (N_207,N_80,N_166);
and U208 (N_208,In_498,In_154);
xnor U209 (N_209,In_410,N_126);
and U210 (N_210,N_74,In_35);
and U211 (N_211,N_100,N_13);
and U212 (N_212,N_82,N_122);
nand U213 (N_213,N_103,In_326);
nand U214 (N_214,In_438,In_10);
xor U215 (N_215,In_329,In_144);
xnor U216 (N_216,N_118,In_98);
or U217 (N_217,N_146,In_201);
nor U218 (N_218,N_105,In_17);
nand U219 (N_219,In_39,N_137);
nor U220 (N_220,In_101,In_322);
and U221 (N_221,N_140,N_79);
or U222 (N_222,In_455,In_124);
xor U223 (N_223,In_374,N_179);
and U224 (N_224,N_102,N_88);
nor U225 (N_225,In_219,N_26);
or U226 (N_226,In_228,N_21);
or U227 (N_227,N_65,In_393);
nand U228 (N_228,N_9,In_3);
nand U229 (N_229,N_22,In_345);
and U230 (N_230,In_313,In_203);
and U231 (N_231,In_261,In_356);
xor U232 (N_232,In_196,In_320);
nand U233 (N_233,N_124,In_1);
and U234 (N_234,N_10,N_99);
nand U235 (N_235,N_156,In_315);
nand U236 (N_236,N_68,N_125);
nand U237 (N_237,In_276,In_433);
nand U238 (N_238,N_162,In_444);
or U239 (N_239,N_95,In_297);
nand U240 (N_240,N_160,N_186);
nand U241 (N_241,N_131,In_310);
nand U242 (N_242,N_224,In_99);
or U243 (N_243,In_172,In_59);
nand U244 (N_244,N_190,N_3);
or U245 (N_245,In_347,N_235);
nor U246 (N_246,N_201,N_114);
or U247 (N_247,N_239,In_145);
and U248 (N_248,N_157,In_300);
nand U249 (N_249,N_143,N_116);
nor U250 (N_250,In_109,In_357);
xor U251 (N_251,N_130,In_275);
nand U252 (N_252,N_217,In_451);
nor U253 (N_253,N_227,In_36);
or U254 (N_254,In_318,N_76);
nand U255 (N_255,N_236,In_77);
nor U256 (N_256,In_304,In_25);
and U257 (N_257,In_391,In_170);
xnor U258 (N_258,In_285,N_208);
and U259 (N_259,N_98,In_217);
or U260 (N_260,In_404,N_192);
and U261 (N_261,In_290,N_232);
nand U262 (N_262,N_178,In_62);
nor U263 (N_263,In_136,In_311);
nand U264 (N_264,N_61,N_238);
nor U265 (N_265,In_363,N_191);
or U266 (N_266,N_182,N_188);
nor U267 (N_267,N_48,In_338);
nor U268 (N_268,N_71,In_270);
nand U269 (N_269,N_198,N_168);
xor U270 (N_270,N_119,In_231);
nor U271 (N_271,N_110,N_207);
nor U272 (N_272,N_73,N_225);
xnor U273 (N_273,In_75,N_237);
nand U274 (N_274,N_53,N_212);
nand U275 (N_275,In_128,In_56);
and U276 (N_276,In_221,In_442);
nand U277 (N_277,In_495,In_323);
nor U278 (N_278,N_4,N_58);
and U279 (N_279,N_194,In_319);
or U280 (N_280,N_195,In_420);
or U281 (N_281,In_492,In_389);
or U282 (N_282,N_144,N_229);
or U283 (N_283,In_82,In_118);
nand U284 (N_284,N_133,N_230);
or U285 (N_285,N_214,N_215);
nand U286 (N_286,In_437,N_142);
and U287 (N_287,In_205,In_121);
xnor U288 (N_288,N_210,In_58);
and U289 (N_289,N_181,In_123);
xnor U290 (N_290,N_89,N_211);
and U291 (N_291,In_368,In_398);
nand U292 (N_292,N_121,N_128);
xor U293 (N_293,In_162,N_204);
or U294 (N_294,In_399,N_127);
and U295 (N_295,In_468,N_30);
or U296 (N_296,In_359,In_188);
or U297 (N_297,In_198,In_92);
nor U298 (N_298,In_483,N_174);
nand U299 (N_299,In_191,N_197);
or U300 (N_300,In_386,In_28);
and U301 (N_301,N_72,N_187);
and U302 (N_302,N_281,In_182);
nor U303 (N_303,N_163,In_142);
xor U304 (N_304,In_173,N_97);
and U305 (N_305,N_250,In_291);
nand U306 (N_306,N_280,N_171);
and U307 (N_307,N_193,In_284);
and U308 (N_308,N_289,N_298);
nand U309 (N_309,N_96,In_384);
nor U310 (N_310,N_252,N_245);
or U311 (N_311,N_284,N_297);
and U312 (N_312,N_249,N_203);
nor U313 (N_313,In_308,In_298);
and U314 (N_314,N_172,In_312);
xnor U315 (N_315,N_136,N_129);
or U316 (N_316,In_388,N_205);
xor U317 (N_317,N_282,N_81);
and U318 (N_318,N_57,N_279);
or U319 (N_319,N_180,N_287);
nor U320 (N_320,In_143,In_412);
nor U321 (N_321,In_479,In_63);
nor U322 (N_322,N_138,N_169);
or U323 (N_323,N_164,In_387);
nand U324 (N_324,N_111,N_233);
nand U325 (N_325,N_220,N_285);
nor U326 (N_326,N_202,N_256);
nand U327 (N_327,N_216,In_371);
and U328 (N_328,In_100,In_274);
xor U329 (N_329,N_199,In_240);
nand U330 (N_330,In_407,N_242);
nor U331 (N_331,N_196,N_243);
xor U332 (N_332,In_41,In_126);
xor U333 (N_333,In_416,N_254);
nand U334 (N_334,N_228,N_148);
nor U335 (N_335,N_52,N_176);
and U336 (N_336,N_231,In_351);
and U337 (N_337,In_46,N_290);
nor U338 (N_338,In_4,N_135);
nor U339 (N_339,In_54,N_286);
and U340 (N_340,N_253,N_261);
nand U341 (N_341,N_273,In_376);
nor U342 (N_342,In_213,N_184);
nand U343 (N_343,N_183,N_167);
or U344 (N_344,In_242,N_161);
and U345 (N_345,N_267,In_156);
nand U346 (N_346,N_266,N_264);
and U347 (N_347,N_278,N_132);
nor U348 (N_348,In_64,N_222);
xnor U349 (N_349,N_173,N_270);
and U350 (N_350,N_218,N_275);
or U351 (N_351,N_283,In_403);
and U352 (N_352,N_200,N_259);
nor U353 (N_353,In_457,N_291);
nor U354 (N_354,N_296,N_288);
nand U355 (N_355,N_206,In_282);
nand U356 (N_356,N_293,In_91);
nor U357 (N_357,N_113,N_147);
xor U358 (N_358,N_134,N_139);
nor U359 (N_359,N_299,N_59);
nor U360 (N_360,N_265,N_226);
nor U361 (N_361,N_46,In_131);
and U362 (N_362,In_370,In_277);
nor U363 (N_363,In_413,N_348);
nor U364 (N_364,N_274,N_347);
nand U365 (N_365,N_340,N_294);
or U366 (N_366,In_337,N_349);
and U367 (N_367,N_342,N_336);
and U368 (N_368,N_268,N_316);
nor U369 (N_369,In_460,N_170);
nand U370 (N_370,In_452,N_159);
nand U371 (N_371,N_241,N_328);
or U372 (N_372,N_25,N_258);
nand U373 (N_373,N_359,N_120);
nor U374 (N_374,N_346,N_326);
nand U375 (N_375,N_318,N_272);
or U376 (N_376,N_27,N_248);
and U377 (N_377,N_308,In_52);
and U378 (N_378,N_317,In_342);
nand U379 (N_379,N_123,N_300);
and U380 (N_380,N_78,N_86);
nand U381 (N_381,N_93,N_337);
nand U382 (N_382,N_358,N_304);
nand U383 (N_383,N_330,N_309);
or U384 (N_384,In_482,N_312);
or U385 (N_385,In_149,N_83);
and U386 (N_386,In_472,N_177);
and U387 (N_387,N_314,N_351);
nand U388 (N_388,N_315,N_246);
nand U389 (N_389,N_276,N_352);
nor U390 (N_390,N_310,N_319);
and U391 (N_391,In_336,N_321);
or U392 (N_392,N_354,In_248);
xnor U393 (N_393,N_175,N_357);
xor U394 (N_394,N_247,N_185);
nor U395 (N_395,N_341,N_292);
nor U396 (N_396,N_353,N_257);
and U397 (N_397,N_165,N_344);
xnor U398 (N_398,In_235,N_302);
and U399 (N_399,N_311,N_271);
nand U400 (N_400,N_145,N_322);
or U401 (N_401,N_221,N_189);
nor U402 (N_402,N_334,N_307);
nand U403 (N_403,In_163,N_305);
and U404 (N_404,N_327,N_223);
nor U405 (N_405,In_236,N_295);
nor U406 (N_406,N_18,N_269);
nand U407 (N_407,N_255,N_325);
and U408 (N_408,N_338,N_350);
nor U409 (N_409,N_356,N_219);
xor U410 (N_410,N_0,N_277);
nor U411 (N_411,N_151,N_244);
nor U412 (N_412,In_260,In_474);
nor U413 (N_413,N_115,N_234);
or U414 (N_414,N_306,N_333);
or U415 (N_415,N_332,N_262);
and U416 (N_416,N_343,N_6);
nor U417 (N_417,N_339,N_263);
nor U418 (N_418,N_320,N_303);
nor U419 (N_419,N_301,N_50);
xnor U420 (N_420,N_401,N_395);
nor U421 (N_421,N_406,N_376);
and U422 (N_422,N_384,In_37);
or U423 (N_423,In_24,N_209);
xnor U424 (N_424,N_407,N_411);
nand U425 (N_425,N_355,N_398);
or U426 (N_426,N_417,N_367);
nand U427 (N_427,N_372,N_380);
and U428 (N_428,N_331,N_360);
and U429 (N_429,N_324,N_379);
nor U430 (N_430,N_385,N_368);
or U431 (N_431,N_418,N_397);
nand U432 (N_432,N_390,N_388);
and U433 (N_433,N_365,N_323);
or U434 (N_434,In_44,N_394);
nand U435 (N_435,N_329,N_313);
nand U436 (N_436,N_412,N_260);
and U437 (N_437,N_369,N_362);
and U438 (N_438,N_387,N_382);
nor U439 (N_439,N_374,N_363);
nor U440 (N_440,N_371,N_345);
or U441 (N_441,N_213,N_392);
nand U442 (N_442,N_383,N_240);
nor U443 (N_443,N_378,N_419);
and U444 (N_444,N_409,N_400);
and U445 (N_445,N_405,In_206);
or U446 (N_446,N_381,N_396);
nor U447 (N_447,N_415,N_361);
nand U448 (N_448,N_391,N_377);
and U449 (N_449,N_251,N_410);
and U450 (N_450,N_69,N_402);
nor U451 (N_451,N_404,N_389);
or U452 (N_452,In_80,N_403);
or U453 (N_453,N_375,N_366);
and U454 (N_454,N_370,N_413);
xor U455 (N_455,N_364,N_335);
xor U456 (N_456,N_416,N_393);
xor U457 (N_457,N_386,N_399);
or U458 (N_458,N_408,N_373);
nor U459 (N_459,In_29,N_414);
xnor U460 (N_460,N_392,N_406);
nand U461 (N_461,N_379,N_373);
nor U462 (N_462,N_394,N_390);
nand U463 (N_463,N_389,N_393);
xnor U464 (N_464,N_368,N_362);
or U465 (N_465,N_383,N_412);
and U466 (N_466,N_313,N_386);
or U467 (N_467,N_386,N_390);
or U468 (N_468,In_206,N_213);
and U469 (N_469,N_375,N_323);
nand U470 (N_470,N_390,N_360);
or U471 (N_471,N_403,N_382);
and U472 (N_472,N_401,N_393);
nor U473 (N_473,N_380,N_403);
nand U474 (N_474,N_418,N_400);
or U475 (N_475,In_24,N_394);
or U476 (N_476,N_360,N_371);
and U477 (N_477,In_80,N_410);
nor U478 (N_478,N_366,N_398);
nand U479 (N_479,N_260,N_415);
or U480 (N_480,N_432,N_473);
nand U481 (N_481,N_428,N_467);
and U482 (N_482,N_475,N_457);
or U483 (N_483,N_466,N_460);
nor U484 (N_484,N_453,N_440);
and U485 (N_485,N_459,N_436);
nand U486 (N_486,N_464,N_465);
xnor U487 (N_487,N_423,N_433);
nand U488 (N_488,N_437,N_448);
nand U489 (N_489,N_449,N_450);
or U490 (N_490,N_420,N_471);
nor U491 (N_491,N_474,N_458);
nand U492 (N_492,N_454,N_421);
and U493 (N_493,N_463,N_447);
nand U494 (N_494,N_429,N_435);
nand U495 (N_495,N_442,N_426);
nor U496 (N_496,N_476,N_446);
xor U497 (N_497,N_456,N_430);
nor U498 (N_498,N_439,N_472);
nand U499 (N_499,N_431,N_427);
and U500 (N_500,N_478,N_477);
nand U501 (N_501,N_443,N_424);
nor U502 (N_502,N_468,N_438);
nor U503 (N_503,N_441,N_455);
nor U504 (N_504,N_434,N_444);
nor U505 (N_505,N_479,N_461);
or U506 (N_506,N_451,N_470);
or U507 (N_507,N_469,N_445);
nand U508 (N_508,N_452,N_462);
and U509 (N_509,N_422,N_425);
nor U510 (N_510,N_434,N_445);
and U511 (N_511,N_439,N_465);
and U512 (N_512,N_460,N_444);
or U513 (N_513,N_438,N_456);
nand U514 (N_514,N_457,N_449);
or U515 (N_515,N_466,N_421);
nand U516 (N_516,N_444,N_458);
xor U517 (N_517,N_428,N_433);
or U518 (N_518,N_420,N_472);
nand U519 (N_519,N_433,N_425);
or U520 (N_520,N_469,N_436);
xnor U521 (N_521,N_451,N_469);
xor U522 (N_522,N_434,N_452);
or U523 (N_523,N_426,N_479);
nor U524 (N_524,N_465,N_444);
or U525 (N_525,N_474,N_444);
or U526 (N_526,N_458,N_455);
and U527 (N_527,N_472,N_436);
or U528 (N_528,N_462,N_461);
xnor U529 (N_529,N_440,N_425);
and U530 (N_530,N_443,N_461);
nand U531 (N_531,N_444,N_424);
and U532 (N_532,N_423,N_424);
nor U533 (N_533,N_475,N_474);
and U534 (N_534,N_456,N_440);
nand U535 (N_535,N_447,N_474);
xor U536 (N_536,N_450,N_476);
nand U537 (N_537,N_434,N_473);
and U538 (N_538,N_461,N_424);
nor U539 (N_539,N_456,N_461);
nor U540 (N_540,N_515,N_513);
or U541 (N_541,N_534,N_537);
nand U542 (N_542,N_539,N_494);
nand U543 (N_543,N_503,N_530);
nand U544 (N_544,N_493,N_521);
nand U545 (N_545,N_505,N_499);
or U546 (N_546,N_510,N_520);
nor U547 (N_547,N_526,N_514);
nand U548 (N_548,N_496,N_490);
nor U549 (N_549,N_538,N_501);
or U550 (N_550,N_532,N_516);
and U551 (N_551,N_535,N_506);
xnor U552 (N_552,N_487,N_500);
nor U553 (N_553,N_507,N_486);
or U554 (N_554,N_517,N_483);
nand U555 (N_555,N_485,N_480);
nor U556 (N_556,N_528,N_529);
xnor U557 (N_557,N_533,N_504);
nor U558 (N_558,N_482,N_492);
xor U559 (N_559,N_523,N_495);
or U560 (N_560,N_509,N_488);
or U561 (N_561,N_511,N_525);
or U562 (N_562,N_481,N_522);
or U563 (N_563,N_518,N_508);
or U564 (N_564,N_519,N_531);
nor U565 (N_565,N_536,N_498);
or U566 (N_566,N_491,N_497);
xnor U567 (N_567,N_524,N_512);
nand U568 (N_568,N_527,N_489);
or U569 (N_569,N_484,N_502);
nand U570 (N_570,N_507,N_504);
nor U571 (N_571,N_526,N_500);
or U572 (N_572,N_532,N_510);
nand U573 (N_573,N_520,N_533);
nor U574 (N_574,N_493,N_494);
nand U575 (N_575,N_494,N_496);
nand U576 (N_576,N_514,N_535);
nor U577 (N_577,N_528,N_539);
nor U578 (N_578,N_493,N_517);
xnor U579 (N_579,N_494,N_513);
or U580 (N_580,N_486,N_537);
nand U581 (N_581,N_516,N_529);
nor U582 (N_582,N_518,N_486);
and U583 (N_583,N_517,N_484);
nor U584 (N_584,N_499,N_487);
nand U585 (N_585,N_529,N_489);
or U586 (N_586,N_539,N_495);
nor U587 (N_587,N_493,N_524);
and U588 (N_588,N_511,N_488);
or U589 (N_589,N_496,N_518);
xor U590 (N_590,N_480,N_513);
nand U591 (N_591,N_535,N_526);
nand U592 (N_592,N_502,N_486);
or U593 (N_593,N_487,N_484);
or U594 (N_594,N_519,N_503);
or U595 (N_595,N_494,N_500);
and U596 (N_596,N_496,N_516);
and U597 (N_597,N_510,N_538);
or U598 (N_598,N_497,N_488);
nor U599 (N_599,N_490,N_513);
xnor U600 (N_600,N_561,N_593);
or U601 (N_601,N_568,N_596);
and U602 (N_602,N_544,N_583);
nor U603 (N_603,N_577,N_575);
or U604 (N_604,N_548,N_592);
nor U605 (N_605,N_584,N_550);
nor U606 (N_606,N_576,N_570);
nand U607 (N_607,N_557,N_552);
or U608 (N_608,N_573,N_572);
nor U609 (N_609,N_541,N_587);
nor U610 (N_610,N_569,N_595);
or U611 (N_611,N_560,N_566);
nand U612 (N_612,N_597,N_551);
or U613 (N_613,N_554,N_546);
or U614 (N_614,N_574,N_591);
or U615 (N_615,N_564,N_571);
nand U616 (N_616,N_599,N_565);
nand U617 (N_617,N_578,N_567);
or U618 (N_618,N_553,N_562);
xor U619 (N_619,N_549,N_594);
nor U620 (N_620,N_590,N_589);
or U621 (N_621,N_547,N_563);
nor U622 (N_622,N_585,N_588);
nand U623 (N_623,N_582,N_542);
nor U624 (N_624,N_586,N_545);
nor U625 (N_625,N_543,N_581);
or U626 (N_626,N_558,N_556);
or U627 (N_627,N_555,N_598);
or U628 (N_628,N_579,N_580);
xnor U629 (N_629,N_559,N_540);
nor U630 (N_630,N_589,N_542);
or U631 (N_631,N_579,N_581);
and U632 (N_632,N_576,N_598);
nor U633 (N_633,N_567,N_575);
and U634 (N_634,N_547,N_551);
or U635 (N_635,N_555,N_552);
and U636 (N_636,N_545,N_548);
nand U637 (N_637,N_591,N_571);
nand U638 (N_638,N_562,N_550);
xnor U639 (N_639,N_558,N_551);
xor U640 (N_640,N_561,N_560);
nor U641 (N_641,N_556,N_549);
or U642 (N_642,N_572,N_562);
or U643 (N_643,N_594,N_558);
nand U644 (N_644,N_594,N_593);
or U645 (N_645,N_560,N_542);
and U646 (N_646,N_578,N_545);
nand U647 (N_647,N_566,N_555);
or U648 (N_648,N_583,N_553);
xnor U649 (N_649,N_551,N_580);
nand U650 (N_650,N_544,N_592);
nand U651 (N_651,N_553,N_599);
or U652 (N_652,N_577,N_593);
or U653 (N_653,N_542,N_550);
or U654 (N_654,N_563,N_579);
and U655 (N_655,N_594,N_578);
nor U656 (N_656,N_574,N_575);
and U657 (N_657,N_549,N_563);
or U658 (N_658,N_564,N_543);
nor U659 (N_659,N_562,N_589);
nor U660 (N_660,N_637,N_631);
or U661 (N_661,N_656,N_622);
or U662 (N_662,N_620,N_629);
xnor U663 (N_663,N_623,N_614);
and U664 (N_664,N_601,N_638);
nor U665 (N_665,N_617,N_618);
nand U666 (N_666,N_652,N_628);
nor U667 (N_667,N_605,N_610);
or U668 (N_668,N_619,N_654);
or U669 (N_669,N_602,N_609);
and U670 (N_670,N_648,N_657);
nand U671 (N_671,N_607,N_604);
nor U672 (N_672,N_646,N_659);
and U673 (N_673,N_608,N_645);
nor U674 (N_674,N_634,N_653);
or U675 (N_675,N_635,N_658);
nand U676 (N_676,N_616,N_650);
or U677 (N_677,N_651,N_643);
and U678 (N_678,N_642,N_632);
and U679 (N_679,N_621,N_649);
nand U680 (N_680,N_647,N_611);
nor U681 (N_681,N_600,N_644);
and U682 (N_682,N_615,N_606);
nor U683 (N_683,N_639,N_633);
or U684 (N_684,N_655,N_613);
nand U685 (N_685,N_626,N_627);
nor U686 (N_686,N_625,N_603);
and U687 (N_687,N_641,N_630);
xnor U688 (N_688,N_612,N_636);
or U689 (N_689,N_624,N_640);
or U690 (N_690,N_600,N_654);
nand U691 (N_691,N_650,N_654);
and U692 (N_692,N_655,N_645);
nor U693 (N_693,N_636,N_656);
and U694 (N_694,N_611,N_639);
nand U695 (N_695,N_625,N_657);
nand U696 (N_696,N_625,N_616);
and U697 (N_697,N_625,N_628);
nand U698 (N_698,N_613,N_659);
xnor U699 (N_699,N_602,N_612);
and U700 (N_700,N_632,N_646);
nor U701 (N_701,N_609,N_647);
nand U702 (N_702,N_625,N_645);
or U703 (N_703,N_631,N_610);
or U704 (N_704,N_655,N_650);
nand U705 (N_705,N_633,N_648);
nor U706 (N_706,N_602,N_652);
and U707 (N_707,N_611,N_654);
nor U708 (N_708,N_610,N_601);
and U709 (N_709,N_637,N_634);
or U710 (N_710,N_647,N_618);
nor U711 (N_711,N_626,N_657);
nand U712 (N_712,N_648,N_656);
nor U713 (N_713,N_650,N_606);
nand U714 (N_714,N_621,N_628);
nand U715 (N_715,N_618,N_606);
and U716 (N_716,N_647,N_629);
xor U717 (N_717,N_611,N_613);
or U718 (N_718,N_639,N_600);
and U719 (N_719,N_628,N_611);
nand U720 (N_720,N_667,N_684);
and U721 (N_721,N_710,N_686);
nand U722 (N_722,N_707,N_692);
and U723 (N_723,N_680,N_699);
nor U724 (N_724,N_674,N_683);
nor U725 (N_725,N_678,N_719);
nor U726 (N_726,N_698,N_660);
and U727 (N_727,N_677,N_671);
or U728 (N_728,N_704,N_670);
or U729 (N_729,N_688,N_718);
xor U730 (N_730,N_664,N_702);
or U731 (N_731,N_703,N_666);
nand U732 (N_732,N_714,N_690);
nand U733 (N_733,N_705,N_717);
nand U734 (N_734,N_691,N_685);
xnor U735 (N_735,N_715,N_661);
nand U736 (N_736,N_687,N_700);
and U737 (N_737,N_713,N_712);
nor U738 (N_738,N_663,N_708);
nand U739 (N_739,N_701,N_716);
nor U740 (N_740,N_711,N_706);
or U741 (N_741,N_693,N_681);
nor U742 (N_742,N_669,N_668);
and U743 (N_743,N_665,N_689);
xnor U744 (N_744,N_695,N_675);
and U745 (N_745,N_662,N_697);
nand U746 (N_746,N_679,N_696);
or U747 (N_747,N_676,N_682);
or U748 (N_748,N_709,N_672);
or U749 (N_749,N_673,N_694);
xor U750 (N_750,N_700,N_675);
and U751 (N_751,N_711,N_705);
nand U752 (N_752,N_689,N_668);
nand U753 (N_753,N_675,N_660);
or U754 (N_754,N_669,N_679);
xnor U755 (N_755,N_710,N_661);
and U756 (N_756,N_687,N_694);
nand U757 (N_757,N_716,N_672);
xnor U758 (N_758,N_717,N_703);
and U759 (N_759,N_706,N_697);
or U760 (N_760,N_711,N_698);
and U761 (N_761,N_692,N_718);
nor U762 (N_762,N_704,N_676);
nor U763 (N_763,N_663,N_660);
and U764 (N_764,N_709,N_682);
or U765 (N_765,N_662,N_667);
and U766 (N_766,N_705,N_703);
or U767 (N_767,N_686,N_674);
nand U768 (N_768,N_690,N_677);
nor U769 (N_769,N_682,N_693);
nand U770 (N_770,N_677,N_685);
nand U771 (N_771,N_677,N_694);
nand U772 (N_772,N_718,N_691);
nor U773 (N_773,N_712,N_663);
nand U774 (N_774,N_702,N_697);
nand U775 (N_775,N_706,N_687);
and U776 (N_776,N_679,N_695);
and U777 (N_777,N_701,N_679);
xor U778 (N_778,N_663,N_686);
nor U779 (N_779,N_665,N_675);
and U780 (N_780,N_765,N_762);
or U781 (N_781,N_774,N_734);
and U782 (N_782,N_771,N_777);
nor U783 (N_783,N_773,N_729);
nand U784 (N_784,N_741,N_730);
nor U785 (N_785,N_721,N_749);
nor U786 (N_786,N_767,N_740);
xor U787 (N_787,N_776,N_779);
or U788 (N_788,N_723,N_739);
and U789 (N_789,N_770,N_733);
nand U790 (N_790,N_735,N_768);
nor U791 (N_791,N_759,N_750);
or U792 (N_792,N_736,N_756);
or U793 (N_793,N_752,N_772);
nand U794 (N_794,N_763,N_743);
or U795 (N_795,N_764,N_722);
nand U796 (N_796,N_720,N_747);
and U797 (N_797,N_737,N_742);
and U798 (N_798,N_744,N_758);
nor U799 (N_799,N_754,N_766);
nor U800 (N_800,N_755,N_724);
nand U801 (N_801,N_728,N_727);
nand U802 (N_802,N_731,N_753);
nor U803 (N_803,N_748,N_760);
xor U804 (N_804,N_726,N_746);
and U805 (N_805,N_757,N_732);
nand U806 (N_806,N_769,N_745);
xnor U807 (N_807,N_778,N_738);
xnor U808 (N_808,N_775,N_751);
and U809 (N_809,N_725,N_761);
and U810 (N_810,N_745,N_755);
and U811 (N_811,N_742,N_731);
and U812 (N_812,N_729,N_762);
nor U813 (N_813,N_765,N_731);
or U814 (N_814,N_776,N_772);
nand U815 (N_815,N_779,N_771);
or U816 (N_816,N_748,N_750);
and U817 (N_817,N_730,N_751);
nand U818 (N_818,N_721,N_728);
or U819 (N_819,N_778,N_763);
nand U820 (N_820,N_720,N_778);
and U821 (N_821,N_735,N_772);
nor U822 (N_822,N_766,N_749);
or U823 (N_823,N_729,N_730);
nor U824 (N_824,N_774,N_732);
nand U825 (N_825,N_761,N_757);
and U826 (N_826,N_727,N_766);
or U827 (N_827,N_756,N_723);
nand U828 (N_828,N_761,N_763);
and U829 (N_829,N_736,N_721);
nand U830 (N_830,N_752,N_736);
nand U831 (N_831,N_739,N_770);
nor U832 (N_832,N_758,N_771);
xor U833 (N_833,N_754,N_748);
and U834 (N_834,N_751,N_733);
and U835 (N_835,N_779,N_732);
or U836 (N_836,N_752,N_723);
nor U837 (N_837,N_724,N_749);
or U838 (N_838,N_745,N_743);
nand U839 (N_839,N_774,N_751);
or U840 (N_840,N_786,N_789);
nand U841 (N_841,N_821,N_785);
nand U842 (N_842,N_835,N_819);
and U843 (N_843,N_802,N_823);
or U844 (N_844,N_797,N_799);
or U845 (N_845,N_811,N_836);
xor U846 (N_846,N_814,N_804);
nor U847 (N_847,N_818,N_801);
nand U848 (N_848,N_792,N_787);
and U849 (N_849,N_817,N_838);
or U850 (N_850,N_834,N_810);
or U851 (N_851,N_830,N_820);
or U852 (N_852,N_798,N_808);
nor U853 (N_853,N_793,N_809);
or U854 (N_854,N_782,N_780);
or U855 (N_855,N_783,N_828);
nor U856 (N_856,N_832,N_784);
nand U857 (N_857,N_800,N_816);
or U858 (N_858,N_812,N_803);
nand U859 (N_859,N_813,N_781);
nand U860 (N_860,N_831,N_790);
nor U861 (N_861,N_824,N_827);
nand U862 (N_862,N_839,N_796);
or U863 (N_863,N_837,N_815);
nor U864 (N_864,N_833,N_806);
or U865 (N_865,N_791,N_807);
or U866 (N_866,N_822,N_794);
and U867 (N_867,N_826,N_805);
and U868 (N_868,N_829,N_825);
nor U869 (N_869,N_795,N_788);
nor U870 (N_870,N_801,N_831);
nand U871 (N_871,N_824,N_787);
or U872 (N_872,N_838,N_814);
nand U873 (N_873,N_795,N_785);
nor U874 (N_874,N_814,N_832);
and U875 (N_875,N_821,N_791);
and U876 (N_876,N_832,N_798);
or U877 (N_877,N_787,N_786);
nand U878 (N_878,N_815,N_810);
xnor U879 (N_879,N_791,N_825);
or U880 (N_880,N_799,N_800);
or U881 (N_881,N_819,N_801);
nand U882 (N_882,N_827,N_816);
xnor U883 (N_883,N_802,N_820);
nor U884 (N_884,N_827,N_781);
and U885 (N_885,N_798,N_787);
nand U886 (N_886,N_822,N_802);
nor U887 (N_887,N_812,N_824);
or U888 (N_888,N_815,N_790);
or U889 (N_889,N_791,N_798);
and U890 (N_890,N_809,N_827);
xnor U891 (N_891,N_829,N_790);
or U892 (N_892,N_812,N_832);
xor U893 (N_893,N_808,N_829);
and U894 (N_894,N_781,N_828);
nand U895 (N_895,N_828,N_816);
or U896 (N_896,N_788,N_836);
nand U897 (N_897,N_838,N_831);
and U898 (N_898,N_789,N_795);
or U899 (N_899,N_785,N_807);
nand U900 (N_900,N_864,N_848);
or U901 (N_901,N_884,N_855);
nor U902 (N_902,N_897,N_887);
nor U903 (N_903,N_854,N_886);
nor U904 (N_904,N_892,N_893);
or U905 (N_905,N_858,N_845);
xnor U906 (N_906,N_889,N_894);
or U907 (N_907,N_861,N_878);
nand U908 (N_908,N_841,N_843);
and U909 (N_909,N_849,N_865);
and U910 (N_910,N_882,N_871);
and U911 (N_911,N_879,N_862);
nor U912 (N_912,N_860,N_857);
nand U913 (N_913,N_842,N_877);
and U914 (N_914,N_873,N_856);
nor U915 (N_915,N_863,N_880);
nand U916 (N_916,N_866,N_844);
or U917 (N_917,N_840,N_885);
nor U918 (N_918,N_898,N_874);
nor U919 (N_919,N_876,N_896);
and U920 (N_920,N_859,N_853);
xnor U921 (N_921,N_891,N_895);
or U922 (N_922,N_890,N_851);
nand U923 (N_923,N_869,N_870);
xor U924 (N_924,N_850,N_881);
or U925 (N_925,N_868,N_875);
nor U926 (N_926,N_867,N_888);
nand U927 (N_927,N_847,N_852);
and U928 (N_928,N_872,N_883);
or U929 (N_929,N_846,N_899);
nor U930 (N_930,N_878,N_867);
or U931 (N_931,N_862,N_881);
nor U932 (N_932,N_848,N_859);
xor U933 (N_933,N_887,N_851);
nand U934 (N_934,N_886,N_875);
or U935 (N_935,N_872,N_844);
and U936 (N_936,N_882,N_843);
xnor U937 (N_937,N_887,N_850);
or U938 (N_938,N_899,N_890);
or U939 (N_939,N_853,N_840);
and U940 (N_940,N_864,N_865);
xnor U941 (N_941,N_877,N_856);
or U942 (N_942,N_879,N_853);
or U943 (N_943,N_894,N_862);
xor U944 (N_944,N_841,N_863);
nor U945 (N_945,N_847,N_893);
and U946 (N_946,N_840,N_861);
and U947 (N_947,N_866,N_855);
and U948 (N_948,N_848,N_861);
and U949 (N_949,N_861,N_897);
and U950 (N_950,N_897,N_863);
nor U951 (N_951,N_881,N_897);
and U952 (N_952,N_870,N_848);
xor U953 (N_953,N_870,N_881);
nor U954 (N_954,N_875,N_851);
nor U955 (N_955,N_869,N_895);
and U956 (N_956,N_871,N_879);
and U957 (N_957,N_883,N_870);
xor U958 (N_958,N_873,N_878);
nand U959 (N_959,N_853,N_868);
nor U960 (N_960,N_950,N_926);
xor U961 (N_961,N_917,N_915);
xor U962 (N_962,N_906,N_958);
nand U963 (N_963,N_945,N_909);
nor U964 (N_964,N_923,N_913);
and U965 (N_965,N_907,N_928);
or U966 (N_966,N_959,N_904);
and U967 (N_967,N_927,N_911);
or U968 (N_968,N_949,N_908);
or U969 (N_969,N_952,N_942);
or U970 (N_970,N_914,N_916);
nand U971 (N_971,N_919,N_938);
and U972 (N_972,N_944,N_954);
nand U973 (N_973,N_936,N_924);
and U974 (N_974,N_937,N_943);
and U975 (N_975,N_930,N_929);
nor U976 (N_976,N_905,N_921);
xor U977 (N_977,N_939,N_903);
and U978 (N_978,N_918,N_940);
or U979 (N_979,N_941,N_902);
nand U980 (N_980,N_925,N_931);
or U981 (N_981,N_951,N_953);
nor U982 (N_982,N_912,N_955);
nand U983 (N_983,N_933,N_920);
and U984 (N_984,N_901,N_946);
nand U985 (N_985,N_957,N_900);
and U986 (N_986,N_910,N_934);
nor U987 (N_987,N_935,N_948);
xnor U988 (N_988,N_922,N_956);
and U989 (N_989,N_932,N_947);
nor U990 (N_990,N_907,N_906);
nor U991 (N_991,N_905,N_949);
or U992 (N_992,N_901,N_937);
or U993 (N_993,N_945,N_936);
or U994 (N_994,N_918,N_949);
xor U995 (N_995,N_917,N_946);
nor U996 (N_996,N_958,N_950);
or U997 (N_997,N_924,N_955);
nor U998 (N_998,N_937,N_916);
nor U999 (N_999,N_918,N_909);
nand U1000 (N_1000,N_916,N_909);
nor U1001 (N_1001,N_909,N_939);
and U1002 (N_1002,N_952,N_903);
nor U1003 (N_1003,N_945,N_924);
or U1004 (N_1004,N_915,N_923);
nor U1005 (N_1005,N_933,N_958);
or U1006 (N_1006,N_957,N_903);
or U1007 (N_1007,N_908,N_937);
nand U1008 (N_1008,N_921,N_919);
nor U1009 (N_1009,N_954,N_916);
nor U1010 (N_1010,N_918,N_929);
or U1011 (N_1011,N_901,N_924);
xnor U1012 (N_1012,N_932,N_909);
and U1013 (N_1013,N_954,N_918);
and U1014 (N_1014,N_905,N_926);
nand U1015 (N_1015,N_942,N_923);
or U1016 (N_1016,N_942,N_903);
or U1017 (N_1017,N_950,N_941);
and U1018 (N_1018,N_918,N_916);
nor U1019 (N_1019,N_929,N_941);
and U1020 (N_1020,N_975,N_999);
xor U1021 (N_1021,N_984,N_994);
or U1022 (N_1022,N_993,N_1012);
nor U1023 (N_1023,N_973,N_972);
nor U1024 (N_1024,N_1013,N_1019);
nor U1025 (N_1025,N_961,N_1006);
xnor U1026 (N_1026,N_997,N_967);
nor U1027 (N_1027,N_991,N_974);
nand U1028 (N_1028,N_1008,N_964);
nand U1029 (N_1029,N_1003,N_977);
xnor U1030 (N_1030,N_1015,N_996);
and U1031 (N_1031,N_1004,N_980);
or U1032 (N_1032,N_970,N_992);
or U1033 (N_1033,N_963,N_965);
nor U1034 (N_1034,N_990,N_969);
nor U1035 (N_1035,N_978,N_979);
or U1036 (N_1036,N_1005,N_986);
xnor U1037 (N_1037,N_966,N_982);
and U1038 (N_1038,N_987,N_985);
nand U1039 (N_1039,N_962,N_976);
or U1040 (N_1040,N_1017,N_971);
xor U1041 (N_1041,N_1002,N_960);
or U1042 (N_1042,N_968,N_1010);
nand U1043 (N_1043,N_998,N_1011);
nor U1044 (N_1044,N_983,N_1000);
xnor U1045 (N_1045,N_981,N_1007);
nor U1046 (N_1046,N_1014,N_1016);
and U1047 (N_1047,N_1018,N_1009);
nand U1048 (N_1048,N_1001,N_988);
nand U1049 (N_1049,N_989,N_995);
nor U1050 (N_1050,N_990,N_1019);
or U1051 (N_1051,N_991,N_969);
or U1052 (N_1052,N_1007,N_990);
nand U1053 (N_1053,N_974,N_993);
nand U1054 (N_1054,N_973,N_994);
xor U1055 (N_1055,N_1016,N_1005);
and U1056 (N_1056,N_963,N_980);
nor U1057 (N_1057,N_981,N_968);
nor U1058 (N_1058,N_963,N_970);
xor U1059 (N_1059,N_1003,N_1018);
nor U1060 (N_1060,N_1012,N_1018);
nor U1061 (N_1061,N_979,N_1014);
or U1062 (N_1062,N_1010,N_1000);
or U1063 (N_1063,N_966,N_989);
and U1064 (N_1064,N_992,N_1003);
and U1065 (N_1065,N_1016,N_995);
xor U1066 (N_1066,N_978,N_998);
xor U1067 (N_1067,N_975,N_1010);
and U1068 (N_1068,N_1002,N_970);
xnor U1069 (N_1069,N_995,N_1004);
and U1070 (N_1070,N_1007,N_1018);
and U1071 (N_1071,N_965,N_987);
and U1072 (N_1072,N_975,N_1004);
nor U1073 (N_1073,N_967,N_968);
nand U1074 (N_1074,N_996,N_989);
nor U1075 (N_1075,N_993,N_978);
nor U1076 (N_1076,N_1012,N_994);
nand U1077 (N_1077,N_990,N_1008);
and U1078 (N_1078,N_987,N_1000);
nor U1079 (N_1079,N_993,N_962);
nand U1080 (N_1080,N_1068,N_1042);
xnor U1081 (N_1081,N_1020,N_1054);
or U1082 (N_1082,N_1023,N_1067);
xor U1083 (N_1083,N_1027,N_1051);
xor U1084 (N_1084,N_1066,N_1064);
nand U1085 (N_1085,N_1029,N_1073);
nor U1086 (N_1086,N_1037,N_1022);
xnor U1087 (N_1087,N_1070,N_1078);
xor U1088 (N_1088,N_1039,N_1025);
and U1089 (N_1089,N_1062,N_1032);
or U1090 (N_1090,N_1069,N_1035);
nand U1091 (N_1091,N_1034,N_1050);
or U1092 (N_1092,N_1043,N_1033);
and U1093 (N_1093,N_1075,N_1060);
and U1094 (N_1094,N_1076,N_1058);
nor U1095 (N_1095,N_1044,N_1063);
xor U1096 (N_1096,N_1071,N_1057);
nand U1097 (N_1097,N_1055,N_1036);
xnor U1098 (N_1098,N_1074,N_1046);
nand U1099 (N_1099,N_1072,N_1048);
nand U1100 (N_1100,N_1065,N_1056);
nor U1101 (N_1101,N_1047,N_1059);
nor U1102 (N_1102,N_1038,N_1052);
or U1103 (N_1103,N_1040,N_1049);
nand U1104 (N_1104,N_1077,N_1021);
nand U1105 (N_1105,N_1053,N_1045);
nand U1106 (N_1106,N_1024,N_1061);
and U1107 (N_1107,N_1031,N_1041);
or U1108 (N_1108,N_1079,N_1026);
and U1109 (N_1109,N_1028,N_1030);
nor U1110 (N_1110,N_1020,N_1064);
and U1111 (N_1111,N_1023,N_1054);
and U1112 (N_1112,N_1054,N_1042);
and U1113 (N_1113,N_1070,N_1060);
nor U1114 (N_1114,N_1077,N_1034);
and U1115 (N_1115,N_1032,N_1070);
or U1116 (N_1116,N_1045,N_1041);
xnor U1117 (N_1117,N_1034,N_1065);
and U1118 (N_1118,N_1023,N_1038);
nor U1119 (N_1119,N_1030,N_1049);
nor U1120 (N_1120,N_1060,N_1024);
or U1121 (N_1121,N_1072,N_1045);
nand U1122 (N_1122,N_1040,N_1030);
nand U1123 (N_1123,N_1068,N_1051);
xor U1124 (N_1124,N_1042,N_1075);
nand U1125 (N_1125,N_1022,N_1069);
nand U1126 (N_1126,N_1026,N_1054);
nand U1127 (N_1127,N_1068,N_1030);
nor U1128 (N_1128,N_1050,N_1020);
and U1129 (N_1129,N_1060,N_1063);
nor U1130 (N_1130,N_1039,N_1035);
nand U1131 (N_1131,N_1028,N_1063);
and U1132 (N_1132,N_1069,N_1060);
xnor U1133 (N_1133,N_1028,N_1033);
xor U1134 (N_1134,N_1022,N_1060);
or U1135 (N_1135,N_1039,N_1050);
xor U1136 (N_1136,N_1046,N_1037);
and U1137 (N_1137,N_1066,N_1060);
nand U1138 (N_1138,N_1067,N_1056);
or U1139 (N_1139,N_1059,N_1030);
or U1140 (N_1140,N_1112,N_1088);
or U1141 (N_1141,N_1084,N_1138);
nand U1142 (N_1142,N_1101,N_1117);
and U1143 (N_1143,N_1116,N_1093);
nand U1144 (N_1144,N_1114,N_1111);
nor U1145 (N_1145,N_1085,N_1119);
nor U1146 (N_1146,N_1108,N_1098);
or U1147 (N_1147,N_1135,N_1125);
and U1148 (N_1148,N_1100,N_1124);
and U1149 (N_1149,N_1109,N_1090);
nor U1150 (N_1150,N_1106,N_1096);
or U1151 (N_1151,N_1115,N_1120);
and U1152 (N_1152,N_1105,N_1095);
nand U1153 (N_1153,N_1081,N_1134);
xor U1154 (N_1154,N_1122,N_1102);
and U1155 (N_1155,N_1082,N_1107);
nor U1156 (N_1156,N_1113,N_1097);
nor U1157 (N_1157,N_1139,N_1126);
and U1158 (N_1158,N_1123,N_1133);
nor U1159 (N_1159,N_1137,N_1110);
or U1160 (N_1160,N_1131,N_1092);
and U1161 (N_1161,N_1118,N_1087);
or U1162 (N_1162,N_1091,N_1080);
nand U1163 (N_1163,N_1103,N_1132);
or U1164 (N_1164,N_1121,N_1127);
nand U1165 (N_1165,N_1128,N_1130);
nand U1166 (N_1166,N_1136,N_1089);
or U1167 (N_1167,N_1086,N_1094);
or U1168 (N_1168,N_1083,N_1099);
nor U1169 (N_1169,N_1129,N_1104);
and U1170 (N_1170,N_1119,N_1082);
nor U1171 (N_1171,N_1096,N_1139);
and U1172 (N_1172,N_1125,N_1114);
nor U1173 (N_1173,N_1132,N_1133);
and U1174 (N_1174,N_1093,N_1089);
and U1175 (N_1175,N_1117,N_1136);
nand U1176 (N_1176,N_1096,N_1089);
or U1177 (N_1177,N_1109,N_1128);
and U1178 (N_1178,N_1132,N_1129);
or U1179 (N_1179,N_1107,N_1106);
nand U1180 (N_1180,N_1102,N_1112);
and U1181 (N_1181,N_1123,N_1114);
xnor U1182 (N_1182,N_1098,N_1123);
nand U1183 (N_1183,N_1135,N_1115);
nand U1184 (N_1184,N_1138,N_1083);
nor U1185 (N_1185,N_1093,N_1123);
nor U1186 (N_1186,N_1138,N_1130);
and U1187 (N_1187,N_1127,N_1081);
xnor U1188 (N_1188,N_1082,N_1130);
nor U1189 (N_1189,N_1132,N_1107);
and U1190 (N_1190,N_1090,N_1092);
or U1191 (N_1191,N_1116,N_1085);
or U1192 (N_1192,N_1118,N_1098);
or U1193 (N_1193,N_1131,N_1137);
xnor U1194 (N_1194,N_1101,N_1131);
nor U1195 (N_1195,N_1098,N_1135);
and U1196 (N_1196,N_1090,N_1096);
nand U1197 (N_1197,N_1086,N_1132);
nor U1198 (N_1198,N_1087,N_1081);
nand U1199 (N_1199,N_1094,N_1123);
and U1200 (N_1200,N_1159,N_1168);
nor U1201 (N_1201,N_1156,N_1157);
and U1202 (N_1202,N_1175,N_1153);
or U1203 (N_1203,N_1194,N_1191);
nor U1204 (N_1204,N_1185,N_1145);
or U1205 (N_1205,N_1141,N_1154);
and U1206 (N_1206,N_1161,N_1149);
nand U1207 (N_1207,N_1173,N_1140);
nand U1208 (N_1208,N_1162,N_1160);
and U1209 (N_1209,N_1192,N_1195);
nor U1210 (N_1210,N_1147,N_1158);
and U1211 (N_1211,N_1187,N_1193);
nand U1212 (N_1212,N_1178,N_1151);
xor U1213 (N_1213,N_1144,N_1184);
and U1214 (N_1214,N_1163,N_1146);
nand U1215 (N_1215,N_1186,N_1180);
or U1216 (N_1216,N_1189,N_1183);
and U1217 (N_1217,N_1167,N_1142);
xnor U1218 (N_1218,N_1155,N_1171);
nor U1219 (N_1219,N_1174,N_1152);
and U1220 (N_1220,N_1172,N_1164);
nand U1221 (N_1221,N_1199,N_1190);
or U1222 (N_1222,N_1179,N_1150);
and U1223 (N_1223,N_1166,N_1143);
or U1224 (N_1224,N_1198,N_1181);
nor U1225 (N_1225,N_1182,N_1169);
nor U1226 (N_1226,N_1188,N_1197);
nor U1227 (N_1227,N_1148,N_1165);
nor U1228 (N_1228,N_1176,N_1177);
and U1229 (N_1229,N_1170,N_1196);
nand U1230 (N_1230,N_1192,N_1159);
or U1231 (N_1231,N_1181,N_1169);
nor U1232 (N_1232,N_1155,N_1146);
xnor U1233 (N_1233,N_1158,N_1169);
and U1234 (N_1234,N_1154,N_1144);
and U1235 (N_1235,N_1198,N_1180);
nor U1236 (N_1236,N_1162,N_1153);
xnor U1237 (N_1237,N_1149,N_1188);
nor U1238 (N_1238,N_1164,N_1143);
and U1239 (N_1239,N_1146,N_1161);
nand U1240 (N_1240,N_1171,N_1166);
or U1241 (N_1241,N_1190,N_1178);
or U1242 (N_1242,N_1159,N_1189);
and U1243 (N_1243,N_1159,N_1140);
nor U1244 (N_1244,N_1194,N_1170);
and U1245 (N_1245,N_1161,N_1189);
nand U1246 (N_1246,N_1168,N_1183);
nand U1247 (N_1247,N_1175,N_1191);
xnor U1248 (N_1248,N_1193,N_1159);
and U1249 (N_1249,N_1161,N_1144);
nand U1250 (N_1250,N_1182,N_1175);
xnor U1251 (N_1251,N_1199,N_1143);
nor U1252 (N_1252,N_1191,N_1177);
nor U1253 (N_1253,N_1155,N_1163);
nor U1254 (N_1254,N_1153,N_1166);
or U1255 (N_1255,N_1166,N_1199);
nand U1256 (N_1256,N_1183,N_1145);
nand U1257 (N_1257,N_1153,N_1163);
nor U1258 (N_1258,N_1196,N_1181);
nor U1259 (N_1259,N_1180,N_1165);
or U1260 (N_1260,N_1230,N_1238);
and U1261 (N_1261,N_1211,N_1239);
and U1262 (N_1262,N_1233,N_1222);
nor U1263 (N_1263,N_1253,N_1236);
and U1264 (N_1264,N_1256,N_1200);
nand U1265 (N_1265,N_1213,N_1224);
or U1266 (N_1266,N_1225,N_1245);
nor U1267 (N_1267,N_1223,N_1206);
nor U1268 (N_1268,N_1210,N_1227);
nor U1269 (N_1269,N_1244,N_1207);
and U1270 (N_1270,N_1254,N_1234);
nor U1271 (N_1271,N_1220,N_1218);
nand U1272 (N_1272,N_1204,N_1242);
nor U1273 (N_1273,N_1209,N_1205);
nand U1274 (N_1274,N_1214,N_1250);
or U1275 (N_1275,N_1235,N_1246);
nor U1276 (N_1276,N_1240,N_1243);
nor U1277 (N_1277,N_1255,N_1221);
nor U1278 (N_1278,N_1217,N_1215);
or U1279 (N_1279,N_1249,N_1247);
nand U1280 (N_1280,N_1241,N_1231);
nand U1281 (N_1281,N_1203,N_1202);
nor U1282 (N_1282,N_1232,N_1228);
and U1283 (N_1283,N_1258,N_1257);
or U1284 (N_1284,N_1201,N_1226);
and U1285 (N_1285,N_1219,N_1252);
nor U1286 (N_1286,N_1212,N_1248);
xnor U1287 (N_1287,N_1259,N_1216);
or U1288 (N_1288,N_1208,N_1251);
nand U1289 (N_1289,N_1229,N_1237);
nor U1290 (N_1290,N_1202,N_1207);
and U1291 (N_1291,N_1206,N_1202);
or U1292 (N_1292,N_1220,N_1245);
nor U1293 (N_1293,N_1244,N_1252);
and U1294 (N_1294,N_1205,N_1211);
xnor U1295 (N_1295,N_1212,N_1231);
nand U1296 (N_1296,N_1246,N_1245);
or U1297 (N_1297,N_1237,N_1203);
and U1298 (N_1298,N_1256,N_1224);
and U1299 (N_1299,N_1247,N_1250);
and U1300 (N_1300,N_1230,N_1208);
nor U1301 (N_1301,N_1232,N_1204);
or U1302 (N_1302,N_1253,N_1213);
and U1303 (N_1303,N_1242,N_1201);
nand U1304 (N_1304,N_1235,N_1249);
and U1305 (N_1305,N_1255,N_1232);
or U1306 (N_1306,N_1228,N_1252);
nand U1307 (N_1307,N_1227,N_1250);
nand U1308 (N_1308,N_1214,N_1218);
xor U1309 (N_1309,N_1259,N_1219);
or U1310 (N_1310,N_1259,N_1257);
and U1311 (N_1311,N_1254,N_1207);
nand U1312 (N_1312,N_1238,N_1234);
nor U1313 (N_1313,N_1205,N_1223);
nor U1314 (N_1314,N_1236,N_1257);
nor U1315 (N_1315,N_1246,N_1226);
nand U1316 (N_1316,N_1243,N_1208);
nand U1317 (N_1317,N_1230,N_1234);
xor U1318 (N_1318,N_1241,N_1223);
nand U1319 (N_1319,N_1241,N_1253);
nor U1320 (N_1320,N_1271,N_1301);
nand U1321 (N_1321,N_1309,N_1317);
nand U1322 (N_1322,N_1273,N_1267);
nand U1323 (N_1323,N_1296,N_1279);
and U1324 (N_1324,N_1307,N_1261);
nor U1325 (N_1325,N_1306,N_1300);
nand U1326 (N_1326,N_1290,N_1272);
or U1327 (N_1327,N_1313,N_1284);
nand U1328 (N_1328,N_1278,N_1292);
nand U1329 (N_1329,N_1310,N_1285);
nand U1330 (N_1330,N_1299,N_1268);
and U1331 (N_1331,N_1281,N_1270);
nor U1332 (N_1332,N_1303,N_1280);
or U1333 (N_1333,N_1260,N_1276);
or U1334 (N_1334,N_1269,N_1294);
nand U1335 (N_1335,N_1287,N_1293);
nor U1336 (N_1336,N_1263,N_1291);
nor U1337 (N_1337,N_1266,N_1264);
or U1338 (N_1338,N_1286,N_1289);
and U1339 (N_1339,N_1295,N_1298);
nand U1340 (N_1340,N_1283,N_1315);
nor U1341 (N_1341,N_1277,N_1311);
nand U1342 (N_1342,N_1265,N_1304);
nand U1343 (N_1343,N_1282,N_1318);
nor U1344 (N_1344,N_1319,N_1297);
nor U1345 (N_1345,N_1308,N_1262);
and U1346 (N_1346,N_1275,N_1314);
nand U1347 (N_1347,N_1305,N_1288);
nor U1348 (N_1348,N_1274,N_1312);
nand U1349 (N_1349,N_1302,N_1316);
or U1350 (N_1350,N_1311,N_1304);
xor U1351 (N_1351,N_1271,N_1266);
xnor U1352 (N_1352,N_1287,N_1277);
xnor U1353 (N_1353,N_1319,N_1296);
nand U1354 (N_1354,N_1276,N_1297);
nor U1355 (N_1355,N_1312,N_1305);
nand U1356 (N_1356,N_1264,N_1314);
or U1357 (N_1357,N_1260,N_1308);
and U1358 (N_1358,N_1267,N_1263);
nand U1359 (N_1359,N_1287,N_1301);
or U1360 (N_1360,N_1283,N_1308);
nor U1361 (N_1361,N_1271,N_1273);
and U1362 (N_1362,N_1290,N_1285);
and U1363 (N_1363,N_1272,N_1306);
and U1364 (N_1364,N_1302,N_1315);
nand U1365 (N_1365,N_1302,N_1291);
nor U1366 (N_1366,N_1303,N_1284);
nor U1367 (N_1367,N_1311,N_1297);
nor U1368 (N_1368,N_1305,N_1276);
or U1369 (N_1369,N_1315,N_1310);
nor U1370 (N_1370,N_1269,N_1290);
xor U1371 (N_1371,N_1304,N_1294);
nor U1372 (N_1372,N_1275,N_1277);
xnor U1373 (N_1373,N_1285,N_1303);
xor U1374 (N_1374,N_1291,N_1303);
or U1375 (N_1375,N_1274,N_1299);
or U1376 (N_1376,N_1282,N_1280);
nand U1377 (N_1377,N_1289,N_1283);
nand U1378 (N_1378,N_1307,N_1318);
or U1379 (N_1379,N_1283,N_1318);
and U1380 (N_1380,N_1330,N_1361);
xnor U1381 (N_1381,N_1321,N_1365);
xnor U1382 (N_1382,N_1338,N_1335);
nor U1383 (N_1383,N_1372,N_1367);
nor U1384 (N_1384,N_1340,N_1376);
nor U1385 (N_1385,N_1323,N_1355);
nor U1386 (N_1386,N_1337,N_1368);
nand U1387 (N_1387,N_1329,N_1360);
nand U1388 (N_1388,N_1349,N_1356);
nor U1389 (N_1389,N_1366,N_1322);
or U1390 (N_1390,N_1331,N_1357);
or U1391 (N_1391,N_1332,N_1320);
nand U1392 (N_1392,N_1358,N_1325);
nor U1393 (N_1393,N_1344,N_1354);
nand U1394 (N_1394,N_1347,N_1379);
nand U1395 (N_1395,N_1346,N_1375);
and U1396 (N_1396,N_1333,N_1342);
nand U1397 (N_1397,N_1364,N_1377);
nand U1398 (N_1398,N_1369,N_1350);
or U1399 (N_1399,N_1327,N_1378);
nand U1400 (N_1400,N_1341,N_1359);
nand U1401 (N_1401,N_1363,N_1324);
or U1402 (N_1402,N_1370,N_1328);
or U1403 (N_1403,N_1348,N_1362);
or U1404 (N_1404,N_1326,N_1352);
nand U1405 (N_1405,N_1345,N_1339);
or U1406 (N_1406,N_1374,N_1373);
nand U1407 (N_1407,N_1334,N_1343);
nand U1408 (N_1408,N_1336,N_1351);
xnor U1409 (N_1409,N_1371,N_1353);
and U1410 (N_1410,N_1345,N_1321);
and U1411 (N_1411,N_1351,N_1323);
nor U1412 (N_1412,N_1344,N_1338);
or U1413 (N_1413,N_1327,N_1357);
and U1414 (N_1414,N_1360,N_1323);
nand U1415 (N_1415,N_1378,N_1367);
or U1416 (N_1416,N_1373,N_1349);
and U1417 (N_1417,N_1354,N_1322);
xor U1418 (N_1418,N_1327,N_1359);
nand U1419 (N_1419,N_1359,N_1340);
nand U1420 (N_1420,N_1370,N_1335);
and U1421 (N_1421,N_1348,N_1372);
nor U1422 (N_1422,N_1378,N_1329);
nor U1423 (N_1423,N_1321,N_1331);
nand U1424 (N_1424,N_1364,N_1349);
and U1425 (N_1425,N_1332,N_1373);
or U1426 (N_1426,N_1359,N_1371);
and U1427 (N_1427,N_1347,N_1374);
nor U1428 (N_1428,N_1323,N_1370);
and U1429 (N_1429,N_1327,N_1351);
nand U1430 (N_1430,N_1356,N_1370);
nand U1431 (N_1431,N_1333,N_1369);
nand U1432 (N_1432,N_1355,N_1371);
or U1433 (N_1433,N_1329,N_1375);
nor U1434 (N_1434,N_1333,N_1353);
and U1435 (N_1435,N_1342,N_1335);
xnor U1436 (N_1436,N_1349,N_1365);
nor U1437 (N_1437,N_1355,N_1349);
or U1438 (N_1438,N_1364,N_1334);
or U1439 (N_1439,N_1361,N_1377);
or U1440 (N_1440,N_1426,N_1424);
and U1441 (N_1441,N_1417,N_1404);
or U1442 (N_1442,N_1386,N_1427);
nand U1443 (N_1443,N_1414,N_1433);
nand U1444 (N_1444,N_1425,N_1429);
nor U1445 (N_1445,N_1401,N_1393);
nor U1446 (N_1446,N_1435,N_1418);
or U1447 (N_1447,N_1405,N_1389);
nand U1448 (N_1448,N_1410,N_1413);
and U1449 (N_1449,N_1407,N_1394);
nor U1450 (N_1450,N_1387,N_1390);
or U1451 (N_1451,N_1411,N_1391);
xnor U1452 (N_1452,N_1396,N_1419);
nand U1453 (N_1453,N_1412,N_1382);
and U1454 (N_1454,N_1431,N_1439);
nand U1455 (N_1455,N_1432,N_1416);
nand U1456 (N_1456,N_1399,N_1406);
nand U1457 (N_1457,N_1392,N_1388);
nor U1458 (N_1458,N_1408,N_1420);
and U1459 (N_1459,N_1421,N_1436);
or U1460 (N_1460,N_1402,N_1430);
and U1461 (N_1461,N_1415,N_1400);
xnor U1462 (N_1462,N_1380,N_1385);
nand U1463 (N_1463,N_1383,N_1422);
nor U1464 (N_1464,N_1423,N_1438);
or U1465 (N_1465,N_1437,N_1403);
nor U1466 (N_1466,N_1428,N_1409);
nand U1467 (N_1467,N_1395,N_1398);
or U1468 (N_1468,N_1384,N_1381);
nand U1469 (N_1469,N_1434,N_1397);
or U1470 (N_1470,N_1388,N_1391);
nor U1471 (N_1471,N_1390,N_1409);
nor U1472 (N_1472,N_1410,N_1419);
nand U1473 (N_1473,N_1407,N_1416);
nor U1474 (N_1474,N_1439,N_1384);
xor U1475 (N_1475,N_1401,N_1416);
nor U1476 (N_1476,N_1401,N_1387);
and U1477 (N_1477,N_1401,N_1382);
nand U1478 (N_1478,N_1404,N_1409);
and U1479 (N_1479,N_1407,N_1432);
and U1480 (N_1480,N_1408,N_1401);
or U1481 (N_1481,N_1437,N_1430);
nor U1482 (N_1482,N_1387,N_1399);
or U1483 (N_1483,N_1420,N_1399);
and U1484 (N_1484,N_1409,N_1435);
nand U1485 (N_1485,N_1428,N_1386);
nand U1486 (N_1486,N_1436,N_1403);
nand U1487 (N_1487,N_1419,N_1435);
or U1488 (N_1488,N_1403,N_1395);
nand U1489 (N_1489,N_1389,N_1408);
nor U1490 (N_1490,N_1395,N_1419);
nor U1491 (N_1491,N_1431,N_1403);
nand U1492 (N_1492,N_1421,N_1406);
xnor U1493 (N_1493,N_1387,N_1404);
nor U1494 (N_1494,N_1412,N_1391);
or U1495 (N_1495,N_1394,N_1403);
nand U1496 (N_1496,N_1420,N_1391);
or U1497 (N_1497,N_1418,N_1421);
xnor U1498 (N_1498,N_1380,N_1406);
nor U1499 (N_1499,N_1394,N_1439);
or U1500 (N_1500,N_1467,N_1441);
nor U1501 (N_1501,N_1442,N_1443);
nand U1502 (N_1502,N_1478,N_1491);
nand U1503 (N_1503,N_1471,N_1474);
nand U1504 (N_1504,N_1489,N_1454);
or U1505 (N_1505,N_1469,N_1494);
nor U1506 (N_1506,N_1447,N_1496);
or U1507 (N_1507,N_1452,N_1470);
nand U1508 (N_1508,N_1458,N_1464);
and U1509 (N_1509,N_1460,N_1487);
nor U1510 (N_1510,N_1497,N_1493);
nand U1511 (N_1511,N_1492,N_1490);
or U1512 (N_1512,N_1463,N_1477);
nand U1513 (N_1513,N_1480,N_1472);
nor U1514 (N_1514,N_1450,N_1482);
and U1515 (N_1515,N_1453,N_1473);
xor U1516 (N_1516,N_1483,N_1481);
nand U1517 (N_1517,N_1455,N_1461);
and U1518 (N_1518,N_1444,N_1475);
and U1519 (N_1519,N_1465,N_1486);
nor U1520 (N_1520,N_1445,N_1499);
xnor U1521 (N_1521,N_1459,N_1488);
or U1522 (N_1522,N_1468,N_1484);
and U1523 (N_1523,N_1448,N_1457);
and U1524 (N_1524,N_1456,N_1466);
and U1525 (N_1525,N_1485,N_1451);
nand U1526 (N_1526,N_1479,N_1462);
nand U1527 (N_1527,N_1449,N_1440);
nand U1528 (N_1528,N_1476,N_1498);
or U1529 (N_1529,N_1495,N_1446);
nor U1530 (N_1530,N_1476,N_1447);
nor U1531 (N_1531,N_1467,N_1488);
nor U1532 (N_1532,N_1455,N_1489);
and U1533 (N_1533,N_1449,N_1494);
and U1534 (N_1534,N_1479,N_1475);
xor U1535 (N_1535,N_1449,N_1450);
nor U1536 (N_1536,N_1483,N_1479);
or U1537 (N_1537,N_1482,N_1478);
nor U1538 (N_1538,N_1465,N_1455);
nor U1539 (N_1539,N_1447,N_1465);
or U1540 (N_1540,N_1483,N_1444);
and U1541 (N_1541,N_1463,N_1449);
and U1542 (N_1542,N_1468,N_1450);
nor U1543 (N_1543,N_1450,N_1469);
nand U1544 (N_1544,N_1495,N_1499);
or U1545 (N_1545,N_1452,N_1453);
xor U1546 (N_1546,N_1462,N_1449);
or U1547 (N_1547,N_1497,N_1457);
nand U1548 (N_1548,N_1483,N_1461);
and U1549 (N_1549,N_1449,N_1486);
nor U1550 (N_1550,N_1465,N_1484);
or U1551 (N_1551,N_1489,N_1457);
or U1552 (N_1552,N_1486,N_1447);
nor U1553 (N_1553,N_1448,N_1459);
or U1554 (N_1554,N_1444,N_1449);
nor U1555 (N_1555,N_1444,N_1442);
or U1556 (N_1556,N_1456,N_1473);
nor U1557 (N_1557,N_1468,N_1441);
and U1558 (N_1558,N_1480,N_1491);
and U1559 (N_1559,N_1465,N_1473);
nor U1560 (N_1560,N_1504,N_1529);
or U1561 (N_1561,N_1524,N_1517);
and U1562 (N_1562,N_1537,N_1536);
or U1563 (N_1563,N_1515,N_1533);
or U1564 (N_1564,N_1539,N_1527);
nand U1565 (N_1565,N_1505,N_1510);
nand U1566 (N_1566,N_1541,N_1509);
or U1567 (N_1567,N_1500,N_1531);
and U1568 (N_1568,N_1501,N_1556);
and U1569 (N_1569,N_1542,N_1552);
and U1570 (N_1570,N_1518,N_1535);
nand U1571 (N_1571,N_1557,N_1526);
or U1572 (N_1572,N_1547,N_1516);
nor U1573 (N_1573,N_1528,N_1558);
nand U1574 (N_1574,N_1538,N_1503);
nand U1575 (N_1575,N_1508,N_1532);
and U1576 (N_1576,N_1523,N_1512);
nand U1577 (N_1577,N_1520,N_1507);
or U1578 (N_1578,N_1519,N_1530);
and U1579 (N_1579,N_1553,N_1551);
nor U1580 (N_1580,N_1546,N_1549);
or U1581 (N_1581,N_1521,N_1514);
xnor U1582 (N_1582,N_1534,N_1545);
nor U1583 (N_1583,N_1554,N_1559);
or U1584 (N_1584,N_1550,N_1513);
nand U1585 (N_1585,N_1522,N_1506);
or U1586 (N_1586,N_1555,N_1543);
xor U1587 (N_1587,N_1511,N_1502);
nor U1588 (N_1588,N_1548,N_1544);
or U1589 (N_1589,N_1540,N_1525);
nor U1590 (N_1590,N_1522,N_1543);
nor U1591 (N_1591,N_1501,N_1537);
and U1592 (N_1592,N_1502,N_1542);
nor U1593 (N_1593,N_1505,N_1547);
and U1594 (N_1594,N_1558,N_1548);
or U1595 (N_1595,N_1549,N_1502);
or U1596 (N_1596,N_1503,N_1555);
and U1597 (N_1597,N_1535,N_1515);
nand U1598 (N_1598,N_1502,N_1524);
or U1599 (N_1599,N_1516,N_1557);
nand U1600 (N_1600,N_1512,N_1535);
nor U1601 (N_1601,N_1534,N_1520);
nand U1602 (N_1602,N_1504,N_1539);
nor U1603 (N_1603,N_1542,N_1516);
and U1604 (N_1604,N_1500,N_1551);
nand U1605 (N_1605,N_1530,N_1514);
xnor U1606 (N_1606,N_1548,N_1503);
or U1607 (N_1607,N_1517,N_1516);
and U1608 (N_1608,N_1535,N_1505);
and U1609 (N_1609,N_1514,N_1529);
or U1610 (N_1610,N_1528,N_1520);
and U1611 (N_1611,N_1511,N_1544);
and U1612 (N_1612,N_1527,N_1531);
or U1613 (N_1613,N_1518,N_1520);
or U1614 (N_1614,N_1521,N_1552);
or U1615 (N_1615,N_1520,N_1505);
or U1616 (N_1616,N_1525,N_1528);
or U1617 (N_1617,N_1533,N_1500);
xor U1618 (N_1618,N_1551,N_1515);
nand U1619 (N_1619,N_1506,N_1502);
nor U1620 (N_1620,N_1565,N_1613);
or U1621 (N_1621,N_1571,N_1570);
nand U1622 (N_1622,N_1592,N_1583);
and U1623 (N_1623,N_1563,N_1609);
nand U1624 (N_1624,N_1618,N_1579);
nand U1625 (N_1625,N_1597,N_1615);
nand U1626 (N_1626,N_1611,N_1566);
nand U1627 (N_1627,N_1585,N_1578);
nand U1628 (N_1628,N_1586,N_1608);
and U1629 (N_1629,N_1607,N_1590);
nor U1630 (N_1630,N_1605,N_1601);
and U1631 (N_1631,N_1614,N_1617);
nor U1632 (N_1632,N_1577,N_1588);
nand U1633 (N_1633,N_1568,N_1569);
or U1634 (N_1634,N_1561,N_1574);
nor U1635 (N_1635,N_1596,N_1595);
nand U1636 (N_1636,N_1616,N_1593);
nor U1637 (N_1637,N_1564,N_1619);
or U1638 (N_1638,N_1560,N_1589);
and U1639 (N_1639,N_1573,N_1581);
nand U1640 (N_1640,N_1584,N_1587);
nand U1641 (N_1641,N_1599,N_1572);
nor U1642 (N_1642,N_1562,N_1567);
nand U1643 (N_1643,N_1582,N_1576);
nand U1644 (N_1644,N_1600,N_1598);
and U1645 (N_1645,N_1602,N_1606);
and U1646 (N_1646,N_1610,N_1612);
or U1647 (N_1647,N_1580,N_1604);
nor U1648 (N_1648,N_1594,N_1591);
nor U1649 (N_1649,N_1575,N_1603);
and U1650 (N_1650,N_1579,N_1597);
and U1651 (N_1651,N_1600,N_1584);
and U1652 (N_1652,N_1600,N_1610);
nor U1653 (N_1653,N_1569,N_1563);
nor U1654 (N_1654,N_1576,N_1610);
xor U1655 (N_1655,N_1601,N_1572);
or U1656 (N_1656,N_1607,N_1598);
nor U1657 (N_1657,N_1592,N_1571);
and U1658 (N_1658,N_1615,N_1564);
or U1659 (N_1659,N_1591,N_1589);
nand U1660 (N_1660,N_1593,N_1594);
nor U1661 (N_1661,N_1567,N_1596);
nor U1662 (N_1662,N_1581,N_1595);
and U1663 (N_1663,N_1614,N_1565);
nand U1664 (N_1664,N_1619,N_1574);
nand U1665 (N_1665,N_1603,N_1589);
nor U1666 (N_1666,N_1616,N_1586);
or U1667 (N_1667,N_1579,N_1612);
or U1668 (N_1668,N_1610,N_1598);
and U1669 (N_1669,N_1575,N_1617);
nor U1670 (N_1670,N_1578,N_1570);
nor U1671 (N_1671,N_1574,N_1562);
or U1672 (N_1672,N_1599,N_1576);
nor U1673 (N_1673,N_1591,N_1612);
or U1674 (N_1674,N_1602,N_1585);
nor U1675 (N_1675,N_1607,N_1585);
and U1676 (N_1676,N_1613,N_1606);
and U1677 (N_1677,N_1598,N_1585);
nand U1678 (N_1678,N_1572,N_1588);
xnor U1679 (N_1679,N_1607,N_1580);
and U1680 (N_1680,N_1635,N_1675);
or U1681 (N_1681,N_1661,N_1655);
and U1682 (N_1682,N_1644,N_1673);
xor U1683 (N_1683,N_1621,N_1658);
nand U1684 (N_1684,N_1665,N_1632);
xor U1685 (N_1685,N_1654,N_1664);
and U1686 (N_1686,N_1656,N_1666);
or U1687 (N_1687,N_1657,N_1631);
nand U1688 (N_1688,N_1668,N_1650);
or U1689 (N_1689,N_1652,N_1622);
nand U1690 (N_1690,N_1653,N_1660);
nor U1691 (N_1691,N_1674,N_1641);
nor U1692 (N_1692,N_1642,N_1651);
and U1693 (N_1693,N_1676,N_1679);
nor U1694 (N_1694,N_1630,N_1627);
xor U1695 (N_1695,N_1620,N_1649);
or U1696 (N_1696,N_1626,N_1628);
nor U1697 (N_1697,N_1677,N_1634);
nor U1698 (N_1698,N_1643,N_1623);
and U1699 (N_1699,N_1647,N_1637);
nor U1700 (N_1700,N_1645,N_1670);
and U1701 (N_1701,N_1633,N_1671);
and U1702 (N_1702,N_1638,N_1629);
xnor U1703 (N_1703,N_1624,N_1663);
nand U1704 (N_1704,N_1636,N_1639);
or U1705 (N_1705,N_1669,N_1672);
nor U1706 (N_1706,N_1648,N_1640);
xnor U1707 (N_1707,N_1625,N_1646);
nand U1708 (N_1708,N_1678,N_1662);
or U1709 (N_1709,N_1667,N_1659);
and U1710 (N_1710,N_1640,N_1627);
nand U1711 (N_1711,N_1635,N_1652);
xor U1712 (N_1712,N_1666,N_1661);
nand U1713 (N_1713,N_1636,N_1673);
nand U1714 (N_1714,N_1633,N_1665);
nand U1715 (N_1715,N_1650,N_1626);
nand U1716 (N_1716,N_1639,N_1653);
nor U1717 (N_1717,N_1638,N_1663);
and U1718 (N_1718,N_1647,N_1662);
and U1719 (N_1719,N_1645,N_1676);
or U1720 (N_1720,N_1635,N_1668);
and U1721 (N_1721,N_1643,N_1655);
nor U1722 (N_1722,N_1632,N_1639);
nor U1723 (N_1723,N_1663,N_1636);
and U1724 (N_1724,N_1655,N_1640);
and U1725 (N_1725,N_1671,N_1645);
or U1726 (N_1726,N_1676,N_1643);
nand U1727 (N_1727,N_1679,N_1657);
nor U1728 (N_1728,N_1640,N_1674);
nor U1729 (N_1729,N_1667,N_1671);
nand U1730 (N_1730,N_1631,N_1668);
and U1731 (N_1731,N_1654,N_1675);
and U1732 (N_1732,N_1636,N_1620);
or U1733 (N_1733,N_1634,N_1651);
and U1734 (N_1734,N_1667,N_1648);
xnor U1735 (N_1735,N_1669,N_1656);
nand U1736 (N_1736,N_1677,N_1624);
nand U1737 (N_1737,N_1676,N_1652);
nor U1738 (N_1738,N_1631,N_1646);
or U1739 (N_1739,N_1656,N_1675);
nand U1740 (N_1740,N_1699,N_1726);
or U1741 (N_1741,N_1681,N_1711);
or U1742 (N_1742,N_1715,N_1737);
or U1743 (N_1743,N_1694,N_1698);
and U1744 (N_1744,N_1704,N_1707);
or U1745 (N_1745,N_1738,N_1700);
or U1746 (N_1746,N_1733,N_1724);
nor U1747 (N_1747,N_1705,N_1706);
nand U1748 (N_1748,N_1691,N_1683);
or U1749 (N_1749,N_1712,N_1688);
or U1750 (N_1750,N_1696,N_1731);
nor U1751 (N_1751,N_1736,N_1729);
nand U1752 (N_1752,N_1684,N_1739);
nor U1753 (N_1753,N_1695,N_1730);
nand U1754 (N_1754,N_1686,N_1693);
or U1755 (N_1755,N_1735,N_1732);
and U1756 (N_1756,N_1708,N_1719);
and U1757 (N_1757,N_1720,N_1714);
nand U1758 (N_1758,N_1716,N_1723);
nand U1759 (N_1759,N_1727,N_1702);
or U1760 (N_1760,N_1718,N_1721);
nand U1761 (N_1761,N_1703,N_1692);
and U1762 (N_1762,N_1728,N_1689);
and U1763 (N_1763,N_1710,N_1685);
nor U1764 (N_1764,N_1701,N_1690);
nand U1765 (N_1765,N_1722,N_1682);
or U1766 (N_1766,N_1687,N_1709);
nor U1767 (N_1767,N_1713,N_1680);
and U1768 (N_1768,N_1697,N_1725);
and U1769 (N_1769,N_1717,N_1734);
nand U1770 (N_1770,N_1733,N_1721);
and U1771 (N_1771,N_1686,N_1728);
xnor U1772 (N_1772,N_1690,N_1717);
or U1773 (N_1773,N_1687,N_1730);
nor U1774 (N_1774,N_1719,N_1694);
or U1775 (N_1775,N_1700,N_1718);
nor U1776 (N_1776,N_1688,N_1693);
or U1777 (N_1777,N_1707,N_1711);
nor U1778 (N_1778,N_1699,N_1688);
nor U1779 (N_1779,N_1680,N_1718);
and U1780 (N_1780,N_1728,N_1718);
or U1781 (N_1781,N_1727,N_1700);
xor U1782 (N_1782,N_1718,N_1688);
nor U1783 (N_1783,N_1731,N_1738);
or U1784 (N_1784,N_1699,N_1720);
nor U1785 (N_1785,N_1696,N_1727);
nand U1786 (N_1786,N_1724,N_1725);
and U1787 (N_1787,N_1721,N_1722);
nand U1788 (N_1788,N_1682,N_1699);
and U1789 (N_1789,N_1723,N_1703);
nand U1790 (N_1790,N_1701,N_1737);
nor U1791 (N_1791,N_1716,N_1733);
and U1792 (N_1792,N_1688,N_1719);
and U1793 (N_1793,N_1680,N_1720);
and U1794 (N_1794,N_1707,N_1698);
xor U1795 (N_1795,N_1721,N_1734);
nand U1796 (N_1796,N_1710,N_1702);
nor U1797 (N_1797,N_1719,N_1682);
nand U1798 (N_1798,N_1701,N_1708);
and U1799 (N_1799,N_1702,N_1700);
and U1800 (N_1800,N_1797,N_1788);
and U1801 (N_1801,N_1785,N_1778);
and U1802 (N_1802,N_1774,N_1779);
nand U1803 (N_1803,N_1742,N_1762);
xnor U1804 (N_1804,N_1784,N_1782);
nor U1805 (N_1805,N_1771,N_1745);
and U1806 (N_1806,N_1773,N_1768);
nor U1807 (N_1807,N_1765,N_1786);
nand U1808 (N_1808,N_1760,N_1789);
nor U1809 (N_1809,N_1777,N_1767);
nor U1810 (N_1810,N_1770,N_1776);
nor U1811 (N_1811,N_1756,N_1751);
or U1812 (N_1812,N_1755,N_1754);
nand U1813 (N_1813,N_1750,N_1787);
or U1814 (N_1814,N_1758,N_1792);
xor U1815 (N_1815,N_1766,N_1761);
and U1816 (N_1816,N_1799,N_1746);
xor U1817 (N_1817,N_1741,N_1744);
or U1818 (N_1818,N_1763,N_1795);
xnor U1819 (N_1819,N_1794,N_1783);
nor U1820 (N_1820,N_1781,N_1780);
xnor U1821 (N_1821,N_1790,N_1793);
nor U1822 (N_1822,N_1740,N_1769);
or U1823 (N_1823,N_1757,N_1747);
or U1824 (N_1824,N_1796,N_1749);
or U1825 (N_1825,N_1764,N_1791);
nand U1826 (N_1826,N_1743,N_1752);
nand U1827 (N_1827,N_1772,N_1759);
nor U1828 (N_1828,N_1798,N_1753);
xor U1829 (N_1829,N_1748,N_1775);
and U1830 (N_1830,N_1745,N_1746);
or U1831 (N_1831,N_1766,N_1777);
and U1832 (N_1832,N_1754,N_1758);
or U1833 (N_1833,N_1791,N_1774);
or U1834 (N_1834,N_1777,N_1781);
nor U1835 (N_1835,N_1760,N_1763);
nor U1836 (N_1836,N_1794,N_1756);
and U1837 (N_1837,N_1762,N_1758);
and U1838 (N_1838,N_1755,N_1764);
or U1839 (N_1839,N_1780,N_1750);
nor U1840 (N_1840,N_1762,N_1753);
or U1841 (N_1841,N_1793,N_1774);
nor U1842 (N_1842,N_1754,N_1744);
and U1843 (N_1843,N_1750,N_1748);
nand U1844 (N_1844,N_1748,N_1790);
and U1845 (N_1845,N_1771,N_1758);
nand U1846 (N_1846,N_1741,N_1799);
nor U1847 (N_1847,N_1764,N_1769);
and U1848 (N_1848,N_1780,N_1769);
nand U1849 (N_1849,N_1776,N_1788);
and U1850 (N_1850,N_1760,N_1774);
or U1851 (N_1851,N_1747,N_1794);
xnor U1852 (N_1852,N_1780,N_1784);
and U1853 (N_1853,N_1789,N_1748);
nor U1854 (N_1854,N_1765,N_1764);
nor U1855 (N_1855,N_1777,N_1760);
xor U1856 (N_1856,N_1758,N_1782);
nor U1857 (N_1857,N_1783,N_1742);
xor U1858 (N_1858,N_1785,N_1765);
or U1859 (N_1859,N_1766,N_1753);
xnor U1860 (N_1860,N_1841,N_1851);
xnor U1861 (N_1861,N_1859,N_1849);
and U1862 (N_1862,N_1850,N_1819);
and U1863 (N_1863,N_1832,N_1822);
and U1864 (N_1864,N_1844,N_1837);
or U1865 (N_1865,N_1829,N_1840);
or U1866 (N_1866,N_1853,N_1815);
xor U1867 (N_1867,N_1802,N_1813);
nand U1868 (N_1868,N_1812,N_1821);
nor U1869 (N_1869,N_1828,N_1843);
nand U1870 (N_1870,N_1852,N_1854);
nor U1871 (N_1871,N_1816,N_1858);
and U1872 (N_1872,N_1817,N_1823);
nor U1873 (N_1873,N_1801,N_1818);
nor U1874 (N_1874,N_1838,N_1836);
or U1875 (N_1875,N_1811,N_1848);
or U1876 (N_1876,N_1809,N_1835);
nor U1877 (N_1877,N_1806,N_1804);
and U1878 (N_1878,N_1824,N_1810);
nor U1879 (N_1879,N_1825,N_1820);
xnor U1880 (N_1880,N_1833,N_1827);
nand U1881 (N_1881,N_1846,N_1855);
or U1882 (N_1882,N_1805,N_1807);
and U1883 (N_1883,N_1834,N_1831);
and U1884 (N_1884,N_1803,N_1830);
nor U1885 (N_1885,N_1847,N_1839);
or U1886 (N_1886,N_1856,N_1842);
nand U1887 (N_1887,N_1814,N_1826);
and U1888 (N_1888,N_1845,N_1857);
or U1889 (N_1889,N_1808,N_1800);
nand U1890 (N_1890,N_1840,N_1847);
nand U1891 (N_1891,N_1859,N_1819);
nor U1892 (N_1892,N_1836,N_1849);
xnor U1893 (N_1893,N_1838,N_1855);
nor U1894 (N_1894,N_1845,N_1834);
nand U1895 (N_1895,N_1821,N_1838);
and U1896 (N_1896,N_1829,N_1808);
or U1897 (N_1897,N_1844,N_1855);
nand U1898 (N_1898,N_1845,N_1821);
nand U1899 (N_1899,N_1856,N_1834);
nand U1900 (N_1900,N_1813,N_1808);
nand U1901 (N_1901,N_1849,N_1817);
or U1902 (N_1902,N_1805,N_1834);
nor U1903 (N_1903,N_1812,N_1835);
nand U1904 (N_1904,N_1828,N_1839);
and U1905 (N_1905,N_1818,N_1803);
and U1906 (N_1906,N_1845,N_1855);
nand U1907 (N_1907,N_1823,N_1808);
or U1908 (N_1908,N_1838,N_1818);
and U1909 (N_1909,N_1855,N_1824);
nor U1910 (N_1910,N_1814,N_1831);
and U1911 (N_1911,N_1838,N_1816);
nand U1912 (N_1912,N_1831,N_1838);
nor U1913 (N_1913,N_1804,N_1811);
nor U1914 (N_1914,N_1833,N_1854);
nand U1915 (N_1915,N_1823,N_1838);
xnor U1916 (N_1916,N_1805,N_1818);
or U1917 (N_1917,N_1855,N_1809);
nor U1918 (N_1918,N_1800,N_1820);
nand U1919 (N_1919,N_1809,N_1814);
nand U1920 (N_1920,N_1914,N_1903);
nor U1921 (N_1921,N_1872,N_1884);
and U1922 (N_1922,N_1889,N_1880);
and U1923 (N_1923,N_1918,N_1892);
and U1924 (N_1924,N_1906,N_1897);
or U1925 (N_1925,N_1912,N_1900);
xor U1926 (N_1926,N_1870,N_1877);
nor U1927 (N_1927,N_1898,N_1891);
nand U1928 (N_1928,N_1890,N_1863);
or U1929 (N_1929,N_1917,N_1869);
xor U1930 (N_1930,N_1881,N_1916);
nor U1931 (N_1931,N_1861,N_1910);
nand U1932 (N_1932,N_1911,N_1878);
and U1933 (N_1933,N_1876,N_1907);
nand U1934 (N_1934,N_1864,N_1886);
xnor U1935 (N_1935,N_1902,N_1887);
or U1936 (N_1936,N_1862,N_1867);
nor U1937 (N_1937,N_1893,N_1883);
nor U1938 (N_1938,N_1909,N_1868);
and U1939 (N_1939,N_1899,N_1882);
nand U1940 (N_1940,N_1874,N_1888);
and U1941 (N_1941,N_1873,N_1908);
and U1942 (N_1942,N_1901,N_1895);
or U1943 (N_1943,N_1875,N_1860);
and U1944 (N_1944,N_1871,N_1879);
nor U1945 (N_1945,N_1905,N_1865);
or U1946 (N_1946,N_1919,N_1894);
nor U1947 (N_1947,N_1913,N_1915);
xor U1948 (N_1948,N_1896,N_1866);
nor U1949 (N_1949,N_1904,N_1885);
and U1950 (N_1950,N_1862,N_1875);
nand U1951 (N_1951,N_1862,N_1899);
and U1952 (N_1952,N_1883,N_1868);
nand U1953 (N_1953,N_1909,N_1866);
or U1954 (N_1954,N_1873,N_1910);
or U1955 (N_1955,N_1896,N_1870);
and U1956 (N_1956,N_1878,N_1877);
and U1957 (N_1957,N_1885,N_1871);
nand U1958 (N_1958,N_1897,N_1904);
xnor U1959 (N_1959,N_1884,N_1889);
and U1960 (N_1960,N_1914,N_1918);
or U1961 (N_1961,N_1885,N_1895);
or U1962 (N_1962,N_1871,N_1883);
and U1963 (N_1963,N_1880,N_1919);
nor U1964 (N_1964,N_1876,N_1896);
nand U1965 (N_1965,N_1910,N_1898);
or U1966 (N_1966,N_1901,N_1902);
and U1967 (N_1967,N_1906,N_1882);
nand U1968 (N_1968,N_1892,N_1861);
nand U1969 (N_1969,N_1888,N_1865);
or U1970 (N_1970,N_1865,N_1899);
nand U1971 (N_1971,N_1874,N_1895);
and U1972 (N_1972,N_1886,N_1911);
nor U1973 (N_1973,N_1888,N_1887);
nand U1974 (N_1974,N_1887,N_1910);
nor U1975 (N_1975,N_1891,N_1916);
nand U1976 (N_1976,N_1916,N_1919);
and U1977 (N_1977,N_1889,N_1862);
and U1978 (N_1978,N_1884,N_1886);
xor U1979 (N_1979,N_1887,N_1899);
or U1980 (N_1980,N_1965,N_1975);
nand U1981 (N_1981,N_1976,N_1932);
or U1982 (N_1982,N_1974,N_1979);
or U1983 (N_1983,N_1946,N_1920);
nand U1984 (N_1984,N_1960,N_1930);
and U1985 (N_1985,N_1937,N_1933);
nor U1986 (N_1986,N_1934,N_1954);
nor U1987 (N_1987,N_1953,N_1944);
and U1988 (N_1988,N_1941,N_1942);
nor U1989 (N_1989,N_1951,N_1977);
nand U1990 (N_1990,N_1931,N_1927);
nor U1991 (N_1991,N_1962,N_1968);
nand U1992 (N_1992,N_1926,N_1972);
and U1993 (N_1993,N_1938,N_1956);
and U1994 (N_1994,N_1961,N_1969);
and U1995 (N_1995,N_1955,N_1967);
and U1996 (N_1996,N_1947,N_1959);
nor U1997 (N_1997,N_1964,N_1921);
and U1998 (N_1998,N_1945,N_1923);
and U1999 (N_1999,N_1948,N_1939);
nand U2000 (N_2000,N_1924,N_1928);
and U2001 (N_2001,N_1958,N_1957);
xor U2002 (N_2002,N_1935,N_1970);
xor U2003 (N_2003,N_1973,N_1925);
or U2004 (N_2004,N_1966,N_1922);
and U2005 (N_2005,N_1971,N_1978);
or U2006 (N_2006,N_1949,N_1936);
and U2007 (N_2007,N_1950,N_1963);
nand U2008 (N_2008,N_1952,N_1940);
or U2009 (N_2009,N_1929,N_1943);
or U2010 (N_2010,N_1920,N_1953);
nand U2011 (N_2011,N_1973,N_1922);
nor U2012 (N_2012,N_1969,N_1921);
nand U2013 (N_2013,N_1960,N_1941);
nand U2014 (N_2014,N_1944,N_1960);
or U2015 (N_2015,N_1920,N_1963);
or U2016 (N_2016,N_1962,N_1951);
or U2017 (N_2017,N_1927,N_1952);
or U2018 (N_2018,N_1955,N_1971);
and U2019 (N_2019,N_1934,N_1971);
or U2020 (N_2020,N_1964,N_1943);
nand U2021 (N_2021,N_1952,N_1979);
nand U2022 (N_2022,N_1946,N_1970);
and U2023 (N_2023,N_1978,N_1954);
and U2024 (N_2024,N_1951,N_1959);
and U2025 (N_2025,N_1926,N_1953);
nand U2026 (N_2026,N_1945,N_1939);
xor U2027 (N_2027,N_1927,N_1955);
or U2028 (N_2028,N_1940,N_1938);
nand U2029 (N_2029,N_1960,N_1925);
nand U2030 (N_2030,N_1964,N_1930);
nor U2031 (N_2031,N_1960,N_1942);
nor U2032 (N_2032,N_1936,N_1946);
or U2033 (N_2033,N_1967,N_1942);
and U2034 (N_2034,N_1929,N_1921);
and U2035 (N_2035,N_1972,N_1947);
xnor U2036 (N_2036,N_1969,N_1970);
nor U2037 (N_2037,N_1931,N_1975);
nand U2038 (N_2038,N_1950,N_1955);
nand U2039 (N_2039,N_1941,N_1939);
nor U2040 (N_2040,N_2038,N_2005);
or U2041 (N_2041,N_1991,N_2006);
nor U2042 (N_2042,N_2015,N_1981);
nand U2043 (N_2043,N_2001,N_2000);
and U2044 (N_2044,N_1984,N_1983);
nor U2045 (N_2045,N_2030,N_1982);
xnor U2046 (N_2046,N_2035,N_1985);
xnor U2047 (N_2047,N_2011,N_2024);
nor U2048 (N_2048,N_1995,N_1988);
or U2049 (N_2049,N_2034,N_2021);
and U2050 (N_2050,N_1996,N_2022);
and U2051 (N_2051,N_1987,N_2014);
or U2052 (N_2052,N_1993,N_2023);
and U2053 (N_2053,N_1990,N_2009);
and U2054 (N_2054,N_1994,N_1989);
or U2055 (N_2055,N_2002,N_2039);
or U2056 (N_2056,N_2032,N_2029);
or U2057 (N_2057,N_1999,N_2025);
xor U2058 (N_2058,N_2037,N_2027);
nor U2059 (N_2059,N_2004,N_1998);
xnor U2060 (N_2060,N_2008,N_2026);
or U2061 (N_2061,N_2031,N_1997);
nor U2062 (N_2062,N_2003,N_2036);
nand U2063 (N_2063,N_2028,N_2010);
or U2064 (N_2064,N_2017,N_2020);
or U2065 (N_2065,N_1986,N_2012);
nand U2066 (N_2066,N_2019,N_2033);
xnor U2067 (N_2067,N_1980,N_2007);
nor U2068 (N_2068,N_2016,N_2013);
and U2069 (N_2069,N_1992,N_2018);
nor U2070 (N_2070,N_2005,N_2007);
or U2071 (N_2071,N_2023,N_2014);
nor U2072 (N_2072,N_1981,N_2028);
or U2073 (N_2073,N_2010,N_1992);
and U2074 (N_2074,N_2010,N_2007);
and U2075 (N_2075,N_1988,N_2012);
or U2076 (N_2076,N_1993,N_2013);
nand U2077 (N_2077,N_1981,N_2018);
or U2078 (N_2078,N_1996,N_2033);
or U2079 (N_2079,N_2001,N_2028);
or U2080 (N_2080,N_2002,N_2021);
and U2081 (N_2081,N_1997,N_2000);
or U2082 (N_2082,N_2021,N_1980);
or U2083 (N_2083,N_2036,N_1998);
or U2084 (N_2084,N_1997,N_2007);
and U2085 (N_2085,N_2020,N_2019);
nor U2086 (N_2086,N_2034,N_1987);
or U2087 (N_2087,N_1986,N_1999);
nand U2088 (N_2088,N_2038,N_2007);
and U2089 (N_2089,N_1988,N_1982);
xnor U2090 (N_2090,N_2032,N_2009);
or U2091 (N_2091,N_2004,N_2025);
xor U2092 (N_2092,N_2007,N_2018);
and U2093 (N_2093,N_1990,N_1981);
nand U2094 (N_2094,N_1989,N_2023);
xor U2095 (N_2095,N_1980,N_1982);
or U2096 (N_2096,N_2021,N_2029);
nor U2097 (N_2097,N_1980,N_1984);
or U2098 (N_2098,N_1996,N_2017);
or U2099 (N_2099,N_1990,N_2034);
nand U2100 (N_2100,N_2040,N_2094);
and U2101 (N_2101,N_2046,N_2044);
and U2102 (N_2102,N_2099,N_2059);
and U2103 (N_2103,N_2070,N_2056);
and U2104 (N_2104,N_2062,N_2081);
nor U2105 (N_2105,N_2093,N_2052);
nor U2106 (N_2106,N_2078,N_2088);
nor U2107 (N_2107,N_2091,N_2050);
nand U2108 (N_2108,N_2041,N_2077);
or U2109 (N_2109,N_2064,N_2048);
or U2110 (N_2110,N_2072,N_2075);
and U2111 (N_2111,N_2061,N_2082);
and U2112 (N_2112,N_2067,N_2085);
nand U2113 (N_2113,N_2066,N_2060);
nand U2114 (N_2114,N_2045,N_2095);
nor U2115 (N_2115,N_2092,N_2084);
nor U2116 (N_2116,N_2053,N_2047);
and U2117 (N_2117,N_2089,N_2058);
xor U2118 (N_2118,N_2096,N_2063);
xor U2119 (N_2119,N_2068,N_2069);
or U2120 (N_2120,N_2086,N_2079);
nand U2121 (N_2121,N_2051,N_2097);
and U2122 (N_2122,N_2055,N_2071);
xor U2123 (N_2123,N_2080,N_2057);
nor U2124 (N_2124,N_2054,N_2074);
and U2125 (N_2125,N_2049,N_2073);
and U2126 (N_2126,N_2043,N_2083);
and U2127 (N_2127,N_2042,N_2098);
and U2128 (N_2128,N_2076,N_2065);
nor U2129 (N_2129,N_2090,N_2087);
and U2130 (N_2130,N_2089,N_2042);
nor U2131 (N_2131,N_2080,N_2067);
or U2132 (N_2132,N_2091,N_2053);
nor U2133 (N_2133,N_2085,N_2083);
or U2134 (N_2134,N_2047,N_2068);
and U2135 (N_2135,N_2058,N_2067);
xor U2136 (N_2136,N_2088,N_2097);
and U2137 (N_2137,N_2067,N_2045);
nor U2138 (N_2138,N_2078,N_2071);
or U2139 (N_2139,N_2085,N_2088);
and U2140 (N_2140,N_2090,N_2081);
nand U2141 (N_2141,N_2049,N_2057);
or U2142 (N_2142,N_2088,N_2046);
or U2143 (N_2143,N_2092,N_2061);
nor U2144 (N_2144,N_2059,N_2053);
or U2145 (N_2145,N_2074,N_2051);
nor U2146 (N_2146,N_2090,N_2091);
nor U2147 (N_2147,N_2069,N_2063);
nor U2148 (N_2148,N_2041,N_2056);
and U2149 (N_2149,N_2082,N_2078);
nor U2150 (N_2150,N_2044,N_2047);
nand U2151 (N_2151,N_2066,N_2046);
nor U2152 (N_2152,N_2049,N_2059);
nand U2153 (N_2153,N_2044,N_2072);
nand U2154 (N_2154,N_2061,N_2081);
or U2155 (N_2155,N_2080,N_2046);
or U2156 (N_2156,N_2044,N_2060);
nor U2157 (N_2157,N_2077,N_2046);
and U2158 (N_2158,N_2083,N_2063);
nand U2159 (N_2159,N_2077,N_2049);
nor U2160 (N_2160,N_2151,N_2112);
nor U2161 (N_2161,N_2149,N_2148);
or U2162 (N_2162,N_2104,N_2159);
xor U2163 (N_2163,N_2126,N_2125);
nand U2164 (N_2164,N_2120,N_2115);
and U2165 (N_2165,N_2155,N_2152);
xnor U2166 (N_2166,N_2106,N_2103);
and U2167 (N_2167,N_2129,N_2135);
nand U2168 (N_2168,N_2145,N_2102);
and U2169 (N_2169,N_2124,N_2131);
xnor U2170 (N_2170,N_2113,N_2146);
or U2171 (N_2171,N_2144,N_2111);
or U2172 (N_2172,N_2110,N_2138);
or U2173 (N_2173,N_2100,N_2107);
nor U2174 (N_2174,N_2157,N_2123);
nor U2175 (N_2175,N_2122,N_2143);
and U2176 (N_2176,N_2117,N_2109);
nand U2177 (N_2177,N_2133,N_2136);
xor U2178 (N_2178,N_2130,N_2101);
nor U2179 (N_2179,N_2105,N_2153);
xor U2180 (N_2180,N_2139,N_2127);
or U2181 (N_2181,N_2158,N_2128);
and U2182 (N_2182,N_2150,N_2116);
nor U2183 (N_2183,N_2118,N_2121);
nor U2184 (N_2184,N_2147,N_2140);
nor U2185 (N_2185,N_2137,N_2134);
or U2186 (N_2186,N_2156,N_2141);
nand U2187 (N_2187,N_2142,N_2108);
or U2188 (N_2188,N_2154,N_2132);
and U2189 (N_2189,N_2119,N_2114);
nor U2190 (N_2190,N_2152,N_2110);
nor U2191 (N_2191,N_2134,N_2147);
and U2192 (N_2192,N_2106,N_2136);
and U2193 (N_2193,N_2116,N_2128);
nor U2194 (N_2194,N_2112,N_2126);
nor U2195 (N_2195,N_2110,N_2136);
nor U2196 (N_2196,N_2103,N_2130);
nor U2197 (N_2197,N_2110,N_2155);
xor U2198 (N_2198,N_2106,N_2121);
xor U2199 (N_2199,N_2140,N_2134);
and U2200 (N_2200,N_2132,N_2131);
and U2201 (N_2201,N_2139,N_2156);
or U2202 (N_2202,N_2143,N_2121);
nand U2203 (N_2203,N_2109,N_2142);
and U2204 (N_2204,N_2138,N_2157);
nand U2205 (N_2205,N_2112,N_2141);
or U2206 (N_2206,N_2116,N_2156);
and U2207 (N_2207,N_2144,N_2153);
or U2208 (N_2208,N_2102,N_2112);
xor U2209 (N_2209,N_2119,N_2103);
and U2210 (N_2210,N_2119,N_2159);
nor U2211 (N_2211,N_2152,N_2139);
nand U2212 (N_2212,N_2103,N_2136);
or U2213 (N_2213,N_2114,N_2151);
nor U2214 (N_2214,N_2130,N_2124);
nand U2215 (N_2215,N_2125,N_2145);
or U2216 (N_2216,N_2154,N_2121);
nand U2217 (N_2217,N_2110,N_2102);
and U2218 (N_2218,N_2146,N_2157);
or U2219 (N_2219,N_2115,N_2127);
or U2220 (N_2220,N_2185,N_2176);
nand U2221 (N_2221,N_2192,N_2164);
xor U2222 (N_2222,N_2194,N_2208);
nand U2223 (N_2223,N_2219,N_2177);
nand U2224 (N_2224,N_2183,N_2211);
nor U2225 (N_2225,N_2165,N_2178);
nand U2226 (N_2226,N_2166,N_2171);
nor U2227 (N_2227,N_2187,N_2170);
nor U2228 (N_2228,N_2213,N_2200);
or U2229 (N_2229,N_2190,N_2169);
and U2230 (N_2230,N_2180,N_2172);
xor U2231 (N_2231,N_2209,N_2174);
or U2232 (N_2232,N_2163,N_2201);
nor U2233 (N_2233,N_2161,N_2212);
nor U2234 (N_2234,N_2195,N_2218);
nor U2235 (N_2235,N_2175,N_2210);
nor U2236 (N_2236,N_2206,N_2217);
or U2237 (N_2237,N_2207,N_2197);
or U2238 (N_2238,N_2189,N_2188);
nor U2239 (N_2239,N_2202,N_2215);
or U2240 (N_2240,N_2199,N_2182);
xor U2241 (N_2241,N_2179,N_2214);
nor U2242 (N_2242,N_2184,N_2204);
nor U2243 (N_2243,N_2160,N_2181);
xor U2244 (N_2244,N_2216,N_2186);
and U2245 (N_2245,N_2205,N_2191);
xnor U2246 (N_2246,N_2168,N_2203);
nand U2247 (N_2247,N_2196,N_2193);
xor U2248 (N_2248,N_2167,N_2173);
nor U2249 (N_2249,N_2162,N_2198);
nor U2250 (N_2250,N_2166,N_2175);
and U2251 (N_2251,N_2183,N_2203);
or U2252 (N_2252,N_2197,N_2215);
xnor U2253 (N_2253,N_2190,N_2185);
or U2254 (N_2254,N_2160,N_2170);
nor U2255 (N_2255,N_2166,N_2207);
nor U2256 (N_2256,N_2204,N_2165);
nand U2257 (N_2257,N_2209,N_2214);
and U2258 (N_2258,N_2197,N_2177);
or U2259 (N_2259,N_2201,N_2196);
or U2260 (N_2260,N_2175,N_2169);
or U2261 (N_2261,N_2167,N_2179);
and U2262 (N_2262,N_2209,N_2189);
xor U2263 (N_2263,N_2192,N_2205);
or U2264 (N_2264,N_2184,N_2181);
or U2265 (N_2265,N_2203,N_2199);
and U2266 (N_2266,N_2191,N_2219);
or U2267 (N_2267,N_2171,N_2213);
nand U2268 (N_2268,N_2214,N_2199);
xor U2269 (N_2269,N_2166,N_2211);
nor U2270 (N_2270,N_2206,N_2219);
nor U2271 (N_2271,N_2172,N_2168);
and U2272 (N_2272,N_2177,N_2212);
nor U2273 (N_2273,N_2199,N_2204);
and U2274 (N_2274,N_2164,N_2169);
nand U2275 (N_2275,N_2196,N_2163);
or U2276 (N_2276,N_2189,N_2218);
nor U2277 (N_2277,N_2166,N_2214);
nand U2278 (N_2278,N_2196,N_2208);
nor U2279 (N_2279,N_2214,N_2185);
xor U2280 (N_2280,N_2243,N_2249);
and U2281 (N_2281,N_2255,N_2226);
nand U2282 (N_2282,N_2244,N_2273);
nand U2283 (N_2283,N_2235,N_2265);
or U2284 (N_2284,N_2271,N_2223);
or U2285 (N_2285,N_2240,N_2261);
or U2286 (N_2286,N_2251,N_2231);
or U2287 (N_2287,N_2245,N_2247);
nor U2288 (N_2288,N_2242,N_2275);
nand U2289 (N_2289,N_2250,N_2246);
nor U2290 (N_2290,N_2279,N_2277);
nor U2291 (N_2291,N_2238,N_2239);
or U2292 (N_2292,N_2264,N_2259);
or U2293 (N_2293,N_2224,N_2260);
nand U2294 (N_2294,N_2272,N_2254);
nand U2295 (N_2295,N_2262,N_2241);
or U2296 (N_2296,N_2268,N_2225);
or U2297 (N_2297,N_2252,N_2221);
nor U2298 (N_2298,N_2236,N_2227);
and U2299 (N_2299,N_2269,N_2270);
nor U2300 (N_2300,N_2248,N_2274);
and U2301 (N_2301,N_2222,N_2253);
and U2302 (N_2302,N_2258,N_2257);
nor U2303 (N_2303,N_2230,N_2229);
and U2304 (N_2304,N_2256,N_2266);
and U2305 (N_2305,N_2228,N_2233);
or U2306 (N_2306,N_2267,N_2234);
xnor U2307 (N_2307,N_2278,N_2220);
nor U2308 (N_2308,N_2232,N_2237);
and U2309 (N_2309,N_2263,N_2276);
nand U2310 (N_2310,N_2255,N_2230);
and U2311 (N_2311,N_2240,N_2239);
or U2312 (N_2312,N_2225,N_2265);
nor U2313 (N_2313,N_2241,N_2278);
or U2314 (N_2314,N_2242,N_2267);
xnor U2315 (N_2315,N_2238,N_2240);
and U2316 (N_2316,N_2258,N_2236);
nand U2317 (N_2317,N_2254,N_2247);
nor U2318 (N_2318,N_2232,N_2243);
and U2319 (N_2319,N_2258,N_2222);
nand U2320 (N_2320,N_2262,N_2274);
nand U2321 (N_2321,N_2229,N_2279);
and U2322 (N_2322,N_2232,N_2249);
nor U2323 (N_2323,N_2258,N_2249);
and U2324 (N_2324,N_2279,N_2240);
nor U2325 (N_2325,N_2235,N_2246);
nor U2326 (N_2326,N_2240,N_2229);
nor U2327 (N_2327,N_2270,N_2232);
or U2328 (N_2328,N_2224,N_2222);
and U2329 (N_2329,N_2248,N_2250);
or U2330 (N_2330,N_2229,N_2246);
or U2331 (N_2331,N_2239,N_2255);
xnor U2332 (N_2332,N_2230,N_2227);
nand U2333 (N_2333,N_2239,N_2279);
nor U2334 (N_2334,N_2255,N_2279);
nand U2335 (N_2335,N_2252,N_2241);
or U2336 (N_2336,N_2247,N_2250);
nand U2337 (N_2337,N_2249,N_2264);
nand U2338 (N_2338,N_2238,N_2233);
and U2339 (N_2339,N_2236,N_2263);
xor U2340 (N_2340,N_2301,N_2287);
nand U2341 (N_2341,N_2336,N_2330);
and U2342 (N_2342,N_2302,N_2296);
and U2343 (N_2343,N_2319,N_2289);
or U2344 (N_2344,N_2324,N_2295);
or U2345 (N_2345,N_2290,N_2305);
nand U2346 (N_2346,N_2299,N_2328);
and U2347 (N_2347,N_2282,N_2292);
nor U2348 (N_2348,N_2313,N_2312);
and U2349 (N_2349,N_2283,N_2280);
or U2350 (N_2350,N_2311,N_2297);
and U2351 (N_2351,N_2318,N_2309);
and U2352 (N_2352,N_2284,N_2285);
and U2353 (N_2353,N_2322,N_2329);
and U2354 (N_2354,N_2288,N_2294);
or U2355 (N_2355,N_2315,N_2326);
xor U2356 (N_2356,N_2335,N_2310);
or U2357 (N_2357,N_2281,N_2331);
and U2358 (N_2358,N_2293,N_2338);
nand U2359 (N_2359,N_2304,N_2325);
nor U2360 (N_2360,N_2306,N_2321);
nand U2361 (N_2361,N_2314,N_2286);
nor U2362 (N_2362,N_2337,N_2320);
nor U2363 (N_2363,N_2291,N_2303);
xnor U2364 (N_2364,N_2332,N_2316);
xnor U2365 (N_2365,N_2307,N_2308);
and U2366 (N_2366,N_2317,N_2339);
xor U2367 (N_2367,N_2334,N_2327);
nor U2368 (N_2368,N_2298,N_2333);
or U2369 (N_2369,N_2300,N_2323);
and U2370 (N_2370,N_2282,N_2324);
nor U2371 (N_2371,N_2329,N_2306);
or U2372 (N_2372,N_2283,N_2314);
nand U2373 (N_2373,N_2338,N_2313);
nand U2374 (N_2374,N_2283,N_2288);
nor U2375 (N_2375,N_2301,N_2319);
nand U2376 (N_2376,N_2280,N_2326);
nand U2377 (N_2377,N_2317,N_2310);
or U2378 (N_2378,N_2321,N_2285);
nor U2379 (N_2379,N_2313,N_2302);
and U2380 (N_2380,N_2305,N_2291);
nand U2381 (N_2381,N_2334,N_2312);
nor U2382 (N_2382,N_2317,N_2333);
and U2383 (N_2383,N_2332,N_2300);
and U2384 (N_2384,N_2303,N_2312);
or U2385 (N_2385,N_2337,N_2284);
or U2386 (N_2386,N_2307,N_2296);
nand U2387 (N_2387,N_2298,N_2338);
nand U2388 (N_2388,N_2335,N_2331);
or U2389 (N_2389,N_2283,N_2292);
and U2390 (N_2390,N_2299,N_2294);
nand U2391 (N_2391,N_2299,N_2298);
nor U2392 (N_2392,N_2329,N_2318);
nand U2393 (N_2393,N_2329,N_2295);
nor U2394 (N_2394,N_2318,N_2333);
nor U2395 (N_2395,N_2282,N_2306);
nand U2396 (N_2396,N_2319,N_2322);
and U2397 (N_2397,N_2300,N_2297);
nor U2398 (N_2398,N_2280,N_2303);
nor U2399 (N_2399,N_2334,N_2304);
xor U2400 (N_2400,N_2346,N_2347);
nand U2401 (N_2401,N_2391,N_2349);
and U2402 (N_2402,N_2350,N_2352);
nand U2403 (N_2403,N_2388,N_2393);
or U2404 (N_2404,N_2390,N_2360);
and U2405 (N_2405,N_2354,N_2387);
nor U2406 (N_2406,N_2340,N_2368);
nor U2407 (N_2407,N_2385,N_2392);
and U2408 (N_2408,N_2364,N_2344);
and U2409 (N_2409,N_2359,N_2365);
or U2410 (N_2410,N_2351,N_2374);
or U2411 (N_2411,N_2372,N_2371);
and U2412 (N_2412,N_2355,N_2343);
nand U2413 (N_2413,N_2397,N_2399);
or U2414 (N_2414,N_2348,N_2353);
nand U2415 (N_2415,N_2361,N_2378);
nand U2416 (N_2416,N_2363,N_2381);
nand U2417 (N_2417,N_2369,N_2376);
or U2418 (N_2418,N_2380,N_2357);
nor U2419 (N_2419,N_2373,N_2377);
nor U2420 (N_2420,N_2362,N_2367);
and U2421 (N_2421,N_2342,N_2382);
nor U2422 (N_2422,N_2395,N_2384);
nor U2423 (N_2423,N_2370,N_2366);
nand U2424 (N_2424,N_2345,N_2398);
nor U2425 (N_2425,N_2389,N_2356);
or U2426 (N_2426,N_2358,N_2394);
and U2427 (N_2427,N_2375,N_2383);
nor U2428 (N_2428,N_2396,N_2379);
and U2429 (N_2429,N_2341,N_2386);
nand U2430 (N_2430,N_2372,N_2350);
nand U2431 (N_2431,N_2380,N_2351);
nand U2432 (N_2432,N_2393,N_2358);
nor U2433 (N_2433,N_2399,N_2345);
and U2434 (N_2434,N_2377,N_2351);
nor U2435 (N_2435,N_2394,N_2393);
and U2436 (N_2436,N_2358,N_2372);
nor U2437 (N_2437,N_2384,N_2387);
and U2438 (N_2438,N_2384,N_2352);
or U2439 (N_2439,N_2384,N_2392);
nor U2440 (N_2440,N_2375,N_2396);
nand U2441 (N_2441,N_2371,N_2380);
and U2442 (N_2442,N_2345,N_2379);
and U2443 (N_2443,N_2368,N_2399);
xnor U2444 (N_2444,N_2346,N_2381);
or U2445 (N_2445,N_2377,N_2399);
or U2446 (N_2446,N_2366,N_2346);
and U2447 (N_2447,N_2363,N_2344);
and U2448 (N_2448,N_2373,N_2346);
xor U2449 (N_2449,N_2347,N_2364);
xnor U2450 (N_2450,N_2374,N_2362);
nand U2451 (N_2451,N_2353,N_2363);
nand U2452 (N_2452,N_2368,N_2374);
and U2453 (N_2453,N_2351,N_2386);
or U2454 (N_2454,N_2385,N_2384);
nor U2455 (N_2455,N_2362,N_2360);
xnor U2456 (N_2456,N_2341,N_2393);
or U2457 (N_2457,N_2390,N_2362);
xnor U2458 (N_2458,N_2343,N_2352);
and U2459 (N_2459,N_2361,N_2372);
and U2460 (N_2460,N_2440,N_2431);
nand U2461 (N_2461,N_2405,N_2439);
and U2462 (N_2462,N_2451,N_2423);
and U2463 (N_2463,N_2419,N_2415);
nor U2464 (N_2464,N_2441,N_2456);
nor U2465 (N_2465,N_2420,N_2442);
and U2466 (N_2466,N_2453,N_2414);
nor U2467 (N_2467,N_2402,N_2455);
nand U2468 (N_2468,N_2412,N_2406);
or U2469 (N_2469,N_2434,N_2404);
xor U2470 (N_2470,N_2408,N_2432);
and U2471 (N_2471,N_2433,N_2435);
nor U2472 (N_2472,N_2413,N_2403);
or U2473 (N_2473,N_2422,N_2409);
nor U2474 (N_2474,N_2416,N_2400);
nand U2475 (N_2475,N_2436,N_2444);
or U2476 (N_2476,N_2430,N_2454);
and U2477 (N_2477,N_2418,N_2428);
and U2478 (N_2478,N_2452,N_2443);
xor U2479 (N_2479,N_2446,N_2410);
and U2480 (N_2480,N_2401,N_2421);
nor U2481 (N_2481,N_2438,N_2458);
nor U2482 (N_2482,N_2429,N_2447);
xnor U2483 (N_2483,N_2457,N_2459);
or U2484 (N_2484,N_2445,N_2437);
and U2485 (N_2485,N_2424,N_2425);
and U2486 (N_2486,N_2449,N_2450);
nand U2487 (N_2487,N_2411,N_2426);
xnor U2488 (N_2488,N_2417,N_2448);
nor U2489 (N_2489,N_2427,N_2407);
xnor U2490 (N_2490,N_2412,N_2414);
nor U2491 (N_2491,N_2416,N_2441);
or U2492 (N_2492,N_2405,N_2422);
nor U2493 (N_2493,N_2431,N_2433);
or U2494 (N_2494,N_2435,N_2432);
nand U2495 (N_2495,N_2402,N_2445);
nand U2496 (N_2496,N_2435,N_2428);
and U2497 (N_2497,N_2435,N_2416);
and U2498 (N_2498,N_2442,N_2407);
nor U2499 (N_2499,N_2404,N_2408);
nand U2500 (N_2500,N_2452,N_2426);
xnor U2501 (N_2501,N_2417,N_2432);
nor U2502 (N_2502,N_2456,N_2415);
nor U2503 (N_2503,N_2433,N_2408);
and U2504 (N_2504,N_2401,N_2406);
or U2505 (N_2505,N_2432,N_2426);
and U2506 (N_2506,N_2443,N_2444);
nand U2507 (N_2507,N_2406,N_2448);
xor U2508 (N_2508,N_2419,N_2405);
or U2509 (N_2509,N_2414,N_2437);
and U2510 (N_2510,N_2427,N_2415);
nor U2511 (N_2511,N_2421,N_2457);
nand U2512 (N_2512,N_2437,N_2424);
nor U2513 (N_2513,N_2414,N_2433);
and U2514 (N_2514,N_2429,N_2453);
and U2515 (N_2515,N_2448,N_2445);
and U2516 (N_2516,N_2411,N_2444);
and U2517 (N_2517,N_2400,N_2422);
or U2518 (N_2518,N_2419,N_2454);
or U2519 (N_2519,N_2452,N_2453);
or U2520 (N_2520,N_2466,N_2472);
nor U2521 (N_2521,N_2479,N_2492);
nor U2522 (N_2522,N_2462,N_2483);
or U2523 (N_2523,N_2486,N_2475);
nand U2524 (N_2524,N_2504,N_2482);
or U2525 (N_2525,N_2495,N_2480);
nand U2526 (N_2526,N_2510,N_2508);
nor U2527 (N_2527,N_2516,N_2471);
or U2528 (N_2528,N_2503,N_2474);
nand U2529 (N_2529,N_2499,N_2481);
or U2530 (N_2530,N_2497,N_2493);
and U2531 (N_2531,N_2476,N_2487);
nand U2532 (N_2532,N_2488,N_2496);
nand U2533 (N_2533,N_2511,N_2512);
nor U2534 (N_2534,N_2498,N_2467);
and U2535 (N_2535,N_2460,N_2478);
nand U2536 (N_2536,N_2517,N_2485);
nand U2537 (N_2537,N_2473,N_2505);
or U2538 (N_2538,N_2464,N_2509);
and U2539 (N_2539,N_2469,N_2489);
or U2540 (N_2540,N_2500,N_2519);
nor U2541 (N_2541,N_2501,N_2513);
nor U2542 (N_2542,N_2490,N_2470);
or U2543 (N_2543,N_2465,N_2518);
xnor U2544 (N_2544,N_2502,N_2491);
and U2545 (N_2545,N_2494,N_2506);
and U2546 (N_2546,N_2507,N_2515);
nor U2547 (N_2547,N_2477,N_2484);
or U2548 (N_2548,N_2461,N_2468);
and U2549 (N_2549,N_2514,N_2463);
and U2550 (N_2550,N_2481,N_2519);
nand U2551 (N_2551,N_2507,N_2513);
and U2552 (N_2552,N_2490,N_2480);
nor U2553 (N_2553,N_2492,N_2500);
or U2554 (N_2554,N_2466,N_2491);
or U2555 (N_2555,N_2483,N_2489);
or U2556 (N_2556,N_2476,N_2519);
nand U2557 (N_2557,N_2474,N_2517);
xnor U2558 (N_2558,N_2483,N_2464);
and U2559 (N_2559,N_2482,N_2515);
and U2560 (N_2560,N_2474,N_2507);
or U2561 (N_2561,N_2470,N_2496);
nor U2562 (N_2562,N_2514,N_2518);
or U2563 (N_2563,N_2491,N_2461);
and U2564 (N_2564,N_2503,N_2462);
xnor U2565 (N_2565,N_2467,N_2472);
and U2566 (N_2566,N_2495,N_2505);
nand U2567 (N_2567,N_2473,N_2501);
nand U2568 (N_2568,N_2517,N_2464);
nand U2569 (N_2569,N_2511,N_2461);
nand U2570 (N_2570,N_2482,N_2502);
nor U2571 (N_2571,N_2475,N_2507);
nand U2572 (N_2572,N_2461,N_2515);
or U2573 (N_2573,N_2516,N_2478);
nand U2574 (N_2574,N_2505,N_2488);
and U2575 (N_2575,N_2468,N_2519);
nor U2576 (N_2576,N_2485,N_2518);
nand U2577 (N_2577,N_2500,N_2468);
and U2578 (N_2578,N_2496,N_2494);
or U2579 (N_2579,N_2484,N_2489);
and U2580 (N_2580,N_2559,N_2538);
xnor U2581 (N_2581,N_2539,N_2526);
nand U2582 (N_2582,N_2577,N_2529);
or U2583 (N_2583,N_2569,N_2530);
nor U2584 (N_2584,N_2543,N_2522);
or U2585 (N_2585,N_2570,N_2557);
nand U2586 (N_2586,N_2561,N_2562);
nor U2587 (N_2587,N_2533,N_2551);
and U2588 (N_2588,N_2524,N_2550);
or U2589 (N_2589,N_2520,N_2531);
nand U2590 (N_2590,N_2536,N_2548);
and U2591 (N_2591,N_2560,N_2556);
nand U2592 (N_2592,N_2571,N_2537);
nand U2593 (N_2593,N_2534,N_2567);
nand U2594 (N_2594,N_2552,N_2549);
and U2595 (N_2595,N_2558,N_2554);
and U2596 (N_2596,N_2523,N_2573);
nand U2597 (N_2597,N_2545,N_2525);
nor U2598 (N_2598,N_2532,N_2544);
nor U2599 (N_2599,N_2574,N_2578);
nand U2600 (N_2600,N_2528,N_2541);
nand U2601 (N_2601,N_2579,N_2568);
nor U2602 (N_2602,N_2542,N_2535);
and U2603 (N_2603,N_2565,N_2566);
nand U2604 (N_2604,N_2572,N_2553);
nand U2605 (N_2605,N_2555,N_2576);
or U2606 (N_2606,N_2540,N_2547);
nand U2607 (N_2607,N_2546,N_2564);
nor U2608 (N_2608,N_2563,N_2575);
nor U2609 (N_2609,N_2521,N_2527);
and U2610 (N_2610,N_2564,N_2522);
or U2611 (N_2611,N_2540,N_2543);
nand U2612 (N_2612,N_2536,N_2539);
nand U2613 (N_2613,N_2556,N_2572);
nand U2614 (N_2614,N_2566,N_2560);
nand U2615 (N_2615,N_2523,N_2549);
nor U2616 (N_2616,N_2527,N_2576);
and U2617 (N_2617,N_2579,N_2555);
xor U2618 (N_2618,N_2561,N_2529);
nand U2619 (N_2619,N_2564,N_2571);
and U2620 (N_2620,N_2526,N_2579);
nor U2621 (N_2621,N_2536,N_2555);
xor U2622 (N_2622,N_2572,N_2574);
or U2623 (N_2623,N_2531,N_2552);
nor U2624 (N_2624,N_2574,N_2522);
nor U2625 (N_2625,N_2530,N_2543);
nand U2626 (N_2626,N_2562,N_2540);
nor U2627 (N_2627,N_2559,N_2560);
or U2628 (N_2628,N_2579,N_2569);
nand U2629 (N_2629,N_2543,N_2525);
nor U2630 (N_2630,N_2567,N_2559);
nor U2631 (N_2631,N_2541,N_2543);
xor U2632 (N_2632,N_2569,N_2574);
and U2633 (N_2633,N_2562,N_2563);
xnor U2634 (N_2634,N_2553,N_2579);
nand U2635 (N_2635,N_2573,N_2567);
or U2636 (N_2636,N_2521,N_2552);
xnor U2637 (N_2637,N_2556,N_2554);
nand U2638 (N_2638,N_2527,N_2575);
nor U2639 (N_2639,N_2568,N_2548);
nand U2640 (N_2640,N_2584,N_2590);
xnor U2641 (N_2641,N_2614,N_2581);
nand U2642 (N_2642,N_2595,N_2600);
or U2643 (N_2643,N_2635,N_2612);
and U2644 (N_2644,N_2637,N_2632);
nor U2645 (N_2645,N_2624,N_2607);
and U2646 (N_2646,N_2628,N_2602);
or U2647 (N_2647,N_2582,N_2620);
and U2648 (N_2648,N_2585,N_2601);
nand U2649 (N_2649,N_2604,N_2605);
nand U2650 (N_2650,N_2588,N_2613);
or U2651 (N_2651,N_2597,N_2610);
nand U2652 (N_2652,N_2603,N_2587);
or U2653 (N_2653,N_2621,N_2591);
nor U2654 (N_2654,N_2625,N_2599);
and U2655 (N_2655,N_2615,N_2611);
or U2656 (N_2656,N_2580,N_2609);
nor U2657 (N_2657,N_2606,N_2638);
nor U2658 (N_2658,N_2633,N_2631);
or U2659 (N_2659,N_2629,N_2636);
nand U2660 (N_2660,N_2619,N_2596);
nand U2661 (N_2661,N_2589,N_2622);
or U2662 (N_2662,N_2594,N_2626);
nand U2663 (N_2663,N_2634,N_2627);
xnor U2664 (N_2664,N_2598,N_2639);
nand U2665 (N_2665,N_2623,N_2617);
and U2666 (N_2666,N_2592,N_2586);
nand U2667 (N_2667,N_2608,N_2616);
and U2668 (N_2668,N_2593,N_2618);
or U2669 (N_2669,N_2583,N_2630);
nor U2670 (N_2670,N_2580,N_2603);
nor U2671 (N_2671,N_2602,N_2638);
nand U2672 (N_2672,N_2592,N_2593);
nand U2673 (N_2673,N_2605,N_2620);
and U2674 (N_2674,N_2636,N_2600);
and U2675 (N_2675,N_2630,N_2636);
and U2676 (N_2676,N_2607,N_2630);
xor U2677 (N_2677,N_2600,N_2617);
or U2678 (N_2678,N_2629,N_2621);
nor U2679 (N_2679,N_2634,N_2605);
nand U2680 (N_2680,N_2583,N_2633);
nor U2681 (N_2681,N_2610,N_2604);
nand U2682 (N_2682,N_2609,N_2615);
nor U2683 (N_2683,N_2613,N_2637);
xnor U2684 (N_2684,N_2600,N_2623);
and U2685 (N_2685,N_2619,N_2632);
or U2686 (N_2686,N_2626,N_2611);
or U2687 (N_2687,N_2618,N_2625);
and U2688 (N_2688,N_2594,N_2580);
nand U2689 (N_2689,N_2619,N_2600);
nand U2690 (N_2690,N_2632,N_2587);
or U2691 (N_2691,N_2617,N_2605);
or U2692 (N_2692,N_2619,N_2605);
nand U2693 (N_2693,N_2612,N_2630);
nand U2694 (N_2694,N_2580,N_2605);
xnor U2695 (N_2695,N_2614,N_2616);
or U2696 (N_2696,N_2623,N_2637);
or U2697 (N_2697,N_2603,N_2625);
nand U2698 (N_2698,N_2639,N_2597);
nor U2699 (N_2699,N_2620,N_2631);
and U2700 (N_2700,N_2642,N_2641);
or U2701 (N_2701,N_2659,N_2675);
or U2702 (N_2702,N_2640,N_2688);
or U2703 (N_2703,N_2644,N_2686);
nor U2704 (N_2704,N_2672,N_2662);
and U2705 (N_2705,N_2690,N_2683);
or U2706 (N_2706,N_2648,N_2696);
or U2707 (N_2707,N_2656,N_2668);
nand U2708 (N_2708,N_2653,N_2670);
or U2709 (N_2709,N_2657,N_2694);
nand U2710 (N_2710,N_2666,N_2681);
nand U2711 (N_2711,N_2677,N_2698);
nand U2712 (N_2712,N_2643,N_2658);
nand U2713 (N_2713,N_2678,N_2660);
xnor U2714 (N_2714,N_2647,N_2693);
or U2715 (N_2715,N_2649,N_2682);
nand U2716 (N_2716,N_2667,N_2671);
nor U2717 (N_2717,N_2679,N_2655);
nand U2718 (N_2718,N_2699,N_2663);
and U2719 (N_2719,N_2680,N_2691);
and U2720 (N_2720,N_2692,N_2651);
or U2721 (N_2721,N_2669,N_2695);
or U2722 (N_2722,N_2650,N_2685);
or U2723 (N_2723,N_2645,N_2673);
and U2724 (N_2724,N_2652,N_2674);
nand U2725 (N_2725,N_2661,N_2676);
or U2726 (N_2726,N_2664,N_2646);
or U2727 (N_2727,N_2689,N_2697);
nor U2728 (N_2728,N_2687,N_2684);
nor U2729 (N_2729,N_2665,N_2654);
nor U2730 (N_2730,N_2652,N_2669);
and U2731 (N_2731,N_2686,N_2699);
or U2732 (N_2732,N_2681,N_2687);
nand U2733 (N_2733,N_2659,N_2646);
xor U2734 (N_2734,N_2648,N_2689);
nor U2735 (N_2735,N_2667,N_2643);
xor U2736 (N_2736,N_2664,N_2694);
and U2737 (N_2737,N_2647,N_2671);
or U2738 (N_2738,N_2693,N_2685);
nand U2739 (N_2739,N_2694,N_2692);
nor U2740 (N_2740,N_2663,N_2652);
nor U2741 (N_2741,N_2663,N_2667);
and U2742 (N_2742,N_2658,N_2697);
nor U2743 (N_2743,N_2678,N_2687);
or U2744 (N_2744,N_2663,N_2666);
nor U2745 (N_2745,N_2640,N_2646);
or U2746 (N_2746,N_2660,N_2659);
or U2747 (N_2747,N_2684,N_2680);
nor U2748 (N_2748,N_2648,N_2656);
nand U2749 (N_2749,N_2668,N_2649);
and U2750 (N_2750,N_2692,N_2697);
nand U2751 (N_2751,N_2653,N_2645);
nand U2752 (N_2752,N_2662,N_2679);
xor U2753 (N_2753,N_2699,N_2696);
nand U2754 (N_2754,N_2694,N_2674);
and U2755 (N_2755,N_2643,N_2647);
nand U2756 (N_2756,N_2690,N_2665);
and U2757 (N_2757,N_2688,N_2690);
and U2758 (N_2758,N_2699,N_2641);
or U2759 (N_2759,N_2641,N_2689);
or U2760 (N_2760,N_2732,N_2740);
or U2761 (N_2761,N_2726,N_2738);
xnor U2762 (N_2762,N_2720,N_2723);
nor U2763 (N_2763,N_2736,N_2753);
and U2764 (N_2764,N_2755,N_2728);
xnor U2765 (N_2765,N_2722,N_2757);
nor U2766 (N_2766,N_2704,N_2701);
nand U2767 (N_2767,N_2705,N_2747);
and U2768 (N_2768,N_2725,N_2733);
or U2769 (N_2769,N_2729,N_2737);
nand U2770 (N_2770,N_2713,N_2739);
nor U2771 (N_2771,N_2719,N_2724);
xor U2772 (N_2772,N_2706,N_2751);
and U2773 (N_2773,N_2748,N_2711);
nand U2774 (N_2774,N_2749,N_2743);
and U2775 (N_2775,N_2718,N_2721);
and U2776 (N_2776,N_2709,N_2744);
or U2777 (N_2777,N_2750,N_2715);
nor U2778 (N_2778,N_2700,N_2730);
or U2779 (N_2779,N_2714,N_2703);
or U2780 (N_2780,N_2734,N_2717);
or U2781 (N_2781,N_2716,N_2746);
nor U2782 (N_2782,N_2708,N_2710);
or U2783 (N_2783,N_2742,N_2735);
or U2784 (N_2784,N_2707,N_2702);
nor U2785 (N_2785,N_2759,N_2745);
nand U2786 (N_2786,N_2752,N_2727);
and U2787 (N_2787,N_2754,N_2712);
xnor U2788 (N_2788,N_2741,N_2731);
and U2789 (N_2789,N_2758,N_2756);
nor U2790 (N_2790,N_2735,N_2723);
nand U2791 (N_2791,N_2714,N_2730);
nand U2792 (N_2792,N_2735,N_2751);
or U2793 (N_2793,N_2753,N_2751);
xnor U2794 (N_2794,N_2714,N_2726);
or U2795 (N_2795,N_2727,N_2700);
xnor U2796 (N_2796,N_2735,N_2713);
or U2797 (N_2797,N_2734,N_2704);
or U2798 (N_2798,N_2743,N_2722);
nand U2799 (N_2799,N_2747,N_2759);
nand U2800 (N_2800,N_2722,N_2730);
and U2801 (N_2801,N_2743,N_2707);
and U2802 (N_2802,N_2710,N_2729);
nand U2803 (N_2803,N_2758,N_2705);
nand U2804 (N_2804,N_2704,N_2709);
nand U2805 (N_2805,N_2728,N_2730);
or U2806 (N_2806,N_2739,N_2726);
nor U2807 (N_2807,N_2736,N_2752);
nand U2808 (N_2808,N_2701,N_2752);
nor U2809 (N_2809,N_2729,N_2705);
or U2810 (N_2810,N_2758,N_2738);
nand U2811 (N_2811,N_2747,N_2728);
nor U2812 (N_2812,N_2728,N_2750);
or U2813 (N_2813,N_2707,N_2710);
nor U2814 (N_2814,N_2747,N_2706);
nand U2815 (N_2815,N_2747,N_2746);
xnor U2816 (N_2816,N_2704,N_2731);
nor U2817 (N_2817,N_2703,N_2731);
and U2818 (N_2818,N_2700,N_2724);
xor U2819 (N_2819,N_2749,N_2710);
and U2820 (N_2820,N_2778,N_2808);
or U2821 (N_2821,N_2772,N_2801);
xor U2822 (N_2822,N_2783,N_2815);
or U2823 (N_2823,N_2760,N_2780);
or U2824 (N_2824,N_2777,N_2797);
and U2825 (N_2825,N_2793,N_2775);
nand U2826 (N_2826,N_2763,N_2802);
nor U2827 (N_2827,N_2794,N_2774);
or U2828 (N_2828,N_2773,N_2795);
and U2829 (N_2829,N_2799,N_2813);
or U2830 (N_2830,N_2761,N_2762);
and U2831 (N_2831,N_2769,N_2786);
or U2832 (N_2832,N_2807,N_2779);
and U2833 (N_2833,N_2781,N_2771);
nor U2834 (N_2834,N_2809,N_2804);
and U2835 (N_2835,N_2782,N_2791);
nor U2836 (N_2836,N_2819,N_2800);
nor U2837 (N_2837,N_2788,N_2798);
or U2838 (N_2838,N_2812,N_2810);
nor U2839 (N_2839,N_2768,N_2803);
and U2840 (N_2840,N_2785,N_2787);
nor U2841 (N_2841,N_2765,N_2770);
and U2842 (N_2842,N_2816,N_2776);
nand U2843 (N_2843,N_2818,N_2814);
nand U2844 (N_2844,N_2796,N_2790);
nor U2845 (N_2845,N_2806,N_2817);
nand U2846 (N_2846,N_2784,N_2764);
and U2847 (N_2847,N_2789,N_2766);
and U2848 (N_2848,N_2805,N_2792);
or U2849 (N_2849,N_2767,N_2811);
xnor U2850 (N_2850,N_2812,N_2785);
nor U2851 (N_2851,N_2805,N_2782);
nor U2852 (N_2852,N_2785,N_2794);
nand U2853 (N_2853,N_2785,N_2772);
nand U2854 (N_2854,N_2810,N_2781);
or U2855 (N_2855,N_2795,N_2777);
and U2856 (N_2856,N_2802,N_2796);
nand U2857 (N_2857,N_2800,N_2775);
nor U2858 (N_2858,N_2768,N_2804);
and U2859 (N_2859,N_2798,N_2773);
xnor U2860 (N_2860,N_2785,N_2803);
or U2861 (N_2861,N_2809,N_2802);
nand U2862 (N_2862,N_2813,N_2819);
nand U2863 (N_2863,N_2773,N_2791);
or U2864 (N_2864,N_2765,N_2812);
nor U2865 (N_2865,N_2818,N_2805);
or U2866 (N_2866,N_2765,N_2817);
nand U2867 (N_2867,N_2761,N_2768);
nand U2868 (N_2868,N_2771,N_2810);
nand U2869 (N_2869,N_2790,N_2769);
or U2870 (N_2870,N_2777,N_2801);
xnor U2871 (N_2871,N_2808,N_2814);
xor U2872 (N_2872,N_2816,N_2763);
or U2873 (N_2873,N_2788,N_2767);
or U2874 (N_2874,N_2812,N_2818);
and U2875 (N_2875,N_2768,N_2777);
and U2876 (N_2876,N_2806,N_2819);
and U2877 (N_2877,N_2792,N_2815);
and U2878 (N_2878,N_2764,N_2769);
or U2879 (N_2879,N_2787,N_2770);
nand U2880 (N_2880,N_2875,N_2833);
nand U2881 (N_2881,N_2867,N_2878);
or U2882 (N_2882,N_2835,N_2841);
or U2883 (N_2883,N_2821,N_2823);
nor U2884 (N_2884,N_2843,N_2859);
or U2885 (N_2885,N_2857,N_2861);
and U2886 (N_2886,N_2824,N_2837);
nor U2887 (N_2887,N_2863,N_2864);
and U2888 (N_2888,N_2851,N_2871);
and U2889 (N_2889,N_2842,N_2827);
and U2890 (N_2890,N_2850,N_2872);
and U2891 (N_2891,N_2825,N_2854);
and U2892 (N_2892,N_2868,N_2862);
nor U2893 (N_2893,N_2829,N_2874);
and U2894 (N_2894,N_2847,N_2838);
or U2895 (N_2895,N_2845,N_2856);
nand U2896 (N_2896,N_2866,N_2852);
nor U2897 (N_2897,N_2826,N_2848);
or U2898 (N_2898,N_2849,N_2865);
and U2899 (N_2899,N_2879,N_2832);
or U2900 (N_2900,N_2840,N_2869);
nor U2901 (N_2901,N_2828,N_2858);
nor U2902 (N_2902,N_2822,N_2876);
or U2903 (N_2903,N_2831,N_2860);
xnor U2904 (N_2904,N_2853,N_2844);
nand U2905 (N_2905,N_2820,N_2834);
xnor U2906 (N_2906,N_2855,N_2873);
nand U2907 (N_2907,N_2846,N_2870);
nand U2908 (N_2908,N_2839,N_2836);
nor U2909 (N_2909,N_2830,N_2877);
nor U2910 (N_2910,N_2877,N_2838);
nor U2911 (N_2911,N_2870,N_2841);
nor U2912 (N_2912,N_2858,N_2830);
or U2913 (N_2913,N_2871,N_2843);
and U2914 (N_2914,N_2822,N_2871);
nand U2915 (N_2915,N_2844,N_2824);
or U2916 (N_2916,N_2829,N_2820);
nor U2917 (N_2917,N_2860,N_2849);
nor U2918 (N_2918,N_2844,N_2855);
or U2919 (N_2919,N_2844,N_2847);
nand U2920 (N_2920,N_2874,N_2849);
and U2921 (N_2921,N_2845,N_2850);
nand U2922 (N_2922,N_2878,N_2825);
or U2923 (N_2923,N_2840,N_2844);
or U2924 (N_2924,N_2844,N_2827);
nor U2925 (N_2925,N_2838,N_2848);
or U2926 (N_2926,N_2854,N_2842);
xor U2927 (N_2927,N_2851,N_2859);
xnor U2928 (N_2928,N_2855,N_2863);
nand U2929 (N_2929,N_2833,N_2874);
and U2930 (N_2930,N_2831,N_2878);
xor U2931 (N_2931,N_2858,N_2863);
nor U2932 (N_2932,N_2823,N_2835);
xor U2933 (N_2933,N_2879,N_2842);
and U2934 (N_2934,N_2862,N_2821);
and U2935 (N_2935,N_2870,N_2871);
xor U2936 (N_2936,N_2847,N_2867);
and U2937 (N_2937,N_2872,N_2844);
xnor U2938 (N_2938,N_2843,N_2844);
nand U2939 (N_2939,N_2830,N_2853);
nor U2940 (N_2940,N_2912,N_2937);
or U2941 (N_2941,N_2927,N_2887);
or U2942 (N_2942,N_2931,N_2921);
and U2943 (N_2943,N_2900,N_2906);
and U2944 (N_2944,N_2885,N_2934);
nand U2945 (N_2945,N_2886,N_2903);
and U2946 (N_2946,N_2895,N_2939);
and U2947 (N_2947,N_2916,N_2896);
nand U2948 (N_2948,N_2929,N_2928);
nor U2949 (N_2949,N_2930,N_2926);
nand U2950 (N_2950,N_2892,N_2883);
or U2951 (N_2951,N_2922,N_2914);
and U2952 (N_2952,N_2938,N_2881);
nor U2953 (N_2953,N_2897,N_2899);
nor U2954 (N_2954,N_2891,N_2890);
nand U2955 (N_2955,N_2904,N_2907);
or U2956 (N_2956,N_2919,N_2902);
xor U2957 (N_2957,N_2888,N_2898);
or U2958 (N_2958,N_2918,N_2905);
and U2959 (N_2959,N_2933,N_2913);
or U2960 (N_2960,N_2932,N_2908);
nand U2961 (N_2961,N_2894,N_2911);
and U2962 (N_2962,N_2910,N_2915);
nor U2963 (N_2963,N_2935,N_2901);
nor U2964 (N_2964,N_2924,N_2917);
nor U2965 (N_2965,N_2889,N_2920);
or U2966 (N_2966,N_2884,N_2923);
nand U2967 (N_2967,N_2893,N_2882);
and U2968 (N_2968,N_2925,N_2909);
nand U2969 (N_2969,N_2936,N_2880);
and U2970 (N_2970,N_2932,N_2892);
and U2971 (N_2971,N_2909,N_2926);
nand U2972 (N_2972,N_2914,N_2929);
nand U2973 (N_2973,N_2906,N_2924);
or U2974 (N_2974,N_2924,N_2893);
nor U2975 (N_2975,N_2916,N_2928);
or U2976 (N_2976,N_2880,N_2935);
and U2977 (N_2977,N_2887,N_2888);
or U2978 (N_2978,N_2891,N_2913);
or U2979 (N_2979,N_2887,N_2926);
or U2980 (N_2980,N_2927,N_2904);
and U2981 (N_2981,N_2911,N_2885);
nand U2982 (N_2982,N_2927,N_2923);
or U2983 (N_2983,N_2898,N_2903);
or U2984 (N_2984,N_2908,N_2893);
or U2985 (N_2985,N_2909,N_2903);
or U2986 (N_2986,N_2917,N_2881);
nand U2987 (N_2987,N_2916,N_2908);
nor U2988 (N_2988,N_2900,N_2893);
nand U2989 (N_2989,N_2938,N_2927);
and U2990 (N_2990,N_2937,N_2909);
nand U2991 (N_2991,N_2929,N_2901);
and U2992 (N_2992,N_2889,N_2883);
nor U2993 (N_2993,N_2938,N_2898);
nand U2994 (N_2994,N_2917,N_2913);
or U2995 (N_2995,N_2907,N_2896);
nor U2996 (N_2996,N_2937,N_2895);
nor U2997 (N_2997,N_2912,N_2891);
nand U2998 (N_2998,N_2925,N_2889);
nand U2999 (N_2999,N_2885,N_2895);
nand UO_0 (O_0,N_2976,N_2966);
or UO_1 (O_1,N_2994,N_2995);
nand UO_2 (O_2,N_2959,N_2961);
or UO_3 (O_3,N_2958,N_2996);
nor UO_4 (O_4,N_2989,N_2974);
xor UO_5 (O_5,N_2949,N_2953);
nand UO_6 (O_6,N_2951,N_2978);
nor UO_7 (O_7,N_2946,N_2977);
nand UO_8 (O_8,N_2988,N_2947);
nor UO_9 (O_9,N_2954,N_2952);
or UO_10 (O_10,N_2971,N_2968);
nand UO_11 (O_11,N_2975,N_2943);
and UO_12 (O_12,N_2987,N_2973);
nor UO_13 (O_13,N_2967,N_2941);
and UO_14 (O_14,N_2948,N_2983);
nand UO_15 (O_15,N_2991,N_2970);
and UO_16 (O_16,N_2997,N_2998);
or UO_17 (O_17,N_2982,N_2985);
or UO_18 (O_18,N_2981,N_2986);
nand UO_19 (O_19,N_2950,N_2999);
nand UO_20 (O_20,N_2993,N_2964);
or UO_21 (O_21,N_2963,N_2992);
nand UO_22 (O_22,N_2965,N_2945);
and UO_23 (O_23,N_2957,N_2942);
nand UO_24 (O_24,N_2960,N_2944);
nand UO_25 (O_25,N_2984,N_2940);
or UO_26 (O_26,N_2972,N_2990);
xor UO_27 (O_27,N_2980,N_2956);
nand UO_28 (O_28,N_2969,N_2979);
nor UO_29 (O_29,N_2955,N_2962);
xnor UO_30 (O_30,N_2972,N_2944);
and UO_31 (O_31,N_2989,N_2953);
or UO_32 (O_32,N_2961,N_2998);
and UO_33 (O_33,N_2971,N_2945);
or UO_34 (O_34,N_2992,N_2983);
or UO_35 (O_35,N_2965,N_2953);
nand UO_36 (O_36,N_2952,N_2955);
nor UO_37 (O_37,N_2984,N_2942);
and UO_38 (O_38,N_2962,N_2970);
and UO_39 (O_39,N_2950,N_2986);
xor UO_40 (O_40,N_2997,N_2962);
and UO_41 (O_41,N_2977,N_2943);
or UO_42 (O_42,N_2966,N_2971);
nand UO_43 (O_43,N_2956,N_2997);
nor UO_44 (O_44,N_2980,N_2961);
or UO_45 (O_45,N_2956,N_2940);
nor UO_46 (O_46,N_2946,N_2991);
nand UO_47 (O_47,N_2966,N_2982);
and UO_48 (O_48,N_2951,N_2962);
nand UO_49 (O_49,N_2976,N_2953);
nand UO_50 (O_50,N_2990,N_2977);
nor UO_51 (O_51,N_2948,N_2960);
or UO_52 (O_52,N_2968,N_2977);
nor UO_53 (O_53,N_2986,N_2994);
nand UO_54 (O_54,N_2942,N_2977);
or UO_55 (O_55,N_2999,N_2967);
and UO_56 (O_56,N_2967,N_2965);
or UO_57 (O_57,N_2967,N_2988);
and UO_58 (O_58,N_2952,N_2940);
or UO_59 (O_59,N_2944,N_2957);
nand UO_60 (O_60,N_2977,N_2982);
or UO_61 (O_61,N_2958,N_2977);
nand UO_62 (O_62,N_2978,N_2998);
nor UO_63 (O_63,N_2992,N_2976);
or UO_64 (O_64,N_2977,N_2985);
xor UO_65 (O_65,N_2992,N_2949);
nor UO_66 (O_66,N_2972,N_2986);
xnor UO_67 (O_67,N_2989,N_2993);
or UO_68 (O_68,N_2943,N_2969);
and UO_69 (O_69,N_2944,N_2959);
or UO_70 (O_70,N_2976,N_2972);
xor UO_71 (O_71,N_2965,N_2981);
nor UO_72 (O_72,N_2955,N_2983);
and UO_73 (O_73,N_2973,N_2953);
or UO_74 (O_74,N_2957,N_2945);
nand UO_75 (O_75,N_2973,N_2996);
xor UO_76 (O_76,N_2964,N_2963);
nor UO_77 (O_77,N_2999,N_2951);
and UO_78 (O_78,N_2991,N_2996);
nand UO_79 (O_79,N_2951,N_2994);
and UO_80 (O_80,N_2972,N_2942);
and UO_81 (O_81,N_2948,N_2973);
nand UO_82 (O_82,N_2986,N_2998);
or UO_83 (O_83,N_2960,N_2982);
and UO_84 (O_84,N_2941,N_2947);
nand UO_85 (O_85,N_2942,N_2973);
nand UO_86 (O_86,N_2994,N_2985);
and UO_87 (O_87,N_2980,N_2944);
and UO_88 (O_88,N_2969,N_2955);
xnor UO_89 (O_89,N_2997,N_2969);
nor UO_90 (O_90,N_2986,N_2955);
and UO_91 (O_91,N_2945,N_2969);
and UO_92 (O_92,N_2963,N_2966);
and UO_93 (O_93,N_2962,N_2980);
nor UO_94 (O_94,N_2954,N_2947);
and UO_95 (O_95,N_2948,N_2996);
xor UO_96 (O_96,N_2975,N_2970);
and UO_97 (O_97,N_2945,N_2958);
or UO_98 (O_98,N_2962,N_2942);
and UO_99 (O_99,N_2991,N_2976);
nor UO_100 (O_100,N_2954,N_2943);
or UO_101 (O_101,N_2983,N_2997);
nor UO_102 (O_102,N_2983,N_2964);
or UO_103 (O_103,N_2957,N_2956);
and UO_104 (O_104,N_2946,N_2998);
nand UO_105 (O_105,N_2959,N_2965);
and UO_106 (O_106,N_2949,N_2940);
nor UO_107 (O_107,N_2994,N_2973);
nand UO_108 (O_108,N_2961,N_2957);
and UO_109 (O_109,N_2977,N_2983);
nand UO_110 (O_110,N_2995,N_2971);
and UO_111 (O_111,N_2948,N_2944);
or UO_112 (O_112,N_2980,N_2999);
or UO_113 (O_113,N_2949,N_2959);
nor UO_114 (O_114,N_2953,N_2992);
nand UO_115 (O_115,N_2940,N_2990);
nand UO_116 (O_116,N_2981,N_2974);
and UO_117 (O_117,N_2983,N_2940);
nor UO_118 (O_118,N_2944,N_2996);
nor UO_119 (O_119,N_2954,N_2983);
or UO_120 (O_120,N_2990,N_2997);
nor UO_121 (O_121,N_2942,N_2943);
nor UO_122 (O_122,N_2985,N_2949);
or UO_123 (O_123,N_2997,N_2980);
xnor UO_124 (O_124,N_2980,N_2978);
or UO_125 (O_125,N_2964,N_2981);
nor UO_126 (O_126,N_2995,N_2984);
nand UO_127 (O_127,N_2971,N_2988);
nand UO_128 (O_128,N_2961,N_2969);
nand UO_129 (O_129,N_2944,N_2999);
or UO_130 (O_130,N_2944,N_2991);
xnor UO_131 (O_131,N_2983,N_2979);
nor UO_132 (O_132,N_2982,N_2955);
xor UO_133 (O_133,N_2945,N_2981);
and UO_134 (O_134,N_2973,N_2983);
and UO_135 (O_135,N_2950,N_2994);
and UO_136 (O_136,N_2999,N_2954);
or UO_137 (O_137,N_2978,N_2967);
and UO_138 (O_138,N_2999,N_2948);
or UO_139 (O_139,N_2945,N_2961);
and UO_140 (O_140,N_2980,N_2992);
xor UO_141 (O_141,N_2974,N_2959);
nand UO_142 (O_142,N_2955,N_2940);
xnor UO_143 (O_143,N_2961,N_2981);
nand UO_144 (O_144,N_2989,N_2943);
nor UO_145 (O_145,N_2958,N_2963);
nand UO_146 (O_146,N_2948,N_2982);
and UO_147 (O_147,N_2982,N_2967);
and UO_148 (O_148,N_2970,N_2993);
or UO_149 (O_149,N_2949,N_2986);
or UO_150 (O_150,N_2984,N_2948);
or UO_151 (O_151,N_2975,N_2977);
or UO_152 (O_152,N_2980,N_2943);
and UO_153 (O_153,N_2997,N_2942);
xor UO_154 (O_154,N_2994,N_2976);
nor UO_155 (O_155,N_2962,N_2993);
xor UO_156 (O_156,N_2977,N_2980);
nand UO_157 (O_157,N_2997,N_2941);
and UO_158 (O_158,N_2952,N_2977);
or UO_159 (O_159,N_2945,N_2992);
and UO_160 (O_160,N_2981,N_2962);
nand UO_161 (O_161,N_2990,N_2973);
or UO_162 (O_162,N_2998,N_2966);
nor UO_163 (O_163,N_2949,N_2950);
nand UO_164 (O_164,N_2949,N_2972);
or UO_165 (O_165,N_2970,N_2941);
and UO_166 (O_166,N_2956,N_2954);
or UO_167 (O_167,N_2957,N_2972);
nor UO_168 (O_168,N_2955,N_2951);
and UO_169 (O_169,N_2996,N_2943);
nor UO_170 (O_170,N_2961,N_2987);
nand UO_171 (O_171,N_2964,N_2966);
nand UO_172 (O_172,N_2981,N_2976);
nor UO_173 (O_173,N_2954,N_2988);
nand UO_174 (O_174,N_2972,N_2961);
and UO_175 (O_175,N_2963,N_2954);
or UO_176 (O_176,N_2949,N_2982);
nor UO_177 (O_177,N_2994,N_2998);
nand UO_178 (O_178,N_2948,N_2980);
nor UO_179 (O_179,N_2978,N_2966);
nor UO_180 (O_180,N_2959,N_2984);
nor UO_181 (O_181,N_2982,N_2996);
nand UO_182 (O_182,N_2968,N_2947);
or UO_183 (O_183,N_2984,N_2950);
and UO_184 (O_184,N_2977,N_2991);
nand UO_185 (O_185,N_2947,N_2964);
and UO_186 (O_186,N_2991,N_2982);
or UO_187 (O_187,N_2941,N_2944);
nor UO_188 (O_188,N_2975,N_2959);
xor UO_189 (O_189,N_2960,N_2945);
or UO_190 (O_190,N_2980,N_2975);
xor UO_191 (O_191,N_2971,N_2978);
nor UO_192 (O_192,N_2968,N_2984);
or UO_193 (O_193,N_2960,N_2951);
or UO_194 (O_194,N_2990,N_2992);
or UO_195 (O_195,N_2990,N_2994);
and UO_196 (O_196,N_2980,N_2940);
or UO_197 (O_197,N_2966,N_2999);
nor UO_198 (O_198,N_2946,N_2970);
xnor UO_199 (O_199,N_2977,N_2966);
nand UO_200 (O_200,N_2940,N_2947);
nor UO_201 (O_201,N_2985,N_2961);
and UO_202 (O_202,N_2997,N_2999);
or UO_203 (O_203,N_2974,N_2956);
nand UO_204 (O_204,N_2942,N_2985);
nand UO_205 (O_205,N_2990,N_2946);
and UO_206 (O_206,N_2952,N_2942);
and UO_207 (O_207,N_2989,N_2998);
or UO_208 (O_208,N_2974,N_2991);
or UO_209 (O_209,N_2970,N_2964);
nor UO_210 (O_210,N_2974,N_2963);
nor UO_211 (O_211,N_2985,N_2993);
nand UO_212 (O_212,N_2967,N_2975);
and UO_213 (O_213,N_2948,N_2997);
nor UO_214 (O_214,N_2973,N_2985);
nand UO_215 (O_215,N_2979,N_2996);
xnor UO_216 (O_216,N_2943,N_2978);
and UO_217 (O_217,N_2991,N_2972);
and UO_218 (O_218,N_2943,N_2974);
and UO_219 (O_219,N_2999,N_2975);
or UO_220 (O_220,N_2971,N_2941);
xnor UO_221 (O_221,N_2996,N_2980);
or UO_222 (O_222,N_2987,N_2993);
nand UO_223 (O_223,N_2961,N_2964);
or UO_224 (O_224,N_2975,N_2964);
nor UO_225 (O_225,N_2979,N_2980);
xor UO_226 (O_226,N_2973,N_2950);
nand UO_227 (O_227,N_2974,N_2995);
or UO_228 (O_228,N_2981,N_2979);
nand UO_229 (O_229,N_2959,N_2947);
or UO_230 (O_230,N_2949,N_2946);
and UO_231 (O_231,N_2994,N_2960);
and UO_232 (O_232,N_2995,N_2969);
nor UO_233 (O_233,N_2956,N_2975);
or UO_234 (O_234,N_2943,N_2960);
or UO_235 (O_235,N_2966,N_2955);
xnor UO_236 (O_236,N_2965,N_2941);
nor UO_237 (O_237,N_2946,N_2957);
xnor UO_238 (O_238,N_2943,N_2971);
or UO_239 (O_239,N_2991,N_2983);
nand UO_240 (O_240,N_2992,N_2973);
or UO_241 (O_241,N_2985,N_2941);
nand UO_242 (O_242,N_2943,N_2981);
or UO_243 (O_243,N_2942,N_2989);
and UO_244 (O_244,N_2971,N_2951);
or UO_245 (O_245,N_2998,N_2942);
nor UO_246 (O_246,N_2993,N_2982);
and UO_247 (O_247,N_2962,N_2972);
nor UO_248 (O_248,N_2991,N_2971);
nor UO_249 (O_249,N_2978,N_2957);
and UO_250 (O_250,N_2949,N_2943);
nor UO_251 (O_251,N_2941,N_2959);
and UO_252 (O_252,N_2983,N_2999);
and UO_253 (O_253,N_2954,N_2973);
xnor UO_254 (O_254,N_2954,N_2955);
nand UO_255 (O_255,N_2992,N_2971);
nand UO_256 (O_256,N_2982,N_2959);
xor UO_257 (O_257,N_2988,N_2966);
nor UO_258 (O_258,N_2998,N_2951);
and UO_259 (O_259,N_2970,N_2972);
nand UO_260 (O_260,N_2948,N_2989);
and UO_261 (O_261,N_2996,N_2983);
and UO_262 (O_262,N_2994,N_2981);
nor UO_263 (O_263,N_2985,N_2945);
and UO_264 (O_264,N_2987,N_2959);
nor UO_265 (O_265,N_2974,N_2973);
and UO_266 (O_266,N_2981,N_2954);
or UO_267 (O_267,N_2961,N_2948);
nand UO_268 (O_268,N_2957,N_2981);
or UO_269 (O_269,N_2951,N_2968);
nand UO_270 (O_270,N_2980,N_2988);
nor UO_271 (O_271,N_2965,N_2996);
nor UO_272 (O_272,N_2965,N_2991);
nand UO_273 (O_273,N_2960,N_2946);
nor UO_274 (O_274,N_2965,N_2960);
nor UO_275 (O_275,N_2963,N_2986);
and UO_276 (O_276,N_2968,N_2979);
nor UO_277 (O_277,N_2984,N_2965);
or UO_278 (O_278,N_2944,N_2986);
nor UO_279 (O_279,N_2960,N_2976);
or UO_280 (O_280,N_2942,N_2953);
or UO_281 (O_281,N_2940,N_2946);
nand UO_282 (O_282,N_2966,N_2944);
and UO_283 (O_283,N_2944,N_2997);
nand UO_284 (O_284,N_2956,N_2984);
and UO_285 (O_285,N_2961,N_2982);
or UO_286 (O_286,N_2963,N_2988);
and UO_287 (O_287,N_2988,N_2975);
or UO_288 (O_288,N_2952,N_2979);
nor UO_289 (O_289,N_2951,N_2964);
nor UO_290 (O_290,N_2998,N_2960);
or UO_291 (O_291,N_2964,N_2944);
and UO_292 (O_292,N_2996,N_2972);
nand UO_293 (O_293,N_2943,N_2963);
xnor UO_294 (O_294,N_2979,N_2985);
or UO_295 (O_295,N_2972,N_2974);
nor UO_296 (O_296,N_2973,N_2976);
xor UO_297 (O_297,N_2970,N_2976);
nor UO_298 (O_298,N_2962,N_2961);
or UO_299 (O_299,N_2949,N_2984);
nor UO_300 (O_300,N_2987,N_2976);
xnor UO_301 (O_301,N_2977,N_2988);
nand UO_302 (O_302,N_2982,N_2994);
nor UO_303 (O_303,N_2971,N_2970);
nand UO_304 (O_304,N_2990,N_2948);
nand UO_305 (O_305,N_2954,N_2995);
or UO_306 (O_306,N_2943,N_2993);
and UO_307 (O_307,N_2957,N_2974);
or UO_308 (O_308,N_2995,N_2987);
or UO_309 (O_309,N_2983,N_2974);
or UO_310 (O_310,N_2978,N_2954);
nand UO_311 (O_311,N_2954,N_2951);
nor UO_312 (O_312,N_2980,N_2968);
nand UO_313 (O_313,N_2984,N_2953);
nand UO_314 (O_314,N_2969,N_2964);
nand UO_315 (O_315,N_2952,N_2999);
or UO_316 (O_316,N_2993,N_2963);
xor UO_317 (O_317,N_2961,N_2994);
nand UO_318 (O_318,N_2947,N_2944);
nand UO_319 (O_319,N_2991,N_2953);
or UO_320 (O_320,N_2941,N_2981);
and UO_321 (O_321,N_2960,N_2940);
xnor UO_322 (O_322,N_2975,N_2973);
and UO_323 (O_323,N_2987,N_2945);
nor UO_324 (O_324,N_2985,N_2946);
and UO_325 (O_325,N_2994,N_2974);
and UO_326 (O_326,N_2990,N_2986);
nand UO_327 (O_327,N_2982,N_2990);
nand UO_328 (O_328,N_2966,N_2957);
or UO_329 (O_329,N_2994,N_2968);
nand UO_330 (O_330,N_2940,N_2976);
and UO_331 (O_331,N_2958,N_2992);
nand UO_332 (O_332,N_2986,N_2940);
or UO_333 (O_333,N_2974,N_2990);
or UO_334 (O_334,N_2944,N_2956);
nand UO_335 (O_335,N_2960,N_2956);
or UO_336 (O_336,N_2943,N_2992);
or UO_337 (O_337,N_2975,N_2965);
nor UO_338 (O_338,N_2946,N_2961);
and UO_339 (O_339,N_2996,N_2946);
or UO_340 (O_340,N_2956,N_2983);
or UO_341 (O_341,N_2997,N_2995);
or UO_342 (O_342,N_2962,N_2966);
nand UO_343 (O_343,N_2966,N_2983);
or UO_344 (O_344,N_2963,N_2952);
nor UO_345 (O_345,N_2968,N_2983);
and UO_346 (O_346,N_2993,N_2959);
nand UO_347 (O_347,N_2967,N_2948);
xnor UO_348 (O_348,N_2978,N_2946);
or UO_349 (O_349,N_2967,N_2993);
and UO_350 (O_350,N_2989,N_2940);
xnor UO_351 (O_351,N_2990,N_2981);
nand UO_352 (O_352,N_2941,N_2966);
nand UO_353 (O_353,N_2978,N_2975);
and UO_354 (O_354,N_2940,N_2957);
nor UO_355 (O_355,N_2947,N_2989);
and UO_356 (O_356,N_2987,N_2985);
and UO_357 (O_357,N_2994,N_2943);
or UO_358 (O_358,N_2957,N_2955);
or UO_359 (O_359,N_2990,N_2953);
xor UO_360 (O_360,N_2951,N_2989);
xor UO_361 (O_361,N_2969,N_2948);
or UO_362 (O_362,N_2987,N_2970);
nor UO_363 (O_363,N_2954,N_2969);
nor UO_364 (O_364,N_2956,N_2989);
nand UO_365 (O_365,N_2992,N_2968);
nand UO_366 (O_366,N_2950,N_2975);
xnor UO_367 (O_367,N_2951,N_2945);
or UO_368 (O_368,N_2940,N_2996);
nand UO_369 (O_369,N_2945,N_2988);
or UO_370 (O_370,N_2954,N_2960);
and UO_371 (O_371,N_2987,N_2942);
nand UO_372 (O_372,N_2983,N_2946);
and UO_373 (O_373,N_2993,N_2956);
and UO_374 (O_374,N_2963,N_2975);
and UO_375 (O_375,N_2942,N_2982);
and UO_376 (O_376,N_2961,N_2971);
xnor UO_377 (O_377,N_2998,N_2953);
and UO_378 (O_378,N_2979,N_2974);
or UO_379 (O_379,N_2987,N_2988);
nor UO_380 (O_380,N_2951,N_2950);
nor UO_381 (O_381,N_2983,N_2962);
or UO_382 (O_382,N_2962,N_2982);
and UO_383 (O_383,N_2942,N_2950);
nor UO_384 (O_384,N_2982,N_2979);
nor UO_385 (O_385,N_2991,N_2978);
nor UO_386 (O_386,N_2974,N_2977);
and UO_387 (O_387,N_2999,N_2961);
nor UO_388 (O_388,N_2961,N_2995);
nand UO_389 (O_389,N_2992,N_2960);
and UO_390 (O_390,N_2954,N_2977);
nor UO_391 (O_391,N_2972,N_2948);
nor UO_392 (O_392,N_2950,N_2969);
and UO_393 (O_393,N_2950,N_2960);
or UO_394 (O_394,N_2977,N_2950);
nor UO_395 (O_395,N_2965,N_2964);
and UO_396 (O_396,N_2962,N_2988);
and UO_397 (O_397,N_2942,N_2956);
nand UO_398 (O_398,N_2978,N_2973);
xor UO_399 (O_399,N_2977,N_2970);
or UO_400 (O_400,N_2991,N_2943);
nand UO_401 (O_401,N_2965,N_2993);
and UO_402 (O_402,N_2968,N_2945);
nand UO_403 (O_403,N_2981,N_2969);
or UO_404 (O_404,N_2946,N_2945);
or UO_405 (O_405,N_2971,N_2975);
or UO_406 (O_406,N_2956,N_2995);
or UO_407 (O_407,N_2941,N_2987);
xor UO_408 (O_408,N_2977,N_2996);
nand UO_409 (O_409,N_2956,N_2973);
nand UO_410 (O_410,N_2988,N_2949);
nand UO_411 (O_411,N_2965,N_2962);
and UO_412 (O_412,N_2999,N_2962);
xnor UO_413 (O_413,N_2976,N_2971);
nor UO_414 (O_414,N_2982,N_2970);
xnor UO_415 (O_415,N_2976,N_2967);
and UO_416 (O_416,N_2972,N_2947);
nand UO_417 (O_417,N_2945,N_2948);
and UO_418 (O_418,N_2966,N_2987);
or UO_419 (O_419,N_2988,N_2996);
nor UO_420 (O_420,N_2984,N_2955);
nand UO_421 (O_421,N_2969,N_2965);
nand UO_422 (O_422,N_2969,N_2949);
nand UO_423 (O_423,N_2988,N_2982);
or UO_424 (O_424,N_2942,N_2986);
and UO_425 (O_425,N_2965,N_2961);
or UO_426 (O_426,N_2962,N_2946);
or UO_427 (O_427,N_2965,N_2998);
xor UO_428 (O_428,N_2947,N_2979);
nor UO_429 (O_429,N_2992,N_2952);
and UO_430 (O_430,N_2980,N_2998);
nor UO_431 (O_431,N_2988,N_2978);
or UO_432 (O_432,N_2979,N_2967);
xor UO_433 (O_433,N_2982,N_2972);
nor UO_434 (O_434,N_2961,N_2986);
nor UO_435 (O_435,N_2997,N_2979);
xor UO_436 (O_436,N_2951,N_2957);
nor UO_437 (O_437,N_2988,N_2957);
and UO_438 (O_438,N_2971,N_2994);
or UO_439 (O_439,N_2979,N_2948);
or UO_440 (O_440,N_2970,N_2960);
and UO_441 (O_441,N_2944,N_2990);
xnor UO_442 (O_442,N_2977,N_2960);
and UO_443 (O_443,N_2974,N_2985);
nand UO_444 (O_444,N_2970,N_2949);
nor UO_445 (O_445,N_2955,N_2999);
or UO_446 (O_446,N_2963,N_2981);
nor UO_447 (O_447,N_2999,N_2968);
nor UO_448 (O_448,N_2967,N_2971);
nor UO_449 (O_449,N_2958,N_2989);
nor UO_450 (O_450,N_2991,N_2973);
nor UO_451 (O_451,N_2947,N_2955);
nand UO_452 (O_452,N_2964,N_2992);
or UO_453 (O_453,N_2967,N_2945);
nand UO_454 (O_454,N_2949,N_2956);
nand UO_455 (O_455,N_2988,N_2961);
xor UO_456 (O_456,N_2995,N_2953);
nor UO_457 (O_457,N_2967,N_2974);
and UO_458 (O_458,N_2970,N_2992);
and UO_459 (O_459,N_2940,N_2994);
and UO_460 (O_460,N_2998,N_2988);
nand UO_461 (O_461,N_2999,N_2956);
nor UO_462 (O_462,N_2968,N_2956);
nor UO_463 (O_463,N_2979,N_2971);
or UO_464 (O_464,N_2961,N_2974);
or UO_465 (O_465,N_2984,N_2997);
nor UO_466 (O_466,N_2956,N_2994);
and UO_467 (O_467,N_2961,N_2989);
nand UO_468 (O_468,N_2950,N_2966);
nor UO_469 (O_469,N_2976,N_2998);
nor UO_470 (O_470,N_2943,N_2958);
nand UO_471 (O_471,N_2953,N_2969);
and UO_472 (O_472,N_2958,N_2966);
nand UO_473 (O_473,N_2964,N_2999);
and UO_474 (O_474,N_2950,N_2989);
nor UO_475 (O_475,N_2949,N_2998);
or UO_476 (O_476,N_2958,N_2982);
and UO_477 (O_477,N_2948,N_2959);
and UO_478 (O_478,N_2955,N_2998);
or UO_479 (O_479,N_2961,N_2990);
nor UO_480 (O_480,N_2961,N_2954);
or UO_481 (O_481,N_2969,N_2974);
and UO_482 (O_482,N_2959,N_2971);
and UO_483 (O_483,N_2988,N_2976);
nor UO_484 (O_484,N_2990,N_2985);
nor UO_485 (O_485,N_2990,N_2966);
or UO_486 (O_486,N_2998,N_2975);
nor UO_487 (O_487,N_2949,N_2971);
nor UO_488 (O_488,N_2974,N_2948);
or UO_489 (O_489,N_2944,N_2982);
nand UO_490 (O_490,N_2969,N_2947);
or UO_491 (O_491,N_2959,N_2951);
nand UO_492 (O_492,N_2989,N_2955);
nand UO_493 (O_493,N_2943,N_2983);
nor UO_494 (O_494,N_2996,N_2959);
nor UO_495 (O_495,N_2981,N_2982);
nand UO_496 (O_496,N_2988,N_2960);
nor UO_497 (O_497,N_2952,N_2993);
or UO_498 (O_498,N_2947,N_2974);
nor UO_499 (O_499,N_2964,N_2987);
endmodule