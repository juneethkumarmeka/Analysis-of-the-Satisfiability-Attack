module basic_500_3000_500_60_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_336,In_97);
and U1 (N_1,In_465,In_257);
or U2 (N_2,In_18,In_246);
nand U3 (N_3,In_149,In_395);
and U4 (N_4,In_310,In_84);
or U5 (N_5,In_114,In_202);
nand U6 (N_6,In_16,In_463);
nand U7 (N_7,In_230,In_394);
nand U8 (N_8,In_214,In_220);
and U9 (N_9,In_113,In_19);
or U10 (N_10,In_91,In_212);
nand U11 (N_11,In_377,In_355);
or U12 (N_12,In_101,In_450);
and U13 (N_13,In_140,In_129);
or U14 (N_14,In_262,In_15);
nand U15 (N_15,In_49,In_311);
nand U16 (N_16,In_444,In_486);
and U17 (N_17,In_156,In_415);
and U18 (N_18,In_418,In_61);
nand U19 (N_19,In_436,In_164);
or U20 (N_20,In_191,In_72);
nand U21 (N_21,In_335,In_48);
or U22 (N_22,In_75,In_357);
nor U23 (N_23,In_85,In_272);
nor U24 (N_24,In_458,In_152);
or U25 (N_25,In_44,In_5);
and U26 (N_26,In_365,In_118);
nand U27 (N_27,In_494,In_0);
nand U28 (N_28,In_263,In_204);
nand U29 (N_29,In_349,In_95);
or U30 (N_30,In_8,In_332);
and U31 (N_31,In_322,In_136);
nor U32 (N_32,In_51,In_177);
nand U33 (N_33,In_242,In_386);
and U34 (N_34,In_217,In_475);
nand U35 (N_35,In_182,In_40);
nand U36 (N_36,In_430,In_338);
nor U37 (N_37,In_170,In_356);
or U38 (N_38,In_438,In_34);
xnor U39 (N_39,In_427,In_209);
or U40 (N_40,In_329,In_150);
or U41 (N_41,In_396,In_65);
nor U42 (N_42,In_260,In_341);
or U43 (N_43,In_304,In_483);
nand U44 (N_44,In_478,In_171);
xnor U45 (N_45,In_408,In_172);
or U46 (N_46,In_31,In_146);
nor U47 (N_47,In_142,In_23);
nand U48 (N_48,In_71,In_208);
nor U49 (N_49,In_412,In_120);
and U50 (N_50,In_218,N_42);
nand U51 (N_51,In_42,In_62);
or U52 (N_52,In_441,In_487);
nor U53 (N_53,N_4,N_41);
nand U54 (N_54,In_434,In_312);
and U55 (N_55,In_473,In_24);
nand U56 (N_56,In_378,In_155);
nor U57 (N_57,In_265,In_213);
and U58 (N_58,N_31,In_173);
nor U59 (N_59,N_10,In_169);
xnor U60 (N_60,In_374,In_20);
xnor U61 (N_61,In_184,In_132);
or U62 (N_62,N_29,In_210);
nand U63 (N_63,In_145,In_227);
nand U64 (N_64,In_433,In_47);
nand U65 (N_65,In_89,In_411);
or U66 (N_66,In_404,N_25);
nor U67 (N_67,In_4,In_92);
nor U68 (N_68,In_285,In_387);
nand U69 (N_69,In_66,N_46);
or U70 (N_70,In_470,In_327);
and U71 (N_71,In_313,In_30);
nor U72 (N_72,In_316,N_17);
or U73 (N_73,In_485,In_130);
nor U74 (N_74,In_471,In_122);
nand U75 (N_75,In_498,In_160);
and U76 (N_76,In_350,In_141);
nand U77 (N_77,In_426,In_307);
or U78 (N_78,In_368,In_10);
nand U79 (N_79,In_370,In_440);
nor U80 (N_80,In_296,In_109);
and U81 (N_81,In_73,In_369);
nand U82 (N_82,In_28,In_309);
or U83 (N_83,In_86,In_385);
nor U84 (N_84,In_39,In_479);
nand U85 (N_85,In_64,In_36);
nor U86 (N_86,N_38,In_253);
or U87 (N_87,In_446,In_12);
nand U88 (N_88,In_466,N_7);
xnor U89 (N_89,In_148,In_45);
nor U90 (N_90,In_139,In_106);
nor U91 (N_91,In_468,In_424);
xor U92 (N_92,In_105,In_244);
or U93 (N_93,N_33,N_44);
nor U94 (N_94,In_428,In_302);
or U95 (N_95,In_480,In_460);
or U96 (N_96,In_94,In_381);
nor U97 (N_97,In_207,In_358);
or U98 (N_98,In_27,N_35);
nand U99 (N_99,In_180,In_442);
xnor U100 (N_100,N_70,In_81);
or U101 (N_101,N_54,In_401);
or U102 (N_102,In_351,In_281);
nor U103 (N_103,In_174,In_299);
xnor U104 (N_104,In_420,In_491);
xor U105 (N_105,In_371,In_407);
and U106 (N_106,In_195,In_205);
nor U107 (N_107,In_168,In_294);
nand U108 (N_108,N_1,In_287);
or U109 (N_109,In_163,In_477);
or U110 (N_110,In_157,In_80);
nand U111 (N_111,In_111,In_280);
nor U112 (N_112,In_421,In_297);
or U113 (N_113,In_211,N_80);
nor U114 (N_114,N_96,In_413);
nor U115 (N_115,In_186,In_429);
nand U116 (N_116,In_423,In_151);
or U117 (N_117,N_95,In_288);
xor U118 (N_118,In_258,In_376);
or U119 (N_119,In_78,In_321);
nand U120 (N_120,N_57,In_324);
nand U121 (N_121,In_254,In_189);
or U122 (N_122,In_58,In_372);
or U123 (N_123,In_128,In_46);
nor U124 (N_124,In_448,In_289);
and U125 (N_125,N_55,In_226);
nor U126 (N_126,N_15,In_380);
or U127 (N_127,In_459,In_451);
and U128 (N_128,In_190,In_419);
nor U129 (N_129,In_241,In_279);
nor U130 (N_130,In_293,In_138);
nor U131 (N_131,In_476,In_41);
or U132 (N_132,In_422,In_306);
and U133 (N_133,In_482,In_431);
and U134 (N_134,In_320,In_445);
nor U135 (N_135,In_382,In_29);
nor U136 (N_136,In_390,In_499);
or U137 (N_137,In_99,N_26);
or U138 (N_138,In_2,In_250);
and U139 (N_139,In_67,In_154);
nand U140 (N_140,In_53,In_112);
nand U141 (N_141,In_266,In_222);
nor U142 (N_142,In_193,In_117);
or U143 (N_143,In_88,In_219);
nand U144 (N_144,N_98,In_247);
xor U145 (N_145,N_11,In_22);
or U146 (N_146,In_269,In_496);
nand U147 (N_147,N_92,In_277);
nand U148 (N_148,N_28,In_389);
xor U149 (N_149,N_30,N_83);
nor U150 (N_150,N_116,N_58);
or U151 (N_151,In_215,In_185);
xor U152 (N_152,In_410,In_308);
nor U153 (N_153,In_198,N_132);
or U154 (N_154,N_137,In_314);
nor U155 (N_155,In_437,In_38);
or U156 (N_156,N_88,In_249);
nor U157 (N_157,In_133,In_323);
nand U158 (N_158,N_19,In_236);
or U159 (N_159,N_133,N_45);
nand U160 (N_160,N_52,In_96);
or U161 (N_161,N_74,In_60);
or U162 (N_162,In_238,In_290);
xnor U163 (N_163,In_178,In_9);
and U164 (N_164,N_142,N_117);
xnor U165 (N_165,N_146,N_134);
or U166 (N_166,In_181,N_89);
nand U167 (N_167,N_147,In_397);
nand U168 (N_168,In_367,In_301);
nand U169 (N_169,In_197,N_21);
or U170 (N_170,In_384,In_143);
nand U171 (N_171,N_6,In_334);
nand U172 (N_172,In_98,In_409);
nand U173 (N_173,In_93,In_1);
xnor U174 (N_174,In_449,In_467);
nand U175 (N_175,In_119,In_282);
nand U176 (N_176,N_69,In_347);
nand U177 (N_177,N_13,In_158);
nand U178 (N_178,In_489,In_57);
or U179 (N_179,In_255,In_239);
xnor U180 (N_180,In_35,N_102);
and U181 (N_181,In_402,In_264);
nor U182 (N_182,In_11,N_101);
xor U183 (N_183,In_317,In_50);
nand U184 (N_184,N_90,In_417);
or U185 (N_185,In_267,N_62);
or U186 (N_186,N_20,In_276);
nand U187 (N_187,N_149,N_36);
nor U188 (N_188,In_360,N_139);
nand U189 (N_189,N_143,N_126);
or U190 (N_190,In_175,In_388);
and U191 (N_191,In_333,In_464);
and U192 (N_192,N_59,In_56);
nor U193 (N_193,N_127,In_79);
or U194 (N_194,In_32,N_68);
or U195 (N_195,N_85,N_12);
or U196 (N_196,In_90,In_278);
nand U197 (N_197,In_3,N_99);
and U198 (N_198,In_108,N_107);
or U199 (N_199,N_14,N_71);
or U200 (N_200,In_188,In_456);
xor U201 (N_201,N_154,N_135);
nor U202 (N_202,In_492,N_97);
nand U203 (N_203,In_472,In_74);
or U204 (N_204,N_27,N_186);
or U205 (N_205,N_179,N_199);
xnor U206 (N_206,N_118,In_147);
xnor U207 (N_207,N_136,In_361);
nor U208 (N_208,In_425,In_363);
nand U209 (N_209,N_24,N_173);
and U210 (N_210,N_86,N_108);
nand U211 (N_211,N_16,In_121);
and U212 (N_212,In_87,N_104);
or U213 (N_213,In_447,In_196);
and U214 (N_214,N_131,N_73);
and U215 (N_215,N_3,N_67);
nor U216 (N_216,N_171,In_252);
or U217 (N_217,N_188,In_59);
nor U218 (N_218,N_140,In_457);
nand U219 (N_219,In_286,In_194);
or U220 (N_220,In_391,In_201);
and U221 (N_221,N_100,In_76);
nor U222 (N_222,N_119,In_298);
nor U223 (N_223,N_77,In_179);
nand U224 (N_224,In_319,N_176);
and U225 (N_225,In_134,N_60);
xor U226 (N_226,N_115,In_439);
nand U227 (N_227,In_344,In_127);
nor U228 (N_228,N_32,N_56);
nor U229 (N_229,In_153,In_100);
or U230 (N_230,N_180,N_128);
or U231 (N_231,In_490,In_271);
or U232 (N_232,N_122,In_70);
nand U233 (N_233,N_111,In_229);
and U234 (N_234,In_162,In_137);
nor U235 (N_235,In_115,In_453);
and U236 (N_236,N_159,In_256);
nor U237 (N_237,N_114,In_455);
nor U238 (N_238,In_305,In_52);
nor U239 (N_239,N_125,In_176);
xor U240 (N_240,N_61,N_191);
or U241 (N_241,In_495,In_346);
nor U242 (N_242,N_2,N_184);
nand U243 (N_243,In_461,N_112);
xnor U244 (N_244,N_79,In_77);
and U245 (N_245,In_234,N_81);
and U246 (N_246,In_63,N_187);
nand U247 (N_247,N_103,In_37);
and U248 (N_248,N_39,N_198);
nand U249 (N_249,In_318,N_22);
nand U250 (N_250,N_47,N_144);
and U251 (N_251,In_343,N_123);
or U252 (N_252,In_144,N_206);
nand U253 (N_253,N_168,N_156);
and U254 (N_254,N_222,N_232);
and U255 (N_255,N_192,In_125);
nand U256 (N_256,N_201,N_43);
or U257 (N_257,N_214,In_224);
nor U258 (N_258,N_121,In_235);
and U259 (N_259,N_167,In_295);
and U260 (N_260,In_399,N_233);
and U261 (N_261,N_219,N_0);
and U262 (N_262,N_160,In_192);
nor U263 (N_263,N_158,N_174);
and U264 (N_264,In_400,In_107);
and U265 (N_265,N_82,N_150);
or U266 (N_266,In_126,N_65);
and U267 (N_267,N_212,N_76);
and U268 (N_268,In_379,In_452);
or U269 (N_269,N_157,N_249);
nand U270 (N_270,N_172,In_116);
and U271 (N_271,N_48,In_26);
nand U272 (N_272,In_291,In_359);
or U273 (N_273,N_197,N_246);
nor U274 (N_274,N_9,In_484);
nor U275 (N_275,In_21,In_221);
nor U276 (N_276,N_64,In_497);
or U277 (N_277,N_205,In_366);
nand U278 (N_278,In_166,N_189);
nand U279 (N_279,N_181,N_243);
xor U280 (N_280,N_215,In_82);
and U281 (N_281,N_130,N_213);
nand U282 (N_282,N_218,N_202);
and U283 (N_283,N_161,In_69);
nor U284 (N_284,N_109,In_104);
xnor U285 (N_285,In_303,N_164);
and U286 (N_286,N_242,N_53);
nor U287 (N_287,N_216,In_273);
nor U288 (N_288,N_34,N_138);
nor U289 (N_289,N_225,In_469);
nand U290 (N_290,N_182,In_414);
and U291 (N_291,N_145,N_245);
xor U292 (N_292,In_330,N_178);
or U293 (N_293,N_195,N_110);
and U294 (N_294,In_167,In_454);
and U295 (N_295,In_200,In_232);
and U296 (N_296,In_340,N_204);
nor U297 (N_297,In_352,In_223);
xnor U298 (N_298,In_432,N_223);
nor U299 (N_299,In_259,In_435);
xor U300 (N_300,N_170,N_23);
nor U301 (N_301,N_37,N_165);
xor U302 (N_302,N_129,In_6);
nor U303 (N_303,N_239,N_40);
nor U304 (N_304,In_131,N_63);
or U305 (N_305,In_345,In_348);
nor U306 (N_306,In_233,In_275);
nand U307 (N_307,In_54,N_237);
and U308 (N_308,N_105,N_280);
and U309 (N_309,N_238,N_166);
xnor U310 (N_310,N_235,In_102);
or U311 (N_311,N_155,N_279);
or U312 (N_312,N_203,In_123);
and U313 (N_313,In_199,N_281);
or U314 (N_314,N_262,In_161);
or U315 (N_315,In_362,N_271);
and U316 (N_316,N_257,In_268);
nor U317 (N_317,N_87,N_296);
or U318 (N_318,In_110,In_315);
nand U319 (N_319,N_220,In_326);
or U320 (N_320,N_175,N_261);
nor U321 (N_321,N_51,N_268);
and U322 (N_322,N_228,N_190);
or U323 (N_323,In_274,In_245);
or U324 (N_324,N_211,In_216);
or U325 (N_325,N_236,N_231);
nor U326 (N_326,N_113,In_231);
or U327 (N_327,N_124,N_94);
or U328 (N_328,N_278,In_398);
and U329 (N_329,In_13,N_292);
nand U330 (N_330,N_153,N_252);
nor U331 (N_331,In_474,N_208);
nand U332 (N_332,N_291,In_261);
nand U333 (N_333,N_224,N_287);
and U334 (N_334,N_260,N_8);
nor U335 (N_335,N_256,In_353);
and U336 (N_336,N_162,In_392);
or U337 (N_337,N_66,N_200);
nand U338 (N_338,N_194,In_25);
and U339 (N_339,N_244,In_124);
nand U340 (N_340,N_251,In_393);
nor U341 (N_341,In_183,In_481);
nand U342 (N_342,N_286,N_298);
nand U343 (N_343,In_292,In_55);
or U344 (N_344,N_248,In_243);
nor U345 (N_345,N_295,N_290);
or U346 (N_346,N_230,In_225);
and U347 (N_347,In_187,In_339);
and U348 (N_348,In_300,In_43);
nand U349 (N_349,In_203,N_283);
nand U350 (N_350,N_319,N_285);
xor U351 (N_351,N_310,N_265);
nand U352 (N_352,In_462,N_207);
and U353 (N_353,N_183,N_339);
nor U354 (N_354,In_493,N_333);
xor U355 (N_355,N_301,N_317);
nand U356 (N_356,In_159,N_169);
nor U357 (N_357,N_315,N_196);
and U358 (N_358,N_309,N_277);
nor U359 (N_359,N_330,N_331);
nand U360 (N_360,N_84,N_273);
nor U361 (N_361,N_141,N_163);
xnor U362 (N_362,N_328,N_151);
xor U363 (N_363,N_348,N_50);
xor U364 (N_364,In_443,N_253);
nor U365 (N_365,N_193,In_325);
nor U366 (N_366,N_318,N_272);
and U367 (N_367,N_259,N_346);
xor U368 (N_368,N_342,In_373);
nand U369 (N_369,N_241,N_324);
and U370 (N_370,In_240,N_276);
xnor U371 (N_371,In_403,N_314);
nand U372 (N_372,N_263,N_210);
or U373 (N_373,N_18,N_217);
and U374 (N_374,In_17,N_326);
and U375 (N_375,N_282,In_68);
and U376 (N_376,In_135,N_307);
and U377 (N_377,N_78,N_322);
xnor U378 (N_378,In_83,N_267);
or U379 (N_379,In_375,N_247);
or U380 (N_380,In_354,N_335);
and U381 (N_381,N_270,N_288);
nor U382 (N_382,In_488,N_349);
or U383 (N_383,N_226,In_251);
and U384 (N_384,N_294,N_341);
nor U385 (N_385,N_152,N_289);
or U386 (N_386,N_5,N_269);
or U387 (N_387,N_240,N_254);
and U388 (N_388,In_416,N_308);
nor U389 (N_389,In_228,N_327);
nor U390 (N_390,In_405,N_302);
nor U391 (N_391,In_331,In_165);
xnor U392 (N_392,N_325,N_320);
and U393 (N_393,N_227,N_340);
or U394 (N_394,In_284,N_229);
nor U395 (N_395,N_250,In_337);
nand U396 (N_396,N_72,N_293);
and U397 (N_397,In_33,In_270);
nand U398 (N_398,N_148,N_323);
nor U399 (N_399,N_305,N_332);
and U400 (N_400,N_388,N_177);
and U401 (N_401,In_383,N_360);
nor U402 (N_402,In_328,N_364);
nand U403 (N_403,N_372,N_363);
nand U404 (N_404,N_356,N_395);
xnor U405 (N_405,N_106,In_248);
and U406 (N_406,N_338,N_329);
and U407 (N_407,N_397,N_382);
or U408 (N_408,N_300,N_361);
and U409 (N_409,N_367,N_384);
nand U410 (N_410,N_390,N_377);
and U411 (N_411,N_368,N_347);
nor U412 (N_412,N_396,N_185);
nand U413 (N_413,N_389,N_264);
or U414 (N_414,N_120,N_355);
nand U415 (N_415,N_378,N_334);
nor U416 (N_416,N_297,N_303);
and U417 (N_417,N_391,N_91);
nand U418 (N_418,In_406,N_383);
nor U419 (N_419,N_221,N_337);
nand U420 (N_420,N_312,N_234);
and U421 (N_421,N_387,N_375);
or U422 (N_422,N_93,N_275);
or U423 (N_423,N_371,N_392);
nand U424 (N_424,In_283,N_385);
and U425 (N_425,In_14,N_304);
and U426 (N_426,N_354,N_374);
xor U427 (N_427,N_266,N_386);
xnor U428 (N_428,N_370,N_353);
or U429 (N_429,N_357,N_352);
and U430 (N_430,N_380,N_362);
nand U431 (N_431,N_255,N_316);
and U432 (N_432,N_365,N_381);
xor U433 (N_433,N_258,N_351);
nor U434 (N_434,In_342,N_336);
or U435 (N_435,N_369,N_284);
nor U436 (N_436,N_358,In_364);
or U437 (N_437,N_299,N_366);
or U438 (N_438,N_394,In_206);
and U439 (N_439,N_398,In_7);
or U440 (N_440,N_379,N_344);
and U441 (N_441,N_343,N_209);
nor U442 (N_442,N_274,N_313);
and U443 (N_443,N_345,N_311);
or U444 (N_444,N_350,N_321);
nand U445 (N_445,N_399,N_376);
nand U446 (N_446,N_359,N_373);
and U447 (N_447,In_237,In_103);
nor U448 (N_448,N_393,N_75);
or U449 (N_449,N_306,N_49);
and U450 (N_450,N_428,N_400);
and U451 (N_451,N_410,N_409);
xor U452 (N_452,N_421,N_441);
nor U453 (N_453,N_425,N_437);
and U454 (N_454,N_445,N_419);
nor U455 (N_455,N_422,N_440);
nand U456 (N_456,N_402,N_408);
nor U457 (N_457,N_430,N_413);
nand U458 (N_458,N_424,N_411);
nor U459 (N_459,N_423,N_414);
xor U460 (N_460,N_449,N_403);
nand U461 (N_461,N_417,N_420);
nand U462 (N_462,N_446,N_433);
and U463 (N_463,N_447,N_429);
and U464 (N_464,N_416,N_436);
or U465 (N_465,N_442,N_444);
or U466 (N_466,N_438,N_405);
nand U467 (N_467,N_406,N_443);
or U468 (N_468,N_426,N_439);
xor U469 (N_469,N_418,N_434);
nor U470 (N_470,N_412,N_404);
nand U471 (N_471,N_401,N_407);
nor U472 (N_472,N_431,N_448);
nor U473 (N_473,N_415,N_427);
nor U474 (N_474,N_432,N_435);
nor U475 (N_475,N_408,N_426);
and U476 (N_476,N_445,N_440);
and U477 (N_477,N_426,N_407);
or U478 (N_478,N_401,N_400);
and U479 (N_479,N_421,N_419);
nand U480 (N_480,N_417,N_439);
nor U481 (N_481,N_448,N_446);
or U482 (N_482,N_413,N_429);
nor U483 (N_483,N_403,N_439);
and U484 (N_484,N_404,N_437);
nand U485 (N_485,N_426,N_402);
and U486 (N_486,N_428,N_415);
or U487 (N_487,N_427,N_416);
nor U488 (N_488,N_423,N_434);
nand U489 (N_489,N_417,N_442);
and U490 (N_490,N_409,N_430);
nand U491 (N_491,N_446,N_413);
nor U492 (N_492,N_402,N_432);
xnor U493 (N_493,N_413,N_419);
or U494 (N_494,N_448,N_440);
xnor U495 (N_495,N_443,N_416);
nand U496 (N_496,N_443,N_432);
and U497 (N_497,N_428,N_405);
and U498 (N_498,N_420,N_444);
xnor U499 (N_499,N_416,N_449);
nor U500 (N_500,N_454,N_460);
or U501 (N_501,N_461,N_476);
nor U502 (N_502,N_463,N_484);
or U503 (N_503,N_490,N_492);
or U504 (N_504,N_462,N_481);
nor U505 (N_505,N_453,N_477);
and U506 (N_506,N_475,N_471);
and U507 (N_507,N_459,N_496);
and U508 (N_508,N_467,N_486);
nor U509 (N_509,N_487,N_489);
nand U510 (N_510,N_455,N_479);
and U511 (N_511,N_499,N_465);
nand U512 (N_512,N_485,N_483);
or U513 (N_513,N_464,N_452);
and U514 (N_514,N_498,N_472);
nand U515 (N_515,N_451,N_457);
or U516 (N_516,N_474,N_470);
nand U517 (N_517,N_469,N_495);
and U518 (N_518,N_497,N_491);
or U519 (N_519,N_488,N_480);
nand U520 (N_520,N_482,N_458);
and U521 (N_521,N_494,N_493);
or U522 (N_522,N_450,N_456);
or U523 (N_523,N_466,N_478);
nand U524 (N_524,N_468,N_473);
or U525 (N_525,N_459,N_454);
or U526 (N_526,N_451,N_484);
and U527 (N_527,N_478,N_474);
or U528 (N_528,N_466,N_455);
or U529 (N_529,N_477,N_455);
or U530 (N_530,N_466,N_467);
nand U531 (N_531,N_480,N_455);
and U532 (N_532,N_493,N_482);
nor U533 (N_533,N_493,N_472);
nor U534 (N_534,N_465,N_453);
or U535 (N_535,N_457,N_483);
nand U536 (N_536,N_465,N_497);
nor U537 (N_537,N_493,N_469);
or U538 (N_538,N_499,N_466);
nand U539 (N_539,N_494,N_457);
nor U540 (N_540,N_457,N_467);
or U541 (N_541,N_488,N_466);
or U542 (N_542,N_471,N_473);
or U543 (N_543,N_497,N_478);
nor U544 (N_544,N_494,N_465);
nand U545 (N_545,N_478,N_472);
nor U546 (N_546,N_460,N_473);
nor U547 (N_547,N_470,N_464);
nor U548 (N_548,N_498,N_461);
nand U549 (N_549,N_470,N_493);
xor U550 (N_550,N_527,N_532);
nor U551 (N_551,N_520,N_521);
or U552 (N_552,N_531,N_545);
and U553 (N_553,N_544,N_534);
nand U554 (N_554,N_543,N_547);
nor U555 (N_555,N_514,N_530);
nand U556 (N_556,N_502,N_522);
or U557 (N_557,N_507,N_503);
and U558 (N_558,N_542,N_541);
xor U559 (N_559,N_510,N_508);
and U560 (N_560,N_537,N_500);
and U561 (N_561,N_539,N_549);
and U562 (N_562,N_525,N_501);
nand U563 (N_563,N_519,N_511);
or U564 (N_564,N_528,N_506);
xor U565 (N_565,N_512,N_517);
or U566 (N_566,N_509,N_535);
nor U567 (N_567,N_523,N_540);
nand U568 (N_568,N_548,N_533);
and U569 (N_569,N_513,N_518);
or U570 (N_570,N_524,N_536);
or U571 (N_571,N_504,N_515);
nor U572 (N_572,N_505,N_526);
xor U573 (N_573,N_529,N_516);
xor U574 (N_574,N_546,N_538);
nor U575 (N_575,N_500,N_517);
nand U576 (N_576,N_514,N_541);
and U577 (N_577,N_524,N_522);
and U578 (N_578,N_502,N_540);
and U579 (N_579,N_530,N_545);
xnor U580 (N_580,N_500,N_512);
or U581 (N_581,N_538,N_545);
or U582 (N_582,N_520,N_522);
xor U583 (N_583,N_536,N_534);
nand U584 (N_584,N_546,N_507);
nor U585 (N_585,N_530,N_529);
nor U586 (N_586,N_525,N_510);
nand U587 (N_587,N_531,N_519);
and U588 (N_588,N_542,N_546);
nor U589 (N_589,N_539,N_522);
or U590 (N_590,N_515,N_525);
nor U591 (N_591,N_535,N_528);
nand U592 (N_592,N_522,N_544);
nor U593 (N_593,N_523,N_541);
xor U594 (N_594,N_549,N_513);
or U595 (N_595,N_525,N_532);
and U596 (N_596,N_528,N_522);
nor U597 (N_597,N_528,N_505);
nor U598 (N_598,N_548,N_518);
and U599 (N_599,N_539,N_531);
nand U600 (N_600,N_597,N_588);
nor U601 (N_601,N_574,N_596);
xor U602 (N_602,N_561,N_575);
nor U603 (N_603,N_580,N_587);
nor U604 (N_604,N_591,N_567);
nand U605 (N_605,N_555,N_595);
nor U606 (N_606,N_584,N_570);
or U607 (N_607,N_572,N_585);
or U608 (N_608,N_566,N_556);
xnor U609 (N_609,N_550,N_593);
or U610 (N_610,N_573,N_583);
xor U611 (N_611,N_581,N_551);
and U612 (N_612,N_565,N_586);
and U613 (N_613,N_578,N_599);
or U614 (N_614,N_568,N_552);
nor U615 (N_615,N_598,N_554);
or U616 (N_616,N_592,N_553);
or U617 (N_617,N_594,N_576);
nor U618 (N_618,N_560,N_579);
and U619 (N_619,N_569,N_559);
xnor U620 (N_620,N_571,N_558);
nand U621 (N_621,N_590,N_562);
and U622 (N_622,N_589,N_582);
xor U623 (N_623,N_577,N_557);
and U624 (N_624,N_564,N_563);
and U625 (N_625,N_550,N_567);
nor U626 (N_626,N_558,N_567);
and U627 (N_627,N_552,N_597);
nand U628 (N_628,N_565,N_562);
or U629 (N_629,N_574,N_581);
xnor U630 (N_630,N_598,N_560);
and U631 (N_631,N_578,N_566);
nor U632 (N_632,N_560,N_576);
and U633 (N_633,N_595,N_556);
nor U634 (N_634,N_553,N_550);
or U635 (N_635,N_598,N_590);
nand U636 (N_636,N_577,N_568);
or U637 (N_637,N_555,N_591);
or U638 (N_638,N_576,N_552);
or U639 (N_639,N_577,N_554);
and U640 (N_640,N_560,N_589);
and U641 (N_641,N_585,N_554);
nand U642 (N_642,N_564,N_560);
and U643 (N_643,N_574,N_573);
nand U644 (N_644,N_576,N_587);
or U645 (N_645,N_569,N_588);
and U646 (N_646,N_561,N_571);
nand U647 (N_647,N_559,N_573);
nand U648 (N_648,N_583,N_553);
nand U649 (N_649,N_596,N_563);
nand U650 (N_650,N_606,N_636);
or U651 (N_651,N_601,N_635);
or U652 (N_652,N_618,N_648);
xnor U653 (N_653,N_649,N_626);
nor U654 (N_654,N_615,N_639);
or U655 (N_655,N_611,N_642);
xnor U656 (N_656,N_616,N_620);
xnor U657 (N_657,N_628,N_614);
nor U658 (N_658,N_631,N_625);
and U659 (N_659,N_629,N_634);
xnor U660 (N_660,N_641,N_612);
nor U661 (N_661,N_644,N_605);
and U662 (N_662,N_640,N_617);
and U663 (N_663,N_632,N_643);
nand U664 (N_664,N_603,N_624);
nand U665 (N_665,N_621,N_630);
nand U666 (N_666,N_610,N_647);
or U667 (N_667,N_604,N_607);
or U668 (N_668,N_613,N_622);
nand U669 (N_669,N_638,N_608);
xor U670 (N_670,N_600,N_645);
and U671 (N_671,N_623,N_609);
or U672 (N_672,N_627,N_646);
or U673 (N_673,N_619,N_602);
nand U674 (N_674,N_633,N_637);
nand U675 (N_675,N_611,N_643);
or U676 (N_676,N_607,N_612);
or U677 (N_677,N_646,N_606);
nor U678 (N_678,N_627,N_600);
and U679 (N_679,N_624,N_640);
or U680 (N_680,N_635,N_640);
nand U681 (N_681,N_614,N_625);
or U682 (N_682,N_649,N_624);
and U683 (N_683,N_610,N_621);
or U684 (N_684,N_641,N_622);
nor U685 (N_685,N_605,N_640);
and U686 (N_686,N_607,N_611);
nor U687 (N_687,N_623,N_631);
nand U688 (N_688,N_627,N_620);
nand U689 (N_689,N_614,N_644);
nand U690 (N_690,N_617,N_608);
or U691 (N_691,N_602,N_608);
and U692 (N_692,N_622,N_649);
and U693 (N_693,N_635,N_609);
or U694 (N_694,N_622,N_624);
or U695 (N_695,N_643,N_626);
and U696 (N_696,N_604,N_602);
and U697 (N_697,N_630,N_624);
or U698 (N_698,N_644,N_606);
or U699 (N_699,N_607,N_642);
nor U700 (N_700,N_661,N_673);
nand U701 (N_701,N_685,N_678);
nor U702 (N_702,N_657,N_674);
nand U703 (N_703,N_658,N_654);
nand U704 (N_704,N_692,N_695);
or U705 (N_705,N_688,N_671);
xor U706 (N_706,N_656,N_683);
and U707 (N_707,N_689,N_690);
and U708 (N_708,N_681,N_694);
or U709 (N_709,N_665,N_659);
nand U710 (N_710,N_651,N_660);
xnor U711 (N_711,N_664,N_663);
nand U712 (N_712,N_693,N_672);
nand U713 (N_713,N_650,N_668);
nand U714 (N_714,N_680,N_652);
nor U715 (N_715,N_699,N_677);
or U716 (N_716,N_698,N_675);
and U717 (N_717,N_697,N_666);
and U718 (N_718,N_687,N_686);
or U719 (N_719,N_667,N_676);
and U720 (N_720,N_696,N_684);
nand U721 (N_721,N_662,N_670);
and U722 (N_722,N_669,N_691);
nand U723 (N_723,N_682,N_679);
nand U724 (N_724,N_653,N_655);
nor U725 (N_725,N_661,N_653);
nor U726 (N_726,N_687,N_673);
and U727 (N_727,N_696,N_661);
or U728 (N_728,N_654,N_684);
or U729 (N_729,N_677,N_675);
nand U730 (N_730,N_681,N_668);
nand U731 (N_731,N_674,N_688);
or U732 (N_732,N_665,N_685);
nor U733 (N_733,N_696,N_692);
nand U734 (N_734,N_654,N_668);
nor U735 (N_735,N_680,N_656);
and U736 (N_736,N_654,N_671);
xnor U737 (N_737,N_690,N_660);
nand U738 (N_738,N_662,N_680);
nand U739 (N_739,N_675,N_671);
and U740 (N_740,N_692,N_666);
nor U741 (N_741,N_697,N_686);
nand U742 (N_742,N_698,N_678);
and U743 (N_743,N_681,N_660);
nand U744 (N_744,N_664,N_673);
xnor U745 (N_745,N_697,N_674);
nand U746 (N_746,N_694,N_671);
or U747 (N_747,N_667,N_692);
or U748 (N_748,N_675,N_678);
and U749 (N_749,N_657,N_677);
nor U750 (N_750,N_714,N_732);
xor U751 (N_751,N_720,N_712);
nand U752 (N_752,N_723,N_737);
nand U753 (N_753,N_748,N_703);
nor U754 (N_754,N_722,N_729);
nand U755 (N_755,N_702,N_711);
nand U756 (N_756,N_721,N_718);
nor U757 (N_757,N_733,N_704);
or U758 (N_758,N_717,N_710);
nor U759 (N_759,N_716,N_719);
or U760 (N_760,N_707,N_736);
nand U761 (N_761,N_724,N_713);
nor U762 (N_762,N_725,N_706);
xnor U763 (N_763,N_708,N_746);
xnor U764 (N_764,N_700,N_739);
nor U765 (N_765,N_747,N_745);
nor U766 (N_766,N_705,N_743);
nor U767 (N_767,N_740,N_701);
nor U768 (N_768,N_726,N_727);
or U769 (N_769,N_741,N_749);
or U770 (N_770,N_734,N_730);
and U771 (N_771,N_735,N_728);
and U772 (N_772,N_742,N_709);
nand U773 (N_773,N_744,N_738);
and U774 (N_774,N_731,N_715);
nand U775 (N_775,N_723,N_705);
nor U776 (N_776,N_724,N_749);
xnor U777 (N_777,N_742,N_721);
nand U778 (N_778,N_730,N_724);
nor U779 (N_779,N_719,N_714);
xor U780 (N_780,N_717,N_723);
or U781 (N_781,N_747,N_718);
nand U782 (N_782,N_708,N_709);
or U783 (N_783,N_734,N_722);
xnor U784 (N_784,N_742,N_710);
and U785 (N_785,N_714,N_720);
and U786 (N_786,N_740,N_723);
nor U787 (N_787,N_718,N_733);
nor U788 (N_788,N_701,N_736);
and U789 (N_789,N_733,N_711);
xor U790 (N_790,N_730,N_702);
nand U791 (N_791,N_727,N_729);
and U792 (N_792,N_717,N_724);
or U793 (N_793,N_723,N_716);
and U794 (N_794,N_703,N_709);
xor U795 (N_795,N_749,N_710);
or U796 (N_796,N_737,N_743);
xor U797 (N_797,N_710,N_730);
or U798 (N_798,N_736,N_733);
or U799 (N_799,N_721,N_711);
nand U800 (N_800,N_784,N_774);
nand U801 (N_801,N_795,N_769);
or U802 (N_802,N_751,N_791);
or U803 (N_803,N_776,N_777);
nand U804 (N_804,N_764,N_799);
nand U805 (N_805,N_787,N_792);
and U806 (N_806,N_770,N_782);
nor U807 (N_807,N_762,N_786);
nor U808 (N_808,N_759,N_775);
and U809 (N_809,N_797,N_785);
nor U810 (N_810,N_798,N_761);
nand U811 (N_811,N_789,N_768);
nor U812 (N_812,N_790,N_779);
nor U813 (N_813,N_781,N_778);
or U814 (N_814,N_760,N_771);
nand U815 (N_815,N_783,N_750);
nand U816 (N_816,N_788,N_758);
nor U817 (N_817,N_765,N_766);
nor U818 (N_818,N_772,N_756);
and U819 (N_819,N_757,N_763);
and U820 (N_820,N_794,N_767);
and U821 (N_821,N_752,N_754);
nand U822 (N_822,N_753,N_773);
nand U823 (N_823,N_780,N_755);
nand U824 (N_824,N_796,N_793);
nor U825 (N_825,N_781,N_750);
nor U826 (N_826,N_786,N_792);
or U827 (N_827,N_798,N_751);
xor U828 (N_828,N_750,N_757);
or U829 (N_829,N_774,N_762);
or U830 (N_830,N_794,N_760);
nand U831 (N_831,N_791,N_769);
nand U832 (N_832,N_750,N_759);
or U833 (N_833,N_792,N_779);
and U834 (N_834,N_781,N_774);
or U835 (N_835,N_770,N_761);
or U836 (N_836,N_762,N_755);
and U837 (N_837,N_752,N_769);
nor U838 (N_838,N_764,N_773);
and U839 (N_839,N_760,N_786);
nand U840 (N_840,N_788,N_772);
and U841 (N_841,N_753,N_781);
nor U842 (N_842,N_786,N_797);
nor U843 (N_843,N_771,N_769);
nand U844 (N_844,N_771,N_782);
nor U845 (N_845,N_761,N_793);
nor U846 (N_846,N_799,N_768);
and U847 (N_847,N_793,N_780);
xor U848 (N_848,N_786,N_780);
nor U849 (N_849,N_798,N_791);
nor U850 (N_850,N_849,N_801);
nand U851 (N_851,N_808,N_840);
nor U852 (N_852,N_802,N_817);
nand U853 (N_853,N_833,N_838);
and U854 (N_854,N_848,N_821);
and U855 (N_855,N_824,N_827);
and U856 (N_856,N_845,N_829);
xnor U857 (N_857,N_823,N_807);
nand U858 (N_858,N_814,N_815);
or U859 (N_859,N_803,N_818);
nand U860 (N_860,N_806,N_813);
nand U861 (N_861,N_800,N_836);
nor U862 (N_862,N_837,N_844);
nor U863 (N_863,N_846,N_842);
or U864 (N_864,N_828,N_826);
or U865 (N_865,N_822,N_839);
nor U866 (N_866,N_825,N_809);
nand U867 (N_867,N_804,N_812);
or U868 (N_868,N_805,N_843);
xor U869 (N_869,N_831,N_820);
nand U870 (N_870,N_819,N_835);
nor U871 (N_871,N_830,N_810);
xor U872 (N_872,N_811,N_816);
nand U873 (N_873,N_841,N_834);
and U874 (N_874,N_832,N_847);
and U875 (N_875,N_846,N_809);
and U876 (N_876,N_841,N_825);
nand U877 (N_877,N_801,N_839);
and U878 (N_878,N_828,N_816);
nor U879 (N_879,N_849,N_848);
xnor U880 (N_880,N_817,N_800);
or U881 (N_881,N_821,N_845);
or U882 (N_882,N_848,N_810);
nor U883 (N_883,N_835,N_804);
nand U884 (N_884,N_819,N_811);
and U885 (N_885,N_821,N_835);
nand U886 (N_886,N_822,N_801);
or U887 (N_887,N_824,N_801);
or U888 (N_888,N_846,N_823);
nor U889 (N_889,N_832,N_840);
xnor U890 (N_890,N_833,N_822);
nor U891 (N_891,N_819,N_821);
or U892 (N_892,N_822,N_849);
nor U893 (N_893,N_820,N_848);
nor U894 (N_894,N_832,N_810);
nor U895 (N_895,N_841,N_810);
and U896 (N_896,N_836,N_818);
nand U897 (N_897,N_846,N_821);
xor U898 (N_898,N_842,N_813);
xnor U899 (N_899,N_823,N_837);
nand U900 (N_900,N_871,N_878);
nor U901 (N_901,N_885,N_892);
and U902 (N_902,N_883,N_880);
nand U903 (N_903,N_874,N_890);
nor U904 (N_904,N_867,N_881);
and U905 (N_905,N_891,N_884);
xnor U906 (N_906,N_886,N_852);
or U907 (N_907,N_856,N_855);
nor U908 (N_908,N_862,N_877);
or U909 (N_909,N_894,N_876);
xor U910 (N_910,N_869,N_860);
nor U911 (N_911,N_872,N_858);
nand U912 (N_912,N_864,N_863);
nor U913 (N_913,N_893,N_896);
or U914 (N_914,N_861,N_865);
nand U915 (N_915,N_875,N_859);
and U916 (N_916,N_850,N_873);
nor U917 (N_917,N_870,N_898);
nand U918 (N_918,N_851,N_888);
nor U919 (N_919,N_879,N_857);
nor U920 (N_920,N_868,N_895);
or U921 (N_921,N_854,N_889);
or U922 (N_922,N_853,N_899);
or U923 (N_923,N_897,N_866);
or U924 (N_924,N_887,N_882);
nand U925 (N_925,N_856,N_887);
or U926 (N_926,N_893,N_850);
xor U927 (N_927,N_873,N_877);
nor U928 (N_928,N_877,N_869);
nor U929 (N_929,N_890,N_857);
or U930 (N_930,N_850,N_887);
nor U931 (N_931,N_881,N_877);
nand U932 (N_932,N_898,N_878);
nand U933 (N_933,N_858,N_874);
nand U934 (N_934,N_854,N_865);
nand U935 (N_935,N_899,N_855);
and U936 (N_936,N_892,N_850);
or U937 (N_937,N_884,N_863);
and U938 (N_938,N_886,N_867);
and U939 (N_939,N_896,N_881);
or U940 (N_940,N_868,N_890);
or U941 (N_941,N_880,N_870);
nand U942 (N_942,N_858,N_886);
or U943 (N_943,N_866,N_882);
nor U944 (N_944,N_884,N_868);
nor U945 (N_945,N_880,N_869);
nor U946 (N_946,N_874,N_899);
or U947 (N_947,N_850,N_890);
and U948 (N_948,N_877,N_887);
and U949 (N_949,N_854,N_879);
and U950 (N_950,N_928,N_922);
nand U951 (N_951,N_939,N_924);
and U952 (N_952,N_907,N_945);
nand U953 (N_953,N_940,N_944);
nand U954 (N_954,N_916,N_908);
nand U955 (N_955,N_925,N_936);
and U956 (N_956,N_927,N_919);
nor U957 (N_957,N_903,N_937);
nor U958 (N_958,N_909,N_933);
or U959 (N_959,N_910,N_949);
nor U960 (N_960,N_911,N_920);
nor U961 (N_961,N_912,N_946);
xor U962 (N_962,N_902,N_906);
nand U963 (N_963,N_943,N_904);
nand U964 (N_964,N_929,N_921);
nand U965 (N_965,N_947,N_914);
xnor U966 (N_966,N_935,N_942);
nor U967 (N_967,N_915,N_917);
or U968 (N_968,N_932,N_901);
nand U969 (N_969,N_948,N_905);
and U970 (N_970,N_918,N_934);
and U971 (N_971,N_923,N_913);
and U972 (N_972,N_900,N_930);
and U973 (N_973,N_938,N_941);
or U974 (N_974,N_926,N_931);
and U975 (N_975,N_930,N_925);
or U976 (N_976,N_922,N_907);
or U977 (N_977,N_935,N_945);
nor U978 (N_978,N_942,N_939);
nand U979 (N_979,N_943,N_906);
or U980 (N_980,N_949,N_922);
nand U981 (N_981,N_924,N_900);
or U982 (N_982,N_927,N_909);
nor U983 (N_983,N_936,N_912);
nand U984 (N_984,N_926,N_906);
or U985 (N_985,N_941,N_902);
or U986 (N_986,N_927,N_913);
and U987 (N_987,N_922,N_929);
and U988 (N_988,N_909,N_911);
nor U989 (N_989,N_908,N_902);
and U990 (N_990,N_916,N_918);
nand U991 (N_991,N_921,N_916);
or U992 (N_992,N_902,N_922);
or U993 (N_993,N_920,N_916);
xor U994 (N_994,N_942,N_944);
and U995 (N_995,N_915,N_902);
or U996 (N_996,N_921,N_939);
nand U997 (N_997,N_939,N_930);
nor U998 (N_998,N_937,N_948);
and U999 (N_999,N_938,N_946);
nor U1000 (N_1000,N_953,N_957);
or U1001 (N_1001,N_978,N_955);
nor U1002 (N_1002,N_991,N_998);
and U1003 (N_1003,N_976,N_983);
nand U1004 (N_1004,N_999,N_971);
or U1005 (N_1005,N_975,N_974);
or U1006 (N_1006,N_958,N_965);
or U1007 (N_1007,N_981,N_962);
xor U1008 (N_1008,N_970,N_964);
nor U1009 (N_1009,N_973,N_985);
and U1010 (N_1010,N_996,N_995);
nand U1011 (N_1011,N_950,N_988);
nand U1012 (N_1012,N_972,N_986);
nand U1013 (N_1013,N_967,N_963);
and U1014 (N_1014,N_960,N_987);
nand U1015 (N_1015,N_989,N_990);
xor U1016 (N_1016,N_968,N_980);
nand U1017 (N_1017,N_984,N_969);
nand U1018 (N_1018,N_994,N_992);
and U1019 (N_1019,N_997,N_951);
nand U1020 (N_1020,N_952,N_966);
and U1021 (N_1021,N_961,N_982);
nand U1022 (N_1022,N_979,N_954);
or U1023 (N_1023,N_993,N_959);
nand U1024 (N_1024,N_956,N_977);
or U1025 (N_1025,N_968,N_997);
or U1026 (N_1026,N_997,N_995);
and U1027 (N_1027,N_953,N_989);
nor U1028 (N_1028,N_994,N_968);
nor U1029 (N_1029,N_959,N_998);
or U1030 (N_1030,N_993,N_989);
and U1031 (N_1031,N_956,N_961);
nor U1032 (N_1032,N_986,N_980);
nor U1033 (N_1033,N_967,N_957);
xnor U1034 (N_1034,N_964,N_965);
nor U1035 (N_1035,N_997,N_987);
and U1036 (N_1036,N_956,N_975);
or U1037 (N_1037,N_999,N_966);
nand U1038 (N_1038,N_975,N_961);
xnor U1039 (N_1039,N_972,N_989);
nand U1040 (N_1040,N_966,N_956);
nand U1041 (N_1041,N_969,N_972);
or U1042 (N_1042,N_978,N_960);
and U1043 (N_1043,N_973,N_969);
nand U1044 (N_1044,N_977,N_998);
and U1045 (N_1045,N_968,N_993);
nor U1046 (N_1046,N_989,N_991);
and U1047 (N_1047,N_981,N_974);
nor U1048 (N_1048,N_981,N_967);
nor U1049 (N_1049,N_968,N_984);
and U1050 (N_1050,N_1030,N_1045);
or U1051 (N_1051,N_1012,N_1001);
nand U1052 (N_1052,N_1021,N_1013);
nand U1053 (N_1053,N_1004,N_1016);
nor U1054 (N_1054,N_1000,N_1024);
or U1055 (N_1055,N_1039,N_1022);
nor U1056 (N_1056,N_1031,N_1017);
nor U1057 (N_1057,N_1032,N_1041);
and U1058 (N_1058,N_1009,N_1033);
nor U1059 (N_1059,N_1020,N_1008);
nor U1060 (N_1060,N_1038,N_1046);
nor U1061 (N_1061,N_1010,N_1026);
nor U1062 (N_1062,N_1036,N_1005);
and U1063 (N_1063,N_1042,N_1027);
nor U1064 (N_1064,N_1029,N_1018);
or U1065 (N_1065,N_1034,N_1002);
nand U1066 (N_1066,N_1006,N_1040);
or U1067 (N_1067,N_1028,N_1049);
nand U1068 (N_1068,N_1025,N_1035);
and U1069 (N_1069,N_1003,N_1023);
nor U1070 (N_1070,N_1019,N_1015);
nor U1071 (N_1071,N_1007,N_1048);
and U1072 (N_1072,N_1037,N_1044);
or U1073 (N_1073,N_1014,N_1043);
nor U1074 (N_1074,N_1047,N_1011);
nor U1075 (N_1075,N_1031,N_1036);
nor U1076 (N_1076,N_1042,N_1013);
and U1077 (N_1077,N_1048,N_1019);
xor U1078 (N_1078,N_1010,N_1035);
xor U1079 (N_1079,N_1006,N_1023);
nand U1080 (N_1080,N_1018,N_1009);
and U1081 (N_1081,N_1048,N_1003);
and U1082 (N_1082,N_1018,N_1048);
or U1083 (N_1083,N_1028,N_1037);
nand U1084 (N_1084,N_1032,N_1026);
nand U1085 (N_1085,N_1041,N_1030);
nor U1086 (N_1086,N_1044,N_1018);
and U1087 (N_1087,N_1049,N_1010);
and U1088 (N_1088,N_1035,N_1036);
xor U1089 (N_1089,N_1020,N_1029);
and U1090 (N_1090,N_1033,N_1035);
nand U1091 (N_1091,N_1046,N_1041);
and U1092 (N_1092,N_1009,N_1032);
and U1093 (N_1093,N_1028,N_1009);
xnor U1094 (N_1094,N_1047,N_1006);
and U1095 (N_1095,N_1031,N_1025);
xnor U1096 (N_1096,N_1015,N_1037);
or U1097 (N_1097,N_1041,N_1040);
nand U1098 (N_1098,N_1006,N_1008);
xor U1099 (N_1099,N_1015,N_1023);
or U1100 (N_1100,N_1082,N_1074);
xor U1101 (N_1101,N_1097,N_1070);
nor U1102 (N_1102,N_1085,N_1072);
nor U1103 (N_1103,N_1093,N_1062);
nor U1104 (N_1104,N_1054,N_1058);
and U1105 (N_1105,N_1091,N_1096);
or U1106 (N_1106,N_1090,N_1063);
nand U1107 (N_1107,N_1092,N_1061);
nor U1108 (N_1108,N_1056,N_1051);
or U1109 (N_1109,N_1077,N_1084);
nor U1110 (N_1110,N_1081,N_1059);
nor U1111 (N_1111,N_1087,N_1078);
nor U1112 (N_1112,N_1053,N_1064);
and U1113 (N_1113,N_1076,N_1073);
xnor U1114 (N_1114,N_1069,N_1080);
and U1115 (N_1115,N_1098,N_1068);
or U1116 (N_1116,N_1088,N_1075);
or U1117 (N_1117,N_1094,N_1095);
nand U1118 (N_1118,N_1060,N_1086);
or U1119 (N_1119,N_1083,N_1071);
and U1120 (N_1120,N_1050,N_1066);
nand U1121 (N_1121,N_1089,N_1067);
nor U1122 (N_1122,N_1099,N_1052);
nor U1123 (N_1123,N_1065,N_1055);
and U1124 (N_1124,N_1079,N_1057);
nand U1125 (N_1125,N_1057,N_1074);
xor U1126 (N_1126,N_1068,N_1077);
nor U1127 (N_1127,N_1094,N_1070);
nor U1128 (N_1128,N_1069,N_1087);
and U1129 (N_1129,N_1063,N_1095);
or U1130 (N_1130,N_1099,N_1086);
or U1131 (N_1131,N_1082,N_1077);
and U1132 (N_1132,N_1098,N_1086);
nand U1133 (N_1133,N_1056,N_1057);
or U1134 (N_1134,N_1078,N_1099);
xor U1135 (N_1135,N_1088,N_1062);
xnor U1136 (N_1136,N_1062,N_1052);
xor U1137 (N_1137,N_1072,N_1076);
or U1138 (N_1138,N_1085,N_1057);
or U1139 (N_1139,N_1066,N_1077);
and U1140 (N_1140,N_1098,N_1069);
nor U1141 (N_1141,N_1092,N_1080);
nand U1142 (N_1142,N_1055,N_1074);
or U1143 (N_1143,N_1067,N_1065);
or U1144 (N_1144,N_1090,N_1050);
nor U1145 (N_1145,N_1065,N_1054);
or U1146 (N_1146,N_1064,N_1076);
or U1147 (N_1147,N_1079,N_1084);
xnor U1148 (N_1148,N_1078,N_1090);
nor U1149 (N_1149,N_1059,N_1077);
and U1150 (N_1150,N_1108,N_1113);
xnor U1151 (N_1151,N_1123,N_1126);
or U1152 (N_1152,N_1111,N_1122);
and U1153 (N_1153,N_1118,N_1101);
and U1154 (N_1154,N_1100,N_1148);
nand U1155 (N_1155,N_1144,N_1137);
nand U1156 (N_1156,N_1119,N_1125);
nor U1157 (N_1157,N_1115,N_1141);
or U1158 (N_1158,N_1104,N_1116);
nand U1159 (N_1159,N_1105,N_1102);
nor U1160 (N_1160,N_1147,N_1129);
or U1161 (N_1161,N_1107,N_1140);
or U1162 (N_1162,N_1143,N_1136);
xor U1163 (N_1163,N_1127,N_1103);
and U1164 (N_1164,N_1142,N_1134);
nand U1165 (N_1165,N_1114,N_1117);
or U1166 (N_1166,N_1124,N_1145);
xnor U1167 (N_1167,N_1135,N_1132);
and U1168 (N_1168,N_1131,N_1120);
nand U1169 (N_1169,N_1109,N_1128);
nand U1170 (N_1170,N_1138,N_1110);
or U1171 (N_1171,N_1112,N_1130);
or U1172 (N_1172,N_1121,N_1146);
and U1173 (N_1173,N_1149,N_1139);
nand U1174 (N_1174,N_1133,N_1106);
or U1175 (N_1175,N_1149,N_1109);
or U1176 (N_1176,N_1137,N_1125);
xnor U1177 (N_1177,N_1113,N_1139);
or U1178 (N_1178,N_1104,N_1112);
nand U1179 (N_1179,N_1118,N_1146);
and U1180 (N_1180,N_1101,N_1115);
and U1181 (N_1181,N_1145,N_1140);
or U1182 (N_1182,N_1105,N_1100);
nand U1183 (N_1183,N_1146,N_1101);
or U1184 (N_1184,N_1125,N_1106);
nor U1185 (N_1185,N_1118,N_1140);
nand U1186 (N_1186,N_1109,N_1103);
nand U1187 (N_1187,N_1132,N_1146);
and U1188 (N_1188,N_1100,N_1106);
or U1189 (N_1189,N_1105,N_1114);
nand U1190 (N_1190,N_1101,N_1145);
or U1191 (N_1191,N_1134,N_1147);
and U1192 (N_1192,N_1108,N_1127);
nand U1193 (N_1193,N_1134,N_1146);
nor U1194 (N_1194,N_1133,N_1108);
nor U1195 (N_1195,N_1147,N_1121);
nand U1196 (N_1196,N_1133,N_1128);
and U1197 (N_1197,N_1146,N_1106);
nor U1198 (N_1198,N_1112,N_1143);
nor U1199 (N_1199,N_1107,N_1121);
xnor U1200 (N_1200,N_1190,N_1150);
or U1201 (N_1201,N_1194,N_1188);
nor U1202 (N_1202,N_1170,N_1153);
and U1203 (N_1203,N_1155,N_1185);
or U1204 (N_1204,N_1189,N_1173);
xnor U1205 (N_1205,N_1193,N_1159);
xor U1206 (N_1206,N_1179,N_1199);
nand U1207 (N_1207,N_1186,N_1184);
xor U1208 (N_1208,N_1161,N_1175);
nor U1209 (N_1209,N_1168,N_1177);
and U1210 (N_1210,N_1192,N_1157);
nor U1211 (N_1211,N_1187,N_1195);
and U1212 (N_1212,N_1196,N_1191);
nand U1213 (N_1213,N_1198,N_1167);
nand U1214 (N_1214,N_1154,N_1166);
nor U1215 (N_1215,N_1156,N_1152);
nor U1216 (N_1216,N_1174,N_1171);
and U1217 (N_1217,N_1165,N_1183);
nor U1218 (N_1218,N_1176,N_1151);
or U1219 (N_1219,N_1182,N_1172);
nor U1220 (N_1220,N_1163,N_1197);
xnor U1221 (N_1221,N_1181,N_1160);
nand U1222 (N_1222,N_1158,N_1162);
and U1223 (N_1223,N_1180,N_1178);
nand U1224 (N_1224,N_1164,N_1169);
or U1225 (N_1225,N_1176,N_1177);
nand U1226 (N_1226,N_1177,N_1199);
nor U1227 (N_1227,N_1173,N_1179);
nor U1228 (N_1228,N_1154,N_1171);
nor U1229 (N_1229,N_1197,N_1176);
or U1230 (N_1230,N_1151,N_1152);
xnor U1231 (N_1231,N_1157,N_1188);
nor U1232 (N_1232,N_1166,N_1191);
nand U1233 (N_1233,N_1170,N_1152);
nor U1234 (N_1234,N_1170,N_1150);
nand U1235 (N_1235,N_1152,N_1173);
nand U1236 (N_1236,N_1190,N_1155);
nand U1237 (N_1237,N_1169,N_1170);
or U1238 (N_1238,N_1152,N_1158);
nand U1239 (N_1239,N_1179,N_1171);
nand U1240 (N_1240,N_1167,N_1158);
nor U1241 (N_1241,N_1173,N_1154);
nor U1242 (N_1242,N_1190,N_1192);
or U1243 (N_1243,N_1172,N_1152);
or U1244 (N_1244,N_1167,N_1173);
nand U1245 (N_1245,N_1187,N_1184);
nor U1246 (N_1246,N_1196,N_1189);
or U1247 (N_1247,N_1168,N_1183);
or U1248 (N_1248,N_1167,N_1199);
nand U1249 (N_1249,N_1189,N_1192);
nand U1250 (N_1250,N_1228,N_1226);
nor U1251 (N_1251,N_1229,N_1237);
or U1252 (N_1252,N_1217,N_1204);
and U1253 (N_1253,N_1219,N_1205);
nand U1254 (N_1254,N_1209,N_1222);
nand U1255 (N_1255,N_1244,N_1234);
and U1256 (N_1256,N_1206,N_1200);
and U1257 (N_1257,N_1227,N_1215);
nor U1258 (N_1258,N_1242,N_1203);
and U1259 (N_1259,N_1238,N_1207);
nor U1260 (N_1260,N_1201,N_1212);
nand U1261 (N_1261,N_1239,N_1249);
nor U1262 (N_1262,N_1240,N_1218);
and U1263 (N_1263,N_1232,N_1223);
nand U1264 (N_1264,N_1247,N_1211);
or U1265 (N_1265,N_1231,N_1246);
and U1266 (N_1266,N_1216,N_1208);
and U1267 (N_1267,N_1224,N_1245);
nor U1268 (N_1268,N_1230,N_1233);
nor U1269 (N_1269,N_1236,N_1221);
and U1270 (N_1270,N_1225,N_1243);
or U1271 (N_1271,N_1241,N_1235);
and U1272 (N_1272,N_1213,N_1214);
and U1273 (N_1273,N_1248,N_1202);
nand U1274 (N_1274,N_1220,N_1210);
and U1275 (N_1275,N_1231,N_1229);
and U1276 (N_1276,N_1243,N_1235);
or U1277 (N_1277,N_1209,N_1249);
and U1278 (N_1278,N_1207,N_1216);
nor U1279 (N_1279,N_1223,N_1241);
nor U1280 (N_1280,N_1212,N_1233);
nor U1281 (N_1281,N_1228,N_1238);
nor U1282 (N_1282,N_1233,N_1216);
or U1283 (N_1283,N_1222,N_1232);
nor U1284 (N_1284,N_1248,N_1200);
nor U1285 (N_1285,N_1211,N_1235);
and U1286 (N_1286,N_1205,N_1201);
or U1287 (N_1287,N_1201,N_1222);
nand U1288 (N_1288,N_1219,N_1221);
nor U1289 (N_1289,N_1209,N_1220);
nor U1290 (N_1290,N_1227,N_1248);
nand U1291 (N_1291,N_1200,N_1227);
and U1292 (N_1292,N_1249,N_1222);
or U1293 (N_1293,N_1205,N_1202);
or U1294 (N_1294,N_1223,N_1230);
nor U1295 (N_1295,N_1203,N_1208);
or U1296 (N_1296,N_1229,N_1210);
or U1297 (N_1297,N_1236,N_1235);
nand U1298 (N_1298,N_1207,N_1215);
nor U1299 (N_1299,N_1203,N_1230);
and U1300 (N_1300,N_1298,N_1280);
and U1301 (N_1301,N_1294,N_1289);
xor U1302 (N_1302,N_1275,N_1296);
or U1303 (N_1303,N_1299,N_1254);
and U1304 (N_1304,N_1293,N_1291);
and U1305 (N_1305,N_1252,N_1277);
nand U1306 (N_1306,N_1251,N_1284);
nand U1307 (N_1307,N_1255,N_1272);
nand U1308 (N_1308,N_1253,N_1273);
nand U1309 (N_1309,N_1297,N_1282);
nor U1310 (N_1310,N_1290,N_1269);
nand U1311 (N_1311,N_1281,N_1286);
nor U1312 (N_1312,N_1264,N_1256);
nor U1313 (N_1313,N_1283,N_1288);
or U1314 (N_1314,N_1274,N_1265);
nor U1315 (N_1315,N_1260,N_1270);
xor U1316 (N_1316,N_1279,N_1278);
nand U1317 (N_1317,N_1250,N_1261);
nor U1318 (N_1318,N_1268,N_1262);
xnor U1319 (N_1319,N_1285,N_1276);
and U1320 (N_1320,N_1292,N_1259);
nor U1321 (N_1321,N_1266,N_1263);
xor U1322 (N_1322,N_1295,N_1257);
nor U1323 (N_1323,N_1287,N_1271);
or U1324 (N_1324,N_1258,N_1267);
nand U1325 (N_1325,N_1253,N_1269);
nand U1326 (N_1326,N_1273,N_1297);
nand U1327 (N_1327,N_1257,N_1297);
xnor U1328 (N_1328,N_1272,N_1270);
nand U1329 (N_1329,N_1293,N_1296);
nor U1330 (N_1330,N_1268,N_1290);
nand U1331 (N_1331,N_1274,N_1291);
and U1332 (N_1332,N_1278,N_1296);
and U1333 (N_1333,N_1277,N_1264);
or U1334 (N_1334,N_1285,N_1264);
nor U1335 (N_1335,N_1251,N_1291);
nand U1336 (N_1336,N_1299,N_1262);
and U1337 (N_1337,N_1270,N_1299);
or U1338 (N_1338,N_1251,N_1264);
xnor U1339 (N_1339,N_1298,N_1288);
nor U1340 (N_1340,N_1257,N_1258);
nand U1341 (N_1341,N_1296,N_1280);
nor U1342 (N_1342,N_1285,N_1282);
nand U1343 (N_1343,N_1292,N_1269);
nand U1344 (N_1344,N_1268,N_1254);
and U1345 (N_1345,N_1265,N_1252);
and U1346 (N_1346,N_1260,N_1297);
xnor U1347 (N_1347,N_1294,N_1256);
and U1348 (N_1348,N_1277,N_1285);
nor U1349 (N_1349,N_1260,N_1294);
or U1350 (N_1350,N_1306,N_1331);
nor U1351 (N_1351,N_1303,N_1339);
nand U1352 (N_1352,N_1349,N_1300);
xor U1353 (N_1353,N_1341,N_1333);
nor U1354 (N_1354,N_1310,N_1322);
and U1355 (N_1355,N_1334,N_1343);
nor U1356 (N_1356,N_1348,N_1313);
or U1357 (N_1357,N_1315,N_1318);
and U1358 (N_1358,N_1338,N_1328);
and U1359 (N_1359,N_1305,N_1337);
or U1360 (N_1360,N_1340,N_1324);
and U1361 (N_1361,N_1301,N_1335);
and U1362 (N_1362,N_1347,N_1336);
or U1363 (N_1363,N_1329,N_1320);
nand U1364 (N_1364,N_1330,N_1345);
nand U1365 (N_1365,N_1344,N_1346);
nand U1366 (N_1366,N_1319,N_1323);
or U1367 (N_1367,N_1325,N_1321);
nand U1368 (N_1368,N_1309,N_1316);
or U1369 (N_1369,N_1314,N_1326);
or U1370 (N_1370,N_1302,N_1332);
nor U1371 (N_1371,N_1311,N_1308);
xor U1372 (N_1372,N_1327,N_1312);
and U1373 (N_1373,N_1307,N_1342);
nor U1374 (N_1374,N_1317,N_1304);
nor U1375 (N_1375,N_1314,N_1340);
or U1376 (N_1376,N_1325,N_1333);
or U1377 (N_1377,N_1338,N_1345);
and U1378 (N_1378,N_1339,N_1342);
or U1379 (N_1379,N_1300,N_1302);
nand U1380 (N_1380,N_1342,N_1334);
nand U1381 (N_1381,N_1301,N_1321);
or U1382 (N_1382,N_1346,N_1314);
xor U1383 (N_1383,N_1320,N_1317);
nand U1384 (N_1384,N_1326,N_1320);
and U1385 (N_1385,N_1304,N_1344);
or U1386 (N_1386,N_1333,N_1313);
nor U1387 (N_1387,N_1333,N_1335);
and U1388 (N_1388,N_1347,N_1313);
nand U1389 (N_1389,N_1309,N_1321);
and U1390 (N_1390,N_1344,N_1300);
or U1391 (N_1391,N_1301,N_1308);
nand U1392 (N_1392,N_1304,N_1345);
nand U1393 (N_1393,N_1332,N_1313);
or U1394 (N_1394,N_1316,N_1313);
and U1395 (N_1395,N_1316,N_1307);
and U1396 (N_1396,N_1345,N_1310);
nor U1397 (N_1397,N_1311,N_1301);
nand U1398 (N_1398,N_1346,N_1327);
nor U1399 (N_1399,N_1323,N_1320);
nor U1400 (N_1400,N_1351,N_1382);
xnor U1401 (N_1401,N_1386,N_1389);
and U1402 (N_1402,N_1367,N_1352);
and U1403 (N_1403,N_1365,N_1376);
nor U1404 (N_1404,N_1356,N_1358);
or U1405 (N_1405,N_1388,N_1384);
nand U1406 (N_1406,N_1395,N_1374);
or U1407 (N_1407,N_1394,N_1387);
or U1408 (N_1408,N_1359,N_1363);
nand U1409 (N_1409,N_1371,N_1381);
or U1410 (N_1410,N_1391,N_1393);
or U1411 (N_1411,N_1364,N_1357);
nor U1412 (N_1412,N_1362,N_1383);
nand U1413 (N_1413,N_1377,N_1373);
or U1414 (N_1414,N_1390,N_1370);
nor U1415 (N_1415,N_1375,N_1369);
nand U1416 (N_1416,N_1399,N_1379);
nand U1417 (N_1417,N_1353,N_1354);
and U1418 (N_1418,N_1360,N_1355);
nand U1419 (N_1419,N_1372,N_1361);
and U1420 (N_1420,N_1397,N_1350);
and U1421 (N_1421,N_1380,N_1378);
nand U1422 (N_1422,N_1385,N_1366);
nand U1423 (N_1423,N_1392,N_1368);
nand U1424 (N_1424,N_1396,N_1398);
xnor U1425 (N_1425,N_1381,N_1380);
nand U1426 (N_1426,N_1363,N_1378);
nand U1427 (N_1427,N_1379,N_1361);
nand U1428 (N_1428,N_1384,N_1374);
nor U1429 (N_1429,N_1369,N_1372);
and U1430 (N_1430,N_1372,N_1354);
nand U1431 (N_1431,N_1378,N_1394);
and U1432 (N_1432,N_1393,N_1354);
and U1433 (N_1433,N_1356,N_1383);
xnor U1434 (N_1434,N_1356,N_1397);
xor U1435 (N_1435,N_1384,N_1356);
nor U1436 (N_1436,N_1389,N_1359);
nor U1437 (N_1437,N_1373,N_1363);
and U1438 (N_1438,N_1363,N_1354);
nor U1439 (N_1439,N_1391,N_1352);
nor U1440 (N_1440,N_1351,N_1387);
nor U1441 (N_1441,N_1360,N_1389);
nor U1442 (N_1442,N_1361,N_1350);
and U1443 (N_1443,N_1380,N_1392);
or U1444 (N_1444,N_1392,N_1399);
nor U1445 (N_1445,N_1381,N_1350);
nor U1446 (N_1446,N_1375,N_1364);
and U1447 (N_1447,N_1379,N_1388);
xor U1448 (N_1448,N_1353,N_1352);
xnor U1449 (N_1449,N_1392,N_1377);
or U1450 (N_1450,N_1402,N_1427);
or U1451 (N_1451,N_1433,N_1432);
nor U1452 (N_1452,N_1401,N_1403);
or U1453 (N_1453,N_1431,N_1425);
nor U1454 (N_1454,N_1426,N_1412);
nand U1455 (N_1455,N_1438,N_1440);
or U1456 (N_1456,N_1430,N_1405);
nand U1457 (N_1457,N_1423,N_1441);
nand U1458 (N_1458,N_1413,N_1437);
or U1459 (N_1459,N_1447,N_1429);
or U1460 (N_1460,N_1404,N_1406);
or U1461 (N_1461,N_1421,N_1411);
or U1462 (N_1462,N_1448,N_1410);
or U1463 (N_1463,N_1419,N_1434);
nand U1464 (N_1464,N_1414,N_1409);
and U1465 (N_1465,N_1443,N_1400);
xnor U1466 (N_1466,N_1408,N_1420);
nor U1467 (N_1467,N_1417,N_1435);
and U1468 (N_1468,N_1428,N_1418);
nand U1469 (N_1469,N_1439,N_1422);
and U1470 (N_1470,N_1449,N_1424);
nor U1471 (N_1471,N_1436,N_1444);
or U1472 (N_1472,N_1407,N_1416);
nand U1473 (N_1473,N_1446,N_1415);
nor U1474 (N_1474,N_1442,N_1445);
xor U1475 (N_1475,N_1446,N_1414);
or U1476 (N_1476,N_1439,N_1401);
xor U1477 (N_1477,N_1427,N_1448);
nor U1478 (N_1478,N_1415,N_1437);
nor U1479 (N_1479,N_1412,N_1443);
and U1480 (N_1480,N_1415,N_1408);
nor U1481 (N_1481,N_1427,N_1411);
nand U1482 (N_1482,N_1445,N_1439);
and U1483 (N_1483,N_1439,N_1435);
xor U1484 (N_1484,N_1424,N_1405);
and U1485 (N_1485,N_1413,N_1418);
or U1486 (N_1486,N_1424,N_1419);
nand U1487 (N_1487,N_1443,N_1445);
nor U1488 (N_1488,N_1426,N_1435);
xor U1489 (N_1489,N_1429,N_1406);
nor U1490 (N_1490,N_1409,N_1407);
or U1491 (N_1491,N_1415,N_1428);
and U1492 (N_1492,N_1407,N_1440);
or U1493 (N_1493,N_1415,N_1400);
and U1494 (N_1494,N_1400,N_1425);
and U1495 (N_1495,N_1419,N_1420);
nand U1496 (N_1496,N_1443,N_1449);
nand U1497 (N_1497,N_1443,N_1413);
nor U1498 (N_1498,N_1420,N_1437);
nor U1499 (N_1499,N_1445,N_1405);
nand U1500 (N_1500,N_1468,N_1471);
nor U1501 (N_1501,N_1497,N_1477);
nand U1502 (N_1502,N_1452,N_1458);
or U1503 (N_1503,N_1464,N_1461);
nand U1504 (N_1504,N_1456,N_1476);
or U1505 (N_1505,N_1457,N_1475);
and U1506 (N_1506,N_1481,N_1491);
nand U1507 (N_1507,N_1480,N_1473);
xor U1508 (N_1508,N_1495,N_1492);
nor U1509 (N_1509,N_1472,N_1490);
and U1510 (N_1510,N_1493,N_1496);
or U1511 (N_1511,N_1488,N_1487);
xor U1512 (N_1512,N_1485,N_1489);
xor U1513 (N_1513,N_1463,N_1454);
nor U1514 (N_1514,N_1455,N_1467);
nor U1515 (N_1515,N_1474,N_1478);
nand U1516 (N_1516,N_1479,N_1459);
nor U1517 (N_1517,N_1470,N_1451);
or U1518 (N_1518,N_1465,N_1453);
and U1519 (N_1519,N_1483,N_1469);
nor U1520 (N_1520,N_1494,N_1466);
xor U1521 (N_1521,N_1486,N_1499);
xor U1522 (N_1522,N_1498,N_1450);
or U1523 (N_1523,N_1484,N_1460);
or U1524 (N_1524,N_1462,N_1482);
nand U1525 (N_1525,N_1460,N_1477);
xor U1526 (N_1526,N_1452,N_1488);
or U1527 (N_1527,N_1456,N_1464);
and U1528 (N_1528,N_1496,N_1469);
or U1529 (N_1529,N_1450,N_1456);
or U1530 (N_1530,N_1476,N_1497);
and U1531 (N_1531,N_1462,N_1456);
and U1532 (N_1532,N_1480,N_1472);
and U1533 (N_1533,N_1450,N_1451);
nand U1534 (N_1534,N_1471,N_1466);
xor U1535 (N_1535,N_1463,N_1493);
xor U1536 (N_1536,N_1463,N_1476);
xor U1537 (N_1537,N_1475,N_1487);
nor U1538 (N_1538,N_1461,N_1472);
nand U1539 (N_1539,N_1460,N_1466);
and U1540 (N_1540,N_1485,N_1466);
and U1541 (N_1541,N_1474,N_1466);
and U1542 (N_1542,N_1498,N_1495);
nand U1543 (N_1543,N_1493,N_1480);
xor U1544 (N_1544,N_1463,N_1488);
nand U1545 (N_1545,N_1475,N_1498);
nor U1546 (N_1546,N_1455,N_1463);
nor U1547 (N_1547,N_1450,N_1494);
or U1548 (N_1548,N_1469,N_1472);
and U1549 (N_1549,N_1491,N_1494);
nor U1550 (N_1550,N_1531,N_1517);
nand U1551 (N_1551,N_1547,N_1500);
and U1552 (N_1552,N_1524,N_1513);
and U1553 (N_1553,N_1521,N_1545);
nand U1554 (N_1554,N_1536,N_1532);
nand U1555 (N_1555,N_1523,N_1502);
nand U1556 (N_1556,N_1546,N_1549);
or U1557 (N_1557,N_1512,N_1520);
or U1558 (N_1558,N_1519,N_1526);
nor U1559 (N_1559,N_1505,N_1544);
or U1560 (N_1560,N_1516,N_1525);
nand U1561 (N_1561,N_1543,N_1535);
and U1562 (N_1562,N_1510,N_1538);
or U1563 (N_1563,N_1507,N_1530);
nand U1564 (N_1564,N_1548,N_1514);
nor U1565 (N_1565,N_1542,N_1533);
nand U1566 (N_1566,N_1515,N_1540);
nor U1567 (N_1567,N_1522,N_1509);
and U1568 (N_1568,N_1511,N_1534);
nor U1569 (N_1569,N_1527,N_1539);
and U1570 (N_1570,N_1508,N_1537);
nor U1571 (N_1571,N_1506,N_1528);
xor U1572 (N_1572,N_1529,N_1541);
or U1573 (N_1573,N_1503,N_1501);
xor U1574 (N_1574,N_1504,N_1518);
nor U1575 (N_1575,N_1541,N_1507);
or U1576 (N_1576,N_1541,N_1520);
and U1577 (N_1577,N_1538,N_1512);
nand U1578 (N_1578,N_1540,N_1530);
and U1579 (N_1579,N_1503,N_1520);
or U1580 (N_1580,N_1538,N_1528);
nand U1581 (N_1581,N_1535,N_1538);
nor U1582 (N_1582,N_1521,N_1520);
or U1583 (N_1583,N_1541,N_1535);
nand U1584 (N_1584,N_1518,N_1513);
nor U1585 (N_1585,N_1519,N_1538);
or U1586 (N_1586,N_1507,N_1548);
nand U1587 (N_1587,N_1531,N_1532);
or U1588 (N_1588,N_1527,N_1514);
or U1589 (N_1589,N_1535,N_1530);
nor U1590 (N_1590,N_1538,N_1532);
or U1591 (N_1591,N_1528,N_1511);
and U1592 (N_1592,N_1529,N_1527);
nor U1593 (N_1593,N_1506,N_1532);
nor U1594 (N_1594,N_1534,N_1535);
nand U1595 (N_1595,N_1523,N_1514);
and U1596 (N_1596,N_1503,N_1543);
xnor U1597 (N_1597,N_1539,N_1547);
or U1598 (N_1598,N_1511,N_1531);
or U1599 (N_1599,N_1524,N_1543);
and U1600 (N_1600,N_1596,N_1593);
nor U1601 (N_1601,N_1592,N_1569);
nand U1602 (N_1602,N_1591,N_1572);
nor U1603 (N_1603,N_1568,N_1574);
nand U1604 (N_1604,N_1579,N_1594);
xor U1605 (N_1605,N_1578,N_1581);
or U1606 (N_1606,N_1563,N_1550);
or U1607 (N_1607,N_1558,N_1555);
nand U1608 (N_1608,N_1571,N_1587);
or U1609 (N_1609,N_1580,N_1595);
xnor U1610 (N_1610,N_1590,N_1561);
and U1611 (N_1611,N_1564,N_1585);
or U1612 (N_1612,N_1566,N_1575);
nand U1613 (N_1613,N_1562,N_1583);
nand U1614 (N_1614,N_1573,N_1565);
nand U1615 (N_1615,N_1588,N_1567);
nor U1616 (N_1616,N_1570,N_1551);
and U1617 (N_1617,N_1576,N_1553);
nor U1618 (N_1618,N_1556,N_1554);
and U1619 (N_1619,N_1589,N_1552);
or U1620 (N_1620,N_1598,N_1557);
or U1621 (N_1621,N_1577,N_1586);
and U1622 (N_1622,N_1597,N_1599);
nand U1623 (N_1623,N_1582,N_1584);
or U1624 (N_1624,N_1559,N_1560);
or U1625 (N_1625,N_1575,N_1578);
nor U1626 (N_1626,N_1593,N_1566);
or U1627 (N_1627,N_1578,N_1592);
or U1628 (N_1628,N_1561,N_1592);
nor U1629 (N_1629,N_1559,N_1573);
nor U1630 (N_1630,N_1563,N_1565);
nor U1631 (N_1631,N_1554,N_1561);
nand U1632 (N_1632,N_1584,N_1557);
or U1633 (N_1633,N_1572,N_1558);
nand U1634 (N_1634,N_1581,N_1552);
and U1635 (N_1635,N_1596,N_1566);
or U1636 (N_1636,N_1586,N_1599);
xor U1637 (N_1637,N_1557,N_1553);
xnor U1638 (N_1638,N_1595,N_1568);
nand U1639 (N_1639,N_1587,N_1560);
nor U1640 (N_1640,N_1565,N_1550);
nor U1641 (N_1641,N_1550,N_1564);
or U1642 (N_1642,N_1555,N_1553);
or U1643 (N_1643,N_1556,N_1575);
nand U1644 (N_1644,N_1592,N_1577);
or U1645 (N_1645,N_1555,N_1571);
xnor U1646 (N_1646,N_1557,N_1550);
or U1647 (N_1647,N_1561,N_1553);
xnor U1648 (N_1648,N_1591,N_1569);
or U1649 (N_1649,N_1555,N_1585);
nor U1650 (N_1650,N_1644,N_1647);
nand U1651 (N_1651,N_1643,N_1646);
or U1652 (N_1652,N_1639,N_1635);
or U1653 (N_1653,N_1613,N_1638);
or U1654 (N_1654,N_1617,N_1632);
and U1655 (N_1655,N_1600,N_1619);
nor U1656 (N_1656,N_1618,N_1641);
or U1657 (N_1657,N_1604,N_1620);
or U1658 (N_1658,N_1616,N_1607);
and U1659 (N_1659,N_1623,N_1609);
or U1660 (N_1660,N_1608,N_1649);
nand U1661 (N_1661,N_1636,N_1602);
nand U1662 (N_1662,N_1630,N_1605);
or U1663 (N_1663,N_1603,N_1640);
nor U1664 (N_1664,N_1634,N_1648);
nor U1665 (N_1665,N_1601,N_1628);
nand U1666 (N_1666,N_1631,N_1633);
nor U1667 (N_1667,N_1614,N_1626);
xnor U1668 (N_1668,N_1611,N_1624);
or U1669 (N_1669,N_1606,N_1629);
nor U1670 (N_1670,N_1637,N_1621);
nand U1671 (N_1671,N_1612,N_1625);
nand U1672 (N_1672,N_1610,N_1642);
or U1673 (N_1673,N_1615,N_1622);
or U1674 (N_1674,N_1645,N_1627);
or U1675 (N_1675,N_1607,N_1615);
nor U1676 (N_1676,N_1608,N_1604);
xnor U1677 (N_1677,N_1607,N_1632);
xnor U1678 (N_1678,N_1605,N_1637);
and U1679 (N_1679,N_1623,N_1614);
nor U1680 (N_1680,N_1648,N_1617);
and U1681 (N_1681,N_1642,N_1614);
or U1682 (N_1682,N_1641,N_1605);
nand U1683 (N_1683,N_1606,N_1625);
and U1684 (N_1684,N_1648,N_1606);
or U1685 (N_1685,N_1631,N_1635);
or U1686 (N_1686,N_1614,N_1647);
nand U1687 (N_1687,N_1626,N_1640);
nor U1688 (N_1688,N_1603,N_1628);
or U1689 (N_1689,N_1640,N_1642);
and U1690 (N_1690,N_1621,N_1605);
and U1691 (N_1691,N_1624,N_1643);
nand U1692 (N_1692,N_1644,N_1612);
nand U1693 (N_1693,N_1646,N_1647);
nor U1694 (N_1694,N_1628,N_1627);
or U1695 (N_1695,N_1601,N_1646);
and U1696 (N_1696,N_1605,N_1638);
xnor U1697 (N_1697,N_1615,N_1611);
nor U1698 (N_1698,N_1611,N_1633);
nand U1699 (N_1699,N_1606,N_1626);
or U1700 (N_1700,N_1683,N_1674);
and U1701 (N_1701,N_1652,N_1654);
and U1702 (N_1702,N_1662,N_1677);
xnor U1703 (N_1703,N_1681,N_1696);
nand U1704 (N_1704,N_1673,N_1680);
xnor U1705 (N_1705,N_1661,N_1651);
and U1706 (N_1706,N_1664,N_1655);
nand U1707 (N_1707,N_1689,N_1675);
or U1708 (N_1708,N_1659,N_1698);
and U1709 (N_1709,N_1693,N_1685);
nand U1710 (N_1710,N_1690,N_1665);
nor U1711 (N_1711,N_1684,N_1686);
nor U1712 (N_1712,N_1691,N_1697);
xor U1713 (N_1713,N_1688,N_1667);
nand U1714 (N_1714,N_1671,N_1687);
xnor U1715 (N_1715,N_1672,N_1670);
and U1716 (N_1716,N_1695,N_1657);
or U1717 (N_1717,N_1653,N_1676);
xnor U1718 (N_1718,N_1682,N_1669);
nand U1719 (N_1719,N_1666,N_1679);
nand U1720 (N_1720,N_1692,N_1663);
nand U1721 (N_1721,N_1699,N_1660);
nand U1722 (N_1722,N_1656,N_1668);
or U1723 (N_1723,N_1678,N_1694);
or U1724 (N_1724,N_1658,N_1650);
and U1725 (N_1725,N_1688,N_1693);
and U1726 (N_1726,N_1693,N_1668);
or U1727 (N_1727,N_1682,N_1675);
nand U1728 (N_1728,N_1664,N_1650);
nor U1729 (N_1729,N_1655,N_1674);
or U1730 (N_1730,N_1665,N_1669);
or U1731 (N_1731,N_1656,N_1655);
nor U1732 (N_1732,N_1654,N_1694);
or U1733 (N_1733,N_1680,N_1686);
xnor U1734 (N_1734,N_1674,N_1681);
xor U1735 (N_1735,N_1689,N_1695);
or U1736 (N_1736,N_1677,N_1681);
or U1737 (N_1737,N_1678,N_1672);
or U1738 (N_1738,N_1687,N_1676);
and U1739 (N_1739,N_1694,N_1664);
or U1740 (N_1740,N_1654,N_1685);
nor U1741 (N_1741,N_1673,N_1698);
nor U1742 (N_1742,N_1676,N_1699);
or U1743 (N_1743,N_1665,N_1675);
or U1744 (N_1744,N_1673,N_1653);
nor U1745 (N_1745,N_1688,N_1677);
nor U1746 (N_1746,N_1691,N_1666);
xnor U1747 (N_1747,N_1655,N_1695);
xor U1748 (N_1748,N_1650,N_1695);
nand U1749 (N_1749,N_1662,N_1683);
and U1750 (N_1750,N_1707,N_1710);
or U1751 (N_1751,N_1702,N_1726);
nand U1752 (N_1752,N_1706,N_1738);
nand U1753 (N_1753,N_1746,N_1708);
nor U1754 (N_1754,N_1720,N_1714);
or U1755 (N_1755,N_1709,N_1722);
nor U1756 (N_1756,N_1716,N_1705);
nand U1757 (N_1757,N_1723,N_1739);
nand U1758 (N_1758,N_1711,N_1740);
xor U1759 (N_1759,N_1743,N_1730);
nor U1760 (N_1760,N_1704,N_1747);
and U1761 (N_1761,N_1748,N_1734);
nor U1762 (N_1762,N_1724,N_1719);
and U1763 (N_1763,N_1735,N_1731);
or U1764 (N_1764,N_1745,N_1727);
or U1765 (N_1765,N_1736,N_1725);
and U1766 (N_1766,N_1733,N_1718);
nor U1767 (N_1767,N_1744,N_1742);
and U1768 (N_1768,N_1715,N_1703);
nand U1769 (N_1769,N_1737,N_1713);
or U1770 (N_1770,N_1717,N_1728);
nor U1771 (N_1771,N_1749,N_1712);
nand U1772 (N_1772,N_1732,N_1701);
nor U1773 (N_1773,N_1741,N_1721);
or U1774 (N_1774,N_1729,N_1700);
nand U1775 (N_1775,N_1740,N_1713);
nand U1776 (N_1776,N_1713,N_1708);
or U1777 (N_1777,N_1744,N_1724);
and U1778 (N_1778,N_1733,N_1702);
or U1779 (N_1779,N_1704,N_1706);
or U1780 (N_1780,N_1742,N_1733);
nand U1781 (N_1781,N_1701,N_1734);
xnor U1782 (N_1782,N_1743,N_1727);
and U1783 (N_1783,N_1709,N_1705);
and U1784 (N_1784,N_1737,N_1731);
nand U1785 (N_1785,N_1726,N_1724);
nor U1786 (N_1786,N_1737,N_1720);
xnor U1787 (N_1787,N_1737,N_1732);
nor U1788 (N_1788,N_1709,N_1720);
and U1789 (N_1789,N_1749,N_1731);
nand U1790 (N_1790,N_1734,N_1730);
nand U1791 (N_1791,N_1732,N_1743);
and U1792 (N_1792,N_1736,N_1708);
nor U1793 (N_1793,N_1728,N_1742);
xor U1794 (N_1794,N_1736,N_1714);
xor U1795 (N_1795,N_1746,N_1715);
xnor U1796 (N_1796,N_1709,N_1726);
xnor U1797 (N_1797,N_1719,N_1733);
or U1798 (N_1798,N_1747,N_1716);
nand U1799 (N_1799,N_1719,N_1749);
xor U1800 (N_1800,N_1789,N_1783);
nor U1801 (N_1801,N_1759,N_1798);
nor U1802 (N_1802,N_1782,N_1784);
and U1803 (N_1803,N_1750,N_1754);
nor U1804 (N_1804,N_1758,N_1792);
and U1805 (N_1805,N_1767,N_1778);
nor U1806 (N_1806,N_1771,N_1772);
nor U1807 (N_1807,N_1756,N_1774);
nor U1808 (N_1808,N_1777,N_1799);
and U1809 (N_1809,N_1790,N_1766);
nor U1810 (N_1810,N_1795,N_1768);
nor U1811 (N_1811,N_1781,N_1787);
nand U1812 (N_1812,N_1765,N_1776);
nand U1813 (N_1813,N_1757,N_1764);
and U1814 (N_1814,N_1780,N_1753);
nor U1815 (N_1815,N_1791,N_1793);
and U1816 (N_1816,N_1763,N_1761);
or U1817 (N_1817,N_1796,N_1770);
or U1818 (N_1818,N_1794,N_1760);
xnor U1819 (N_1819,N_1786,N_1752);
or U1820 (N_1820,N_1755,N_1769);
and U1821 (N_1821,N_1751,N_1788);
and U1822 (N_1822,N_1762,N_1797);
and U1823 (N_1823,N_1775,N_1785);
and U1824 (N_1824,N_1779,N_1773);
or U1825 (N_1825,N_1759,N_1776);
or U1826 (N_1826,N_1765,N_1798);
xor U1827 (N_1827,N_1770,N_1771);
and U1828 (N_1828,N_1752,N_1758);
and U1829 (N_1829,N_1756,N_1762);
nor U1830 (N_1830,N_1769,N_1775);
nor U1831 (N_1831,N_1789,N_1795);
nor U1832 (N_1832,N_1799,N_1784);
nor U1833 (N_1833,N_1758,N_1788);
nand U1834 (N_1834,N_1751,N_1765);
and U1835 (N_1835,N_1764,N_1752);
and U1836 (N_1836,N_1752,N_1780);
or U1837 (N_1837,N_1795,N_1757);
xor U1838 (N_1838,N_1762,N_1776);
or U1839 (N_1839,N_1765,N_1771);
and U1840 (N_1840,N_1765,N_1775);
nand U1841 (N_1841,N_1753,N_1754);
nor U1842 (N_1842,N_1778,N_1755);
nor U1843 (N_1843,N_1797,N_1795);
nand U1844 (N_1844,N_1783,N_1796);
xor U1845 (N_1845,N_1796,N_1788);
and U1846 (N_1846,N_1794,N_1755);
and U1847 (N_1847,N_1768,N_1798);
and U1848 (N_1848,N_1753,N_1750);
nor U1849 (N_1849,N_1750,N_1776);
and U1850 (N_1850,N_1831,N_1826);
and U1851 (N_1851,N_1810,N_1802);
nand U1852 (N_1852,N_1822,N_1848);
nor U1853 (N_1853,N_1806,N_1815);
and U1854 (N_1854,N_1829,N_1800);
xnor U1855 (N_1855,N_1845,N_1842);
nand U1856 (N_1856,N_1837,N_1817);
nand U1857 (N_1857,N_1834,N_1841);
nand U1858 (N_1858,N_1819,N_1813);
nand U1859 (N_1859,N_1816,N_1830);
nor U1860 (N_1860,N_1832,N_1812);
nand U1861 (N_1861,N_1828,N_1808);
or U1862 (N_1862,N_1805,N_1839);
nand U1863 (N_1863,N_1847,N_1821);
xor U1864 (N_1864,N_1820,N_1838);
nand U1865 (N_1865,N_1803,N_1849);
or U1866 (N_1866,N_1843,N_1824);
and U1867 (N_1867,N_1801,N_1823);
and U1868 (N_1868,N_1833,N_1840);
xnor U1869 (N_1869,N_1836,N_1825);
nand U1870 (N_1870,N_1835,N_1844);
and U1871 (N_1871,N_1818,N_1827);
or U1872 (N_1872,N_1814,N_1807);
nor U1873 (N_1873,N_1811,N_1846);
or U1874 (N_1874,N_1809,N_1804);
or U1875 (N_1875,N_1803,N_1848);
or U1876 (N_1876,N_1830,N_1809);
and U1877 (N_1877,N_1829,N_1835);
xor U1878 (N_1878,N_1810,N_1818);
nor U1879 (N_1879,N_1822,N_1847);
nand U1880 (N_1880,N_1826,N_1833);
xor U1881 (N_1881,N_1808,N_1818);
nor U1882 (N_1882,N_1809,N_1829);
and U1883 (N_1883,N_1814,N_1816);
and U1884 (N_1884,N_1805,N_1822);
nand U1885 (N_1885,N_1807,N_1844);
nand U1886 (N_1886,N_1841,N_1808);
xor U1887 (N_1887,N_1847,N_1824);
and U1888 (N_1888,N_1815,N_1809);
or U1889 (N_1889,N_1843,N_1834);
or U1890 (N_1890,N_1813,N_1803);
or U1891 (N_1891,N_1845,N_1841);
nor U1892 (N_1892,N_1840,N_1834);
nand U1893 (N_1893,N_1837,N_1831);
or U1894 (N_1894,N_1837,N_1814);
nand U1895 (N_1895,N_1803,N_1819);
and U1896 (N_1896,N_1800,N_1807);
nand U1897 (N_1897,N_1840,N_1810);
nand U1898 (N_1898,N_1815,N_1804);
or U1899 (N_1899,N_1840,N_1807);
xnor U1900 (N_1900,N_1873,N_1878);
nor U1901 (N_1901,N_1899,N_1863);
nand U1902 (N_1902,N_1880,N_1897);
nand U1903 (N_1903,N_1891,N_1870);
nor U1904 (N_1904,N_1898,N_1883);
and U1905 (N_1905,N_1862,N_1851);
or U1906 (N_1906,N_1890,N_1857);
or U1907 (N_1907,N_1858,N_1855);
or U1908 (N_1908,N_1872,N_1894);
xnor U1909 (N_1909,N_1867,N_1874);
and U1910 (N_1910,N_1860,N_1884);
or U1911 (N_1911,N_1889,N_1856);
nand U1912 (N_1912,N_1881,N_1859);
nand U1913 (N_1913,N_1854,N_1875);
and U1914 (N_1914,N_1868,N_1886);
xor U1915 (N_1915,N_1895,N_1866);
and U1916 (N_1916,N_1871,N_1876);
or U1917 (N_1917,N_1864,N_1887);
nand U1918 (N_1918,N_1861,N_1852);
and U1919 (N_1919,N_1896,N_1882);
xor U1920 (N_1920,N_1879,N_1865);
and U1921 (N_1921,N_1885,N_1892);
and U1922 (N_1922,N_1888,N_1877);
and U1923 (N_1923,N_1893,N_1869);
nor U1924 (N_1924,N_1850,N_1853);
xnor U1925 (N_1925,N_1886,N_1888);
nand U1926 (N_1926,N_1884,N_1858);
or U1927 (N_1927,N_1896,N_1883);
nand U1928 (N_1928,N_1888,N_1885);
and U1929 (N_1929,N_1852,N_1896);
or U1930 (N_1930,N_1877,N_1872);
nand U1931 (N_1931,N_1895,N_1879);
nor U1932 (N_1932,N_1850,N_1862);
nor U1933 (N_1933,N_1889,N_1870);
and U1934 (N_1934,N_1882,N_1869);
nand U1935 (N_1935,N_1855,N_1872);
or U1936 (N_1936,N_1887,N_1872);
and U1937 (N_1937,N_1886,N_1860);
nor U1938 (N_1938,N_1897,N_1871);
xnor U1939 (N_1939,N_1875,N_1881);
and U1940 (N_1940,N_1887,N_1883);
or U1941 (N_1941,N_1884,N_1889);
and U1942 (N_1942,N_1868,N_1860);
nand U1943 (N_1943,N_1899,N_1889);
and U1944 (N_1944,N_1888,N_1874);
nand U1945 (N_1945,N_1850,N_1851);
and U1946 (N_1946,N_1879,N_1891);
nand U1947 (N_1947,N_1883,N_1875);
xnor U1948 (N_1948,N_1885,N_1893);
or U1949 (N_1949,N_1896,N_1899);
and U1950 (N_1950,N_1948,N_1901);
and U1951 (N_1951,N_1914,N_1920);
or U1952 (N_1952,N_1910,N_1922);
and U1953 (N_1953,N_1930,N_1949);
or U1954 (N_1954,N_1931,N_1919);
nor U1955 (N_1955,N_1928,N_1926);
and U1956 (N_1956,N_1904,N_1916);
and U1957 (N_1957,N_1902,N_1900);
and U1958 (N_1958,N_1929,N_1912);
nor U1959 (N_1959,N_1946,N_1938);
and U1960 (N_1960,N_1918,N_1943);
and U1961 (N_1961,N_1939,N_1944);
or U1962 (N_1962,N_1924,N_1925);
or U1963 (N_1963,N_1940,N_1936);
nand U1964 (N_1964,N_1915,N_1903);
nor U1965 (N_1965,N_1927,N_1905);
nor U1966 (N_1966,N_1913,N_1909);
nor U1967 (N_1967,N_1947,N_1906);
and U1968 (N_1968,N_1935,N_1908);
nand U1969 (N_1969,N_1921,N_1923);
and U1970 (N_1970,N_1933,N_1917);
or U1971 (N_1971,N_1907,N_1934);
or U1972 (N_1972,N_1945,N_1942);
and U1973 (N_1973,N_1937,N_1932);
and U1974 (N_1974,N_1941,N_1911);
and U1975 (N_1975,N_1918,N_1949);
and U1976 (N_1976,N_1917,N_1910);
nor U1977 (N_1977,N_1934,N_1915);
and U1978 (N_1978,N_1911,N_1949);
nand U1979 (N_1979,N_1921,N_1901);
and U1980 (N_1980,N_1932,N_1948);
or U1981 (N_1981,N_1903,N_1914);
nand U1982 (N_1982,N_1915,N_1932);
nand U1983 (N_1983,N_1925,N_1913);
xnor U1984 (N_1984,N_1946,N_1940);
or U1985 (N_1985,N_1918,N_1907);
nor U1986 (N_1986,N_1945,N_1913);
nor U1987 (N_1987,N_1943,N_1948);
and U1988 (N_1988,N_1944,N_1949);
nor U1989 (N_1989,N_1941,N_1910);
nand U1990 (N_1990,N_1906,N_1907);
or U1991 (N_1991,N_1935,N_1945);
nor U1992 (N_1992,N_1934,N_1921);
nand U1993 (N_1993,N_1946,N_1900);
nand U1994 (N_1994,N_1920,N_1929);
or U1995 (N_1995,N_1945,N_1924);
nor U1996 (N_1996,N_1916,N_1933);
xor U1997 (N_1997,N_1938,N_1934);
and U1998 (N_1998,N_1935,N_1901);
xnor U1999 (N_1999,N_1928,N_1921);
or U2000 (N_2000,N_1980,N_1992);
nor U2001 (N_2001,N_1996,N_1963);
nand U2002 (N_2002,N_1972,N_1984);
nor U2003 (N_2003,N_1969,N_1970);
nor U2004 (N_2004,N_1994,N_1950);
nor U2005 (N_2005,N_1986,N_1967);
nor U2006 (N_2006,N_1957,N_1958);
and U2007 (N_2007,N_1993,N_1978);
nor U2008 (N_2008,N_1962,N_1965);
or U2009 (N_2009,N_1985,N_1988);
xnor U2010 (N_2010,N_1977,N_1998);
or U2011 (N_2011,N_1954,N_1971);
nor U2012 (N_2012,N_1976,N_1951);
nand U2013 (N_2013,N_1973,N_1953);
and U2014 (N_2014,N_1952,N_1960);
nor U2015 (N_2015,N_1982,N_1981);
nor U2016 (N_2016,N_1975,N_1990);
xnor U2017 (N_2017,N_1983,N_1955);
or U2018 (N_2018,N_1997,N_1956);
nand U2019 (N_2019,N_1964,N_1995);
nor U2020 (N_2020,N_1989,N_1961);
nand U2021 (N_2021,N_1987,N_1999);
nor U2022 (N_2022,N_1974,N_1959);
and U2023 (N_2023,N_1966,N_1968);
and U2024 (N_2024,N_1979,N_1991);
nand U2025 (N_2025,N_1967,N_1987);
xor U2026 (N_2026,N_1996,N_1990);
nor U2027 (N_2027,N_1977,N_1990);
and U2028 (N_2028,N_1954,N_1961);
or U2029 (N_2029,N_1973,N_1970);
nand U2030 (N_2030,N_1968,N_1961);
nor U2031 (N_2031,N_1953,N_1951);
or U2032 (N_2032,N_1981,N_1953);
nand U2033 (N_2033,N_1957,N_1998);
nor U2034 (N_2034,N_1951,N_1981);
nor U2035 (N_2035,N_1995,N_1959);
nor U2036 (N_2036,N_1978,N_1987);
or U2037 (N_2037,N_1990,N_1966);
or U2038 (N_2038,N_1954,N_1963);
xnor U2039 (N_2039,N_1984,N_1956);
nand U2040 (N_2040,N_1980,N_1964);
and U2041 (N_2041,N_1981,N_1993);
nand U2042 (N_2042,N_1989,N_1980);
nor U2043 (N_2043,N_1961,N_1979);
nand U2044 (N_2044,N_1958,N_1997);
nor U2045 (N_2045,N_1998,N_1967);
nor U2046 (N_2046,N_1974,N_1992);
xnor U2047 (N_2047,N_1961,N_1964);
and U2048 (N_2048,N_1978,N_1954);
or U2049 (N_2049,N_1987,N_1961);
nand U2050 (N_2050,N_2031,N_2034);
nand U2051 (N_2051,N_2045,N_2023);
xor U2052 (N_2052,N_2008,N_2015);
nor U2053 (N_2053,N_2021,N_2044);
or U2054 (N_2054,N_2014,N_2001);
nor U2055 (N_2055,N_2022,N_2027);
xor U2056 (N_2056,N_2004,N_2037);
nand U2057 (N_2057,N_2010,N_2043);
nor U2058 (N_2058,N_2035,N_2042);
or U2059 (N_2059,N_2017,N_2013);
and U2060 (N_2060,N_2046,N_2003);
and U2061 (N_2061,N_2047,N_2040);
nand U2062 (N_2062,N_2029,N_2018);
nor U2063 (N_2063,N_2048,N_2024);
or U2064 (N_2064,N_2025,N_2011);
nor U2065 (N_2065,N_2007,N_2020);
and U2066 (N_2066,N_2000,N_2028);
xor U2067 (N_2067,N_2016,N_2030);
or U2068 (N_2068,N_2049,N_2041);
nor U2069 (N_2069,N_2002,N_2032);
nand U2070 (N_2070,N_2039,N_2005);
and U2071 (N_2071,N_2036,N_2019);
xnor U2072 (N_2072,N_2009,N_2038);
nand U2073 (N_2073,N_2012,N_2033);
or U2074 (N_2074,N_2006,N_2026);
nand U2075 (N_2075,N_2012,N_2029);
and U2076 (N_2076,N_2039,N_2044);
nand U2077 (N_2077,N_2029,N_2004);
nor U2078 (N_2078,N_2011,N_2017);
or U2079 (N_2079,N_2038,N_2003);
or U2080 (N_2080,N_2011,N_2030);
and U2081 (N_2081,N_2004,N_2000);
nand U2082 (N_2082,N_2025,N_2031);
xnor U2083 (N_2083,N_2012,N_2037);
nor U2084 (N_2084,N_2027,N_2020);
nand U2085 (N_2085,N_2024,N_2017);
or U2086 (N_2086,N_2022,N_2005);
or U2087 (N_2087,N_2044,N_2011);
nand U2088 (N_2088,N_2046,N_2024);
xor U2089 (N_2089,N_2044,N_2015);
nor U2090 (N_2090,N_2019,N_2013);
and U2091 (N_2091,N_2033,N_2007);
and U2092 (N_2092,N_2018,N_2031);
nor U2093 (N_2093,N_2015,N_2009);
nor U2094 (N_2094,N_2005,N_2026);
or U2095 (N_2095,N_2018,N_2045);
and U2096 (N_2096,N_2006,N_2030);
xor U2097 (N_2097,N_2049,N_2044);
or U2098 (N_2098,N_2003,N_2035);
nor U2099 (N_2099,N_2000,N_2021);
nor U2100 (N_2100,N_2050,N_2052);
and U2101 (N_2101,N_2053,N_2096);
nand U2102 (N_2102,N_2061,N_2064);
nor U2103 (N_2103,N_2057,N_2083);
nor U2104 (N_2104,N_2062,N_2084);
nor U2105 (N_2105,N_2054,N_2081);
nand U2106 (N_2106,N_2051,N_2065);
and U2107 (N_2107,N_2093,N_2069);
nor U2108 (N_2108,N_2079,N_2070);
nand U2109 (N_2109,N_2092,N_2072);
nor U2110 (N_2110,N_2056,N_2059);
nor U2111 (N_2111,N_2071,N_2067);
and U2112 (N_2112,N_2097,N_2076);
xnor U2113 (N_2113,N_2073,N_2085);
or U2114 (N_2114,N_2094,N_2090);
and U2115 (N_2115,N_2080,N_2098);
nor U2116 (N_2116,N_2066,N_2074);
nand U2117 (N_2117,N_2078,N_2060);
nand U2118 (N_2118,N_2055,N_2091);
xor U2119 (N_2119,N_2087,N_2086);
nor U2120 (N_2120,N_2068,N_2077);
nor U2121 (N_2121,N_2089,N_2095);
and U2122 (N_2122,N_2082,N_2088);
nand U2123 (N_2123,N_2063,N_2075);
nand U2124 (N_2124,N_2058,N_2099);
nor U2125 (N_2125,N_2070,N_2072);
and U2126 (N_2126,N_2052,N_2084);
and U2127 (N_2127,N_2059,N_2090);
xnor U2128 (N_2128,N_2058,N_2053);
and U2129 (N_2129,N_2056,N_2050);
and U2130 (N_2130,N_2071,N_2063);
or U2131 (N_2131,N_2061,N_2074);
and U2132 (N_2132,N_2069,N_2094);
nor U2133 (N_2133,N_2096,N_2089);
and U2134 (N_2134,N_2055,N_2083);
nand U2135 (N_2135,N_2081,N_2075);
or U2136 (N_2136,N_2081,N_2058);
xnor U2137 (N_2137,N_2059,N_2092);
nor U2138 (N_2138,N_2071,N_2069);
nor U2139 (N_2139,N_2058,N_2051);
or U2140 (N_2140,N_2060,N_2097);
nor U2141 (N_2141,N_2076,N_2066);
and U2142 (N_2142,N_2064,N_2071);
nand U2143 (N_2143,N_2052,N_2057);
and U2144 (N_2144,N_2070,N_2094);
nor U2145 (N_2145,N_2058,N_2062);
or U2146 (N_2146,N_2051,N_2080);
xnor U2147 (N_2147,N_2052,N_2056);
nor U2148 (N_2148,N_2091,N_2061);
or U2149 (N_2149,N_2062,N_2053);
nor U2150 (N_2150,N_2125,N_2136);
nor U2151 (N_2151,N_2115,N_2123);
nand U2152 (N_2152,N_2107,N_2147);
nand U2153 (N_2153,N_2146,N_2100);
nand U2154 (N_2154,N_2126,N_2114);
and U2155 (N_2155,N_2149,N_2145);
or U2156 (N_2156,N_2130,N_2119);
nor U2157 (N_2157,N_2122,N_2121);
nor U2158 (N_2158,N_2148,N_2134);
or U2159 (N_2159,N_2132,N_2108);
and U2160 (N_2160,N_2137,N_2112);
and U2161 (N_2161,N_2139,N_2111);
nand U2162 (N_2162,N_2120,N_2128);
nor U2163 (N_2163,N_2110,N_2129);
or U2164 (N_2164,N_2106,N_2109);
xor U2165 (N_2165,N_2143,N_2144);
and U2166 (N_2166,N_2131,N_2105);
and U2167 (N_2167,N_2141,N_2124);
or U2168 (N_2168,N_2142,N_2127);
nand U2169 (N_2169,N_2102,N_2116);
nor U2170 (N_2170,N_2101,N_2133);
nand U2171 (N_2171,N_2103,N_2140);
nand U2172 (N_2172,N_2118,N_2138);
and U2173 (N_2173,N_2117,N_2135);
nor U2174 (N_2174,N_2104,N_2113);
or U2175 (N_2175,N_2143,N_2127);
nand U2176 (N_2176,N_2132,N_2145);
nand U2177 (N_2177,N_2142,N_2117);
xnor U2178 (N_2178,N_2112,N_2108);
nand U2179 (N_2179,N_2114,N_2147);
and U2180 (N_2180,N_2136,N_2143);
nor U2181 (N_2181,N_2111,N_2101);
and U2182 (N_2182,N_2126,N_2117);
or U2183 (N_2183,N_2111,N_2102);
and U2184 (N_2184,N_2130,N_2148);
nand U2185 (N_2185,N_2143,N_2149);
and U2186 (N_2186,N_2138,N_2134);
nor U2187 (N_2187,N_2142,N_2121);
nand U2188 (N_2188,N_2147,N_2122);
or U2189 (N_2189,N_2111,N_2109);
nand U2190 (N_2190,N_2108,N_2139);
nor U2191 (N_2191,N_2140,N_2106);
nor U2192 (N_2192,N_2140,N_2112);
nand U2193 (N_2193,N_2102,N_2104);
nand U2194 (N_2194,N_2115,N_2132);
and U2195 (N_2195,N_2134,N_2110);
nor U2196 (N_2196,N_2148,N_2143);
xor U2197 (N_2197,N_2127,N_2122);
or U2198 (N_2198,N_2146,N_2116);
nand U2199 (N_2199,N_2118,N_2113);
nand U2200 (N_2200,N_2193,N_2172);
and U2201 (N_2201,N_2192,N_2157);
nor U2202 (N_2202,N_2158,N_2150);
nand U2203 (N_2203,N_2155,N_2161);
nor U2204 (N_2204,N_2183,N_2188);
or U2205 (N_2205,N_2175,N_2167);
nor U2206 (N_2206,N_2154,N_2180);
xnor U2207 (N_2207,N_2198,N_2156);
or U2208 (N_2208,N_2151,N_2165);
or U2209 (N_2209,N_2181,N_2166);
nand U2210 (N_2210,N_2194,N_2162);
nand U2211 (N_2211,N_2152,N_2174);
nor U2212 (N_2212,N_2163,N_2168);
or U2213 (N_2213,N_2169,N_2186);
or U2214 (N_2214,N_2179,N_2191);
or U2215 (N_2215,N_2189,N_2196);
nor U2216 (N_2216,N_2199,N_2195);
nand U2217 (N_2217,N_2187,N_2173);
nor U2218 (N_2218,N_2185,N_2176);
xor U2219 (N_2219,N_2164,N_2177);
xnor U2220 (N_2220,N_2182,N_2190);
xor U2221 (N_2221,N_2159,N_2178);
nor U2222 (N_2222,N_2170,N_2153);
nor U2223 (N_2223,N_2197,N_2171);
and U2224 (N_2224,N_2160,N_2184);
and U2225 (N_2225,N_2153,N_2181);
nand U2226 (N_2226,N_2171,N_2152);
and U2227 (N_2227,N_2190,N_2194);
nor U2228 (N_2228,N_2161,N_2174);
nand U2229 (N_2229,N_2173,N_2190);
nand U2230 (N_2230,N_2189,N_2177);
and U2231 (N_2231,N_2153,N_2184);
or U2232 (N_2232,N_2163,N_2171);
and U2233 (N_2233,N_2191,N_2198);
and U2234 (N_2234,N_2168,N_2169);
and U2235 (N_2235,N_2191,N_2195);
nand U2236 (N_2236,N_2198,N_2189);
nor U2237 (N_2237,N_2154,N_2181);
nor U2238 (N_2238,N_2187,N_2185);
or U2239 (N_2239,N_2156,N_2184);
xnor U2240 (N_2240,N_2159,N_2179);
nand U2241 (N_2241,N_2190,N_2185);
and U2242 (N_2242,N_2168,N_2178);
xor U2243 (N_2243,N_2192,N_2180);
and U2244 (N_2244,N_2186,N_2184);
xor U2245 (N_2245,N_2194,N_2172);
or U2246 (N_2246,N_2163,N_2151);
nand U2247 (N_2247,N_2187,N_2157);
or U2248 (N_2248,N_2151,N_2190);
nand U2249 (N_2249,N_2190,N_2174);
nand U2250 (N_2250,N_2212,N_2232);
and U2251 (N_2251,N_2242,N_2226);
or U2252 (N_2252,N_2211,N_2248);
or U2253 (N_2253,N_2204,N_2233);
nor U2254 (N_2254,N_2216,N_2206);
and U2255 (N_2255,N_2202,N_2225);
nand U2256 (N_2256,N_2231,N_2240);
xor U2257 (N_2257,N_2222,N_2229);
xor U2258 (N_2258,N_2220,N_2228);
or U2259 (N_2259,N_2238,N_2236);
nand U2260 (N_2260,N_2223,N_2210);
nor U2261 (N_2261,N_2208,N_2217);
nand U2262 (N_2262,N_2203,N_2246);
or U2263 (N_2263,N_2218,N_2221);
nand U2264 (N_2264,N_2205,N_2200);
xnor U2265 (N_2265,N_2213,N_2237);
xnor U2266 (N_2266,N_2230,N_2239);
nand U2267 (N_2267,N_2241,N_2245);
nor U2268 (N_2268,N_2215,N_2227);
or U2269 (N_2269,N_2234,N_2244);
nor U2270 (N_2270,N_2219,N_2243);
or U2271 (N_2271,N_2235,N_2249);
nand U2272 (N_2272,N_2214,N_2247);
nand U2273 (N_2273,N_2201,N_2224);
and U2274 (N_2274,N_2209,N_2207);
xnor U2275 (N_2275,N_2237,N_2203);
nand U2276 (N_2276,N_2213,N_2239);
nor U2277 (N_2277,N_2207,N_2227);
nor U2278 (N_2278,N_2232,N_2207);
or U2279 (N_2279,N_2204,N_2210);
nor U2280 (N_2280,N_2232,N_2248);
nand U2281 (N_2281,N_2245,N_2243);
nand U2282 (N_2282,N_2226,N_2245);
or U2283 (N_2283,N_2218,N_2246);
nor U2284 (N_2284,N_2203,N_2209);
nor U2285 (N_2285,N_2228,N_2219);
or U2286 (N_2286,N_2230,N_2232);
nand U2287 (N_2287,N_2224,N_2210);
nand U2288 (N_2288,N_2226,N_2231);
or U2289 (N_2289,N_2231,N_2235);
or U2290 (N_2290,N_2228,N_2222);
nor U2291 (N_2291,N_2211,N_2220);
nand U2292 (N_2292,N_2212,N_2240);
or U2293 (N_2293,N_2247,N_2216);
and U2294 (N_2294,N_2208,N_2247);
or U2295 (N_2295,N_2237,N_2227);
nor U2296 (N_2296,N_2200,N_2240);
nand U2297 (N_2297,N_2216,N_2226);
and U2298 (N_2298,N_2245,N_2221);
nand U2299 (N_2299,N_2235,N_2238);
and U2300 (N_2300,N_2256,N_2280);
nor U2301 (N_2301,N_2252,N_2274);
xor U2302 (N_2302,N_2250,N_2261);
and U2303 (N_2303,N_2253,N_2255);
or U2304 (N_2304,N_2299,N_2259);
or U2305 (N_2305,N_2297,N_2263);
and U2306 (N_2306,N_2295,N_2290);
and U2307 (N_2307,N_2270,N_2266);
and U2308 (N_2308,N_2279,N_2282);
nand U2309 (N_2309,N_2296,N_2284);
nor U2310 (N_2310,N_2294,N_2276);
and U2311 (N_2311,N_2281,N_2283);
xnor U2312 (N_2312,N_2271,N_2298);
and U2313 (N_2313,N_2268,N_2289);
xor U2314 (N_2314,N_2293,N_2278);
and U2315 (N_2315,N_2257,N_2273);
nor U2316 (N_2316,N_2275,N_2288);
nor U2317 (N_2317,N_2286,N_2260);
and U2318 (N_2318,N_2272,N_2262);
nand U2319 (N_2319,N_2292,N_2291);
nor U2320 (N_2320,N_2254,N_2269);
nand U2321 (N_2321,N_2285,N_2251);
xor U2322 (N_2322,N_2287,N_2258);
nor U2323 (N_2323,N_2277,N_2267);
nor U2324 (N_2324,N_2265,N_2264);
and U2325 (N_2325,N_2296,N_2265);
nor U2326 (N_2326,N_2298,N_2297);
nand U2327 (N_2327,N_2260,N_2251);
or U2328 (N_2328,N_2278,N_2271);
and U2329 (N_2329,N_2267,N_2294);
nand U2330 (N_2330,N_2296,N_2272);
or U2331 (N_2331,N_2277,N_2276);
and U2332 (N_2332,N_2272,N_2260);
nand U2333 (N_2333,N_2263,N_2299);
nor U2334 (N_2334,N_2251,N_2261);
and U2335 (N_2335,N_2290,N_2287);
xor U2336 (N_2336,N_2262,N_2251);
nor U2337 (N_2337,N_2254,N_2279);
nor U2338 (N_2338,N_2250,N_2274);
nand U2339 (N_2339,N_2250,N_2284);
and U2340 (N_2340,N_2265,N_2273);
nand U2341 (N_2341,N_2250,N_2294);
and U2342 (N_2342,N_2263,N_2250);
or U2343 (N_2343,N_2262,N_2259);
and U2344 (N_2344,N_2282,N_2295);
nand U2345 (N_2345,N_2269,N_2289);
nand U2346 (N_2346,N_2283,N_2261);
or U2347 (N_2347,N_2250,N_2258);
and U2348 (N_2348,N_2263,N_2289);
nor U2349 (N_2349,N_2261,N_2293);
nor U2350 (N_2350,N_2324,N_2328);
nand U2351 (N_2351,N_2319,N_2311);
or U2352 (N_2352,N_2342,N_2339);
xnor U2353 (N_2353,N_2303,N_2308);
xnor U2354 (N_2354,N_2300,N_2335);
and U2355 (N_2355,N_2332,N_2316);
nor U2356 (N_2356,N_2337,N_2330);
xnor U2357 (N_2357,N_2315,N_2336);
nand U2358 (N_2358,N_2325,N_2304);
nor U2359 (N_2359,N_2323,N_2318);
and U2360 (N_2360,N_2321,N_2331);
and U2361 (N_2361,N_2341,N_2344);
nor U2362 (N_2362,N_2326,N_2334);
or U2363 (N_2363,N_2320,N_2313);
nand U2364 (N_2364,N_2322,N_2343);
and U2365 (N_2365,N_2346,N_2347);
nand U2366 (N_2366,N_2301,N_2314);
or U2367 (N_2367,N_2338,N_2349);
nand U2368 (N_2368,N_2329,N_2345);
nor U2369 (N_2369,N_2317,N_2310);
or U2370 (N_2370,N_2306,N_2312);
nand U2371 (N_2371,N_2327,N_2340);
nor U2372 (N_2372,N_2309,N_2307);
or U2373 (N_2373,N_2305,N_2333);
xnor U2374 (N_2374,N_2302,N_2348);
nor U2375 (N_2375,N_2347,N_2324);
xor U2376 (N_2376,N_2312,N_2300);
and U2377 (N_2377,N_2324,N_2334);
nand U2378 (N_2378,N_2322,N_2321);
and U2379 (N_2379,N_2343,N_2310);
nand U2380 (N_2380,N_2343,N_2341);
and U2381 (N_2381,N_2315,N_2346);
nor U2382 (N_2382,N_2309,N_2324);
and U2383 (N_2383,N_2315,N_2306);
and U2384 (N_2384,N_2306,N_2340);
nand U2385 (N_2385,N_2307,N_2335);
nand U2386 (N_2386,N_2323,N_2322);
and U2387 (N_2387,N_2321,N_2336);
or U2388 (N_2388,N_2325,N_2307);
or U2389 (N_2389,N_2316,N_2310);
xor U2390 (N_2390,N_2332,N_2317);
nor U2391 (N_2391,N_2313,N_2341);
nor U2392 (N_2392,N_2335,N_2316);
nand U2393 (N_2393,N_2341,N_2312);
nor U2394 (N_2394,N_2323,N_2330);
or U2395 (N_2395,N_2315,N_2305);
nand U2396 (N_2396,N_2329,N_2327);
or U2397 (N_2397,N_2315,N_2343);
nand U2398 (N_2398,N_2307,N_2326);
and U2399 (N_2399,N_2312,N_2316);
nand U2400 (N_2400,N_2358,N_2351);
and U2401 (N_2401,N_2385,N_2381);
xnor U2402 (N_2402,N_2398,N_2366);
or U2403 (N_2403,N_2373,N_2387);
and U2404 (N_2404,N_2367,N_2393);
or U2405 (N_2405,N_2375,N_2374);
or U2406 (N_2406,N_2353,N_2380);
nor U2407 (N_2407,N_2378,N_2363);
xor U2408 (N_2408,N_2362,N_2392);
and U2409 (N_2409,N_2396,N_2355);
nor U2410 (N_2410,N_2364,N_2352);
nand U2411 (N_2411,N_2379,N_2369);
nor U2412 (N_2412,N_2365,N_2388);
and U2413 (N_2413,N_2371,N_2399);
nor U2414 (N_2414,N_2386,N_2350);
nor U2415 (N_2415,N_2394,N_2383);
or U2416 (N_2416,N_2391,N_2390);
nand U2417 (N_2417,N_2377,N_2356);
and U2418 (N_2418,N_2397,N_2357);
nand U2419 (N_2419,N_2382,N_2359);
or U2420 (N_2420,N_2376,N_2354);
and U2421 (N_2421,N_2372,N_2389);
or U2422 (N_2422,N_2370,N_2384);
nor U2423 (N_2423,N_2361,N_2360);
and U2424 (N_2424,N_2368,N_2395);
or U2425 (N_2425,N_2385,N_2360);
nor U2426 (N_2426,N_2394,N_2374);
and U2427 (N_2427,N_2352,N_2393);
nor U2428 (N_2428,N_2381,N_2364);
nand U2429 (N_2429,N_2392,N_2354);
nor U2430 (N_2430,N_2352,N_2358);
or U2431 (N_2431,N_2394,N_2385);
or U2432 (N_2432,N_2385,N_2376);
or U2433 (N_2433,N_2358,N_2397);
or U2434 (N_2434,N_2373,N_2376);
nor U2435 (N_2435,N_2384,N_2385);
or U2436 (N_2436,N_2354,N_2372);
nor U2437 (N_2437,N_2359,N_2352);
nor U2438 (N_2438,N_2389,N_2356);
and U2439 (N_2439,N_2355,N_2381);
nor U2440 (N_2440,N_2371,N_2370);
xor U2441 (N_2441,N_2368,N_2365);
or U2442 (N_2442,N_2352,N_2390);
nor U2443 (N_2443,N_2351,N_2353);
xor U2444 (N_2444,N_2389,N_2354);
nand U2445 (N_2445,N_2361,N_2353);
or U2446 (N_2446,N_2378,N_2356);
nor U2447 (N_2447,N_2369,N_2386);
and U2448 (N_2448,N_2374,N_2355);
and U2449 (N_2449,N_2373,N_2386);
nand U2450 (N_2450,N_2420,N_2438);
or U2451 (N_2451,N_2444,N_2418);
and U2452 (N_2452,N_2421,N_2417);
or U2453 (N_2453,N_2430,N_2407);
nor U2454 (N_2454,N_2432,N_2423);
nand U2455 (N_2455,N_2448,N_2412);
nor U2456 (N_2456,N_2413,N_2443);
or U2457 (N_2457,N_2446,N_2411);
xor U2458 (N_2458,N_2433,N_2439);
nand U2459 (N_2459,N_2447,N_2429);
and U2460 (N_2460,N_2449,N_2406);
nor U2461 (N_2461,N_2441,N_2422);
nor U2462 (N_2462,N_2425,N_2435);
and U2463 (N_2463,N_2419,N_2437);
xnor U2464 (N_2464,N_2401,N_2445);
or U2465 (N_2465,N_2440,N_2405);
and U2466 (N_2466,N_2428,N_2431);
or U2467 (N_2467,N_2404,N_2442);
or U2468 (N_2468,N_2414,N_2409);
nand U2469 (N_2469,N_2403,N_2434);
nand U2470 (N_2470,N_2426,N_2427);
and U2471 (N_2471,N_2416,N_2424);
nand U2472 (N_2472,N_2436,N_2402);
and U2473 (N_2473,N_2400,N_2408);
nor U2474 (N_2474,N_2410,N_2415);
nor U2475 (N_2475,N_2429,N_2414);
or U2476 (N_2476,N_2416,N_2446);
nor U2477 (N_2477,N_2441,N_2427);
xnor U2478 (N_2478,N_2441,N_2430);
and U2479 (N_2479,N_2425,N_2439);
nor U2480 (N_2480,N_2420,N_2424);
xor U2481 (N_2481,N_2403,N_2423);
and U2482 (N_2482,N_2431,N_2409);
and U2483 (N_2483,N_2446,N_2428);
and U2484 (N_2484,N_2449,N_2425);
and U2485 (N_2485,N_2412,N_2429);
nor U2486 (N_2486,N_2432,N_2403);
nand U2487 (N_2487,N_2402,N_2428);
nor U2488 (N_2488,N_2401,N_2407);
nand U2489 (N_2489,N_2427,N_2437);
and U2490 (N_2490,N_2449,N_2415);
and U2491 (N_2491,N_2445,N_2448);
or U2492 (N_2492,N_2412,N_2446);
or U2493 (N_2493,N_2409,N_2410);
xnor U2494 (N_2494,N_2401,N_2448);
nand U2495 (N_2495,N_2403,N_2428);
nor U2496 (N_2496,N_2410,N_2405);
nor U2497 (N_2497,N_2430,N_2417);
nor U2498 (N_2498,N_2417,N_2424);
and U2499 (N_2499,N_2415,N_2438);
and U2500 (N_2500,N_2481,N_2463);
and U2501 (N_2501,N_2499,N_2483);
and U2502 (N_2502,N_2461,N_2478);
nor U2503 (N_2503,N_2490,N_2452);
xnor U2504 (N_2504,N_2458,N_2489);
or U2505 (N_2505,N_2497,N_2454);
or U2506 (N_2506,N_2459,N_2469);
or U2507 (N_2507,N_2475,N_2486);
and U2508 (N_2508,N_2492,N_2484);
or U2509 (N_2509,N_2470,N_2491);
nor U2510 (N_2510,N_2476,N_2487);
or U2511 (N_2511,N_2460,N_2455);
nand U2512 (N_2512,N_2473,N_2453);
nand U2513 (N_2513,N_2493,N_2474);
or U2514 (N_2514,N_2456,N_2472);
nand U2515 (N_2515,N_2465,N_2488);
nand U2516 (N_2516,N_2457,N_2466);
nor U2517 (N_2517,N_2482,N_2480);
nor U2518 (N_2518,N_2467,N_2471);
or U2519 (N_2519,N_2451,N_2496);
nand U2520 (N_2520,N_2485,N_2477);
nand U2521 (N_2521,N_2494,N_2450);
nor U2522 (N_2522,N_2495,N_2468);
nand U2523 (N_2523,N_2498,N_2462);
nand U2524 (N_2524,N_2479,N_2464);
nor U2525 (N_2525,N_2452,N_2478);
or U2526 (N_2526,N_2472,N_2495);
and U2527 (N_2527,N_2456,N_2498);
and U2528 (N_2528,N_2490,N_2497);
and U2529 (N_2529,N_2460,N_2486);
or U2530 (N_2530,N_2492,N_2461);
xnor U2531 (N_2531,N_2450,N_2484);
nand U2532 (N_2532,N_2476,N_2489);
nand U2533 (N_2533,N_2478,N_2487);
and U2534 (N_2534,N_2484,N_2459);
nor U2535 (N_2535,N_2468,N_2492);
or U2536 (N_2536,N_2475,N_2461);
and U2537 (N_2537,N_2455,N_2465);
nor U2538 (N_2538,N_2469,N_2455);
and U2539 (N_2539,N_2468,N_2487);
nand U2540 (N_2540,N_2486,N_2462);
nor U2541 (N_2541,N_2471,N_2483);
or U2542 (N_2542,N_2454,N_2480);
nor U2543 (N_2543,N_2485,N_2499);
nand U2544 (N_2544,N_2497,N_2494);
nand U2545 (N_2545,N_2472,N_2479);
nor U2546 (N_2546,N_2466,N_2475);
nor U2547 (N_2547,N_2468,N_2464);
and U2548 (N_2548,N_2457,N_2459);
nand U2549 (N_2549,N_2490,N_2468);
nand U2550 (N_2550,N_2524,N_2538);
nand U2551 (N_2551,N_2545,N_2502);
xnor U2552 (N_2552,N_2540,N_2534);
or U2553 (N_2553,N_2546,N_2531);
nor U2554 (N_2554,N_2541,N_2514);
or U2555 (N_2555,N_2507,N_2505);
or U2556 (N_2556,N_2535,N_2522);
nor U2557 (N_2557,N_2513,N_2516);
xnor U2558 (N_2558,N_2519,N_2527);
nand U2559 (N_2559,N_2533,N_2504);
and U2560 (N_2560,N_2508,N_2529);
xor U2561 (N_2561,N_2547,N_2501);
and U2562 (N_2562,N_2511,N_2530);
or U2563 (N_2563,N_2506,N_2549);
and U2564 (N_2564,N_2515,N_2509);
and U2565 (N_2565,N_2542,N_2503);
nor U2566 (N_2566,N_2548,N_2517);
or U2567 (N_2567,N_2525,N_2543);
and U2568 (N_2568,N_2536,N_2526);
nor U2569 (N_2569,N_2520,N_2512);
nor U2570 (N_2570,N_2523,N_2518);
or U2571 (N_2571,N_2510,N_2528);
xor U2572 (N_2572,N_2544,N_2532);
nor U2573 (N_2573,N_2500,N_2539);
nand U2574 (N_2574,N_2521,N_2537);
and U2575 (N_2575,N_2516,N_2536);
nor U2576 (N_2576,N_2544,N_2530);
or U2577 (N_2577,N_2525,N_2547);
and U2578 (N_2578,N_2531,N_2518);
or U2579 (N_2579,N_2519,N_2505);
nand U2580 (N_2580,N_2543,N_2505);
and U2581 (N_2581,N_2539,N_2523);
nand U2582 (N_2582,N_2533,N_2508);
or U2583 (N_2583,N_2542,N_2531);
or U2584 (N_2584,N_2512,N_2523);
and U2585 (N_2585,N_2532,N_2515);
nor U2586 (N_2586,N_2537,N_2515);
nor U2587 (N_2587,N_2533,N_2500);
or U2588 (N_2588,N_2506,N_2547);
and U2589 (N_2589,N_2546,N_2541);
and U2590 (N_2590,N_2543,N_2541);
and U2591 (N_2591,N_2549,N_2520);
or U2592 (N_2592,N_2549,N_2540);
and U2593 (N_2593,N_2543,N_2516);
or U2594 (N_2594,N_2508,N_2506);
or U2595 (N_2595,N_2521,N_2548);
or U2596 (N_2596,N_2542,N_2516);
nand U2597 (N_2597,N_2514,N_2525);
nand U2598 (N_2598,N_2536,N_2508);
nand U2599 (N_2599,N_2507,N_2523);
nand U2600 (N_2600,N_2589,N_2594);
xor U2601 (N_2601,N_2550,N_2560);
and U2602 (N_2602,N_2571,N_2559);
and U2603 (N_2603,N_2577,N_2573);
nor U2604 (N_2604,N_2593,N_2553);
nor U2605 (N_2605,N_2581,N_2570);
nand U2606 (N_2606,N_2557,N_2579);
nor U2607 (N_2607,N_2578,N_2563);
nand U2608 (N_2608,N_2552,N_2592);
nor U2609 (N_2609,N_2569,N_2586);
nand U2610 (N_2610,N_2590,N_2572);
and U2611 (N_2611,N_2558,N_2583);
nor U2612 (N_2612,N_2596,N_2576);
xnor U2613 (N_2613,N_2554,N_2595);
or U2614 (N_2614,N_2584,N_2551);
and U2615 (N_2615,N_2555,N_2598);
and U2616 (N_2616,N_2582,N_2574);
and U2617 (N_2617,N_2567,N_2566);
nor U2618 (N_2618,N_2564,N_2580);
or U2619 (N_2619,N_2575,N_2561);
nand U2620 (N_2620,N_2597,N_2587);
and U2621 (N_2621,N_2599,N_2565);
nand U2622 (N_2622,N_2562,N_2591);
nand U2623 (N_2623,N_2588,N_2556);
xnor U2624 (N_2624,N_2585,N_2568);
nor U2625 (N_2625,N_2593,N_2565);
nor U2626 (N_2626,N_2596,N_2558);
nand U2627 (N_2627,N_2598,N_2593);
nor U2628 (N_2628,N_2585,N_2553);
nor U2629 (N_2629,N_2567,N_2564);
nor U2630 (N_2630,N_2550,N_2556);
or U2631 (N_2631,N_2578,N_2587);
and U2632 (N_2632,N_2576,N_2595);
xnor U2633 (N_2633,N_2562,N_2583);
or U2634 (N_2634,N_2587,N_2560);
or U2635 (N_2635,N_2572,N_2594);
or U2636 (N_2636,N_2593,N_2577);
nand U2637 (N_2637,N_2589,N_2592);
nor U2638 (N_2638,N_2561,N_2590);
xnor U2639 (N_2639,N_2559,N_2573);
and U2640 (N_2640,N_2577,N_2574);
nor U2641 (N_2641,N_2575,N_2551);
or U2642 (N_2642,N_2566,N_2571);
or U2643 (N_2643,N_2575,N_2595);
or U2644 (N_2644,N_2578,N_2582);
nand U2645 (N_2645,N_2568,N_2573);
and U2646 (N_2646,N_2558,N_2570);
and U2647 (N_2647,N_2583,N_2575);
nor U2648 (N_2648,N_2594,N_2560);
and U2649 (N_2649,N_2562,N_2578);
or U2650 (N_2650,N_2608,N_2616);
nor U2651 (N_2651,N_2622,N_2605);
or U2652 (N_2652,N_2603,N_2618);
and U2653 (N_2653,N_2640,N_2625);
and U2654 (N_2654,N_2606,N_2648);
nor U2655 (N_2655,N_2636,N_2634);
nand U2656 (N_2656,N_2629,N_2617);
and U2657 (N_2657,N_2632,N_2637);
or U2658 (N_2658,N_2643,N_2635);
and U2659 (N_2659,N_2627,N_2626);
or U2660 (N_2660,N_2620,N_2614);
and U2661 (N_2661,N_2641,N_2610);
and U2662 (N_2662,N_2630,N_2628);
nand U2663 (N_2663,N_2644,N_2646);
or U2664 (N_2664,N_2621,N_2615);
or U2665 (N_2665,N_2647,N_2645);
nand U2666 (N_2666,N_2639,N_2604);
nand U2667 (N_2667,N_2600,N_2611);
xor U2668 (N_2668,N_2638,N_2601);
and U2669 (N_2669,N_2624,N_2631);
nand U2670 (N_2670,N_2602,N_2609);
nor U2671 (N_2671,N_2642,N_2619);
xnor U2672 (N_2672,N_2607,N_2649);
or U2673 (N_2673,N_2623,N_2633);
nor U2674 (N_2674,N_2613,N_2612);
and U2675 (N_2675,N_2647,N_2648);
or U2676 (N_2676,N_2639,N_2620);
or U2677 (N_2677,N_2631,N_2649);
nor U2678 (N_2678,N_2634,N_2644);
nor U2679 (N_2679,N_2638,N_2619);
nand U2680 (N_2680,N_2630,N_2618);
or U2681 (N_2681,N_2638,N_2622);
or U2682 (N_2682,N_2633,N_2614);
and U2683 (N_2683,N_2608,N_2634);
nand U2684 (N_2684,N_2622,N_2625);
and U2685 (N_2685,N_2643,N_2626);
or U2686 (N_2686,N_2612,N_2649);
nand U2687 (N_2687,N_2649,N_2604);
nand U2688 (N_2688,N_2613,N_2649);
xnor U2689 (N_2689,N_2622,N_2632);
nand U2690 (N_2690,N_2631,N_2603);
nor U2691 (N_2691,N_2647,N_2634);
or U2692 (N_2692,N_2604,N_2605);
and U2693 (N_2693,N_2636,N_2631);
nor U2694 (N_2694,N_2620,N_2606);
and U2695 (N_2695,N_2638,N_2639);
nand U2696 (N_2696,N_2648,N_2630);
or U2697 (N_2697,N_2637,N_2610);
and U2698 (N_2698,N_2623,N_2621);
nor U2699 (N_2699,N_2611,N_2649);
nor U2700 (N_2700,N_2671,N_2664);
nand U2701 (N_2701,N_2673,N_2665);
and U2702 (N_2702,N_2669,N_2699);
nor U2703 (N_2703,N_2675,N_2676);
nand U2704 (N_2704,N_2685,N_2666);
nor U2705 (N_2705,N_2662,N_2659);
nand U2706 (N_2706,N_2652,N_2678);
xnor U2707 (N_2707,N_2680,N_2663);
nor U2708 (N_2708,N_2679,N_2651);
and U2709 (N_2709,N_2672,N_2668);
nand U2710 (N_2710,N_2653,N_2667);
and U2711 (N_2711,N_2689,N_2670);
and U2712 (N_2712,N_2695,N_2660);
nor U2713 (N_2713,N_2687,N_2654);
or U2714 (N_2714,N_2682,N_2686);
nor U2715 (N_2715,N_2693,N_2658);
nand U2716 (N_2716,N_2694,N_2657);
or U2717 (N_2717,N_2650,N_2698);
nand U2718 (N_2718,N_2688,N_2677);
nor U2719 (N_2719,N_2690,N_2683);
nand U2720 (N_2720,N_2696,N_2681);
nand U2721 (N_2721,N_2674,N_2697);
and U2722 (N_2722,N_2661,N_2691);
nand U2723 (N_2723,N_2684,N_2656);
and U2724 (N_2724,N_2655,N_2692);
nor U2725 (N_2725,N_2672,N_2681);
xnor U2726 (N_2726,N_2651,N_2695);
or U2727 (N_2727,N_2654,N_2691);
nor U2728 (N_2728,N_2697,N_2671);
and U2729 (N_2729,N_2683,N_2697);
and U2730 (N_2730,N_2678,N_2685);
nand U2731 (N_2731,N_2690,N_2673);
and U2732 (N_2732,N_2686,N_2650);
xnor U2733 (N_2733,N_2675,N_2666);
nor U2734 (N_2734,N_2659,N_2668);
or U2735 (N_2735,N_2662,N_2671);
or U2736 (N_2736,N_2674,N_2686);
and U2737 (N_2737,N_2660,N_2677);
or U2738 (N_2738,N_2698,N_2696);
nand U2739 (N_2739,N_2680,N_2674);
nand U2740 (N_2740,N_2676,N_2668);
nand U2741 (N_2741,N_2698,N_2669);
and U2742 (N_2742,N_2667,N_2655);
or U2743 (N_2743,N_2683,N_2664);
xnor U2744 (N_2744,N_2676,N_2696);
nor U2745 (N_2745,N_2694,N_2684);
or U2746 (N_2746,N_2676,N_2656);
nor U2747 (N_2747,N_2699,N_2698);
and U2748 (N_2748,N_2692,N_2651);
nor U2749 (N_2749,N_2679,N_2674);
nor U2750 (N_2750,N_2746,N_2717);
or U2751 (N_2751,N_2734,N_2732);
nor U2752 (N_2752,N_2731,N_2735);
nor U2753 (N_2753,N_2730,N_2712);
nand U2754 (N_2754,N_2739,N_2716);
nor U2755 (N_2755,N_2710,N_2700);
xnor U2756 (N_2756,N_2738,N_2708);
or U2757 (N_2757,N_2714,N_2742);
and U2758 (N_2758,N_2725,N_2729);
and U2759 (N_2759,N_2715,N_2748);
nor U2760 (N_2760,N_2745,N_2740);
or U2761 (N_2761,N_2724,N_2720);
and U2762 (N_2762,N_2707,N_2744);
nor U2763 (N_2763,N_2718,N_2727);
and U2764 (N_2764,N_2709,N_2728);
and U2765 (N_2765,N_2702,N_2721);
nand U2766 (N_2766,N_2704,N_2749);
and U2767 (N_2767,N_2747,N_2722);
nor U2768 (N_2768,N_2713,N_2733);
xnor U2769 (N_2769,N_2723,N_2719);
or U2770 (N_2770,N_2705,N_2701);
and U2771 (N_2771,N_2741,N_2726);
xor U2772 (N_2772,N_2706,N_2736);
and U2773 (N_2773,N_2743,N_2703);
or U2774 (N_2774,N_2737,N_2711);
and U2775 (N_2775,N_2747,N_2738);
xnor U2776 (N_2776,N_2746,N_2704);
and U2777 (N_2777,N_2735,N_2713);
nor U2778 (N_2778,N_2746,N_2708);
nand U2779 (N_2779,N_2711,N_2746);
nor U2780 (N_2780,N_2744,N_2725);
or U2781 (N_2781,N_2731,N_2743);
and U2782 (N_2782,N_2716,N_2727);
and U2783 (N_2783,N_2732,N_2723);
nand U2784 (N_2784,N_2720,N_2736);
nand U2785 (N_2785,N_2727,N_2739);
nor U2786 (N_2786,N_2723,N_2702);
nand U2787 (N_2787,N_2704,N_2700);
nand U2788 (N_2788,N_2720,N_2746);
and U2789 (N_2789,N_2712,N_2714);
nor U2790 (N_2790,N_2721,N_2731);
and U2791 (N_2791,N_2724,N_2700);
xnor U2792 (N_2792,N_2742,N_2726);
and U2793 (N_2793,N_2749,N_2706);
nand U2794 (N_2794,N_2702,N_2705);
and U2795 (N_2795,N_2719,N_2703);
nand U2796 (N_2796,N_2732,N_2722);
and U2797 (N_2797,N_2711,N_2725);
nor U2798 (N_2798,N_2740,N_2741);
or U2799 (N_2799,N_2735,N_2715);
nand U2800 (N_2800,N_2786,N_2766);
or U2801 (N_2801,N_2777,N_2751);
or U2802 (N_2802,N_2798,N_2762);
nand U2803 (N_2803,N_2767,N_2797);
and U2804 (N_2804,N_2773,N_2796);
xnor U2805 (N_2805,N_2760,N_2763);
and U2806 (N_2806,N_2793,N_2799);
and U2807 (N_2807,N_2770,N_2755);
nand U2808 (N_2808,N_2789,N_2781);
or U2809 (N_2809,N_2778,N_2776);
and U2810 (N_2810,N_2779,N_2750);
or U2811 (N_2811,N_2787,N_2782);
nand U2812 (N_2812,N_2765,N_2756);
and U2813 (N_2813,N_2788,N_2791);
xnor U2814 (N_2814,N_2783,N_2780);
nand U2815 (N_2815,N_2761,N_2792);
nor U2816 (N_2816,N_2769,N_2752);
or U2817 (N_2817,N_2753,N_2775);
nand U2818 (N_2818,N_2759,N_2785);
or U2819 (N_2819,N_2794,N_2772);
xnor U2820 (N_2820,N_2758,N_2768);
or U2821 (N_2821,N_2764,N_2790);
or U2822 (N_2822,N_2784,N_2754);
nand U2823 (N_2823,N_2774,N_2757);
or U2824 (N_2824,N_2771,N_2795);
or U2825 (N_2825,N_2778,N_2771);
nor U2826 (N_2826,N_2757,N_2792);
or U2827 (N_2827,N_2758,N_2776);
nor U2828 (N_2828,N_2787,N_2784);
nor U2829 (N_2829,N_2799,N_2777);
nand U2830 (N_2830,N_2752,N_2758);
nand U2831 (N_2831,N_2753,N_2751);
or U2832 (N_2832,N_2798,N_2761);
nand U2833 (N_2833,N_2755,N_2785);
or U2834 (N_2834,N_2782,N_2772);
and U2835 (N_2835,N_2771,N_2791);
or U2836 (N_2836,N_2793,N_2794);
nor U2837 (N_2837,N_2793,N_2796);
nor U2838 (N_2838,N_2763,N_2759);
or U2839 (N_2839,N_2756,N_2750);
nand U2840 (N_2840,N_2782,N_2752);
nand U2841 (N_2841,N_2796,N_2783);
nand U2842 (N_2842,N_2798,N_2793);
and U2843 (N_2843,N_2759,N_2760);
and U2844 (N_2844,N_2776,N_2796);
xor U2845 (N_2845,N_2786,N_2781);
and U2846 (N_2846,N_2794,N_2751);
and U2847 (N_2847,N_2755,N_2750);
nand U2848 (N_2848,N_2753,N_2773);
nand U2849 (N_2849,N_2785,N_2750);
or U2850 (N_2850,N_2844,N_2827);
xor U2851 (N_2851,N_2825,N_2819);
nand U2852 (N_2852,N_2807,N_2833);
or U2853 (N_2853,N_2848,N_2816);
nand U2854 (N_2854,N_2808,N_2802);
and U2855 (N_2855,N_2806,N_2846);
nand U2856 (N_2856,N_2847,N_2817);
and U2857 (N_2857,N_2839,N_2810);
and U2858 (N_2858,N_2840,N_2820);
nand U2859 (N_2859,N_2800,N_2831);
xor U2860 (N_2860,N_2835,N_2841);
nand U2861 (N_2861,N_2849,N_2818);
nor U2862 (N_2862,N_2836,N_2824);
nand U2863 (N_2863,N_2837,N_2815);
and U2864 (N_2864,N_2826,N_2838);
nor U2865 (N_2865,N_2829,N_2823);
nand U2866 (N_2866,N_2842,N_2822);
nand U2867 (N_2867,N_2830,N_2811);
and U2868 (N_2868,N_2813,N_2804);
nand U2869 (N_2869,N_2812,N_2832);
and U2870 (N_2870,N_2801,N_2805);
and U2871 (N_2871,N_2821,N_2809);
nor U2872 (N_2872,N_2803,N_2845);
nand U2873 (N_2873,N_2814,N_2843);
nand U2874 (N_2874,N_2828,N_2834);
and U2875 (N_2875,N_2833,N_2804);
and U2876 (N_2876,N_2847,N_2824);
nand U2877 (N_2877,N_2829,N_2820);
nand U2878 (N_2878,N_2821,N_2842);
and U2879 (N_2879,N_2838,N_2832);
and U2880 (N_2880,N_2803,N_2819);
or U2881 (N_2881,N_2829,N_2842);
nor U2882 (N_2882,N_2836,N_2803);
and U2883 (N_2883,N_2831,N_2801);
and U2884 (N_2884,N_2803,N_2801);
and U2885 (N_2885,N_2845,N_2831);
nand U2886 (N_2886,N_2837,N_2835);
or U2887 (N_2887,N_2801,N_2820);
and U2888 (N_2888,N_2849,N_2842);
nand U2889 (N_2889,N_2830,N_2802);
and U2890 (N_2890,N_2847,N_2848);
nor U2891 (N_2891,N_2807,N_2809);
nand U2892 (N_2892,N_2823,N_2835);
nand U2893 (N_2893,N_2843,N_2842);
or U2894 (N_2894,N_2845,N_2818);
and U2895 (N_2895,N_2830,N_2813);
nand U2896 (N_2896,N_2837,N_2826);
nand U2897 (N_2897,N_2801,N_2829);
nand U2898 (N_2898,N_2848,N_2810);
xnor U2899 (N_2899,N_2846,N_2802);
nand U2900 (N_2900,N_2868,N_2872);
or U2901 (N_2901,N_2878,N_2894);
or U2902 (N_2902,N_2865,N_2851);
and U2903 (N_2903,N_2895,N_2864);
nand U2904 (N_2904,N_2882,N_2869);
or U2905 (N_2905,N_2890,N_2880);
nand U2906 (N_2906,N_2856,N_2853);
nand U2907 (N_2907,N_2886,N_2898);
nor U2908 (N_2908,N_2862,N_2874);
or U2909 (N_2909,N_2891,N_2875);
xor U2910 (N_2910,N_2896,N_2870);
nor U2911 (N_2911,N_2855,N_2852);
nand U2912 (N_2912,N_2857,N_2867);
or U2913 (N_2913,N_2888,N_2889);
and U2914 (N_2914,N_2860,N_2897);
and U2915 (N_2915,N_2858,N_2861);
and U2916 (N_2916,N_2893,N_2854);
xnor U2917 (N_2917,N_2866,N_2876);
or U2918 (N_2918,N_2892,N_2899);
nand U2919 (N_2919,N_2887,N_2881);
nor U2920 (N_2920,N_2873,N_2871);
and U2921 (N_2921,N_2859,N_2877);
and U2922 (N_2922,N_2850,N_2884);
and U2923 (N_2923,N_2883,N_2879);
and U2924 (N_2924,N_2885,N_2863);
or U2925 (N_2925,N_2873,N_2899);
or U2926 (N_2926,N_2890,N_2865);
or U2927 (N_2927,N_2869,N_2892);
xor U2928 (N_2928,N_2852,N_2873);
xor U2929 (N_2929,N_2861,N_2892);
or U2930 (N_2930,N_2896,N_2873);
and U2931 (N_2931,N_2898,N_2875);
nand U2932 (N_2932,N_2858,N_2870);
nor U2933 (N_2933,N_2860,N_2896);
nand U2934 (N_2934,N_2863,N_2873);
or U2935 (N_2935,N_2892,N_2886);
xor U2936 (N_2936,N_2873,N_2872);
and U2937 (N_2937,N_2851,N_2894);
or U2938 (N_2938,N_2893,N_2898);
or U2939 (N_2939,N_2881,N_2863);
and U2940 (N_2940,N_2865,N_2866);
and U2941 (N_2941,N_2874,N_2876);
nand U2942 (N_2942,N_2894,N_2890);
nand U2943 (N_2943,N_2882,N_2853);
or U2944 (N_2944,N_2872,N_2898);
nand U2945 (N_2945,N_2892,N_2867);
or U2946 (N_2946,N_2875,N_2885);
or U2947 (N_2947,N_2894,N_2895);
and U2948 (N_2948,N_2883,N_2893);
or U2949 (N_2949,N_2883,N_2890);
or U2950 (N_2950,N_2923,N_2947);
and U2951 (N_2951,N_2945,N_2946);
xnor U2952 (N_2952,N_2937,N_2914);
nor U2953 (N_2953,N_2938,N_2918);
or U2954 (N_2954,N_2915,N_2928);
nand U2955 (N_2955,N_2901,N_2939);
or U2956 (N_2956,N_2920,N_2930);
nor U2957 (N_2957,N_2924,N_2943);
nor U2958 (N_2958,N_2935,N_2902);
and U2959 (N_2959,N_2907,N_2941);
and U2960 (N_2960,N_2927,N_2916);
nand U2961 (N_2961,N_2936,N_2904);
and U2962 (N_2962,N_2922,N_2944);
nor U2963 (N_2963,N_2934,N_2913);
xnor U2964 (N_2964,N_2929,N_2949);
nand U2965 (N_2965,N_2912,N_2942);
nand U2966 (N_2966,N_2925,N_2909);
or U2967 (N_2967,N_2933,N_2921);
nor U2968 (N_2968,N_2917,N_2903);
nand U2969 (N_2969,N_2911,N_2908);
nor U2970 (N_2970,N_2926,N_2900);
nor U2971 (N_2971,N_2940,N_2905);
nand U2972 (N_2972,N_2919,N_2910);
or U2973 (N_2973,N_2931,N_2932);
or U2974 (N_2974,N_2906,N_2948);
or U2975 (N_2975,N_2900,N_2949);
or U2976 (N_2976,N_2917,N_2936);
or U2977 (N_2977,N_2907,N_2942);
or U2978 (N_2978,N_2908,N_2907);
nand U2979 (N_2979,N_2928,N_2913);
xnor U2980 (N_2980,N_2933,N_2948);
xor U2981 (N_2981,N_2923,N_2904);
nand U2982 (N_2982,N_2925,N_2924);
or U2983 (N_2983,N_2941,N_2913);
and U2984 (N_2984,N_2939,N_2915);
or U2985 (N_2985,N_2917,N_2928);
nand U2986 (N_2986,N_2908,N_2943);
nor U2987 (N_2987,N_2921,N_2916);
nor U2988 (N_2988,N_2940,N_2927);
and U2989 (N_2989,N_2900,N_2927);
or U2990 (N_2990,N_2927,N_2914);
xor U2991 (N_2991,N_2929,N_2907);
nand U2992 (N_2992,N_2913,N_2912);
and U2993 (N_2993,N_2908,N_2948);
nor U2994 (N_2994,N_2911,N_2904);
and U2995 (N_2995,N_2922,N_2935);
nand U2996 (N_2996,N_2924,N_2940);
nand U2997 (N_2997,N_2913,N_2946);
nand U2998 (N_2998,N_2937,N_2921);
nor U2999 (N_2999,N_2910,N_2933);
nor UO_0 (O_0,N_2971,N_2961);
nand UO_1 (O_1,N_2982,N_2998);
nor UO_2 (O_2,N_2969,N_2987);
and UO_3 (O_3,N_2989,N_2956);
xnor UO_4 (O_4,N_2996,N_2975);
and UO_5 (O_5,N_2991,N_2963);
and UO_6 (O_6,N_2988,N_2999);
nor UO_7 (O_7,N_2964,N_2993);
and UO_8 (O_8,N_2972,N_2968);
and UO_9 (O_9,N_2980,N_2997);
nand UO_10 (O_10,N_2952,N_2986);
or UO_11 (O_11,N_2977,N_2959);
nand UO_12 (O_12,N_2984,N_2979);
or UO_13 (O_13,N_2974,N_2990);
nor UO_14 (O_14,N_2973,N_2970);
nor UO_15 (O_15,N_2976,N_2981);
nor UO_16 (O_16,N_2966,N_2960);
and UO_17 (O_17,N_2983,N_2950);
and UO_18 (O_18,N_2985,N_2967);
or UO_19 (O_19,N_2957,N_2954);
or UO_20 (O_20,N_2962,N_2953);
or UO_21 (O_21,N_2992,N_2951);
nor UO_22 (O_22,N_2965,N_2955);
and UO_23 (O_23,N_2995,N_2994);
or UO_24 (O_24,N_2978,N_2958);
or UO_25 (O_25,N_2979,N_2989);
and UO_26 (O_26,N_2960,N_2955);
or UO_27 (O_27,N_2985,N_2980);
and UO_28 (O_28,N_2995,N_2979);
nand UO_29 (O_29,N_2953,N_2970);
and UO_30 (O_30,N_2992,N_2965);
and UO_31 (O_31,N_2988,N_2955);
nand UO_32 (O_32,N_2981,N_2996);
nand UO_33 (O_33,N_2970,N_2974);
nand UO_34 (O_34,N_2991,N_2950);
nand UO_35 (O_35,N_2977,N_2950);
nand UO_36 (O_36,N_2968,N_2956);
xnor UO_37 (O_37,N_2988,N_2958);
or UO_38 (O_38,N_2979,N_2998);
nand UO_39 (O_39,N_2995,N_2969);
nor UO_40 (O_40,N_2986,N_2980);
nand UO_41 (O_41,N_2986,N_2955);
or UO_42 (O_42,N_2979,N_2982);
nand UO_43 (O_43,N_2968,N_2975);
nor UO_44 (O_44,N_2958,N_2992);
nand UO_45 (O_45,N_2965,N_2963);
or UO_46 (O_46,N_2986,N_2994);
nand UO_47 (O_47,N_2990,N_2972);
xor UO_48 (O_48,N_2967,N_2995);
and UO_49 (O_49,N_2963,N_2987);
or UO_50 (O_50,N_2991,N_2982);
xnor UO_51 (O_51,N_2960,N_2961);
nor UO_52 (O_52,N_2989,N_2980);
xnor UO_53 (O_53,N_2988,N_2976);
nor UO_54 (O_54,N_2977,N_2981);
or UO_55 (O_55,N_2987,N_2954);
and UO_56 (O_56,N_2985,N_2999);
or UO_57 (O_57,N_2967,N_2952);
or UO_58 (O_58,N_2997,N_2983);
nor UO_59 (O_59,N_2976,N_2965);
or UO_60 (O_60,N_2962,N_2995);
or UO_61 (O_61,N_2958,N_2961);
nand UO_62 (O_62,N_2993,N_2958);
or UO_63 (O_63,N_2950,N_2965);
and UO_64 (O_64,N_2967,N_2979);
xnor UO_65 (O_65,N_2985,N_2981);
and UO_66 (O_66,N_2990,N_2966);
nand UO_67 (O_67,N_2970,N_2956);
nor UO_68 (O_68,N_2993,N_2980);
nor UO_69 (O_69,N_2966,N_2955);
nor UO_70 (O_70,N_2984,N_2951);
and UO_71 (O_71,N_2982,N_2960);
nor UO_72 (O_72,N_2960,N_2956);
or UO_73 (O_73,N_2957,N_2970);
nand UO_74 (O_74,N_2979,N_2961);
or UO_75 (O_75,N_2971,N_2991);
nand UO_76 (O_76,N_2952,N_2995);
nand UO_77 (O_77,N_2955,N_2963);
nand UO_78 (O_78,N_2970,N_2984);
and UO_79 (O_79,N_2998,N_2994);
nor UO_80 (O_80,N_2955,N_2985);
or UO_81 (O_81,N_2981,N_2956);
nand UO_82 (O_82,N_2999,N_2976);
xor UO_83 (O_83,N_2956,N_2972);
nand UO_84 (O_84,N_2998,N_2968);
nor UO_85 (O_85,N_2983,N_2978);
nor UO_86 (O_86,N_2995,N_2959);
or UO_87 (O_87,N_2978,N_2969);
and UO_88 (O_88,N_2952,N_2988);
or UO_89 (O_89,N_2962,N_2997);
nand UO_90 (O_90,N_2975,N_2958);
nand UO_91 (O_91,N_2962,N_2984);
nor UO_92 (O_92,N_2975,N_2990);
nor UO_93 (O_93,N_2978,N_2964);
nor UO_94 (O_94,N_2973,N_2959);
nand UO_95 (O_95,N_2994,N_2969);
nand UO_96 (O_96,N_2976,N_2974);
or UO_97 (O_97,N_2981,N_2950);
or UO_98 (O_98,N_2969,N_2977);
and UO_99 (O_99,N_2963,N_2961);
xor UO_100 (O_100,N_2981,N_2954);
or UO_101 (O_101,N_2990,N_2983);
xor UO_102 (O_102,N_2993,N_2994);
xor UO_103 (O_103,N_2964,N_2968);
nand UO_104 (O_104,N_2957,N_2950);
or UO_105 (O_105,N_2969,N_2972);
xor UO_106 (O_106,N_2954,N_2956);
and UO_107 (O_107,N_2954,N_2951);
or UO_108 (O_108,N_2956,N_2993);
and UO_109 (O_109,N_2966,N_2995);
and UO_110 (O_110,N_2959,N_2989);
or UO_111 (O_111,N_2971,N_2986);
and UO_112 (O_112,N_2965,N_2969);
nor UO_113 (O_113,N_2994,N_2976);
nor UO_114 (O_114,N_2995,N_2972);
nand UO_115 (O_115,N_2981,N_2967);
and UO_116 (O_116,N_2953,N_2967);
and UO_117 (O_117,N_2957,N_2976);
nor UO_118 (O_118,N_2964,N_2970);
nor UO_119 (O_119,N_2991,N_2969);
or UO_120 (O_120,N_2959,N_2966);
nor UO_121 (O_121,N_2960,N_2954);
or UO_122 (O_122,N_2950,N_2959);
or UO_123 (O_123,N_2985,N_2953);
nand UO_124 (O_124,N_2959,N_2969);
xor UO_125 (O_125,N_2997,N_2998);
nand UO_126 (O_126,N_2999,N_2982);
nand UO_127 (O_127,N_2983,N_2993);
nor UO_128 (O_128,N_2990,N_2960);
or UO_129 (O_129,N_2961,N_2981);
nor UO_130 (O_130,N_2956,N_2997);
nor UO_131 (O_131,N_2979,N_2954);
nor UO_132 (O_132,N_2970,N_2951);
or UO_133 (O_133,N_2988,N_2990);
nor UO_134 (O_134,N_2951,N_2952);
nand UO_135 (O_135,N_2959,N_2999);
nand UO_136 (O_136,N_2950,N_2989);
nand UO_137 (O_137,N_2959,N_2967);
or UO_138 (O_138,N_2992,N_2954);
nand UO_139 (O_139,N_2961,N_2954);
xnor UO_140 (O_140,N_2956,N_2952);
and UO_141 (O_141,N_2990,N_2993);
nor UO_142 (O_142,N_2953,N_2963);
nand UO_143 (O_143,N_2958,N_2989);
nand UO_144 (O_144,N_2971,N_2993);
nor UO_145 (O_145,N_2963,N_2964);
and UO_146 (O_146,N_2975,N_2970);
nor UO_147 (O_147,N_2965,N_2991);
nand UO_148 (O_148,N_2993,N_2976);
nor UO_149 (O_149,N_2980,N_2983);
nor UO_150 (O_150,N_2995,N_2981);
or UO_151 (O_151,N_2983,N_2977);
and UO_152 (O_152,N_2960,N_2970);
and UO_153 (O_153,N_2953,N_2974);
and UO_154 (O_154,N_2959,N_2954);
or UO_155 (O_155,N_2963,N_2984);
nand UO_156 (O_156,N_2961,N_2992);
or UO_157 (O_157,N_2972,N_2978);
nor UO_158 (O_158,N_2994,N_2973);
and UO_159 (O_159,N_2986,N_2979);
nor UO_160 (O_160,N_2985,N_2990);
and UO_161 (O_161,N_2980,N_2978);
and UO_162 (O_162,N_2993,N_2985);
nand UO_163 (O_163,N_2953,N_2989);
nand UO_164 (O_164,N_2994,N_2950);
xor UO_165 (O_165,N_2956,N_2950);
or UO_166 (O_166,N_2989,N_2951);
and UO_167 (O_167,N_2952,N_2983);
and UO_168 (O_168,N_2967,N_2988);
or UO_169 (O_169,N_2989,N_2982);
or UO_170 (O_170,N_2952,N_2997);
nand UO_171 (O_171,N_2977,N_2963);
nand UO_172 (O_172,N_2991,N_2962);
nand UO_173 (O_173,N_2980,N_2982);
and UO_174 (O_174,N_2967,N_2978);
nand UO_175 (O_175,N_2981,N_2984);
xnor UO_176 (O_176,N_2996,N_2967);
or UO_177 (O_177,N_2956,N_2980);
nor UO_178 (O_178,N_2983,N_2991);
nand UO_179 (O_179,N_2989,N_2957);
and UO_180 (O_180,N_2957,N_2962);
and UO_181 (O_181,N_2980,N_2969);
nor UO_182 (O_182,N_2954,N_2991);
and UO_183 (O_183,N_2962,N_2985);
nand UO_184 (O_184,N_2957,N_2984);
nor UO_185 (O_185,N_2952,N_2971);
and UO_186 (O_186,N_2974,N_2984);
nor UO_187 (O_187,N_2983,N_2961);
and UO_188 (O_188,N_2983,N_2968);
nand UO_189 (O_189,N_2978,N_2996);
nor UO_190 (O_190,N_2975,N_2994);
and UO_191 (O_191,N_2963,N_2962);
or UO_192 (O_192,N_2997,N_2978);
nand UO_193 (O_193,N_2977,N_2970);
and UO_194 (O_194,N_2983,N_2984);
nand UO_195 (O_195,N_2955,N_2959);
and UO_196 (O_196,N_2989,N_2964);
nand UO_197 (O_197,N_2967,N_2999);
or UO_198 (O_198,N_2968,N_2957);
nor UO_199 (O_199,N_2992,N_2976);
xnor UO_200 (O_200,N_2991,N_2990);
nor UO_201 (O_201,N_2961,N_2984);
nand UO_202 (O_202,N_2992,N_2973);
xnor UO_203 (O_203,N_2978,N_2982);
or UO_204 (O_204,N_2964,N_2999);
and UO_205 (O_205,N_2997,N_2969);
nand UO_206 (O_206,N_2993,N_2974);
nand UO_207 (O_207,N_2988,N_2965);
and UO_208 (O_208,N_2994,N_2958);
and UO_209 (O_209,N_2978,N_2961);
or UO_210 (O_210,N_2951,N_2981);
nor UO_211 (O_211,N_2954,N_2955);
nor UO_212 (O_212,N_2955,N_2983);
xnor UO_213 (O_213,N_2995,N_2999);
nor UO_214 (O_214,N_2984,N_2980);
or UO_215 (O_215,N_2996,N_2974);
or UO_216 (O_216,N_2967,N_2963);
nor UO_217 (O_217,N_2996,N_2957);
and UO_218 (O_218,N_2958,N_2991);
or UO_219 (O_219,N_2967,N_2997);
nand UO_220 (O_220,N_2983,N_2999);
nor UO_221 (O_221,N_2997,N_2964);
and UO_222 (O_222,N_2974,N_2969);
nand UO_223 (O_223,N_2986,N_2982);
nand UO_224 (O_224,N_2981,N_2991);
xnor UO_225 (O_225,N_2998,N_2975);
nand UO_226 (O_226,N_2966,N_2992);
and UO_227 (O_227,N_2963,N_2983);
and UO_228 (O_228,N_2999,N_2961);
and UO_229 (O_229,N_2950,N_2976);
nand UO_230 (O_230,N_2975,N_2957);
nor UO_231 (O_231,N_2958,N_2962);
and UO_232 (O_232,N_2952,N_2987);
nor UO_233 (O_233,N_2951,N_2977);
nand UO_234 (O_234,N_2979,N_2963);
nand UO_235 (O_235,N_2951,N_2962);
nand UO_236 (O_236,N_2962,N_2955);
nor UO_237 (O_237,N_2980,N_2996);
and UO_238 (O_238,N_2971,N_2992);
xor UO_239 (O_239,N_2960,N_2974);
nor UO_240 (O_240,N_2980,N_2990);
nand UO_241 (O_241,N_2953,N_2964);
and UO_242 (O_242,N_2979,N_2992);
xnor UO_243 (O_243,N_2981,N_2960);
nor UO_244 (O_244,N_2974,N_2971);
nand UO_245 (O_245,N_2973,N_2997);
xor UO_246 (O_246,N_2991,N_2987);
xnor UO_247 (O_247,N_2974,N_2998);
and UO_248 (O_248,N_2964,N_2985);
and UO_249 (O_249,N_2986,N_2976);
or UO_250 (O_250,N_2995,N_2980);
nand UO_251 (O_251,N_2953,N_2976);
and UO_252 (O_252,N_2981,N_2983);
and UO_253 (O_253,N_2950,N_2974);
or UO_254 (O_254,N_2990,N_2992);
or UO_255 (O_255,N_2980,N_2972);
xnor UO_256 (O_256,N_2962,N_2952);
nand UO_257 (O_257,N_2986,N_2950);
xnor UO_258 (O_258,N_2997,N_2976);
and UO_259 (O_259,N_2990,N_2963);
xor UO_260 (O_260,N_2993,N_2966);
nand UO_261 (O_261,N_2973,N_2950);
xor UO_262 (O_262,N_2971,N_2983);
nand UO_263 (O_263,N_2968,N_2982);
and UO_264 (O_264,N_2999,N_2977);
and UO_265 (O_265,N_2982,N_2976);
nand UO_266 (O_266,N_2983,N_2975);
or UO_267 (O_267,N_2960,N_2986);
nand UO_268 (O_268,N_2996,N_2966);
or UO_269 (O_269,N_2990,N_2979);
nand UO_270 (O_270,N_2958,N_2999);
nor UO_271 (O_271,N_2969,N_2966);
nand UO_272 (O_272,N_2969,N_2993);
or UO_273 (O_273,N_2968,N_2994);
nor UO_274 (O_274,N_2975,N_2963);
or UO_275 (O_275,N_2984,N_2982);
and UO_276 (O_276,N_2985,N_2989);
nand UO_277 (O_277,N_2985,N_2984);
or UO_278 (O_278,N_2990,N_2999);
nor UO_279 (O_279,N_2958,N_2972);
and UO_280 (O_280,N_2967,N_2983);
nor UO_281 (O_281,N_2965,N_2996);
or UO_282 (O_282,N_2950,N_2978);
nand UO_283 (O_283,N_2953,N_2998);
nand UO_284 (O_284,N_2971,N_2994);
nand UO_285 (O_285,N_2961,N_2989);
or UO_286 (O_286,N_2989,N_2972);
nand UO_287 (O_287,N_2953,N_2990);
nor UO_288 (O_288,N_2981,N_2966);
and UO_289 (O_289,N_2984,N_2958);
nand UO_290 (O_290,N_2982,N_2962);
nand UO_291 (O_291,N_2995,N_2964);
nor UO_292 (O_292,N_2986,N_2997);
nor UO_293 (O_293,N_2985,N_2976);
nor UO_294 (O_294,N_2967,N_2960);
nand UO_295 (O_295,N_2963,N_2950);
and UO_296 (O_296,N_2968,N_2960);
and UO_297 (O_297,N_2965,N_2985);
nand UO_298 (O_298,N_2966,N_2962);
nand UO_299 (O_299,N_2972,N_2961);
and UO_300 (O_300,N_2966,N_2956);
and UO_301 (O_301,N_2950,N_2997);
or UO_302 (O_302,N_2963,N_2999);
or UO_303 (O_303,N_2988,N_2993);
and UO_304 (O_304,N_2980,N_2965);
nand UO_305 (O_305,N_2965,N_2982);
nor UO_306 (O_306,N_2953,N_2994);
nand UO_307 (O_307,N_2950,N_2961);
and UO_308 (O_308,N_2965,N_2959);
nand UO_309 (O_309,N_2954,N_2977);
nand UO_310 (O_310,N_2965,N_2958);
nand UO_311 (O_311,N_2965,N_2961);
and UO_312 (O_312,N_2974,N_2991);
xnor UO_313 (O_313,N_2974,N_2985);
and UO_314 (O_314,N_2992,N_2993);
nand UO_315 (O_315,N_2976,N_2951);
nand UO_316 (O_316,N_2976,N_2960);
nor UO_317 (O_317,N_2976,N_2971);
and UO_318 (O_318,N_2983,N_2992);
nand UO_319 (O_319,N_2963,N_2996);
and UO_320 (O_320,N_2973,N_2965);
nor UO_321 (O_321,N_2973,N_2951);
or UO_322 (O_322,N_2968,N_2999);
or UO_323 (O_323,N_2991,N_2978);
xor UO_324 (O_324,N_2998,N_2984);
or UO_325 (O_325,N_2989,N_2963);
nor UO_326 (O_326,N_2978,N_2963);
and UO_327 (O_327,N_2987,N_2972);
and UO_328 (O_328,N_2966,N_2978);
nor UO_329 (O_329,N_2972,N_2953);
nor UO_330 (O_330,N_2956,N_2975);
or UO_331 (O_331,N_2967,N_2971);
or UO_332 (O_332,N_2975,N_2967);
nor UO_333 (O_333,N_2971,N_2999);
nor UO_334 (O_334,N_2956,N_2986);
nor UO_335 (O_335,N_2998,N_2991);
nor UO_336 (O_336,N_2986,N_2953);
or UO_337 (O_337,N_2999,N_2979);
nand UO_338 (O_338,N_2974,N_2999);
nand UO_339 (O_339,N_2978,N_2955);
nor UO_340 (O_340,N_2969,N_2957);
and UO_341 (O_341,N_2999,N_2978);
or UO_342 (O_342,N_2964,N_2955);
and UO_343 (O_343,N_2990,N_2964);
and UO_344 (O_344,N_2997,N_2960);
and UO_345 (O_345,N_2957,N_2971);
nand UO_346 (O_346,N_2999,N_2950);
xor UO_347 (O_347,N_2981,N_2982);
xnor UO_348 (O_348,N_2957,N_2958);
nand UO_349 (O_349,N_2960,N_2951);
xor UO_350 (O_350,N_2957,N_2991);
and UO_351 (O_351,N_2995,N_2968);
or UO_352 (O_352,N_2960,N_2980);
and UO_353 (O_353,N_2986,N_2993);
nand UO_354 (O_354,N_2956,N_2969);
and UO_355 (O_355,N_2975,N_2973);
and UO_356 (O_356,N_2952,N_2950);
nor UO_357 (O_357,N_2976,N_2955);
nand UO_358 (O_358,N_2971,N_2996);
or UO_359 (O_359,N_2970,N_2986);
or UO_360 (O_360,N_2955,N_2999);
and UO_361 (O_361,N_2960,N_2964);
and UO_362 (O_362,N_2959,N_2978);
nor UO_363 (O_363,N_2995,N_2954);
nand UO_364 (O_364,N_2984,N_2993);
nor UO_365 (O_365,N_2950,N_2988);
and UO_366 (O_366,N_2986,N_2958);
nor UO_367 (O_367,N_2963,N_2952);
nor UO_368 (O_368,N_2983,N_2986);
and UO_369 (O_369,N_2995,N_2978);
nor UO_370 (O_370,N_2993,N_2968);
and UO_371 (O_371,N_2968,N_2973);
nand UO_372 (O_372,N_2953,N_2968);
or UO_373 (O_373,N_2950,N_2998);
nor UO_374 (O_374,N_2989,N_2969);
nand UO_375 (O_375,N_2957,N_2998);
or UO_376 (O_376,N_2961,N_2993);
or UO_377 (O_377,N_2982,N_2971);
nand UO_378 (O_378,N_2983,N_2956);
nor UO_379 (O_379,N_2962,N_2973);
nor UO_380 (O_380,N_2982,N_2993);
nor UO_381 (O_381,N_2975,N_2984);
nor UO_382 (O_382,N_2967,N_2968);
nor UO_383 (O_383,N_2964,N_2987);
or UO_384 (O_384,N_2980,N_2955);
nand UO_385 (O_385,N_2977,N_2975);
nor UO_386 (O_386,N_2961,N_2969);
or UO_387 (O_387,N_2994,N_2966);
or UO_388 (O_388,N_2951,N_2950);
nor UO_389 (O_389,N_2972,N_2957);
or UO_390 (O_390,N_2953,N_2955);
or UO_391 (O_391,N_2954,N_2986);
nand UO_392 (O_392,N_2978,N_2990);
nand UO_393 (O_393,N_2959,N_2968);
nand UO_394 (O_394,N_2995,N_2982);
and UO_395 (O_395,N_2986,N_2988);
nand UO_396 (O_396,N_2973,N_2969);
xnor UO_397 (O_397,N_2988,N_2998);
or UO_398 (O_398,N_2996,N_2997);
and UO_399 (O_399,N_2998,N_2969);
nand UO_400 (O_400,N_2971,N_2975);
nand UO_401 (O_401,N_2987,N_2976);
or UO_402 (O_402,N_2991,N_2952);
nand UO_403 (O_403,N_2960,N_2975);
nor UO_404 (O_404,N_2979,N_2988);
or UO_405 (O_405,N_2985,N_2966);
nor UO_406 (O_406,N_2968,N_2992);
nor UO_407 (O_407,N_2963,N_2971);
nand UO_408 (O_408,N_2960,N_2987);
nand UO_409 (O_409,N_2998,N_2996);
or UO_410 (O_410,N_2950,N_2968);
nand UO_411 (O_411,N_2968,N_2996);
nor UO_412 (O_412,N_2961,N_2975);
or UO_413 (O_413,N_2964,N_2951);
or UO_414 (O_414,N_2987,N_2994);
nor UO_415 (O_415,N_2999,N_2986);
and UO_416 (O_416,N_2957,N_2987);
xnor UO_417 (O_417,N_2979,N_2962);
or UO_418 (O_418,N_2970,N_2989);
nand UO_419 (O_419,N_2950,N_2960);
or UO_420 (O_420,N_2951,N_2975);
nand UO_421 (O_421,N_2973,N_2960);
nand UO_422 (O_422,N_2993,N_2987);
and UO_423 (O_423,N_2970,N_2996);
nand UO_424 (O_424,N_2996,N_2958);
nor UO_425 (O_425,N_2991,N_2968);
or UO_426 (O_426,N_2975,N_2950);
and UO_427 (O_427,N_2982,N_2973);
or UO_428 (O_428,N_2970,N_2980);
nor UO_429 (O_429,N_2995,N_2992);
nor UO_430 (O_430,N_2982,N_2996);
nor UO_431 (O_431,N_2996,N_2950);
and UO_432 (O_432,N_2985,N_2988);
nand UO_433 (O_433,N_2981,N_2953);
or UO_434 (O_434,N_2977,N_2995);
nor UO_435 (O_435,N_2972,N_2967);
nand UO_436 (O_436,N_2958,N_2987);
xnor UO_437 (O_437,N_2976,N_2964);
or UO_438 (O_438,N_2967,N_2950);
nor UO_439 (O_439,N_2997,N_2971);
and UO_440 (O_440,N_2984,N_2950);
nand UO_441 (O_441,N_2997,N_2958);
and UO_442 (O_442,N_2953,N_2997);
and UO_443 (O_443,N_2988,N_2975);
xnor UO_444 (O_444,N_2951,N_2994);
or UO_445 (O_445,N_2953,N_2950);
and UO_446 (O_446,N_2984,N_2972);
and UO_447 (O_447,N_2952,N_2975);
nor UO_448 (O_448,N_2990,N_2967);
nand UO_449 (O_449,N_2968,N_2978);
and UO_450 (O_450,N_2995,N_2983);
xor UO_451 (O_451,N_2965,N_2981);
xnor UO_452 (O_452,N_2956,N_2990);
nor UO_453 (O_453,N_2973,N_2956);
nand UO_454 (O_454,N_2990,N_2969);
nand UO_455 (O_455,N_2977,N_2978);
nor UO_456 (O_456,N_2956,N_2951);
nor UO_457 (O_457,N_2979,N_2987);
nand UO_458 (O_458,N_2952,N_2994);
or UO_459 (O_459,N_2956,N_2996);
or UO_460 (O_460,N_2978,N_2979);
and UO_461 (O_461,N_2951,N_2968);
xor UO_462 (O_462,N_2953,N_2959);
or UO_463 (O_463,N_2972,N_2971);
or UO_464 (O_464,N_2980,N_2954);
nand UO_465 (O_465,N_2968,N_2965);
nand UO_466 (O_466,N_2975,N_2993);
nor UO_467 (O_467,N_2972,N_2966);
nand UO_468 (O_468,N_2960,N_2972);
nand UO_469 (O_469,N_2997,N_2963);
nand UO_470 (O_470,N_2967,N_2974);
or UO_471 (O_471,N_2983,N_2966);
or UO_472 (O_472,N_2981,N_2992);
nand UO_473 (O_473,N_2956,N_2971);
xnor UO_474 (O_474,N_2994,N_2985);
nor UO_475 (O_475,N_2962,N_2954);
and UO_476 (O_476,N_2964,N_2967);
nor UO_477 (O_477,N_2975,N_2992);
nor UO_478 (O_478,N_2999,N_2975);
and UO_479 (O_479,N_2964,N_2961);
nor UO_480 (O_480,N_2988,N_2973);
or UO_481 (O_481,N_2986,N_2972);
xnor UO_482 (O_482,N_2981,N_2972);
or UO_483 (O_483,N_2953,N_2952);
and UO_484 (O_484,N_2999,N_2973);
and UO_485 (O_485,N_2973,N_2980);
nand UO_486 (O_486,N_2954,N_2998);
nor UO_487 (O_487,N_2997,N_2961);
and UO_488 (O_488,N_2994,N_2965);
or UO_489 (O_489,N_2982,N_2974);
nor UO_490 (O_490,N_2981,N_2974);
or UO_491 (O_491,N_2987,N_2973);
nor UO_492 (O_492,N_2968,N_2970);
and UO_493 (O_493,N_2975,N_2997);
or UO_494 (O_494,N_2997,N_2974);
and UO_495 (O_495,N_2980,N_2967);
and UO_496 (O_496,N_2957,N_2983);
nand UO_497 (O_497,N_2978,N_2956);
xnor UO_498 (O_498,N_2958,N_2959);
nor UO_499 (O_499,N_2954,N_2968);
endmodule