module basic_1500_15000_2000_10_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_64,In_979);
xor U1 (N_1,In_870,In_688);
or U2 (N_2,In_1111,In_588);
nand U3 (N_3,In_1484,In_1029);
and U4 (N_4,In_860,In_74);
nand U5 (N_5,In_674,In_1239);
nor U6 (N_6,In_1322,In_887);
or U7 (N_7,In_1491,In_1082);
xnor U8 (N_8,In_166,In_607);
nor U9 (N_9,In_625,In_1237);
nor U10 (N_10,In_1370,In_1247);
and U11 (N_11,In_1466,In_1285);
or U12 (N_12,In_150,In_444);
or U13 (N_13,In_72,In_1019);
nor U14 (N_14,In_512,In_120);
xor U15 (N_15,In_646,In_1451);
nor U16 (N_16,In_541,In_1292);
nand U17 (N_17,In_1289,In_857);
nor U18 (N_18,In_1261,In_172);
nor U19 (N_19,In_429,In_766);
xor U20 (N_20,In_119,In_827);
nand U21 (N_21,In_1226,In_296);
nor U22 (N_22,In_579,In_148);
nand U23 (N_23,In_1450,In_194);
nor U24 (N_24,In_542,In_775);
nand U25 (N_25,In_585,In_754);
nand U26 (N_26,In_1079,In_87);
and U27 (N_27,In_483,In_480);
nand U28 (N_28,In_1447,In_25);
and U29 (N_29,In_143,In_390);
and U30 (N_30,In_1075,In_1481);
nand U31 (N_31,In_938,In_156);
or U32 (N_32,In_1165,In_1469);
nor U33 (N_33,In_1015,In_1053);
or U34 (N_34,In_339,In_1166);
nand U35 (N_35,In_196,In_812);
and U36 (N_36,In_1021,In_1406);
nand U37 (N_37,In_971,In_245);
and U38 (N_38,In_696,In_170);
xor U39 (N_39,In_42,In_933);
and U40 (N_40,In_1255,In_1238);
nand U41 (N_41,In_69,In_1148);
or U42 (N_42,In_387,In_935);
or U43 (N_43,In_185,In_654);
nand U44 (N_44,In_879,In_1030);
and U45 (N_45,In_1182,In_729);
nand U46 (N_46,In_1337,In_1319);
and U47 (N_47,In_433,In_1036);
xnor U48 (N_48,In_1023,In_1426);
and U49 (N_49,In_1206,In_976);
and U50 (N_50,In_1124,In_792);
xnor U51 (N_51,In_604,In_389);
nand U52 (N_52,In_941,In_1225);
nand U53 (N_53,In_1175,In_551);
nor U54 (N_54,In_1326,In_670);
nand U55 (N_55,In_1083,In_278);
and U56 (N_56,In_716,In_371);
nand U57 (N_57,In_1099,In_325);
nand U58 (N_58,In_104,In_1091);
nand U59 (N_59,In_1186,In_1061);
xor U60 (N_60,In_580,In_1108);
or U61 (N_61,In_748,In_732);
and U62 (N_62,In_651,In_533);
and U63 (N_63,In_566,In_822);
and U64 (N_64,In_849,In_1095);
and U65 (N_65,In_277,In_690);
xnor U66 (N_66,In_543,In_1009);
nor U67 (N_67,In_1402,In_452);
and U68 (N_68,In_586,In_920);
nand U69 (N_69,In_727,In_491);
and U70 (N_70,In_1432,In_1412);
nor U71 (N_71,In_1440,In_873);
nor U72 (N_72,In_269,In_774);
and U73 (N_73,In_1336,In_1194);
and U74 (N_74,In_1134,In_81);
nor U75 (N_75,In_1313,In_1263);
or U76 (N_76,In_854,In_1390);
and U77 (N_77,In_254,In_2);
or U78 (N_78,In_461,In_1127);
nand U79 (N_79,In_693,In_340);
nor U80 (N_80,In_430,In_758);
and U81 (N_81,In_584,In_1100);
nand U82 (N_82,In_1477,In_73);
and U83 (N_83,In_1136,In_96);
nor U84 (N_84,In_1475,In_815);
or U85 (N_85,In_1131,In_610);
and U86 (N_86,In_374,In_515);
nand U87 (N_87,In_628,In_1328);
nor U88 (N_88,In_1153,In_1064);
nand U89 (N_89,In_455,In_145);
or U90 (N_90,In_486,In_439);
or U91 (N_91,In_83,In_821);
or U92 (N_92,In_1032,In_307);
nor U93 (N_93,In_1035,In_710);
nor U94 (N_94,In_924,In_1042);
and U95 (N_95,In_292,In_1094);
and U96 (N_96,In_475,In_1202);
or U97 (N_97,In_1380,In_1383);
and U98 (N_98,In_1275,In_1459);
and U99 (N_99,In_833,In_351);
nor U100 (N_100,In_1014,In_1245);
nor U101 (N_101,In_1274,In_846);
and U102 (N_102,In_568,In_989);
or U103 (N_103,In_823,In_71);
or U104 (N_104,In_410,In_407);
xor U105 (N_105,In_233,In_1462);
or U106 (N_106,In_1102,In_1010);
and U107 (N_107,In_1096,In_1057);
nand U108 (N_108,In_1220,In_788);
nor U109 (N_109,In_1222,In_713);
or U110 (N_110,In_1417,In_505);
or U111 (N_111,In_332,In_612);
and U112 (N_112,In_851,In_671);
and U113 (N_113,In_1437,In_153);
nand U114 (N_114,In_1104,In_503);
nor U115 (N_115,In_52,In_304);
nor U116 (N_116,In_311,In_930);
or U117 (N_117,In_1154,In_1086);
or U118 (N_118,In_248,In_892);
nand U119 (N_119,In_883,In_1283);
or U120 (N_120,In_814,In_1286);
and U121 (N_121,In_965,In_927);
and U122 (N_122,In_776,In_1210);
or U123 (N_123,In_19,In_1138);
nor U124 (N_124,In_1244,In_835);
and U125 (N_125,In_1217,In_319);
nor U126 (N_126,In_582,In_1321);
and U127 (N_127,In_911,In_313);
and U128 (N_128,In_522,In_1146);
nand U129 (N_129,In_745,In_592);
and U130 (N_130,In_418,In_1428);
nand U131 (N_131,In_1080,In_441);
or U132 (N_132,In_1456,In_859);
and U133 (N_133,In_962,In_1498);
xor U134 (N_134,In_1007,In_697);
nor U135 (N_135,In_1158,In_1366);
xnor U136 (N_136,In_523,In_1199);
and U137 (N_137,In_449,In_1427);
nand U138 (N_138,In_225,In_162);
or U139 (N_139,In_228,In_1435);
xor U140 (N_140,In_202,In_717);
nand U141 (N_141,In_1125,In_482);
and U142 (N_142,In_1,In_321);
or U143 (N_143,In_567,In_715);
and U144 (N_144,In_1250,In_1157);
nor U145 (N_145,In_560,In_126);
nand U146 (N_146,In_536,In_63);
or U147 (N_147,In_286,In_676);
nor U148 (N_148,In_234,In_23);
nor U149 (N_149,In_1468,In_1395);
nor U150 (N_150,In_921,In_498);
or U151 (N_151,In_681,In_521);
or U152 (N_152,In_333,In_487);
xor U153 (N_153,In_70,In_1218);
xnor U154 (N_154,In_127,In_1101);
nand U155 (N_155,In_1103,In_288);
nor U156 (N_156,In_850,In_876);
nand U157 (N_157,In_1304,In_231);
and U158 (N_158,In_250,In_94);
or U159 (N_159,In_10,In_1284);
xnor U160 (N_160,In_722,In_905);
nand U161 (N_161,In_1271,In_1020);
nand U162 (N_162,In_513,In_624);
nor U163 (N_163,In_45,In_587);
nor U164 (N_164,In_317,In_1008);
or U165 (N_165,In_1480,In_326);
nor U166 (N_166,In_1438,In_92);
nor U167 (N_167,In_1130,In_1232);
and U168 (N_168,In_144,In_844);
nand U169 (N_169,In_200,In_440);
nand U170 (N_170,In_699,In_1087);
nand U171 (N_171,In_620,In_1122);
and U172 (N_172,In_878,In_644);
nor U173 (N_173,In_838,In_347);
nand U174 (N_174,In_1031,In_392);
xnor U175 (N_175,In_330,In_1041);
and U176 (N_176,In_589,In_537);
and U177 (N_177,In_272,In_1351);
nor U178 (N_178,In_1329,In_217);
or U179 (N_179,In_1170,In_1482);
and U180 (N_180,In_755,In_581);
xnor U181 (N_181,In_1325,In_479);
or U182 (N_182,In_7,In_763);
nor U183 (N_183,In_1419,In_805);
and U184 (N_184,In_1397,In_502);
and U185 (N_185,In_1295,In_203);
nand U186 (N_186,In_1270,In_1294);
or U187 (N_187,In_847,In_600);
xnor U188 (N_188,In_1107,In_664);
or U189 (N_189,In_672,In_558);
nor U190 (N_190,In_204,In_982);
nor U191 (N_191,In_926,In_456);
nor U192 (N_192,In_53,In_1110);
or U193 (N_193,In_386,In_1056);
nor U194 (N_194,In_826,In_1002);
and U195 (N_195,In_1205,In_695);
or U196 (N_196,In_861,In_362);
xor U197 (N_197,In_290,In_401);
or U198 (N_198,In_1078,In_1347);
nand U199 (N_199,In_310,In_1115);
nor U200 (N_200,In_159,In_358);
nand U201 (N_201,In_1463,In_149);
and U202 (N_202,In_673,In_28);
nand U203 (N_203,In_540,In_1376);
nor U204 (N_204,In_771,In_723);
nand U205 (N_205,In_1051,In_416);
and U206 (N_206,In_497,In_394);
xnor U207 (N_207,In_124,In_952);
and U208 (N_208,In_20,In_1369);
nand U209 (N_209,In_779,In_252);
nor U210 (N_210,In_214,In_1132);
nand U211 (N_211,In_1401,In_1072);
nor U212 (N_212,In_1109,In_1488);
xnor U213 (N_213,In_1393,In_561);
xnor U214 (N_214,In_1092,In_241);
and U215 (N_215,In_8,In_256);
nor U216 (N_216,In_1256,In_685);
xor U217 (N_217,In_431,In_1327);
or U218 (N_218,In_1389,In_557);
xnor U219 (N_219,In_934,In_575);
or U220 (N_220,In_728,In_725);
and U221 (N_221,In_504,In_785);
nand U222 (N_222,In_154,In_527);
and U223 (N_223,In_552,In_419);
nand U224 (N_224,In_229,In_947);
nand U225 (N_225,In_1142,In_443);
or U226 (N_226,In_135,In_608);
and U227 (N_227,In_174,In_897);
nand U228 (N_228,In_1416,In_1400);
nor U229 (N_229,In_1464,In_21);
nand U230 (N_230,In_1037,In_261);
and U231 (N_231,In_186,In_216);
and U232 (N_232,In_632,In_1490);
nor U233 (N_233,In_400,In_51);
nor U234 (N_234,In_1171,In_413);
or U235 (N_235,In_79,In_791);
nand U236 (N_236,In_142,In_1240);
or U237 (N_237,In_100,In_1167);
nor U238 (N_238,In_473,In_1215);
and U239 (N_239,In_1229,In_1024);
nand U240 (N_240,In_741,In_97);
or U241 (N_241,In_460,In_466);
xnor U242 (N_242,In_308,In_160);
or U243 (N_243,In_9,In_117);
nand U244 (N_244,In_1346,In_649);
or U245 (N_245,In_1180,In_187);
and U246 (N_246,In_1121,In_315);
nor U247 (N_247,In_738,In_331);
nand U248 (N_248,In_1373,In_1430);
xnor U249 (N_249,In_1299,In_47);
nor U250 (N_250,In_939,In_909);
nand U251 (N_251,In_1183,In_240);
and U252 (N_252,In_855,In_516);
nor U253 (N_253,In_1128,In_901);
and U254 (N_254,In_432,In_1422);
nand U255 (N_255,In_244,In_613);
or U256 (N_256,In_1161,In_434);
and U257 (N_257,In_1118,In_134);
xnor U258 (N_258,In_1331,In_147);
xor U259 (N_259,In_291,In_735);
or U260 (N_260,In_334,In_305);
or U261 (N_261,In_597,In_376);
xor U262 (N_262,In_556,In_488);
and U263 (N_263,In_743,In_871);
or U264 (N_264,In_1272,In_423);
and U265 (N_265,In_968,In_1474);
xnor U266 (N_266,In_571,In_1214);
nor U267 (N_267,In_427,In_843);
nand U268 (N_268,In_1106,In_856);
nand U269 (N_269,In_1173,In_809);
nor U270 (N_270,In_271,In_642);
and U271 (N_271,In_555,In_1404);
or U272 (N_272,In_1352,In_1185);
and U273 (N_273,In_62,In_877);
and U274 (N_274,In_891,In_631);
or U275 (N_275,In_1190,In_88);
nor U276 (N_276,In_633,In_1068);
xnor U277 (N_277,In_1266,In_1418);
xnor U278 (N_278,In_155,In_188);
xor U279 (N_279,In_559,In_1431);
nor U280 (N_280,In_798,In_377);
or U281 (N_281,In_975,In_226);
and U282 (N_282,In_1378,In_958);
or U283 (N_283,In_1409,In_235);
and U284 (N_284,In_603,In_573);
nor U285 (N_285,In_1381,In_1209);
or U286 (N_286,In_707,In_110);
nor U287 (N_287,In_1155,In_837);
xnor U288 (N_288,In_824,In_1040);
xnor U289 (N_289,In_1357,In_853);
or U290 (N_290,In_1461,In_596);
nor U291 (N_291,In_611,In_866);
or U292 (N_292,In_1140,In_266);
nor U293 (N_293,In_1398,In_60);
and U294 (N_294,In_622,In_1353);
and U295 (N_295,In_641,In_1273);
xor U296 (N_296,In_1059,In_1333);
or U297 (N_297,In_263,In_661);
nand U298 (N_298,In_886,In_1066);
nor U299 (N_299,In_141,In_687);
or U300 (N_300,In_1457,In_819);
nor U301 (N_301,In_1489,In_918);
nand U302 (N_302,In_114,In_50);
and U303 (N_303,In_1358,In_1034);
nand U304 (N_304,In_570,In_499);
xnor U305 (N_305,In_1043,In_535);
or U306 (N_306,In_795,In_509);
or U307 (N_307,In_260,In_1311);
and U308 (N_308,In_56,In_1258);
or U309 (N_309,In_282,In_1359);
or U310 (N_310,In_719,In_1143);
nand U311 (N_311,In_906,In_564);
nand U312 (N_312,In_82,In_289);
xnor U313 (N_313,In_1268,In_205);
nand U314 (N_314,In_1211,In_128);
or U315 (N_315,In_1297,In_253);
or U316 (N_316,In_818,In_1062);
nand U317 (N_317,In_804,In_1307);
or U318 (N_318,In_1442,In_1309);
or U319 (N_319,In_737,In_1387);
nor U320 (N_320,In_329,In_964);
nor U321 (N_321,In_1097,In_550);
and U322 (N_322,In_974,In_639);
or U323 (N_323,In_1340,In_1159);
or U324 (N_324,In_565,In_972);
and U325 (N_325,In_184,In_1163);
nor U326 (N_326,In_361,In_1470);
nand U327 (N_327,In_1446,In_1476);
or U328 (N_328,In_297,In_662);
nor U329 (N_329,In_6,In_506);
or U330 (N_330,In_1179,In_1288);
and U331 (N_331,In_274,In_369);
or U332 (N_332,In_1384,In_1133);
xnor U333 (N_333,In_784,In_1213);
nand U334 (N_334,In_655,In_1071);
nand U335 (N_335,In_199,In_181);
and U336 (N_336,In_1203,In_786);
nor U337 (N_337,In_708,In_1196);
nand U338 (N_338,In_796,In_1473);
or U339 (N_339,In_593,In_230);
or U340 (N_340,In_5,In_481);
nor U341 (N_341,In_669,In_222);
nor U342 (N_342,In_1291,In_1415);
and U343 (N_343,In_992,In_395);
or U344 (N_344,In_1499,In_869);
or U345 (N_345,In_1379,In_948);
and U346 (N_346,In_1223,In_1160);
nand U347 (N_347,In_30,In_1172);
and U348 (N_348,In_1151,In_730);
or U349 (N_349,In_415,In_946);
or U350 (N_350,In_652,In_345);
nor U351 (N_351,In_137,In_1077);
or U352 (N_352,In_3,In_700);
and U353 (N_353,In_1063,In_138);
and U354 (N_354,In_459,In_109);
or U355 (N_355,In_470,In_437);
or U356 (N_356,In_1221,In_336);
or U357 (N_357,In_287,In_295);
and U358 (N_358,In_1181,In_1269);
nor U359 (N_359,In_764,In_882);
nor U360 (N_360,In_380,In_528);
or U361 (N_361,In_55,In_1039);
and U362 (N_362,In_1486,In_1197);
nand U363 (N_363,In_963,In_1184);
and U364 (N_364,In_477,In_1375);
nand U365 (N_365,In_842,In_1135);
nand U366 (N_366,In_684,In_1334);
and U367 (N_367,In_169,In_967);
and U368 (N_368,In_890,In_381);
nand U369 (N_369,In_465,In_797);
nor U370 (N_370,In_1018,In_751);
and U371 (N_371,In_312,In_1259);
nor U372 (N_372,In_950,In_1028);
nor U373 (N_373,In_977,In_731);
and U374 (N_374,In_26,In_686);
and U375 (N_375,In_102,In_1305);
xnor U376 (N_376,In_945,In_1368);
nand U377 (N_377,In_84,In_91);
xor U378 (N_378,In_341,In_820);
nor U379 (N_379,In_817,In_894);
or U380 (N_380,In_116,In_283);
xor U381 (N_381,In_501,In_1162);
xor U382 (N_382,In_206,In_1081);
nor U383 (N_383,In_178,In_85);
nor U384 (N_384,In_1105,In_1433);
nor U385 (N_385,In_17,In_635);
and U386 (N_386,In_151,In_1436);
or U387 (N_387,In_354,In_1385);
nor U388 (N_388,In_985,In_46);
xor U389 (N_389,In_406,In_399);
and U390 (N_390,In_1314,In_973);
nand U391 (N_391,In_492,In_1241);
xnor U392 (N_392,In_1455,In_1332);
or U393 (N_393,In_1296,In_1348);
xnor U394 (N_394,In_667,In_609);
nor U395 (N_395,In_238,In_469);
nand U396 (N_396,In_384,In_960);
and U397 (N_397,In_98,In_1058);
and U398 (N_398,In_1495,In_813);
or U399 (N_399,In_1371,In_1123);
and U400 (N_400,In_220,In_1405);
or U401 (N_401,In_1382,In_29);
or U402 (N_402,In_1342,In_760);
xnor U403 (N_403,In_285,In_1248);
nor U404 (N_404,In_1301,In_606);
or U405 (N_405,In_834,In_683);
xor U406 (N_406,In_675,In_40);
nor U407 (N_407,In_490,In_1207);
nand U408 (N_408,In_595,In_425);
nand U409 (N_409,In_529,In_1208);
nand U410 (N_410,In_41,In_1413);
or U411 (N_411,In_1147,In_408);
or U412 (N_412,In_1277,In_75);
nor U413 (N_413,In_829,In_753);
or U414 (N_414,In_500,In_1339);
or U415 (N_415,In_414,In_1388);
nor U416 (N_416,In_761,In_176);
nor U417 (N_417,In_18,In_320);
nor U418 (N_418,In_382,In_1046);
or U419 (N_419,In_299,In_209);
nor U420 (N_420,In_211,In_526);
and U421 (N_421,In_790,In_893);
nor U422 (N_422,In_177,In_424);
and U423 (N_423,In_643,In_778);
and U424 (N_424,In_33,In_1361);
or U425 (N_425,In_212,In_1191);
and U426 (N_426,In_136,In_616);
nor U427 (N_427,In_146,In_396);
xnor U428 (N_428,In_990,In_420);
nand U429 (N_429,In_167,In_1493);
and U430 (N_430,In_300,In_808);
nor U431 (N_431,In_335,In_1187);
xor U432 (N_432,In_1324,In_511);
nor U433 (N_433,In_316,In_703);
and U434 (N_434,In_1204,In_507);
xnor U435 (N_435,In_1164,In_1224);
nor U436 (N_436,In_981,In_1414);
nor U437 (N_437,In_412,In_198);
nor U438 (N_438,In_1126,In_765);
or U439 (N_439,In_1047,In_769);
and U440 (N_440,In_698,In_617);
nor U441 (N_441,In_615,In_388);
and U442 (N_442,In_734,In_66);
or U443 (N_443,In_265,In_1093);
nor U444 (N_444,In_1065,In_880);
or U445 (N_445,In_1374,In_1454);
or U446 (N_446,In_1243,In_489);
xor U447 (N_447,In_553,In_458);
and U448 (N_448,In_1200,In_656);
or U449 (N_449,In_298,In_1227);
and U450 (N_450,In_125,In_706);
and U451 (N_451,In_157,In_378);
or U452 (N_452,In_1025,In_322);
xor U453 (N_453,In_807,In_1335);
or U454 (N_454,In_36,In_547);
nor U455 (N_455,In_1090,In_665);
nor U456 (N_456,In_984,In_421);
or U457 (N_457,In_344,In_1290);
and U458 (N_458,In_12,In_576);
xnor U459 (N_459,In_464,In_14);
and U460 (N_460,In_1189,In_726);
nand U461 (N_461,In_1033,In_262);
and U462 (N_462,In_363,In_907);
and U463 (N_463,In_1098,In_1483);
or U464 (N_464,In_77,In_1408);
and U465 (N_465,In_944,In_268);
or U466 (N_466,In_1038,In_1312);
nor U467 (N_467,In_1487,In_357);
and U468 (N_468,In_991,In_996);
and U469 (N_469,In_1302,In_379);
or U470 (N_470,In_712,In_742);
and U471 (N_471,In_32,In_447);
or U472 (N_472,In_409,In_1386);
xnor U473 (N_473,In_1156,In_862);
xor U474 (N_474,In_689,In_577);
or U475 (N_475,In_759,In_636);
nor U476 (N_476,In_121,In_1177);
nor U477 (N_477,In_746,In_1235);
and U478 (N_478,In_1168,In_875);
nand U479 (N_479,In_1228,In_747);
or U480 (N_480,In_1049,In_375);
nor U481 (N_481,In_539,In_1216);
xor U482 (N_482,In_1350,In_966);
xor U483 (N_483,In_1253,In_640);
nand U484 (N_484,In_1303,In_995);
and U485 (N_485,In_448,In_158);
xnor U486 (N_486,In_484,In_563);
and U487 (N_487,In_630,In_1152);
and U488 (N_488,In_619,In_101);
and U489 (N_489,In_89,In_599);
xor U490 (N_490,In_1377,In_825);
nor U491 (N_491,In_1201,In_249);
nand U492 (N_492,In_1279,In_1013);
or U493 (N_493,In_442,In_711);
nand U494 (N_494,In_997,In_267);
and U495 (N_495,In_1349,In_457);
nand U496 (N_496,In_534,In_393);
or U497 (N_497,In_1055,In_634);
and U498 (N_498,In_1372,In_113);
nand U499 (N_499,In_720,In_1254);
nand U500 (N_500,In_1212,In_925);
nor U501 (N_501,In_323,In_701);
nand U502 (N_502,In_658,In_35);
xnor U503 (N_503,In_175,In_197);
or U504 (N_504,In_402,In_1219);
and U505 (N_505,In_931,In_1452);
or U506 (N_506,In_1293,In_239);
nor U507 (N_507,In_1174,In_1421);
nand U508 (N_508,In_1257,In_663);
nor U509 (N_509,In_1392,In_899);
nor U510 (N_510,In_270,In_195);
xnor U511 (N_511,In_476,In_598);
and U512 (N_512,In_132,In_768);
xor U513 (N_513,In_152,In_954);
and U514 (N_514,In_496,In_405);
and U515 (N_515,In_95,In_213);
nor U516 (N_516,In_218,In_445);
or U517 (N_517,In_328,In_1193);
or U518 (N_518,In_1150,In_1429);
xor U519 (N_519,In_1298,In_841);
nor U520 (N_520,In_980,In_919);
or U521 (N_521,In_90,In_802);
xnor U522 (N_522,In_1320,In_1485);
or U523 (N_523,In_545,In_721);
and U524 (N_524,In_546,In_227);
nand U525 (N_525,In_1396,In_783);
nand U526 (N_526,In_359,In_1306);
nor U527 (N_527,In_1280,In_811);
or U528 (N_528,In_1076,In_327);
nor U529 (N_529,In_78,In_1341);
and U530 (N_530,In_803,In_355);
nor U531 (N_531,In_451,In_590);
and U532 (N_532,In_161,In_24);
or U533 (N_533,In_538,In_739);
nor U534 (N_534,In_349,In_858);
or U535 (N_535,In_583,In_895);
nor U536 (N_536,In_1262,In_709);
or U537 (N_537,In_1264,In_1444);
and U538 (N_538,In_1022,In_961);
or U539 (N_539,In_1231,In_530);
nand U540 (N_540,In_446,In_224);
nor U541 (N_541,In_182,In_1249);
nor U542 (N_542,In_367,In_627);
nor U543 (N_543,In_1281,In_385);
xnor U544 (N_544,In_1112,In_1027);
nand U545 (N_545,In_1497,In_767);
and U546 (N_546,In_428,In_436);
nand U547 (N_547,In_383,In_957);
nand U548 (N_548,In_183,In_391);
xor U549 (N_549,In_1439,In_1425);
nor U550 (N_550,In_621,In_884);
nand U551 (N_551,In_370,In_44);
nand U552 (N_552,In_780,In_131);
nand U553 (N_553,In_1252,In_549);
and U554 (N_554,In_902,In_936);
and U555 (N_555,In_831,In_193);
xnor U556 (N_556,In_1114,In_998);
and U557 (N_557,In_626,In_532);
nand U558 (N_558,In_912,In_605);
or U559 (N_559,In_682,In_848);
nand U560 (N_560,In_1496,In_903);
and U561 (N_561,In_691,In_789);
and U562 (N_562,In_454,In_368);
nor U563 (N_563,In_810,In_601);
nor U564 (N_564,In_799,In_68);
nor U565 (N_565,In_569,In_163);
xnor U566 (N_566,In_932,In_1403);
or U567 (N_567,In_544,In_524);
or U568 (N_568,In_836,In_191);
nor U569 (N_569,In_852,In_302);
nor U570 (N_570,In_1354,In_171);
and U571 (N_571,In_1394,In_112);
and U572 (N_572,In_80,In_970);
nand U573 (N_573,In_494,In_324);
nor U574 (N_574,In_1236,In_660);
or U575 (N_575,In_772,In_1411);
nor U576 (N_576,In_180,In_485);
or U577 (N_577,In_915,In_404);
nor U578 (N_578,In_937,In_647);
and U579 (N_579,In_1448,In_874);
nand U580 (N_580,In_236,In_48);
or U581 (N_581,In_1084,In_54);
and U582 (N_582,In_348,In_940);
and U583 (N_583,In_750,In_923);
nand U584 (N_584,In_221,In_910);
or U585 (N_585,In_1067,In_309);
and U586 (N_586,In_1434,In_956);
nor U587 (N_587,In_718,In_190);
xnor U588 (N_588,In_749,In_108);
and U589 (N_589,In_752,In_832);
xor U590 (N_590,In_450,In_1282);
nor U591 (N_591,In_1265,In_463);
and U592 (N_592,In_900,In_338);
and U593 (N_593,In_1026,In_133);
nand U594 (N_594,In_1001,In_864);
nor U595 (N_595,In_680,In_951);
nor U596 (N_596,In_365,In_1089);
xnor U597 (N_597,In_872,In_215);
nor U598 (N_598,In_714,In_574);
nor U599 (N_599,In_257,In_519);
nand U600 (N_600,In_1242,In_111);
and U601 (N_601,In_86,In_1141);
and U602 (N_602,In_694,In_107);
nand U603 (N_603,In_904,In_13);
xor U604 (N_604,In_987,In_259);
xnor U605 (N_605,In_493,In_189);
and U606 (N_606,In_801,In_922);
nand U607 (N_607,In_1230,In_1367);
nand U608 (N_608,In_1074,In_885);
and U609 (N_609,In_360,In_281);
and U610 (N_610,In_591,In_303);
or U611 (N_611,In_1000,In_943);
or U612 (N_612,In_1052,In_840);
nand U613 (N_613,In_422,In_1472);
and U614 (N_614,In_637,In_913);
or U615 (N_615,In_1017,In_294);
and U616 (N_616,In_306,In_917);
xnor U617 (N_617,In_1330,In_255);
nand U618 (N_618,In_397,In_959);
nor U619 (N_619,In_61,In_57);
or U620 (N_620,In_398,In_1044);
or U621 (N_621,In_638,In_472);
and U622 (N_622,In_756,In_1169);
and U623 (N_623,In_517,In_275);
and U624 (N_624,In_978,In_1362);
and U625 (N_625,In_740,In_1145);
and U626 (N_626,In_411,In_929);
nor U627 (N_627,In_372,In_179);
and U628 (N_628,In_562,In_578);
nand U629 (N_629,In_828,In_208);
or U630 (N_630,In_207,In_246);
nand U631 (N_631,In_366,In_993);
and U632 (N_632,In_467,In_1178);
nand U633 (N_633,In_1085,In_1016);
nor U634 (N_634,In_602,In_704);
and U635 (N_635,In_237,In_38);
nand U636 (N_636,In_666,In_733);
nand U637 (N_637,In_1355,In_314);
nor U638 (N_638,In_164,In_1139);
or U639 (N_639,In_99,In_242);
nor U640 (N_640,In_76,In_353);
and U641 (N_641,In_129,In_1467);
and U642 (N_642,In_1188,In_22);
nand U643 (N_643,In_115,In_510);
xnor U644 (N_644,In_762,In_103);
and U645 (N_645,In_478,In_39);
nand U646 (N_646,In_648,In_67);
nand U647 (N_647,In_705,In_1006);
and U648 (N_648,In_1233,In_736);
nand U649 (N_649,In_279,In_123);
nand U650 (N_650,In_949,In_373);
nand U651 (N_651,In_1420,In_782);
nand U652 (N_652,In_1410,In_1045);
nor U653 (N_653,In_1050,In_514);
nand U654 (N_654,In_118,In_1278);
and U655 (N_655,In_1391,In_165);
nand U656 (N_656,In_1494,In_724);
or U657 (N_657,In_1004,In_668);
and U658 (N_658,In_27,In_816);
nor U659 (N_659,In_657,In_1144);
or U660 (N_660,In_1479,In_692);
xor U661 (N_661,In_1360,In_1070);
or U662 (N_662,In_983,In_806);
nor U663 (N_663,In_800,In_37);
or U664 (N_664,In_350,In_928);
nor U665 (N_665,In_1458,In_251);
xnor U666 (N_666,In_122,In_508);
nand U667 (N_667,In_276,In_679);
and U668 (N_668,In_1246,In_1344);
nand U669 (N_669,In_106,In_1251);
and U670 (N_670,In_1119,In_677);
and U671 (N_671,In_1198,In_1343);
and U672 (N_672,In_168,In_1407);
nand U673 (N_673,In_364,In_468);
or U674 (N_674,In_518,In_618);
or U675 (N_675,In_525,In_273);
and U676 (N_676,In_232,In_49);
nor U677 (N_677,In_614,In_462);
nand U678 (N_678,In_34,In_11);
nand U679 (N_679,In_438,In_865);
and U680 (N_680,In_1460,In_223);
and U681 (N_681,In_1365,In_1060);
nand U682 (N_682,In_301,In_192);
nand U683 (N_683,In_986,In_219);
or U684 (N_684,In_139,In_868);
nand U685 (N_685,In_1195,In_343);
xnor U686 (N_686,In_889,In_520);
nor U687 (N_687,In_105,In_280);
xor U688 (N_688,In_777,In_264);
or U689 (N_689,In_1356,In_863);
and U690 (N_690,In_623,In_93);
and U691 (N_691,In_1471,In_1445);
nand U692 (N_692,In_757,In_988);
nor U693 (N_693,In_258,In_346);
and U694 (N_694,In_1316,In_1323);
xnor U695 (N_695,In_770,In_426);
nand U696 (N_696,In_1424,In_4);
nand U697 (N_697,In_773,In_1443);
and U698 (N_698,In_845,In_830);
nor U699 (N_699,In_1073,In_403);
nor U700 (N_700,In_867,In_888);
and U701 (N_701,In_1300,In_781);
or U702 (N_702,In_1117,In_1441);
and U703 (N_703,In_594,In_1116);
nand U704 (N_704,In_130,In_1267);
and U705 (N_705,In_1120,In_201);
or U706 (N_706,In_1315,In_1465);
or U707 (N_707,In_702,In_794);
and U708 (N_708,In_1276,In_15);
xor U709 (N_709,In_1137,In_58);
xor U710 (N_710,In_896,In_914);
xor U711 (N_711,In_1287,In_678);
xor U712 (N_712,In_572,In_352);
and U713 (N_713,In_1399,In_1345);
or U714 (N_714,In_247,In_969);
and U715 (N_715,In_342,In_1449);
xor U716 (N_716,In_1492,In_881);
xor U717 (N_717,In_1088,In_43);
nand U718 (N_718,In_1318,In_453);
or U719 (N_719,In_554,In_908);
nand U720 (N_720,In_65,In_471);
and U721 (N_721,In_1338,In_1317);
nand U722 (N_722,In_1363,In_417);
xor U723 (N_723,In_1011,In_1478);
and U724 (N_724,In_1192,In_531);
nor U725 (N_725,In_1003,In_1260);
or U726 (N_726,In_1176,In_1310);
nand U727 (N_727,In_337,In_140);
and U728 (N_728,In_0,In_898);
or U729 (N_729,In_356,In_942);
xor U730 (N_730,In_1048,In_1423);
or U731 (N_731,In_1005,In_744);
or U732 (N_732,In_793,In_953);
nor U733 (N_733,In_1234,In_435);
nor U734 (N_734,In_787,In_59);
nand U735 (N_735,In_994,In_1129);
and U736 (N_736,In_1012,In_284);
nand U737 (N_737,In_629,In_548);
nor U738 (N_738,In_243,In_1054);
nand U739 (N_739,In_659,In_474);
nand U740 (N_740,In_16,In_653);
nor U741 (N_741,In_210,In_1453);
or U742 (N_742,In_645,In_173);
nand U743 (N_743,In_955,In_1308);
nand U744 (N_744,In_495,In_839);
nand U745 (N_745,In_999,In_916);
or U746 (N_746,In_1364,In_1113);
or U747 (N_747,In_318,In_1149);
nor U748 (N_748,In_31,In_293);
xnor U749 (N_749,In_650,In_1069);
nor U750 (N_750,In_516,In_239);
or U751 (N_751,In_165,In_737);
and U752 (N_752,In_1043,In_279);
or U753 (N_753,In_1297,In_185);
nor U754 (N_754,In_1442,In_1083);
or U755 (N_755,In_1303,In_84);
or U756 (N_756,In_1081,In_1469);
or U757 (N_757,In_1467,In_492);
nand U758 (N_758,In_410,In_919);
or U759 (N_759,In_1035,In_503);
or U760 (N_760,In_1058,In_1466);
and U761 (N_761,In_62,In_654);
nor U762 (N_762,In_805,In_244);
nand U763 (N_763,In_1197,In_1388);
and U764 (N_764,In_689,In_1035);
nor U765 (N_765,In_987,In_1337);
nor U766 (N_766,In_1124,In_1296);
and U767 (N_767,In_295,In_1055);
nand U768 (N_768,In_1418,In_882);
nor U769 (N_769,In_539,In_789);
nand U770 (N_770,In_516,In_925);
nand U771 (N_771,In_280,In_982);
and U772 (N_772,In_1366,In_132);
or U773 (N_773,In_301,In_879);
xor U774 (N_774,In_130,In_1435);
or U775 (N_775,In_467,In_59);
nand U776 (N_776,In_1304,In_1196);
or U777 (N_777,In_956,In_1253);
or U778 (N_778,In_662,In_23);
and U779 (N_779,In_678,In_265);
or U780 (N_780,In_1132,In_1441);
nand U781 (N_781,In_733,In_696);
or U782 (N_782,In_1116,In_773);
nor U783 (N_783,In_1293,In_1408);
nand U784 (N_784,In_997,In_1332);
nand U785 (N_785,In_1186,In_399);
or U786 (N_786,In_1186,In_1195);
and U787 (N_787,In_1248,In_15);
or U788 (N_788,In_888,In_407);
and U789 (N_789,In_1010,In_1238);
and U790 (N_790,In_1346,In_379);
nand U791 (N_791,In_730,In_74);
and U792 (N_792,In_1100,In_1428);
or U793 (N_793,In_854,In_485);
nor U794 (N_794,In_138,In_847);
nor U795 (N_795,In_743,In_940);
or U796 (N_796,In_1216,In_119);
nor U797 (N_797,In_501,In_1076);
and U798 (N_798,In_214,In_501);
nor U799 (N_799,In_897,In_377);
or U800 (N_800,In_1042,In_363);
and U801 (N_801,In_508,In_1266);
nor U802 (N_802,In_1319,In_1155);
or U803 (N_803,In_224,In_1472);
or U804 (N_804,In_1196,In_1207);
nor U805 (N_805,In_1277,In_34);
nand U806 (N_806,In_650,In_112);
and U807 (N_807,In_1405,In_449);
nand U808 (N_808,In_339,In_724);
or U809 (N_809,In_461,In_1462);
nand U810 (N_810,In_415,In_596);
nand U811 (N_811,In_1130,In_546);
or U812 (N_812,In_528,In_878);
nor U813 (N_813,In_221,In_659);
nand U814 (N_814,In_812,In_190);
or U815 (N_815,In_89,In_100);
nor U816 (N_816,In_410,In_258);
and U817 (N_817,In_1372,In_968);
nand U818 (N_818,In_125,In_428);
nand U819 (N_819,In_903,In_1454);
nor U820 (N_820,In_1438,In_353);
nor U821 (N_821,In_430,In_283);
and U822 (N_822,In_895,In_1062);
nor U823 (N_823,In_646,In_1257);
or U824 (N_824,In_926,In_512);
and U825 (N_825,In_1442,In_778);
xor U826 (N_826,In_231,In_1072);
or U827 (N_827,In_1418,In_21);
or U828 (N_828,In_883,In_1449);
nand U829 (N_829,In_431,In_619);
nand U830 (N_830,In_340,In_890);
and U831 (N_831,In_918,In_265);
nor U832 (N_832,In_197,In_378);
and U833 (N_833,In_997,In_145);
and U834 (N_834,In_1260,In_1107);
and U835 (N_835,In_1451,In_744);
xnor U836 (N_836,In_970,In_366);
and U837 (N_837,In_530,In_119);
and U838 (N_838,In_550,In_744);
nand U839 (N_839,In_674,In_578);
nor U840 (N_840,In_1484,In_852);
or U841 (N_841,In_1457,In_386);
or U842 (N_842,In_1019,In_195);
or U843 (N_843,In_841,In_1364);
nand U844 (N_844,In_510,In_452);
or U845 (N_845,In_599,In_1451);
or U846 (N_846,In_1467,In_1227);
nor U847 (N_847,In_929,In_1184);
nand U848 (N_848,In_225,In_1492);
and U849 (N_849,In_804,In_770);
nand U850 (N_850,In_1031,In_243);
or U851 (N_851,In_459,In_201);
or U852 (N_852,In_602,In_189);
and U853 (N_853,In_1483,In_42);
and U854 (N_854,In_32,In_56);
nand U855 (N_855,In_1153,In_1256);
nor U856 (N_856,In_981,In_1124);
nor U857 (N_857,In_968,In_1048);
nand U858 (N_858,In_1442,In_421);
nor U859 (N_859,In_271,In_880);
and U860 (N_860,In_285,In_1467);
xnor U861 (N_861,In_413,In_744);
xor U862 (N_862,In_1228,In_1314);
or U863 (N_863,In_610,In_161);
nand U864 (N_864,In_359,In_952);
nor U865 (N_865,In_834,In_136);
nand U866 (N_866,In_719,In_292);
nor U867 (N_867,In_420,In_741);
xor U868 (N_868,In_1242,In_1377);
nand U869 (N_869,In_662,In_1456);
nand U870 (N_870,In_1229,In_918);
and U871 (N_871,In_933,In_1192);
nor U872 (N_872,In_1332,In_1028);
xor U873 (N_873,In_633,In_647);
or U874 (N_874,In_1194,In_1185);
and U875 (N_875,In_408,In_538);
xor U876 (N_876,In_16,In_1134);
nor U877 (N_877,In_206,In_1348);
or U878 (N_878,In_1454,In_539);
or U879 (N_879,In_1420,In_1101);
nand U880 (N_880,In_249,In_48);
or U881 (N_881,In_380,In_873);
xnor U882 (N_882,In_573,In_845);
and U883 (N_883,In_511,In_558);
or U884 (N_884,In_1262,In_180);
nand U885 (N_885,In_1080,In_1077);
and U886 (N_886,In_433,In_1433);
nor U887 (N_887,In_756,In_1223);
nor U888 (N_888,In_1441,In_1216);
nor U889 (N_889,In_634,In_1401);
and U890 (N_890,In_732,In_648);
and U891 (N_891,In_505,In_231);
or U892 (N_892,In_1397,In_72);
or U893 (N_893,In_960,In_1340);
or U894 (N_894,In_141,In_729);
or U895 (N_895,In_1126,In_381);
nor U896 (N_896,In_1096,In_1317);
nand U897 (N_897,In_282,In_915);
and U898 (N_898,In_1352,In_0);
xor U899 (N_899,In_790,In_61);
or U900 (N_900,In_938,In_682);
and U901 (N_901,In_1242,In_91);
or U902 (N_902,In_410,In_859);
xnor U903 (N_903,In_304,In_765);
nor U904 (N_904,In_640,In_952);
nor U905 (N_905,In_1038,In_229);
nand U906 (N_906,In_304,In_910);
or U907 (N_907,In_1273,In_418);
xor U908 (N_908,In_28,In_1030);
and U909 (N_909,In_1141,In_62);
nand U910 (N_910,In_769,In_762);
nand U911 (N_911,In_752,In_999);
or U912 (N_912,In_138,In_1077);
or U913 (N_913,In_100,In_694);
nand U914 (N_914,In_1449,In_108);
and U915 (N_915,In_54,In_221);
xor U916 (N_916,In_97,In_512);
and U917 (N_917,In_521,In_138);
nand U918 (N_918,In_473,In_959);
or U919 (N_919,In_975,In_156);
nor U920 (N_920,In_731,In_821);
nor U921 (N_921,In_713,In_1);
nor U922 (N_922,In_201,In_1127);
and U923 (N_923,In_841,In_1272);
nor U924 (N_924,In_243,In_413);
or U925 (N_925,In_801,In_1346);
xor U926 (N_926,In_786,In_677);
xor U927 (N_927,In_885,In_807);
or U928 (N_928,In_694,In_545);
xnor U929 (N_929,In_1014,In_689);
nand U930 (N_930,In_201,In_970);
nor U931 (N_931,In_1033,In_443);
and U932 (N_932,In_910,In_1264);
nand U933 (N_933,In_1200,In_588);
and U934 (N_934,In_548,In_293);
and U935 (N_935,In_373,In_1307);
nor U936 (N_936,In_435,In_164);
nand U937 (N_937,In_662,In_1060);
nand U938 (N_938,In_281,In_28);
nand U939 (N_939,In_989,In_1417);
or U940 (N_940,In_366,In_1152);
or U941 (N_941,In_462,In_65);
nor U942 (N_942,In_719,In_582);
xnor U943 (N_943,In_46,In_807);
xor U944 (N_944,In_512,In_1006);
nand U945 (N_945,In_945,In_1378);
or U946 (N_946,In_348,In_681);
nor U947 (N_947,In_216,In_1277);
nand U948 (N_948,In_911,In_475);
and U949 (N_949,In_949,In_59);
and U950 (N_950,In_1377,In_939);
nand U951 (N_951,In_106,In_354);
nand U952 (N_952,In_320,In_690);
xor U953 (N_953,In_581,In_1242);
nor U954 (N_954,In_839,In_291);
nand U955 (N_955,In_1029,In_1041);
nand U956 (N_956,In_1132,In_184);
or U957 (N_957,In_809,In_1005);
or U958 (N_958,In_1054,In_558);
and U959 (N_959,In_907,In_669);
nor U960 (N_960,In_1156,In_413);
nor U961 (N_961,In_458,In_375);
nand U962 (N_962,In_1202,In_703);
nor U963 (N_963,In_851,In_1464);
nand U964 (N_964,In_526,In_600);
nand U965 (N_965,In_141,In_1213);
xor U966 (N_966,In_38,In_106);
or U967 (N_967,In_1199,In_15);
nor U968 (N_968,In_284,In_729);
and U969 (N_969,In_1241,In_899);
xnor U970 (N_970,In_548,In_485);
or U971 (N_971,In_1087,In_1349);
and U972 (N_972,In_685,In_1097);
xnor U973 (N_973,In_16,In_22);
nand U974 (N_974,In_903,In_406);
xor U975 (N_975,In_155,In_1139);
nor U976 (N_976,In_130,In_494);
or U977 (N_977,In_570,In_72);
nand U978 (N_978,In_590,In_1394);
nor U979 (N_979,In_1366,In_145);
nand U980 (N_980,In_188,In_173);
nor U981 (N_981,In_965,In_1154);
or U982 (N_982,In_373,In_484);
nor U983 (N_983,In_1442,In_987);
or U984 (N_984,In_339,In_981);
or U985 (N_985,In_684,In_569);
nand U986 (N_986,In_1224,In_590);
nand U987 (N_987,In_1440,In_1046);
or U988 (N_988,In_908,In_1160);
nand U989 (N_989,In_240,In_834);
or U990 (N_990,In_929,In_1059);
nand U991 (N_991,In_1388,In_793);
nor U992 (N_992,In_1199,In_80);
nor U993 (N_993,In_557,In_1410);
nor U994 (N_994,In_434,In_176);
nor U995 (N_995,In_1031,In_551);
xor U996 (N_996,In_691,In_809);
and U997 (N_997,In_998,In_406);
nor U998 (N_998,In_303,In_194);
nor U999 (N_999,In_307,In_956);
nand U1000 (N_1000,In_1326,In_758);
or U1001 (N_1001,In_300,In_1078);
nor U1002 (N_1002,In_306,In_609);
or U1003 (N_1003,In_1130,In_719);
or U1004 (N_1004,In_762,In_1289);
nand U1005 (N_1005,In_92,In_858);
and U1006 (N_1006,In_1251,In_165);
and U1007 (N_1007,In_1496,In_889);
nor U1008 (N_1008,In_819,In_466);
nor U1009 (N_1009,In_150,In_175);
nand U1010 (N_1010,In_242,In_498);
nand U1011 (N_1011,In_698,In_643);
nand U1012 (N_1012,In_800,In_1135);
and U1013 (N_1013,In_349,In_766);
nand U1014 (N_1014,In_895,In_381);
nand U1015 (N_1015,In_528,In_754);
and U1016 (N_1016,In_354,In_805);
and U1017 (N_1017,In_673,In_1061);
nand U1018 (N_1018,In_392,In_1115);
nand U1019 (N_1019,In_1225,In_1223);
and U1020 (N_1020,In_307,In_814);
and U1021 (N_1021,In_810,In_1406);
nor U1022 (N_1022,In_116,In_414);
or U1023 (N_1023,In_410,In_399);
nor U1024 (N_1024,In_1206,In_1386);
nand U1025 (N_1025,In_962,In_1358);
or U1026 (N_1026,In_438,In_1045);
nand U1027 (N_1027,In_243,In_429);
nand U1028 (N_1028,In_84,In_1240);
and U1029 (N_1029,In_127,In_1179);
and U1030 (N_1030,In_733,In_681);
nor U1031 (N_1031,In_161,In_537);
and U1032 (N_1032,In_583,In_215);
nand U1033 (N_1033,In_1469,In_1093);
nor U1034 (N_1034,In_532,In_1373);
or U1035 (N_1035,In_481,In_195);
or U1036 (N_1036,In_1406,In_184);
or U1037 (N_1037,In_1260,In_843);
nor U1038 (N_1038,In_800,In_761);
and U1039 (N_1039,In_1116,In_1089);
and U1040 (N_1040,In_101,In_213);
and U1041 (N_1041,In_328,In_1410);
nand U1042 (N_1042,In_1393,In_1469);
or U1043 (N_1043,In_1039,In_54);
nand U1044 (N_1044,In_684,In_281);
or U1045 (N_1045,In_323,In_1096);
nand U1046 (N_1046,In_784,In_1252);
nor U1047 (N_1047,In_955,In_75);
or U1048 (N_1048,In_1425,In_1336);
xor U1049 (N_1049,In_292,In_609);
or U1050 (N_1050,In_1054,In_292);
or U1051 (N_1051,In_1073,In_709);
or U1052 (N_1052,In_1451,In_543);
and U1053 (N_1053,In_240,In_5);
nand U1054 (N_1054,In_540,In_377);
nor U1055 (N_1055,In_168,In_1022);
and U1056 (N_1056,In_1361,In_196);
or U1057 (N_1057,In_104,In_617);
and U1058 (N_1058,In_285,In_484);
and U1059 (N_1059,In_450,In_1025);
or U1060 (N_1060,In_359,In_421);
nor U1061 (N_1061,In_629,In_606);
and U1062 (N_1062,In_1307,In_126);
nor U1063 (N_1063,In_1451,In_308);
or U1064 (N_1064,In_1026,In_1296);
nor U1065 (N_1065,In_616,In_892);
nand U1066 (N_1066,In_177,In_492);
nor U1067 (N_1067,In_818,In_228);
xor U1068 (N_1068,In_451,In_424);
nand U1069 (N_1069,In_943,In_1044);
nor U1070 (N_1070,In_576,In_147);
nand U1071 (N_1071,In_953,In_1349);
nand U1072 (N_1072,In_531,In_718);
and U1073 (N_1073,In_303,In_501);
and U1074 (N_1074,In_161,In_1396);
or U1075 (N_1075,In_548,In_1403);
nor U1076 (N_1076,In_561,In_302);
nor U1077 (N_1077,In_179,In_425);
nand U1078 (N_1078,In_365,In_241);
and U1079 (N_1079,In_50,In_1203);
nand U1080 (N_1080,In_184,In_648);
and U1081 (N_1081,In_110,In_830);
or U1082 (N_1082,In_1205,In_381);
nand U1083 (N_1083,In_1266,In_567);
nor U1084 (N_1084,In_1162,In_227);
nor U1085 (N_1085,In_241,In_1210);
and U1086 (N_1086,In_1305,In_389);
xor U1087 (N_1087,In_483,In_482);
nor U1088 (N_1088,In_1250,In_821);
nor U1089 (N_1089,In_1034,In_705);
or U1090 (N_1090,In_1481,In_131);
and U1091 (N_1091,In_410,In_681);
and U1092 (N_1092,In_1229,In_798);
or U1093 (N_1093,In_731,In_544);
or U1094 (N_1094,In_1196,In_1499);
and U1095 (N_1095,In_1364,In_1470);
nand U1096 (N_1096,In_698,In_688);
xnor U1097 (N_1097,In_1206,In_222);
and U1098 (N_1098,In_1094,In_793);
and U1099 (N_1099,In_965,In_964);
nor U1100 (N_1100,In_431,In_1162);
or U1101 (N_1101,In_1431,In_1484);
nand U1102 (N_1102,In_866,In_1097);
or U1103 (N_1103,In_533,In_851);
or U1104 (N_1104,In_843,In_1020);
nand U1105 (N_1105,In_1218,In_747);
nand U1106 (N_1106,In_1094,In_1373);
nor U1107 (N_1107,In_1082,In_745);
or U1108 (N_1108,In_574,In_688);
nand U1109 (N_1109,In_740,In_519);
nor U1110 (N_1110,In_474,In_1147);
nor U1111 (N_1111,In_539,In_482);
nand U1112 (N_1112,In_907,In_777);
nor U1113 (N_1113,In_471,In_881);
and U1114 (N_1114,In_581,In_1129);
or U1115 (N_1115,In_1390,In_277);
or U1116 (N_1116,In_1365,In_274);
nor U1117 (N_1117,In_1043,In_237);
nor U1118 (N_1118,In_1120,In_895);
xor U1119 (N_1119,In_1497,In_625);
nor U1120 (N_1120,In_169,In_1417);
and U1121 (N_1121,In_571,In_1289);
and U1122 (N_1122,In_943,In_1348);
nand U1123 (N_1123,In_1155,In_1079);
or U1124 (N_1124,In_960,In_1311);
and U1125 (N_1125,In_995,In_960);
or U1126 (N_1126,In_694,In_367);
and U1127 (N_1127,In_126,In_727);
nand U1128 (N_1128,In_477,In_1160);
xor U1129 (N_1129,In_776,In_12);
and U1130 (N_1130,In_1349,In_3);
or U1131 (N_1131,In_1083,In_689);
or U1132 (N_1132,In_302,In_212);
nor U1133 (N_1133,In_190,In_592);
and U1134 (N_1134,In_171,In_1352);
and U1135 (N_1135,In_558,In_501);
nand U1136 (N_1136,In_73,In_224);
xnor U1137 (N_1137,In_951,In_38);
nor U1138 (N_1138,In_476,In_168);
xor U1139 (N_1139,In_67,In_17);
xnor U1140 (N_1140,In_1003,In_687);
nand U1141 (N_1141,In_750,In_831);
nand U1142 (N_1142,In_1477,In_1299);
nand U1143 (N_1143,In_1104,In_1360);
nor U1144 (N_1144,In_509,In_630);
or U1145 (N_1145,In_1204,In_1251);
nand U1146 (N_1146,In_1023,In_1060);
and U1147 (N_1147,In_724,In_303);
nand U1148 (N_1148,In_70,In_156);
nor U1149 (N_1149,In_423,In_1067);
or U1150 (N_1150,In_78,In_1189);
nand U1151 (N_1151,In_947,In_387);
or U1152 (N_1152,In_83,In_1051);
nand U1153 (N_1153,In_123,In_412);
or U1154 (N_1154,In_726,In_1468);
nand U1155 (N_1155,In_784,In_240);
nor U1156 (N_1156,In_1006,In_620);
and U1157 (N_1157,In_990,In_1394);
or U1158 (N_1158,In_22,In_501);
or U1159 (N_1159,In_221,In_1466);
nor U1160 (N_1160,In_748,In_1395);
or U1161 (N_1161,In_1491,In_1200);
or U1162 (N_1162,In_1279,In_59);
nand U1163 (N_1163,In_1029,In_526);
or U1164 (N_1164,In_627,In_518);
nor U1165 (N_1165,In_1321,In_617);
nor U1166 (N_1166,In_408,In_456);
nand U1167 (N_1167,In_285,In_781);
nor U1168 (N_1168,In_1265,In_1207);
and U1169 (N_1169,In_695,In_1060);
nand U1170 (N_1170,In_998,In_172);
and U1171 (N_1171,In_918,In_1289);
or U1172 (N_1172,In_247,In_1170);
or U1173 (N_1173,In_989,In_29);
xor U1174 (N_1174,In_932,In_373);
xnor U1175 (N_1175,In_211,In_425);
nor U1176 (N_1176,In_1266,In_1483);
and U1177 (N_1177,In_320,In_893);
nand U1178 (N_1178,In_895,In_404);
nor U1179 (N_1179,In_644,In_856);
nor U1180 (N_1180,In_1288,In_1189);
or U1181 (N_1181,In_849,In_1128);
nor U1182 (N_1182,In_819,In_943);
nand U1183 (N_1183,In_464,In_1299);
or U1184 (N_1184,In_1111,In_1359);
xnor U1185 (N_1185,In_1490,In_552);
or U1186 (N_1186,In_1212,In_926);
or U1187 (N_1187,In_1283,In_966);
nand U1188 (N_1188,In_1427,In_1325);
and U1189 (N_1189,In_1143,In_521);
nand U1190 (N_1190,In_859,In_1075);
or U1191 (N_1191,In_1150,In_1350);
or U1192 (N_1192,In_1305,In_582);
nand U1193 (N_1193,In_1263,In_1228);
nor U1194 (N_1194,In_431,In_1193);
nor U1195 (N_1195,In_202,In_549);
and U1196 (N_1196,In_567,In_1059);
nand U1197 (N_1197,In_578,In_1385);
xnor U1198 (N_1198,In_972,In_629);
or U1199 (N_1199,In_955,In_1479);
nor U1200 (N_1200,In_387,In_437);
nand U1201 (N_1201,In_890,In_900);
or U1202 (N_1202,In_1234,In_853);
nor U1203 (N_1203,In_1153,In_745);
nor U1204 (N_1204,In_1228,In_987);
or U1205 (N_1205,In_1225,In_692);
and U1206 (N_1206,In_313,In_1219);
and U1207 (N_1207,In_1403,In_498);
nand U1208 (N_1208,In_31,In_744);
or U1209 (N_1209,In_1181,In_467);
or U1210 (N_1210,In_1444,In_378);
nor U1211 (N_1211,In_1219,In_1192);
nor U1212 (N_1212,In_63,In_923);
or U1213 (N_1213,In_1198,In_462);
nor U1214 (N_1214,In_832,In_391);
nor U1215 (N_1215,In_1398,In_840);
nand U1216 (N_1216,In_551,In_55);
and U1217 (N_1217,In_296,In_1112);
or U1218 (N_1218,In_694,In_211);
and U1219 (N_1219,In_385,In_416);
nand U1220 (N_1220,In_255,In_1216);
and U1221 (N_1221,In_50,In_186);
nand U1222 (N_1222,In_598,In_1042);
and U1223 (N_1223,In_974,In_1152);
and U1224 (N_1224,In_1245,In_590);
nand U1225 (N_1225,In_275,In_298);
nor U1226 (N_1226,In_1136,In_1201);
nor U1227 (N_1227,In_801,In_418);
or U1228 (N_1228,In_575,In_1058);
or U1229 (N_1229,In_903,In_1292);
or U1230 (N_1230,In_118,In_31);
nand U1231 (N_1231,In_473,In_1186);
or U1232 (N_1232,In_1294,In_616);
or U1233 (N_1233,In_664,In_252);
nand U1234 (N_1234,In_891,In_1175);
nor U1235 (N_1235,In_976,In_718);
nand U1236 (N_1236,In_1438,In_1058);
nand U1237 (N_1237,In_83,In_327);
nor U1238 (N_1238,In_1365,In_326);
xnor U1239 (N_1239,In_195,In_871);
and U1240 (N_1240,In_405,In_1278);
or U1241 (N_1241,In_430,In_125);
nor U1242 (N_1242,In_389,In_1261);
nor U1243 (N_1243,In_1380,In_148);
or U1244 (N_1244,In_652,In_636);
nand U1245 (N_1245,In_435,In_626);
or U1246 (N_1246,In_577,In_636);
or U1247 (N_1247,In_208,In_1423);
nand U1248 (N_1248,In_250,In_1235);
nor U1249 (N_1249,In_51,In_1080);
nor U1250 (N_1250,In_1095,In_302);
and U1251 (N_1251,In_822,In_602);
nand U1252 (N_1252,In_1406,In_520);
nand U1253 (N_1253,In_163,In_1100);
nand U1254 (N_1254,In_183,In_1304);
nand U1255 (N_1255,In_679,In_1250);
xnor U1256 (N_1256,In_470,In_851);
xnor U1257 (N_1257,In_1195,In_1494);
nor U1258 (N_1258,In_569,In_887);
nor U1259 (N_1259,In_126,In_760);
xor U1260 (N_1260,In_1174,In_598);
or U1261 (N_1261,In_58,In_1286);
xnor U1262 (N_1262,In_1470,In_1023);
and U1263 (N_1263,In_136,In_626);
nand U1264 (N_1264,In_320,In_365);
or U1265 (N_1265,In_60,In_576);
nor U1266 (N_1266,In_807,In_882);
nand U1267 (N_1267,In_1308,In_1063);
nor U1268 (N_1268,In_615,In_646);
nand U1269 (N_1269,In_739,In_256);
nor U1270 (N_1270,In_511,In_349);
xnor U1271 (N_1271,In_1127,In_782);
or U1272 (N_1272,In_890,In_1478);
and U1273 (N_1273,In_290,In_345);
xnor U1274 (N_1274,In_1308,In_88);
nand U1275 (N_1275,In_415,In_1440);
nand U1276 (N_1276,In_1058,In_630);
and U1277 (N_1277,In_1280,In_211);
nor U1278 (N_1278,In_589,In_582);
nor U1279 (N_1279,In_1301,In_58);
or U1280 (N_1280,In_323,In_1276);
nor U1281 (N_1281,In_1371,In_511);
xnor U1282 (N_1282,In_919,In_111);
and U1283 (N_1283,In_562,In_1495);
xnor U1284 (N_1284,In_1063,In_675);
nor U1285 (N_1285,In_385,In_654);
xnor U1286 (N_1286,In_431,In_449);
nor U1287 (N_1287,In_762,In_1378);
nor U1288 (N_1288,In_227,In_819);
nor U1289 (N_1289,In_1033,In_1018);
nor U1290 (N_1290,In_1271,In_161);
nand U1291 (N_1291,In_1156,In_1124);
and U1292 (N_1292,In_502,In_932);
nand U1293 (N_1293,In_943,In_117);
nor U1294 (N_1294,In_268,In_919);
nand U1295 (N_1295,In_1241,In_1022);
nand U1296 (N_1296,In_58,In_1026);
nor U1297 (N_1297,In_1300,In_363);
and U1298 (N_1298,In_896,In_348);
or U1299 (N_1299,In_605,In_993);
or U1300 (N_1300,In_916,In_202);
nor U1301 (N_1301,In_857,In_315);
nand U1302 (N_1302,In_1176,In_994);
and U1303 (N_1303,In_151,In_1245);
and U1304 (N_1304,In_1028,In_507);
nor U1305 (N_1305,In_952,In_206);
nor U1306 (N_1306,In_508,In_52);
or U1307 (N_1307,In_163,In_545);
nor U1308 (N_1308,In_735,In_515);
and U1309 (N_1309,In_676,In_591);
xnor U1310 (N_1310,In_145,In_612);
or U1311 (N_1311,In_319,In_761);
nor U1312 (N_1312,In_1064,In_634);
nor U1313 (N_1313,In_343,In_389);
and U1314 (N_1314,In_74,In_46);
nand U1315 (N_1315,In_1388,In_221);
nand U1316 (N_1316,In_1494,In_1079);
nand U1317 (N_1317,In_1102,In_1397);
xor U1318 (N_1318,In_899,In_172);
and U1319 (N_1319,In_848,In_10);
xor U1320 (N_1320,In_1026,In_132);
nor U1321 (N_1321,In_1040,In_1176);
nor U1322 (N_1322,In_32,In_318);
and U1323 (N_1323,In_1440,In_1392);
xor U1324 (N_1324,In_792,In_481);
or U1325 (N_1325,In_265,In_1469);
nor U1326 (N_1326,In_37,In_633);
nor U1327 (N_1327,In_689,In_411);
nor U1328 (N_1328,In_176,In_403);
and U1329 (N_1329,In_260,In_335);
nor U1330 (N_1330,In_969,In_960);
or U1331 (N_1331,In_867,In_689);
or U1332 (N_1332,In_91,In_154);
nand U1333 (N_1333,In_515,In_1063);
nor U1334 (N_1334,In_1092,In_1006);
nor U1335 (N_1335,In_1462,In_992);
xnor U1336 (N_1336,In_997,In_1259);
xnor U1337 (N_1337,In_37,In_948);
xor U1338 (N_1338,In_99,In_1115);
xnor U1339 (N_1339,In_1407,In_428);
and U1340 (N_1340,In_1078,In_626);
nand U1341 (N_1341,In_1235,In_1373);
nor U1342 (N_1342,In_1344,In_46);
nand U1343 (N_1343,In_1462,In_591);
nor U1344 (N_1344,In_116,In_222);
or U1345 (N_1345,In_672,In_271);
nor U1346 (N_1346,In_291,In_249);
and U1347 (N_1347,In_1185,In_207);
nor U1348 (N_1348,In_982,In_689);
or U1349 (N_1349,In_85,In_1438);
nor U1350 (N_1350,In_1148,In_670);
nor U1351 (N_1351,In_57,In_1023);
nand U1352 (N_1352,In_177,In_721);
xnor U1353 (N_1353,In_951,In_977);
nand U1354 (N_1354,In_1193,In_248);
nor U1355 (N_1355,In_97,In_1165);
nand U1356 (N_1356,In_74,In_1172);
and U1357 (N_1357,In_264,In_472);
and U1358 (N_1358,In_783,In_247);
and U1359 (N_1359,In_821,In_438);
or U1360 (N_1360,In_717,In_447);
nand U1361 (N_1361,In_235,In_658);
nor U1362 (N_1362,In_610,In_15);
and U1363 (N_1363,In_1272,In_637);
and U1364 (N_1364,In_267,In_1401);
nand U1365 (N_1365,In_249,In_702);
and U1366 (N_1366,In_1065,In_440);
or U1367 (N_1367,In_1071,In_1152);
nor U1368 (N_1368,In_1391,In_1267);
xor U1369 (N_1369,In_237,In_1004);
nand U1370 (N_1370,In_1302,In_273);
and U1371 (N_1371,In_444,In_1259);
nand U1372 (N_1372,In_1327,In_1402);
and U1373 (N_1373,In_1470,In_665);
nor U1374 (N_1374,In_114,In_907);
xnor U1375 (N_1375,In_914,In_25);
nor U1376 (N_1376,In_364,In_56);
nand U1377 (N_1377,In_1486,In_1343);
and U1378 (N_1378,In_895,In_736);
and U1379 (N_1379,In_950,In_361);
and U1380 (N_1380,In_959,In_981);
or U1381 (N_1381,In_846,In_703);
and U1382 (N_1382,In_268,In_1441);
and U1383 (N_1383,In_1430,In_51);
and U1384 (N_1384,In_757,In_382);
or U1385 (N_1385,In_769,In_747);
and U1386 (N_1386,In_935,In_565);
xnor U1387 (N_1387,In_346,In_700);
nor U1388 (N_1388,In_745,In_789);
nor U1389 (N_1389,In_98,In_629);
and U1390 (N_1390,In_1465,In_1044);
or U1391 (N_1391,In_325,In_1368);
or U1392 (N_1392,In_452,In_975);
or U1393 (N_1393,In_983,In_221);
or U1394 (N_1394,In_1237,In_1370);
and U1395 (N_1395,In_194,In_61);
nand U1396 (N_1396,In_1146,In_499);
xnor U1397 (N_1397,In_673,In_922);
nand U1398 (N_1398,In_94,In_1258);
nor U1399 (N_1399,In_729,In_643);
or U1400 (N_1400,In_718,In_999);
nor U1401 (N_1401,In_827,In_768);
or U1402 (N_1402,In_961,In_1109);
nor U1403 (N_1403,In_38,In_448);
nand U1404 (N_1404,In_1266,In_1181);
and U1405 (N_1405,In_1017,In_1167);
nand U1406 (N_1406,In_1045,In_183);
and U1407 (N_1407,In_1210,In_904);
or U1408 (N_1408,In_1105,In_556);
nor U1409 (N_1409,In_1038,In_1139);
and U1410 (N_1410,In_184,In_1320);
nand U1411 (N_1411,In_307,In_80);
nor U1412 (N_1412,In_865,In_617);
xnor U1413 (N_1413,In_495,In_509);
nand U1414 (N_1414,In_14,In_612);
or U1415 (N_1415,In_1417,In_1307);
nor U1416 (N_1416,In_1210,In_1269);
or U1417 (N_1417,In_312,In_1268);
nor U1418 (N_1418,In_1074,In_954);
and U1419 (N_1419,In_479,In_82);
and U1420 (N_1420,In_1283,In_866);
nand U1421 (N_1421,In_1370,In_1416);
or U1422 (N_1422,In_1144,In_862);
xnor U1423 (N_1423,In_1298,In_772);
nor U1424 (N_1424,In_467,In_144);
and U1425 (N_1425,In_133,In_181);
or U1426 (N_1426,In_379,In_162);
nor U1427 (N_1427,In_41,In_788);
and U1428 (N_1428,In_703,In_875);
and U1429 (N_1429,In_432,In_962);
nor U1430 (N_1430,In_899,In_538);
nand U1431 (N_1431,In_290,In_1462);
xor U1432 (N_1432,In_241,In_572);
and U1433 (N_1433,In_1049,In_141);
nand U1434 (N_1434,In_695,In_1129);
nand U1435 (N_1435,In_1167,In_287);
nand U1436 (N_1436,In_1103,In_189);
or U1437 (N_1437,In_1456,In_305);
nor U1438 (N_1438,In_250,In_587);
nor U1439 (N_1439,In_480,In_219);
nor U1440 (N_1440,In_429,In_1424);
or U1441 (N_1441,In_1035,In_128);
nor U1442 (N_1442,In_764,In_303);
or U1443 (N_1443,In_836,In_862);
nor U1444 (N_1444,In_1289,In_667);
or U1445 (N_1445,In_324,In_784);
nor U1446 (N_1446,In_1312,In_54);
xor U1447 (N_1447,In_1346,In_641);
nor U1448 (N_1448,In_162,In_1214);
and U1449 (N_1449,In_1483,In_257);
nand U1450 (N_1450,In_358,In_1242);
or U1451 (N_1451,In_1084,In_22);
or U1452 (N_1452,In_1358,In_597);
and U1453 (N_1453,In_1329,In_1281);
or U1454 (N_1454,In_413,In_1063);
nand U1455 (N_1455,In_260,In_1221);
nand U1456 (N_1456,In_149,In_1088);
or U1457 (N_1457,In_1339,In_639);
nand U1458 (N_1458,In_80,In_993);
xnor U1459 (N_1459,In_857,In_35);
or U1460 (N_1460,In_1260,In_967);
xor U1461 (N_1461,In_366,In_1031);
and U1462 (N_1462,In_265,In_110);
or U1463 (N_1463,In_416,In_1055);
nor U1464 (N_1464,In_1034,In_464);
or U1465 (N_1465,In_423,In_298);
nand U1466 (N_1466,In_305,In_802);
nand U1467 (N_1467,In_819,In_208);
nor U1468 (N_1468,In_863,In_239);
and U1469 (N_1469,In_875,In_1195);
or U1470 (N_1470,In_576,In_1051);
nor U1471 (N_1471,In_686,In_1462);
and U1472 (N_1472,In_1280,In_1416);
nand U1473 (N_1473,In_320,In_800);
nor U1474 (N_1474,In_1417,In_583);
nor U1475 (N_1475,In_905,In_357);
nand U1476 (N_1476,In_650,In_1317);
nand U1477 (N_1477,In_294,In_934);
nand U1478 (N_1478,In_449,In_1124);
or U1479 (N_1479,In_1471,In_720);
or U1480 (N_1480,In_1200,In_502);
or U1481 (N_1481,In_327,In_1020);
and U1482 (N_1482,In_792,In_638);
or U1483 (N_1483,In_277,In_345);
nor U1484 (N_1484,In_1372,In_1248);
nor U1485 (N_1485,In_967,In_1041);
nand U1486 (N_1486,In_1450,In_618);
and U1487 (N_1487,In_1462,In_1146);
nand U1488 (N_1488,In_890,In_1042);
and U1489 (N_1489,In_1260,In_629);
or U1490 (N_1490,In_747,In_415);
nor U1491 (N_1491,In_1224,In_917);
xor U1492 (N_1492,In_1280,In_1043);
or U1493 (N_1493,In_299,In_619);
nor U1494 (N_1494,In_405,In_1233);
and U1495 (N_1495,In_1412,In_38);
and U1496 (N_1496,In_1436,In_339);
and U1497 (N_1497,In_1166,In_382);
and U1498 (N_1498,In_138,In_228);
or U1499 (N_1499,In_1322,In_587);
or U1500 (N_1500,N_1273,N_91);
nand U1501 (N_1501,N_1350,N_64);
and U1502 (N_1502,N_1044,N_541);
and U1503 (N_1503,N_770,N_160);
and U1504 (N_1504,N_885,N_533);
and U1505 (N_1505,N_1051,N_1149);
nor U1506 (N_1506,N_406,N_1302);
nor U1507 (N_1507,N_810,N_520);
nand U1508 (N_1508,N_1128,N_558);
nand U1509 (N_1509,N_838,N_466);
nand U1510 (N_1510,N_60,N_288);
nor U1511 (N_1511,N_1385,N_419);
nand U1512 (N_1512,N_1216,N_1112);
nor U1513 (N_1513,N_526,N_76);
and U1514 (N_1514,N_129,N_229);
and U1515 (N_1515,N_472,N_185);
or U1516 (N_1516,N_826,N_556);
nand U1517 (N_1517,N_470,N_1248);
xnor U1518 (N_1518,N_336,N_342);
or U1519 (N_1519,N_878,N_223);
and U1520 (N_1520,N_719,N_1133);
xor U1521 (N_1521,N_1214,N_80);
nand U1522 (N_1522,N_124,N_1146);
nand U1523 (N_1523,N_150,N_1315);
nand U1524 (N_1524,N_148,N_18);
nor U1525 (N_1525,N_230,N_371);
or U1526 (N_1526,N_1353,N_509);
and U1527 (N_1527,N_999,N_169);
nor U1528 (N_1528,N_1262,N_337);
and U1529 (N_1529,N_659,N_487);
nor U1530 (N_1530,N_334,N_1161);
or U1531 (N_1531,N_784,N_711);
nor U1532 (N_1532,N_1108,N_820);
or U1533 (N_1533,N_521,N_1032);
and U1534 (N_1534,N_311,N_614);
or U1535 (N_1535,N_671,N_1278);
nor U1536 (N_1536,N_1176,N_1284);
xor U1537 (N_1537,N_324,N_1489);
nand U1538 (N_1538,N_530,N_641);
nand U1539 (N_1539,N_465,N_836);
nor U1540 (N_1540,N_847,N_1289);
nor U1541 (N_1541,N_1387,N_738);
nand U1542 (N_1542,N_1317,N_1480);
nor U1543 (N_1543,N_226,N_1107);
or U1544 (N_1544,N_849,N_574);
and U1545 (N_1545,N_1467,N_207);
nor U1546 (N_1546,N_271,N_1265);
nand U1547 (N_1547,N_1338,N_709);
nor U1548 (N_1548,N_1346,N_568);
xnor U1549 (N_1549,N_3,N_412);
nor U1550 (N_1550,N_1141,N_218);
and U1551 (N_1551,N_636,N_1300);
or U1552 (N_1552,N_1193,N_834);
xnor U1553 (N_1553,N_189,N_537);
nand U1554 (N_1554,N_1170,N_612);
and U1555 (N_1555,N_1293,N_1089);
and U1556 (N_1556,N_1426,N_536);
nor U1557 (N_1557,N_1410,N_1144);
nor U1558 (N_1558,N_903,N_1490);
nor U1559 (N_1559,N_260,N_173);
nor U1560 (N_1560,N_984,N_134);
nor U1561 (N_1561,N_908,N_759);
xor U1562 (N_1562,N_831,N_590);
and U1563 (N_1563,N_1336,N_1160);
nor U1564 (N_1564,N_430,N_339);
and U1565 (N_1565,N_1428,N_1279);
nand U1566 (N_1566,N_85,N_151);
or U1567 (N_1567,N_504,N_289);
xor U1568 (N_1568,N_186,N_962);
xnor U1569 (N_1569,N_159,N_750);
or U1570 (N_1570,N_544,N_1227);
xor U1571 (N_1571,N_23,N_691);
and U1572 (N_1572,N_437,N_771);
and U1573 (N_1573,N_615,N_548);
nand U1574 (N_1574,N_296,N_110);
and U1575 (N_1575,N_843,N_588);
nor U1576 (N_1576,N_1377,N_1168);
nor U1577 (N_1577,N_2,N_1482);
xor U1578 (N_1578,N_88,N_1013);
nor U1579 (N_1579,N_1126,N_47);
xor U1580 (N_1580,N_469,N_1362);
xor U1581 (N_1581,N_1328,N_667);
nand U1582 (N_1582,N_1201,N_506);
nor U1583 (N_1583,N_1424,N_354);
nand U1584 (N_1584,N_1186,N_1460);
and U1585 (N_1585,N_193,N_922);
and U1586 (N_1586,N_212,N_247);
nor U1587 (N_1587,N_1406,N_261);
xor U1588 (N_1588,N_255,N_792);
nor U1589 (N_1589,N_462,N_499);
nor U1590 (N_1590,N_741,N_475);
or U1591 (N_1591,N_1115,N_1469);
and U1592 (N_1592,N_917,N_603);
or U1593 (N_1593,N_886,N_190);
xor U1594 (N_1594,N_1208,N_914);
or U1595 (N_1595,N_344,N_1202);
nand U1596 (N_1596,N_935,N_726);
and U1597 (N_1597,N_263,N_1091);
nor U1598 (N_1598,N_1435,N_206);
nand U1599 (N_1599,N_1322,N_915);
nand U1600 (N_1600,N_477,N_73);
or U1601 (N_1601,N_292,N_880);
and U1602 (N_1602,N_1466,N_1197);
nor U1603 (N_1603,N_822,N_388);
nor U1604 (N_1604,N_158,N_303);
or U1605 (N_1605,N_454,N_168);
or U1606 (N_1606,N_593,N_366);
nand U1607 (N_1607,N_86,N_276);
nor U1608 (N_1608,N_1207,N_128);
or U1609 (N_1609,N_748,N_974);
nand U1610 (N_1610,N_500,N_1403);
xnor U1611 (N_1611,N_1233,N_1283);
or U1612 (N_1612,N_1188,N_635);
xor U1613 (N_1613,N_712,N_1026);
xor U1614 (N_1614,N_1349,N_936);
nand U1615 (N_1615,N_425,N_595);
and U1616 (N_1616,N_54,N_702);
and U1617 (N_1617,N_932,N_877);
nor U1618 (N_1618,N_449,N_1347);
nor U1619 (N_1619,N_845,N_1156);
nor U1620 (N_1620,N_460,N_217);
nor U1621 (N_1621,N_1306,N_902);
nor U1622 (N_1622,N_390,N_731);
nor U1623 (N_1623,N_569,N_524);
and U1624 (N_1624,N_1251,N_357);
nand U1625 (N_1625,N_258,N_1035);
and U1626 (N_1626,N_241,N_1166);
or U1627 (N_1627,N_468,N_823);
nand U1628 (N_1628,N_14,N_51);
nand U1629 (N_1629,N_347,N_685);
or U1630 (N_1630,N_201,N_282);
nand U1631 (N_1631,N_1028,N_543);
nand U1632 (N_1632,N_1185,N_1454);
nand U1633 (N_1633,N_1183,N_340);
nand U1634 (N_1634,N_815,N_1020);
and U1635 (N_1635,N_889,N_1354);
or U1636 (N_1636,N_1103,N_627);
or U1637 (N_1637,N_651,N_862);
or U1638 (N_1638,N_179,N_1021);
and U1639 (N_1639,N_853,N_16);
or U1640 (N_1640,N_1043,N_798);
nand U1641 (N_1641,N_243,N_571);
nor U1642 (N_1642,N_278,N_1179);
nand U1643 (N_1643,N_1461,N_944);
and U1644 (N_1644,N_1215,N_431);
nor U1645 (N_1645,N_1340,N_961);
nor U1646 (N_1646,N_1364,N_538);
and U1647 (N_1647,N_5,N_140);
nand U1648 (N_1648,N_1030,N_417);
nor U1649 (N_1649,N_507,N_1450);
nor U1650 (N_1650,N_1255,N_341);
nor U1651 (N_1651,N_989,N_1079);
or U1652 (N_1652,N_988,N_1039);
nor U1653 (N_1653,N_529,N_52);
or U1654 (N_1654,N_916,N_154);
or U1655 (N_1655,N_29,N_827);
and U1656 (N_1656,N_1453,N_65);
nand U1657 (N_1657,N_428,N_482);
nand U1658 (N_1658,N_1199,N_355);
or U1659 (N_1659,N_319,N_503);
nor U1660 (N_1660,N_1427,N_152);
nand U1661 (N_1661,N_1298,N_1105);
nor U1662 (N_1662,N_1037,N_6);
nand U1663 (N_1663,N_1145,N_391);
nor U1664 (N_1664,N_1131,N_952);
and U1665 (N_1665,N_597,N_800);
or U1666 (N_1666,N_1059,N_325);
nor U1667 (N_1667,N_1368,N_739);
and U1668 (N_1668,N_767,N_581);
or U1669 (N_1669,N_1154,N_403);
or U1670 (N_1670,N_839,N_683);
and U1671 (N_1671,N_634,N_705);
nand U1672 (N_1672,N_1433,N_970);
nor U1673 (N_1673,N_921,N_385);
and U1674 (N_1674,N_1425,N_8);
or U1675 (N_1675,N_138,N_755);
and U1676 (N_1676,N_119,N_649);
and U1677 (N_1677,N_644,N_560);
or U1678 (N_1678,N_1080,N_1174);
or U1679 (N_1679,N_424,N_931);
nand U1680 (N_1680,N_133,N_1242);
and U1681 (N_1681,N_760,N_1012);
or U1682 (N_1682,N_182,N_1111);
nor U1683 (N_1683,N_98,N_455);
and U1684 (N_1684,N_298,N_1083);
nand U1685 (N_1685,N_225,N_807);
or U1686 (N_1686,N_1061,N_1240);
and U1687 (N_1687,N_638,N_584);
nand U1688 (N_1688,N_7,N_1003);
and U1689 (N_1689,N_415,N_1439);
nor U1690 (N_1690,N_1132,N_632);
nand U1691 (N_1691,N_1245,N_155);
xnor U1692 (N_1692,N_1150,N_1184);
xor U1693 (N_1693,N_491,N_768);
nand U1694 (N_1694,N_576,N_686);
nand U1695 (N_1695,N_959,N_1191);
xor U1696 (N_1696,N_732,N_1415);
nor U1697 (N_1697,N_549,N_411);
or U1698 (N_1698,N_1041,N_1475);
nand U1699 (N_1699,N_1281,N_1253);
xor U1700 (N_1700,N_97,N_1110);
xnor U1701 (N_1701,N_617,N_62);
and U1702 (N_1702,N_82,N_979);
nand U1703 (N_1703,N_214,N_1238);
nand U1704 (N_1704,N_299,N_71);
nand U1705 (N_1705,N_601,N_332);
or U1706 (N_1706,N_219,N_343);
nor U1707 (N_1707,N_435,N_1206);
or U1708 (N_1708,N_1429,N_1065);
nand U1709 (N_1709,N_523,N_1046);
nand U1710 (N_1710,N_1437,N_1153);
xnor U1711 (N_1711,N_443,N_28);
and U1712 (N_1712,N_493,N_892);
or U1713 (N_1713,N_1499,N_697);
or U1714 (N_1714,N_1396,N_251);
nor U1715 (N_1715,N_400,N_335);
nor U1716 (N_1716,N_934,N_1481);
nor U1717 (N_1717,N_473,N_266);
nand U1718 (N_1718,N_871,N_1177);
and U1719 (N_1719,N_898,N_284);
nand U1720 (N_1720,N_1224,N_640);
nor U1721 (N_1721,N_866,N_814);
and U1722 (N_1722,N_444,N_1304);
or U1723 (N_1723,N_84,N_525);
nor U1724 (N_1724,N_135,N_825);
nand U1725 (N_1725,N_1102,N_832);
and U1726 (N_1726,N_893,N_897);
xor U1727 (N_1727,N_1363,N_972);
nand U1728 (N_1728,N_202,N_293);
nor U1729 (N_1729,N_680,N_253);
nor U1730 (N_1730,N_211,N_375);
or U1731 (N_1731,N_381,N_1143);
xor U1732 (N_1732,N_365,N_658);
nand U1733 (N_1733,N_1130,N_1001);
nand U1734 (N_1734,N_1351,N_410);
xor U1735 (N_1735,N_174,N_1383);
and U1736 (N_1736,N_378,N_1282);
and U1737 (N_1737,N_130,N_793);
and U1738 (N_1738,N_1477,N_1222);
or U1739 (N_1739,N_256,N_68);
nand U1740 (N_1740,N_653,N_254);
or U1741 (N_1741,N_801,N_1334);
and U1742 (N_1742,N_1098,N_824);
nand U1743 (N_1743,N_306,N_108);
or U1744 (N_1744,N_512,N_180);
and U1745 (N_1745,N_1123,N_362);
xnor U1746 (N_1746,N_539,N_89);
nand U1747 (N_1747,N_348,N_1458);
nor U1748 (N_1748,N_166,N_598);
nand U1749 (N_1749,N_439,N_1264);
or U1750 (N_1750,N_1250,N_372);
or U1751 (N_1751,N_684,N_716);
and U1752 (N_1752,N_352,N_811);
or U1753 (N_1753,N_162,N_111);
or U1754 (N_1754,N_1449,N_1371);
and U1755 (N_1755,N_237,N_1373);
nand U1756 (N_1756,N_95,N_1189);
nor U1757 (N_1757,N_657,N_1388);
nor U1758 (N_1758,N_83,N_1063);
or U1759 (N_1759,N_923,N_232);
and U1760 (N_1760,N_43,N_224);
nand U1761 (N_1761,N_890,N_446);
or U1762 (N_1762,N_115,N_244);
and U1763 (N_1763,N_604,N_474);
nand U1764 (N_1764,N_1088,N_136);
and U1765 (N_1765,N_331,N_1087);
nor U1766 (N_1766,N_1023,N_1301);
nor U1767 (N_1767,N_114,N_1448);
nor U1768 (N_1768,N_891,N_478);
or U1769 (N_1769,N_874,N_580);
and U1770 (N_1770,N_183,N_854);
or U1771 (N_1771,N_208,N_1212);
or U1772 (N_1772,N_220,N_476);
nand U1773 (N_1773,N_1078,N_955);
nand U1774 (N_1774,N_1047,N_630);
and U1775 (N_1775,N_1198,N_656);
and U1776 (N_1776,N_888,N_859);
xor U1777 (N_1777,N_730,N_295);
and U1778 (N_1778,N_949,N_1162);
and U1779 (N_1779,N_101,N_575);
or U1780 (N_1780,N_639,N_401);
or U1781 (N_1781,N_1033,N_1122);
and U1782 (N_1782,N_1099,N_1071);
or U1783 (N_1783,N_106,N_1280);
or U1784 (N_1784,N_673,N_534);
and U1785 (N_1785,N_1288,N_953);
and U1786 (N_1786,N_925,N_678);
and U1787 (N_1787,N_429,N_1465);
or U1788 (N_1788,N_389,N_620);
nand U1789 (N_1789,N_395,N_882);
or U1790 (N_1790,N_228,N_297);
nor U1791 (N_1791,N_420,N_699);
and U1792 (N_1792,N_690,N_0);
nor U1793 (N_1793,N_1005,N_484);
nand U1794 (N_1794,N_143,N_1101);
nor U1795 (N_1795,N_78,N_1268);
nor U1796 (N_1796,N_1297,N_1405);
and U1797 (N_1797,N_992,N_734);
and U1798 (N_1798,N_817,N_833);
or U1799 (N_1799,N_291,N_1374);
xnor U1800 (N_1800,N_1230,N_1400);
and U1801 (N_1801,N_1231,N_535);
and U1802 (N_1802,N_1002,N_1256);
and U1803 (N_1803,N_104,N_561);
and U1804 (N_1804,N_1492,N_49);
or U1805 (N_1805,N_585,N_518);
and U1806 (N_1806,N_579,N_1243);
or U1807 (N_1807,N_1380,N_830);
nor U1808 (N_1808,N_876,N_1022);
or U1809 (N_1809,N_756,N_38);
or U1810 (N_1810,N_307,N_710);
and U1811 (N_1811,N_589,N_144);
nand U1812 (N_1812,N_829,N_1048);
nand U1813 (N_1813,N_488,N_1129);
nor U1814 (N_1814,N_1075,N_252);
xnor U1815 (N_1815,N_1029,N_1137);
and U1816 (N_1816,N_776,N_294);
or U1817 (N_1817,N_812,N_433);
nor U1818 (N_1818,N_1342,N_851);
and U1819 (N_1819,N_1488,N_56);
or U1820 (N_1820,N_1470,N_281);
or U1821 (N_1821,N_930,N_199);
nand U1822 (N_1822,N_963,N_275);
nor U1823 (N_1823,N_1332,N_747);
or U1824 (N_1824,N_1444,N_39);
nand U1825 (N_1825,N_946,N_167);
xor U1826 (N_1826,N_528,N_459);
or U1827 (N_1827,N_187,N_125);
or U1828 (N_1828,N_1225,N_648);
xor U1829 (N_1829,N_577,N_996);
or U1830 (N_1830,N_321,N_1138);
or U1831 (N_1831,N_1018,N_1299);
nand U1832 (N_1832,N_868,N_971);
nand U1833 (N_1833,N_157,N_682);
and U1834 (N_1834,N_1459,N_464);
xnor U1835 (N_1835,N_704,N_1274);
and U1836 (N_1836,N_326,N_346);
nor U1837 (N_1837,N_1053,N_1010);
or U1838 (N_1838,N_987,N_1181);
nor U1839 (N_1839,N_951,N_1375);
nor U1840 (N_1840,N_272,N_485);
nor U1841 (N_1841,N_1422,N_610);
nor U1842 (N_1842,N_715,N_345);
or U1843 (N_1843,N_765,N_744);
nor U1844 (N_1844,N_15,N_50);
and U1845 (N_1845,N_1267,N_1117);
or U1846 (N_1846,N_761,N_1052);
xor U1847 (N_1847,N_1398,N_1476);
or U1848 (N_1848,N_677,N_943);
and U1849 (N_1849,N_178,N_668);
or U1850 (N_1850,N_1495,N_1257);
nand U1851 (N_1851,N_242,N_165);
or U1852 (N_1852,N_661,N_513);
nand U1853 (N_1853,N_669,N_41);
nor U1854 (N_1854,N_844,N_61);
nor U1855 (N_1855,N_63,N_234);
or U1856 (N_1856,N_1209,N_1235);
and U1857 (N_1857,N_495,N_727);
xor U1858 (N_1858,N_647,N_1443);
nand U1859 (N_1859,N_1163,N_545);
or U1860 (N_1860,N_377,N_586);
or U1861 (N_1861,N_990,N_522);
nand U1862 (N_1862,N_457,N_1182);
nand U1863 (N_1863,N_196,N_205);
nor U1864 (N_1864,N_985,N_591);
or U1865 (N_1865,N_494,N_370);
or U1866 (N_1866,N_783,N_414);
nor U1867 (N_1867,N_821,N_1218);
or U1868 (N_1868,N_613,N_1407);
and U1869 (N_1869,N_1271,N_1345);
nor U1870 (N_1870,N_947,N_1462);
xor U1871 (N_1871,N_940,N_426);
and U1872 (N_1872,N_386,N_1485);
nor U1873 (N_1873,N_1095,N_248);
and U1874 (N_1874,N_442,N_808);
xnor U1875 (N_1875,N_422,N_1077);
nor U1876 (N_1876,N_1445,N_1178);
or U1877 (N_1877,N_650,N_1436);
or U1878 (N_1878,N_856,N_164);
or U1879 (N_1879,N_479,N_156);
xnor U1880 (N_1880,N_1472,N_757);
or U1881 (N_1881,N_210,N_1430);
xnor U1882 (N_1882,N_175,N_1344);
nand U1883 (N_1883,N_1159,N_13);
or U1884 (N_1884,N_1127,N_440);
xnor U1885 (N_1885,N_1402,N_34);
xor U1886 (N_1886,N_1064,N_666);
or U1887 (N_1887,N_725,N_21);
nor U1888 (N_1888,N_624,N_583);
nand U1889 (N_1889,N_1084,N_94);
or U1890 (N_1890,N_1254,N_75);
or U1891 (N_1891,N_384,N_622);
nand U1892 (N_1892,N_1074,N_374);
or U1893 (N_1893,N_587,N_942);
nand U1894 (N_1894,N_1210,N_763);
nand U1895 (N_1895,N_799,N_599);
or U1896 (N_1896,N_787,N_803);
nand U1897 (N_1897,N_200,N_447);
nand U1898 (N_1898,N_563,N_1446);
and U1899 (N_1899,N_816,N_177);
nor U1900 (N_1900,N_10,N_122);
or U1901 (N_1901,N_899,N_141);
nand U1902 (N_1902,N_333,N_872);
and U1903 (N_1903,N_69,N_968);
nand U1904 (N_1904,N_142,N_879);
and U1905 (N_1905,N_769,N_1312);
nand U1906 (N_1906,N_161,N_112);
nand U1907 (N_1907,N_692,N_36);
nor U1908 (N_1908,N_637,N_1258);
nor U1909 (N_1909,N_689,N_1479);
nor U1910 (N_1910,N_250,N_928);
nand U1911 (N_1911,N_277,N_616);
or U1912 (N_1912,N_302,N_1038);
nor U1913 (N_1913,N_969,N_107);
and U1914 (N_1914,N_4,N_204);
or U1915 (N_1915,N_609,N_305);
nand U1916 (N_1916,N_626,N_222);
nand U1917 (N_1917,N_722,N_1329);
nand U1918 (N_1918,N_721,N_551);
nor U1919 (N_1919,N_100,N_858);
nand U1920 (N_1920,N_1416,N_53);
nor U1921 (N_1921,N_1165,N_919);
or U1922 (N_1922,N_611,N_758);
nand U1923 (N_1923,N_310,N_1211);
or U1924 (N_1924,N_498,N_910);
or U1925 (N_1925,N_766,N_1014);
and U1926 (N_1926,N_249,N_1220);
and U1927 (N_1927,N_1484,N_1316);
and U1928 (N_1928,N_1341,N_960);
or U1929 (N_1929,N_121,N_1171);
or U1930 (N_1930,N_1270,N_330);
nor U1931 (N_1931,N_1019,N_1070);
nand U1932 (N_1932,N_1434,N_35);
nor U1933 (N_1933,N_751,N_1379);
or U1934 (N_1934,N_1204,N_806);
and U1935 (N_1935,N_1008,N_1097);
or U1936 (N_1936,N_1408,N_458);
or U1937 (N_1937,N_707,N_486);
or U1938 (N_1938,N_245,N_688);
nor U1939 (N_1939,N_1333,N_1308);
or U1940 (N_1940,N_1195,N_117);
and U1941 (N_1941,N_1432,N_1239);
nor U1942 (N_1942,N_909,N_1440);
and U1943 (N_1943,N_1395,N_215);
nand U1944 (N_1944,N_287,N_663);
xnor U1945 (N_1945,N_777,N_309);
and U1946 (N_1946,N_965,N_1323);
nor U1947 (N_1947,N_1082,N_1468);
xor U1948 (N_1948,N_1229,N_981);
and U1949 (N_1949,N_954,N_1359);
or U1950 (N_1950,N_861,N_323);
nand U1951 (N_1951,N_1121,N_1324);
nor U1952 (N_1952,N_840,N_789);
and U1953 (N_1953,N_557,N_1348);
nand U1954 (N_1954,N_570,N_918);
nor U1955 (N_1955,N_818,N_280);
nor U1956 (N_1956,N_1247,N_1100);
and U1957 (N_1957,N_745,N_841);
xor U1958 (N_1958,N_933,N_813);
and U1959 (N_1959,N_701,N_116);
or U1960 (N_1960,N_132,N_1139);
nand U1961 (N_1961,N_857,N_1384);
and U1962 (N_1962,N_301,N_467);
xor U1963 (N_1963,N_1417,N_184);
xor U1964 (N_1964,N_300,N_360);
and U1965 (N_1965,N_1196,N_329);
xor U1966 (N_1966,N_67,N_1173);
nor U1967 (N_1967,N_1054,N_1420);
and U1968 (N_1968,N_399,N_1483);
nor U1969 (N_1969,N_1118,N_788);
or U1970 (N_1970,N_1090,N_267);
or U1971 (N_1971,N_700,N_1275);
xnor U1972 (N_1972,N_227,N_1114);
nand U1973 (N_1973,N_1120,N_42);
or U1974 (N_1974,N_1277,N_92);
nor U1975 (N_1975,N_779,N_957);
nor U1976 (N_1976,N_188,N_559);
nor U1977 (N_1977,N_269,N_749);
xnor U1978 (N_1978,N_976,N_735);
xnor U1979 (N_1979,N_1081,N_964);
xnor U1980 (N_1980,N_1116,N_894);
or U1981 (N_1981,N_920,N_1069);
and U1982 (N_1982,N_754,N_672);
and U1983 (N_1983,N_90,N_527);
or U1984 (N_1984,N_1187,N_316);
nand U1985 (N_1985,N_181,N_718);
nand U1986 (N_1986,N_1269,N_314);
xnor U1987 (N_1987,N_1004,N_884);
and U1988 (N_1988,N_1296,N_471);
or U1989 (N_1989,N_131,N_48);
and U1990 (N_1990,N_674,N_646);
or U1991 (N_1991,N_32,N_804);
nor U1992 (N_1992,N_983,N_693);
and U1993 (N_1993,N_772,N_553);
nand U1994 (N_1994,N_191,N_982);
nor U1995 (N_1995,N_363,N_1164);
or U1996 (N_1996,N_413,N_221);
and U1997 (N_1997,N_397,N_264);
nand U1998 (N_1998,N_552,N_358);
nor U1999 (N_1999,N_448,N_1167);
or U2000 (N_2000,N_432,N_1134);
and U2001 (N_2001,N_887,N_1140);
or U2002 (N_2002,N_995,N_1326);
nor U2003 (N_2003,N_1473,N_1357);
or U2004 (N_2004,N_665,N_550);
and U2005 (N_2005,N_285,N_147);
nand U2006 (N_2006,N_436,N_369);
nand U2007 (N_2007,N_72,N_1232);
or U2008 (N_2008,N_736,N_213);
or U2009 (N_2009,N_681,N_1025);
and U2010 (N_2010,N_592,N_194);
and U2011 (N_2011,N_1085,N_742);
or U2012 (N_2012,N_1062,N_864);
or U2013 (N_2013,N_379,N_393);
or U2014 (N_2014,N_404,N_775);
nor U2015 (N_2015,N_322,N_350);
xor U2016 (N_2016,N_975,N_1337);
nand U2017 (N_2017,N_231,N_728);
nor U2018 (N_2018,N_881,N_664);
nand U2019 (N_2019,N_1221,N_1050);
nor U2020 (N_2020,N_860,N_145);
nand U2021 (N_2021,N_1431,N_1321);
or U2022 (N_2022,N_1367,N_567);
nand U2023 (N_2023,N_1027,N_1223);
nand U2024 (N_2024,N_913,N_40);
xnor U2025 (N_2025,N_113,N_30);
and U2026 (N_2026,N_1180,N_1493);
xor U2027 (N_2027,N_44,N_1011);
or U2028 (N_2028,N_290,N_1017);
and U2029 (N_2029,N_794,N_514);
or U2030 (N_2030,N_991,N_1007);
nor U2031 (N_2031,N_24,N_1318);
nand U2032 (N_2032,N_1276,N_515);
or U2033 (N_2033,N_1066,N_58);
nor U2034 (N_2034,N_773,N_1382);
or U2035 (N_2035,N_1310,N_203);
nand U2036 (N_2036,N_835,N_746);
nor U2037 (N_2037,N_1414,N_163);
or U2038 (N_2038,N_368,N_1213);
or U2039 (N_2039,N_501,N_1190);
nand U2040 (N_2040,N_602,N_1266);
nor U2041 (N_2041,N_396,N_1366);
nor U2042 (N_2042,N_1136,N_216);
nor U2043 (N_2043,N_1192,N_1057);
nor U2044 (N_2044,N_320,N_96);
or U2045 (N_2045,N_1260,N_1313);
or U2046 (N_2046,N_895,N_555);
and U2047 (N_2047,N_1263,N_351);
or U2048 (N_2048,N_1356,N_273);
nand U2049 (N_2049,N_850,N_676);
or U2050 (N_2050,N_941,N_392);
nand U2051 (N_2051,N_505,N_1155);
nor U2052 (N_2052,N_780,N_945);
nand U2053 (N_2053,N_79,N_1327);
xor U2054 (N_2054,N_566,N_318);
nand U2055 (N_2055,N_197,N_643);
nand U2056 (N_2056,N_238,N_642);
or U2057 (N_2057,N_408,N_463);
nand U2058 (N_2058,N_896,N_480);
and U2059 (N_2059,N_828,N_367);
and U2060 (N_2060,N_628,N_1236);
nand U2061 (N_2061,N_937,N_502);
or U2062 (N_2062,N_279,N_1452);
and U2063 (N_2063,N_20,N_172);
and U2064 (N_2064,N_1352,N_578);
nor U2065 (N_2065,N_233,N_621);
nand U2066 (N_2066,N_376,N_623);
nor U2067 (N_2067,N_662,N_1096);
nor U2068 (N_2068,N_1113,N_59);
or U2069 (N_2069,N_1157,N_373);
nor U2070 (N_2070,N_993,N_364);
nand U2071 (N_2071,N_547,N_127);
or U2072 (N_2072,N_905,N_313);
or U2073 (N_2073,N_1401,N_11);
xnor U2074 (N_2074,N_619,N_1320);
and U2075 (N_2075,N_327,N_511);
nand U2076 (N_2076,N_46,N_540);
nor U2077 (N_2077,N_1378,N_1093);
and U2078 (N_2078,N_137,N_265);
or U2079 (N_2079,N_394,N_268);
or U2080 (N_2080,N_451,N_582);
nor U2081 (N_2081,N_805,N_338);
nand U2082 (N_2082,N_209,N_1290);
nor U2083 (N_2083,N_1272,N_631);
and U2084 (N_2084,N_1169,N_9);
and U2085 (N_2085,N_382,N_240);
and U2086 (N_2086,N_1365,N_416);
nor U2087 (N_2087,N_70,N_863);
nor U2088 (N_2088,N_171,N_1413);
xnor U2089 (N_2089,N_1152,N_126);
xnor U2090 (N_2090,N_1024,N_283);
nor U2091 (N_2091,N_508,N_192);
or U2092 (N_2092,N_790,N_418);
nor U2093 (N_2093,N_450,N_809);
nor U2094 (N_2094,N_956,N_1358);
and U2095 (N_2095,N_270,N_869);
xnor U2096 (N_2096,N_1175,N_139);
and U2097 (N_2097,N_262,N_1104);
nand U2098 (N_2098,N_87,N_239);
and U2099 (N_2099,N_25,N_1056);
or U2100 (N_2100,N_865,N_1335);
nand U2101 (N_2101,N_774,N_785);
nand U2102 (N_2102,N_1447,N_762);
or U2103 (N_2103,N_675,N_904);
nor U2104 (N_2104,N_737,N_149);
nor U2105 (N_2105,N_55,N_875);
and U2106 (N_2106,N_153,N_516);
nor U2107 (N_2107,N_315,N_1307);
and U2108 (N_2108,N_312,N_235);
and U2109 (N_2109,N_1497,N_906);
and U2110 (N_2110,N_1135,N_1076);
or U2111 (N_2111,N_1194,N_170);
and U2112 (N_2112,N_57,N_1092);
nor U2113 (N_2113,N_198,N_625);
and U2114 (N_2114,N_1376,N_1147);
and U2115 (N_2115,N_546,N_1471);
and U2116 (N_2116,N_383,N_1151);
nand U2117 (N_2117,N_713,N_929);
nand U2118 (N_2118,N_967,N_328);
or U2119 (N_2119,N_977,N_1331);
and U2120 (N_2120,N_842,N_12);
nor U2121 (N_2121,N_380,N_572);
nor U2122 (N_2122,N_565,N_883);
and U2123 (N_2123,N_966,N_74);
and U2124 (N_2124,N_1200,N_1285);
or U2125 (N_2125,N_510,N_706);
and U2126 (N_2126,N_1438,N_438);
xnor U2127 (N_2127,N_1464,N_600);
and U2128 (N_2128,N_1261,N_1498);
nor U2129 (N_2129,N_1397,N_1303);
nand U2130 (N_2130,N_1486,N_998);
nor U2131 (N_2131,N_786,N_489);
or U2132 (N_2132,N_1086,N_1252);
or U2133 (N_2133,N_1042,N_1399);
and U2134 (N_2134,N_1072,N_1040);
and U2135 (N_2135,N_1217,N_1419);
or U2136 (N_2136,N_1241,N_1009);
nor U2137 (N_2137,N_633,N_1494);
nand U2138 (N_2138,N_77,N_724);
nor U2139 (N_2139,N_1291,N_398);
or U2140 (N_2140,N_948,N_1246);
and U2141 (N_2141,N_409,N_720);
or U2142 (N_2142,N_1369,N_1421);
and U2143 (N_2143,N_986,N_1314);
or U2144 (N_2144,N_308,N_1474);
and U2145 (N_2145,N_246,N_434);
or U2146 (N_2146,N_1244,N_1158);
xnor U2147 (N_2147,N_1124,N_973);
nand U2148 (N_2148,N_618,N_938);
and U2149 (N_2149,N_645,N_1309);
nor U2150 (N_2150,N_1343,N_926);
nand U2151 (N_2151,N_1058,N_1016);
xnor U2152 (N_2152,N_778,N_37);
xnor U2153 (N_2153,N_698,N_402);
or U2154 (N_2154,N_723,N_532);
nand U2155 (N_2155,N_1325,N_870);
nand U2156 (N_2156,N_1404,N_1172);
and U2157 (N_2157,N_461,N_407);
xor U2158 (N_2158,N_900,N_1456);
xnor U2159 (N_2159,N_708,N_1478);
nand U2160 (N_2160,N_912,N_257);
and U2161 (N_2161,N_1287,N_441);
nand U2162 (N_2162,N_1036,N_66);
nand U2163 (N_2163,N_105,N_517);
nand U2164 (N_2164,N_1237,N_1361);
nand U2165 (N_2165,N_606,N_490);
xnor U2166 (N_2166,N_349,N_361);
nor U2167 (N_2167,N_703,N_740);
nor U2168 (N_2168,N_1073,N_195);
or U2169 (N_2169,N_99,N_1049);
nand U2170 (N_2170,N_573,N_1409);
and U2171 (N_2171,N_1045,N_1451);
xnor U2172 (N_2172,N_1249,N_1034);
nand U2173 (N_2173,N_958,N_1106);
xor U2174 (N_2174,N_1394,N_274);
nand U2175 (N_2175,N_605,N_1496);
and U2176 (N_2176,N_445,N_554);
nor U2177 (N_2177,N_1330,N_1423);
nand U2178 (N_2178,N_629,N_873);
nand U2179 (N_2179,N_717,N_236);
and U2180 (N_2180,N_427,N_492);
nor U2181 (N_2181,N_687,N_837);
nand U2182 (N_2182,N_19,N_753);
nand U2183 (N_2183,N_1418,N_542);
nand U2184 (N_2184,N_846,N_950);
or U2185 (N_2185,N_1219,N_259);
xor U2186 (N_2186,N_103,N_1148);
or U2187 (N_2187,N_608,N_1);
nand U2188 (N_2188,N_733,N_1412);
nand U2189 (N_2189,N_1390,N_696);
nor U2190 (N_2190,N_901,N_1311);
nand U2191 (N_2191,N_1372,N_796);
and U2192 (N_2192,N_26,N_1226);
or U2193 (N_2193,N_109,N_531);
xnor U2194 (N_2194,N_353,N_519);
nand U2195 (N_2195,N_654,N_1000);
xnor U2196 (N_2196,N_286,N_120);
nor U2197 (N_2197,N_782,N_1463);
or U2198 (N_2198,N_1228,N_997);
and U2199 (N_2199,N_481,N_1339);
and U2200 (N_2200,N_848,N_729);
xnor U2201 (N_2201,N_781,N_1360);
nor U2202 (N_2202,N_1491,N_655);
and U2203 (N_2203,N_1142,N_45);
or U2204 (N_2204,N_22,N_27);
nor U2205 (N_2205,N_802,N_855);
nand U2206 (N_2206,N_978,N_1295);
and U2207 (N_2207,N_1031,N_1442);
and U2208 (N_2208,N_123,N_867);
nor U2209 (N_2209,N_31,N_795);
nor U2210 (N_2210,N_660,N_1391);
nor U2211 (N_2211,N_819,N_1015);
or U2212 (N_2212,N_1060,N_927);
nor U2213 (N_2213,N_907,N_93);
nand U2214 (N_2214,N_452,N_118);
nand U2215 (N_2215,N_1370,N_317);
or U2216 (N_2216,N_652,N_359);
nor U2217 (N_2217,N_453,N_1286);
or U2218 (N_2218,N_497,N_102);
and U2219 (N_2219,N_679,N_1203);
or U2220 (N_2220,N_81,N_496);
and U2221 (N_2221,N_911,N_176);
nor U2222 (N_2222,N_1487,N_1455);
or U2223 (N_2223,N_939,N_564);
or U2224 (N_2224,N_1386,N_1441);
nand U2225 (N_2225,N_1068,N_1109);
and U2226 (N_2226,N_17,N_1305);
and U2227 (N_2227,N_1234,N_1355);
nor U2228 (N_2228,N_852,N_1006);
and U2229 (N_2229,N_1094,N_33);
or U2230 (N_2230,N_483,N_1381);
nor U2231 (N_2231,N_1125,N_1259);
or U2232 (N_2232,N_607,N_1205);
and U2233 (N_2233,N_1389,N_980);
nand U2234 (N_2234,N_994,N_1294);
nand U2235 (N_2235,N_670,N_714);
and U2236 (N_2236,N_421,N_387);
nor U2237 (N_2237,N_1392,N_1457);
nand U2238 (N_2238,N_1119,N_694);
or U2239 (N_2239,N_356,N_146);
xor U2240 (N_2240,N_304,N_594);
or U2241 (N_2241,N_764,N_1319);
xor U2242 (N_2242,N_405,N_562);
or U2243 (N_2243,N_797,N_423);
nor U2244 (N_2244,N_752,N_1067);
nor U2245 (N_2245,N_1393,N_743);
and U2246 (N_2246,N_695,N_596);
and U2247 (N_2247,N_924,N_456);
xor U2248 (N_2248,N_791,N_1292);
nor U2249 (N_2249,N_1055,N_1411);
and U2250 (N_2250,N_1448,N_961);
nand U2251 (N_2251,N_751,N_1387);
or U2252 (N_2252,N_54,N_650);
or U2253 (N_2253,N_950,N_1106);
nor U2254 (N_2254,N_46,N_1256);
xor U2255 (N_2255,N_655,N_972);
and U2256 (N_2256,N_952,N_169);
nand U2257 (N_2257,N_95,N_418);
xor U2258 (N_2258,N_1243,N_813);
xnor U2259 (N_2259,N_254,N_1383);
and U2260 (N_2260,N_383,N_1328);
and U2261 (N_2261,N_1058,N_1417);
nand U2262 (N_2262,N_1329,N_407);
xnor U2263 (N_2263,N_6,N_446);
nand U2264 (N_2264,N_261,N_460);
and U2265 (N_2265,N_150,N_380);
nand U2266 (N_2266,N_1065,N_45);
and U2267 (N_2267,N_663,N_1363);
and U2268 (N_2268,N_501,N_1062);
xnor U2269 (N_2269,N_1399,N_1464);
and U2270 (N_2270,N_672,N_339);
or U2271 (N_2271,N_1301,N_914);
and U2272 (N_2272,N_467,N_963);
or U2273 (N_2273,N_1486,N_1496);
and U2274 (N_2274,N_81,N_1432);
xor U2275 (N_2275,N_577,N_508);
or U2276 (N_2276,N_1021,N_44);
nand U2277 (N_2277,N_480,N_556);
nand U2278 (N_2278,N_693,N_590);
and U2279 (N_2279,N_889,N_509);
or U2280 (N_2280,N_914,N_1076);
or U2281 (N_2281,N_483,N_735);
and U2282 (N_2282,N_260,N_345);
and U2283 (N_2283,N_1479,N_9);
or U2284 (N_2284,N_269,N_850);
and U2285 (N_2285,N_1223,N_4);
xor U2286 (N_2286,N_963,N_1009);
nand U2287 (N_2287,N_846,N_612);
nor U2288 (N_2288,N_1226,N_1094);
nor U2289 (N_2289,N_588,N_497);
nand U2290 (N_2290,N_1368,N_1046);
or U2291 (N_2291,N_194,N_920);
and U2292 (N_2292,N_388,N_869);
nor U2293 (N_2293,N_1076,N_1172);
and U2294 (N_2294,N_226,N_1301);
or U2295 (N_2295,N_107,N_729);
xnor U2296 (N_2296,N_857,N_1349);
and U2297 (N_2297,N_563,N_458);
nor U2298 (N_2298,N_1320,N_569);
nor U2299 (N_2299,N_911,N_748);
and U2300 (N_2300,N_1243,N_849);
nor U2301 (N_2301,N_35,N_1135);
or U2302 (N_2302,N_1433,N_248);
nor U2303 (N_2303,N_1436,N_1157);
or U2304 (N_2304,N_493,N_160);
nor U2305 (N_2305,N_326,N_208);
nand U2306 (N_2306,N_908,N_1034);
nor U2307 (N_2307,N_1048,N_213);
or U2308 (N_2308,N_1480,N_666);
nand U2309 (N_2309,N_1247,N_863);
nor U2310 (N_2310,N_83,N_79);
nand U2311 (N_2311,N_931,N_377);
and U2312 (N_2312,N_610,N_165);
or U2313 (N_2313,N_346,N_117);
nor U2314 (N_2314,N_636,N_872);
or U2315 (N_2315,N_1482,N_959);
and U2316 (N_2316,N_0,N_341);
and U2317 (N_2317,N_613,N_0);
nand U2318 (N_2318,N_1497,N_935);
nand U2319 (N_2319,N_29,N_879);
nor U2320 (N_2320,N_335,N_243);
nand U2321 (N_2321,N_1018,N_1219);
nor U2322 (N_2322,N_531,N_1094);
nor U2323 (N_2323,N_1488,N_1012);
nand U2324 (N_2324,N_182,N_604);
or U2325 (N_2325,N_158,N_1138);
nand U2326 (N_2326,N_1041,N_252);
nor U2327 (N_2327,N_313,N_247);
xnor U2328 (N_2328,N_1022,N_1206);
nor U2329 (N_2329,N_1376,N_1052);
xor U2330 (N_2330,N_1111,N_1334);
or U2331 (N_2331,N_857,N_1449);
or U2332 (N_2332,N_1037,N_837);
nor U2333 (N_2333,N_161,N_947);
nand U2334 (N_2334,N_921,N_1301);
or U2335 (N_2335,N_937,N_932);
or U2336 (N_2336,N_1361,N_1208);
nand U2337 (N_2337,N_1385,N_828);
nor U2338 (N_2338,N_528,N_1058);
and U2339 (N_2339,N_907,N_71);
and U2340 (N_2340,N_1083,N_778);
nand U2341 (N_2341,N_963,N_964);
and U2342 (N_2342,N_1397,N_526);
or U2343 (N_2343,N_731,N_148);
nor U2344 (N_2344,N_288,N_510);
nor U2345 (N_2345,N_152,N_247);
or U2346 (N_2346,N_1486,N_507);
nor U2347 (N_2347,N_1107,N_1075);
and U2348 (N_2348,N_1432,N_529);
nor U2349 (N_2349,N_270,N_1131);
nor U2350 (N_2350,N_1076,N_673);
nand U2351 (N_2351,N_430,N_14);
and U2352 (N_2352,N_223,N_47);
nor U2353 (N_2353,N_1158,N_984);
xor U2354 (N_2354,N_572,N_192);
nand U2355 (N_2355,N_675,N_204);
or U2356 (N_2356,N_378,N_435);
or U2357 (N_2357,N_583,N_1395);
nor U2358 (N_2358,N_40,N_99);
nand U2359 (N_2359,N_998,N_393);
nor U2360 (N_2360,N_764,N_1381);
and U2361 (N_2361,N_734,N_1249);
or U2362 (N_2362,N_341,N_2);
or U2363 (N_2363,N_619,N_267);
nand U2364 (N_2364,N_375,N_1174);
xor U2365 (N_2365,N_130,N_524);
and U2366 (N_2366,N_203,N_157);
and U2367 (N_2367,N_1481,N_995);
or U2368 (N_2368,N_1037,N_849);
nor U2369 (N_2369,N_15,N_1067);
nor U2370 (N_2370,N_40,N_1403);
nand U2371 (N_2371,N_1418,N_738);
or U2372 (N_2372,N_121,N_150);
nand U2373 (N_2373,N_1213,N_1464);
and U2374 (N_2374,N_88,N_43);
and U2375 (N_2375,N_576,N_144);
or U2376 (N_2376,N_1289,N_925);
nand U2377 (N_2377,N_1264,N_629);
nand U2378 (N_2378,N_831,N_51);
and U2379 (N_2379,N_940,N_331);
or U2380 (N_2380,N_262,N_689);
nand U2381 (N_2381,N_741,N_986);
or U2382 (N_2382,N_170,N_1421);
nand U2383 (N_2383,N_1427,N_1400);
nand U2384 (N_2384,N_3,N_768);
and U2385 (N_2385,N_763,N_180);
and U2386 (N_2386,N_462,N_144);
nor U2387 (N_2387,N_968,N_207);
xnor U2388 (N_2388,N_52,N_455);
nand U2389 (N_2389,N_1182,N_498);
nor U2390 (N_2390,N_1073,N_404);
nor U2391 (N_2391,N_237,N_1041);
nand U2392 (N_2392,N_259,N_332);
or U2393 (N_2393,N_775,N_1173);
nand U2394 (N_2394,N_1311,N_342);
nor U2395 (N_2395,N_19,N_748);
or U2396 (N_2396,N_795,N_691);
and U2397 (N_2397,N_154,N_1371);
xnor U2398 (N_2398,N_1236,N_204);
xor U2399 (N_2399,N_2,N_472);
nand U2400 (N_2400,N_1325,N_512);
or U2401 (N_2401,N_93,N_11);
nor U2402 (N_2402,N_5,N_1);
and U2403 (N_2403,N_1324,N_165);
nand U2404 (N_2404,N_1233,N_492);
nand U2405 (N_2405,N_834,N_903);
and U2406 (N_2406,N_46,N_1269);
xnor U2407 (N_2407,N_518,N_962);
nand U2408 (N_2408,N_377,N_1175);
nor U2409 (N_2409,N_572,N_628);
nor U2410 (N_2410,N_1330,N_1203);
xnor U2411 (N_2411,N_139,N_46);
xnor U2412 (N_2412,N_803,N_80);
nand U2413 (N_2413,N_769,N_1363);
nor U2414 (N_2414,N_117,N_1430);
nand U2415 (N_2415,N_763,N_1365);
or U2416 (N_2416,N_558,N_1018);
and U2417 (N_2417,N_491,N_539);
nor U2418 (N_2418,N_98,N_174);
nor U2419 (N_2419,N_345,N_1007);
nand U2420 (N_2420,N_630,N_504);
nand U2421 (N_2421,N_133,N_96);
and U2422 (N_2422,N_337,N_1497);
nor U2423 (N_2423,N_184,N_1303);
nor U2424 (N_2424,N_1074,N_1359);
and U2425 (N_2425,N_1067,N_1407);
nor U2426 (N_2426,N_417,N_1388);
or U2427 (N_2427,N_483,N_442);
nand U2428 (N_2428,N_164,N_387);
nand U2429 (N_2429,N_659,N_1473);
and U2430 (N_2430,N_1448,N_692);
nand U2431 (N_2431,N_304,N_559);
and U2432 (N_2432,N_441,N_1161);
nand U2433 (N_2433,N_1211,N_766);
and U2434 (N_2434,N_925,N_1290);
xor U2435 (N_2435,N_1176,N_1151);
and U2436 (N_2436,N_990,N_165);
and U2437 (N_2437,N_324,N_676);
xor U2438 (N_2438,N_566,N_401);
or U2439 (N_2439,N_211,N_607);
and U2440 (N_2440,N_599,N_1171);
or U2441 (N_2441,N_1300,N_1339);
or U2442 (N_2442,N_891,N_208);
nand U2443 (N_2443,N_696,N_59);
nor U2444 (N_2444,N_1441,N_651);
and U2445 (N_2445,N_850,N_897);
nand U2446 (N_2446,N_1432,N_412);
or U2447 (N_2447,N_1356,N_1289);
nor U2448 (N_2448,N_375,N_652);
xnor U2449 (N_2449,N_937,N_1038);
nand U2450 (N_2450,N_123,N_128);
nand U2451 (N_2451,N_1063,N_359);
nand U2452 (N_2452,N_262,N_87);
or U2453 (N_2453,N_207,N_789);
and U2454 (N_2454,N_293,N_680);
or U2455 (N_2455,N_860,N_598);
or U2456 (N_2456,N_639,N_1220);
nor U2457 (N_2457,N_375,N_278);
xnor U2458 (N_2458,N_0,N_908);
or U2459 (N_2459,N_478,N_264);
or U2460 (N_2460,N_1001,N_1046);
nor U2461 (N_2461,N_241,N_413);
and U2462 (N_2462,N_473,N_1062);
and U2463 (N_2463,N_860,N_576);
nor U2464 (N_2464,N_497,N_607);
nor U2465 (N_2465,N_1193,N_583);
or U2466 (N_2466,N_1011,N_40);
or U2467 (N_2467,N_548,N_985);
or U2468 (N_2468,N_149,N_181);
nor U2469 (N_2469,N_251,N_1033);
xor U2470 (N_2470,N_1057,N_1033);
or U2471 (N_2471,N_1002,N_1242);
nand U2472 (N_2472,N_217,N_1250);
or U2473 (N_2473,N_630,N_536);
or U2474 (N_2474,N_884,N_765);
nand U2475 (N_2475,N_166,N_66);
or U2476 (N_2476,N_1405,N_1018);
nand U2477 (N_2477,N_516,N_1394);
or U2478 (N_2478,N_735,N_791);
nor U2479 (N_2479,N_1257,N_547);
nand U2480 (N_2480,N_684,N_1490);
nor U2481 (N_2481,N_1368,N_974);
and U2482 (N_2482,N_686,N_536);
and U2483 (N_2483,N_84,N_802);
nand U2484 (N_2484,N_559,N_773);
or U2485 (N_2485,N_740,N_1225);
or U2486 (N_2486,N_770,N_983);
nand U2487 (N_2487,N_1359,N_184);
and U2488 (N_2488,N_908,N_191);
nor U2489 (N_2489,N_202,N_380);
nand U2490 (N_2490,N_629,N_91);
nand U2491 (N_2491,N_1097,N_719);
and U2492 (N_2492,N_1445,N_934);
or U2493 (N_2493,N_812,N_962);
nand U2494 (N_2494,N_1039,N_1090);
nor U2495 (N_2495,N_1471,N_636);
nor U2496 (N_2496,N_951,N_601);
and U2497 (N_2497,N_613,N_246);
or U2498 (N_2498,N_840,N_780);
and U2499 (N_2499,N_223,N_314);
or U2500 (N_2500,N_583,N_330);
and U2501 (N_2501,N_876,N_1164);
or U2502 (N_2502,N_839,N_209);
and U2503 (N_2503,N_1157,N_129);
and U2504 (N_2504,N_224,N_792);
and U2505 (N_2505,N_387,N_1235);
nor U2506 (N_2506,N_948,N_831);
xor U2507 (N_2507,N_543,N_1326);
nor U2508 (N_2508,N_230,N_398);
and U2509 (N_2509,N_284,N_715);
nand U2510 (N_2510,N_633,N_1340);
nor U2511 (N_2511,N_1429,N_30);
nor U2512 (N_2512,N_1448,N_30);
nand U2513 (N_2513,N_1038,N_558);
and U2514 (N_2514,N_723,N_1236);
or U2515 (N_2515,N_612,N_396);
nand U2516 (N_2516,N_785,N_1323);
and U2517 (N_2517,N_1497,N_226);
and U2518 (N_2518,N_942,N_357);
nand U2519 (N_2519,N_13,N_1269);
nor U2520 (N_2520,N_1162,N_942);
nor U2521 (N_2521,N_1138,N_1039);
nor U2522 (N_2522,N_505,N_1132);
nor U2523 (N_2523,N_502,N_635);
and U2524 (N_2524,N_378,N_381);
or U2525 (N_2525,N_5,N_1323);
and U2526 (N_2526,N_735,N_462);
nand U2527 (N_2527,N_544,N_765);
nand U2528 (N_2528,N_285,N_876);
nor U2529 (N_2529,N_1221,N_317);
nor U2530 (N_2530,N_1263,N_844);
or U2531 (N_2531,N_1275,N_49);
or U2532 (N_2532,N_868,N_364);
nor U2533 (N_2533,N_899,N_355);
or U2534 (N_2534,N_494,N_1451);
nor U2535 (N_2535,N_401,N_1314);
or U2536 (N_2536,N_901,N_622);
and U2537 (N_2537,N_1036,N_562);
and U2538 (N_2538,N_693,N_17);
or U2539 (N_2539,N_838,N_835);
nor U2540 (N_2540,N_441,N_342);
or U2541 (N_2541,N_60,N_1106);
and U2542 (N_2542,N_330,N_233);
nand U2543 (N_2543,N_1062,N_447);
and U2544 (N_2544,N_1037,N_1301);
or U2545 (N_2545,N_572,N_325);
nor U2546 (N_2546,N_530,N_128);
nand U2547 (N_2547,N_1427,N_862);
and U2548 (N_2548,N_482,N_119);
nor U2549 (N_2549,N_333,N_1336);
nand U2550 (N_2550,N_1098,N_614);
or U2551 (N_2551,N_858,N_78);
nand U2552 (N_2552,N_334,N_352);
nand U2553 (N_2553,N_1363,N_492);
or U2554 (N_2554,N_795,N_1316);
or U2555 (N_2555,N_708,N_1068);
nor U2556 (N_2556,N_122,N_1376);
or U2557 (N_2557,N_734,N_1420);
and U2558 (N_2558,N_1372,N_1299);
nor U2559 (N_2559,N_1127,N_326);
nand U2560 (N_2560,N_597,N_922);
nor U2561 (N_2561,N_1420,N_1381);
nand U2562 (N_2562,N_285,N_1181);
nor U2563 (N_2563,N_1381,N_499);
nand U2564 (N_2564,N_538,N_1014);
or U2565 (N_2565,N_1365,N_579);
or U2566 (N_2566,N_155,N_258);
nor U2567 (N_2567,N_1258,N_1464);
nand U2568 (N_2568,N_933,N_1480);
or U2569 (N_2569,N_506,N_788);
and U2570 (N_2570,N_1433,N_88);
nand U2571 (N_2571,N_699,N_1104);
and U2572 (N_2572,N_1279,N_193);
or U2573 (N_2573,N_1274,N_800);
nor U2574 (N_2574,N_792,N_739);
and U2575 (N_2575,N_729,N_186);
or U2576 (N_2576,N_996,N_1457);
or U2577 (N_2577,N_784,N_527);
xor U2578 (N_2578,N_782,N_1019);
or U2579 (N_2579,N_811,N_264);
and U2580 (N_2580,N_1315,N_66);
nor U2581 (N_2581,N_162,N_315);
and U2582 (N_2582,N_45,N_22);
and U2583 (N_2583,N_1052,N_677);
and U2584 (N_2584,N_445,N_633);
or U2585 (N_2585,N_1489,N_1330);
and U2586 (N_2586,N_377,N_907);
and U2587 (N_2587,N_1171,N_1434);
xnor U2588 (N_2588,N_1403,N_285);
nor U2589 (N_2589,N_1072,N_1344);
nand U2590 (N_2590,N_469,N_970);
and U2591 (N_2591,N_1382,N_512);
or U2592 (N_2592,N_100,N_107);
nor U2593 (N_2593,N_894,N_1386);
nor U2594 (N_2594,N_166,N_123);
nor U2595 (N_2595,N_1253,N_1115);
or U2596 (N_2596,N_702,N_281);
nand U2597 (N_2597,N_1175,N_1414);
and U2598 (N_2598,N_333,N_1169);
or U2599 (N_2599,N_1370,N_1168);
nand U2600 (N_2600,N_524,N_906);
xor U2601 (N_2601,N_820,N_1290);
nor U2602 (N_2602,N_1469,N_1350);
nand U2603 (N_2603,N_836,N_890);
nand U2604 (N_2604,N_240,N_1099);
nor U2605 (N_2605,N_1456,N_1280);
and U2606 (N_2606,N_403,N_76);
or U2607 (N_2607,N_1135,N_1439);
nand U2608 (N_2608,N_144,N_532);
or U2609 (N_2609,N_566,N_1142);
nand U2610 (N_2610,N_40,N_42);
xnor U2611 (N_2611,N_886,N_90);
nor U2612 (N_2612,N_636,N_159);
xor U2613 (N_2613,N_726,N_649);
nand U2614 (N_2614,N_257,N_100);
xnor U2615 (N_2615,N_221,N_669);
nand U2616 (N_2616,N_1321,N_1059);
nor U2617 (N_2617,N_283,N_1202);
or U2618 (N_2618,N_479,N_690);
xor U2619 (N_2619,N_346,N_1169);
nand U2620 (N_2620,N_533,N_486);
nor U2621 (N_2621,N_1362,N_189);
or U2622 (N_2622,N_424,N_806);
nor U2623 (N_2623,N_478,N_1397);
or U2624 (N_2624,N_1237,N_72);
or U2625 (N_2625,N_290,N_1452);
xor U2626 (N_2626,N_683,N_1154);
nor U2627 (N_2627,N_1073,N_1445);
xnor U2628 (N_2628,N_715,N_323);
nand U2629 (N_2629,N_779,N_145);
nand U2630 (N_2630,N_1196,N_684);
nor U2631 (N_2631,N_364,N_1044);
nand U2632 (N_2632,N_23,N_459);
nand U2633 (N_2633,N_988,N_771);
nand U2634 (N_2634,N_367,N_971);
xor U2635 (N_2635,N_961,N_88);
nor U2636 (N_2636,N_1317,N_609);
nand U2637 (N_2637,N_1248,N_1061);
nor U2638 (N_2638,N_1243,N_101);
nor U2639 (N_2639,N_1249,N_545);
xor U2640 (N_2640,N_1317,N_565);
or U2641 (N_2641,N_1043,N_616);
nor U2642 (N_2642,N_326,N_671);
and U2643 (N_2643,N_771,N_1422);
and U2644 (N_2644,N_187,N_788);
or U2645 (N_2645,N_499,N_1452);
xnor U2646 (N_2646,N_256,N_940);
nor U2647 (N_2647,N_1042,N_1405);
nand U2648 (N_2648,N_876,N_740);
nand U2649 (N_2649,N_1281,N_119);
and U2650 (N_2650,N_922,N_1114);
and U2651 (N_2651,N_1356,N_730);
or U2652 (N_2652,N_1429,N_355);
nand U2653 (N_2653,N_742,N_485);
and U2654 (N_2654,N_105,N_659);
and U2655 (N_2655,N_1275,N_635);
nand U2656 (N_2656,N_1299,N_1435);
nand U2657 (N_2657,N_12,N_1141);
nor U2658 (N_2658,N_802,N_324);
xor U2659 (N_2659,N_1058,N_1336);
and U2660 (N_2660,N_101,N_920);
or U2661 (N_2661,N_1266,N_832);
xor U2662 (N_2662,N_107,N_461);
and U2663 (N_2663,N_887,N_287);
nor U2664 (N_2664,N_887,N_316);
nand U2665 (N_2665,N_325,N_25);
xor U2666 (N_2666,N_1499,N_1218);
and U2667 (N_2667,N_1183,N_411);
nand U2668 (N_2668,N_264,N_871);
or U2669 (N_2669,N_260,N_1170);
nor U2670 (N_2670,N_1130,N_1039);
nor U2671 (N_2671,N_488,N_69);
and U2672 (N_2672,N_1195,N_258);
nand U2673 (N_2673,N_722,N_1100);
and U2674 (N_2674,N_1291,N_297);
xnor U2675 (N_2675,N_441,N_13);
nor U2676 (N_2676,N_677,N_524);
nand U2677 (N_2677,N_397,N_1425);
and U2678 (N_2678,N_42,N_1053);
nor U2679 (N_2679,N_635,N_719);
and U2680 (N_2680,N_949,N_969);
xor U2681 (N_2681,N_94,N_10);
nor U2682 (N_2682,N_1020,N_385);
nand U2683 (N_2683,N_1040,N_907);
nand U2684 (N_2684,N_440,N_419);
nand U2685 (N_2685,N_1147,N_1209);
or U2686 (N_2686,N_638,N_933);
nand U2687 (N_2687,N_1133,N_1288);
nor U2688 (N_2688,N_832,N_250);
xnor U2689 (N_2689,N_1444,N_1390);
nand U2690 (N_2690,N_450,N_701);
and U2691 (N_2691,N_241,N_487);
xor U2692 (N_2692,N_1418,N_372);
nand U2693 (N_2693,N_1303,N_261);
nor U2694 (N_2694,N_693,N_635);
and U2695 (N_2695,N_992,N_548);
nor U2696 (N_2696,N_731,N_283);
and U2697 (N_2697,N_1318,N_790);
nand U2698 (N_2698,N_847,N_1164);
and U2699 (N_2699,N_675,N_743);
xor U2700 (N_2700,N_750,N_1274);
nor U2701 (N_2701,N_498,N_1304);
nand U2702 (N_2702,N_341,N_1495);
and U2703 (N_2703,N_880,N_389);
or U2704 (N_2704,N_1368,N_1045);
nand U2705 (N_2705,N_302,N_161);
nand U2706 (N_2706,N_1018,N_340);
and U2707 (N_2707,N_422,N_1024);
and U2708 (N_2708,N_1120,N_609);
nand U2709 (N_2709,N_818,N_851);
nand U2710 (N_2710,N_21,N_1479);
or U2711 (N_2711,N_47,N_1259);
nand U2712 (N_2712,N_1255,N_704);
and U2713 (N_2713,N_675,N_586);
and U2714 (N_2714,N_374,N_370);
or U2715 (N_2715,N_1140,N_1450);
nand U2716 (N_2716,N_696,N_1461);
nor U2717 (N_2717,N_78,N_1032);
and U2718 (N_2718,N_376,N_531);
nand U2719 (N_2719,N_1317,N_479);
nor U2720 (N_2720,N_802,N_913);
and U2721 (N_2721,N_870,N_386);
and U2722 (N_2722,N_59,N_951);
xor U2723 (N_2723,N_21,N_95);
nand U2724 (N_2724,N_1314,N_1229);
nor U2725 (N_2725,N_1430,N_599);
or U2726 (N_2726,N_364,N_1184);
nand U2727 (N_2727,N_739,N_1108);
nand U2728 (N_2728,N_930,N_1420);
nand U2729 (N_2729,N_741,N_425);
or U2730 (N_2730,N_696,N_382);
or U2731 (N_2731,N_811,N_477);
and U2732 (N_2732,N_516,N_365);
and U2733 (N_2733,N_141,N_831);
nor U2734 (N_2734,N_847,N_246);
xnor U2735 (N_2735,N_862,N_1129);
nor U2736 (N_2736,N_1413,N_612);
and U2737 (N_2737,N_135,N_696);
nand U2738 (N_2738,N_635,N_295);
or U2739 (N_2739,N_1187,N_1228);
or U2740 (N_2740,N_209,N_536);
or U2741 (N_2741,N_705,N_209);
or U2742 (N_2742,N_355,N_523);
nand U2743 (N_2743,N_369,N_1471);
or U2744 (N_2744,N_459,N_261);
or U2745 (N_2745,N_220,N_379);
and U2746 (N_2746,N_1166,N_636);
or U2747 (N_2747,N_299,N_312);
xor U2748 (N_2748,N_799,N_1192);
and U2749 (N_2749,N_39,N_667);
nand U2750 (N_2750,N_1311,N_502);
xor U2751 (N_2751,N_90,N_731);
xor U2752 (N_2752,N_1079,N_472);
or U2753 (N_2753,N_917,N_28);
and U2754 (N_2754,N_1304,N_869);
and U2755 (N_2755,N_816,N_737);
nor U2756 (N_2756,N_554,N_1126);
nor U2757 (N_2757,N_1358,N_418);
or U2758 (N_2758,N_1047,N_484);
nor U2759 (N_2759,N_21,N_467);
nand U2760 (N_2760,N_302,N_371);
and U2761 (N_2761,N_887,N_1252);
nand U2762 (N_2762,N_647,N_1449);
nand U2763 (N_2763,N_87,N_1188);
or U2764 (N_2764,N_889,N_40);
nor U2765 (N_2765,N_881,N_272);
nand U2766 (N_2766,N_835,N_1048);
nor U2767 (N_2767,N_850,N_857);
nand U2768 (N_2768,N_737,N_718);
or U2769 (N_2769,N_386,N_1404);
or U2770 (N_2770,N_402,N_148);
nand U2771 (N_2771,N_422,N_870);
nand U2772 (N_2772,N_900,N_231);
or U2773 (N_2773,N_536,N_961);
and U2774 (N_2774,N_420,N_451);
nand U2775 (N_2775,N_1026,N_18);
xnor U2776 (N_2776,N_888,N_960);
or U2777 (N_2777,N_1197,N_170);
or U2778 (N_2778,N_500,N_92);
and U2779 (N_2779,N_341,N_1106);
and U2780 (N_2780,N_953,N_613);
and U2781 (N_2781,N_799,N_698);
nand U2782 (N_2782,N_462,N_709);
nor U2783 (N_2783,N_356,N_127);
nand U2784 (N_2784,N_959,N_510);
nor U2785 (N_2785,N_790,N_1140);
and U2786 (N_2786,N_350,N_1427);
nand U2787 (N_2787,N_258,N_871);
or U2788 (N_2788,N_1150,N_590);
or U2789 (N_2789,N_652,N_1336);
and U2790 (N_2790,N_343,N_1310);
and U2791 (N_2791,N_95,N_1269);
and U2792 (N_2792,N_443,N_491);
xor U2793 (N_2793,N_203,N_635);
or U2794 (N_2794,N_1143,N_598);
nand U2795 (N_2795,N_162,N_400);
nand U2796 (N_2796,N_132,N_1365);
xnor U2797 (N_2797,N_809,N_1285);
or U2798 (N_2798,N_136,N_929);
nand U2799 (N_2799,N_1408,N_1012);
or U2800 (N_2800,N_1152,N_35);
nand U2801 (N_2801,N_499,N_1241);
and U2802 (N_2802,N_729,N_630);
xnor U2803 (N_2803,N_640,N_144);
nand U2804 (N_2804,N_624,N_415);
xor U2805 (N_2805,N_1198,N_624);
and U2806 (N_2806,N_1439,N_37);
and U2807 (N_2807,N_1353,N_1155);
or U2808 (N_2808,N_546,N_828);
nand U2809 (N_2809,N_940,N_1387);
nor U2810 (N_2810,N_440,N_1172);
or U2811 (N_2811,N_191,N_70);
nor U2812 (N_2812,N_884,N_1058);
nand U2813 (N_2813,N_391,N_644);
nand U2814 (N_2814,N_1289,N_126);
nor U2815 (N_2815,N_1462,N_1327);
xnor U2816 (N_2816,N_122,N_1220);
nand U2817 (N_2817,N_840,N_130);
nand U2818 (N_2818,N_1278,N_45);
or U2819 (N_2819,N_494,N_1234);
and U2820 (N_2820,N_711,N_1030);
or U2821 (N_2821,N_1485,N_232);
or U2822 (N_2822,N_1497,N_1128);
and U2823 (N_2823,N_1030,N_1416);
nand U2824 (N_2824,N_1426,N_997);
and U2825 (N_2825,N_619,N_683);
and U2826 (N_2826,N_590,N_584);
or U2827 (N_2827,N_401,N_1339);
or U2828 (N_2828,N_1344,N_575);
xnor U2829 (N_2829,N_462,N_792);
nor U2830 (N_2830,N_387,N_1442);
nand U2831 (N_2831,N_1359,N_1236);
nor U2832 (N_2832,N_1430,N_558);
nand U2833 (N_2833,N_630,N_1433);
nor U2834 (N_2834,N_1340,N_1271);
nand U2835 (N_2835,N_66,N_788);
nor U2836 (N_2836,N_773,N_820);
nand U2837 (N_2837,N_782,N_1257);
nor U2838 (N_2838,N_207,N_1288);
and U2839 (N_2839,N_634,N_1348);
or U2840 (N_2840,N_226,N_1089);
nand U2841 (N_2841,N_837,N_282);
xor U2842 (N_2842,N_1291,N_432);
nand U2843 (N_2843,N_572,N_1117);
or U2844 (N_2844,N_32,N_1425);
nand U2845 (N_2845,N_70,N_121);
nor U2846 (N_2846,N_1035,N_308);
nand U2847 (N_2847,N_835,N_120);
nor U2848 (N_2848,N_577,N_928);
or U2849 (N_2849,N_1370,N_1441);
or U2850 (N_2850,N_992,N_1413);
nand U2851 (N_2851,N_1064,N_803);
and U2852 (N_2852,N_299,N_727);
and U2853 (N_2853,N_388,N_538);
xnor U2854 (N_2854,N_1075,N_272);
nand U2855 (N_2855,N_663,N_1040);
or U2856 (N_2856,N_1318,N_1060);
and U2857 (N_2857,N_297,N_1499);
nor U2858 (N_2858,N_1120,N_955);
or U2859 (N_2859,N_590,N_507);
xor U2860 (N_2860,N_1054,N_166);
nor U2861 (N_2861,N_9,N_805);
nor U2862 (N_2862,N_30,N_600);
nor U2863 (N_2863,N_413,N_1123);
and U2864 (N_2864,N_1011,N_1060);
or U2865 (N_2865,N_1009,N_1304);
nor U2866 (N_2866,N_831,N_1074);
nor U2867 (N_2867,N_1042,N_1204);
or U2868 (N_2868,N_357,N_1018);
nand U2869 (N_2869,N_621,N_1242);
nor U2870 (N_2870,N_842,N_1168);
nand U2871 (N_2871,N_984,N_901);
nand U2872 (N_2872,N_1255,N_1190);
and U2873 (N_2873,N_585,N_361);
and U2874 (N_2874,N_683,N_657);
and U2875 (N_2875,N_410,N_104);
or U2876 (N_2876,N_663,N_1277);
or U2877 (N_2877,N_533,N_246);
and U2878 (N_2878,N_32,N_50);
or U2879 (N_2879,N_219,N_569);
nand U2880 (N_2880,N_1254,N_216);
nor U2881 (N_2881,N_670,N_6);
or U2882 (N_2882,N_855,N_1012);
or U2883 (N_2883,N_1413,N_897);
nor U2884 (N_2884,N_1426,N_1380);
or U2885 (N_2885,N_1282,N_1278);
nand U2886 (N_2886,N_257,N_1036);
and U2887 (N_2887,N_1396,N_36);
or U2888 (N_2888,N_508,N_827);
nor U2889 (N_2889,N_973,N_665);
xnor U2890 (N_2890,N_1411,N_1014);
or U2891 (N_2891,N_965,N_1154);
and U2892 (N_2892,N_15,N_1357);
or U2893 (N_2893,N_287,N_148);
or U2894 (N_2894,N_0,N_965);
or U2895 (N_2895,N_1272,N_357);
or U2896 (N_2896,N_1120,N_1160);
and U2897 (N_2897,N_568,N_720);
or U2898 (N_2898,N_892,N_15);
nand U2899 (N_2899,N_454,N_316);
or U2900 (N_2900,N_375,N_1182);
or U2901 (N_2901,N_992,N_352);
or U2902 (N_2902,N_1494,N_641);
and U2903 (N_2903,N_822,N_86);
and U2904 (N_2904,N_1271,N_11);
nor U2905 (N_2905,N_481,N_580);
or U2906 (N_2906,N_902,N_938);
nor U2907 (N_2907,N_896,N_554);
and U2908 (N_2908,N_1215,N_394);
nand U2909 (N_2909,N_731,N_1262);
nor U2910 (N_2910,N_237,N_1186);
nor U2911 (N_2911,N_438,N_1081);
xnor U2912 (N_2912,N_423,N_515);
and U2913 (N_2913,N_835,N_1039);
xnor U2914 (N_2914,N_219,N_629);
and U2915 (N_2915,N_380,N_1376);
nor U2916 (N_2916,N_275,N_211);
or U2917 (N_2917,N_206,N_1236);
and U2918 (N_2918,N_1052,N_1218);
or U2919 (N_2919,N_903,N_1001);
xnor U2920 (N_2920,N_1301,N_543);
and U2921 (N_2921,N_137,N_899);
or U2922 (N_2922,N_231,N_642);
nand U2923 (N_2923,N_56,N_8);
nand U2924 (N_2924,N_1198,N_560);
or U2925 (N_2925,N_1302,N_911);
and U2926 (N_2926,N_60,N_661);
nor U2927 (N_2927,N_56,N_593);
nor U2928 (N_2928,N_348,N_693);
or U2929 (N_2929,N_547,N_442);
and U2930 (N_2930,N_980,N_414);
and U2931 (N_2931,N_318,N_1031);
and U2932 (N_2932,N_1271,N_716);
nand U2933 (N_2933,N_276,N_982);
nor U2934 (N_2934,N_631,N_107);
nor U2935 (N_2935,N_425,N_59);
nand U2936 (N_2936,N_1123,N_688);
nor U2937 (N_2937,N_190,N_208);
and U2938 (N_2938,N_112,N_1478);
or U2939 (N_2939,N_1109,N_266);
and U2940 (N_2940,N_669,N_223);
nand U2941 (N_2941,N_260,N_321);
xor U2942 (N_2942,N_562,N_322);
or U2943 (N_2943,N_909,N_957);
and U2944 (N_2944,N_203,N_1467);
xor U2945 (N_2945,N_772,N_103);
xor U2946 (N_2946,N_1452,N_1042);
and U2947 (N_2947,N_1132,N_379);
and U2948 (N_2948,N_78,N_300);
and U2949 (N_2949,N_580,N_722);
nor U2950 (N_2950,N_555,N_1390);
nand U2951 (N_2951,N_1278,N_700);
and U2952 (N_2952,N_1100,N_778);
nor U2953 (N_2953,N_34,N_952);
and U2954 (N_2954,N_1454,N_1384);
and U2955 (N_2955,N_790,N_1150);
or U2956 (N_2956,N_947,N_1199);
nor U2957 (N_2957,N_591,N_1153);
nor U2958 (N_2958,N_1055,N_708);
nor U2959 (N_2959,N_19,N_579);
and U2960 (N_2960,N_77,N_846);
xor U2961 (N_2961,N_1323,N_996);
or U2962 (N_2962,N_809,N_885);
or U2963 (N_2963,N_803,N_391);
nor U2964 (N_2964,N_335,N_877);
and U2965 (N_2965,N_573,N_357);
nand U2966 (N_2966,N_604,N_1271);
or U2967 (N_2967,N_1315,N_912);
and U2968 (N_2968,N_1268,N_338);
and U2969 (N_2969,N_474,N_187);
nor U2970 (N_2970,N_1216,N_8);
nand U2971 (N_2971,N_995,N_58);
nor U2972 (N_2972,N_871,N_1141);
and U2973 (N_2973,N_391,N_523);
nand U2974 (N_2974,N_1165,N_387);
xnor U2975 (N_2975,N_211,N_319);
nand U2976 (N_2976,N_580,N_1414);
or U2977 (N_2977,N_162,N_171);
nand U2978 (N_2978,N_633,N_1079);
and U2979 (N_2979,N_417,N_423);
and U2980 (N_2980,N_71,N_309);
nor U2981 (N_2981,N_570,N_937);
nand U2982 (N_2982,N_743,N_868);
and U2983 (N_2983,N_99,N_399);
and U2984 (N_2984,N_308,N_597);
nor U2985 (N_2985,N_1401,N_1092);
and U2986 (N_2986,N_435,N_1184);
or U2987 (N_2987,N_1277,N_933);
and U2988 (N_2988,N_370,N_680);
and U2989 (N_2989,N_1495,N_535);
or U2990 (N_2990,N_287,N_1208);
and U2991 (N_2991,N_625,N_481);
or U2992 (N_2992,N_663,N_1396);
or U2993 (N_2993,N_704,N_502);
and U2994 (N_2994,N_479,N_1028);
nor U2995 (N_2995,N_772,N_1169);
nor U2996 (N_2996,N_260,N_39);
nor U2997 (N_2997,N_729,N_3);
nand U2998 (N_2998,N_30,N_324);
and U2999 (N_2999,N_679,N_834);
nand U3000 (N_3000,N_1985,N_2095);
and U3001 (N_3001,N_1918,N_2531);
nand U3002 (N_3002,N_2639,N_2084);
and U3003 (N_3003,N_2678,N_1696);
and U3004 (N_3004,N_2263,N_2010);
and U3005 (N_3005,N_1811,N_2922);
nor U3006 (N_3006,N_1856,N_1686);
xnor U3007 (N_3007,N_2816,N_2865);
nand U3008 (N_3008,N_1887,N_2723);
or U3009 (N_3009,N_1870,N_1847);
nand U3010 (N_3010,N_1627,N_1898);
nand U3011 (N_3011,N_1653,N_2251);
or U3012 (N_3012,N_2204,N_2536);
or U3013 (N_3013,N_2641,N_2066);
and U3014 (N_3014,N_2079,N_2601);
or U3015 (N_3015,N_2710,N_2008);
nor U3016 (N_3016,N_1867,N_2684);
nand U3017 (N_3017,N_2174,N_2383);
nor U3018 (N_3018,N_1664,N_2895);
nor U3019 (N_3019,N_1668,N_2915);
or U3020 (N_3020,N_2602,N_2725);
or U3021 (N_3021,N_2056,N_2506);
nand U3022 (N_3022,N_2041,N_2157);
or U3023 (N_3023,N_1950,N_2683);
nor U3024 (N_3024,N_2435,N_2075);
or U3025 (N_3025,N_1961,N_1715);
nand U3026 (N_3026,N_2637,N_1901);
or U3027 (N_3027,N_2061,N_1842);
or U3028 (N_3028,N_2447,N_2403);
or U3029 (N_3029,N_2134,N_1877);
or U3030 (N_3030,N_2476,N_1701);
xnor U3031 (N_3031,N_1769,N_2722);
and U3032 (N_3032,N_2546,N_2200);
and U3033 (N_3033,N_1751,N_1885);
or U3034 (N_3034,N_2630,N_2610);
or U3035 (N_3035,N_2269,N_2230);
or U3036 (N_3036,N_1682,N_2800);
and U3037 (N_3037,N_2340,N_2194);
or U3038 (N_3038,N_2677,N_2966);
or U3039 (N_3039,N_1576,N_1991);
and U3040 (N_3040,N_2648,N_2358);
xnor U3041 (N_3041,N_2125,N_2616);
or U3042 (N_3042,N_1880,N_1927);
nand U3043 (N_3043,N_2645,N_2604);
nor U3044 (N_3044,N_2261,N_1922);
xnor U3045 (N_3045,N_2647,N_2117);
or U3046 (N_3046,N_2283,N_2381);
nor U3047 (N_3047,N_1539,N_2896);
nor U3048 (N_3048,N_2523,N_2394);
nor U3049 (N_3049,N_2555,N_2595);
nor U3050 (N_3050,N_2196,N_1772);
nor U3051 (N_3051,N_1655,N_2003);
nand U3052 (N_3052,N_2092,N_2467);
or U3053 (N_3053,N_1626,N_2989);
or U3054 (N_3054,N_1502,N_1999);
and U3055 (N_3055,N_2369,N_1910);
nand U3056 (N_3056,N_2347,N_1824);
or U3057 (N_3057,N_2797,N_1529);
and U3058 (N_3058,N_2267,N_2016);
and U3059 (N_3059,N_2950,N_2408);
or U3060 (N_3060,N_2191,N_1896);
and U3061 (N_3061,N_1695,N_2480);
and U3062 (N_3062,N_1526,N_1992);
xor U3063 (N_3063,N_1959,N_2748);
xor U3064 (N_3064,N_2671,N_2691);
nor U3065 (N_3065,N_2132,N_2022);
or U3066 (N_3066,N_2605,N_2786);
nor U3067 (N_3067,N_2873,N_2741);
xnor U3068 (N_3068,N_1524,N_2568);
and U3069 (N_3069,N_2809,N_2757);
xor U3070 (N_3070,N_2736,N_2864);
or U3071 (N_3071,N_2378,N_2057);
nand U3072 (N_3072,N_1625,N_2212);
nand U3073 (N_3073,N_2571,N_2695);
nor U3074 (N_3074,N_1844,N_2799);
and U3075 (N_3075,N_1796,N_2238);
and U3076 (N_3076,N_2493,N_2301);
or U3077 (N_3077,N_2428,N_2640);
and U3078 (N_3078,N_1749,N_2789);
and U3079 (N_3079,N_2747,N_1754);
xnor U3080 (N_3080,N_2072,N_2588);
or U3081 (N_3081,N_2030,N_1591);
xnor U3082 (N_3082,N_2686,N_1638);
and U3083 (N_3083,N_2193,N_2430);
and U3084 (N_3084,N_2367,N_2221);
or U3085 (N_3085,N_2266,N_1702);
nand U3086 (N_3086,N_1672,N_1786);
and U3087 (N_3087,N_2004,N_2107);
nor U3088 (N_3088,N_2356,N_2908);
nand U3089 (N_3089,N_1601,N_1590);
nand U3090 (N_3090,N_1639,N_1814);
xnor U3091 (N_3091,N_2877,N_2416);
and U3092 (N_3092,N_2206,N_1719);
and U3093 (N_3093,N_1736,N_2670);
xnor U3094 (N_3094,N_1859,N_2622);
and U3095 (N_3095,N_2051,N_1596);
or U3096 (N_3096,N_2243,N_1516);
or U3097 (N_3097,N_2456,N_2275);
nor U3098 (N_3098,N_1511,N_2596);
nand U3099 (N_3099,N_2763,N_2461);
nand U3100 (N_3100,N_2302,N_2071);
and U3101 (N_3101,N_1865,N_2594);
nor U3102 (N_3102,N_2669,N_2364);
nand U3103 (N_3103,N_2629,N_2309);
or U3104 (N_3104,N_2838,N_2498);
nand U3105 (N_3105,N_1504,N_2374);
or U3106 (N_3106,N_2017,N_2912);
and U3107 (N_3107,N_2697,N_1544);
and U3108 (N_3108,N_1651,N_2389);
nand U3109 (N_3109,N_2516,N_2188);
and U3110 (N_3110,N_1892,N_1712);
nand U3111 (N_3111,N_2563,N_1911);
and U3112 (N_3112,N_1734,N_2177);
and U3113 (N_3113,N_1611,N_1993);
and U3114 (N_3114,N_2636,N_2661);
nor U3115 (N_3115,N_2527,N_2070);
and U3116 (N_3116,N_2719,N_1650);
nand U3117 (N_3117,N_2611,N_2796);
or U3118 (N_3118,N_2119,N_2808);
nand U3119 (N_3119,N_2828,N_2603);
and U3120 (N_3120,N_2933,N_2110);
xor U3121 (N_3121,N_2843,N_1642);
or U3122 (N_3122,N_2772,N_1602);
or U3123 (N_3123,N_1966,N_2449);
or U3124 (N_3124,N_2305,N_2291);
nand U3125 (N_3125,N_1727,N_2703);
nor U3126 (N_3126,N_1753,N_2240);
nor U3127 (N_3127,N_2373,N_1723);
xnor U3128 (N_3128,N_1989,N_2902);
nand U3129 (N_3129,N_1967,N_2341);
nand U3130 (N_3130,N_1775,N_2500);
nand U3131 (N_3131,N_1770,N_2566);
or U3132 (N_3132,N_1570,N_2730);
and U3133 (N_3133,N_2939,N_2286);
nand U3134 (N_3134,N_2402,N_1803);
or U3135 (N_3135,N_2100,N_2623);
nor U3136 (N_3136,N_2790,N_2054);
nand U3137 (N_3137,N_2372,N_2544);
or U3138 (N_3138,N_2984,N_2466);
nand U3139 (N_3139,N_1660,N_1534);
nand U3140 (N_3140,N_1584,N_2149);
nand U3141 (N_3141,N_2040,N_1517);
nor U3142 (N_3142,N_2087,N_2929);
or U3143 (N_3143,N_2650,N_2998);
and U3144 (N_3144,N_1899,N_1538);
and U3145 (N_3145,N_1741,N_2781);
nand U3146 (N_3146,N_2919,N_1860);
and U3147 (N_3147,N_1799,N_1748);
nor U3148 (N_3148,N_2976,N_2580);
nand U3149 (N_3149,N_1681,N_1585);
or U3150 (N_3150,N_1980,N_1873);
nand U3151 (N_3151,N_2482,N_2672);
or U3152 (N_3152,N_1781,N_2205);
nor U3153 (N_3153,N_1560,N_2570);
and U3154 (N_3154,N_1667,N_2752);
nor U3155 (N_3155,N_2209,N_1757);
and U3156 (N_3156,N_2438,N_2533);
nand U3157 (N_3157,N_2012,N_1863);
nand U3158 (N_3158,N_2437,N_2944);
or U3159 (N_3159,N_2208,N_1931);
xor U3160 (N_3160,N_2158,N_2459);
or U3161 (N_3161,N_2176,N_1872);
and U3162 (N_3162,N_2185,N_2658);
and U3163 (N_3163,N_2285,N_2328);
nand U3164 (N_3164,N_2577,N_2478);
nand U3165 (N_3165,N_2281,N_2143);
nor U3166 (N_3166,N_2962,N_2551);
nand U3167 (N_3167,N_2241,N_2236);
nor U3168 (N_3168,N_1735,N_2052);
or U3169 (N_3169,N_1850,N_1548);
or U3170 (N_3170,N_2019,N_2308);
nand U3171 (N_3171,N_2558,N_2928);
nand U3172 (N_3172,N_2625,N_2830);
nor U3173 (N_3173,N_2848,N_2810);
or U3174 (N_3174,N_1646,N_2632);
nand U3175 (N_3175,N_1595,N_2044);
xor U3176 (N_3176,N_1909,N_1661);
nor U3177 (N_3177,N_1897,N_2363);
nand U3178 (N_3178,N_1503,N_2918);
or U3179 (N_3179,N_1636,N_2298);
nand U3180 (N_3180,N_2831,N_2885);
nor U3181 (N_3181,N_1780,N_2979);
and U3182 (N_3182,N_2218,N_2349);
and U3183 (N_3183,N_2362,N_1588);
nand U3184 (N_3184,N_2982,N_2264);
and U3185 (N_3185,N_1614,N_1834);
nand U3186 (N_3186,N_1798,N_2954);
or U3187 (N_3187,N_2643,N_2320);
nor U3188 (N_3188,N_1641,N_2495);
nand U3189 (N_3189,N_2699,N_1849);
nand U3190 (N_3190,N_2122,N_1935);
nand U3191 (N_3191,N_2901,N_2295);
nor U3192 (N_3192,N_2313,N_1581);
or U3193 (N_3193,N_1916,N_2652);
and U3194 (N_3194,N_1890,N_2225);
and U3195 (N_3195,N_1843,N_1518);
nor U3196 (N_3196,N_2762,N_1706);
or U3197 (N_3197,N_1527,N_1658);
and U3198 (N_3198,N_1501,N_2910);
or U3199 (N_3199,N_1688,N_1903);
nand U3200 (N_3200,N_2554,N_2080);
nand U3201 (N_3201,N_2514,N_2888);
and U3202 (N_3202,N_2897,N_2376);
and U3203 (N_3203,N_2862,N_2742);
nand U3204 (N_3204,N_2379,N_1981);
and U3205 (N_3205,N_1963,N_2573);
xor U3206 (N_3206,N_1833,N_1506);
and U3207 (N_3207,N_2951,N_1571);
nand U3208 (N_3208,N_2245,N_1854);
and U3209 (N_3209,N_1866,N_1561);
nand U3210 (N_3210,N_1808,N_2469);
and U3211 (N_3211,N_1505,N_2065);
nor U3212 (N_3212,N_1851,N_2835);
nand U3213 (N_3213,N_2525,N_1716);
and U3214 (N_3214,N_1731,N_1820);
and U3215 (N_3215,N_2222,N_2260);
and U3216 (N_3216,N_2685,N_2673);
nand U3217 (N_3217,N_2971,N_2322);
and U3218 (N_3218,N_2869,N_2314);
nand U3219 (N_3219,N_2633,N_2593);
or U3220 (N_3220,N_2986,N_1553);
or U3221 (N_3221,N_2534,N_2708);
nor U3222 (N_3222,N_2776,N_1745);
and U3223 (N_3223,N_2907,N_2964);
or U3224 (N_3224,N_2987,N_2583);
nand U3225 (N_3225,N_2854,N_2598);
nor U3226 (N_3226,N_2088,N_1635);
nor U3227 (N_3227,N_2352,N_2168);
nor U3228 (N_3228,N_2137,N_1816);
and U3229 (N_3229,N_2473,N_2696);
and U3230 (N_3230,N_1746,N_2935);
nand U3231 (N_3231,N_2837,N_2660);
nor U3232 (N_3232,N_1829,N_1938);
or U3233 (N_3233,N_1965,N_1555);
and U3234 (N_3234,N_1940,N_2359);
nand U3235 (N_3235,N_2009,N_2280);
nor U3236 (N_3236,N_2769,N_2543);
xor U3237 (N_3237,N_2759,N_1827);
or U3238 (N_3238,N_2900,N_2425);
or U3239 (N_3239,N_2423,N_1879);
nor U3240 (N_3240,N_1633,N_1687);
xor U3241 (N_3241,N_1519,N_2475);
or U3242 (N_3242,N_2248,N_2300);
or U3243 (N_3243,N_2572,N_2845);
nand U3244 (N_3244,N_2945,N_2199);
nor U3245 (N_3245,N_2892,N_2085);
or U3246 (N_3246,N_1637,N_2733);
nand U3247 (N_3247,N_1883,N_2999);
xnor U3248 (N_3248,N_2180,N_1670);
xnor U3249 (N_3249,N_2136,N_2909);
and U3250 (N_3250,N_2409,N_2496);
nor U3251 (N_3251,N_1825,N_2932);
or U3252 (N_3252,N_2289,N_2734);
or U3253 (N_3253,N_1747,N_1709);
and U3254 (N_3254,N_2846,N_1648);
xnor U3255 (N_3255,N_1975,N_2181);
and U3256 (N_3256,N_1738,N_2528);
nand U3257 (N_3257,N_2344,N_1693);
nor U3258 (N_3258,N_2689,N_2756);
or U3259 (N_3259,N_2118,N_1703);
nor U3260 (N_3260,N_2224,N_2411);
nand U3261 (N_3261,N_2779,N_1623);
xor U3262 (N_3262,N_2483,N_1630);
or U3263 (N_3263,N_2728,N_2624);
xor U3264 (N_3264,N_2538,N_2096);
or U3265 (N_3265,N_1926,N_1948);
xor U3266 (N_3266,N_2537,N_1766);
or U3267 (N_3267,N_2668,N_2780);
nand U3268 (N_3268,N_2532,N_2899);
nand U3269 (N_3269,N_2863,N_2774);
nor U3270 (N_3270,N_2812,N_2975);
and U3271 (N_3271,N_1944,N_1868);
nand U3272 (N_3272,N_1783,N_2413);
nor U3273 (N_3273,N_2342,N_2766);
nand U3274 (N_3274,N_2278,N_1592);
nand U3275 (N_3275,N_1606,N_2764);
nor U3276 (N_3276,N_2294,N_1970);
and U3277 (N_3277,N_1572,N_2709);
or U3278 (N_3278,N_2424,N_2108);
and U3279 (N_3279,N_1542,N_2114);
nor U3280 (N_3280,N_2046,N_2343);
xor U3281 (N_3281,N_2323,N_2020);
nor U3282 (N_3282,N_2244,N_2214);
or U3283 (N_3283,N_2631,N_2141);
nand U3284 (N_3284,N_1855,N_2621);
nor U3285 (N_3285,N_2913,N_1562);
and U3286 (N_3286,N_1713,N_1628);
or U3287 (N_3287,N_1612,N_1622);
nand U3288 (N_3288,N_2327,N_2128);
nand U3289 (N_3289,N_2732,N_2811);
and U3290 (N_3290,N_2740,N_2911);
nor U3291 (N_3291,N_2013,N_2524);
and U3292 (N_3292,N_2421,N_1724);
nor U3293 (N_3293,N_2518,N_2513);
or U3294 (N_3294,N_2607,N_2189);
nand U3295 (N_3295,N_2242,N_1788);
nand U3296 (N_3296,N_2564,N_2914);
nor U3297 (N_3297,N_2960,N_2023);
and U3298 (N_3298,N_2250,N_2958);
and U3299 (N_3299,N_2039,N_2981);
nand U3300 (N_3300,N_2649,N_2167);
xnor U3301 (N_3301,N_2693,N_1752);
or U3302 (N_3302,N_2934,N_2113);
nor U3303 (N_3303,N_2098,N_1894);
nand U3304 (N_3304,N_1604,N_2959);
xor U3305 (N_3305,N_1558,N_1976);
or U3306 (N_3306,N_2211,N_2827);
nand U3307 (N_3307,N_1832,N_2824);
xnor U3308 (N_3308,N_2879,N_2656);
nand U3309 (N_3309,N_1846,N_2161);
and U3310 (N_3310,N_2777,N_2317);
or U3311 (N_3311,N_2116,N_2585);
and U3312 (N_3312,N_2600,N_2968);
nor U3313 (N_3313,N_2850,N_2706);
or U3314 (N_3314,N_2399,N_1669);
and U3315 (N_3315,N_2694,N_2952);
and U3316 (N_3316,N_2169,N_2599);
or U3317 (N_3317,N_1972,N_2985);
and U3318 (N_3318,N_1678,N_2924);
nand U3319 (N_3319,N_2179,N_1822);
nand U3320 (N_3320,N_2081,N_2657);
nand U3321 (N_3321,N_2626,N_2817);
nor U3322 (N_3322,N_2454,N_1861);
nor U3323 (N_3323,N_1684,N_2529);
nor U3324 (N_3324,N_2111,N_1705);
nor U3325 (N_3325,N_1760,N_1968);
nor U3326 (N_3326,N_1500,N_2035);
xor U3327 (N_3327,N_1891,N_2923);
or U3328 (N_3328,N_1522,N_2388);
or U3329 (N_3329,N_1532,N_2487);
and U3330 (N_3330,N_1521,N_1722);
nor U3331 (N_3331,N_2033,N_2679);
nand U3332 (N_3332,N_1513,N_2059);
or U3333 (N_3333,N_1986,N_2450);
and U3334 (N_3334,N_2953,N_2802);
or U3335 (N_3335,N_1563,N_1996);
or U3336 (N_3336,N_1895,N_1552);
or U3337 (N_3337,N_2463,N_2511);
nand U3338 (N_3338,N_1593,N_2228);
or U3339 (N_3339,N_2018,N_1815);
nand U3340 (N_3340,N_1728,N_1774);
and U3341 (N_3341,N_1654,N_2472);
nor U3342 (N_3342,N_1945,N_2468);
or U3343 (N_3343,N_2332,N_2721);
and U3344 (N_3344,N_1919,N_2880);
or U3345 (N_3345,N_2775,N_2943);
and U3346 (N_3346,N_2874,N_1512);
nand U3347 (N_3347,N_1920,N_1946);
nand U3348 (N_3348,N_1974,N_2026);
or U3349 (N_3349,N_2284,N_1644);
and U3350 (N_3350,N_2821,N_2099);
and U3351 (N_3351,N_2891,N_2234);
or U3352 (N_3352,N_2159,N_2872);
or U3353 (N_3353,N_2584,N_2271);
nor U3354 (N_3354,N_2589,N_1795);
nand U3355 (N_3355,N_1762,N_2505);
and U3356 (N_3356,N_1589,N_2047);
xor U3357 (N_3357,N_2431,N_2484);
and U3358 (N_3358,N_2833,N_2963);
and U3359 (N_3359,N_2094,N_2702);
or U3360 (N_3360,N_1862,N_1685);
nor U3361 (N_3361,N_2207,N_2638);
and U3362 (N_3362,N_1771,N_2990);
nand U3363 (N_3363,N_2792,N_2049);
nand U3364 (N_3364,N_1597,N_1507);
and U3365 (N_3365,N_2414,N_2365);
xnor U3366 (N_3366,N_1573,N_2839);
and U3367 (N_3367,N_2793,N_1806);
and U3368 (N_3368,N_1928,N_1907);
and U3369 (N_3369,N_2028,N_2307);
or U3370 (N_3370,N_2938,N_2876);
nor U3371 (N_3371,N_1789,N_2445);
and U3372 (N_3372,N_1740,N_2692);
nand U3373 (N_3373,N_1540,N_2665);
or U3374 (N_3374,N_1836,N_1982);
or U3375 (N_3375,N_2078,N_1971);
nor U3376 (N_3376,N_2259,N_2510);
and U3377 (N_3377,N_2502,N_2316);
or U3378 (N_3378,N_2973,N_1707);
and U3379 (N_3379,N_2813,N_2994);
and U3380 (N_3380,N_1881,N_1657);
nand U3381 (N_3381,N_1805,N_2898);
or U3382 (N_3382,N_2074,N_2716);
or U3383 (N_3383,N_2273,N_2216);
xnor U3384 (N_3384,N_1690,N_2714);
or U3385 (N_3385,N_2509,N_2060);
nand U3386 (N_3386,N_2458,N_1675);
or U3387 (N_3387,N_2457,N_1952);
xnor U3388 (N_3388,N_2097,N_2612);
and U3389 (N_3389,N_1726,N_2045);
nand U3390 (N_3390,N_2252,N_1624);
or U3391 (N_3391,N_2247,N_2642);
or U3392 (N_3392,N_2745,N_1776);
and U3393 (N_3393,N_2042,N_2920);
and U3394 (N_3394,N_1810,N_1694);
nor U3395 (N_3395,N_1878,N_1797);
nand U3396 (N_3396,N_2488,N_2257);
and U3397 (N_3397,N_1720,N_2822);
nand U3398 (N_3398,N_2718,N_2319);
or U3399 (N_3399,N_2115,N_2829);
and U3400 (N_3400,N_1621,N_2031);
nor U3401 (N_3401,N_2350,N_1765);
nand U3402 (N_3402,N_2520,N_2836);
or U3403 (N_3403,N_1759,N_2265);
nand U3404 (N_3404,N_2007,N_1857);
nor U3405 (N_3405,N_2490,N_1826);
or U3406 (N_3406,N_2858,N_2682);
and U3407 (N_3407,N_1932,N_1665);
nand U3408 (N_3408,N_2299,N_2552);
nor U3409 (N_3409,N_1768,N_2120);
and U3410 (N_3410,N_2217,N_2256);
nand U3411 (N_3411,N_1886,N_1676);
and U3412 (N_3412,N_2597,N_2991);
nand U3413 (N_3413,N_2674,N_2337);
nor U3414 (N_3414,N_1575,N_2417);
nand U3415 (N_3415,N_2315,N_2700);
nand U3416 (N_3416,N_2942,N_2561);
nand U3417 (N_3417,N_2375,N_2470);
or U3418 (N_3418,N_1912,N_1947);
or U3419 (N_3419,N_2330,N_1997);
nand U3420 (N_3420,N_1779,N_2288);
and U3421 (N_3421,N_2794,N_1750);
and U3422 (N_3422,N_2492,N_2698);
nand U3423 (N_3423,N_2878,N_1618);
or U3424 (N_3424,N_1742,N_1547);
nand U3425 (N_3425,N_2530,N_1743);
nand U3426 (N_3426,N_2883,N_2832);
nand U3427 (N_3427,N_1608,N_1787);
nand U3428 (N_3428,N_1848,N_1988);
nor U3429 (N_3429,N_1958,N_2032);
or U3430 (N_3430,N_2894,N_1537);
nor U3431 (N_3431,N_2983,N_2433);
and U3432 (N_3432,N_1594,N_2972);
xor U3433 (N_3433,N_1730,N_2329);
nor U3434 (N_3434,N_2659,N_1884);
nor U3435 (N_3435,N_1964,N_1640);
nand U3436 (N_3436,N_1845,N_1755);
xnor U3437 (N_3437,N_2170,N_1804);
nand U3438 (N_3438,N_1613,N_1528);
xnor U3439 (N_3439,N_2961,N_1793);
xor U3440 (N_3440,N_2936,N_2773);
and U3441 (N_3441,N_2575,N_2574);
and U3442 (N_3442,N_1807,N_2644);
nand U3443 (N_3443,N_2664,N_1679);
xnor U3444 (N_3444,N_2608,N_1582);
xnor U3445 (N_3445,N_2171,N_1875);
nand U3446 (N_3446,N_2420,N_2014);
or U3447 (N_3447,N_1744,N_2549);
nand U3448 (N_3448,N_1869,N_2705);
nor U3449 (N_3449,N_2771,N_2393);
xnor U3450 (N_3450,N_2153,N_1689);
or U3451 (N_3451,N_2744,N_1782);
nand U3452 (N_3452,N_2321,N_2582);
or U3453 (N_3453,N_1605,N_2784);
and U3454 (N_3454,N_2460,N_2548);
and U3455 (N_3455,N_2162,N_2881);
nor U3456 (N_3456,N_1671,N_2064);
and U3457 (N_3457,N_2750,N_1990);
xor U3458 (N_3458,N_2034,N_2201);
nor U3459 (N_3459,N_2615,N_2351);
and U3460 (N_3460,N_1794,N_2226);
and U3461 (N_3461,N_2814,N_2729);
nor U3462 (N_3462,N_1510,N_2390);
and U3463 (N_3463,N_1554,N_2819);
xor U3464 (N_3464,N_2334,N_2795);
xnor U3465 (N_3465,N_2818,N_1737);
or U3466 (N_3466,N_1652,N_1680);
or U3467 (N_3467,N_2720,N_2142);
or U3468 (N_3468,N_2178,N_2727);
or U3469 (N_3469,N_1580,N_2852);
or U3470 (N_3470,N_2997,N_2905);
nor U3471 (N_3471,N_2290,N_2105);
nand U3472 (N_3472,N_1837,N_1923);
xor U3473 (N_3473,N_1564,N_2474);
nor U3474 (N_3474,N_1556,N_2195);
and U3475 (N_3475,N_2426,N_2804);
and U3476 (N_3476,N_2823,N_1545);
nor U3477 (N_3477,N_2190,N_1821);
and U3478 (N_3478,N_2724,N_2387);
and U3479 (N_3479,N_2444,N_2002);
or U3480 (N_3480,N_1708,N_2377);
and U3481 (N_3481,N_2385,N_2182);
nand U3482 (N_3482,N_2073,N_2540);
xor U3483 (N_3483,N_2613,N_2521);
or U3484 (N_3484,N_1525,N_1934);
nand U3485 (N_3485,N_2735,N_2653);
nand U3486 (N_3486,N_1536,N_1508);
or U3487 (N_3487,N_2941,N_2210);
nand U3488 (N_3488,N_2688,N_1914);
nor U3489 (N_3489,N_2133,N_2738);
and U3490 (N_3490,N_2627,N_2917);
or U3491 (N_3491,N_2834,N_2371);
nand U3492 (N_3492,N_1721,N_2277);
or U3493 (N_3493,N_1913,N_2336);
nor U3494 (N_3494,N_1809,N_2076);
and U3495 (N_3495,N_2712,N_1578);
nand U3496 (N_3496,N_2711,N_1586);
and U3497 (N_3497,N_2067,N_2274);
or U3498 (N_3498,N_2089,N_2324);
or U3499 (N_3499,N_2464,N_1643);
nand U3500 (N_3500,N_2384,N_1520);
and U3501 (N_3501,N_1790,N_2215);
and U3502 (N_3502,N_2586,N_1647);
nand U3503 (N_3503,N_2499,N_1831);
nand U3504 (N_3504,N_2654,N_1714);
or U3505 (N_3505,N_2889,N_1813);
xnor U3506 (N_3506,N_2011,N_1733);
nor U3507 (N_3507,N_1541,N_2893);
nand U3508 (N_3508,N_2392,N_2859);
nand U3509 (N_3509,N_1951,N_1515);
or U3510 (N_3510,N_2556,N_2036);
xor U3511 (N_3511,N_2440,N_2494);
or U3512 (N_3512,N_1607,N_2992);
nor U3513 (N_3513,N_2198,N_1761);
or U3514 (N_3514,N_2931,N_2760);
and U3515 (N_3515,N_1792,N_2853);
or U3516 (N_3516,N_2000,N_1549);
nand U3517 (N_3517,N_1939,N_1929);
and U3518 (N_3518,N_2788,N_1864);
nand U3519 (N_3519,N_2481,N_1717);
xnor U3520 (N_3520,N_2262,N_2995);
nor U3521 (N_3521,N_2522,N_2292);
and U3522 (N_3522,N_1523,N_2121);
nor U3523 (N_3523,N_2357,N_2006);
nand U3524 (N_3524,N_1533,N_2753);
nand U3525 (N_3525,N_2184,N_2380);
xnor U3526 (N_3526,N_2948,N_1530);
nor U3527 (N_3527,N_2965,N_2847);
and U3528 (N_3528,N_2152,N_2254);
nor U3529 (N_3529,N_1603,N_2579);
or U3530 (N_3530,N_2326,N_2310);
or U3531 (N_3531,N_2197,N_1632);
nand U3532 (N_3532,N_2366,N_2957);
or U3533 (N_3533,N_2485,N_2055);
nor U3534 (N_3534,N_1711,N_2400);
nor U3535 (N_3535,N_2857,N_1874);
or U3536 (N_3536,N_2628,N_2842);
and U3537 (N_3537,N_2717,N_2591);
or U3538 (N_3538,N_1677,N_2993);
nor U3539 (N_3539,N_1819,N_2526);
nor U3540 (N_3540,N_2758,N_2050);
nand U3541 (N_3541,N_1620,N_2930);
nor U3542 (N_3542,N_2446,N_2884);
nand U3543 (N_3543,N_1942,N_1773);
and U3544 (N_3544,N_2969,N_1882);
nor U3545 (N_3545,N_2429,N_2109);
nand U3546 (N_3546,N_2124,N_2501);
nor U3547 (N_3547,N_1917,N_2560);
nand U3548 (N_3548,N_2354,N_1767);
and U3549 (N_3549,N_1609,N_2015);
and U3550 (N_3550,N_2229,N_2681);
nand U3551 (N_3551,N_2436,N_2826);
nand U3552 (N_3552,N_2726,N_2663);
nand U3553 (N_3553,N_2123,N_2077);
nor U3554 (N_3554,N_2606,N_1998);
nor U3555 (N_3555,N_2233,N_1598);
nor U3556 (N_3556,N_1756,N_2068);
or U3557 (N_3557,N_2441,N_2707);
and U3558 (N_3558,N_1656,N_2849);
nor U3559 (N_3559,N_2249,N_2785);
and U3560 (N_3560,N_2967,N_2844);
and U3561 (N_3561,N_2338,N_2970);
nor U3562 (N_3562,N_1583,N_2557);
and U3563 (N_3563,N_1900,N_2140);
nand U3564 (N_3564,N_1888,N_1784);
or U3565 (N_3565,N_2186,N_2882);
nand U3566 (N_3566,N_1777,N_2940);
or U3567 (N_3567,N_1994,N_1666);
and U3568 (N_3568,N_1710,N_2618);
or U3569 (N_3569,N_2988,N_2405);
nand U3570 (N_3570,N_2279,N_1969);
xor U3571 (N_3571,N_2861,N_2386);
or U3572 (N_3572,N_2553,N_2739);
xor U3573 (N_3573,N_2422,N_2025);
nand U3574 (N_3574,N_2956,N_2165);
and U3575 (N_3575,N_1764,N_2287);
nor U3576 (N_3576,N_2325,N_1812);
nor U3577 (N_3577,N_1852,N_2801);
xor U3578 (N_3578,N_2255,N_2173);
nand U3579 (N_3579,N_2253,N_2304);
or U3580 (N_3580,N_2127,N_1839);
nand U3581 (N_3581,N_1718,N_2239);
xnor U3582 (N_3582,N_2227,N_1841);
and U3583 (N_3583,N_1871,N_2946);
and U3584 (N_3584,N_1908,N_2667);
nor U3585 (N_3585,N_1941,N_2130);
or U3586 (N_3586,N_2559,N_2955);
nand U3587 (N_3587,N_2886,N_2086);
nand U3588 (N_3588,N_2419,N_2980);
or U3589 (N_3589,N_2401,N_2160);
nor U3590 (N_3590,N_2761,N_2486);
nor U3591 (N_3591,N_2192,N_2112);
nand U3592 (N_3592,N_2448,N_1791);
and U3593 (N_3593,N_1698,N_1763);
nand U3594 (N_3594,N_2138,N_1566);
and U3595 (N_3595,N_2868,N_1954);
and U3596 (N_3596,N_1957,N_2974);
nand U3597 (N_3597,N_1995,N_2455);
nand U3598 (N_3598,N_2101,N_1587);
or U3599 (N_3599,N_1631,N_1984);
nand U3600 (N_3600,N_2038,N_1739);
and U3601 (N_3601,N_2815,N_2202);
xor U3602 (N_3602,N_2432,N_2798);
or U3603 (N_3603,N_2479,N_2001);
and U3604 (N_3604,N_2272,N_1983);
nand U3605 (N_3605,N_2183,N_2154);
or U3606 (N_3606,N_2751,N_2787);
nand U3607 (N_3607,N_1617,N_2451);
nand U3608 (N_3608,N_2415,N_1629);
nor U3609 (N_3609,N_2303,N_2144);
nand U3610 (N_3610,N_2737,N_2690);
and U3611 (N_3611,N_1559,N_1943);
nand U3612 (N_3612,N_2867,N_1692);
and U3613 (N_3613,N_2148,N_2102);
nand U3614 (N_3614,N_2806,N_2395);
and U3615 (N_3615,N_2512,N_1557);
or U3616 (N_3616,N_2620,N_2172);
and U3617 (N_3617,N_2397,N_2765);
and U3618 (N_3618,N_1823,N_2361);
nand U3619 (N_3619,N_2231,N_1785);
nand U3620 (N_3620,N_2021,N_1978);
and U3621 (N_3621,N_2545,N_2335);
or U3622 (N_3622,N_1933,N_2043);
nand U3623 (N_3623,N_2346,N_1579);
and U3624 (N_3624,N_2609,N_1725);
or U3625 (N_3625,N_1616,N_2410);
nand U3626 (N_3626,N_2567,N_2145);
nor U3627 (N_3627,N_2398,N_2701);
nand U3628 (N_3628,N_1691,N_2825);
nand U3629 (N_3629,N_2462,N_2687);
or U3630 (N_3630,N_2519,N_1700);
xnor U3631 (N_3631,N_2662,N_2855);
nand U3632 (N_3632,N_2311,N_2333);
nand U3633 (N_3633,N_2048,N_2949);
nand U3634 (N_3634,N_2666,N_1550);
nand U3635 (N_3635,N_2535,N_2407);
nand U3636 (N_3636,N_1830,N_2005);
and U3637 (N_3637,N_2617,N_1645);
nand U3638 (N_3638,N_2166,N_2439);
or U3639 (N_3639,N_2542,N_1904);
xnor U3640 (N_3640,N_2477,N_2406);
nand U3641 (N_3641,N_1853,N_2927);
and U3642 (N_3642,N_2270,N_2465);
nor U3643 (N_3643,N_1924,N_2651);
xor U3644 (N_3644,N_2820,N_2619);
or U3645 (N_3645,N_2508,N_2676);
nor U3646 (N_3646,N_2581,N_2871);
nand U3647 (N_3647,N_2541,N_1568);
or U3648 (N_3648,N_2937,N_2947);
and U3649 (N_3649,N_1659,N_1577);
nor U3650 (N_3650,N_2090,N_2550);
or U3651 (N_3651,N_2306,N_2807);
nand U3652 (N_3652,N_1915,N_1949);
and U3653 (N_3653,N_2587,N_1921);
nand U3654 (N_3654,N_1535,N_2515);
nand U3655 (N_3655,N_2053,N_2770);
nand U3656 (N_3656,N_2246,N_2749);
nand U3657 (N_3657,N_2370,N_2353);
and U3658 (N_3658,N_2547,N_1663);
xnor U3659 (N_3659,N_2187,N_1930);
and U3660 (N_3660,N_2063,N_2783);
and U3661 (N_3661,N_2147,N_2029);
nor U3662 (N_3662,N_1960,N_2360);
nor U3663 (N_3663,N_2404,N_2565);
and U3664 (N_3664,N_1987,N_2903);
nor U3665 (N_3665,N_1599,N_2146);
nor U3666 (N_3666,N_1697,N_2916);
nand U3667 (N_3667,N_1610,N_1973);
nor U3668 (N_3668,N_2675,N_2396);
and U3669 (N_3669,N_1674,N_2743);
nor U3670 (N_3670,N_2805,N_1600);
nor U3671 (N_3671,N_2276,N_2368);
nand U3672 (N_3672,N_1543,N_2887);
nand U3673 (N_3673,N_2680,N_1906);
xor U3674 (N_3674,N_1615,N_2655);
nand U3675 (N_3675,N_2539,N_2318);
nand U3676 (N_3676,N_2856,N_2704);
and U3677 (N_3677,N_2452,N_2782);
xnor U3678 (N_3678,N_2135,N_1565);
and U3679 (N_3679,N_1876,N_2803);
nand U3680 (N_3680,N_1858,N_1514);
and U3681 (N_3681,N_2219,N_2203);
nand U3682 (N_3682,N_1955,N_1509);
and U3683 (N_3683,N_2921,N_2517);
and U3684 (N_3684,N_2223,N_1699);
and U3685 (N_3685,N_1893,N_2106);
nor U3686 (N_3686,N_2027,N_2978);
or U3687 (N_3687,N_2875,N_2104);
and U3688 (N_3688,N_2427,N_1802);
and U3689 (N_3689,N_2297,N_2083);
and U3690 (N_3690,N_1889,N_2926);
nor U3691 (N_3691,N_2348,N_2150);
nand U3692 (N_3692,N_2037,N_1531);
and U3693 (N_3693,N_1758,N_2069);
nor U3694 (N_3694,N_2232,N_2755);
or U3695 (N_3695,N_1662,N_1649);
nand U3696 (N_3696,N_1567,N_2562);
and U3697 (N_3697,N_2890,N_2576);
xor U3698 (N_3698,N_2175,N_2491);
or U3699 (N_3699,N_2412,N_1835);
nand U3700 (N_3700,N_2453,N_1569);
nand U3701 (N_3701,N_2592,N_1778);
or U3702 (N_3702,N_2860,N_2355);
nand U3703 (N_3703,N_2434,N_1574);
nand U3704 (N_3704,N_2151,N_2768);
nand U3705 (N_3705,N_1956,N_2870);
or U3706 (N_3706,N_2129,N_1936);
nand U3707 (N_3707,N_2139,N_2906);
nand U3708 (N_3708,N_2213,N_1925);
nor U3709 (N_3709,N_2503,N_2569);
and U3710 (N_3710,N_2996,N_2382);
nor U3711 (N_3711,N_1979,N_2345);
nand U3712 (N_3712,N_1704,N_1732);
and U3713 (N_3713,N_1953,N_2058);
nand U3714 (N_3714,N_1673,N_2715);
and U3715 (N_3715,N_2391,N_2635);
nor U3716 (N_3716,N_2746,N_2507);
xnor U3717 (N_3717,N_1683,N_2293);
nand U3718 (N_3718,N_2578,N_2103);
nand U3719 (N_3719,N_2331,N_1817);
or U3720 (N_3720,N_2282,N_1937);
or U3721 (N_3721,N_2504,N_2778);
and U3722 (N_3722,N_1619,N_2164);
nand U3723 (N_3723,N_1977,N_2754);
or U3724 (N_3724,N_2024,N_2904);
or U3725 (N_3725,N_2418,N_2258);
nor U3726 (N_3726,N_2471,N_1905);
nor U3727 (N_3727,N_2296,N_2851);
and U3728 (N_3728,N_2925,N_1551);
or U3729 (N_3729,N_2791,N_2126);
and U3730 (N_3730,N_1729,N_2312);
or U3731 (N_3731,N_2062,N_1840);
nand U3732 (N_3732,N_2268,N_2731);
or U3733 (N_3733,N_2497,N_2156);
or U3734 (N_3734,N_2713,N_2093);
and U3735 (N_3735,N_2977,N_1818);
and U3736 (N_3736,N_1838,N_1634);
xnor U3737 (N_3737,N_2155,N_1962);
nor U3738 (N_3738,N_2220,N_1800);
nand U3739 (N_3739,N_2237,N_1902);
and U3740 (N_3740,N_2866,N_2767);
nand U3741 (N_3741,N_2082,N_1546);
or U3742 (N_3742,N_2489,N_2634);
or U3743 (N_3743,N_2646,N_1801);
nand U3744 (N_3744,N_1828,N_2131);
and U3745 (N_3745,N_2339,N_2443);
or U3746 (N_3746,N_2590,N_2163);
nand U3747 (N_3747,N_2840,N_2614);
and U3748 (N_3748,N_2235,N_2442);
and U3749 (N_3749,N_2091,N_2841);
and U3750 (N_3750,N_2158,N_2616);
nand U3751 (N_3751,N_2909,N_2191);
xnor U3752 (N_3752,N_2257,N_2360);
or U3753 (N_3753,N_1946,N_2920);
and U3754 (N_3754,N_1584,N_2196);
nor U3755 (N_3755,N_2517,N_1550);
nor U3756 (N_3756,N_2704,N_2435);
nor U3757 (N_3757,N_2975,N_2924);
or U3758 (N_3758,N_1590,N_2344);
nor U3759 (N_3759,N_2343,N_2789);
and U3760 (N_3760,N_2919,N_1596);
nand U3761 (N_3761,N_2767,N_1685);
nor U3762 (N_3762,N_2290,N_2975);
nor U3763 (N_3763,N_2200,N_1524);
nand U3764 (N_3764,N_2316,N_2461);
nand U3765 (N_3765,N_1554,N_2302);
nor U3766 (N_3766,N_2460,N_1525);
xnor U3767 (N_3767,N_1846,N_2724);
and U3768 (N_3768,N_2768,N_2033);
xor U3769 (N_3769,N_2629,N_2435);
nor U3770 (N_3770,N_2706,N_2124);
nor U3771 (N_3771,N_1651,N_1702);
nor U3772 (N_3772,N_2794,N_1929);
nor U3773 (N_3773,N_2716,N_2578);
nand U3774 (N_3774,N_1922,N_2762);
or U3775 (N_3775,N_2743,N_2804);
nor U3776 (N_3776,N_2941,N_2196);
or U3777 (N_3777,N_2533,N_1740);
nor U3778 (N_3778,N_2664,N_1568);
nand U3779 (N_3779,N_2897,N_2326);
and U3780 (N_3780,N_2824,N_2294);
or U3781 (N_3781,N_1987,N_1996);
xnor U3782 (N_3782,N_2754,N_2156);
nor U3783 (N_3783,N_2415,N_2190);
xnor U3784 (N_3784,N_1829,N_2078);
or U3785 (N_3785,N_1505,N_2824);
or U3786 (N_3786,N_1808,N_2914);
nand U3787 (N_3787,N_2536,N_2755);
nand U3788 (N_3788,N_2728,N_1868);
nor U3789 (N_3789,N_2147,N_2152);
nand U3790 (N_3790,N_2989,N_2999);
nor U3791 (N_3791,N_2720,N_2032);
and U3792 (N_3792,N_2500,N_1960);
or U3793 (N_3793,N_2711,N_1624);
or U3794 (N_3794,N_2240,N_2645);
or U3795 (N_3795,N_2100,N_2944);
nand U3796 (N_3796,N_2158,N_2718);
and U3797 (N_3797,N_2647,N_1732);
and U3798 (N_3798,N_2780,N_1557);
nor U3799 (N_3799,N_1765,N_2596);
nand U3800 (N_3800,N_1576,N_1512);
nand U3801 (N_3801,N_2832,N_2028);
nand U3802 (N_3802,N_1656,N_1529);
nand U3803 (N_3803,N_1652,N_2299);
or U3804 (N_3804,N_2549,N_1776);
nor U3805 (N_3805,N_2985,N_1945);
or U3806 (N_3806,N_2749,N_2819);
and U3807 (N_3807,N_2677,N_2347);
nand U3808 (N_3808,N_2010,N_2239);
nor U3809 (N_3809,N_2284,N_1868);
nor U3810 (N_3810,N_1946,N_2384);
and U3811 (N_3811,N_2193,N_2133);
xor U3812 (N_3812,N_1716,N_2638);
nand U3813 (N_3813,N_1820,N_2567);
nand U3814 (N_3814,N_2283,N_1933);
and U3815 (N_3815,N_1528,N_2665);
or U3816 (N_3816,N_2792,N_2898);
nand U3817 (N_3817,N_1838,N_2793);
and U3818 (N_3818,N_2718,N_2824);
and U3819 (N_3819,N_1641,N_2185);
or U3820 (N_3820,N_1971,N_2393);
and U3821 (N_3821,N_2650,N_2941);
and U3822 (N_3822,N_2516,N_1564);
nor U3823 (N_3823,N_2859,N_2876);
nor U3824 (N_3824,N_2054,N_2833);
nor U3825 (N_3825,N_1953,N_2255);
and U3826 (N_3826,N_2735,N_2707);
nor U3827 (N_3827,N_2193,N_1832);
and U3828 (N_3828,N_2386,N_2669);
nor U3829 (N_3829,N_2289,N_2437);
nor U3830 (N_3830,N_2430,N_2063);
or U3831 (N_3831,N_2669,N_2717);
nor U3832 (N_3832,N_2165,N_2442);
or U3833 (N_3833,N_1624,N_2952);
and U3834 (N_3834,N_1838,N_2693);
xor U3835 (N_3835,N_2099,N_2396);
nand U3836 (N_3836,N_2161,N_2450);
nor U3837 (N_3837,N_2086,N_2119);
nor U3838 (N_3838,N_1742,N_2218);
nor U3839 (N_3839,N_2618,N_2066);
nor U3840 (N_3840,N_2266,N_2069);
and U3841 (N_3841,N_2769,N_2781);
and U3842 (N_3842,N_1591,N_2483);
nand U3843 (N_3843,N_2922,N_1544);
and U3844 (N_3844,N_2070,N_2574);
and U3845 (N_3845,N_2745,N_2753);
or U3846 (N_3846,N_1987,N_2753);
xor U3847 (N_3847,N_2965,N_2958);
or U3848 (N_3848,N_2101,N_2620);
nor U3849 (N_3849,N_2838,N_2481);
xnor U3850 (N_3850,N_2657,N_2301);
and U3851 (N_3851,N_2388,N_1721);
nand U3852 (N_3852,N_2110,N_2546);
and U3853 (N_3853,N_2774,N_2022);
or U3854 (N_3854,N_2486,N_1940);
nor U3855 (N_3855,N_1892,N_2882);
nor U3856 (N_3856,N_2504,N_1513);
and U3857 (N_3857,N_2095,N_2857);
and U3858 (N_3858,N_1791,N_1681);
and U3859 (N_3859,N_2815,N_1676);
xor U3860 (N_3860,N_1653,N_1986);
nor U3861 (N_3861,N_2845,N_2890);
nand U3862 (N_3862,N_2833,N_2911);
xor U3863 (N_3863,N_2752,N_2776);
or U3864 (N_3864,N_1652,N_2787);
xor U3865 (N_3865,N_1859,N_1721);
xnor U3866 (N_3866,N_2201,N_2912);
or U3867 (N_3867,N_2059,N_1593);
xnor U3868 (N_3868,N_2504,N_2311);
nor U3869 (N_3869,N_2386,N_2605);
xor U3870 (N_3870,N_1862,N_2817);
and U3871 (N_3871,N_2833,N_1750);
nor U3872 (N_3872,N_1990,N_2708);
nor U3873 (N_3873,N_1760,N_2743);
or U3874 (N_3874,N_2820,N_2439);
xnor U3875 (N_3875,N_2124,N_2731);
xor U3876 (N_3876,N_2272,N_2505);
and U3877 (N_3877,N_2910,N_1978);
nor U3878 (N_3878,N_2851,N_1859);
nor U3879 (N_3879,N_2783,N_2221);
or U3880 (N_3880,N_2623,N_2869);
xor U3881 (N_3881,N_2251,N_2243);
nor U3882 (N_3882,N_2870,N_2966);
nor U3883 (N_3883,N_2323,N_2799);
nand U3884 (N_3884,N_2509,N_2339);
and U3885 (N_3885,N_1857,N_2931);
and U3886 (N_3886,N_2400,N_1917);
xnor U3887 (N_3887,N_2236,N_2323);
or U3888 (N_3888,N_2682,N_2803);
and U3889 (N_3889,N_2620,N_2007);
or U3890 (N_3890,N_1708,N_2021);
nand U3891 (N_3891,N_1612,N_1578);
nand U3892 (N_3892,N_2271,N_1789);
or U3893 (N_3893,N_1775,N_2832);
nand U3894 (N_3894,N_2153,N_1578);
nand U3895 (N_3895,N_2663,N_1979);
or U3896 (N_3896,N_2533,N_2121);
nand U3897 (N_3897,N_1515,N_2368);
and U3898 (N_3898,N_2367,N_1889);
or U3899 (N_3899,N_1882,N_2257);
nor U3900 (N_3900,N_2458,N_2154);
and U3901 (N_3901,N_1707,N_2169);
nor U3902 (N_3902,N_2659,N_1945);
nor U3903 (N_3903,N_1714,N_2254);
and U3904 (N_3904,N_2737,N_2153);
xor U3905 (N_3905,N_2550,N_2445);
nand U3906 (N_3906,N_2944,N_2892);
nand U3907 (N_3907,N_2331,N_2443);
nand U3908 (N_3908,N_2536,N_1697);
nor U3909 (N_3909,N_2391,N_2158);
and U3910 (N_3910,N_2876,N_2259);
xor U3911 (N_3911,N_2452,N_2275);
nor U3912 (N_3912,N_2551,N_2802);
or U3913 (N_3913,N_2629,N_2433);
nor U3914 (N_3914,N_2744,N_2522);
nand U3915 (N_3915,N_2654,N_2793);
xor U3916 (N_3916,N_2598,N_2764);
or U3917 (N_3917,N_2218,N_1666);
or U3918 (N_3918,N_1779,N_1941);
nand U3919 (N_3919,N_2791,N_1789);
and U3920 (N_3920,N_2817,N_2886);
and U3921 (N_3921,N_2461,N_2916);
nand U3922 (N_3922,N_1573,N_2071);
nor U3923 (N_3923,N_2322,N_1711);
or U3924 (N_3924,N_1642,N_2095);
nand U3925 (N_3925,N_2653,N_1846);
xor U3926 (N_3926,N_2931,N_2203);
nand U3927 (N_3927,N_2495,N_2214);
nand U3928 (N_3928,N_2006,N_2531);
or U3929 (N_3929,N_1549,N_2217);
or U3930 (N_3930,N_2634,N_1922);
or U3931 (N_3931,N_1623,N_2313);
or U3932 (N_3932,N_2173,N_2920);
or U3933 (N_3933,N_2825,N_2491);
xor U3934 (N_3934,N_1614,N_1618);
nand U3935 (N_3935,N_1504,N_2780);
and U3936 (N_3936,N_2900,N_2228);
or U3937 (N_3937,N_2943,N_1884);
or U3938 (N_3938,N_1615,N_2928);
and U3939 (N_3939,N_2036,N_1712);
and U3940 (N_3940,N_2691,N_1598);
nand U3941 (N_3941,N_1647,N_2219);
and U3942 (N_3942,N_2942,N_1808);
and U3943 (N_3943,N_2713,N_2858);
and U3944 (N_3944,N_1822,N_2654);
xnor U3945 (N_3945,N_2382,N_2125);
nand U3946 (N_3946,N_2386,N_2113);
or U3947 (N_3947,N_1933,N_2107);
nand U3948 (N_3948,N_2142,N_1970);
nor U3949 (N_3949,N_2691,N_1986);
or U3950 (N_3950,N_2594,N_1812);
and U3951 (N_3951,N_2357,N_2653);
xnor U3952 (N_3952,N_2494,N_2197);
and U3953 (N_3953,N_2903,N_2051);
nor U3954 (N_3954,N_2096,N_2210);
nor U3955 (N_3955,N_2914,N_2104);
or U3956 (N_3956,N_2227,N_2765);
nand U3957 (N_3957,N_2129,N_2974);
nor U3958 (N_3958,N_2102,N_1615);
nor U3959 (N_3959,N_1819,N_2231);
or U3960 (N_3960,N_1789,N_2794);
and U3961 (N_3961,N_2006,N_1630);
or U3962 (N_3962,N_2176,N_2762);
xnor U3963 (N_3963,N_2809,N_1812);
nand U3964 (N_3964,N_2919,N_2857);
nor U3965 (N_3965,N_1798,N_1561);
nor U3966 (N_3966,N_2924,N_2399);
nand U3967 (N_3967,N_1613,N_2653);
nor U3968 (N_3968,N_1955,N_1949);
nand U3969 (N_3969,N_1946,N_1758);
nor U3970 (N_3970,N_2671,N_2943);
or U3971 (N_3971,N_2332,N_1738);
and U3972 (N_3972,N_2938,N_1670);
and U3973 (N_3973,N_2501,N_2349);
or U3974 (N_3974,N_1849,N_1832);
xor U3975 (N_3975,N_1648,N_2711);
xor U3976 (N_3976,N_2137,N_2161);
xor U3977 (N_3977,N_2378,N_2617);
or U3978 (N_3978,N_1914,N_2899);
nor U3979 (N_3979,N_2677,N_1982);
xnor U3980 (N_3980,N_2167,N_2722);
nand U3981 (N_3981,N_1893,N_2247);
nand U3982 (N_3982,N_1858,N_2099);
nor U3983 (N_3983,N_1672,N_2753);
nor U3984 (N_3984,N_2730,N_1523);
or U3985 (N_3985,N_1684,N_2375);
xnor U3986 (N_3986,N_2331,N_1883);
or U3987 (N_3987,N_1792,N_1794);
or U3988 (N_3988,N_2073,N_2716);
nand U3989 (N_3989,N_1902,N_2177);
or U3990 (N_3990,N_1886,N_1731);
nand U3991 (N_3991,N_2562,N_1730);
or U3992 (N_3992,N_1627,N_2387);
and U3993 (N_3993,N_2844,N_2608);
or U3994 (N_3994,N_2188,N_2920);
nand U3995 (N_3995,N_2664,N_2253);
nor U3996 (N_3996,N_2747,N_2785);
nand U3997 (N_3997,N_2092,N_2121);
nor U3998 (N_3998,N_2807,N_1817);
or U3999 (N_3999,N_2087,N_2506);
and U4000 (N_4000,N_2107,N_2724);
and U4001 (N_4001,N_2690,N_1797);
or U4002 (N_4002,N_2848,N_2866);
xor U4003 (N_4003,N_1694,N_1611);
and U4004 (N_4004,N_2992,N_2683);
nand U4005 (N_4005,N_2125,N_1638);
nor U4006 (N_4006,N_1653,N_1632);
nand U4007 (N_4007,N_2527,N_2433);
nor U4008 (N_4008,N_2475,N_1924);
nand U4009 (N_4009,N_2474,N_2208);
or U4010 (N_4010,N_1791,N_2935);
nor U4011 (N_4011,N_1706,N_2954);
nor U4012 (N_4012,N_2226,N_1525);
or U4013 (N_4013,N_1671,N_2952);
and U4014 (N_4014,N_2015,N_2355);
nand U4015 (N_4015,N_1966,N_2228);
nor U4016 (N_4016,N_2654,N_2413);
and U4017 (N_4017,N_2483,N_2668);
nand U4018 (N_4018,N_2779,N_2846);
nand U4019 (N_4019,N_1739,N_1980);
nand U4020 (N_4020,N_2964,N_1771);
and U4021 (N_4021,N_2217,N_2492);
xnor U4022 (N_4022,N_2174,N_2942);
and U4023 (N_4023,N_2454,N_1893);
and U4024 (N_4024,N_2390,N_1843);
nor U4025 (N_4025,N_1855,N_1567);
and U4026 (N_4026,N_1762,N_2408);
or U4027 (N_4027,N_2072,N_2640);
nand U4028 (N_4028,N_2975,N_1969);
xor U4029 (N_4029,N_2127,N_2501);
or U4030 (N_4030,N_2808,N_1839);
nor U4031 (N_4031,N_1894,N_1653);
nor U4032 (N_4032,N_1515,N_2438);
and U4033 (N_4033,N_2242,N_2942);
and U4034 (N_4034,N_1985,N_2159);
and U4035 (N_4035,N_1560,N_2384);
nand U4036 (N_4036,N_2401,N_1959);
nor U4037 (N_4037,N_1699,N_1750);
or U4038 (N_4038,N_1850,N_2788);
and U4039 (N_4039,N_1725,N_1850);
or U4040 (N_4040,N_2326,N_2675);
and U4041 (N_4041,N_2012,N_2621);
and U4042 (N_4042,N_2349,N_1766);
xnor U4043 (N_4043,N_2421,N_1709);
nand U4044 (N_4044,N_2208,N_1844);
nor U4045 (N_4045,N_1889,N_2726);
and U4046 (N_4046,N_1737,N_1957);
nand U4047 (N_4047,N_2404,N_1758);
nand U4048 (N_4048,N_2069,N_1868);
or U4049 (N_4049,N_2789,N_1737);
nor U4050 (N_4050,N_2054,N_2294);
nand U4051 (N_4051,N_2983,N_2638);
nand U4052 (N_4052,N_2863,N_2199);
nand U4053 (N_4053,N_2616,N_2562);
or U4054 (N_4054,N_2971,N_2978);
xnor U4055 (N_4055,N_2317,N_2934);
nor U4056 (N_4056,N_1518,N_2286);
or U4057 (N_4057,N_2987,N_1811);
and U4058 (N_4058,N_2218,N_2816);
nand U4059 (N_4059,N_2882,N_1724);
nor U4060 (N_4060,N_2454,N_2730);
and U4061 (N_4061,N_1800,N_2423);
nand U4062 (N_4062,N_1697,N_1603);
and U4063 (N_4063,N_2072,N_1565);
or U4064 (N_4064,N_2224,N_2136);
and U4065 (N_4065,N_2844,N_2202);
nor U4066 (N_4066,N_2476,N_1516);
xnor U4067 (N_4067,N_2778,N_2605);
or U4068 (N_4068,N_2254,N_2664);
xnor U4069 (N_4069,N_1960,N_1594);
nand U4070 (N_4070,N_1550,N_2614);
and U4071 (N_4071,N_2410,N_2639);
or U4072 (N_4072,N_2573,N_2717);
and U4073 (N_4073,N_2390,N_1832);
or U4074 (N_4074,N_2723,N_1557);
xor U4075 (N_4075,N_1626,N_2722);
nand U4076 (N_4076,N_2561,N_1795);
nand U4077 (N_4077,N_2257,N_2120);
xor U4078 (N_4078,N_2868,N_2535);
and U4079 (N_4079,N_2785,N_2076);
nand U4080 (N_4080,N_2482,N_2533);
or U4081 (N_4081,N_2623,N_2642);
nand U4082 (N_4082,N_2693,N_2911);
nand U4083 (N_4083,N_2741,N_2054);
and U4084 (N_4084,N_2045,N_2626);
or U4085 (N_4085,N_2691,N_2073);
and U4086 (N_4086,N_1886,N_2854);
or U4087 (N_4087,N_2250,N_1569);
nand U4088 (N_4088,N_2269,N_2442);
and U4089 (N_4089,N_1515,N_2846);
nor U4090 (N_4090,N_2225,N_2030);
nand U4091 (N_4091,N_1779,N_1618);
and U4092 (N_4092,N_2847,N_1979);
xor U4093 (N_4093,N_2093,N_1637);
or U4094 (N_4094,N_2351,N_2118);
and U4095 (N_4095,N_2952,N_1676);
or U4096 (N_4096,N_1707,N_2646);
nand U4097 (N_4097,N_2733,N_2625);
nand U4098 (N_4098,N_2087,N_2328);
and U4099 (N_4099,N_2465,N_2733);
nor U4100 (N_4100,N_1603,N_2486);
or U4101 (N_4101,N_2670,N_2235);
nand U4102 (N_4102,N_2820,N_1505);
or U4103 (N_4103,N_2077,N_2101);
and U4104 (N_4104,N_2143,N_2808);
nand U4105 (N_4105,N_2937,N_1768);
or U4106 (N_4106,N_2861,N_1694);
nor U4107 (N_4107,N_1757,N_2384);
nand U4108 (N_4108,N_2235,N_2073);
and U4109 (N_4109,N_1891,N_2687);
and U4110 (N_4110,N_2888,N_1987);
nor U4111 (N_4111,N_2781,N_2446);
nand U4112 (N_4112,N_1528,N_2875);
and U4113 (N_4113,N_2693,N_2155);
nor U4114 (N_4114,N_2258,N_2149);
or U4115 (N_4115,N_2736,N_2632);
and U4116 (N_4116,N_2174,N_2828);
and U4117 (N_4117,N_1602,N_2504);
nor U4118 (N_4118,N_2720,N_1515);
and U4119 (N_4119,N_2532,N_2648);
or U4120 (N_4120,N_2501,N_2576);
or U4121 (N_4121,N_1646,N_2634);
and U4122 (N_4122,N_1506,N_1556);
nor U4123 (N_4123,N_2965,N_1653);
and U4124 (N_4124,N_1539,N_2983);
nor U4125 (N_4125,N_2742,N_2413);
nand U4126 (N_4126,N_2549,N_2684);
nor U4127 (N_4127,N_2486,N_2153);
nand U4128 (N_4128,N_1901,N_2685);
or U4129 (N_4129,N_1628,N_2952);
or U4130 (N_4130,N_2321,N_2166);
nand U4131 (N_4131,N_2688,N_2863);
nand U4132 (N_4132,N_2886,N_2393);
and U4133 (N_4133,N_2410,N_2792);
or U4134 (N_4134,N_2407,N_1600);
or U4135 (N_4135,N_2700,N_2042);
nor U4136 (N_4136,N_1643,N_1803);
or U4137 (N_4137,N_2598,N_2615);
or U4138 (N_4138,N_2109,N_2117);
nand U4139 (N_4139,N_2914,N_2319);
or U4140 (N_4140,N_2728,N_2648);
xnor U4141 (N_4141,N_2848,N_2898);
xnor U4142 (N_4142,N_2864,N_1938);
nand U4143 (N_4143,N_1833,N_2302);
and U4144 (N_4144,N_2237,N_1684);
nand U4145 (N_4145,N_1588,N_1835);
nand U4146 (N_4146,N_2626,N_2422);
or U4147 (N_4147,N_1561,N_2821);
or U4148 (N_4148,N_1519,N_1510);
and U4149 (N_4149,N_2977,N_1945);
and U4150 (N_4150,N_2367,N_2657);
xor U4151 (N_4151,N_1645,N_2593);
and U4152 (N_4152,N_2212,N_1727);
nand U4153 (N_4153,N_2314,N_2653);
and U4154 (N_4154,N_2389,N_2482);
or U4155 (N_4155,N_1813,N_1896);
xor U4156 (N_4156,N_2255,N_2656);
xor U4157 (N_4157,N_1561,N_1727);
and U4158 (N_4158,N_1746,N_2376);
nand U4159 (N_4159,N_2757,N_2812);
nor U4160 (N_4160,N_1697,N_1769);
and U4161 (N_4161,N_1805,N_1733);
nand U4162 (N_4162,N_2898,N_1563);
and U4163 (N_4163,N_1775,N_1792);
or U4164 (N_4164,N_2182,N_2691);
and U4165 (N_4165,N_2371,N_2982);
and U4166 (N_4166,N_1607,N_1783);
nand U4167 (N_4167,N_1895,N_2252);
or U4168 (N_4168,N_2326,N_1843);
and U4169 (N_4169,N_2502,N_2625);
nand U4170 (N_4170,N_1554,N_2053);
and U4171 (N_4171,N_2475,N_2514);
nand U4172 (N_4172,N_2067,N_1674);
xnor U4173 (N_4173,N_2157,N_1823);
nor U4174 (N_4174,N_2710,N_2293);
and U4175 (N_4175,N_2112,N_2409);
nor U4176 (N_4176,N_2873,N_1545);
nand U4177 (N_4177,N_1773,N_1931);
nor U4178 (N_4178,N_2281,N_2566);
and U4179 (N_4179,N_2199,N_1786);
nor U4180 (N_4180,N_2118,N_2373);
and U4181 (N_4181,N_1851,N_2403);
nand U4182 (N_4182,N_1754,N_2643);
nor U4183 (N_4183,N_2446,N_2673);
nand U4184 (N_4184,N_2944,N_2225);
nor U4185 (N_4185,N_2489,N_1567);
nand U4186 (N_4186,N_1512,N_2669);
and U4187 (N_4187,N_1958,N_2031);
xor U4188 (N_4188,N_2238,N_2289);
nor U4189 (N_4189,N_2040,N_2393);
or U4190 (N_4190,N_2929,N_2009);
or U4191 (N_4191,N_2865,N_2876);
and U4192 (N_4192,N_1816,N_2508);
nand U4193 (N_4193,N_2925,N_1801);
nand U4194 (N_4194,N_2519,N_1839);
nand U4195 (N_4195,N_2471,N_2066);
nand U4196 (N_4196,N_2298,N_2537);
xor U4197 (N_4197,N_2260,N_2809);
nor U4198 (N_4198,N_2314,N_1511);
nand U4199 (N_4199,N_2430,N_2749);
nor U4200 (N_4200,N_2645,N_1992);
and U4201 (N_4201,N_2911,N_2818);
or U4202 (N_4202,N_2059,N_2171);
nor U4203 (N_4203,N_2601,N_1765);
or U4204 (N_4204,N_1554,N_1861);
nor U4205 (N_4205,N_2551,N_1589);
or U4206 (N_4206,N_2334,N_2309);
xnor U4207 (N_4207,N_1812,N_2669);
nand U4208 (N_4208,N_1989,N_2975);
or U4209 (N_4209,N_1744,N_1988);
or U4210 (N_4210,N_1679,N_2097);
and U4211 (N_4211,N_2273,N_2246);
nor U4212 (N_4212,N_1613,N_2436);
xor U4213 (N_4213,N_2248,N_2473);
or U4214 (N_4214,N_2072,N_2272);
nand U4215 (N_4215,N_2297,N_2312);
xnor U4216 (N_4216,N_1562,N_2366);
or U4217 (N_4217,N_2368,N_2663);
nand U4218 (N_4218,N_2102,N_2903);
xor U4219 (N_4219,N_1602,N_1510);
nor U4220 (N_4220,N_2599,N_2506);
nand U4221 (N_4221,N_2416,N_2139);
nand U4222 (N_4222,N_2041,N_2474);
or U4223 (N_4223,N_1870,N_1769);
nor U4224 (N_4224,N_1534,N_2294);
nand U4225 (N_4225,N_1658,N_2771);
nand U4226 (N_4226,N_1685,N_2146);
nand U4227 (N_4227,N_2462,N_1620);
nor U4228 (N_4228,N_2874,N_2735);
and U4229 (N_4229,N_2416,N_1734);
nand U4230 (N_4230,N_1743,N_2558);
and U4231 (N_4231,N_2032,N_2164);
nand U4232 (N_4232,N_1739,N_1661);
and U4233 (N_4233,N_1590,N_1694);
or U4234 (N_4234,N_1559,N_2131);
and U4235 (N_4235,N_2846,N_2491);
xnor U4236 (N_4236,N_2743,N_2369);
xor U4237 (N_4237,N_2479,N_2275);
and U4238 (N_4238,N_2577,N_1847);
nand U4239 (N_4239,N_1849,N_2890);
or U4240 (N_4240,N_2539,N_2636);
or U4241 (N_4241,N_2173,N_2566);
and U4242 (N_4242,N_2444,N_2442);
nand U4243 (N_4243,N_1894,N_2239);
nor U4244 (N_4244,N_1628,N_1651);
or U4245 (N_4245,N_1715,N_2579);
nand U4246 (N_4246,N_2069,N_2937);
and U4247 (N_4247,N_1592,N_2507);
nor U4248 (N_4248,N_2190,N_2049);
and U4249 (N_4249,N_2274,N_2361);
nand U4250 (N_4250,N_2692,N_2237);
and U4251 (N_4251,N_2337,N_1891);
nand U4252 (N_4252,N_2451,N_1782);
nand U4253 (N_4253,N_2022,N_2018);
nand U4254 (N_4254,N_2152,N_1522);
and U4255 (N_4255,N_2601,N_2005);
nor U4256 (N_4256,N_2012,N_1952);
and U4257 (N_4257,N_2395,N_2803);
or U4258 (N_4258,N_1545,N_2682);
and U4259 (N_4259,N_1645,N_1711);
nor U4260 (N_4260,N_1948,N_2662);
or U4261 (N_4261,N_1880,N_2074);
nand U4262 (N_4262,N_1704,N_1983);
and U4263 (N_4263,N_1520,N_2968);
or U4264 (N_4264,N_1842,N_1898);
and U4265 (N_4265,N_2774,N_2613);
and U4266 (N_4266,N_1984,N_1513);
and U4267 (N_4267,N_1810,N_1638);
nand U4268 (N_4268,N_2439,N_2064);
nor U4269 (N_4269,N_2435,N_2852);
and U4270 (N_4270,N_2376,N_2108);
and U4271 (N_4271,N_2462,N_2853);
and U4272 (N_4272,N_2223,N_2116);
and U4273 (N_4273,N_2161,N_2147);
nand U4274 (N_4274,N_2284,N_2242);
nand U4275 (N_4275,N_2346,N_2310);
nor U4276 (N_4276,N_1717,N_1923);
nor U4277 (N_4277,N_1505,N_1726);
or U4278 (N_4278,N_2405,N_2242);
and U4279 (N_4279,N_1703,N_2311);
nor U4280 (N_4280,N_2356,N_1594);
xor U4281 (N_4281,N_1741,N_2450);
nor U4282 (N_4282,N_2593,N_2115);
nor U4283 (N_4283,N_1720,N_2321);
or U4284 (N_4284,N_2626,N_1931);
and U4285 (N_4285,N_1863,N_2353);
nor U4286 (N_4286,N_2628,N_2164);
and U4287 (N_4287,N_2289,N_1948);
or U4288 (N_4288,N_2960,N_1820);
and U4289 (N_4289,N_1862,N_2374);
and U4290 (N_4290,N_2552,N_1653);
and U4291 (N_4291,N_1778,N_1650);
or U4292 (N_4292,N_2867,N_2095);
nand U4293 (N_4293,N_2176,N_1743);
and U4294 (N_4294,N_2567,N_2415);
xor U4295 (N_4295,N_2024,N_1712);
and U4296 (N_4296,N_1533,N_2567);
nand U4297 (N_4297,N_1613,N_2083);
nor U4298 (N_4298,N_1751,N_2854);
nand U4299 (N_4299,N_2537,N_1833);
and U4300 (N_4300,N_2484,N_2669);
nand U4301 (N_4301,N_2666,N_1793);
nor U4302 (N_4302,N_1894,N_2187);
nor U4303 (N_4303,N_2929,N_2619);
and U4304 (N_4304,N_2009,N_1876);
and U4305 (N_4305,N_2583,N_2574);
xnor U4306 (N_4306,N_1636,N_1574);
or U4307 (N_4307,N_2465,N_1639);
or U4308 (N_4308,N_2538,N_2051);
nand U4309 (N_4309,N_1922,N_1593);
and U4310 (N_4310,N_2298,N_2259);
and U4311 (N_4311,N_2729,N_1559);
nand U4312 (N_4312,N_1690,N_2296);
nand U4313 (N_4313,N_2141,N_2403);
xor U4314 (N_4314,N_2917,N_2225);
or U4315 (N_4315,N_1750,N_2003);
nand U4316 (N_4316,N_2496,N_1797);
xnor U4317 (N_4317,N_2344,N_1602);
nor U4318 (N_4318,N_2500,N_1999);
nor U4319 (N_4319,N_1821,N_2129);
or U4320 (N_4320,N_1747,N_2267);
nor U4321 (N_4321,N_2706,N_1508);
or U4322 (N_4322,N_2985,N_1831);
nand U4323 (N_4323,N_2128,N_2623);
or U4324 (N_4324,N_1806,N_2700);
nand U4325 (N_4325,N_2829,N_2333);
nor U4326 (N_4326,N_1680,N_2694);
and U4327 (N_4327,N_2030,N_1924);
nand U4328 (N_4328,N_2382,N_2635);
nand U4329 (N_4329,N_1608,N_2636);
nand U4330 (N_4330,N_2181,N_1527);
and U4331 (N_4331,N_1634,N_2726);
or U4332 (N_4332,N_1933,N_1994);
and U4333 (N_4333,N_1622,N_1739);
nor U4334 (N_4334,N_1991,N_2369);
nor U4335 (N_4335,N_1944,N_1991);
nor U4336 (N_4336,N_2252,N_1761);
nand U4337 (N_4337,N_1947,N_2170);
nand U4338 (N_4338,N_2772,N_1591);
xnor U4339 (N_4339,N_1749,N_2435);
and U4340 (N_4340,N_1871,N_2513);
nor U4341 (N_4341,N_2726,N_2227);
or U4342 (N_4342,N_2524,N_1533);
or U4343 (N_4343,N_2000,N_2031);
nand U4344 (N_4344,N_1913,N_2408);
or U4345 (N_4345,N_2003,N_1729);
nand U4346 (N_4346,N_1630,N_2895);
nor U4347 (N_4347,N_2683,N_2643);
or U4348 (N_4348,N_1909,N_2494);
and U4349 (N_4349,N_2209,N_1837);
and U4350 (N_4350,N_2231,N_2137);
and U4351 (N_4351,N_2672,N_2569);
nand U4352 (N_4352,N_2519,N_2201);
nand U4353 (N_4353,N_1670,N_1845);
and U4354 (N_4354,N_1913,N_2042);
nor U4355 (N_4355,N_2969,N_2759);
or U4356 (N_4356,N_2988,N_2660);
or U4357 (N_4357,N_2083,N_1724);
or U4358 (N_4358,N_2784,N_1961);
and U4359 (N_4359,N_2320,N_2008);
and U4360 (N_4360,N_2285,N_2207);
and U4361 (N_4361,N_2691,N_1958);
or U4362 (N_4362,N_2134,N_2990);
and U4363 (N_4363,N_2154,N_2529);
and U4364 (N_4364,N_1783,N_2720);
and U4365 (N_4365,N_2625,N_2385);
or U4366 (N_4366,N_2896,N_2287);
nor U4367 (N_4367,N_2907,N_2137);
nand U4368 (N_4368,N_2466,N_2217);
nor U4369 (N_4369,N_2064,N_2688);
or U4370 (N_4370,N_2334,N_1932);
nand U4371 (N_4371,N_2624,N_2008);
or U4372 (N_4372,N_2435,N_2166);
or U4373 (N_4373,N_2268,N_1855);
xnor U4374 (N_4374,N_2894,N_2083);
and U4375 (N_4375,N_1653,N_2583);
xnor U4376 (N_4376,N_2182,N_2594);
nand U4377 (N_4377,N_2304,N_1575);
or U4378 (N_4378,N_2311,N_1709);
xor U4379 (N_4379,N_2414,N_1694);
nand U4380 (N_4380,N_2489,N_2100);
or U4381 (N_4381,N_1870,N_1887);
nor U4382 (N_4382,N_2259,N_1540);
nand U4383 (N_4383,N_2778,N_2133);
or U4384 (N_4384,N_1981,N_2061);
nand U4385 (N_4385,N_2293,N_1909);
nand U4386 (N_4386,N_2657,N_1820);
and U4387 (N_4387,N_2218,N_2667);
and U4388 (N_4388,N_1671,N_2729);
and U4389 (N_4389,N_1948,N_2480);
and U4390 (N_4390,N_1625,N_1641);
or U4391 (N_4391,N_2062,N_2353);
and U4392 (N_4392,N_1504,N_1760);
nand U4393 (N_4393,N_2699,N_1534);
nand U4394 (N_4394,N_2693,N_1725);
nor U4395 (N_4395,N_2142,N_2288);
nor U4396 (N_4396,N_2185,N_2828);
or U4397 (N_4397,N_1703,N_1763);
nor U4398 (N_4398,N_2821,N_1524);
nor U4399 (N_4399,N_2326,N_1855);
or U4400 (N_4400,N_2491,N_2632);
nor U4401 (N_4401,N_2602,N_1619);
or U4402 (N_4402,N_1852,N_2872);
nor U4403 (N_4403,N_2512,N_1725);
nor U4404 (N_4404,N_1996,N_2300);
nand U4405 (N_4405,N_1501,N_2614);
nor U4406 (N_4406,N_1606,N_2782);
and U4407 (N_4407,N_2673,N_2587);
nor U4408 (N_4408,N_2766,N_2290);
xor U4409 (N_4409,N_1854,N_2164);
or U4410 (N_4410,N_2570,N_1888);
and U4411 (N_4411,N_2112,N_2854);
or U4412 (N_4412,N_2805,N_2412);
and U4413 (N_4413,N_2347,N_2033);
and U4414 (N_4414,N_2359,N_2460);
and U4415 (N_4415,N_1981,N_2380);
and U4416 (N_4416,N_2862,N_1517);
and U4417 (N_4417,N_1826,N_2426);
nor U4418 (N_4418,N_2369,N_2715);
nand U4419 (N_4419,N_2111,N_2535);
and U4420 (N_4420,N_1831,N_1674);
or U4421 (N_4421,N_2177,N_2981);
nand U4422 (N_4422,N_1547,N_2195);
or U4423 (N_4423,N_2520,N_2545);
xor U4424 (N_4424,N_2884,N_1835);
nor U4425 (N_4425,N_2513,N_2932);
nor U4426 (N_4426,N_1781,N_2925);
and U4427 (N_4427,N_1851,N_1542);
xnor U4428 (N_4428,N_1505,N_2602);
and U4429 (N_4429,N_1542,N_2423);
or U4430 (N_4430,N_1928,N_1523);
nor U4431 (N_4431,N_2679,N_2690);
and U4432 (N_4432,N_2237,N_2705);
or U4433 (N_4433,N_2937,N_2283);
or U4434 (N_4434,N_2352,N_2188);
xnor U4435 (N_4435,N_2195,N_2614);
nand U4436 (N_4436,N_1909,N_2083);
nor U4437 (N_4437,N_2501,N_2540);
or U4438 (N_4438,N_1923,N_1682);
nand U4439 (N_4439,N_1895,N_2930);
nand U4440 (N_4440,N_2804,N_1659);
nand U4441 (N_4441,N_1846,N_2404);
or U4442 (N_4442,N_2603,N_2797);
and U4443 (N_4443,N_1982,N_2254);
or U4444 (N_4444,N_1596,N_2408);
nor U4445 (N_4445,N_2479,N_2077);
or U4446 (N_4446,N_2345,N_2682);
nor U4447 (N_4447,N_2515,N_2054);
and U4448 (N_4448,N_2668,N_2984);
and U4449 (N_4449,N_2081,N_2006);
nand U4450 (N_4450,N_2881,N_1719);
nor U4451 (N_4451,N_2968,N_2693);
or U4452 (N_4452,N_2027,N_2500);
or U4453 (N_4453,N_2716,N_2010);
nor U4454 (N_4454,N_2115,N_2932);
nand U4455 (N_4455,N_1993,N_2932);
and U4456 (N_4456,N_1694,N_2839);
nand U4457 (N_4457,N_1978,N_2384);
and U4458 (N_4458,N_2968,N_2566);
xnor U4459 (N_4459,N_2279,N_2016);
nor U4460 (N_4460,N_2390,N_2885);
or U4461 (N_4461,N_2840,N_2200);
or U4462 (N_4462,N_1871,N_2523);
nor U4463 (N_4463,N_2323,N_2775);
nor U4464 (N_4464,N_2494,N_1573);
nor U4465 (N_4465,N_2075,N_2615);
nand U4466 (N_4466,N_2767,N_2261);
nand U4467 (N_4467,N_1756,N_2759);
nor U4468 (N_4468,N_2189,N_1819);
nor U4469 (N_4469,N_2425,N_2989);
nor U4470 (N_4470,N_2936,N_1720);
nand U4471 (N_4471,N_1980,N_1675);
nor U4472 (N_4472,N_1795,N_2983);
nor U4473 (N_4473,N_2209,N_1654);
xnor U4474 (N_4474,N_2688,N_2368);
xor U4475 (N_4475,N_2602,N_2722);
xor U4476 (N_4476,N_2260,N_2052);
nand U4477 (N_4477,N_2621,N_2958);
nor U4478 (N_4478,N_2310,N_2939);
nor U4479 (N_4479,N_2762,N_2571);
nand U4480 (N_4480,N_2267,N_1610);
nor U4481 (N_4481,N_2721,N_1723);
xor U4482 (N_4482,N_1892,N_1541);
or U4483 (N_4483,N_2081,N_2014);
nor U4484 (N_4484,N_2151,N_2103);
or U4485 (N_4485,N_2963,N_1756);
or U4486 (N_4486,N_1930,N_1990);
xor U4487 (N_4487,N_2263,N_2345);
and U4488 (N_4488,N_1708,N_1751);
or U4489 (N_4489,N_1684,N_2878);
nor U4490 (N_4490,N_2612,N_1983);
and U4491 (N_4491,N_2126,N_2349);
and U4492 (N_4492,N_1915,N_2673);
xnor U4493 (N_4493,N_2085,N_1509);
nand U4494 (N_4494,N_2835,N_1615);
xnor U4495 (N_4495,N_2463,N_2372);
nand U4496 (N_4496,N_1523,N_2781);
or U4497 (N_4497,N_2736,N_2307);
or U4498 (N_4498,N_2579,N_1573);
and U4499 (N_4499,N_2516,N_1725);
xnor U4500 (N_4500,N_4272,N_4273);
and U4501 (N_4501,N_3311,N_3653);
nand U4502 (N_4502,N_3290,N_4023);
nand U4503 (N_4503,N_4177,N_4071);
nand U4504 (N_4504,N_4133,N_4097);
xor U4505 (N_4505,N_3016,N_4395);
and U4506 (N_4506,N_3272,N_3728);
nor U4507 (N_4507,N_3708,N_4078);
and U4508 (N_4508,N_3264,N_4022);
nand U4509 (N_4509,N_3136,N_3424);
or U4510 (N_4510,N_4457,N_4283);
nand U4511 (N_4511,N_3148,N_3224);
and U4512 (N_4512,N_3001,N_3748);
and U4513 (N_4513,N_3484,N_4460);
nor U4514 (N_4514,N_3785,N_3569);
and U4515 (N_4515,N_3204,N_3262);
nand U4516 (N_4516,N_3798,N_3092);
nor U4517 (N_4517,N_3236,N_3182);
and U4518 (N_4518,N_3763,N_3945);
and U4519 (N_4519,N_4226,N_3494);
and U4520 (N_4520,N_3574,N_3333);
or U4521 (N_4521,N_3385,N_3808);
or U4522 (N_4522,N_3852,N_3939);
and U4523 (N_4523,N_3379,N_3274);
and U4524 (N_4524,N_4346,N_3602);
and U4525 (N_4525,N_3742,N_3160);
and U4526 (N_4526,N_3523,N_4215);
nand U4527 (N_4527,N_3519,N_4277);
xor U4528 (N_4528,N_4330,N_3230);
nand U4529 (N_4529,N_3138,N_3587);
or U4530 (N_4530,N_4038,N_4275);
nor U4531 (N_4531,N_3793,N_3952);
or U4532 (N_4532,N_3556,N_4455);
or U4533 (N_4533,N_3943,N_3083);
or U4534 (N_4534,N_3848,N_4216);
or U4535 (N_4535,N_4483,N_4179);
nor U4536 (N_4536,N_3542,N_3752);
nor U4537 (N_4537,N_4051,N_3563);
and U4538 (N_4538,N_3759,N_3298);
nor U4539 (N_4539,N_3522,N_3816);
or U4540 (N_4540,N_3391,N_3723);
and U4541 (N_4541,N_3437,N_3051);
nand U4542 (N_4542,N_3745,N_3195);
and U4543 (N_4543,N_4012,N_4404);
nand U4544 (N_4544,N_3971,N_3303);
nand U4545 (N_4545,N_3454,N_4109);
xnor U4546 (N_4546,N_3143,N_4056);
nor U4547 (N_4547,N_4076,N_3782);
nand U4548 (N_4548,N_3972,N_4037);
nand U4549 (N_4549,N_3367,N_4142);
nand U4550 (N_4550,N_3826,N_3471);
nor U4551 (N_4551,N_4295,N_3447);
nand U4552 (N_4552,N_4421,N_3913);
and U4553 (N_4553,N_3020,N_4384);
nand U4554 (N_4554,N_3406,N_3549);
nor U4555 (N_4555,N_3661,N_3888);
and U4556 (N_4556,N_3117,N_4093);
nor U4557 (N_4557,N_4242,N_3606);
nor U4558 (N_4558,N_4351,N_3637);
nor U4559 (N_4559,N_3273,N_4017);
nor U4560 (N_4560,N_3674,N_3318);
or U4561 (N_4561,N_3356,N_3807);
and U4562 (N_4562,N_3854,N_3427);
or U4563 (N_4563,N_3104,N_3799);
or U4564 (N_4564,N_3300,N_3886);
nor U4565 (N_4565,N_4227,N_3968);
nand U4566 (N_4566,N_3255,N_4143);
or U4567 (N_4567,N_3439,N_3070);
nor U4568 (N_4568,N_4259,N_4009);
nor U4569 (N_4569,N_3038,N_4468);
and U4570 (N_4570,N_4372,N_3166);
nor U4571 (N_4571,N_3260,N_3875);
nand U4572 (N_4572,N_3977,N_3696);
nand U4573 (N_4573,N_3097,N_3192);
and U4574 (N_4574,N_4059,N_3850);
nand U4575 (N_4575,N_3281,N_4393);
or U4576 (N_4576,N_3149,N_3150);
nor U4577 (N_4577,N_3052,N_4293);
or U4578 (N_4578,N_3261,N_3455);
or U4579 (N_4579,N_3517,N_4223);
and U4580 (N_4580,N_3716,N_3414);
or U4581 (N_4581,N_4181,N_3488);
nand U4582 (N_4582,N_3256,N_3177);
and U4583 (N_4583,N_3172,N_3113);
nand U4584 (N_4584,N_3304,N_3492);
or U4585 (N_4585,N_3720,N_3937);
and U4586 (N_4586,N_4434,N_3753);
and U4587 (N_4587,N_4247,N_3105);
nand U4588 (N_4588,N_3701,N_3677);
xor U4589 (N_4589,N_3757,N_3331);
nand U4590 (N_4590,N_3110,N_3515);
nor U4591 (N_4591,N_3783,N_4328);
or U4592 (N_4592,N_3657,N_4180);
and U4593 (N_4593,N_3338,N_3328);
nor U4594 (N_4594,N_3532,N_3432);
nand U4595 (N_4595,N_3299,N_4386);
or U4596 (N_4596,N_3842,N_4001);
nand U4597 (N_4597,N_3060,N_3251);
or U4598 (N_4598,N_4053,N_3171);
nor U4599 (N_4599,N_4324,N_3025);
or U4600 (N_4600,N_3654,N_4229);
nor U4601 (N_4601,N_4007,N_3246);
nor U4602 (N_4602,N_4061,N_3946);
and U4603 (N_4603,N_3124,N_3646);
nand U4604 (N_4604,N_3226,N_4199);
nor U4605 (N_4605,N_4251,N_3368);
and U4606 (N_4606,N_3837,N_3714);
nor U4607 (N_4607,N_4108,N_4044);
and U4608 (N_4608,N_3578,N_3619);
or U4609 (N_4609,N_3209,N_3374);
nand U4610 (N_4610,N_3847,N_4090);
and U4611 (N_4611,N_3451,N_4183);
and U4612 (N_4612,N_3903,N_3965);
xor U4613 (N_4613,N_3866,N_3649);
nand U4614 (N_4614,N_4452,N_4371);
xor U4615 (N_4615,N_3651,N_3295);
or U4616 (N_4616,N_3932,N_3404);
nand U4617 (N_4617,N_3790,N_3593);
and U4618 (N_4618,N_3530,N_4363);
nand U4619 (N_4619,N_4075,N_3116);
and U4620 (N_4620,N_3675,N_3539);
nor U4621 (N_4621,N_3648,N_3108);
and U4622 (N_4622,N_3553,N_3292);
or U4623 (N_4623,N_4024,N_4124);
nand U4624 (N_4624,N_3480,N_4250);
or U4625 (N_4625,N_3620,N_3729);
and U4626 (N_4626,N_4203,N_3312);
or U4627 (N_4627,N_3141,N_3803);
nor U4628 (N_4628,N_4474,N_3947);
or U4629 (N_4629,N_3313,N_4305);
nand U4630 (N_4630,N_3555,N_4381);
or U4631 (N_4631,N_3764,N_4499);
nor U4632 (N_4632,N_4067,N_3055);
or U4633 (N_4633,N_4299,N_4112);
nand U4634 (N_4634,N_4266,N_3341);
or U4635 (N_4635,N_3395,N_3078);
xnor U4636 (N_4636,N_3794,N_3878);
nand U4637 (N_4637,N_3832,N_3389);
nand U4638 (N_4638,N_3853,N_3122);
xnor U4639 (N_4639,N_3760,N_4362);
nor U4640 (N_4640,N_3652,N_3397);
nand U4641 (N_4641,N_3217,N_4463);
nand U4642 (N_4642,N_3981,N_3769);
nor U4643 (N_4643,N_3375,N_3302);
and U4644 (N_4644,N_3685,N_3678);
nand U4645 (N_4645,N_4361,N_4368);
and U4646 (N_4646,N_3585,N_4397);
or U4647 (N_4647,N_3183,N_4354);
or U4648 (N_4648,N_3372,N_3071);
or U4649 (N_4649,N_3908,N_3282);
and U4650 (N_4650,N_4274,N_3895);
and U4651 (N_4651,N_3394,N_4193);
or U4652 (N_4652,N_4118,N_3431);
or U4653 (N_4653,N_3128,N_3420);
and U4654 (N_4654,N_3373,N_3505);
nor U4655 (N_4655,N_3018,N_3980);
xor U4656 (N_4656,N_3293,N_4425);
nand U4657 (N_4657,N_4288,N_4198);
nor U4658 (N_4658,N_3450,N_3777);
nand U4659 (N_4659,N_3636,N_4125);
or U4660 (N_4660,N_3986,N_3901);
nand U4661 (N_4661,N_3681,N_3030);
and U4662 (N_4662,N_3682,N_3989);
and U4663 (N_4663,N_4427,N_4070);
nor U4664 (N_4664,N_3547,N_3087);
and U4665 (N_4665,N_3332,N_4132);
nand U4666 (N_4666,N_3604,N_3687);
nor U4667 (N_4667,N_3325,N_3448);
nor U4668 (N_4668,N_3434,N_4348);
nand U4669 (N_4669,N_3827,N_3383);
nand U4670 (N_4670,N_4413,N_4429);
xor U4671 (N_4671,N_3558,N_3573);
and U4672 (N_4672,N_4207,N_4428);
and U4673 (N_4673,N_4159,N_3275);
and U4674 (N_4674,N_3684,N_4082);
nand U4675 (N_4675,N_3041,N_3934);
xor U4676 (N_4676,N_4016,N_4212);
or U4677 (N_4677,N_3710,N_4206);
nand U4678 (N_4678,N_3403,N_4360);
xnor U4679 (N_4679,N_3914,N_3964);
or U4680 (N_4680,N_3796,N_3643);
nor U4681 (N_4681,N_3543,N_4326);
and U4682 (N_4682,N_4334,N_3017);
nor U4683 (N_4683,N_4400,N_4015);
or U4684 (N_4684,N_4020,N_4475);
xnor U4685 (N_4685,N_4158,N_3100);
nor U4686 (N_4686,N_3507,N_3398);
and U4687 (N_4687,N_4151,N_3514);
or U4688 (N_4688,N_3381,N_3916);
and U4689 (N_4689,N_4111,N_4103);
and U4690 (N_4690,N_4147,N_3887);
nor U4691 (N_4691,N_3098,N_4278);
xor U4692 (N_4692,N_3548,N_3266);
or U4693 (N_4693,N_3402,N_3039);
and U4694 (N_4694,N_3057,N_3608);
nand U4695 (N_4695,N_3533,N_3787);
nor U4696 (N_4696,N_4482,N_4052);
or U4697 (N_4697,N_3452,N_4058);
nand U4698 (N_4698,N_3059,N_3771);
or U4699 (N_4699,N_4149,N_4213);
or U4700 (N_4700,N_4034,N_3112);
nand U4701 (N_4701,N_3773,N_3546);
or U4702 (N_4702,N_3605,N_4013);
or U4703 (N_4703,N_3446,N_3344);
and U4704 (N_4704,N_4257,N_3525);
nand U4705 (N_4705,N_3711,N_3744);
or U4706 (N_4706,N_3287,N_4126);
nand U4707 (N_4707,N_3475,N_4376);
and U4708 (N_4708,N_3029,N_3072);
and U4709 (N_4709,N_4117,N_3933);
or U4710 (N_4710,N_3929,N_3000);
nand U4711 (N_4711,N_3234,N_3856);
and U4712 (N_4712,N_3921,N_3702);
or U4713 (N_4713,N_3890,N_4217);
nor U4714 (N_4714,N_3993,N_3580);
or U4715 (N_4715,N_3056,N_3865);
nand U4716 (N_4716,N_3985,N_3671);
nand U4717 (N_4717,N_3305,N_4319);
or U4718 (N_4718,N_3090,N_3504);
or U4719 (N_4719,N_3706,N_3317);
and U4720 (N_4720,N_3703,N_3963);
nor U4721 (N_4721,N_3936,N_3429);
or U4722 (N_4722,N_3241,N_4234);
and U4723 (N_4723,N_3984,N_3167);
nor U4724 (N_4724,N_3500,N_3962);
and U4725 (N_4725,N_4420,N_3902);
or U4726 (N_4726,N_4487,N_3709);
nand U4727 (N_4727,N_4336,N_3046);
nor U4728 (N_4728,N_3258,N_4191);
nor U4729 (N_4729,N_3487,N_4172);
nand U4730 (N_4730,N_3622,N_4091);
or U4731 (N_4731,N_4359,N_3225);
or U4732 (N_4732,N_4138,N_3067);
nor U4733 (N_4733,N_3874,N_3600);
nand U4734 (N_4734,N_3770,N_4446);
or U4735 (N_4735,N_3592,N_3283);
nor U4736 (N_4736,N_3238,N_4355);
or U4737 (N_4737,N_4441,N_3726);
nand U4738 (N_4738,N_3893,N_3843);
and U4739 (N_4739,N_3747,N_3307);
nand U4740 (N_4740,N_4261,N_3954);
nand U4741 (N_4741,N_3075,N_4104);
or U4742 (N_4742,N_3468,N_3322);
or U4743 (N_4743,N_3125,N_3876);
nand U4744 (N_4744,N_3179,N_4011);
nand U4745 (N_4745,N_3101,N_4380);
xnor U4746 (N_4746,N_4029,N_4205);
xnor U4747 (N_4747,N_3062,N_3526);
nand U4748 (N_4748,N_3203,N_4136);
nor U4749 (N_4749,N_3023,N_4163);
or U4750 (N_4750,N_4155,N_3491);
xnor U4751 (N_4751,N_4235,N_3221);
and U4752 (N_4752,N_3695,N_4344);
or U4753 (N_4753,N_3516,N_3970);
nor U4754 (N_4754,N_3944,N_3582);
and U4755 (N_4755,N_4315,N_3905);
nand U4756 (N_4756,N_3662,N_3310);
nand U4757 (N_4757,N_4264,N_3165);
xor U4758 (N_4758,N_3297,N_3387);
or U4759 (N_4759,N_3616,N_3650);
xnor U4760 (N_4760,N_3359,N_3880);
or U4761 (N_4761,N_4262,N_4298);
and U4762 (N_4762,N_3680,N_4043);
and U4763 (N_4763,N_3715,N_4102);
nand U4764 (N_4764,N_3570,N_3076);
and U4765 (N_4765,N_4035,N_3169);
or U4766 (N_4766,N_3428,N_3979);
nand U4767 (N_4767,N_4050,N_3214);
or U4768 (N_4768,N_4100,N_3178);
nand U4769 (N_4769,N_3694,N_3134);
and U4770 (N_4770,N_3871,N_3733);
nand U4771 (N_4771,N_3206,N_3673);
nand U4772 (N_4772,N_4208,N_3257);
nor U4773 (N_4773,N_3289,N_3967);
nand U4774 (N_4774,N_3957,N_3707);
and U4775 (N_4775,N_3629,N_3109);
nand U4776 (N_4776,N_4340,N_4160);
or U4777 (N_4777,N_3002,N_4409);
xnor U4778 (N_4778,N_3705,N_4174);
nand U4779 (N_4779,N_3909,N_3614);
xnor U4780 (N_4780,N_4454,N_4048);
and U4781 (N_4781,N_3973,N_3974);
or U4782 (N_4782,N_4440,N_3354);
or U4783 (N_4783,N_3800,N_3811);
and U4784 (N_4784,N_3478,N_4122);
nand U4785 (N_4785,N_4169,N_3380);
nor U4786 (N_4786,N_3786,N_4347);
or U4787 (N_4787,N_3915,N_4327);
or U4788 (N_4788,N_3249,N_3676);
nand U4789 (N_4789,N_4239,N_4433);
or U4790 (N_4790,N_3482,N_3425);
xor U4791 (N_4791,N_3315,N_3340);
nand U4792 (N_4792,N_3635,N_4436);
nor U4793 (N_4793,N_3123,N_3743);
nor U4794 (N_4794,N_3316,N_3469);
nor U4795 (N_4795,N_3551,N_3640);
nand U4796 (N_4796,N_3513,N_3013);
xnor U4797 (N_4797,N_4105,N_3035);
or U4798 (N_4798,N_3527,N_3554);
or U4799 (N_4799,N_3598,N_3806);
and U4800 (N_4800,N_3584,N_3645);
and U4801 (N_4801,N_3173,N_4088);
nand U4802 (N_4802,N_4481,N_4335);
nor U4803 (N_4803,N_3308,N_4025);
nor U4804 (N_4804,N_3334,N_4453);
nor U4805 (N_4805,N_3269,N_3863);
and U4806 (N_4806,N_3867,N_4042);
nor U4807 (N_4807,N_4403,N_3704);
nand U4808 (N_4808,N_3529,N_3762);
nor U4809 (N_4809,N_3781,N_4290);
and U4810 (N_4810,N_3831,N_4480);
and U4811 (N_4811,N_3008,N_4431);
or U4812 (N_4812,N_3725,N_3336);
or U4813 (N_4813,N_4284,N_3919);
nor U4814 (N_4814,N_3474,N_3641);
and U4815 (N_4815,N_4443,N_3268);
nor U4816 (N_4816,N_3626,N_4130);
nand U4817 (N_4817,N_3463,N_3926);
or U4818 (N_4818,N_3858,N_3363);
or U4819 (N_4819,N_4026,N_4406);
nand U4820 (N_4820,N_4137,N_3817);
or U4821 (N_4821,N_3021,N_3756);
nor U4822 (N_4822,N_3692,N_3667);
nor U4823 (N_4823,N_3288,N_3278);
or U4824 (N_4824,N_3309,N_4300);
or U4825 (N_4825,N_4402,N_4072);
nor U4826 (N_4826,N_4218,N_4003);
and U4827 (N_4827,N_3479,N_4369);
and U4828 (N_4828,N_3889,N_4085);
and U4829 (N_4829,N_4031,N_3982);
nand U4830 (N_4830,N_3294,N_3423);
nand U4831 (N_4831,N_3459,N_3306);
nor U4832 (N_4832,N_3955,N_3462);
and U4833 (N_4833,N_3106,N_3658);
nor U4834 (N_4834,N_3417,N_3618);
xnor U4835 (N_4835,N_3821,N_4129);
and U4836 (N_4836,N_4260,N_3263);
xnor U4837 (N_4837,N_3855,N_3412);
and U4838 (N_4838,N_4069,N_3460);
nor U4839 (N_4839,N_3839,N_4349);
nor U4840 (N_4840,N_3885,N_3066);
and U4841 (N_4841,N_3207,N_3024);
nand U4842 (N_4842,N_3058,N_4279);
xnor U4843 (N_4843,N_4370,N_4128);
nand U4844 (N_4844,N_4080,N_3642);
and U4845 (N_4845,N_3321,N_3201);
nor U4846 (N_4846,N_3577,N_3006);
nor U4847 (N_4847,N_4173,N_4219);
nand U4848 (N_4848,N_3992,N_4418);
or U4849 (N_4849,N_4342,N_4352);
and U4850 (N_4850,N_4150,N_3416);
xnor U4851 (N_4851,N_3976,N_4492);
or U4852 (N_4852,N_3319,N_4196);
and U4853 (N_4853,N_4435,N_3664);
nor U4854 (N_4854,N_3153,N_3765);
or U4855 (N_4855,N_4055,N_4323);
nor U4856 (N_4856,N_4225,N_3126);
or U4857 (N_4857,N_3019,N_3660);
xor U4858 (N_4858,N_3879,N_4077);
nor U4859 (N_4859,N_4379,N_3524);
or U4860 (N_4860,N_3481,N_3761);
nand U4861 (N_4861,N_4276,N_3647);
or U4862 (N_4862,N_3027,N_4398);
or U4863 (N_4863,N_3210,N_3730);
nor U4864 (N_4864,N_4365,N_3638);
or U4865 (N_4865,N_3749,N_4243);
nor U4866 (N_4866,N_4232,N_3047);
and U4867 (N_4867,N_3697,N_4407);
or U4868 (N_4868,N_4253,N_4411);
or U4869 (N_4869,N_4157,N_4116);
and U4870 (N_4870,N_4186,N_3518);
nor U4871 (N_4871,N_3998,N_3330);
and U4872 (N_4872,N_3912,N_3501);
nand U4873 (N_4873,N_3511,N_3034);
or U4874 (N_4874,N_3624,N_4139);
nand U4875 (N_4875,N_3668,N_3438);
nand U4876 (N_4876,N_3228,N_4060);
nand U4877 (N_4877,N_3588,N_3615);
nor U4878 (N_4878,N_3253,N_3994);
xnor U4879 (N_4879,N_4014,N_3346);
or U4880 (N_4880,N_3069,N_4332);
or U4881 (N_4881,N_3869,N_4282);
nor U4882 (N_4882,N_4146,N_3528);
or U4883 (N_4883,N_3343,N_3746);
nand U4884 (N_4884,N_4202,N_3736);
xnor U4885 (N_4885,N_3795,N_3894);
nor U4886 (N_4886,N_4000,N_3413);
and U4887 (N_4887,N_4459,N_3951);
xor U4888 (N_4888,N_4367,N_3457);
nand U4889 (N_4889,N_3776,N_3096);
nand U4890 (N_4890,N_3922,N_4064);
xnor U4891 (N_4891,N_3433,N_3004);
nor U4892 (N_4892,N_3734,N_4461);
nor U4893 (N_4893,N_3158,N_4491);
nand U4894 (N_4894,N_3011,N_3031);
xnor U4895 (N_4895,N_3930,N_4092);
nor U4896 (N_4896,N_3223,N_3564);
and U4897 (N_4897,N_4066,N_4466);
nor U4898 (N_4898,N_3559,N_3928);
and U4899 (N_4899,N_4417,N_4280);
and U4900 (N_4900,N_3859,N_3441);
and U4901 (N_4901,N_4063,N_3738);
and U4902 (N_4902,N_3613,N_3983);
nor U4903 (N_4903,N_4165,N_3227);
nand U4904 (N_4904,N_4045,N_4479);
or U4905 (N_4905,N_4170,N_3222);
or U4906 (N_4906,N_3162,N_3579);
and U4907 (N_4907,N_4374,N_3335);
nor U4908 (N_4908,N_3426,N_3621);
nor U4909 (N_4909,N_3857,N_4099);
nor U4910 (N_4910,N_3483,N_4438);
or U4911 (N_4911,N_4473,N_3846);
and U4912 (N_4912,N_4033,N_3314);
nor U4913 (N_4913,N_3639,N_3844);
nand U4914 (N_4914,N_3566,N_3891);
nand U4915 (N_4915,N_4345,N_3155);
nor U4916 (N_4916,N_4465,N_3499);
or U4917 (N_4917,N_4079,N_3093);
or U4918 (N_4918,N_3400,N_3672);
nor U4919 (N_4919,N_4490,N_4008);
nor U4920 (N_4920,N_4030,N_3683);
nor U4921 (N_4921,N_3610,N_3044);
or U4922 (N_4922,N_3157,N_3139);
or U4923 (N_4923,N_4110,N_3498);
nor U4924 (N_4924,N_4176,N_4236);
xor U4925 (N_4925,N_3541,N_3243);
nor U4926 (N_4926,N_3823,N_4311);
nand U4927 (N_4927,N_3927,N_4375);
or U4928 (N_4928,N_3472,N_4113);
nor U4929 (N_4929,N_3737,N_3247);
or U4930 (N_4930,N_3812,N_4422);
xnor U4931 (N_4931,N_3323,N_4287);
or U4932 (N_4932,N_3828,N_3599);
nand U4933 (N_4933,N_3731,N_3280);
and U4934 (N_4934,N_3917,N_3655);
nor U4935 (N_4935,N_4047,N_3495);
xor U4936 (N_4936,N_4152,N_3037);
and U4937 (N_4937,N_4382,N_3819);
nand U4938 (N_4938,N_3248,N_4306);
nand U4939 (N_4939,N_3301,N_3252);
and U4940 (N_4940,N_3216,N_4096);
nand U4941 (N_4941,N_4220,N_4333);
or U4942 (N_4942,N_3497,N_3825);
xor U4943 (N_4943,N_3200,N_3213);
nor U4944 (N_4944,N_4145,N_3767);
nor U4945 (N_4945,N_3665,N_3012);
and U4946 (N_4946,N_4387,N_4241);
and U4947 (N_4947,N_4094,N_3630);
xor U4948 (N_4948,N_3371,N_3538);
nor U4949 (N_4949,N_3085,N_3899);
and U4950 (N_4950,N_3277,N_3187);
and U4951 (N_4951,N_3208,N_4123);
nor U4952 (N_4952,N_4210,N_3445);
and U4953 (N_4953,N_4144,N_3634);
nor U4954 (N_4954,N_4357,N_4494);
or U4955 (N_4955,N_4039,N_4073);
nor U4956 (N_4956,N_4401,N_3068);
nand U4957 (N_4957,N_4211,N_3014);
or U4958 (N_4958,N_3239,N_4263);
nand U4959 (N_4959,N_3244,N_3127);
and U4960 (N_4960,N_3135,N_4054);
or U4961 (N_4961,N_3199,N_3405);
nand U4962 (N_4962,N_4358,N_4303);
and U4963 (N_4963,N_4204,N_3215);
nand U4964 (N_4964,N_3833,N_3789);
and U4965 (N_4965,N_3061,N_4390);
nand U4966 (N_4966,N_3991,N_3232);
or U4967 (N_4967,N_4294,N_4098);
and U4968 (N_4968,N_3073,N_4343);
or U4969 (N_4969,N_3851,N_3911);
or U4970 (N_4970,N_3237,N_4254);
and U4971 (N_4971,N_3140,N_4495);
and U4972 (N_4972,N_4320,N_3152);
nand U4973 (N_4973,N_3419,N_4255);
nand U4974 (N_4974,N_3609,N_3146);
and U4975 (N_4975,N_3461,N_3137);
nor U4976 (N_4976,N_3033,N_3370);
xor U4977 (N_4977,N_3987,N_3797);
nand U4978 (N_4978,N_3382,N_4028);
nand U4979 (N_4979,N_3267,N_3727);
nor U4980 (N_4980,N_3102,N_3352);
nand U4981 (N_4981,N_3510,N_4231);
and U4982 (N_4982,N_4245,N_3925);
nand U4983 (N_4983,N_3360,N_3537);
or U4984 (N_4984,N_3205,N_3193);
nand U4985 (N_4985,N_3410,N_3089);
nor U4986 (N_4986,N_3809,N_4233);
or U4987 (N_4987,N_3502,N_4189);
nor U4988 (N_4988,N_3476,N_3220);
xnor U4989 (N_4989,N_3521,N_4101);
xor U4990 (N_4990,N_4339,N_4184);
and U4991 (N_4991,N_3386,N_3603);
nand U4992 (N_4992,N_3611,N_3935);
or U4993 (N_4993,N_4107,N_3408);
or U4994 (N_4994,N_4424,N_3589);
nand U4995 (N_4995,N_4366,N_3923);
or U4996 (N_4996,N_3082,N_3486);
xor U4997 (N_4997,N_3586,N_4271);
nor U4998 (N_4998,N_4307,N_3357);
nor U4999 (N_4999,N_3361,N_4214);
nor U5000 (N_5000,N_4464,N_4391);
nor U5001 (N_5001,N_3801,N_3378);
and U5002 (N_5002,N_4171,N_4415);
and U5003 (N_5003,N_3633,N_3975);
xnor U5004 (N_5004,N_4267,N_3119);
nand U5005 (N_5005,N_3594,N_3401);
or U5006 (N_5006,N_3938,N_3990);
nand U5007 (N_5007,N_3644,N_3250);
nor U5008 (N_5008,N_4086,N_3184);
nor U5009 (N_5009,N_4430,N_3722);
and U5010 (N_5010,N_3411,N_3751);
nor U5011 (N_5011,N_3063,N_4246);
or U5012 (N_5012,N_4156,N_3095);
or U5013 (N_5013,N_3918,N_3339);
or U5014 (N_5014,N_4062,N_3818);
or U5015 (N_5015,N_4310,N_4018);
nand U5016 (N_5016,N_4040,N_4197);
nand U5017 (N_5017,N_3873,N_3689);
and U5018 (N_5018,N_4444,N_4377);
nor U5019 (N_5019,N_4192,N_3596);
or U5020 (N_5020,N_3534,N_3393);
nor U5021 (N_5021,N_4471,N_3351);
nor U5022 (N_5022,N_3042,N_3154);
nand U5023 (N_5023,N_4432,N_3103);
nor U5024 (N_5024,N_3233,N_3444);
nand U5025 (N_5025,N_3270,N_3477);
nand U5026 (N_5026,N_3181,N_4353);
and U5027 (N_5027,N_4161,N_3575);
or U5028 (N_5028,N_4412,N_3822);
nand U5029 (N_5029,N_3180,N_4269);
or U5030 (N_5030,N_3191,N_3849);
and U5031 (N_5031,N_4478,N_3049);
nand U5032 (N_5032,N_4341,N_3036);
or U5033 (N_5033,N_3048,N_4410);
or U5034 (N_5034,N_3086,N_4281);
nand U5035 (N_5035,N_4312,N_4114);
and U5036 (N_5036,N_4230,N_3324);
nor U5037 (N_5037,N_4074,N_3490);
nor U5038 (N_5038,N_3485,N_3571);
nand U5039 (N_5039,N_3422,N_4489);
or U5040 (N_5040,N_3456,N_3536);
xor U5041 (N_5041,N_3007,N_3130);
nor U5042 (N_5042,N_3557,N_4394);
xor U5043 (N_5043,N_3920,N_3719);
and U5044 (N_5044,N_3870,N_3583);
nand U5045 (N_5045,N_3435,N_3161);
and U5046 (N_5046,N_4304,N_4442);
xor U5047 (N_5047,N_3326,N_4337);
and U5048 (N_5048,N_3296,N_3834);
or U5049 (N_5049,N_3835,N_3779);
nand U5050 (N_5050,N_4195,N_4238);
xnor U5051 (N_5051,N_4488,N_4081);
xor U5052 (N_5052,N_3802,N_3168);
nand U5053 (N_5053,N_3698,N_3094);
and U5054 (N_5054,N_3453,N_3118);
nor U5055 (N_5055,N_3824,N_4087);
and U5056 (N_5056,N_4285,N_4224);
xnor U5057 (N_5057,N_4244,N_3791);
or U5058 (N_5058,N_3631,N_3940);
and U5059 (N_5059,N_4496,N_3601);
or U5060 (N_5060,N_4021,N_3219);
xnor U5061 (N_5061,N_4162,N_3064);
nand U5062 (N_5062,N_3520,N_4252);
xor U5063 (N_5063,N_3960,N_3159);
xnor U5064 (N_5064,N_3107,N_3470);
xor U5065 (N_5065,N_3700,N_3996);
nand U5066 (N_5066,N_4472,N_3329);
and U5067 (N_5067,N_3953,N_3882);
and U5068 (N_5068,N_4006,N_3612);
nand U5069 (N_5069,N_4497,N_3320);
and U5070 (N_5070,N_3473,N_3390);
and U5071 (N_5071,N_3229,N_3788);
nand U5072 (N_5072,N_3544,N_4309);
or U5073 (N_5073,N_3081,N_3956);
and U5074 (N_5074,N_3132,N_3810);
or U5075 (N_5075,N_4115,N_3415);
and U5076 (N_5076,N_3545,N_4068);
and U5077 (N_5077,N_3958,N_3732);
or U5078 (N_5078,N_4256,N_3813);
and U5079 (N_5079,N_3860,N_3623);
nor U5080 (N_5080,N_3659,N_4325);
nand U5081 (N_5081,N_3778,N_3396);
or U5082 (N_5082,N_3999,N_4154);
nor U5083 (N_5083,N_4190,N_3625);
xor U5084 (N_5084,N_4485,N_3022);
and U5085 (N_5085,N_3868,N_3493);
xnor U5086 (N_5086,N_3881,N_3713);
xnor U5087 (N_5087,N_4164,N_3080);
nor U5088 (N_5088,N_3775,N_3884);
and U5089 (N_5089,N_3197,N_3276);
nand U5090 (N_5090,N_3906,N_3561);
nand U5091 (N_5091,N_4027,N_3376);
nor U5092 (N_5092,N_3348,N_3185);
nand U5093 (N_5093,N_4399,N_4317);
nand U5094 (N_5094,N_4209,N_3814);
and U5095 (N_5095,N_3366,N_3353);
or U5096 (N_5096,N_3627,N_3053);
and U5097 (N_5097,N_3688,N_4338);
and U5098 (N_5098,N_4331,N_3286);
xor U5099 (N_5099,N_4416,N_4291);
nand U5100 (N_5100,N_4356,N_3111);
or U5101 (N_5101,N_3830,N_4083);
nand U5102 (N_5102,N_3591,N_3691);
nand U5103 (N_5103,N_3496,N_3355);
or U5104 (N_5104,N_3581,N_4032);
and U5105 (N_5105,N_4002,N_3196);
or U5106 (N_5106,N_4383,N_3512);
nand U5107 (N_5107,N_4270,N_4166);
and U5108 (N_5108,N_3345,N_3190);
nor U5109 (N_5109,N_3679,N_4036);
xnor U5110 (N_5110,N_3271,N_4041);
or U5111 (N_5111,N_3898,N_4450);
nand U5112 (N_5112,N_3562,N_3079);
and U5113 (N_5113,N_3240,N_3900);
nand U5114 (N_5114,N_3467,N_3883);
nand U5115 (N_5115,N_4414,N_3443);
nor U5116 (N_5116,N_4188,N_3758);
xor U5117 (N_5117,N_4467,N_3907);
nand U5118 (N_5118,N_3669,N_4405);
nor U5119 (N_5119,N_4408,N_3506);
nand U5120 (N_5120,N_4194,N_4378);
nor U5121 (N_5121,N_3792,N_4318);
or U5122 (N_5122,N_4127,N_3568);
xnor U5123 (N_5123,N_3768,N_3699);
nor U5124 (N_5124,N_3820,N_3077);
nand U5125 (N_5125,N_4131,N_3174);
nor U5126 (N_5126,N_3724,N_3065);
nand U5127 (N_5127,N_3508,N_3032);
nor U5128 (N_5128,N_3489,N_3074);
nor U5129 (N_5129,N_3254,N_3088);
nand U5130 (N_5130,N_4141,N_4292);
xor U5131 (N_5131,N_4389,N_3176);
nand U5132 (N_5132,N_3349,N_4265);
nand U5133 (N_5133,N_4228,N_4140);
or U5134 (N_5134,N_4004,N_4248);
xnor U5135 (N_5135,N_3838,N_3961);
nand U5136 (N_5136,N_3897,N_4065);
nor U5137 (N_5137,N_4426,N_4095);
or U5138 (N_5138,N_4364,N_3449);
nor U5139 (N_5139,N_3337,N_3231);
nand U5140 (N_5140,N_3531,N_3131);
or U5141 (N_5141,N_4419,N_3156);
nand U5142 (N_5142,N_3284,N_3690);
and U5143 (N_5143,N_3509,N_3211);
nor U5144 (N_5144,N_3265,N_4178);
or U5145 (N_5145,N_3997,N_3750);
or U5146 (N_5146,N_3949,N_4135);
nor U5147 (N_5147,N_4240,N_4498);
or U5148 (N_5148,N_3347,N_4249);
nand U5149 (N_5149,N_3099,N_4134);
or U5150 (N_5150,N_3218,N_4493);
or U5151 (N_5151,N_3291,N_3567);
nor U5152 (N_5152,N_3784,N_3774);
and U5153 (N_5153,N_3804,N_3458);
nor U5154 (N_5154,N_4049,N_3418);
or U5155 (N_5155,N_3145,N_3151);
nand U5156 (N_5156,N_4106,N_3656);
or U5157 (N_5157,N_3815,N_3693);
or U5158 (N_5158,N_3632,N_3739);
xor U5159 (N_5159,N_4296,N_3590);
nor U5160 (N_5160,N_3377,N_4462);
or U5161 (N_5161,N_3840,N_3364);
nand U5162 (N_5162,N_4329,N_4289);
and U5163 (N_5163,N_3430,N_3466);
nand U5164 (N_5164,N_4451,N_4297);
nor U5165 (N_5165,N_3628,N_3503);
or U5166 (N_5166,N_3163,N_3666);
nor U5167 (N_5167,N_4477,N_3259);
nor U5168 (N_5168,N_3862,N_3362);
xor U5169 (N_5169,N_4302,N_3147);
and U5170 (N_5170,N_3966,N_3242);
nor U5171 (N_5171,N_4200,N_4392);
nand U5172 (N_5172,N_3388,N_3597);
and U5173 (N_5173,N_3861,N_3845);
nand U5174 (N_5174,N_3565,N_3931);
or U5175 (N_5175,N_3617,N_4187);
xor U5176 (N_5176,N_3959,N_3028);
xor U5177 (N_5177,N_3245,N_3358);
nor U5178 (N_5178,N_4476,N_3133);
and U5179 (N_5179,N_3988,N_3924);
or U5180 (N_5180,N_3084,N_3175);
nor U5181 (N_5181,N_3829,N_3941);
xnor U5182 (N_5182,N_4321,N_4148);
nor U5183 (N_5183,N_4010,N_3392);
and U5184 (N_5184,N_3550,N_3121);
nor U5185 (N_5185,N_3285,N_3576);
and U5186 (N_5186,N_4222,N_3686);
and U5187 (N_5187,N_4121,N_4185);
and U5188 (N_5188,N_4182,N_3772);
nor U5189 (N_5189,N_3043,N_3327);
nand U5190 (N_5190,N_4316,N_3040);
or U5191 (N_5191,N_4373,N_3995);
and U5192 (N_5192,N_4388,N_3670);
nand U5193 (N_5193,N_4286,N_3050);
xnor U5194 (N_5194,N_4301,N_4470);
and U5195 (N_5195,N_3342,N_4484);
and U5196 (N_5196,N_3164,N_3663);
or U5197 (N_5197,N_3129,N_3552);
xnor U5198 (N_5198,N_3740,N_4385);
nand U5199 (N_5199,N_3721,N_3188);
xnor U5200 (N_5200,N_3170,N_4445);
xnor U5201 (N_5201,N_3892,N_3115);
or U5202 (N_5202,N_4458,N_3754);
or U5203 (N_5203,N_3026,N_3235);
nand U5204 (N_5204,N_4313,N_3896);
nor U5205 (N_5205,N_3755,N_4449);
xor U5206 (N_5206,N_3010,N_4447);
or U5207 (N_5207,N_4448,N_3540);
nand U5208 (N_5208,N_4308,N_3780);
or U5209 (N_5209,N_3279,N_3120);
nand U5210 (N_5210,N_4314,N_3114);
nand U5211 (N_5211,N_4486,N_3950);
nand U5212 (N_5212,N_3009,N_3872);
nor U5213 (N_5213,N_3718,N_3841);
nand U5214 (N_5214,N_3054,N_3717);
or U5215 (N_5215,N_4168,N_4221);
nand U5216 (N_5216,N_4005,N_3969);
and U5217 (N_5217,N_3045,N_3198);
nor U5218 (N_5218,N_4456,N_3948);
nand U5219 (N_5219,N_3142,N_4167);
nand U5220 (N_5220,N_3442,N_3978);
or U5221 (N_5221,N_3864,N_3535);
nand U5222 (N_5222,N_3766,N_3741);
and U5223 (N_5223,N_4153,N_3399);
nand U5224 (N_5224,N_3186,N_3607);
xnor U5225 (N_5225,N_4258,N_3877);
and U5226 (N_5226,N_4120,N_4350);
nand U5227 (N_5227,N_3189,N_4439);
xnor U5228 (N_5228,N_4119,N_3560);
xnor U5229 (N_5229,N_3005,N_3910);
or U5230 (N_5230,N_3194,N_3202);
or U5231 (N_5231,N_3409,N_3440);
nand U5232 (N_5232,N_3904,N_3465);
or U5233 (N_5233,N_3407,N_4322);
or U5234 (N_5234,N_4089,N_3942);
and U5235 (N_5235,N_4469,N_3735);
xnor U5236 (N_5236,N_3369,N_4268);
nor U5237 (N_5237,N_3595,N_3836);
nand U5238 (N_5238,N_3350,N_3712);
nor U5239 (N_5239,N_4175,N_4437);
or U5240 (N_5240,N_4396,N_3436);
xor U5241 (N_5241,N_3464,N_3421);
nor U5242 (N_5242,N_4237,N_3384);
nand U5243 (N_5243,N_3091,N_3015);
or U5244 (N_5244,N_4019,N_3572);
nand U5245 (N_5245,N_4201,N_3365);
or U5246 (N_5246,N_4423,N_3144);
or U5247 (N_5247,N_3212,N_4057);
or U5248 (N_5248,N_3805,N_3003);
or U5249 (N_5249,N_4084,N_4046);
nor U5250 (N_5250,N_3881,N_3322);
nor U5251 (N_5251,N_4134,N_3076);
and U5252 (N_5252,N_3490,N_4297);
or U5253 (N_5253,N_4269,N_3203);
or U5254 (N_5254,N_4494,N_3666);
nor U5255 (N_5255,N_3474,N_3884);
nor U5256 (N_5256,N_3760,N_3553);
nor U5257 (N_5257,N_3363,N_3843);
nor U5258 (N_5258,N_3689,N_3964);
xnor U5259 (N_5259,N_4082,N_3383);
nor U5260 (N_5260,N_4456,N_4209);
nor U5261 (N_5261,N_3476,N_3693);
xnor U5262 (N_5262,N_4233,N_3175);
or U5263 (N_5263,N_3485,N_3089);
nor U5264 (N_5264,N_3025,N_4219);
nand U5265 (N_5265,N_3412,N_4040);
and U5266 (N_5266,N_4000,N_3737);
and U5267 (N_5267,N_3098,N_3264);
nand U5268 (N_5268,N_3103,N_4127);
or U5269 (N_5269,N_3733,N_3021);
nand U5270 (N_5270,N_3452,N_3588);
nor U5271 (N_5271,N_3532,N_3330);
nor U5272 (N_5272,N_3627,N_4368);
and U5273 (N_5273,N_4105,N_3791);
nor U5274 (N_5274,N_4307,N_3913);
and U5275 (N_5275,N_3197,N_4165);
and U5276 (N_5276,N_3513,N_4402);
nand U5277 (N_5277,N_4457,N_4007);
and U5278 (N_5278,N_4494,N_4148);
and U5279 (N_5279,N_3710,N_3319);
nor U5280 (N_5280,N_4269,N_3045);
and U5281 (N_5281,N_4482,N_4264);
or U5282 (N_5282,N_3446,N_3444);
nand U5283 (N_5283,N_3314,N_3402);
nor U5284 (N_5284,N_4154,N_4005);
nor U5285 (N_5285,N_3684,N_4474);
nand U5286 (N_5286,N_3060,N_3353);
nand U5287 (N_5287,N_4304,N_4140);
and U5288 (N_5288,N_4465,N_4083);
nor U5289 (N_5289,N_3666,N_3994);
and U5290 (N_5290,N_3044,N_4453);
nand U5291 (N_5291,N_3794,N_4328);
nand U5292 (N_5292,N_3659,N_3984);
xor U5293 (N_5293,N_3817,N_3652);
and U5294 (N_5294,N_3056,N_4437);
nor U5295 (N_5295,N_3628,N_3966);
nand U5296 (N_5296,N_3341,N_3805);
or U5297 (N_5297,N_3773,N_3022);
xnor U5298 (N_5298,N_4116,N_3696);
and U5299 (N_5299,N_4046,N_4025);
nor U5300 (N_5300,N_3237,N_4344);
and U5301 (N_5301,N_4357,N_3685);
and U5302 (N_5302,N_4213,N_3447);
or U5303 (N_5303,N_4014,N_4486);
and U5304 (N_5304,N_3093,N_4045);
nand U5305 (N_5305,N_4296,N_3719);
xor U5306 (N_5306,N_3265,N_4382);
nor U5307 (N_5307,N_3854,N_3790);
nor U5308 (N_5308,N_3992,N_4359);
or U5309 (N_5309,N_3368,N_3188);
nor U5310 (N_5310,N_3019,N_3005);
nand U5311 (N_5311,N_4049,N_3780);
or U5312 (N_5312,N_4203,N_3776);
nor U5313 (N_5313,N_4175,N_3659);
nand U5314 (N_5314,N_3968,N_3147);
and U5315 (N_5315,N_3667,N_3373);
nor U5316 (N_5316,N_3833,N_4375);
nor U5317 (N_5317,N_3761,N_3013);
or U5318 (N_5318,N_3948,N_3219);
and U5319 (N_5319,N_4060,N_3490);
nand U5320 (N_5320,N_3820,N_4365);
xnor U5321 (N_5321,N_3395,N_4355);
or U5322 (N_5322,N_3584,N_4043);
nand U5323 (N_5323,N_4240,N_4053);
or U5324 (N_5324,N_3686,N_3143);
and U5325 (N_5325,N_3282,N_4499);
or U5326 (N_5326,N_3698,N_4444);
or U5327 (N_5327,N_4400,N_4448);
nor U5328 (N_5328,N_3337,N_4314);
nand U5329 (N_5329,N_3576,N_3910);
or U5330 (N_5330,N_4185,N_3206);
nand U5331 (N_5331,N_4056,N_3903);
nor U5332 (N_5332,N_3915,N_3896);
and U5333 (N_5333,N_3229,N_3156);
nor U5334 (N_5334,N_4348,N_3143);
and U5335 (N_5335,N_3073,N_4488);
and U5336 (N_5336,N_3410,N_3458);
or U5337 (N_5337,N_3346,N_3601);
xnor U5338 (N_5338,N_3858,N_3287);
and U5339 (N_5339,N_3326,N_3051);
or U5340 (N_5340,N_3511,N_3590);
or U5341 (N_5341,N_3876,N_4228);
nand U5342 (N_5342,N_3596,N_3475);
nor U5343 (N_5343,N_3788,N_4003);
and U5344 (N_5344,N_4208,N_4467);
nor U5345 (N_5345,N_3775,N_3050);
nand U5346 (N_5346,N_3336,N_3378);
or U5347 (N_5347,N_4157,N_3281);
nor U5348 (N_5348,N_3635,N_3702);
or U5349 (N_5349,N_4337,N_3085);
nand U5350 (N_5350,N_4286,N_3963);
or U5351 (N_5351,N_4251,N_3924);
or U5352 (N_5352,N_3563,N_4418);
and U5353 (N_5353,N_3888,N_3289);
or U5354 (N_5354,N_3794,N_3900);
or U5355 (N_5355,N_4015,N_4231);
xnor U5356 (N_5356,N_4321,N_4391);
nor U5357 (N_5357,N_3434,N_4055);
nand U5358 (N_5358,N_4496,N_4107);
nor U5359 (N_5359,N_4424,N_3981);
and U5360 (N_5360,N_4435,N_4196);
nor U5361 (N_5361,N_3238,N_3850);
nand U5362 (N_5362,N_4031,N_3556);
or U5363 (N_5363,N_4173,N_3211);
nor U5364 (N_5364,N_4432,N_4183);
nor U5365 (N_5365,N_4120,N_3943);
or U5366 (N_5366,N_4252,N_4276);
nand U5367 (N_5367,N_4329,N_3133);
nand U5368 (N_5368,N_4461,N_4124);
or U5369 (N_5369,N_3627,N_3203);
xor U5370 (N_5370,N_3779,N_3063);
nand U5371 (N_5371,N_3764,N_4158);
nand U5372 (N_5372,N_3393,N_4312);
nand U5373 (N_5373,N_3137,N_4477);
and U5374 (N_5374,N_3551,N_3451);
xnor U5375 (N_5375,N_3856,N_4344);
or U5376 (N_5376,N_4309,N_3697);
xnor U5377 (N_5377,N_3258,N_4044);
and U5378 (N_5378,N_3071,N_3250);
and U5379 (N_5379,N_3658,N_3433);
and U5380 (N_5380,N_3169,N_3183);
nor U5381 (N_5381,N_3558,N_4034);
nor U5382 (N_5382,N_3326,N_3327);
or U5383 (N_5383,N_4299,N_4073);
and U5384 (N_5384,N_3628,N_3116);
xor U5385 (N_5385,N_4333,N_4436);
nor U5386 (N_5386,N_3017,N_4301);
nor U5387 (N_5387,N_4057,N_4107);
nand U5388 (N_5388,N_3634,N_3251);
or U5389 (N_5389,N_3802,N_3061);
or U5390 (N_5390,N_3504,N_4483);
nand U5391 (N_5391,N_3059,N_4418);
nor U5392 (N_5392,N_3882,N_3912);
and U5393 (N_5393,N_4457,N_3665);
and U5394 (N_5394,N_3512,N_3706);
nor U5395 (N_5395,N_3019,N_4239);
and U5396 (N_5396,N_4462,N_3856);
nor U5397 (N_5397,N_3032,N_4068);
nand U5398 (N_5398,N_4325,N_3999);
or U5399 (N_5399,N_3641,N_3841);
and U5400 (N_5400,N_3627,N_4479);
or U5401 (N_5401,N_3562,N_4245);
or U5402 (N_5402,N_3112,N_3683);
xnor U5403 (N_5403,N_3311,N_4284);
or U5404 (N_5404,N_3615,N_3000);
or U5405 (N_5405,N_4388,N_4035);
nand U5406 (N_5406,N_4291,N_3180);
nand U5407 (N_5407,N_4249,N_3060);
nand U5408 (N_5408,N_4361,N_3094);
and U5409 (N_5409,N_3258,N_3713);
nor U5410 (N_5410,N_3952,N_3889);
and U5411 (N_5411,N_3578,N_3841);
nor U5412 (N_5412,N_3763,N_3518);
xor U5413 (N_5413,N_3000,N_4310);
and U5414 (N_5414,N_3176,N_3497);
and U5415 (N_5415,N_3249,N_3157);
nor U5416 (N_5416,N_4420,N_3279);
or U5417 (N_5417,N_3865,N_4090);
nand U5418 (N_5418,N_3134,N_3747);
or U5419 (N_5419,N_4192,N_4203);
xor U5420 (N_5420,N_3142,N_3376);
and U5421 (N_5421,N_3756,N_3555);
nor U5422 (N_5422,N_3040,N_3947);
nor U5423 (N_5423,N_3025,N_4365);
nor U5424 (N_5424,N_4432,N_4171);
xor U5425 (N_5425,N_4395,N_3982);
nor U5426 (N_5426,N_3590,N_4151);
nor U5427 (N_5427,N_3823,N_4279);
and U5428 (N_5428,N_3990,N_4210);
or U5429 (N_5429,N_4007,N_3301);
nand U5430 (N_5430,N_3783,N_4148);
nor U5431 (N_5431,N_3415,N_3251);
nor U5432 (N_5432,N_3245,N_3808);
and U5433 (N_5433,N_3037,N_4131);
and U5434 (N_5434,N_4347,N_3478);
and U5435 (N_5435,N_3085,N_4212);
nor U5436 (N_5436,N_3885,N_3926);
nand U5437 (N_5437,N_4093,N_4281);
nand U5438 (N_5438,N_4219,N_3508);
xnor U5439 (N_5439,N_3120,N_3655);
or U5440 (N_5440,N_4035,N_4392);
or U5441 (N_5441,N_4283,N_4291);
nand U5442 (N_5442,N_3395,N_3975);
nand U5443 (N_5443,N_3357,N_3085);
nand U5444 (N_5444,N_3106,N_4080);
and U5445 (N_5445,N_4094,N_4286);
nand U5446 (N_5446,N_3082,N_4447);
and U5447 (N_5447,N_4381,N_3056);
nor U5448 (N_5448,N_3299,N_3717);
nor U5449 (N_5449,N_4078,N_3242);
or U5450 (N_5450,N_3887,N_3209);
nand U5451 (N_5451,N_3838,N_3754);
and U5452 (N_5452,N_3815,N_3618);
or U5453 (N_5453,N_3891,N_3586);
and U5454 (N_5454,N_3501,N_4444);
nand U5455 (N_5455,N_3788,N_3495);
and U5456 (N_5456,N_3671,N_4180);
nand U5457 (N_5457,N_3029,N_3739);
nand U5458 (N_5458,N_3622,N_3212);
nand U5459 (N_5459,N_3597,N_3515);
nand U5460 (N_5460,N_4006,N_3366);
nor U5461 (N_5461,N_3576,N_3198);
xor U5462 (N_5462,N_3619,N_3309);
nand U5463 (N_5463,N_3516,N_3754);
and U5464 (N_5464,N_3737,N_3013);
xor U5465 (N_5465,N_4096,N_3269);
and U5466 (N_5466,N_3091,N_3469);
nand U5467 (N_5467,N_3454,N_4112);
or U5468 (N_5468,N_3608,N_3686);
or U5469 (N_5469,N_3789,N_3961);
xnor U5470 (N_5470,N_3637,N_3229);
nor U5471 (N_5471,N_3715,N_3674);
and U5472 (N_5472,N_3311,N_3994);
or U5473 (N_5473,N_4319,N_4187);
nand U5474 (N_5474,N_4466,N_4385);
nor U5475 (N_5475,N_4310,N_3769);
nor U5476 (N_5476,N_3324,N_3198);
and U5477 (N_5477,N_3573,N_3770);
nor U5478 (N_5478,N_3645,N_3407);
and U5479 (N_5479,N_3511,N_3354);
and U5480 (N_5480,N_3387,N_3370);
and U5481 (N_5481,N_3331,N_3871);
and U5482 (N_5482,N_3204,N_4389);
and U5483 (N_5483,N_4206,N_3292);
nor U5484 (N_5484,N_3230,N_3457);
nand U5485 (N_5485,N_4171,N_3357);
or U5486 (N_5486,N_3407,N_3014);
nand U5487 (N_5487,N_3626,N_4281);
or U5488 (N_5488,N_3677,N_3503);
or U5489 (N_5489,N_3986,N_3079);
nand U5490 (N_5490,N_3745,N_4018);
nor U5491 (N_5491,N_3448,N_3096);
or U5492 (N_5492,N_3495,N_3156);
and U5493 (N_5493,N_3192,N_3634);
nor U5494 (N_5494,N_4245,N_3389);
or U5495 (N_5495,N_4295,N_3918);
nand U5496 (N_5496,N_3040,N_3113);
xor U5497 (N_5497,N_3700,N_4337);
and U5498 (N_5498,N_3779,N_4197);
and U5499 (N_5499,N_3900,N_4164);
or U5500 (N_5500,N_3621,N_3058);
nand U5501 (N_5501,N_4413,N_3657);
and U5502 (N_5502,N_3339,N_3634);
and U5503 (N_5503,N_3333,N_3025);
nor U5504 (N_5504,N_3189,N_3758);
xor U5505 (N_5505,N_3032,N_4478);
and U5506 (N_5506,N_3444,N_4067);
nor U5507 (N_5507,N_3573,N_3819);
or U5508 (N_5508,N_4365,N_4078);
or U5509 (N_5509,N_3111,N_4215);
nor U5510 (N_5510,N_4190,N_4161);
nand U5511 (N_5511,N_4040,N_4253);
nand U5512 (N_5512,N_3920,N_3832);
nand U5513 (N_5513,N_3618,N_4148);
or U5514 (N_5514,N_3475,N_3751);
nand U5515 (N_5515,N_3540,N_4493);
nor U5516 (N_5516,N_3848,N_3709);
or U5517 (N_5517,N_3286,N_3209);
and U5518 (N_5518,N_4366,N_4027);
xnor U5519 (N_5519,N_3314,N_3155);
nand U5520 (N_5520,N_3450,N_3599);
and U5521 (N_5521,N_4050,N_4146);
and U5522 (N_5522,N_3278,N_4427);
xor U5523 (N_5523,N_3936,N_3407);
or U5524 (N_5524,N_3292,N_4086);
or U5525 (N_5525,N_3080,N_3287);
and U5526 (N_5526,N_3278,N_3368);
and U5527 (N_5527,N_4067,N_3209);
nand U5528 (N_5528,N_4064,N_3779);
xor U5529 (N_5529,N_3901,N_3302);
xor U5530 (N_5530,N_4494,N_3123);
or U5531 (N_5531,N_3430,N_4364);
xnor U5532 (N_5532,N_3756,N_4387);
nor U5533 (N_5533,N_4053,N_3628);
or U5534 (N_5534,N_3915,N_4172);
nor U5535 (N_5535,N_3202,N_4113);
or U5536 (N_5536,N_4277,N_3300);
nand U5537 (N_5537,N_4076,N_4156);
nand U5538 (N_5538,N_3656,N_3619);
xnor U5539 (N_5539,N_3979,N_3440);
and U5540 (N_5540,N_3432,N_4429);
or U5541 (N_5541,N_3907,N_3470);
nand U5542 (N_5542,N_3244,N_3853);
and U5543 (N_5543,N_4362,N_3116);
or U5544 (N_5544,N_4389,N_3113);
or U5545 (N_5545,N_3827,N_3989);
nand U5546 (N_5546,N_3600,N_4440);
xnor U5547 (N_5547,N_4161,N_3775);
nand U5548 (N_5548,N_4421,N_4109);
xnor U5549 (N_5549,N_3348,N_3497);
and U5550 (N_5550,N_3639,N_3976);
and U5551 (N_5551,N_3249,N_3455);
nand U5552 (N_5552,N_3099,N_3387);
or U5553 (N_5553,N_3053,N_3034);
and U5554 (N_5554,N_3542,N_3498);
nand U5555 (N_5555,N_3153,N_4036);
and U5556 (N_5556,N_4060,N_3590);
or U5557 (N_5557,N_4287,N_4011);
nor U5558 (N_5558,N_3728,N_4234);
xnor U5559 (N_5559,N_3377,N_3837);
and U5560 (N_5560,N_3107,N_4033);
or U5561 (N_5561,N_4336,N_3527);
nor U5562 (N_5562,N_4165,N_3451);
or U5563 (N_5563,N_4089,N_3705);
xor U5564 (N_5564,N_4430,N_3688);
nand U5565 (N_5565,N_4490,N_3962);
xnor U5566 (N_5566,N_4114,N_3721);
or U5567 (N_5567,N_4147,N_4266);
and U5568 (N_5568,N_4183,N_3099);
or U5569 (N_5569,N_3853,N_3001);
nor U5570 (N_5570,N_3460,N_3406);
nor U5571 (N_5571,N_3190,N_4160);
or U5572 (N_5572,N_3751,N_3333);
or U5573 (N_5573,N_3483,N_3745);
nand U5574 (N_5574,N_3035,N_3943);
or U5575 (N_5575,N_3937,N_3638);
or U5576 (N_5576,N_4106,N_3551);
and U5577 (N_5577,N_3152,N_3226);
xor U5578 (N_5578,N_4218,N_3908);
or U5579 (N_5579,N_3799,N_3319);
nand U5580 (N_5580,N_3978,N_3719);
and U5581 (N_5581,N_4441,N_4467);
or U5582 (N_5582,N_3912,N_3578);
nor U5583 (N_5583,N_3963,N_3445);
nor U5584 (N_5584,N_3945,N_3883);
or U5585 (N_5585,N_4077,N_3975);
nor U5586 (N_5586,N_3490,N_3556);
and U5587 (N_5587,N_3447,N_3503);
nand U5588 (N_5588,N_3267,N_3141);
xor U5589 (N_5589,N_3061,N_4195);
xnor U5590 (N_5590,N_3911,N_4107);
nand U5591 (N_5591,N_3117,N_4396);
nand U5592 (N_5592,N_4408,N_3082);
nand U5593 (N_5593,N_4063,N_3499);
or U5594 (N_5594,N_4337,N_3207);
xor U5595 (N_5595,N_3480,N_3980);
or U5596 (N_5596,N_3766,N_3299);
nor U5597 (N_5597,N_3862,N_3510);
and U5598 (N_5598,N_3053,N_4183);
and U5599 (N_5599,N_4253,N_3557);
nor U5600 (N_5600,N_4173,N_4321);
nand U5601 (N_5601,N_4004,N_4195);
or U5602 (N_5602,N_3282,N_4038);
nor U5603 (N_5603,N_3839,N_3288);
or U5604 (N_5604,N_3222,N_4205);
xnor U5605 (N_5605,N_3162,N_4278);
and U5606 (N_5606,N_3029,N_3535);
nand U5607 (N_5607,N_3828,N_4491);
or U5608 (N_5608,N_3902,N_3276);
nor U5609 (N_5609,N_4263,N_4196);
nand U5610 (N_5610,N_4385,N_4361);
or U5611 (N_5611,N_3660,N_3721);
and U5612 (N_5612,N_4252,N_3085);
and U5613 (N_5613,N_3968,N_3107);
or U5614 (N_5614,N_4084,N_3201);
and U5615 (N_5615,N_3941,N_3085);
nor U5616 (N_5616,N_3690,N_3344);
and U5617 (N_5617,N_3400,N_3992);
and U5618 (N_5618,N_3681,N_4293);
and U5619 (N_5619,N_3339,N_3761);
xnor U5620 (N_5620,N_4457,N_3382);
nor U5621 (N_5621,N_3691,N_4409);
nor U5622 (N_5622,N_3248,N_3585);
nor U5623 (N_5623,N_3467,N_4117);
and U5624 (N_5624,N_4219,N_3708);
and U5625 (N_5625,N_3705,N_3370);
or U5626 (N_5626,N_4425,N_4274);
nand U5627 (N_5627,N_4425,N_4348);
nand U5628 (N_5628,N_4444,N_4055);
nor U5629 (N_5629,N_4472,N_3024);
nor U5630 (N_5630,N_3670,N_4297);
and U5631 (N_5631,N_3564,N_3533);
nor U5632 (N_5632,N_3700,N_3831);
and U5633 (N_5633,N_3386,N_3673);
and U5634 (N_5634,N_3549,N_4077);
and U5635 (N_5635,N_4247,N_4323);
nand U5636 (N_5636,N_3239,N_3444);
and U5637 (N_5637,N_4317,N_4446);
nand U5638 (N_5638,N_4122,N_3105);
and U5639 (N_5639,N_3877,N_3360);
or U5640 (N_5640,N_4047,N_4195);
and U5641 (N_5641,N_3439,N_3051);
nand U5642 (N_5642,N_3127,N_3487);
nand U5643 (N_5643,N_3119,N_4299);
nand U5644 (N_5644,N_4192,N_3202);
nor U5645 (N_5645,N_3159,N_3105);
nand U5646 (N_5646,N_3253,N_4012);
and U5647 (N_5647,N_3922,N_4259);
xor U5648 (N_5648,N_3892,N_3651);
nand U5649 (N_5649,N_4305,N_3893);
and U5650 (N_5650,N_3589,N_3707);
nor U5651 (N_5651,N_3053,N_4048);
nor U5652 (N_5652,N_4121,N_3365);
nor U5653 (N_5653,N_3033,N_3447);
nor U5654 (N_5654,N_4087,N_3068);
or U5655 (N_5655,N_4360,N_3650);
nand U5656 (N_5656,N_3794,N_4450);
nand U5657 (N_5657,N_3833,N_4449);
nor U5658 (N_5658,N_4091,N_4428);
or U5659 (N_5659,N_3372,N_3594);
or U5660 (N_5660,N_3007,N_3171);
nor U5661 (N_5661,N_3328,N_4054);
nand U5662 (N_5662,N_3053,N_3327);
nor U5663 (N_5663,N_4338,N_3642);
or U5664 (N_5664,N_4189,N_3452);
nor U5665 (N_5665,N_3927,N_4040);
nand U5666 (N_5666,N_3544,N_3587);
and U5667 (N_5667,N_4231,N_3367);
nand U5668 (N_5668,N_3510,N_4002);
or U5669 (N_5669,N_4361,N_4430);
or U5670 (N_5670,N_3752,N_4124);
nor U5671 (N_5671,N_4112,N_4453);
nor U5672 (N_5672,N_4385,N_4320);
nor U5673 (N_5673,N_4132,N_3461);
nand U5674 (N_5674,N_3589,N_4144);
and U5675 (N_5675,N_3106,N_3831);
xnor U5676 (N_5676,N_3131,N_3911);
and U5677 (N_5677,N_4068,N_3882);
and U5678 (N_5678,N_4158,N_3612);
nor U5679 (N_5679,N_3253,N_3415);
nand U5680 (N_5680,N_3777,N_3673);
nor U5681 (N_5681,N_4029,N_3036);
or U5682 (N_5682,N_3448,N_4380);
nand U5683 (N_5683,N_4295,N_4104);
or U5684 (N_5684,N_4487,N_4383);
nor U5685 (N_5685,N_3581,N_3091);
and U5686 (N_5686,N_3135,N_4041);
nor U5687 (N_5687,N_3322,N_3192);
or U5688 (N_5688,N_4311,N_3081);
nand U5689 (N_5689,N_4332,N_3777);
and U5690 (N_5690,N_4451,N_3331);
nor U5691 (N_5691,N_3141,N_3891);
xor U5692 (N_5692,N_3648,N_3389);
nor U5693 (N_5693,N_3874,N_3179);
and U5694 (N_5694,N_3411,N_3819);
xnor U5695 (N_5695,N_3922,N_3215);
and U5696 (N_5696,N_3546,N_3815);
or U5697 (N_5697,N_3150,N_4465);
and U5698 (N_5698,N_4150,N_3246);
nor U5699 (N_5699,N_3237,N_3513);
or U5700 (N_5700,N_3144,N_3550);
and U5701 (N_5701,N_3846,N_3693);
nor U5702 (N_5702,N_3745,N_3284);
nand U5703 (N_5703,N_3119,N_3061);
and U5704 (N_5704,N_4062,N_4114);
nand U5705 (N_5705,N_4373,N_4140);
nor U5706 (N_5706,N_3860,N_3640);
nor U5707 (N_5707,N_4366,N_3447);
nand U5708 (N_5708,N_3397,N_3065);
nand U5709 (N_5709,N_3123,N_3610);
nand U5710 (N_5710,N_4490,N_3759);
nand U5711 (N_5711,N_4467,N_4050);
xnor U5712 (N_5712,N_4278,N_3373);
nor U5713 (N_5713,N_4120,N_3440);
nand U5714 (N_5714,N_3903,N_3830);
nand U5715 (N_5715,N_3190,N_3975);
and U5716 (N_5716,N_3415,N_3748);
and U5717 (N_5717,N_3993,N_3247);
or U5718 (N_5718,N_4229,N_3169);
nand U5719 (N_5719,N_4419,N_3205);
or U5720 (N_5720,N_4466,N_4136);
nand U5721 (N_5721,N_3757,N_3669);
nor U5722 (N_5722,N_4162,N_3197);
xor U5723 (N_5723,N_3589,N_4153);
xor U5724 (N_5724,N_4179,N_3227);
nor U5725 (N_5725,N_3110,N_4310);
nor U5726 (N_5726,N_3686,N_4302);
nor U5727 (N_5727,N_4123,N_4232);
and U5728 (N_5728,N_3309,N_4172);
or U5729 (N_5729,N_3291,N_3469);
or U5730 (N_5730,N_4495,N_3655);
or U5731 (N_5731,N_3456,N_3814);
and U5732 (N_5732,N_3025,N_3861);
xor U5733 (N_5733,N_3178,N_4181);
nand U5734 (N_5734,N_3143,N_4253);
xnor U5735 (N_5735,N_3504,N_3601);
and U5736 (N_5736,N_3807,N_3610);
and U5737 (N_5737,N_3935,N_3530);
nand U5738 (N_5738,N_4488,N_3588);
nor U5739 (N_5739,N_3667,N_4042);
nand U5740 (N_5740,N_3542,N_3437);
nand U5741 (N_5741,N_3669,N_3506);
and U5742 (N_5742,N_3431,N_4017);
nand U5743 (N_5743,N_3647,N_4407);
xor U5744 (N_5744,N_4253,N_4098);
or U5745 (N_5745,N_4313,N_3016);
or U5746 (N_5746,N_3187,N_4213);
nor U5747 (N_5747,N_3608,N_3434);
nor U5748 (N_5748,N_4231,N_4205);
nor U5749 (N_5749,N_3942,N_3550);
nand U5750 (N_5750,N_4017,N_3176);
and U5751 (N_5751,N_3610,N_3122);
and U5752 (N_5752,N_3661,N_4371);
nand U5753 (N_5753,N_3996,N_3288);
nand U5754 (N_5754,N_4149,N_3689);
and U5755 (N_5755,N_3968,N_3738);
and U5756 (N_5756,N_3918,N_3331);
or U5757 (N_5757,N_3821,N_3510);
nor U5758 (N_5758,N_4100,N_4243);
nor U5759 (N_5759,N_3099,N_3100);
nand U5760 (N_5760,N_3991,N_4387);
xnor U5761 (N_5761,N_3110,N_3750);
and U5762 (N_5762,N_3107,N_3211);
nand U5763 (N_5763,N_4498,N_3756);
nor U5764 (N_5764,N_3886,N_3435);
or U5765 (N_5765,N_3020,N_3357);
xnor U5766 (N_5766,N_4333,N_3431);
or U5767 (N_5767,N_4370,N_4235);
nand U5768 (N_5768,N_3124,N_3992);
and U5769 (N_5769,N_3006,N_4287);
and U5770 (N_5770,N_3936,N_3658);
or U5771 (N_5771,N_3985,N_4487);
or U5772 (N_5772,N_3905,N_3688);
and U5773 (N_5773,N_3035,N_3791);
xnor U5774 (N_5774,N_3258,N_3222);
or U5775 (N_5775,N_3059,N_3412);
and U5776 (N_5776,N_3191,N_3082);
or U5777 (N_5777,N_3355,N_4493);
and U5778 (N_5778,N_3877,N_3626);
and U5779 (N_5779,N_3808,N_4405);
and U5780 (N_5780,N_4200,N_3980);
and U5781 (N_5781,N_3048,N_4240);
nand U5782 (N_5782,N_3853,N_3234);
nor U5783 (N_5783,N_3578,N_4265);
xor U5784 (N_5784,N_3618,N_4028);
nor U5785 (N_5785,N_4257,N_3557);
and U5786 (N_5786,N_3253,N_3096);
and U5787 (N_5787,N_4362,N_3674);
nand U5788 (N_5788,N_3167,N_3146);
xor U5789 (N_5789,N_4084,N_3548);
xor U5790 (N_5790,N_3221,N_3552);
nor U5791 (N_5791,N_4266,N_4227);
nand U5792 (N_5792,N_4163,N_3484);
and U5793 (N_5793,N_3353,N_3377);
nand U5794 (N_5794,N_4439,N_3422);
nand U5795 (N_5795,N_3567,N_4144);
xnor U5796 (N_5796,N_3268,N_4241);
and U5797 (N_5797,N_3770,N_3387);
or U5798 (N_5798,N_3805,N_3978);
and U5799 (N_5799,N_4258,N_3901);
nor U5800 (N_5800,N_3371,N_4298);
nor U5801 (N_5801,N_3966,N_3311);
nand U5802 (N_5802,N_4242,N_3879);
or U5803 (N_5803,N_4081,N_3259);
nand U5804 (N_5804,N_3705,N_3115);
or U5805 (N_5805,N_3063,N_4154);
nand U5806 (N_5806,N_3954,N_3071);
or U5807 (N_5807,N_3959,N_3146);
nand U5808 (N_5808,N_3241,N_3119);
or U5809 (N_5809,N_3377,N_3554);
xor U5810 (N_5810,N_3906,N_3898);
or U5811 (N_5811,N_4263,N_3567);
and U5812 (N_5812,N_4423,N_4256);
nor U5813 (N_5813,N_3418,N_3914);
and U5814 (N_5814,N_4398,N_3938);
and U5815 (N_5815,N_4126,N_3062);
xor U5816 (N_5816,N_3712,N_3819);
nand U5817 (N_5817,N_3671,N_3723);
nand U5818 (N_5818,N_3303,N_4138);
nor U5819 (N_5819,N_3959,N_3756);
nor U5820 (N_5820,N_3749,N_3274);
nor U5821 (N_5821,N_3651,N_3452);
and U5822 (N_5822,N_4178,N_3458);
nor U5823 (N_5823,N_3350,N_3229);
nand U5824 (N_5824,N_3142,N_3923);
xor U5825 (N_5825,N_3642,N_4387);
nand U5826 (N_5826,N_4010,N_3229);
nand U5827 (N_5827,N_3564,N_4420);
and U5828 (N_5828,N_4154,N_4110);
nand U5829 (N_5829,N_3050,N_3180);
nand U5830 (N_5830,N_3452,N_3015);
nand U5831 (N_5831,N_3731,N_4264);
nor U5832 (N_5832,N_3999,N_4125);
or U5833 (N_5833,N_3593,N_3199);
nor U5834 (N_5834,N_3481,N_3083);
and U5835 (N_5835,N_3424,N_3748);
nor U5836 (N_5836,N_4445,N_3054);
nor U5837 (N_5837,N_4400,N_3503);
nand U5838 (N_5838,N_3695,N_3654);
nand U5839 (N_5839,N_3817,N_3569);
nor U5840 (N_5840,N_3338,N_4155);
xor U5841 (N_5841,N_4300,N_3918);
nand U5842 (N_5842,N_4157,N_3944);
or U5843 (N_5843,N_4084,N_3561);
or U5844 (N_5844,N_3497,N_4392);
and U5845 (N_5845,N_3137,N_3498);
or U5846 (N_5846,N_4043,N_3183);
and U5847 (N_5847,N_3460,N_3009);
nor U5848 (N_5848,N_4380,N_3574);
nand U5849 (N_5849,N_4229,N_3017);
or U5850 (N_5850,N_4051,N_4447);
and U5851 (N_5851,N_4255,N_3844);
nand U5852 (N_5852,N_3060,N_4267);
or U5853 (N_5853,N_3782,N_3539);
and U5854 (N_5854,N_4250,N_3379);
nand U5855 (N_5855,N_3177,N_3616);
nor U5856 (N_5856,N_3362,N_4377);
nor U5857 (N_5857,N_4416,N_3671);
nand U5858 (N_5858,N_4192,N_4074);
and U5859 (N_5859,N_3920,N_3179);
or U5860 (N_5860,N_3519,N_4366);
and U5861 (N_5861,N_3488,N_3102);
nand U5862 (N_5862,N_3170,N_3756);
nor U5863 (N_5863,N_3909,N_3343);
or U5864 (N_5864,N_3633,N_3642);
and U5865 (N_5865,N_3918,N_4410);
nor U5866 (N_5866,N_4462,N_3485);
or U5867 (N_5867,N_3109,N_3318);
nand U5868 (N_5868,N_4254,N_4190);
nand U5869 (N_5869,N_4142,N_3346);
nor U5870 (N_5870,N_4087,N_3540);
xor U5871 (N_5871,N_3948,N_4127);
nor U5872 (N_5872,N_3442,N_3167);
nand U5873 (N_5873,N_4376,N_4126);
or U5874 (N_5874,N_3041,N_3505);
nor U5875 (N_5875,N_3873,N_4097);
or U5876 (N_5876,N_3405,N_4415);
nor U5877 (N_5877,N_4216,N_3916);
and U5878 (N_5878,N_3929,N_4379);
and U5879 (N_5879,N_3831,N_3218);
nor U5880 (N_5880,N_3832,N_4464);
or U5881 (N_5881,N_3491,N_3378);
or U5882 (N_5882,N_4347,N_3704);
nor U5883 (N_5883,N_3974,N_3882);
or U5884 (N_5884,N_3914,N_3690);
or U5885 (N_5885,N_4383,N_3269);
nor U5886 (N_5886,N_3048,N_4273);
nand U5887 (N_5887,N_3033,N_3421);
nor U5888 (N_5888,N_3000,N_4015);
nand U5889 (N_5889,N_4414,N_3660);
nor U5890 (N_5890,N_3841,N_3741);
nor U5891 (N_5891,N_3574,N_3311);
or U5892 (N_5892,N_3381,N_4327);
and U5893 (N_5893,N_3520,N_3371);
nand U5894 (N_5894,N_3553,N_4127);
or U5895 (N_5895,N_3113,N_3203);
or U5896 (N_5896,N_3112,N_3720);
xnor U5897 (N_5897,N_3239,N_4012);
nand U5898 (N_5898,N_3519,N_3476);
xnor U5899 (N_5899,N_4458,N_3902);
and U5900 (N_5900,N_3398,N_3901);
and U5901 (N_5901,N_3495,N_4178);
nand U5902 (N_5902,N_3581,N_4361);
nand U5903 (N_5903,N_4335,N_4118);
and U5904 (N_5904,N_3154,N_3802);
xor U5905 (N_5905,N_4203,N_4031);
and U5906 (N_5906,N_3344,N_3655);
or U5907 (N_5907,N_3267,N_3332);
or U5908 (N_5908,N_3564,N_4464);
xnor U5909 (N_5909,N_4186,N_4257);
or U5910 (N_5910,N_3809,N_3428);
nand U5911 (N_5911,N_3060,N_3392);
or U5912 (N_5912,N_4389,N_4303);
xor U5913 (N_5913,N_4003,N_3514);
or U5914 (N_5914,N_4043,N_4285);
xnor U5915 (N_5915,N_3885,N_3861);
nand U5916 (N_5916,N_3839,N_3802);
nand U5917 (N_5917,N_4362,N_3873);
and U5918 (N_5918,N_4243,N_4199);
nor U5919 (N_5919,N_3118,N_3029);
or U5920 (N_5920,N_3694,N_3913);
nand U5921 (N_5921,N_3071,N_3571);
or U5922 (N_5922,N_3587,N_3784);
nand U5923 (N_5923,N_3043,N_3651);
and U5924 (N_5924,N_4001,N_4382);
xnor U5925 (N_5925,N_4072,N_3706);
nand U5926 (N_5926,N_3601,N_3018);
nand U5927 (N_5927,N_4017,N_4354);
nand U5928 (N_5928,N_3665,N_3120);
xor U5929 (N_5929,N_3579,N_3336);
or U5930 (N_5930,N_3067,N_4272);
or U5931 (N_5931,N_3737,N_4406);
nor U5932 (N_5932,N_4127,N_3680);
or U5933 (N_5933,N_3221,N_3029);
or U5934 (N_5934,N_4349,N_3105);
or U5935 (N_5935,N_3998,N_3048);
nor U5936 (N_5936,N_4307,N_3852);
or U5937 (N_5937,N_3310,N_3595);
nand U5938 (N_5938,N_4339,N_4454);
and U5939 (N_5939,N_3158,N_4447);
nand U5940 (N_5940,N_3834,N_3494);
nand U5941 (N_5941,N_3479,N_3614);
or U5942 (N_5942,N_3836,N_3315);
and U5943 (N_5943,N_3640,N_3562);
nand U5944 (N_5944,N_4345,N_3221);
nand U5945 (N_5945,N_3801,N_4072);
nand U5946 (N_5946,N_4349,N_3463);
nor U5947 (N_5947,N_3092,N_4278);
or U5948 (N_5948,N_4309,N_3402);
and U5949 (N_5949,N_3403,N_4280);
nor U5950 (N_5950,N_3650,N_4441);
and U5951 (N_5951,N_3542,N_4062);
or U5952 (N_5952,N_3492,N_3155);
nor U5953 (N_5953,N_4161,N_3382);
nor U5954 (N_5954,N_4253,N_3519);
nand U5955 (N_5955,N_3356,N_4256);
or U5956 (N_5956,N_4031,N_3524);
and U5957 (N_5957,N_4064,N_4356);
nor U5958 (N_5958,N_3670,N_3517);
nor U5959 (N_5959,N_3998,N_3074);
and U5960 (N_5960,N_3282,N_3919);
or U5961 (N_5961,N_4360,N_3620);
nor U5962 (N_5962,N_3808,N_3459);
or U5963 (N_5963,N_3713,N_3855);
or U5964 (N_5964,N_3676,N_3773);
and U5965 (N_5965,N_4337,N_3453);
xnor U5966 (N_5966,N_4221,N_3840);
or U5967 (N_5967,N_4063,N_4011);
nand U5968 (N_5968,N_3694,N_3155);
or U5969 (N_5969,N_3316,N_4469);
xnor U5970 (N_5970,N_4262,N_3708);
nor U5971 (N_5971,N_4304,N_4182);
or U5972 (N_5972,N_4364,N_4157);
or U5973 (N_5973,N_4173,N_4253);
and U5974 (N_5974,N_4403,N_4084);
nand U5975 (N_5975,N_4058,N_3129);
or U5976 (N_5976,N_3393,N_3814);
or U5977 (N_5977,N_4351,N_4406);
nand U5978 (N_5978,N_3456,N_3342);
xor U5979 (N_5979,N_4080,N_3946);
or U5980 (N_5980,N_3053,N_3841);
or U5981 (N_5981,N_3383,N_3710);
nor U5982 (N_5982,N_3948,N_3376);
nor U5983 (N_5983,N_4059,N_3099);
nand U5984 (N_5984,N_4325,N_3370);
nor U5985 (N_5985,N_3778,N_3857);
and U5986 (N_5986,N_3028,N_4143);
nand U5987 (N_5987,N_3569,N_3414);
nor U5988 (N_5988,N_3969,N_3132);
or U5989 (N_5989,N_4336,N_3442);
or U5990 (N_5990,N_3465,N_3982);
xor U5991 (N_5991,N_3796,N_3215);
nor U5992 (N_5992,N_3046,N_3245);
nor U5993 (N_5993,N_4253,N_3495);
nand U5994 (N_5994,N_3038,N_3873);
nand U5995 (N_5995,N_4305,N_3193);
or U5996 (N_5996,N_3312,N_3913);
nor U5997 (N_5997,N_3878,N_3520);
and U5998 (N_5998,N_4210,N_4237);
xnor U5999 (N_5999,N_4208,N_4381);
nor U6000 (N_6000,N_4591,N_4867);
nand U6001 (N_6001,N_4948,N_5313);
nor U6002 (N_6002,N_4702,N_4806);
or U6003 (N_6003,N_5139,N_4882);
and U6004 (N_6004,N_4568,N_5672);
or U6005 (N_6005,N_5453,N_5853);
or U6006 (N_6006,N_5185,N_5641);
nor U6007 (N_6007,N_4707,N_4743);
nand U6008 (N_6008,N_4661,N_5946);
and U6009 (N_6009,N_4723,N_5892);
or U6010 (N_6010,N_5642,N_5747);
and U6011 (N_6011,N_4842,N_5310);
xor U6012 (N_6012,N_5999,N_5883);
nor U6013 (N_6013,N_5937,N_5989);
nand U6014 (N_6014,N_5228,N_5863);
nand U6015 (N_6015,N_5502,N_5318);
nor U6016 (N_6016,N_5830,N_5521);
and U6017 (N_6017,N_4925,N_5197);
and U6018 (N_6018,N_5106,N_5528);
nand U6019 (N_6019,N_5013,N_5136);
and U6020 (N_6020,N_5748,N_5257);
and U6021 (N_6021,N_4839,N_5524);
nor U6022 (N_6022,N_4998,N_4576);
or U6023 (N_6023,N_4750,N_5950);
or U6024 (N_6024,N_4895,N_5683);
nand U6025 (N_6025,N_5527,N_5994);
nand U6026 (N_6026,N_5809,N_4663);
nand U6027 (N_6027,N_4994,N_4542);
nand U6028 (N_6028,N_5295,N_4772);
nand U6029 (N_6029,N_5008,N_4567);
or U6030 (N_6030,N_5045,N_5691);
or U6031 (N_6031,N_4958,N_5601);
or U6032 (N_6032,N_5358,N_5949);
or U6033 (N_6033,N_5836,N_5915);
nand U6034 (N_6034,N_4524,N_4960);
and U6035 (N_6035,N_5783,N_4820);
or U6036 (N_6036,N_5213,N_5977);
nor U6037 (N_6037,N_4980,N_5418);
and U6038 (N_6038,N_5895,N_4582);
or U6039 (N_6039,N_5269,N_5708);
or U6040 (N_6040,N_5653,N_5099);
nor U6041 (N_6041,N_5169,N_5694);
xor U6042 (N_6042,N_5459,N_5823);
or U6043 (N_6043,N_5334,N_4504);
nor U6044 (N_6044,N_5877,N_4651);
nand U6045 (N_6045,N_5759,N_4778);
or U6046 (N_6046,N_4982,N_5623);
and U6047 (N_6047,N_5888,N_4607);
and U6048 (N_6048,N_5561,N_5542);
nor U6049 (N_6049,N_5464,N_5326);
and U6050 (N_6050,N_4846,N_5961);
xor U6051 (N_6051,N_5223,N_5535);
and U6052 (N_6052,N_5763,N_5983);
nand U6053 (N_6053,N_5161,N_4747);
or U6054 (N_6054,N_5725,N_5074);
or U6055 (N_6055,N_5309,N_4506);
xnor U6056 (N_6056,N_5323,N_4672);
or U6057 (N_6057,N_5674,N_5673);
or U6058 (N_6058,N_4503,N_4790);
or U6059 (N_6059,N_4652,N_4717);
and U6060 (N_6060,N_5934,N_5077);
and U6061 (N_6061,N_5935,N_4755);
nor U6062 (N_6062,N_5285,N_4648);
xor U6063 (N_6063,N_4650,N_5354);
and U6064 (N_6064,N_4615,N_4543);
nor U6065 (N_6065,N_5907,N_5476);
nor U6066 (N_6066,N_4619,N_4821);
or U6067 (N_6067,N_5982,N_4632);
or U6068 (N_6068,N_4602,N_5756);
nand U6069 (N_6069,N_5945,N_4997);
or U6070 (N_6070,N_4813,N_5104);
and U6071 (N_6071,N_4984,N_4890);
or U6072 (N_6072,N_5485,N_5889);
and U6073 (N_6073,N_5781,N_4612);
nor U6074 (N_6074,N_4872,N_5216);
nand U6075 (N_6075,N_5205,N_5974);
or U6076 (N_6076,N_4517,N_5014);
nand U6077 (N_6077,N_5882,N_4570);
xnor U6078 (N_6078,N_5327,N_5990);
and U6079 (N_6079,N_4978,N_5833);
xnor U6080 (N_6080,N_5308,N_4713);
nand U6081 (N_6081,N_5779,N_4934);
and U6082 (N_6082,N_5630,N_5152);
nand U6083 (N_6083,N_5339,N_5163);
or U6084 (N_6084,N_5168,N_5585);
or U6085 (N_6085,N_4848,N_5852);
nor U6086 (N_6086,N_5773,N_5143);
or U6087 (N_6087,N_5736,N_5194);
nor U6088 (N_6088,N_5238,N_4843);
nor U6089 (N_6089,N_5279,N_5525);
nand U6090 (N_6090,N_4566,N_5956);
and U6091 (N_6091,N_5622,N_5423);
and U6092 (N_6092,N_5862,N_5256);
nand U6093 (N_6093,N_5936,N_5117);
nand U6094 (N_6094,N_5968,N_5322);
and U6095 (N_6095,N_5398,N_5193);
nor U6096 (N_6096,N_5344,N_5491);
and U6097 (N_6097,N_5910,N_4871);
and U6098 (N_6098,N_4887,N_5411);
nor U6099 (N_6099,N_5407,N_5717);
xor U6100 (N_6100,N_5345,N_5178);
and U6101 (N_6101,N_5132,N_5390);
or U6102 (N_6102,N_5359,N_5890);
or U6103 (N_6103,N_4611,N_5504);
nor U6104 (N_6104,N_5245,N_5370);
and U6105 (N_6105,N_4924,N_5599);
nand U6106 (N_6106,N_5925,N_4996);
and U6107 (N_6107,N_5565,N_5383);
xor U6108 (N_6108,N_5131,N_5879);
or U6109 (N_6109,N_5733,N_4509);
nand U6110 (N_6110,N_4667,N_5053);
or U6111 (N_6111,N_4721,N_4683);
xnor U6112 (N_6112,N_4875,N_5079);
and U6113 (N_6113,N_5384,N_5287);
nand U6114 (N_6114,N_5741,N_5769);
nand U6115 (N_6115,N_4770,N_5980);
nor U6116 (N_6116,N_5813,N_5501);
nor U6117 (N_6117,N_5837,N_4622);
nand U6118 (N_6118,N_5495,N_5349);
nor U6119 (N_6119,N_5768,N_5361);
or U6120 (N_6120,N_5162,N_5849);
nand U6121 (N_6121,N_5801,N_4768);
or U6122 (N_6122,N_5094,N_4624);
and U6123 (N_6123,N_5832,N_4527);
nand U6124 (N_6124,N_5722,N_4962);
nand U6125 (N_6125,N_4841,N_5479);
nand U6126 (N_6126,N_5340,N_4722);
and U6127 (N_6127,N_4783,N_4955);
nand U6128 (N_6128,N_5460,N_5775);
or U6129 (N_6129,N_4856,N_5093);
nand U6130 (N_6130,N_5928,N_4754);
nor U6131 (N_6131,N_4815,N_5918);
and U6132 (N_6132,N_4678,N_5843);
and U6133 (N_6133,N_5381,N_5091);
and U6134 (N_6134,N_5329,N_4588);
nor U6135 (N_6135,N_5271,N_5577);
or U6136 (N_6136,N_4729,N_5919);
nor U6137 (N_6137,N_5780,N_4553);
and U6138 (N_6138,N_5078,N_4762);
xnor U6139 (N_6139,N_5087,N_4635);
and U6140 (N_6140,N_4575,N_4851);
nand U6141 (N_6141,N_5207,N_4822);
or U6142 (N_6142,N_5351,N_5067);
xnor U6143 (N_6143,N_5432,N_4947);
and U6144 (N_6144,N_5600,N_5027);
nand U6145 (N_6145,N_5847,N_5002);
xnor U6146 (N_6146,N_4533,N_5229);
and U6147 (N_6147,N_5703,N_5965);
nor U6148 (N_6148,N_5260,N_4928);
and U6149 (N_6149,N_4505,N_5250);
nor U6150 (N_6150,N_5575,N_5239);
nor U6151 (N_6151,N_5729,N_5406);
nand U6152 (N_6152,N_4891,N_5540);
or U6153 (N_6153,N_5015,N_5298);
nor U6154 (N_6154,N_4694,N_5995);
and U6155 (N_6155,N_5803,N_5997);
nor U6156 (N_6156,N_5124,N_4809);
and U6157 (N_6157,N_5859,N_5019);
or U6158 (N_6158,N_5643,N_5389);
nor U6159 (N_6159,N_5878,N_5121);
nand U6160 (N_6160,N_4560,N_4733);
and U6161 (N_6161,N_5566,N_5545);
or U6162 (N_6162,N_5431,N_5408);
and U6163 (N_6163,N_4976,N_4995);
nand U6164 (N_6164,N_4888,N_5312);
or U6165 (N_6165,N_4731,N_4690);
and U6166 (N_6166,N_5115,N_5954);
nand U6167 (N_6167,N_5507,N_4889);
nor U6168 (N_6168,N_4596,N_4555);
and U6169 (N_6169,N_5786,N_5041);
nor U6170 (N_6170,N_5029,N_5166);
nand U6171 (N_6171,N_5249,N_5430);
or U6172 (N_6172,N_5958,N_5973);
and U6173 (N_6173,N_4583,N_5424);
nand U6174 (N_6174,N_4811,N_5613);
nand U6175 (N_6175,N_5710,N_4712);
nor U6176 (N_6176,N_5841,N_4518);
and U6177 (N_6177,N_5544,N_5004);
nand U6178 (N_6178,N_5723,N_5392);
nand U6179 (N_6179,N_5331,N_4645);
nand U6180 (N_6180,N_4520,N_5520);
and U6181 (N_6181,N_5120,N_5160);
or U6182 (N_6182,N_5039,N_4861);
or U6183 (N_6183,N_4860,N_4916);
nor U6184 (N_6184,N_4896,N_5148);
nor U6185 (N_6185,N_5839,N_4742);
and U6186 (N_6186,N_4927,N_5414);
nor U6187 (N_6187,N_5266,N_4883);
nand U6188 (N_6188,N_5861,N_5388);
and U6189 (N_6189,N_4675,N_4579);
nand U6190 (N_6190,N_4515,N_5110);
and U6191 (N_6191,N_4781,N_5401);
nand U6192 (N_6192,N_4938,N_5720);
xor U6193 (N_6193,N_5658,N_5122);
nand U6194 (N_6194,N_4850,N_5224);
xor U6195 (N_6195,N_5665,N_5198);
and U6196 (N_6196,N_5490,N_5556);
nand U6197 (N_6197,N_5069,N_5929);
or U6198 (N_6198,N_4777,N_5259);
nand U6199 (N_6199,N_5288,N_4507);
and U6200 (N_6200,N_5135,N_4625);
nand U6201 (N_6201,N_4913,N_4631);
or U6202 (N_6202,N_5856,N_5868);
xnor U6203 (N_6203,N_5693,N_5206);
nor U6204 (N_6204,N_5367,N_5695);
nand U6205 (N_6205,N_4903,N_5422);
or U6206 (N_6206,N_4764,N_4537);
or U6207 (N_6207,N_5730,N_5043);
nand U6208 (N_6208,N_4565,N_5967);
nand U6209 (N_6209,N_4937,N_4609);
xor U6210 (N_6210,N_5489,N_5119);
or U6211 (N_6211,N_5539,N_5055);
nor U6212 (N_6212,N_5391,N_4544);
nand U6213 (N_6213,N_5416,N_5346);
xnor U6214 (N_6214,N_5712,N_5586);
or U6215 (N_6215,N_5636,N_4597);
and U6216 (N_6216,N_5746,N_4801);
or U6217 (N_6217,N_5241,N_5302);
nand U6218 (N_6218,N_5840,N_5417);
or U6219 (N_6219,N_5042,N_4626);
nor U6220 (N_6220,N_5661,N_4686);
and U6221 (N_6221,N_4677,N_5790);
nor U6222 (N_6222,N_5532,N_4719);
and U6223 (N_6223,N_4840,N_5270);
nor U6224 (N_6224,N_4956,N_5921);
or U6225 (N_6225,N_4808,N_4989);
and U6226 (N_6226,N_4528,N_5443);
nand U6227 (N_6227,N_5278,N_5896);
nor U6228 (N_6228,N_5734,N_5360);
nand U6229 (N_6229,N_5210,N_5628);
or U6230 (N_6230,N_5793,N_4618);
and U6231 (N_6231,N_5248,N_5724);
nor U6232 (N_6232,N_4578,N_5153);
nor U6233 (N_6233,N_4866,N_5938);
nand U6234 (N_6234,N_5705,N_4826);
nor U6235 (N_6235,N_5804,N_4728);
nor U6236 (N_6236,N_5538,N_5264);
xor U6237 (N_6237,N_5713,N_5380);
xnor U6238 (N_6238,N_5175,N_5873);
nand U6239 (N_6239,N_5219,N_5498);
nand U6240 (N_6240,N_4519,N_5851);
nor U6241 (N_6241,N_5650,N_5177);
nor U6242 (N_6242,N_4939,N_4610);
and U6243 (N_6243,N_4914,N_5272);
nor U6244 (N_6244,N_5678,N_5912);
and U6245 (N_6245,N_4824,N_4831);
or U6246 (N_6246,N_5922,N_4899);
and U6247 (N_6247,N_5284,N_5307);
nand U6248 (N_6248,N_4655,N_5735);
or U6249 (N_6249,N_4922,N_5341);
nand U6250 (N_6250,N_5627,N_5588);
or U6251 (N_6251,N_5881,N_5660);
nor U6252 (N_6252,N_5364,N_5581);
or U6253 (N_6253,N_4975,N_5592);
nand U6254 (N_6254,N_5828,N_5046);
or U6255 (N_6255,N_5835,N_5512);
nor U6256 (N_6256,N_5869,N_4658);
nand U6257 (N_6257,N_4745,N_5342);
or U6258 (N_6258,N_5247,N_5728);
nand U6259 (N_6259,N_4911,N_5564);
nor U6260 (N_6260,N_5097,N_4673);
and U6261 (N_6261,N_5992,N_5118);
or U6262 (N_6262,N_4827,N_5058);
or U6263 (N_6263,N_5446,N_5457);
nand U6264 (N_6264,N_5987,N_4541);
or U6265 (N_6265,N_5548,N_4549);
or U6266 (N_6266,N_4556,N_5454);
nor U6267 (N_6267,N_5068,N_5033);
nand U6268 (N_6268,N_4551,N_5951);
and U6269 (N_6269,N_4727,N_4633);
nand U6270 (N_6270,N_5802,N_5006);
and U6271 (N_6271,N_4593,N_4766);
nand U6272 (N_6272,N_5947,N_5984);
nor U6273 (N_6273,N_4585,N_4835);
nand U6274 (N_6274,N_4957,N_5021);
or U6275 (N_6275,N_5620,N_5325);
nand U6276 (N_6276,N_4513,N_5176);
and U6277 (N_6277,N_4697,N_4748);
or U6278 (N_6278,N_5020,N_5294);
nor U6279 (N_6279,N_5552,N_5305);
nor U6280 (N_6280,N_5465,N_5103);
nand U6281 (N_6281,N_5789,N_4548);
and U6282 (N_6282,N_5450,N_4603);
or U6283 (N_6283,N_5814,N_4833);
or U6284 (N_6284,N_5760,N_5582);
nor U6285 (N_6285,N_5433,N_5109);
nand U6286 (N_6286,N_4534,N_5007);
nand U6287 (N_6287,N_5455,N_5807);
or U6288 (N_6288,N_5191,N_5066);
or U6289 (N_6289,N_5514,N_4547);
nand U6290 (N_6290,N_5317,N_4531);
nor U6291 (N_6291,N_5916,N_4680);
nor U6292 (N_6292,N_5884,N_5570);
nor U6293 (N_6293,N_5676,N_4638);
and U6294 (N_6294,N_4501,N_5025);
nand U6295 (N_6295,N_5101,N_5739);
nand U6296 (N_6296,N_5753,N_5679);
or U6297 (N_6297,N_4854,N_5232);
and U6298 (N_6298,N_5222,N_4877);
and U6299 (N_6299,N_5405,N_5001);
nor U6300 (N_6300,N_5605,N_5221);
or U6301 (N_6301,N_4689,N_5111);
or U6302 (N_6302,N_4671,N_4756);
xnor U6303 (N_6303,N_5652,N_5529);
and U6304 (N_6304,N_5865,N_5150);
xnor U6305 (N_6305,N_5274,N_5281);
nor U6306 (N_6306,N_4855,N_5102);
and U6307 (N_6307,N_5214,N_5764);
nor U6308 (N_6308,N_5427,N_4561);
xor U6309 (N_6309,N_5927,N_5083);
nor U6310 (N_6310,N_5410,N_4681);
nor U6311 (N_6311,N_5261,N_5335);
and U6312 (N_6312,N_5440,N_5711);
or U6313 (N_6313,N_4774,N_5463);
or U6314 (N_6314,N_5242,N_4859);
xnor U6315 (N_6315,N_5572,N_5253);
xnor U6316 (N_6316,N_5018,N_5336);
nor U6317 (N_6317,N_5235,N_4940);
nor U6318 (N_6318,N_5023,N_5765);
or U6319 (N_6319,N_5670,N_5766);
nand U6320 (N_6320,N_5755,N_5296);
nor U6321 (N_6321,N_4726,N_5032);
xnor U6322 (N_6322,N_5848,N_5611);
nor U6323 (N_6323,N_5379,N_5726);
or U6324 (N_6324,N_5547,N_4659);
and U6325 (N_6325,N_5064,N_4931);
or U6326 (N_6326,N_5315,N_4695);
xnor U6327 (N_6327,N_5304,N_5061);
xnor U6328 (N_6328,N_4807,N_5822);
nor U6329 (N_6329,N_5209,N_4793);
nand U6330 (N_6330,N_4679,N_5003);
and U6331 (N_6331,N_5744,N_5933);
nand U6332 (N_6332,N_5831,N_4550);
and U6333 (N_6333,N_5821,N_5812);
nand U6334 (N_6334,N_5005,N_5926);
nand U6335 (N_6335,N_4926,N_4894);
nor U6336 (N_6336,N_4688,N_5426);
and U6337 (N_6337,N_5819,N_5902);
nand U6338 (N_6338,N_4758,N_5761);
nand U6339 (N_6339,N_5199,N_5385);
nor U6340 (N_6340,N_5420,N_5378);
nor U6341 (N_6341,N_5030,N_5820);
or U6342 (N_6342,N_5413,N_5147);
and U6343 (N_6343,N_5827,N_5662);
and U6344 (N_6344,N_5128,N_4802);
and U6345 (N_6345,N_4782,N_5603);
and U6346 (N_6346,N_4693,N_4649);
nand U6347 (N_6347,N_5265,N_4572);
nand U6348 (N_6348,N_4961,N_5011);
nand U6349 (N_6349,N_4954,N_5375);
and U6350 (N_6350,N_5772,N_5200);
nor U6351 (N_6351,N_4628,N_5062);
nand U6352 (N_6352,N_4711,N_5844);
nand U6353 (N_6353,N_5034,N_5394);
and U6354 (N_6354,N_5568,N_4732);
nand U6355 (N_6355,N_4682,N_4512);
nor U6356 (N_6356,N_4703,N_5998);
and U6357 (N_6357,N_4963,N_5957);
nand U6358 (N_6358,N_5488,N_5400);
and U6359 (N_6359,N_4740,N_4595);
nor U6360 (N_6360,N_4892,N_4797);
xnor U6361 (N_6361,N_5486,N_5530);
and U6362 (N_6362,N_4941,N_4972);
nor U6363 (N_6363,N_4902,N_4977);
nor U6364 (N_6364,N_5085,N_4910);
xor U6365 (N_6365,N_5964,N_5805);
nor U6366 (N_6366,N_5497,N_5180);
xor U6367 (N_6367,N_4670,N_5971);
or U6368 (N_6368,N_5686,N_5306);
nand U6369 (N_6369,N_4640,N_4921);
or U6370 (N_6370,N_5750,N_5044);
nand U6371 (N_6371,N_5098,N_4880);
nor U6372 (N_6372,N_5645,N_5202);
nor U6373 (N_6373,N_4969,N_4769);
and U6374 (N_6374,N_4776,N_5138);
xnor U6375 (N_6375,N_5505,N_5796);
or U6376 (N_6376,N_4981,N_5886);
xnor U6377 (N_6377,N_4836,N_5518);
nor U6378 (N_6378,N_4852,N_5444);
or U6379 (N_6379,N_5752,N_5573);
and U6380 (N_6380,N_4554,N_4973);
nand U6381 (N_6381,N_4734,N_5614);
or U6382 (N_6382,N_5866,N_4943);
xnor U6383 (N_6383,N_4526,N_4735);
or U6384 (N_6384,N_5519,N_5569);
nor U6385 (N_6385,N_4812,N_5644);
or U6386 (N_6386,N_5084,N_5719);
or U6387 (N_6387,N_5112,N_5787);
nor U6388 (N_6388,N_5395,N_4886);
and U6389 (N_6389,N_5941,N_5439);
nor U6390 (N_6390,N_4825,N_5499);
nor U6391 (N_6391,N_4786,N_5516);
and U6392 (N_6392,N_5009,N_5170);
nor U6393 (N_6393,N_5894,N_5664);
and U6394 (N_6394,N_5049,N_4857);
nand U6395 (N_6395,N_5227,N_5350);
and U6396 (N_6396,N_4918,N_5438);
or U6397 (N_6397,N_4523,N_4799);
and U6398 (N_6398,N_5268,N_5511);
or U6399 (N_6399,N_5409,N_5960);
nand U6400 (N_6400,N_5870,N_5173);
and U6401 (N_6401,N_5610,N_5531);
or U6402 (N_6402,N_5810,N_5468);
and U6403 (N_6403,N_5337,N_5218);
nor U6404 (N_6404,N_5593,N_5419);
or U6405 (N_6405,N_5858,N_4761);
xor U6406 (N_6406,N_5590,N_4828);
and U6407 (N_6407,N_4558,N_5638);
nor U6408 (N_6408,N_5233,N_5404);
nor U6409 (N_6409,N_5523,N_4968);
and U6410 (N_6410,N_5959,N_5421);
nor U6411 (N_6411,N_4909,N_5901);
and U6412 (N_6412,N_5070,N_5942);
nor U6413 (N_6413,N_5762,N_5215);
or U6414 (N_6414,N_5563,N_4992);
or U6415 (N_6415,N_5680,N_5675);
and U6416 (N_6416,N_5010,N_4767);
nor U6417 (N_6417,N_5065,N_4959);
or U6418 (N_6418,N_5681,N_5273);
and U6419 (N_6419,N_5891,N_4908);
nand U6420 (N_6420,N_5275,N_5647);
or U6421 (N_6421,N_4805,N_5595);
nand U6422 (N_6422,N_4864,N_4953);
or U6423 (N_6423,N_5784,N_5633);
and U6424 (N_6424,N_5290,N_5526);
nand U6425 (N_6425,N_5872,N_5026);
nand U6426 (N_6426,N_5096,N_5188);
xor U6427 (N_6427,N_5471,N_4838);
xnor U6428 (N_6428,N_4832,N_5473);
xnor U6429 (N_6429,N_5204,N_5412);
and U6430 (N_6430,N_5666,N_4964);
and U6431 (N_6431,N_5179,N_5157);
and U6432 (N_6432,N_5048,N_5690);
nor U6433 (N_6433,N_5012,N_5038);
nor U6434 (N_6434,N_4616,N_5267);
or U6435 (N_6435,N_5576,N_5151);
or U6436 (N_6436,N_4569,N_4869);
or U6437 (N_6437,N_5616,N_4737);
and U6438 (N_6438,N_5996,N_5187);
or U6439 (N_6439,N_4771,N_5709);
nand U6440 (N_6440,N_5436,N_4944);
nand U6441 (N_6441,N_5758,N_5800);
nor U6442 (N_6442,N_5133,N_4893);
nand U6443 (N_6443,N_5905,N_5081);
or U6444 (N_6444,N_4749,N_5154);
or U6445 (N_6445,N_4614,N_5050);
or U6446 (N_6446,N_4525,N_5167);
and U6447 (N_6447,N_5024,N_5860);
or U6448 (N_6448,N_5190,N_5319);
nand U6449 (N_6449,N_5682,N_4714);
nand U6450 (N_6450,N_4876,N_4798);
and U6451 (N_6451,N_5671,N_4514);
and U6452 (N_6452,N_5792,N_5663);
or U6453 (N_6453,N_5090,N_5040);
and U6454 (N_6454,N_4738,N_4746);
nor U6455 (N_6455,N_4942,N_5551);
or U6456 (N_6456,N_5487,N_5612);
and U6457 (N_6457,N_4521,N_5316);
or U6458 (N_6458,N_5685,N_5470);
nand U6459 (N_6459,N_5054,N_4599);
nor U6460 (N_6460,N_4881,N_5899);
or U6461 (N_6461,N_5931,N_5904);
nor U6462 (N_6462,N_4594,N_5366);
nand U6463 (N_6463,N_4804,N_5126);
or U6464 (N_6464,N_5142,N_5537);
or U6465 (N_6465,N_5494,N_4753);
nor U6466 (N_6466,N_5144,N_5324);
xnor U6467 (N_6467,N_4897,N_5088);
nand U6468 (N_6468,N_5300,N_4539);
nand U6469 (N_6469,N_4929,N_5898);
xnor U6470 (N_6470,N_5757,N_4590);
or U6471 (N_6471,N_5056,N_5435);
or U6472 (N_6472,N_5481,N_5798);
and U6473 (N_6473,N_5037,N_4979);
and U6474 (N_6474,N_5541,N_5754);
or U6475 (N_6475,N_5677,N_5558);
nor U6476 (N_6476,N_5795,N_5333);
and U6477 (N_6477,N_5483,N_5699);
or U6478 (N_6478,N_4692,N_5808);
nor U6479 (N_6479,N_5963,N_5347);
nand U6480 (N_6480,N_5824,N_4589);
xnor U6481 (N_6481,N_5626,N_4630);
or U6482 (N_6482,N_4967,N_4810);
nor U6483 (N_6483,N_5343,N_4571);
or U6484 (N_6484,N_5159,N_4642);
xnor U6485 (N_6485,N_5445,N_5906);
nand U6486 (N_6486,N_4730,N_5818);
and U6487 (N_6487,N_4522,N_5231);
nand U6488 (N_6488,N_5970,N_4718);
nor U6489 (N_6489,N_5509,N_5362);
or U6490 (N_6490,N_5591,N_5788);
and U6491 (N_6491,N_5578,N_5834);
nor U6492 (N_6492,N_4636,N_4511);
and U6493 (N_6493,N_5382,N_5657);
or U6494 (N_6494,N_5437,N_5155);
and U6495 (N_6495,N_5071,N_5738);
nor U6496 (N_6496,N_4946,N_5817);
and U6497 (N_6497,N_5517,N_5129);
or U6498 (N_6498,N_5510,N_5477);
nor U6499 (N_6499,N_5472,N_4653);
nor U6500 (N_6500,N_5778,N_5871);
and U6501 (N_6501,N_4598,N_5687);
and U6502 (N_6502,N_5846,N_4627);
and U6503 (N_6503,N_5036,N_5743);
or U6504 (N_6504,N_4760,N_5893);
and U6505 (N_6505,N_5604,N_5449);
nor U6506 (N_6506,N_4637,N_4700);
and U6507 (N_6507,N_5292,N_5073);
and U6508 (N_6508,N_4985,N_5469);
and U6509 (N_6509,N_4988,N_4991);
nor U6510 (N_6510,N_5580,N_5277);
nand U6511 (N_6511,N_5903,N_5060);
nor U6512 (N_6512,N_5943,N_5914);
nor U6513 (N_6513,N_5885,N_5988);
or U6514 (N_6514,N_5508,N_4999);
and U6515 (N_6515,N_4936,N_4724);
and U6516 (N_6516,N_5283,N_4853);
nand U6517 (N_6517,N_4849,N_5782);
and U6518 (N_6518,N_5377,N_4510);
nor U6519 (N_6519,N_5606,N_4986);
nor U6520 (N_6520,N_5452,N_5716);
xor U6521 (N_6521,N_4739,N_5913);
nor U6522 (N_6522,N_5771,N_5211);
and U6523 (N_6523,N_5195,N_5156);
or U6524 (N_6524,N_4586,N_5924);
or U6525 (N_6525,N_4698,N_5609);
nor U6526 (N_6526,N_5348,N_4660);
nand U6527 (N_6527,N_5165,N_4993);
and U6528 (N_6528,N_5076,N_5522);
or U6529 (N_6529,N_4858,N_5399);
and U6530 (N_6530,N_5017,N_4580);
and U6531 (N_6531,N_5560,N_4600);
xnor U6532 (N_6532,N_5225,N_5461);
and U6533 (N_6533,N_5632,N_4691);
and U6534 (N_6534,N_5631,N_5920);
and U6535 (N_6535,N_5075,N_4562);
and U6536 (N_6536,N_4647,N_5909);
and U6537 (N_6537,N_4701,N_4704);
nand U6538 (N_6538,N_5930,N_5208);
or U6539 (N_6539,N_4604,N_4879);
nand U6540 (N_6540,N_5082,N_5356);
nor U6541 (N_6541,N_4668,N_4536);
nor U6542 (N_6542,N_5655,N_5654);
xor U6543 (N_6543,N_5799,N_4789);
or U6544 (N_6544,N_4862,N_5940);
and U6545 (N_6545,N_4744,N_4644);
and U6546 (N_6546,N_5365,N_4617);
or U6547 (N_6547,N_4935,N_5700);
and U6548 (N_6548,N_5731,N_4932);
and U6549 (N_6549,N_4983,N_5689);
nand U6550 (N_6550,N_5374,N_5776);
or U6551 (N_6551,N_5243,N_5917);
nand U6552 (N_6552,N_4987,N_5767);
nor U6553 (N_6553,N_5651,N_4950);
xnor U6554 (N_6554,N_5258,N_5475);
xor U6555 (N_6555,N_5134,N_5100);
nor U6556 (N_6556,N_5667,N_5353);
and U6557 (N_6557,N_5624,N_5727);
nand U6558 (N_6558,N_5791,N_5000);
and U6559 (N_6559,N_5953,N_4773);
or U6560 (N_6560,N_5252,N_4752);
nor U6561 (N_6561,N_5635,N_4634);
and U6562 (N_6562,N_5701,N_4907);
nand U6563 (N_6563,N_5684,N_4606);
nand U6564 (N_6564,N_4530,N_5867);
nor U6565 (N_6565,N_5328,N_5536);
or U6566 (N_6566,N_4552,N_5372);
and U6567 (N_6567,N_4874,N_5125);
and U6568 (N_6568,N_5543,N_5503);
xnor U6569 (N_6569,N_5864,N_4814);
and U6570 (N_6570,N_5785,N_5583);
or U6571 (N_6571,N_5619,N_5978);
xor U6572 (N_6572,N_5513,N_5559);
and U6573 (N_6573,N_5107,N_5574);
xor U6574 (N_6574,N_5251,N_4878);
or U6575 (N_6575,N_5562,N_5646);
and U6576 (N_6576,N_5467,N_5263);
and U6577 (N_6577,N_4715,N_4676);
or U6578 (N_6578,N_5571,N_4545);
and U6579 (N_6579,N_5816,N_5554);
and U6580 (N_6580,N_5952,N_5607);
or U6581 (N_6581,N_4900,N_4621);
xnor U6582 (N_6582,N_5116,N_4699);
nor U6583 (N_6583,N_4665,N_5149);
and U6584 (N_6584,N_5137,N_5751);
nand U6585 (N_6585,N_5114,N_5875);
nand U6586 (N_6586,N_4546,N_5052);
nor U6587 (N_6587,N_4538,N_5397);
and U6588 (N_6588,N_5145,N_5579);
nand U6589 (N_6589,N_4919,N_4949);
xor U6590 (N_6590,N_5393,N_4791);
or U6591 (N_6591,N_5217,N_5141);
or U6592 (N_6592,N_4564,N_4684);
xor U6593 (N_6593,N_5966,N_4535);
xor U6594 (N_6594,N_4780,N_5113);
nor U6595 (N_6595,N_5189,N_5567);
and U6596 (N_6596,N_5815,N_4800);
or U6597 (N_6597,N_4779,N_5774);
nand U6598 (N_6598,N_5063,N_4870);
xnor U6599 (N_6599,N_5777,N_5047);
and U6600 (N_6600,N_5797,N_5742);
nand U6601 (N_6601,N_4915,N_5311);
nor U6602 (N_6602,N_5286,N_5506);
nand U6603 (N_6603,N_5293,N_4865);
nand U6604 (N_6604,N_5234,N_5991);
nor U6605 (N_6605,N_5466,N_5092);
nand U6606 (N_6606,N_5447,N_5584);
nor U6607 (N_6607,N_5059,N_4629);
or U6608 (N_6608,N_5402,N_4796);
nor U6609 (N_6609,N_5186,N_5975);
or U6610 (N_6610,N_5981,N_4529);
nor U6611 (N_6611,N_5648,N_4662);
and U6612 (N_6612,N_5164,N_5806);
or U6613 (N_6613,N_4775,N_5597);
nor U6614 (N_6614,N_4557,N_4847);
or U6615 (N_6615,N_5972,N_4792);
nor U6616 (N_6616,N_5637,N_5669);
nor U6617 (N_6617,N_4592,N_5594);
or U6618 (N_6618,N_4818,N_5985);
or U6619 (N_6619,N_5911,N_4696);
nor U6620 (N_6620,N_5303,N_5876);
and U6621 (N_6621,N_4904,N_5480);
or U6622 (N_6622,N_5181,N_5900);
nand U6623 (N_6623,N_4945,N_5203);
and U6624 (N_6624,N_5718,N_5442);
or U6625 (N_6625,N_5482,N_5704);
and U6626 (N_6626,N_4516,N_4923);
or U6627 (N_6627,N_5171,N_4794);
nor U6628 (N_6628,N_5668,N_4765);
xor U6629 (N_6629,N_5492,N_4971);
or U6630 (N_6630,N_5086,N_5246);
nand U6631 (N_6631,N_5355,N_5376);
nand U6632 (N_6632,N_5602,N_5254);
or U6633 (N_6633,N_5948,N_5639);
or U6634 (N_6634,N_5979,N_5297);
nand U6635 (N_6635,N_4757,N_4834);
or U6636 (N_6636,N_5908,N_4830);
or U6637 (N_6637,N_4952,N_5456);
nor U6638 (N_6638,N_4920,N_5415);
nor U6639 (N_6639,N_5314,N_5854);
and U6640 (N_6640,N_5589,N_5608);
nand U6641 (N_6641,N_5240,N_5944);
nand U6642 (N_6642,N_5640,N_5553);
nand U6643 (N_6643,N_4666,N_5617);
or U6644 (N_6644,N_5874,N_5811);
nand U6645 (N_6645,N_5534,N_5493);
nor U6646 (N_6646,N_5425,N_4917);
and U6647 (N_6647,N_5192,N_4685);
nor U6648 (N_6648,N_5838,N_5226);
and U6649 (N_6649,N_5707,N_5887);
or U6650 (N_6650,N_5396,N_4710);
xnor U6651 (N_6651,N_5549,N_5237);
or U6652 (N_6652,N_5428,N_5857);
and U6653 (N_6653,N_4608,N_5496);
and U6654 (N_6654,N_5770,N_5371);
and U6655 (N_6655,N_5696,N_5462);
nand U6656 (N_6656,N_4930,N_5184);
or U6657 (N_6657,N_4736,N_4951);
nand U6658 (N_6658,N_5533,N_5649);
or U6659 (N_6659,N_4990,N_5634);
or U6660 (N_6660,N_5140,N_5321);
xor U6661 (N_6661,N_4844,N_5291);
or U6662 (N_6662,N_5474,N_5698);
or U6663 (N_6663,N_5338,N_4906);
and U6664 (N_6664,N_5986,N_5745);
and U6665 (N_6665,N_4584,N_5080);
xnor U6666 (N_6666,N_5289,N_4863);
and U6667 (N_6667,N_5282,N_4620);
nor U6668 (N_6668,N_5478,N_4819);
or U6669 (N_6669,N_5740,N_5749);
nand U6670 (N_6670,N_4705,N_4751);
nor U6671 (N_6671,N_4613,N_5130);
or U6672 (N_6672,N_5976,N_5352);
nand U6673 (N_6673,N_5172,N_4795);
nand U6674 (N_6674,N_5932,N_5016);
nor U6675 (N_6675,N_5955,N_5127);
or U6676 (N_6676,N_4898,N_5236);
and U6677 (N_6677,N_5357,N_5183);
or U6678 (N_6678,N_5108,N_5105);
or U6679 (N_6679,N_5332,N_4816);
and U6680 (N_6680,N_5826,N_5692);
nand U6681 (N_6681,N_4623,N_5451);
nand U6682 (N_6682,N_4581,N_4884);
and U6683 (N_6683,N_4587,N_4933);
and U6684 (N_6684,N_5596,N_5320);
or U6685 (N_6685,N_5429,N_4540);
nand U6686 (N_6686,N_4656,N_5196);
or U6687 (N_6687,N_4763,N_5182);
nand U6688 (N_6688,N_5897,N_5448);
nor U6689 (N_6689,N_5993,N_5028);
and U6690 (N_6690,N_4669,N_4532);
nand U6691 (N_6691,N_5546,N_5688);
xor U6692 (N_6692,N_4574,N_5123);
and U6693 (N_6693,N_5845,N_4965);
or U6694 (N_6694,N_5842,N_5794);
nor U6695 (N_6695,N_4706,N_5825);
nand U6696 (N_6696,N_5276,N_5621);
or U6697 (N_6697,N_5035,N_5697);
nor U6698 (N_6698,N_4508,N_5829);
or U6699 (N_6699,N_5095,N_4829);
nand U6700 (N_6700,N_4741,N_5174);
and U6701 (N_6701,N_5714,N_5201);
nand U6702 (N_6702,N_4502,N_4639);
nor U6703 (N_6703,N_4785,N_5557);
nor U6704 (N_6704,N_5850,N_5369);
or U6705 (N_6705,N_5387,N_5962);
or U6706 (N_6706,N_5363,N_4716);
nand U6707 (N_6707,N_5212,N_5403);
nor U6708 (N_6708,N_5555,N_5615);
nor U6709 (N_6709,N_4823,N_4803);
and U6710 (N_6710,N_4787,N_4563);
or U6711 (N_6711,N_4573,N_5299);
and U6712 (N_6712,N_5855,N_5441);
and U6713 (N_6713,N_5484,N_5702);
and U6714 (N_6714,N_5500,N_5072);
and U6715 (N_6715,N_4654,N_4559);
or U6716 (N_6716,N_5715,N_4759);
or U6717 (N_6717,N_5656,N_4664);
or U6718 (N_6718,N_4646,N_4974);
and U6719 (N_6719,N_4500,N_4708);
or U6720 (N_6720,N_5880,N_4868);
nand U6721 (N_6721,N_4885,N_4687);
or U6722 (N_6722,N_5629,N_5022);
nor U6723 (N_6723,N_5587,N_5220);
nor U6724 (N_6724,N_5280,N_5057);
or U6725 (N_6725,N_5244,N_4970);
nor U6726 (N_6726,N_5923,N_4674);
or U6727 (N_6727,N_4725,N_4966);
xnor U6728 (N_6728,N_5051,N_5434);
and U6729 (N_6729,N_5301,N_5458);
and U6730 (N_6730,N_5158,N_5089);
nor U6731 (N_6731,N_4784,N_4577);
xnor U6732 (N_6732,N_5732,N_5706);
and U6733 (N_6733,N_5737,N_5550);
nand U6734 (N_6734,N_4601,N_5659);
nor U6735 (N_6735,N_5598,N_5368);
nand U6736 (N_6736,N_4817,N_5939);
or U6737 (N_6737,N_4845,N_5625);
or U6738 (N_6738,N_5515,N_5721);
nor U6739 (N_6739,N_5255,N_4905);
xor U6740 (N_6740,N_4788,N_5262);
nor U6741 (N_6741,N_5031,N_5146);
and U6742 (N_6742,N_4912,N_5618);
and U6743 (N_6743,N_4709,N_4873);
nand U6744 (N_6744,N_4657,N_4605);
nor U6745 (N_6745,N_4837,N_4901);
nor U6746 (N_6746,N_5386,N_5330);
nor U6747 (N_6747,N_4641,N_5230);
or U6748 (N_6748,N_5373,N_5969);
xor U6749 (N_6749,N_4720,N_4643);
nand U6750 (N_6750,N_5314,N_4946);
or U6751 (N_6751,N_5241,N_5370);
nor U6752 (N_6752,N_5423,N_4553);
nor U6753 (N_6753,N_5012,N_5579);
xor U6754 (N_6754,N_5244,N_5093);
nand U6755 (N_6755,N_4704,N_5922);
nand U6756 (N_6756,N_5820,N_4617);
nor U6757 (N_6757,N_5982,N_5313);
nor U6758 (N_6758,N_5010,N_4910);
nand U6759 (N_6759,N_5657,N_5413);
and U6760 (N_6760,N_4899,N_5790);
or U6761 (N_6761,N_5569,N_5503);
nor U6762 (N_6762,N_5173,N_4534);
and U6763 (N_6763,N_5258,N_5565);
nand U6764 (N_6764,N_5200,N_5581);
xor U6765 (N_6765,N_5279,N_5666);
nand U6766 (N_6766,N_5219,N_4902);
nand U6767 (N_6767,N_5775,N_5139);
and U6768 (N_6768,N_5346,N_4567);
nand U6769 (N_6769,N_5589,N_4919);
nand U6770 (N_6770,N_5980,N_5299);
nand U6771 (N_6771,N_4943,N_5133);
or U6772 (N_6772,N_5686,N_4870);
nor U6773 (N_6773,N_5916,N_4924);
or U6774 (N_6774,N_5200,N_4645);
nor U6775 (N_6775,N_4523,N_4777);
xor U6776 (N_6776,N_4969,N_5887);
nor U6777 (N_6777,N_4528,N_5514);
or U6778 (N_6778,N_5862,N_5084);
or U6779 (N_6779,N_5906,N_5095);
nand U6780 (N_6780,N_5620,N_5059);
xor U6781 (N_6781,N_5922,N_5446);
or U6782 (N_6782,N_4815,N_5218);
nand U6783 (N_6783,N_4560,N_5497);
and U6784 (N_6784,N_5682,N_5244);
and U6785 (N_6785,N_5209,N_5350);
nand U6786 (N_6786,N_5260,N_4871);
or U6787 (N_6787,N_5651,N_5448);
and U6788 (N_6788,N_5133,N_4867);
xnor U6789 (N_6789,N_4586,N_4880);
or U6790 (N_6790,N_4601,N_5092);
nor U6791 (N_6791,N_5701,N_4920);
and U6792 (N_6792,N_5656,N_4834);
nor U6793 (N_6793,N_4531,N_4909);
nor U6794 (N_6794,N_5861,N_5468);
and U6795 (N_6795,N_4681,N_4750);
nand U6796 (N_6796,N_5547,N_4529);
nor U6797 (N_6797,N_4974,N_4670);
nor U6798 (N_6798,N_4565,N_5046);
nand U6799 (N_6799,N_5554,N_5514);
xnor U6800 (N_6800,N_5912,N_5300);
xor U6801 (N_6801,N_5444,N_5778);
xnor U6802 (N_6802,N_5084,N_4542);
and U6803 (N_6803,N_4719,N_5442);
and U6804 (N_6804,N_4580,N_5314);
or U6805 (N_6805,N_5404,N_5200);
nor U6806 (N_6806,N_4925,N_5329);
nor U6807 (N_6807,N_5058,N_4889);
nand U6808 (N_6808,N_5616,N_4871);
nand U6809 (N_6809,N_4900,N_5436);
nor U6810 (N_6810,N_5624,N_4569);
or U6811 (N_6811,N_5447,N_4944);
and U6812 (N_6812,N_4950,N_4565);
nand U6813 (N_6813,N_5238,N_5847);
xnor U6814 (N_6814,N_5429,N_5707);
nand U6815 (N_6815,N_5822,N_4523);
and U6816 (N_6816,N_4726,N_4553);
and U6817 (N_6817,N_4790,N_5709);
or U6818 (N_6818,N_4634,N_5654);
or U6819 (N_6819,N_5311,N_5877);
or U6820 (N_6820,N_5473,N_5137);
xnor U6821 (N_6821,N_5795,N_4916);
and U6822 (N_6822,N_4957,N_4618);
nand U6823 (N_6823,N_5942,N_5738);
nor U6824 (N_6824,N_5768,N_5931);
and U6825 (N_6825,N_5454,N_4933);
or U6826 (N_6826,N_4548,N_5858);
nor U6827 (N_6827,N_4887,N_5524);
or U6828 (N_6828,N_4529,N_5997);
and U6829 (N_6829,N_5083,N_5657);
and U6830 (N_6830,N_4963,N_5880);
or U6831 (N_6831,N_5733,N_5218);
and U6832 (N_6832,N_5373,N_5474);
or U6833 (N_6833,N_5609,N_5243);
nor U6834 (N_6834,N_5971,N_4938);
or U6835 (N_6835,N_4582,N_5155);
and U6836 (N_6836,N_5582,N_5048);
and U6837 (N_6837,N_5820,N_5683);
or U6838 (N_6838,N_4916,N_5631);
or U6839 (N_6839,N_5161,N_5067);
nand U6840 (N_6840,N_5576,N_4779);
xor U6841 (N_6841,N_4729,N_5640);
nor U6842 (N_6842,N_5351,N_4704);
nor U6843 (N_6843,N_5253,N_4588);
and U6844 (N_6844,N_5988,N_4927);
and U6845 (N_6845,N_5105,N_5898);
and U6846 (N_6846,N_4625,N_4937);
nor U6847 (N_6847,N_5767,N_4613);
or U6848 (N_6848,N_5597,N_5092);
nand U6849 (N_6849,N_5234,N_5633);
or U6850 (N_6850,N_5504,N_4686);
nor U6851 (N_6851,N_4616,N_5961);
and U6852 (N_6852,N_4512,N_5800);
xnor U6853 (N_6853,N_5277,N_5146);
nor U6854 (N_6854,N_5265,N_5031);
nand U6855 (N_6855,N_5988,N_4881);
nor U6856 (N_6856,N_4705,N_5275);
or U6857 (N_6857,N_4747,N_5593);
and U6858 (N_6858,N_5217,N_5043);
nor U6859 (N_6859,N_5418,N_5537);
and U6860 (N_6860,N_5778,N_5780);
and U6861 (N_6861,N_5028,N_5098);
xor U6862 (N_6862,N_4958,N_5239);
nor U6863 (N_6863,N_5640,N_5582);
and U6864 (N_6864,N_4799,N_4876);
or U6865 (N_6865,N_4556,N_5270);
and U6866 (N_6866,N_4665,N_5442);
and U6867 (N_6867,N_5387,N_5424);
nor U6868 (N_6868,N_5536,N_4770);
and U6869 (N_6869,N_4818,N_5346);
nand U6870 (N_6870,N_4516,N_4993);
and U6871 (N_6871,N_5749,N_5282);
and U6872 (N_6872,N_5003,N_5982);
nand U6873 (N_6873,N_4887,N_5077);
nand U6874 (N_6874,N_5842,N_5011);
nor U6875 (N_6875,N_4626,N_5360);
nand U6876 (N_6876,N_4851,N_5927);
nand U6877 (N_6877,N_5540,N_5349);
nor U6878 (N_6878,N_4617,N_4789);
or U6879 (N_6879,N_4797,N_5850);
and U6880 (N_6880,N_5321,N_5666);
and U6881 (N_6881,N_4865,N_4848);
and U6882 (N_6882,N_4637,N_5218);
xnor U6883 (N_6883,N_4928,N_4702);
nand U6884 (N_6884,N_5289,N_4983);
or U6885 (N_6885,N_4898,N_4570);
and U6886 (N_6886,N_5025,N_5188);
nand U6887 (N_6887,N_5518,N_4872);
nand U6888 (N_6888,N_5220,N_5957);
and U6889 (N_6889,N_5779,N_5703);
and U6890 (N_6890,N_5575,N_5794);
xnor U6891 (N_6891,N_5772,N_5622);
nand U6892 (N_6892,N_5040,N_4916);
xnor U6893 (N_6893,N_4863,N_5721);
nor U6894 (N_6894,N_4800,N_4962);
xnor U6895 (N_6895,N_5698,N_5491);
nor U6896 (N_6896,N_4954,N_4579);
nand U6897 (N_6897,N_5573,N_4571);
nor U6898 (N_6898,N_5762,N_4969);
nand U6899 (N_6899,N_5352,N_5782);
or U6900 (N_6900,N_5322,N_5400);
and U6901 (N_6901,N_5707,N_4636);
and U6902 (N_6902,N_5124,N_5174);
or U6903 (N_6903,N_4918,N_4673);
nand U6904 (N_6904,N_4728,N_4986);
and U6905 (N_6905,N_5407,N_5467);
nor U6906 (N_6906,N_5928,N_5898);
nand U6907 (N_6907,N_5998,N_5044);
xnor U6908 (N_6908,N_4877,N_4901);
nand U6909 (N_6909,N_5662,N_5418);
xnor U6910 (N_6910,N_5656,N_5790);
and U6911 (N_6911,N_5422,N_4550);
nor U6912 (N_6912,N_5064,N_4606);
or U6913 (N_6913,N_5385,N_5444);
and U6914 (N_6914,N_5181,N_4551);
nor U6915 (N_6915,N_5592,N_5127);
and U6916 (N_6916,N_4919,N_5769);
or U6917 (N_6917,N_5679,N_5501);
nand U6918 (N_6918,N_5233,N_5636);
nand U6919 (N_6919,N_5669,N_5991);
nor U6920 (N_6920,N_5528,N_5804);
or U6921 (N_6921,N_5120,N_5698);
or U6922 (N_6922,N_5538,N_4969);
nand U6923 (N_6923,N_5886,N_4719);
nor U6924 (N_6924,N_4605,N_5411);
or U6925 (N_6925,N_4609,N_4630);
and U6926 (N_6926,N_5929,N_5868);
nand U6927 (N_6927,N_5069,N_5567);
nor U6928 (N_6928,N_5234,N_5859);
or U6929 (N_6929,N_5301,N_4698);
or U6930 (N_6930,N_5617,N_5293);
nand U6931 (N_6931,N_5170,N_5035);
or U6932 (N_6932,N_5863,N_4510);
nand U6933 (N_6933,N_5631,N_4787);
and U6934 (N_6934,N_4726,N_4625);
and U6935 (N_6935,N_5836,N_4960);
xnor U6936 (N_6936,N_5342,N_5184);
and U6937 (N_6937,N_5569,N_5058);
nor U6938 (N_6938,N_4541,N_5975);
and U6939 (N_6939,N_4660,N_5107);
nand U6940 (N_6940,N_4787,N_4930);
or U6941 (N_6941,N_4925,N_5899);
xnor U6942 (N_6942,N_5142,N_4843);
and U6943 (N_6943,N_5746,N_5990);
and U6944 (N_6944,N_5030,N_5217);
nor U6945 (N_6945,N_5834,N_5797);
nand U6946 (N_6946,N_5408,N_4807);
nor U6947 (N_6947,N_5074,N_5295);
nand U6948 (N_6948,N_5551,N_4511);
nand U6949 (N_6949,N_5879,N_5460);
and U6950 (N_6950,N_5189,N_5824);
nand U6951 (N_6951,N_5984,N_5530);
xor U6952 (N_6952,N_5736,N_5274);
nor U6953 (N_6953,N_4640,N_5741);
or U6954 (N_6954,N_4710,N_4578);
nand U6955 (N_6955,N_4853,N_4970);
nor U6956 (N_6956,N_5191,N_5008);
nand U6957 (N_6957,N_5364,N_5737);
or U6958 (N_6958,N_4685,N_5997);
and U6959 (N_6959,N_5353,N_5317);
xnor U6960 (N_6960,N_4845,N_5540);
and U6961 (N_6961,N_5808,N_5769);
nand U6962 (N_6962,N_5399,N_4579);
or U6963 (N_6963,N_4719,N_5468);
and U6964 (N_6964,N_5179,N_4752);
nand U6965 (N_6965,N_5687,N_5566);
nand U6966 (N_6966,N_4583,N_4804);
or U6967 (N_6967,N_4953,N_4508);
nor U6968 (N_6968,N_5753,N_5813);
nor U6969 (N_6969,N_4915,N_4631);
xor U6970 (N_6970,N_5747,N_5731);
nor U6971 (N_6971,N_5229,N_4508);
and U6972 (N_6972,N_4888,N_4668);
and U6973 (N_6973,N_4957,N_5332);
nand U6974 (N_6974,N_4565,N_4753);
xnor U6975 (N_6975,N_5822,N_5293);
or U6976 (N_6976,N_5427,N_4787);
or U6977 (N_6977,N_5570,N_5043);
xor U6978 (N_6978,N_5342,N_4993);
or U6979 (N_6979,N_5684,N_5027);
nand U6980 (N_6980,N_5844,N_4530);
or U6981 (N_6981,N_5894,N_4702);
or U6982 (N_6982,N_5364,N_4750);
and U6983 (N_6983,N_5565,N_4658);
nor U6984 (N_6984,N_4633,N_5516);
nor U6985 (N_6985,N_4822,N_5451);
nor U6986 (N_6986,N_5958,N_5740);
nand U6987 (N_6987,N_5135,N_5130);
or U6988 (N_6988,N_5443,N_5197);
nor U6989 (N_6989,N_5443,N_5217);
or U6990 (N_6990,N_5422,N_4839);
nor U6991 (N_6991,N_4610,N_4533);
and U6992 (N_6992,N_4869,N_4639);
nand U6993 (N_6993,N_5901,N_5711);
nand U6994 (N_6994,N_5404,N_4705);
xor U6995 (N_6995,N_5395,N_5474);
or U6996 (N_6996,N_5177,N_4671);
or U6997 (N_6997,N_4648,N_5497);
xor U6998 (N_6998,N_5699,N_4647);
nor U6999 (N_6999,N_5017,N_5268);
xor U7000 (N_7000,N_5970,N_5190);
or U7001 (N_7001,N_5299,N_5437);
nand U7002 (N_7002,N_5526,N_5693);
or U7003 (N_7003,N_5408,N_5058);
and U7004 (N_7004,N_5195,N_5053);
nand U7005 (N_7005,N_5198,N_5399);
nor U7006 (N_7006,N_5046,N_4973);
and U7007 (N_7007,N_5527,N_5089);
or U7008 (N_7008,N_5351,N_5261);
or U7009 (N_7009,N_4563,N_5185);
nand U7010 (N_7010,N_5220,N_4605);
xor U7011 (N_7011,N_5918,N_5129);
and U7012 (N_7012,N_5094,N_5509);
nor U7013 (N_7013,N_5941,N_5355);
or U7014 (N_7014,N_5103,N_5293);
and U7015 (N_7015,N_5207,N_5385);
or U7016 (N_7016,N_5213,N_5049);
nand U7017 (N_7017,N_4970,N_5959);
nand U7018 (N_7018,N_5580,N_5717);
or U7019 (N_7019,N_5530,N_5059);
or U7020 (N_7020,N_5401,N_5923);
xnor U7021 (N_7021,N_5385,N_4651);
or U7022 (N_7022,N_5942,N_4856);
nor U7023 (N_7023,N_5672,N_4662);
and U7024 (N_7024,N_5292,N_5683);
nand U7025 (N_7025,N_5949,N_5874);
and U7026 (N_7026,N_5528,N_4585);
xor U7027 (N_7027,N_5379,N_5752);
nand U7028 (N_7028,N_5365,N_5603);
nand U7029 (N_7029,N_4640,N_5668);
and U7030 (N_7030,N_5053,N_4777);
xnor U7031 (N_7031,N_5190,N_5438);
xnor U7032 (N_7032,N_5144,N_5239);
and U7033 (N_7033,N_4597,N_4979);
nor U7034 (N_7034,N_4694,N_4647);
nand U7035 (N_7035,N_4924,N_4547);
nor U7036 (N_7036,N_4959,N_4783);
and U7037 (N_7037,N_5918,N_4961);
or U7038 (N_7038,N_4973,N_5475);
nand U7039 (N_7039,N_5880,N_5367);
nor U7040 (N_7040,N_5164,N_5239);
nand U7041 (N_7041,N_4534,N_5246);
nand U7042 (N_7042,N_5061,N_4575);
nand U7043 (N_7043,N_4534,N_5578);
nand U7044 (N_7044,N_5343,N_5841);
nand U7045 (N_7045,N_5891,N_4728);
and U7046 (N_7046,N_5811,N_5081);
and U7047 (N_7047,N_5613,N_5379);
nor U7048 (N_7048,N_4569,N_4896);
nor U7049 (N_7049,N_5308,N_4937);
nand U7050 (N_7050,N_4531,N_4739);
nor U7051 (N_7051,N_5683,N_4739);
or U7052 (N_7052,N_5149,N_5145);
or U7053 (N_7053,N_4747,N_5695);
and U7054 (N_7054,N_5910,N_5763);
nand U7055 (N_7055,N_4950,N_4817);
nor U7056 (N_7056,N_5789,N_5506);
and U7057 (N_7057,N_5127,N_4955);
and U7058 (N_7058,N_5598,N_5138);
and U7059 (N_7059,N_5350,N_5211);
nand U7060 (N_7060,N_5113,N_5812);
or U7061 (N_7061,N_5733,N_5892);
xnor U7062 (N_7062,N_4815,N_5590);
xor U7063 (N_7063,N_5695,N_5956);
nor U7064 (N_7064,N_5346,N_5866);
or U7065 (N_7065,N_5103,N_5812);
nor U7066 (N_7066,N_5878,N_5416);
xnor U7067 (N_7067,N_4972,N_5846);
nand U7068 (N_7068,N_5711,N_4838);
and U7069 (N_7069,N_5011,N_4512);
nand U7070 (N_7070,N_5608,N_5667);
and U7071 (N_7071,N_5515,N_5398);
or U7072 (N_7072,N_5426,N_5963);
or U7073 (N_7073,N_5941,N_5391);
and U7074 (N_7074,N_5609,N_5904);
and U7075 (N_7075,N_5065,N_5937);
and U7076 (N_7076,N_4538,N_4674);
nor U7077 (N_7077,N_5486,N_5421);
or U7078 (N_7078,N_5499,N_4643);
nor U7079 (N_7079,N_5941,N_5343);
and U7080 (N_7080,N_4949,N_5148);
nand U7081 (N_7081,N_5444,N_5476);
and U7082 (N_7082,N_4564,N_5302);
nand U7083 (N_7083,N_5805,N_5006);
nor U7084 (N_7084,N_5889,N_5418);
and U7085 (N_7085,N_4826,N_5166);
and U7086 (N_7086,N_5867,N_5354);
and U7087 (N_7087,N_5391,N_4967);
nand U7088 (N_7088,N_4905,N_5414);
xor U7089 (N_7089,N_4805,N_4787);
nor U7090 (N_7090,N_5221,N_5202);
nor U7091 (N_7091,N_4915,N_4524);
nor U7092 (N_7092,N_5033,N_4548);
or U7093 (N_7093,N_4906,N_4682);
or U7094 (N_7094,N_5076,N_5376);
nand U7095 (N_7095,N_4550,N_5548);
nor U7096 (N_7096,N_5946,N_5351);
nand U7097 (N_7097,N_5556,N_4716);
nor U7098 (N_7098,N_5835,N_5468);
or U7099 (N_7099,N_4869,N_5891);
and U7100 (N_7100,N_5541,N_5096);
and U7101 (N_7101,N_5197,N_5614);
nor U7102 (N_7102,N_4846,N_5958);
nor U7103 (N_7103,N_5389,N_5117);
nor U7104 (N_7104,N_5220,N_5688);
nor U7105 (N_7105,N_5485,N_5416);
or U7106 (N_7106,N_5252,N_5295);
or U7107 (N_7107,N_5821,N_5178);
nor U7108 (N_7108,N_5205,N_5350);
or U7109 (N_7109,N_5973,N_4920);
nand U7110 (N_7110,N_5347,N_4861);
or U7111 (N_7111,N_5109,N_4534);
nor U7112 (N_7112,N_5559,N_4579);
xor U7113 (N_7113,N_5895,N_4566);
or U7114 (N_7114,N_5215,N_5410);
nor U7115 (N_7115,N_4953,N_5843);
or U7116 (N_7116,N_5391,N_5181);
and U7117 (N_7117,N_5590,N_5666);
xor U7118 (N_7118,N_5395,N_5510);
or U7119 (N_7119,N_5873,N_5220);
and U7120 (N_7120,N_4741,N_5108);
or U7121 (N_7121,N_5647,N_5577);
nand U7122 (N_7122,N_4652,N_4680);
nor U7123 (N_7123,N_5017,N_5285);
nand U7124 (N_7124,N_5165,N_4638);
or U7125 (N_7125,N_5807,N_4725);
nor U7126 (N_7126,N_5177,N_5351);
nand U7127 (N_7127,N_5219,N_4844);
nand U7128 (N_7128,N_4840,N_5624);
nor U7129 (N_7129,N_4933,N_5582);
nand U7130 (N_7130,N_5817,N_5447);
nor U7131 (N_7131,N_5235,N_5356);
nor U7132 (N_7132,N_4636,N_5652);
or U7133 (N_7133,N_5896,N_5349);
and U7134 (N_7134,N_5872,N_4527);
or U7135 (N_7135,N_5575,N_5364);
nor U7136 (N_7136,N_5359,N_5032);
nand U7137 (N_7137,N_4685,N_4743);
nor U7138 (N_7138,N_5050,N_5058);
nor U7139 (N_7139,N_5422,N_5749);
nor U7140 (N_7140,N_4997,N_5970);
nand U7141 (N_7141,N_5187,N_5159);
or U7142 (N_7142,N_5697,N_4556);
nor U7143 (N_7143,N_5025,N_5932);
xnor U7144 (N_7144,N_5528,N_4790);
nor U7145 (N_7145,N_5066,N_5896);
nor U7146 (N_7146,N_5858,N_5129);
xnor U7147 (N_7147,N_5805,N_5228);
and U7148 (N_7148,N_5942,N_4848);
xnor U7149 (N_7149,N_4559,N_5076);
nand U7150 (N_7150,N_5015,N_5643);
nand U7151 (N_7151,N_5740,N_5367);
or U7152 (N_7152,N_4739,N_5922);
or U7153 (N_7153,N_4883,N_5410);
and U7154 (N_7154,N_4544,N_5970);
nor U7155 (N_7155,N_5358,N_4599);
xor U7156 (N_7156,N_5259,N_4644);
or U7157 (N_7157,N_5771,N_4544);
and U7158 (N_7158,N_5565,N_5593);
nor U7159 (N_7159,N_4578,N_5120);
nor U7160 (N_7160,N_4542,N_4736);
xor U7161 (N_7161,N_5288,N_5377);
or U7162 (N_7162,N_4727,N_4748);
nor U7163 (N_7163,N_5973,N_5315);
or U7164 (N_7164,N_5084,N_4593);
nor U7165 (N_7165,N_5177,N_5951);
nor U7166 (N_7166,N_5999,N_5814);
or U7167 (N_7167,N_4953,N_5431);
or U7168 (N_7168,N_5341,N_4872);
and U7169 (N_7169,N_5658,N_5719);
xnor U7170 (N_7170,N_5307,N_5776);
nor U7171 (N_7171,N_4932,N_4945);
nor U7172 (N_7172,N_5820,N_5765);
nor U7173 (N_7173,N_5829,N_5557);
nor U7174 (N_7174,N_5752,N_5727);
or U7175 (N_7175,N_5869,N_5212);
nand U7176 (N_7176,N_5155,N_5712);
nand U7177 (N_7177,N_5428,N_5018);
nand U7178 (N_7178,N_4749,N_4532);
and U7179 (N_7179,N_5014,N_5131);
nor U7180 (N_7180,N_5886,N_5298);
nand U7181 (N_7181,N_5716,N_4924);
nor U7182 (N_7182,N_5673,N_5773);
xnor U7183 (N_7183,N_4844,N_5994);
xnor U7184 (N_7184,N_5588,N_5635);
and U7185 (N_7185,N_5760,N_4544);
nand U7186 (N_7186,N_4763,N_5510);
nand U7187 (N_7187,N_5626,N_4864);
nor U7188 (N_7188,N_5316,N_5882);
and U7189 (N_7189,N_5044,N_5574);
and U7190 (N_7190,N_4620,N_5423);
and U7191 (N_7191,N_4845,N_5177);
nor U7192 (N_7192,N_4973,N_4737);
nor U7193 (N_7193,N_4714,N_4878);
xnor U7194 (N_7194,N_5874,N_5734);
nor U7195 (N_7195,N_5255,N_4538);
xor U7196 (N_7196,N_5830,N_4671);
nand U7197 (N_7197,N_5348,N_5321);
nor U7198 (N_7198,N_4858,N_5182);
nand U7199 (N_7199,N_5368,N_5169);
nand U7200 (N_7200,N_5835,N_5943);
and U7201 (N_7201,N_5163,N_5162);
nand U7202 (N_7202,N_4990,N_5809);
and U7203 (N_7203,N_4561,N_5723);
nand U7204 (N_7204,N_5252,N_5432);
or U7205 (N_7205,N_4653,N_5569);
xnor U7206 (N_7206,N_4607,N_5065);
nand U7207 (N_7207,N_4608,N_5865);
and U7208 (N_7208,N_5546,N_5867);
or U7209 (N_7209,N_5033,N_5593);
or U7210 (N_7210,N_5789,N_5192);
nand U7211 (N_7211,N_5562,N_5793);
and U7212 (N_7212,N_4700,N_5680);
nand U7213 (N_7213,N_5176,N_5120);
nor U7214 (N_7214,N_5088,N_5854);
nor U7215 (N_7215,N_4748,N_5440);
nor U7216 (N_7216,N_5580,N_5850);
xor U7217 (N_7217,N_4601,N_5791);
nor U7218 (N_7218,N_4557,N_4731);
nor U7219 (N_7219,N_5681,N_4628);
and U7220 (N_7220,N_5138,N_5351);
and U7221 (N_7221,N_5557,N_5082);
nand U7222 (N_7222,N_5792,N_5098);
and U7223 (N_7223,N_5697,N_5289);
nand U7224 (N_7224,N_4705,N_4768);
and U7225 (N_7225,N_5472,N_4645);
and U7226 (N_7226,N_5471,N_5551);
nor U7227 (N_7227,N_4545,N_5047);
or U7228 (N_7228,N_5226,N_5959);
nand U7229 (N_7229,N_5039,N_5907);
or U7230 (N_7230,N_5823,N_5262);
nor U7231 (N_7231,N_5266,N_4781);
and U7232 (N_7232,N_4559,N_5455);
or U7233 (N_7233,N_4737,N_4646);
nor U7234 (N_7234,N_4658,N_5604);
nor U7235 (N_7235,N_4689,N_4954);
and U7236 (N_7236,N_5453,N_4750);
and U7237 (N_7237,N_5399,N_5729);
and U7238 (N_7238,N_4607,N_5130);
or U7239 (N_7239,N_5263,N_4908);
or U7240 (N_7240,N_5805,N_5163);
or U7241 (N_7241,N_5434,N_4654);
nor U7242 (N_7242,N_5026,N_5113);
nor U7243 (N_7243,N_4829,N_4855);
and U7244 (N_7244,N_4578,N_5800);
or U7245 (N_7245,N_4731,N_4962);
nand U7246 (N_7246,N_5671,N_5159);
and U7247 (N_7247,N_4683,N_4672);
nand U7248 (N_7248,N_5245,N_4765);
nor U7249 (N_7249,N_5761,N_4532);
or U7250 (N_7250,N_4902,N_5238);
and U7251 (N_7251,N_5635,N_5482);
xor U7252 (N_7252,N_5082,N_5230);
and U7253 (N_7253,N_5460,N_5880);
or U7254 (N_7254,N_5517,N_5059);
nand U7255 (N_7255,N_5784,N_5425);
or U7256 (N_7256,N_5781,N_5066);
nand U7257 (N_7257,N_5537,N_5837);
and U7258 (N_7258,N_5893,N_5159);
nand U7259 (N_7259,N_5890,N_5035);
nand U7260 (N_7260,N_5921,N_5595);
and U7261 (N_7261,N_5601,N_4580);
xnor U7262 (N_7262,N_5329,N_4903);
or U7263 (N_7263,N_5304,N_5756);
and U7264 (N_7264,N_5427,N_4696);
or U7265 (N_7265,N_4715,N_4534);
xor U7266 (N_7266,N_5237,N_5751);
and U7267 (N_7267,N_4894,N_5993);
nand U7268 (N_7268,N_4646,N_4687);
nand U7269 (N_7269,N_5099,N_5572);
nor U7270 (N_7270,N_5056,N_4874);
and U7271 (N_7271,N_4967,N_4658);
nor U7272 (N_7272,N_5012,N_4872);
or U7273 (N_7273,N_5545,N_5229);
nand U7274 (N_7274,N_4713,N_5517);
xnor U7275 (N_7275,N_4539,N_5438);
or U7276 (N_7276,N_4587,N_4838);
and U7277 (N_7277,N_5216,N_5993);
nor U7278 (N_7278,N_5722,N_5850);
xnor U7279 (N_7279,N_5022,N_5259);
nor U7280 (N_7280,N_5888,N_4856);
nor U7281 (N_7281,N_4780,N_5049);
or U7282 (N_7282,N_5818,N_4814);
and U7283 (N_7283,N_4747,N_4816);
or U7284 (N_7284,N_5776,N_5424);
nand U7285 (N_7285,N_5798,N_5265);
nor U7286 (N_7286,N_5794,N_5597);
or U7287 (N_7287,N_4898,N_4760);
nor U7288 (N_7288,N_4931,N_5688);
nand U7289 (N_7289,N_4960,N_5593);
nand U7290 (N_7290,N_5941,N_5886);
or U7291 (N_7291,N_5141,N_5284);
xnor U7292 (N_7292,N_5915,N_5549);
nor U7293 (N_7293,N_5980,N_5254);
and U7294 (N_7294,N_5994,N_5944);
and U7295 (N_7295,N_5644,N_5436);
nor U7296 (N_7296,N_5088,N_4663);
nand U7297 (N_7297,N_5177,N_5767);
and U7298 (N_7298,N_5923,N_5938);
nor U7299 (N_7299,N_5103,N_4515);
and U7300 (N_7300,N_5011,N_5084);
or U7301 (N_7301,N_5514,N_4761);
nand U7302 (N_7302,N_4829,N_5322);
and U7303 (N_7303,N_5144,N_4776);
and U7304 (N_7304,N_4602,N_5482);
or U7305 (N_7305,N_5923,N_5221);
or U7306 (N_7306,N_5264,N_5651);
or U7307 (N_7307,N_5611,N_5594);
nand U7308 (N_7308,N_5325,N_5214);
and U7309 (N_7309,N_5249,N_5234);
or U7310 (N_7310,N_5138,N_5732);
nor U7311 (N_7311,N_5890,N_5698);
nand U7312 (N_7312,N_4562,N_5917);
and U7313 (N_7313,N_4653,N_4588);
xor U7314 (N_7314,N_5521,N_4634);
and U7315 (N_7315,N_5450,N_5472);
nor U7316 (N_7316,N_5162,N_5243);
nand U7317 (N_7317,N_4828,N_5232);
nand U7318 (N_7318,N_5860,N_4589);
or U7319 (N_7319,N_4844,N_5313);
nor U7320 (N_7320,N_5685,N_4553);
xor U7321 (N_7321,N_5717,N_5729);
nor U7322 (N_7322,N_5312,N_4932);
or U7323 (N_7323,N_5931,N_5266);
nor U7324 (N_7324,N_5177,N_5222);
nand U7325 (N_7325,N_4780,N_5213);
and U7326 (N_7326,N_4985,N_5155);
and U7327 (N_7327,N_4543,N_5413);
and U7328 (N_7328,N_5039,N_5297);
nor U7329 (N_7329,N_5465,N_5143);
or U7330 (N_7330,N_4675,N_5027);
nand U7331 (N_7331,N_5213,N_5533);
or U7332 (N_7332,N_4707,N_4936);
and U7333 (N_7333,N_5444,N_5256);
and U7334 (N_7334,N_5245,N_4629);
or U7335 (N_7335,N_5455,N_5940);
or U7336 (N_7336,N_4564,N_5979);
or U7337 (N_7337,N_5639,N_4599);
or U7338 (N_7338,N_5830,N_5829);
or U7339 (N_7339,N_4760,N_5793);
nand U7340 (N_7340,N_5717,N_4565);
nor U7341 (N_7341,N_5530,N_4804);
and U7342 (N_7342,N_5111,N_4556);
or U7343 (N_7343,N_5023,N_5243);
or U7344 (N_7344,N_5221,N_5220);
or U7345 (N_7345,N_5689,N_5017);
nand U7346 (N_7346,N_4512,N_5018);
and U7347 (N_7347,N_5910,N_5395);
nor U7348 (N_7348,N_5178,N_5955);
or U7349 (N_7349,N_5661,N_5471);
or U7350 (N_7350,N_4876,N_5243);
xor U7351 (N_7351,N_4622,N_5983);
nor U7352 (N_7352,N_5552,N_5833);
nand U7353 (N_7353,N_4974,N_4935);
or U7354 (N_7354,N_5232,N_5902);
and U7355 (N_7355,N_4540,N_5045);
or U7356 (N_7356,N_4606,N_5497);
nand U7357 (N_7357,N_5939,N_4769);
nor U7358 (N_7358,N_5580,N_4978);
nand U7359 (N_7359,N_5041,N_5779);
nor U7360 (N_7360,N_5418,N_5954);
and U7361 (N_7361,N_5982,N_4526);
or U7362 (N_7362,N_5075,N_5239);
nand U7363 (N_7363,N_5542,N_5452);
nand U7364 (N_7364,N_5731,N_5481);
or U7365 (N_7365,N_5934,N_4748);
and U7366 (N_7366,N_5742,N_5054);
nand U7367 (N_7367,N_5810,N_5971);
nor U7368 (N_7368,N_5817,N_5633);
nand U7369 (N_7369,N_5969,N_4601);
nand U7370 (N_7370,N_4577,N_5762);
nor U7371 (N_7371,N_4596,N_5927);
xor U7372 (N_7372,N_5075,N_5397);
nor U7373 (N_7373,N_5068,N_5870);
or U7374 (N_7374,N_4822,N_5606);
nand U7375 (N_7375,N_5110,N_5095);
or U7376 (N_7376,N_5383,N_4989);
nor U7377 (N_7377,N_4560,N_5972);
nor U7378 (N_7378,N_5252,N_5450);
or U7379 (N_7379,N_4569,N_5029);
nor U7380 (N_7380,N_5187,N_5270);
nor U7381 (N_7381,N_4558,N_4997);
xnor U7382 (N_7382,N_5984,N_5198);
nor U7383 (N_7383,N_5392,N_5484);
or U7384 (N_7384,N_5048,N_4580);
nand U7385 (N_7385,N_5235,N_4595);
or U7386 (N_7386,N_4568,N_5618);
nor U7387 (N_7387,N_4521,N_5731);
nand U7388 (N_7388,N_5879,N_5852);
or U7389 (N_7389,N_5472,N_4754);
and U7390 (N_7390,N_4570,N_4660);
xnor U7391 (N_7391,N_5766,N_5026);
or U7392 (N_7392,N_5324,N_5503);
nor U7393 (N_7393,N_5244,N_4712);
nand U7394 (N_7394,N_4575,N_5482);
nand U7395 (N_7395,N_4983,N_4716);
or U7396 (N_7396,N_5458,N_4813);
and U7397 (N_7397,N_5530,N_5419);
xnor U7398 (N_7398,N_5524,N_4904);
and U7399 (N_7399,N_4864,N_4514);
nor U7400 (N_7400,N_5115,N_5283);
and U7401 (N_7401,N_5901,N_5846);
and U7402 (N_7402,N_5070,N_5590);
xnor U7403 (N_7403,N_5948,N_4683);
and U7404 (N_7404,N_5973,N_5348);
xor U7405 (N_7405,N_4952,N_5098);
and U7406 (N_7406,N_5088,N_5229);
xnor U7407 (N_7407,N_5959,N_4796);
and U7408 (N_7408,N_5346,N_5255);
nor U7409 (N_7409,N_5446,N_4791);
and U7410 (N_7410,N_5437,N_4898);
and U7411 (N_7411,N_5879,N_5772);
nand U7412 (N_7412,N_5124,N_5422);
and U7413 (N_7413,N_5923,N_5717);
or U7414 (N_7414,N_4990,N_5674);
nand U7415 (N_7415,N_5066,N_4733);
or U7416 (N_7416,N_5908,N_5997);
and U7417 (N_7417,N_4872,N_4508);
or U7418 (N_7418,N_4676,N_5720);
nand U7419 (N_7419,N_5431,N_5239);
and U7420 (N_7420,N_5741,N_4929);
nor U7421 (N_7421,N_5492,N_5176);
nand U7422 (N_7422,N_5783,N_5811);
and U7423 (N_7423,N_5962,N_5028);
nor U7424 (N_7424,N_5428,N_5296);
nand U7425 (N_7425,N_5149,N_5311);
or U7426 (N_7426,N_4765,N_5047);
nor U7427 (N_7427,N_5480,N_5356);
nor U7428 (N_7428,N_5402,N_5642);
nor U7429 (N_7429,N_5140,N_5885);
xor U7430 (N_7430,N_4578,N_4631);
nand U7431 (N_7431,N_5702,N_5613);
nand U7432 (N_7432,N_4740,N_5618);
nand U7433 (N_7433,N_4753,N_5650);
xnor U7434 (N_7434,N_5827,N_5402);
and U7435 (N_7435,N_4739,N_4593);
nand U7436 (N_7436,N_5656,N_5210);
nand U7437 (N_7437,N_4816,N_5997);
or U7438 (N_7438,N_5058,N_5026);
xor U7439 (N_7439,N_4836,N_5374);
or U7440 (N_7440,N_5041,N_5265);
and U7441 (N_7441,N_5101,N_5771);
nand U7442 (N_7442,N_4603,N_5036);
or U7443 (N_7443,N_5608,N_4984);
or U7444 (N_7444,N_5521,N_5177);
nor U7445 (N_7445,N_5360,N_5390);
nand U7446 (N_7446,N_5389,N_5916);
and U7447 (N_7447,N_5038,N_5911);
or U7448 (N_7448,N_4621,N_4656);
and U7449 (N_7449,N_5090,N_4540);
or U7450 (N_7450,N_4609,N_5650);
or U7451 (N_7451,N_4672,N_5486);
xor U7452 (N_7452,N_4562,N_5108);
xor U7453 (N_7453,N_4810,N_4613);
nand U7454 (N_7454,N_4986,N_5924);
or U7455 (N_7455,N_5721,N_5383);
and U7456 (N_7456,N_5226,N_5107);
nor U7457 (N_7457,N_5138,N_5137);
nor U7458 (N_7458,N_5191,N_5303);
nor U7459 (N_7459,N_4560,N_4527);
xor U7460 (N_7460,N_4880,N_4837);
and U7461 (N_7461,N_4923,N_5182);
and U7462 (N_7462,N_4506,N_5006);
nor U7463 (N_7463,N_5027,N_4550);
nand U7464 (N_7464,N_5356,N_5257);
nand U7465 (N_7465,N_5840,N_5876);
nand U7466 (N_7466,N_4786,N_5504);
and U7467 (N_7467,N_4823,N_4744);
nand U7468 (N_7468,N_5818,N_4882);
nand U7469 (N_7469,N_5950,N_4943);
nor U7470 (N_7470,N_5438,N_5685);
xor U7471 (N_7471,N_5556,N_5891);
nand U7472 (N_7472,N_4578,N_5828);
nand U7473 (N_7473,N_5437,N_4600);
or U7474 (N_7474,N_5742,N_5837);
nand U7475 (N_7475,N_5503,N_5853);
and U7476 (N_7476,N_5906,N_5311);
and U7477 (N_7477,N_5762,N_5832);
or U7478 (N_7478,N_5558,N_5074);
and U7479 (N_7479,N_5492,N_5547);
and U7480 (N_7480,N_5945,N_5315);
and U7481 (N_7481,N_5105,N_5299);
or U7482 (N_7482,N_4616,N_5011);
or U7483 (N_7483,N_4985,N_4525);
and U7484 (N_7484,N_5483,N_5292);
and U7485 (N_7485,N_4829,N_4650);
nand U7486 (N_7486,N_4632,N_5423);
nand U7487 (N_7487,N_4934,N_5860);
and U7488 (N_7488,N_4963,N_5823);
and U7489 (N_7489,N_5139,N_5494);
and U7490 (N_7490,N_5086,N_5751);
or U7491 (N_7491,N_5937,N_5845);
nor U7492 (N_7492,N_5320,N_5100);
nor U7493 (N_7493,N_5303,N_4525);
and U7494 (N_7494,N_5163,N_4513);
nor U7495 (N_7495,N_4651,N_4531);
nor U7496 (N_7496,N_5287,N_4617);
or U7497 (N_7497,N_4527,N_5501);
nor U7498 (N_7498,N_5534,N_5830);
nor U7499 (N_7499,N_5861,N_5882);
and U7500 (N_7500,N_6659,N_6350);
and U7501 (N_7501,N_6904,N_6037);
or U7502 (N_7502,N_6406,N_7007);
nor U7503 (N_7503,N_6298,N_6728);
and U7504 (N_7504,N_7334,N_6119);
nand U7505 (N_7505,N_6690,N_6631);
xnor U7506 (N_7506,N_6885,N_6347);
and U7507 (N_7507,N_7248,N_7461);
xnor U7508 (N_7508,N_6460,N_6537);
nand U7509 (N_7509,N_7087,N_6787);
nor U7510 (N_7510,N_6349,N_6292);
nand U7511 (N_7511,N_6984,N_7059);
or U7512 (N_7512,N_6179,N_6687);
nor U7513 (N_7513,N_7285,N_7206);
nor U7514 (N_7514,N_7102,N_7217);
nand U7515 (N_7515,N_6555,N_6838);
nand U7516 (N_7516,N_6772,N_6473);
nand U7517 (N_7517,N_7402,N_6522);
nand U7518 (N_7518,N_7005,N_6265);
nand U7519 (N_7519,N_6260,N_6282);
or U7520 (N_7520,N_7166,N_6870);
nor U7521 (N_7521,N_6222,N_6210);
xnor U7522 (N_7522,N_7481,N_6969);
nor U7523 (N_7523,N_6756,N_6987);
nand U7524 (N_7524,N_6068,N_7260);
xnor U7525 (N_7525,N_6214,N_6344);
and U7526 (N_7526,N_7386,N_7405);
xor U7527 (N_7527,N_6039,N_6516);
nor U7528 (N_7528,N_6193,N_6730);
nand U7529 (N_7529,N_6890,N_7312);
and U7530 (N_7530,N_6353,N_6683);
and U7531 (N_7531,N_7347,N_6285);
nand U7532 (N_7532,N_6189,N_6793);
and U7533 (N_7533,N_7300,N_6733);
and U7534 (N_7534,N_7276,N_6698);
nand U7535 (N_7535,N_6953,N_6767);
nor U7536 (N_7536,N_6238,N_7235);
xnor U7537 (N_7537,N_6174,N_7144);
nand U7538 (N_7538,N_6843,N_7354);
or U7539 (N_7539,N_6655,N_6268);
nor U7540 (N_7540,N_6212,N_7213);
and U7541 (N_7541,N_6942,N_7306);
nor U7542 (N_7542,N_6702,N_6519);
and U7543 (N_7543,N_6610,N_7167);
and U7544 (N_7544,N_6708,N_7198);
nand U7545 (N_7545,N_7298,N_7240);
xnor U7546 (N_7546,N_6133,N_7480);
nand U7547 (N_7547,N_6288,N_6726);
nor U7548 (N_7548,N_6883,N_7370);
nand U7549 (N_7549,N_6939,N_6593);
and U7550 (N_7550,N_6632,N_7228);
and U7551 (N_7551,N_6707,N_6910);
and U7552 (N_7552,N_7001,N_6856);
nand U7553 (N_7553,N_6439,N_7255);
and U7554 (N_7554,N_7262,N_6805);
nor U7555 (N_7555,N_6889,N_6678);
or U7556 (N_7556,N_6499,N_6996);
or U7557 (N_7557,N_6586,N_6542);
or U7558 (N_7558,N_7249,N_6446);
nor U7559 (N_7559,N_6018,N_6782);
and U7560 (N_7560,N_6008,N_6062);
or U7561 (N_7561,N_7449,N_7353);
and U7562 (N_7562,N_6675,N_7436);
and U7563 (N_7563,N_6315,N_6528);
and U7564 (N_7564,N_7281,N_7131);
nor U7565 (N_7565,N_7318,N_6629);
nor U7566 (N_7566,N_6129,N_7054);
xnor U7567 (N_7567,N_6403,N_6228);
nand U7568 (N_7568,N_7315,N_6382);
and U7569 (N_7569,N_7483,N_6845);
or U7570 (N_7570,N_6511,N_6498);
nand U7571 (N_7571,N_6148,N_7208);
nor U7572 (N_7572,N_6633,N_6842);
xor U7573 (N_7573,N_7147,N_6819);
nor U7574 (N_7574,N_7311,N_6386);
nand U7575 (N_7575,N_7134,N_6703);
and U7576 (N_7576,N_6752,N_6034);
or U7577 (N_7577,N_7159,N_6636);
nor U7578 (N_7578,N_7157,N_6035);
and U7579 (N_7579,N_6314,N_7178);
and U7580 (N_7580,N_7388,N_6251);
or U7581 (N_7581,N_6573,N_7321);
and U7582 (N_7582,N_6502,N_7137);
nor U7583 (N_7583,N_7211,N_6147);
nor U7584 (N_7584,N_7006,N_6413);
nor U7585 (N_7585,N_6991,N_6900);
nor U7586 (N_7586,N_6669,N_6024);
or U7587 (N_7587,N_7413,N_6621);
and U7588 (N_7588,N_6967,N_6640);
or U7589 (N_7589,N_6864,N_6836);
xor U7590 (N_7590,N_6426,N_6983);
or U7591 (N_7591,N_7034,N_7109);
nor U7592 (N_7592,N_6358,N_6259);
and U7593 (N_7593,N_6924,N_6012);
or U7594 (N_7594,N_6463,N_6233);
nand U7595 (N_7595,N_6619,N_7485);
and U7596 (N_7596,N_6416,N_7348);
nor U7597 (N_7597,N_6973,N_6695);
nand U7598 (N_7598,N_6146,N_6865);
nand U7599 (N_7599,N_6946,N_6982);
or U7600 (N_7600,N_6396,N_6171);
and U7601 (N_7601,N_6584,N_6764);
nand U7602 (N_7602,N_6735,N_7000);
or U7603 (N_7603,N_6213,N_7045);
nor U7604 (N_7604,N_6951,N_6327);
nor U7605 (N_7605,N_6866,N_7352);
nand U7606 (N_7606,N_6830,N_7030);
nor U7607 (N_7607,N_6393,N_6073);
and U7608 (N_7608,N_6930,N_6097);
or U7609 (N_7609,N_7238,N_6130);
nand U7610 (N_7610,N_7314,N_6091);
or U7611 (N_7611,N_6850,N_7146);
and U7612 (N_7612,N_6820,N_6096);
or U7613 (N_7613,N_6880,N_7075);
or U7614 (N_7614,N_6775,N_6716);
nor U7615 (N_7615,N_6256,N_6369);
or U7616 (N_7616,N_6071,N_6705);
and U7617 (N_7617,N_6668,N_7451);
nor U7618 (N_7618,N_7094,N_7164);
nor U7619 (N_7619,N_6791,N_6602);
nand U7620 (N_7620,N_6624,N_6291);
and U7621 (N_7621,N_6115,N_6554);
nor U7622 (N_7622,N_6231,N_6140);
and U7623 (N_7623,N_7128,N_7371);
nor U7624 (N_7624,N_7303,N_6874);
nor U7625 (N_7625,N_6616,N_6790);
or U7626 (N_7626,N_7310,N_6289);
nand U7627 (N_7627,N_6230,N_6712);
nor U7628 (N_7628,N_6194,N_6411);
or U7629 (N_7629,N_6437,N_7028);
and U7630 (N_7630,N_6641,N_6419);
or U7631 (N_7631,N_6056,N_7283);
or U7632 (N_7632,N_6732,N_7245);
or U7633 (N_7633,N_6400,N_6952);
nand U7634 (N_7634,N_6868,N_6941);
nand U7635 (N_7635,N_7437,N_7170);
and U7636 (N_7636,N_7069,N_6495);
nor U7637 (N_7637,N_6257,N_6753);
nor U7638 (N_7638,N_6267,N_6886);
and U7639 (N_7639,N_6004,N_7287);
and U7640 (N_7640,N_7129,N_7078);
or U7641 (N_7641,N_6184,N_6185);
and U7642 (N_7642,N_6164,N_6774);
or U7643 (N_7643,N_7292,N_6319);
and U7644 (N_7644,N_6679,N_6862);
nand U7645 (N_7645,N_6673,N_7187);
or U7646 (N_7646,N_6553,N_6442);
nor U7647 (N_7647,N_7491,N_6911);
and U7648 (N_7648,N_6970,N_7291);
xnor U7649 (N_7649,N_6438,N_6660);
or U7650 (N_7650,N_6318,N_7191);
nor U7651 (N_7651,N_6622,N_6682);
xnor U7652 (N_7652,N_7038,N_7061);
nor U7653 (N_7653,N_6266,N_7359);
nor U7654 (N_7654,N_6977,N_6643);
nor U7655 (N_7655,N_7395,N_6151);
or U7656 (N_7656,N_6652,N_6468);
and U7657 (N_7657,N_6141,N_6670);
nor U7658 (N_7658,N_6667,N_6860);
nor U7659 (N_7659,N_6645,N_7376);
nand U7660 (N_7660,N_6944,N_6248);
xnor U7661 (N_7661,N_6763,N_6398);
xor U7662 (N_7662,N_6480,N_7203);
nand U7663 (N_7663,N_7339,N_6697);
xor U7664 (N_7664,N_6059,N_6879);
or U7665 (N_7665,N_7080,N_7233);
nor U7666 (N_7666,N_7083,N_6407);
and U7667 (N_7667,N_7017,N_6015);
or U7668 (N_7668,N_6795,N_6055);
nor U7669 (N_7669,N_6471,N_7041);
nor U7670 (N_7670,N_7067,N_6425);
nor U7671 (N_7671,N_6383,N_7169);
nand U7672 (N_7672,N_6773,N_6299);
nand U7673 (N_7673,N_6239,N_6000);
and U7674 (N_7674,N_6453,N_6720);
or U7675 (N_7675,N_6599,N_6340);
nand U7676 (N_7676,N_6770,N_6160);
or U7677 (N_7677,N_6196,N_6409);
and U7678 (N_7678,N_6503,N_7053);
nand U7679 (N_7679,N_7207,N_7122);
nand U7680 (N_7680,N_6558,N_6572);
and U7681 (N_7681,N_6302,N_7390);
nand U7682 (N_7682,N_6907,N_6509);
or U7683 (N_7683,N_7264,N_6966);
and U7684 (N_7684,N_6156,N_7301);
nand U7685 (N_7685,N_6132,N_7358);
nand U7686 (N_7686,N_6143,N_6308);
or U7687 (N_7687,N_7002,N_6075);
nand U7688 (N_7688,N_7297,N_6412);
nor U7689 (N_7689,N_6065,N_6796);
and U7690 (N_7690,N_6818,N_7200);
nand U7691 (N_7691,N_7106,N_6591);
and U7692 (N_7692,N_6053,N_7117);
nor U7693 (N_7693,N_6567,N_6104);
and U7694 (N_7694,N_6069,N_6543);
nor U7695 (N_7695,N_6656,N_7100);
nand U7696 (N_7696,N_6354,N_7060);
and U7697 (N_7697,N_6116,N_6826);
nand U7698 (N_7698,N_6010,N_6063);
nand U7699 (N_7699,N_6792,N_6109);
nand U7700 (N_7700,N_7148,N_6423);
and U7701 (N_7701,N_6410,N_6613);
and U7702 (N_7702,N_6925,N_6825);
and U7703 (N_7703,N_7456,N_6022);
and U7704 (N_7704,N_7445,N_7341);
or U7705 (N_7705,N_7142,N_6514);
nor U7706 (N_7706,N_6481,N_7495);
nor U7707 (N_7707,N_6241,N_7332);
and U7708 (N_7708,N_7265,N_6121);
and U7709 (N_7709,N_6281,N_6070);
or U7710 (N_7710,N_6013,N_7324);
or U7711 (N_7711,N_6727,N_6262);
nand U7712 (N_7712,N_6589,N_7139);
xnor U7713 (N_7713,N_7490,N_7153);
nand U7714 (N_7714,N_6565,N_6131);
nor U7715 (N_7715,N_6313,N_6084);
and U7716 (N_7716,N_7056,N_6661);
nor U7717 (N_7717,N_7120,N_7330);
nand U7718 (N_7718,N_7013,N_6397);
xor U7719 (N_7719,N_6215,N_6334);
nor U7720 (N_7720,N_6863,N_6603);
and U7721 (N_7721,N_6280,N_7021);
or U7722 (N_7722,N_7032,N_6074);
nand U7723 (N_7723,N_7176,N_6666);
and U7724 (N_7724,N_6249,N_7079);
xnor U7725 (N_7725,N_6746,N_6051);
or U7726 (N_7726,N_6723,N_7236);
and U7727 (N_7727,N_6016,N_6744);
nor U7728 (N_7728,N_6391,N_7319);
nor U7729 (N_7729,N_7362,N_6488);
nand U7730 (N_7730,N_6026,N_7464);
nand U7731 (N_7731,N_6149,N_6283);
nand U7732 (N_7732,N_7210,N_7247);
nand U7733 (N_7733,N_7114,N_6336);
nor U7734 (N_7734,N_6855,N_6323);
and U7735 (N_7735,N_6803,N_6837);
and U7736 (N_7736,N_6443,N_6717);
nor U7737 (N_7737,N_6054,N_7316);
and U7738 (N_7738,N_6125,N_6914);
and U7739 (N_7739,N_6303,N_6992);
nand U7740 (N_7740,N_7473,N_7466);
nand U7741 (N_7741,N_6470,N_6552);
and U7742 (N_7742,N_6300,N_6722);
nand U7743 (N_7743,N_7244,N_6680);
nor U7744 (N_7744,N_6548,N_6408);
nor U7745 (N_7745,N_6152,N_7073);
nand U7746 (N_7746,N_6748,N_6533);
nand U7747 (N_7747,N_7047,N_6061);
or U7748 (N_7748,N_6609,N_6541);
or U7749 (N_7749,N_6990,N_6380);
nor U7750 (N_7750,N_6274,N_6840);
and U7751 (N_7751,N_6901,N_6272);
and U7752 (N_7752,N_6896,N_6144);
or U7753 (N_7753,N_7486,N_6330);
or U7754 (N_7754,N_6287,N_7482);
and U7755 (N_7755,N_6738,N_6102);
nand U7756 (N_7756,N_7216,N_6346);
and U7757 (N_7757,N_6405,N_7411);
nand U7758 (N_7758,N_6854,N_7290);
nor U7759 (N_7759,N_7138,N_6145);
nand U7760 (N_7760,N_6508,N_7192);
nand U7761 (N_7761,N_6501,N_7037);
nor U7762 (N_7762,N_6486,N_6235);
and U7763 (N_7763,N_6985,N_6771);
nand U7764 (N_7764,N_6867,N_6312);
xor U7765 (N_7765,N_7331,N_7392);
or U7766 (N_7766,N_7467,N_7003);
or U7767 (N_7767,N_6878,N_6958);
and U7768 (N_7768,N_7010,N_7031);
nor U7769 (N_7769,N_7065,N_6042);
or U7770 (N_7770,N_6120,N_6978);
or U7771 (N_7771,N_6583,N_6596);
and U7772 (N_7772,N_7323,N_6549);
and U7773 (N_7773,N_7012,N_7051);
and U7774 (N_7774,N_6093,N_6768);
or U7775 (N_7775,N_6033,N_6049);
nand U7776 (N_7776,N_7123,N_6653);
xor U7777 (N_7777,N_6812,N_6741);
or U7778 (N_7778,N_7417,N_6557);
and U7779 (N_7779,N_6276,N_6827);
and U7780 (N_7780,N_7035,N_6253);
nand U7781 (N_7781,N_7320,N_6778);
nor U7782 (N_7782,N_7251,N_6066);
or U7783 (N_7783,N_6515,N_6628);
or U7784 (N_7784,N_6875,N_6113);
and U7785 (N_7785,N_6484,N_7072);
nand U7786 (N_7786,N_7181,N_6454);
and U7787 (N_7787,N_6833,N_6255);
nand U7788 (N_7788,N_6536,N_7342);
nand U7789 (N_7789,N_6072,N_7427);
or U7790 (N_7790,N_7416,N_7459);
and U7791 (N_7791,N_6535,N_6713);
nor U7792 (N_7792,N_6388,N_7223);
or U7793 (N_7793,N_6649,N_6821);
nor U7794 (N_7794,N_6112,N_6009);
xor U7795 (N_7795,N_6547,N_6968);
and U7796 (N_7796,N_6003,N_6813);
and U7797 (N_7797,N_7071,N_6834);
nand U7798 (N_7798,N_7355,N_6903);
nor U7799 (N_7799,N_6701,N_6871);
nor U7800 (N_7800,N_6036,N_7136);
nor U7801 (N_7801,N_7068,N_7399);
nand U7802 (N_7802,N_6817,N_7284);
and U7803 (N_7803,N_6433,N_6320);
and U7804 (N_7804,N_6402,N_7112);
nor U7805 (N_7805,N_6365,N_6032);
or U7806 (N_7806,N_6273,N_6451);
nor U7807 (N_7807,N_7452,N_7344);
nor U7808 (N_7808,N_6316,N_7442);
xor U7809 (N_7809,N_6081,N_7337);
nor U7810 (N_7810,N_7175,N_6575);
or U7811 (N_7811,N_7077,N_7243);
or U7812 (N_7812,N_7024,N_7270);
and U7813 (N_7813,N_6157,N_6176);
xor U7814 (N_7814,N_6894,N_6309);
xor U7815 (N_7815,N_6923,N_7018);
nand U7816 (N_7816,N_7462,N_6046);
nor U7817 (N_7817,N_6326,N_7108);
and U7818 (N_7818,N_6906,N_7431);
and U7819 (N_7819,N_6560,N_7225);
and U7820 (N_7820,N_6861,N_6788);
and U7821 (N_7821,N_6154,N_7272);
nand U7822 (N_7822,N_6475,N_7040);
and U7823 (N_7823,N_6296,N_6814);
nor U7824 (N_7824,N_6956,N_6579);
and U7825 (N_7825,N_6852,N_7149);
xor U7826 (N_7826,N_6935,N_7434);
or U7827 (N_7827,N_6674,N_6520);
nor U7828 (N_7828,N_6810,N_6435);
or U7829 (N_7829,N_7161,N_6464);
nor U7830 (N_7830,N_7299,N_6891);
nand U7831 (N_7831,N_7202,N_6279);
xnor U7832 (N_7832,N_7420,N_6823);
or U7833 (N_7833,N_6355,N_6496);
and U7834 (N_7834,N_6092,N_6578);
or U7835 (N_7835,N_6415,N_6479);
or U7836 (N_7836,N_7327,N_6356);
nor U7837 (N_7837,N_6306,N_7224);
or U7838 (N_7838,N_6998,N_7271);
nand U7839 (N_7839,N_6506,N_7458);
xnor U7840 (N_7840,N_7412,N_7160);
and U7841 (N_7841,N_6457,N_6363);
nor U7842 (N_7842,N_6934,N_7326);
nand U7843 (N_7843,N_6218,N_7093);
or U7844 (N_7844,N_6887,N_6582);
xor U7845 (N_7845,N_7400,N_6884);
xor U7846 (N_7846,N_7096,N_7193);
nor U7847 (N_7847,N_6474,N_6339);
nand U7848 (N_7848,N_7130,N_7092);
nor U7849 (N_7849,N_6317,N_7082);
or U7850 (N_7850,N_6098,N_6873);
or U7851 (N_7851,N_6373,N_7429);
xnor U7852 (N_7852,N_6117,N_6384);
and U7853 (N_7853,N_6783,N_7309);
nor U7854 (N_7854,N_6478,N_6006);
or U7855 (N_7855,N_7277,N_6993);
nor U7856 (N_7856,N_6794,N_6580);
xnor U7857 (N_7857,N_6362,N_6044);
nor U7858 (N_7858,N_6324,N_6429);
nor U7859 (N_7859,N_7089,N_6647);
nand U7860 (N_7860,N_6505,N_6374);
nor U7861 (N_7861,N_6761,N_7118);
and U7862 (N_7862,N_6740,N_7226);
xor U7863 (N_7863,N_6108,N_6600);
and U7864 (N_7864,N_6139,N_6882);
nor U7865 (N_7865,N_7457,N_6718);
or U7866 (N_7866,N_6568,N_6684);
nor U7867 (N_7867,N_6079,N_6815);
nor U7868 (N_7868,N_6762,N_7268);
or U7869 (N_7869,N_6607,N_6064);
and U7870 (N_7870,N_6448,N_7062);
nor U7871 (N_7871,N_6829,N_6858);
or U7872 (N_7872,N_7205,N_6913);
and U7873 (N_7873,N_7085,N_7340);
or U7874 (N_7874,N_6310,N_6348);
nand U7875 (N_7875,N_7286,N_6077);
nand U7876 (N_7876,N_6630,N_6472);
or U7877 (N_7877,N_6459,N_7055);
and U7878 (N_7878,N_7057,N_7345);
nor U7879 (N_7879,N_6928,N_6332);
and U7880 (N_7880,N_6811,N_6048);
nand U7881 (N_7881,N_7498,N_6938);
nor U7882 (N_7882,N_6118,N_7184);
nand U7883 (N_7883,N_6912,N_6601);
and U7884 (N_7884,N_7304,N_7052);
nand U7885 (N_7885,N_6394,N_6776);
and U7886 (N_7886,N_7282,N_7070);
or U7887 (N_7887,N_6192,N_7222);
xnor U7888 (N_7888,N_7447,N_6739);
nand U7889 (N_7889,N_7189,N_6665);
or U7890 (N_7890,N_6226,N_7237);
or U7891 (N_7891,N_6963,N_6089);
xor U7892 (N_7892,N_7433,N_6490);
and U7893 (N_7893,N_7302,N_6615);
nand U7894 (N_7894,N_6585,N_6704);
nand U7895 (N_7895,N_7165,N_6662);
nand U7896 (N_7896,N_7378,N_6657);
and U7897 (N_7897,N_6574,N_6694);
and U7898 (N_7898,N_7258,N_6975);
nand U7899 (N_7899,N_6692,N_6234);
nand U7900 (N_7900,N_7081,N_6721);
or U7901 (N_7901,N_6504,N_6205);
nor U7902 (N_7902,N_6876,N_6178);
nor U7903 (N_7903,N_6219,N_6530);
or U7904 (N_7904,N_7194,N_6550);
nor U7905 (N_7905,N_6634,N_6469);
nand U7906 (N_7906,N_6414,N_6769);
nor U7907 (N_7907,N_6808,N_6908);
nor U7908 (N_7908,N_6381,N_7158);
nor U7909 (N_7909,N_6126,N_6221);
and U7910 (N_7910,N_6807,N_6424);
and U7911 (N_7911,N_6040,N_7125);
or U7912 (N_7912,N_7441,N_7022);
and U7913 (N_7913,N_6571,N_7110);
nor U7914 (N_7914,N_7468,N_6625);
nor U7915 (N_7915,N_6007,N_6736);
or U7916 (N_7916,N_6639,N_6421);
nor U7917 (N_7917,N_7197,N_6957);
nor U7918 (N_7918,N_6789,N_6598);
and U7919 (N_7919,N_6087,N_7014);
nor U7920 (N_7920,N_6245,N_6994);
or U7921 (N_7921,N_7463,N_7489);
nand U7922 (N_7922,N_6169,N_6706);
xnor U7923 (N_7923,N_6106,N_7295);
and U7924 (N_7924,N_6019,N_6020);
and U7925 (N_7925,N_7446,N_7177);
xor U7926 (N_7926,N_6620,N_7267);
or U7927 (N_7927,N_6240,N_6745);
and U7928 (N_7928,N_6755,N_6190);
nand U7929 (N_7929,N_6989,N_6592);
and U7930 (N_7930,N_7064,N_6999);
nor U7931 (N_7931,N_7478,N_7214);
nor U7932 (N_7932,N_6798,N_7099);
nand U7933 (N_7933,N_7253,N_6691);
nand U7934 (N_7934,N_6688,N_6859);
nor U7935 (N_7935,N_6338,N_7058);
or U7936 (N_7936,N_6487,N_6569);
and U7937 (N_7937,N_6041,N_7280);
nor U7938 (N_7938,N_6931,N_7409);
nand U7939 (N_7939,N_6085,N_7492);
and U7940 (N_7940,N_6714,N_7043);
xnor U7941 (N_7941,N_6606,N_7050);
or U7942 (N_7942,N_7423,N_7336);
nor U7943 (N_7943,N_7387,N_7116);
or U7944 (N_7944,N_7313,N_7308);
nand U7945 (N_7945,N_7121,N_6321);
or U7946 (N_7946,N_6777,N_6027);
and U7947 (N_7947,N_6962,N_7044);
nand U7948 (N_7948,N_6466,N_6258);
nor U7949 (N_7949,N_6781,N_7430);
nor U7950 (N_7950,N_6638,N_6432);
nand U7951 (N_7951,N_6271,N_6784);
nor U7952 (N_7952,N_6376,N_6014);
nand U7953 (N_7953,N_7410,N_6211);
nand U7954 (N_7954,N_6595,N_7145);
or U7955 (N_7955,N_6758,N_6489);
and U7956 (N_7956,N_7186,N_6031);
and U7957 (N_7957,N_7229,N_6623);
xnor U7958 (N_7958,N_6832,N_6447);
or U7959 (N_7959,N_6370,N_7185);
nor U7960 (N_7960,N_6351,N_6650);
and U7961 (N_7961,N_6177,N_6163);
nor U7962 (N_7962,N_6759,N_7364);
nor U7963 (N_7963,N_6986,N_7168);
nand U7964 (N_7964,N_7263,N_7246);
and U7965 (N_7965,N_6043,N_6220);
nand U7966 (N_7966,N_6948,N_7046);
and U7967 (N_7967,N_7397,N_6372);
and U7968 (N_7968,N_6950,N_7036);
or U7969 (N_7969,N_6025,N_6107);
and U7970 (N_7970,N_6534,N_6809);
xnor U7971 (N_7971,N_6507,N_6430);
or U7972 (N_7972,N_6124,N_6725);
nor U7973 (N_7973,N_7425,N_6869);
and U7974 (N_7974,N_7439,N_6128);
or U7975 (N_7975,N_6750,N_6844);
nand U7976 (N_7976,N_7289,N_6513);
and U7977 (N_7977,N_6899,N_6608);
nor U7978 (N_7978,N_7418,N_6067);
and U7979 (N_7979,N_6857,N_7421);
or U7980 (N_7980,N_6252,N_6441);
and U7981 (N_7981,N_6284,N_6243);
or U7982 (N_7982,N_7151,N_6897);
nand U7983 (N_7983,N_7454,N_6974);
or U7984 (N_7984,N_7443,N_6965);
or U7985 (N_7985,N_6699,N_7333);
nor U7986 (N_7986,N_6919,N_6902);
nor U7987 (N_7987,N_7150,N_6250);
and U7988 (N_7988,N_7152,N_6158);
and U7989 (N_7989,N_7494,N_6170);
nand U7990 (N_7990,N_6626,N_7351);
or U7991 (N_7991,N_6851,N_6021);
nor U7992 (N_7992,N_7173,N_6757);
and U7993 (N_7993,N_6450,N_6960);
xor U7994 (N_7994,N_6893,N_6804);
and U7995 (N_7995,N_6648,N_6577);
or U7996 (N_7996,N_6562,N_7227);
nor U7997 (N_7997,N_6799,N_6590);
nor U7998 (N_7998,N_7363,N_6839);
nor U7999 (N_7999,N_6263,N_7322);
or U8000 (N_8000,N_7188,N_6436);
nor U8001 (N_8001,N_6217,N_6980);
and U8002 (N_8002,N_6926,N_7419);
and U8003 (N_8003,N_6172,N_6526);
nand U8004 (N_8004,N_6331,N_7084);
nand U8005 (N_8005,N_7469,N_6270);
and U8006 (N_8006,N_6920,N_6700);
nand U8007 (N_8007,N_6294,N_7350);
nand U8008 (N_8008,N_7365,N_6637);
nand U8009 (N_8009,N_6207,N_7162);
or U8010 (N_8010,N_6029,N_7234);
nor U8011 (N_8011,N_6444,N_7155);
nand U8012 (N_8012,N_6030,N_6846);
nand U8013 (N_8013,N_6428,N_6045);
nor U8014 (N_8014,N_6083,N_7296);
and U8015 (N_8015,N_6681,N_7141);
nand U8016 (N_8016,N_6088,N_6123);
nor U8017 (N_8017,N_7259,N_7380);
nor U8018 (N_8018,N_7027,N_7346);
and U8019 (N_8019,N_6182,N_6366);
or U8020 (N_8020,N_7241,N_6456);
nor U8021 (N_8021,N_6269,N_7086);
and U8022 (N_8022,N_7098,N_7256);
and U8023 (N_8023,N_6095,N_7444);
xnor U8024 (N_8024,N_6232,N_7472);
nor U8025 (N_8025,N_6001,N_6979);
nor U8026 (N_8026,N_6797,N_7025);
nand U8027 (N_8027,N_6361,N_6824);
nand U8028 (N_8028,N_6976,N_7074);
or U8029 (N_8029,N_6322,N_6802);
or U8030 (N_8030,N_6295,N_6201);
nand U8031 (N_8031,N_6664,N_7349);
or U8032 (N_8032,N_6082,N_7398);
or U8033 (N_8033,N_6165,N_6168);
xor U8034 (N_8034,N_6848,N_6801);
nand U8035 (N_8035,N_6264,N_6835);
nor U8036 (N_8036,N_6929,N_6058);
and U8037 (N_8037,N_6244,N_7063);
and U8038 (N_8038,N_6011,N_6898);
xnor U8039 (N_8039,N_7212,N_6305);
and U8040 (N_8040,N_6559,N_6364);
nor U8041 (N_8041,N_7369,N_6261);
and U8042 (N_8042,N_6047,N_6570);
and U8043 (N_8043,N_6751,N_7140);
nor U8044 (N_8044,N_6195,N_6847);
and U8045 (N_8045,N_6491,N_6995);
or U8046 (N_8046,N_7396,N_6943);
nor U8047 (N_8047,N_6940,N_7432);
and U8048 (N_8048,N_6527,N_7048);
or U8049 (N_8049,N_6378,N_6094);
nand U8050 (N_8050,N_6518,N_6080);
or U8051 (N_8051,N_7132,N_6101);
and U8052 (N_8052,N_6057,N_6872);
and U8053 (N_8053,N_6375,N_7383);
or U8054 (N_8054,N_7273,N_7401);
and U8055 (N_8055,N_7230,N_6418);
xnor U8056 (N_8056,N_6566,N_6137);
and U8057 (N_8057,N_6933,N_6401);
nand U8058 (N_8058,N_7254,N_6892);
nor U8059 (N_8059,N_7438,N_7373);
or U8060 (N_8060,N_6449,N_7391);
nor U8061 (N_8061,N_6604,N_6100);
nand U8062 (N_8062,N_6161,N_6510);
and U8063 (N_8063,N_7368,N_6828);
nor U8064 (N_8064,N_6663,N_7470);
nand U8065 (N_8065,N_7095,N_6524);
nand U8066 (N_8066,N_7361,N_6576);
or U8067 (N_8067,N_6483,N_6311);
and U8068 (N_8068,N_6180,N_7379);
and U8069 (N_8069,N_6086,N_6964);
nand U8070 (N_8070,N_6658,N_7119);
xnor U8071 (N_8071,N_6399,N_7103);
or U8072 (N_8072,N_6462,N_6038);
or U8073 (N_8073,N_6685,N_6617);
nor U8074 (N_8074,N_6523,N_7124);
and U8075 (N_8075,N_7335,N_7252);
and U8076 (N_8076,N_6417,N_6895);
and U8077 (N_8077,N_6492,N_6785);
xor U8078 (N_8078,N_7455,N_6654);
xnor U8079 (N_8079,N_7097,N_7088);
and U8080 (N_8080,N_6563,N_7204);
nand U8081 (N_8081,N_7215,N_6286);
and U8082 (N_8082,N_7465,N_6737);
or U8083 (N_8083,N_7294,N_6997);
nand U8084 (N_8084,N_6597,N_7317);
or U8085 (N_8085,N_6642,N_7477);
xnor U8086 (N_8086,N_7394,N_7221);
and U8087 (N_8087,N_6142,N_6937);
xnor U8088 (N_8088,N_7414,N_6888);
nor U8089 (N_8089,N_7105,N_7448);
and U8090 (N_8090,N_7288,N_6512);
and U8091 (N_8091,N_6760,N_7026);
nor U8092 (N_8092,N_6060,N_7474);
nor U8093 (N_8093,N_6955,N_7435);
nand U8094 (N_8094,N_6114,N_7471);
nor U8095 (N_8095,N_6225,N_6246);
and U8096 (N_8096,N_6465,N_6909);
or U8097 (N_8097,N_6461,N_6359);
nor U8098 (N_8098,N_6766,N_6677);
and U8099 (N_8099,N_7484,N_7171);
or U8100 (N_8100,N_6404,N_6765);
xnor U8101 (N_8101,N_6345,N_6927);
nand U8102 (N_8102,N_7266,N_6175);
or U8103 (N_8103,N_6368,N_6341);
nand U8104 (N_8104,N_7497,N_6500);
nor U8105 (N_8105,N_6540,N_6342);
nand U8106 (N_8106,N_6517,N_7305);
and U8107 (N_8107,N_7163,N_7199);
nor U8108 (N_8108,N_6167,N_7232);
nor U8109 (N_8109,N_6209,N_6395);
nor U8110 (N_8110,N_6482,N_6199);
nand U8111 (N_8111,N_6105,N_6915);
or U8112 (N_8112,N_6275,N_7293);
and U8113 (N_8113,N_7218,N_7460);
nor U8114 (N_8114,N_6689,N_7004);
and U8115 (N_8115,N_6197,N_6961);
or U8116 (N_8116,N_6445,N_7016);
nand U8117 (N_8117,N_6556,N_6076);
and U8118 (N_8118,N_6612,N_7220);
and U8119 (N_8119,N_6103,N_7154);
nor U8120 (N_8120,N_6440,N_7091);
nand U8121 (N_8121,N_7329,N_6605);
nor U8122 (N_8122,N_6099,N_6587);
nand U8123 (N_8123,N_7195,N_6187);
nor U8124 (N_8124,N_6729,N_7242);
or U8125 (N_8125,N_6357,N_6304);
and U8126 (N_8126,N_6434,N_6949);
nand U8127 (N_8127,N_7113,N_7209);
nor U8128 (N_8128,N_6877,N_7126);
nor U8129 (N_8129,N_6254,N_6497);
or U8130 (N_8130,N_6229,N_6538);
and U8131 (N_8131,N_7156,N_6173);
nor U8132 (N_8132,N_7231,N_6191);
or U8133 (N_8133,N_7104,N_6134);
and U8134 (N_8134,N_7450,N_6635);
or U8135 (N_8135,N_7274,N_7111);
or U8136 (N_8136,N_6242,N_7107);
nor U8137 (N_8137,N_7357,N_6545);
and U8138 (N_8138,N_6561,N_7135);
nor U8139 (N_8139,N_6731,N_6452);
or U8140 (N_8140,N_6223,N_6831);
or U8141 (N_8141,N_6581,N_6052);
xnor U8142 (N_8142,N_6477,N_7115);
or U8143 (N_8143,N_6236,N_7307);
nand U8144 (N_8144,N_7372,N_6159);
nor U8145 (N_8145,N_7487,N_7424);
nand U8146 (N_8146,N_7381,N_7279);
nand U8147 (N_8147,N_7407,N_6122);
nor U8148 (N_8148,N_6551,N_6155);
nand U8149 (N_8149,N_6301,N_6127);
nor U8150 (N_8150,N_7172,N_7183);
nor U8151 (N_8151,N_6917,N_6216);
or U8152 (N_8152,N_6186,N_7428);
xor U8153 (N_8153,N_6431,N_6742);
or U8154 (N_8154,N_7042,N_7476);
nand U8155 (N_8155,N_6328,N_6202);
nor U8156 (N_8156,N_6544,N_7389);
xnor U8157 (N_8157,N_7239,N_6005);
nand U8158 (N_8158,N_6277,N_6297);
nor U8159 (N_8159,N_6371,N_6325);
xnor U8160 (N_8160,N_6494,N_7196);
nand U8161 (N_8161,N_6531,N_7403);
nor U8162 (N_8162,N_7493,N_6711);
or U8163 (N_8163,N_6779,N_6816);
nand U8164 (N_8164,N_6110,N_6734);
nor U8165 (N_8165,N_6379,N_6150);
nor U8166 (N_8166,N_7076,N_6078);
or U8167 (N_8167,N_7015,N_7033);
or U8168 (N_8168,N_6420,N_6111);
nand U8169 (N_8169,N_6881,N_6166);
nor U8170 (N_8170,N_6588,N_6337);
or U8171 (N_8171,N_6918,N_6905);
xor U8172 (N_8172,N_6387,N_6676);
xor U8173 (N_8173,N_6936,N_6959);
nand U8174 (N_8174,N_7366,N_6672);
or U8175 (N_8175,N_6247,N_6709);
nand U8176 (N_8176,N_6945,N_7049);
and U8177 (N_8177,N_7039,N_7182);
and U8178 (N_8178,N_7377,N_7343);
and U8179 (N_8179,N_6278,N_6422);
nor U8180 (N_8180,N_6564,N_6525);
nand U8181 (N_8181,N_6686,N_6954);
nor U8182 (N_8182,N_7219,N_6385);
or U8183 (N_8183,N_6208,N_7020);
nand U8184 (N_8184,N_7496,N_7133);
and U8185 (N_8185,N_6162,N_6849);
nand U8186 (N_8186,N_6822,N_6427);
or U8187 (N_8187,N_6611,N_6539);
or U8188 (N_8188,N_7269,N_6307);
xnor U8189 (N_8189,N_7384,N_6916);
nor U8190 (N_8190,N_6719,N_6671);
or U8191 (N_8191,N_7453,N_6485);
or U8192 (N_8192,N_6352,N_6715);
nor U8193 (N_8193,N_7406,N_6343);
nor U8194 (N_8194,N_7488,N_6806);
xor U8195 (N_8195,N_6136,N_6693);
nor U8196 (N_8196,N_6922,N_6971);
xor U8197 (N_8197,N_7499,N_7008);
or U8198 (N_8198,N_7479,N_6932);
nor U8199 (N_8199,N_7374,N_6002);
or U8200 (N_8200,N_6290,N_7367);
nand U8201 (N_8201,N_6458,N_6181);
and U8202 (N_8202,N_6227,N_7278);
nor U8203 (N_8203,N_6644,N_7275);
nand U8204 (N_8204,N_6392,N_6532);
and U8205 (N_8205,N_7179,N_6476);
nand U8206 (N_8206,N_6367,N_7201);
and U8207 (N_8207,N_7393,N_6090);
or U8208 (N_8208,N_6188,N_6455);
or U8209 (N_8209,N_6786,N_7408);
and U8210 (N_8210,N_7325,N_7375);
or U8211 (N_8211,N_6972,N_7180);
or U8212 (N_8212,N_6028,N_6988);
nor U8213 (N_8213,N_6521,N_7101);
xnor U8214 (N_8214,N_6200,N_6529);
nor U8215 (N_8215,N_6546,N_6493);
and U8216 (N_8216,N_7360,N_6198);
nand U8217 (N_8217,N_7404,N_6841);
and U8218 (N_8218,N_6360,N_6696);
and U8219 (N_8219,N_7328,N_6921);
or U8220 (N_8220,N_6594,N_6710);
xnor U8221 (N_8221,N_6017,N_7023);
xnor U8222 (N_8222,N_7090,N_7143);
and U8223 (N_8223,N_7029,N_7127);
and U8224 (N_8224,N_7011,N_6183);
xor U8225 (N_8225,N_7440,N_6853);
nor U8226 (N_8226,N_6023,N_6651);
nor U8227 (N_8227,N_7190,N_7250);
or U8228 (N_8228,N_7475,N_7019);
or U8229 (N_8229,N_7066,N_6947);
nor U8230 (N_8230,N_7382,N_7426);
and U8231 (N_8231,N_6754,N_6389);
xnor U8232 (N_8232,N_7174,N_7385);
xor U8233 (N_8233,N_6050,N_6724);
xnor U8234 (N_8234,N_6749,N_6204);
and U8235 (N_8235,N_6153,N_6390);
and U8236 (N_8236,N_6618,N_6614);
nor U8237 (N_8237,N_6743,N_6329);
nor U8238 (N_8238,N_7257,N_7009);
nor U8239 (N_8239,N_7415,N_6237);
nand U8240 (N_8240,N_7422,N_6335);
xnor U8241 (N_8241,N_6135,N_6646);
or U8242 (N_8242,N_7261,N_6293);
nand U8243 (N_8243,N_7338,N_6377);
and U8244 (N_8244,N_6780,N_6981);
or U8245 (N_8245,N_6467,N_6747);
or U8246 (N_8246,N_6224,N_6333);
and U8247 (N_8247,N_6800,N_6203);
nand U8248 (N_8248,N_7356,N_6627);
nand U8249 (N_8249,N_6138,N_6206);
or U8250 (N_8250,N_6356,N_6730);
nor U8251 (N_8251,N_6127,N_6562);
nand U8252 (N_8252,N_6570,N_6738);
and U8253 (N_8253,N_6326,N_7440);
or U8254 (N_8254,N_6662,N_7280);
and U8255 (N_8255,N_6050,N_6463);
or U8256 (N_8256,N_6034,N_6369);
xnor U8257 (N_8257,N_6697,N_7470);
and U8258 (N_8258,N_7281,N_7091);
nand U8259 (N_8259,N_6240,N_6332);
xor U8260 (N_8260,N_6425,N_6573);
and U8261 (N_8261,N_7008,N_6446);
xnor U8262 (N_8262,N_6672,N_6886);
or U8263 (N_8263,N_6123,N_6297);
and U8264 (N_8264,N_6554,N_7284);
nand U8265 (N_8265,N_7459,N_6111);
nor U8266 (N_8266,N_6575,N_7370);
or U8267 (N_8267,N_6300,N_7045);
nand U8268 (N_8268,N_6990,N_6534);
nor U8269 (N_8269,N_7443,N_6988);
or U8270 (N_8270,N_6096,N_6943);
nand U8271 (N_8271,N_6524,N_6507);
nor U8272 (N_8272,N_6945,N_7199);
or U8273 (N_8273,N_6274,N_6896);
xnor U8274 (N_8274,N_6000,N_6953);
and U8275 (N_8275,N_7471,N_6569);
nor U8276 (N_8276,N_6580,N_7482);
nand U8277 (N_8277,N_6690,N_7198);
xor U8278 (N_8278,N_7189,N_6824);
xor U8279 (N_8279,N_6304,N_6197);
nor U8280 (N_8280,N_6471,N_6309);
and U8281 (N_8281,N_7430,N_6987);
and U8282 (N_8282,N_7403,N_6973);
nand U8283 (N_8283,N_6025,N_6796);
nor U8284 (N_8284,N_6226,N_7099);
nand U8285 (N_8285,N_6634,N_6016);
and U8286 (N_8286,N_7347,N_6536);
or U8287 (N_8287,N_6160,N_7078);
or U8288 (N_8288,N_6643,N_6193);
or U8289 (N_8289,N_6138,N_6088);
nor U8290 (N_8290,N_7308,N_7217);
and U8291 (N_8291,N_7294,N_6772);
nand U8292 (N_8292,N_6443,N_6590);
and U8293 (N_8293,N_6239,N_7492);
or U8294 (N_8294,N_7152,N_7233);
and U8295 (N_8295,N_7381,N_6556);
nand U8296 (N_8296,N_6756,N_7253);
or U8297 (N_8297,N_7396,N_6186);
nor U8298 (N_8298,N_7057,N_6060);
or U8299 (N_8299,N_6824,N_6579);
nand U8300 (N_8300,N_6765,N_6466);
nor U8301 (N_8301,N_6395,N_6021);
and U8302 (N_8302,N_6888,N_7283);
and U8303 (N_8303,N_6817,N_6128);
nor U8304 (N_8304,N_6647,N_6934);
and U8305 (N_8305,N_6192,N_6086);
nand U8306 (N_8306,N_6795,N_6859);
nand U8307 (N_8307,N_6783,N_6230);
nand U8308 (N_8308,N_6844,N_6894);
or U8309 (N_8309,N_6195,N_6733);
nand U8310 (N_8310,N_6992,N_6891);
and U8311 (N_8311,N_7131,N_6086);
or U8312 (N_8312,N_6920,N_7087);
or U8313 (N_8313,N_6357,N_6002);
and U8314 (N_8314,N_7320,N_6359);
nor U8315 (N_8315,N_7305,N_6650);
and U8316 (N_8316,N_6875,N_6456);
or U8317 (N_8317,N_6433,N_6641);
or U8318 (N_8318,N_6462,N_6409);
xor U8319 (N_8319,N_6024,N_7416);
or U8320 (N_8320,N_7356,N_6052);
nor U8321 (N_8321,N_7068,N_6954);
and U8322 (N_8322,N_7156,N_6876);
and U8323 (N_8323,N_6835,N_7411);
and U8324 (N_8324,N_7365,N_7275);
nor U8325 (N_8325,N_7065,N_6090);
nor U8326 (N_8326,N_6805,N_6362);
xor U8327 (N_8327,N_6351,N_7052);
and U8328 (N_8328,N_6533,N_7344);
and U8329 (N_8329,N_7476,N_6855);
nand U8330 (N_8330,N_7190,N_6631);
and U8331 (N_8331,N_7382,N_6739);
xnor U8332 (N_8332,N_7233,N_6385);
nor U8333 (N_8333,N_6664,N_7219);
nor U8334 (N_8334,N_6190,N_6073);
nor U8335 (N_8335,N_6163,N_7405);
nor U8336 (N_8336,N_7287,N_6383);
or U8337 (N_8337,N_7381,N_6635);
xor U8338 (N_8338,N_7323,N_7443);
nand U8339 (N_8339,N_6486,N_6075);
nor U8340 (N_8340,N_6859,N_6900);
nand U8341 (N_8341,N_7466,N_7145);
nand U8342 (N_8342,N_6914,N_7479);
or U8343 (N_8343,N_6107,N_6602);
or U8344 (N_8344,N_6167,N_6320);
or U8345 (N_8345,N_7241,N_7469);
nand U8346 (N_8346,N_6655,N_6963);
or U8347 (N_8347,N_7061,N_6690);
nand U8348 (N_8348,N_7145,N_6037);
nand U8349 (N_8349,N_6345,N_6969);
and U8350 (N_8350,N_6364,N_6702);
xor U8351 (N_8351,N_7017,N_6873);
and U8352 (N_8352,N_7429,N_7029);
or U8353 (N_8353,N_6369,N_6029);
or U8354 (N_8354,N_6480,N_6797);
or U8355 (N_8355,N_6679,N_6727);
nor U8356 (N_8356,N_7469,N_6934);
nor U8357 (N_8357,N_6755,N_7374);
and U8358 (N_8358,N_6939,N_7496);
nand U8359 (N_8359,N_6708,N_6309);
nand U8360 (N_8360,N_6164,N_6602);
xor U8361 (N_8361,N_6525,N_7004);
nor U8362 (N_8362,N_6227,N_6262);
and U8363 (N_8363,N_6073,N_7048);
and U8364 (N_8364,N_6718,N_6755);
nor U8365 (N_8365,N_6422,N_6408);
nand U8366 (N_8366,N_7103,N_6893);
and U8367 (N_8367,N_6667,N_6561);
and U8368 (N_8368,N_6886,N_6728);
and U8369 (N_8369,N_6459,N_6473);
or U8370 (N_8370,N_7354,N_6529);
nand U8371 (N_8371,N_6072,N_6628);
nand U8372 (N_8372,N_7104,N_6229);
nor U8373 (N_8373,N_6255,N_7405);
nand U8374 (N_8374,N_6239,N_6397);
or U8375 (N_8375,N_6677,N_6303);
nand U8376 (N_8376,N_7154,N_7028);
or U8377 (N_8377,N_6191,N_7156);
and U8378 (N_8378,N_6536,N_7217);
and U8379 (N_8379,N_6464,N_6079);
nand U8380 (N_8380,N_6935,N_6436);
and U8381 (N_8381,N_6358,N_6513);
or U8382 (N_8382,N_7182,N_6757);
nand U8383 (N_8383,N_6704,N_6237);
or U8384 (N_8384,N_6403,N_6271);
or U8385 (N_8385,N_6748,N_6579);
or U8386 (N_8386,N_6999,N_6570);
nand U8387 (N_8387,N_6236,N_6483);
nand U8388 (N_8388,N_6721,N_6941);
or U8389 (N_8389,N_6112,N_7108);
nand U8390 (N_8390,N_6330,N_6209);
and U8391 (N_8391,N_6042,N_7349);
or U8392 (N_8392,N_7084,N_6519);
and U8393 (N_8393,N_6357,N_6998);
and U8394 (N_8394,N_6962,N_6529);
and U8395 (N_8395,N_6449,N_7405);
xnor U8396 (N_8396,N_6086,N_7338);
nor U8397 (N_8397,N_7484,N_6111);
nor U8398 (N_8398,N_7250,N_6223);
or U8399 (N_8399,N_7070,N_6608);
nor U8400 (N_8400,N_7403,N_7243);
xor U8401 (N_8401,N_7095,N_6531);
and U8402 (N_8402,N_6932,N_6379);
xor U8403 (N_8403,N_6261,N_6743);
nand U8404 (N_8404,N_6969,N_6126);
xor U8405 (N_8405,N_6116,N_6912);
nand U8406 (N_8406,N_6738,N_6185);
nor U8407 (N_8407,N_6697,N_6986);
nand U8408 (N_8408,N_6501,N_6488);
and U8409 (N_8409,N_6432,N_6303);
nand U8410 (N_8410,N_6930,N_6559);
nor U8411 (N_8411,N_7219,N_6672);
or U8412 (N_8412,N_6142,N_7296);
nor U8413 (N_8413,N_6269,N_6726);
or U8414 (N_8414,N_7309,N_6903);
nand U8415 (N_8415,N_6998,N_6454);
and U8416 (N_8416,N_6329,N_6942);
and U8417 (N_8417,N_6749,N_7264);
or U8418 (N_8418,N_7211,N_7223);
and U8419 (N_8419,N_6060,N_7433);
nand U8420 (N_8420,N_6682,N_6589);
nor U8421 (N_8421,N_7279,N_6420);
and U8422 (N_8422,N_6968,N_6358);
or U8423 (N_8423,N_6367,N_6941);
nand U8424 (N_8424,N_7496,N_6046);
or U8425 (N_8425,N_7335,N_6803);
nor U8426 (N_8426,N_7318,N_6691);
xor U8427 (N_8427,N_7499,N_7443);
or U8428 (N_8428,N_7491,N_7373);
nand U8429 (N_8429,N_6825,N_6442);
xor U8430 (N_8430,N_6934,N_6682);
xor U8431 (N_8431,N_7320,N_6246);
or U8432 (N_8432,N_6932,N_7120);
and U8433 (N_8433,N_6372,N_6226);
nand U8434 (N_8434,N_7098,N_7190);
or U8435 (N_8435,N_7230,N_6366);
and U8436 (N_8436,N_6986,N_6027);
and U8437 (N_8437,N_7122,N_7017);
nor U8438 (N_8438,N_6266,N_6226);
or U8439 (N_8439,N_7031,N_6809);
and U8440 (N_8440,N_6944,N_6567);
nand U8441 (N_8441,N_6261,N_6165);
nand U8442 (N_8442,N_6213,N_7264);
nand U8443 (N_8443,N_6661,N_6070);
nand U8444 (N_8444,N_7143,N_7217);
nor U8445 (N_8445,N_7124,N_7410);
nand U8446 (N_8446,N_6737,N_6395);
and U8447 (N_8447,N_6296,N_7003);
nand U8448 (N_8448,N_6195,N_6334);
or U8449 (N_8449,N_6645,N_6098);
or U8450 (N_8450,N_6860,N_6725);
and U8451 (N_8451,N_7122,N_7466);
nor U8452 (N_8452,N_6403,N_6767);
nand U8453 (N_8453,N_7131,N_7489);
or U8454 (N_8454,N_7225,N_6952);
xnor U8455 (N_8455,N_6570,N_6157);
nor U8456 (N_8456,N_7469,N_6790);
xnor U8457 (N_8457,N_7364,N_6387);
or U8458 (N_8458,N_6342,N_7489);
or U8459 (N_8459,N_6461,N_7145);
nand U8460 (N_8460,N_6417,N_7058);
nor U8461 (N_8461,N_7485,N_7364);
xnor U8462 (N_8462,N_6171,N_6590);
and U8463 (N_8463,N_6797,N_6757);
nand U8464 (N_8464,N_6900,N_7334);
and U8465 (N_8465,N_6032,N_6480);
nand U8466 (N_8466,N_6736,N_7279);
and U8467 (N_8467,N_6473,N_6047);
xor U8468 (N_8468,N_6755,N_6192);
or U8469 (N_8469,N_6849,N_6783);
nand U8470 (N_8470,N_6783,N_6421);
and U8471 (N_8471,N_6127,N_6296);
nand U8472 (N_8472,N_7344,N_6935);
and U8473 (N_8473,N_7003,N_6502);
or U8474 (N_8474,N_7367,N_6456);
or U8475 (N_8475,N_6718,N_6783);
nor U8476 (N_8476,N_6735,N_7405);
nor U8477 (N_8477,N_6692,N_6128);
nand U8478 (N_8478,N_6576,N_7285);
or U8479 (N_8479,N_6426,N_7285);
nand U8480 (N_8480,N_6800,N_6831);
xor U8481 (N_8481,N_6831,N_7470);
and U8482 (N_8482,N_6906,N_6862);
or U8483 (N_8483,N_7144,N_7467);
xor U8484 (N_8484,N_7482,N_7359);
and U8485 (N_8485,N_7033,N_7211);
nor U8486 (N_8486,N_7213,N_6398);
nor U8487 (N_8487,N_6990,N_7486);
nand U8488 (N_8488,N_7381,N_7370);
and U8489 (N_8489,N_6579,N_7185);
nor U8490 (N_8490,N_6288,N_6152);
nor U8491 (N_8491,N_6275,N_6789);
or U8492 (N_8492,N_7478,N_7175);
xnor U8493 (N_8493,N_7335,N_7447);
and U8494 (N_8494,N_6232,N_7465);
and U8495 (N_8495,N_6866,N_6610);
or U8496 (N_8496,N_7014,N_7225);
nand U8497 (N_8497,N_7476,N_7304);
or U8498 (N_8498,N_7300,N_6139);
nor U8499 (N_8499,N_6053,N_6887);
nor U8500 (N_8500,N_6263,N_6615);
nor U8501 (N_8501,N_7080,N_6370);
and U8502 (N_8502,N_6189,N_6929);
nor U8503 (N_8503,N_6462,N_6626);
nand U8504 (N_8504,N_6534,N_6744);
nor U8505 (N_8505,N_6284,N_7459);
nand U8506 (N_8506,N_6896,N_7194);
xnor U8507 (N_8507,N_7272,N_7132);
xnor U8508 (N_8508,N_6204,N_6435);
and U8509 (N_8509,N_7441,N_6063);
nand U8510 (N_8510,N_6356,N_6074);
or U8511 (N_8511,N_7400,N_6690);
nor U8512 (N_8512,N_6891,N_6088);
nand U8513 (N_8513,N_6298,N_6272);
and U8514 (N_8514,N_6186,N_7427);
nand U8515 (N_8515,N_6125,N_6398);
nand U8516 (N_8516,N_6682,N_6539);
and U8517 (N_8517,N_6749,N_6578);
and U8518 (N_8518,N_6884,N_6892);
xnor U8519 (N_8519,N_7313,N_7117);
nand U8520 (N_8520,N_7368,N_6980);
nand U8521 (N_8521,N_7468,N_6391);
or U8522 (N_8522,N_6997,N_6091);
nand U8523 (N_8523,N_6593,N_7361);
or U8524 (N_8524,N_6899,N_6277);
or U8525 (N_8525,N_7496,N_6740);
nor U8526 (N_8526,N_7341,N_7368);
or U8527 (N_8527,N_6977,N_6011);
and U8528 (N_8528,N_6629,N_6134);
and U8529 (N_8529,N_7185,N_6951);
nand U8530 (N_8530,N_7324,N_6391);
nand U8531 (N_8531,N_7123,N_6718);
and U8532 (N_8532,N_6430,N_6829);
nor U8533 (N_8533,N_6986,N_6627);
or U8534 (N_8534,N_6308,N_6125);
nand U8535 (N_8535,N_7293,N_7100);
nor U8536 (N_8536,N_6363,N_7165);
nor U8537 (N_8537,N_6583,N_6234);
nor U8538 (N_8538,N_7298,N_6838);
nand U8539 (N_8539,N_6193,N_6866);
nand U8540 (N_8540,N_7274,N_6023);
or U8541 (N_8541,N_6676,N_7080);
or U8542 (N_8542,N_7211,N_7166);
nor U8543 (N_8543,N_6862,N_6037);
or U8544 (N_8544,N_6765,N_6003);
nor U8545 (N_8545,N_6890,N_6842);
and U8546 (N_8546,N_7447,N_7007);
nor U8547 (N_8547,N_6981,N_6782);
or U8548 (N_8548,N_7101,N_6888);
and U8549 (N_8549,N_6469,N_6153);
or U8550 (N_8550,N_7103,N_7458);
nor U8551 (N_8551,N_6612,N_7119);
nand U8552 (N_8552,N_6792,N_7392);
and U8553 (N_8553,N_6266,N_6999);
nor U8554 (N_8554,N_6052,N_6778);
or U8555 (N_8555,N_6511,N_7124);
and U8556 (N_8556,N_7270,N_7117);
nor U8557 (N_8557,N_6407,N_6698);
and U8558 (N_8558,N_6024,N_6389);
nand U8559 (N_8559,N_7049,N_6383);
nand U8560 (N_8560,N_6366,N_6161);
or U8561 (N_8561,N_6040,N_7168);
and U8562 (N_8562,N_6465,N_6421);
or U8563 (N_8563,N_7002,N_7222);
and U8564 (N_8564,N_7009,N_6142);
and U8565 (N_8565,N_7342,N_6699);
nor U8566 (N_8566,N_6782,N_6033);
nor U8567 (N_8567,N_6373,N_6502);
and U8568 (N_8568,N_6702,N_6104);
and U8569 (N_8569,N_6251,N_6663);
nor U8570 (N_8570,N_7234,N_7325);
nand U8571 (N_8571,N_6994,N_6249);
nand U8572 (N_8572,N_6758,N_6900);
or U8573 (N_8573,N_6630,N_6686);
nand U8574 (N_8574,N_6746,N_6193);
and U8575 (N_8575,N_6533,N_7154);
or U8576 (N_8576,N_6273,N_7266);
or U8577 (N_8577,N_7483,N_6131);
nor U8578 (N_8578,N_7313,N_6189);
and U8579 (N_8579,N_6157,N_6715);
nand U8580 (N_8580,N_7313,N_6317);
nor U8581 (N_8581,N_6475,N_6273);
nor U8582 (N_8582,N_7344,N_6778);
nand U8583 (N_8583,N_7248,N_6557);
and U8584 (N_8584,N_6190,N_6469);
nand U8585 (N_8585,N_6867,N_7336);
and U8586 (N_8586,N_6538,N_7487);
or U8587 (N_8587,N_7329,N_7258);
and U8588 (N_8588,N_6288,N_6830);
and U8589 (N_8589,N_6006,N_7207);
and U8590 (N_8590,N_6327,N_6701);
and U8591 (N_8591,N_7359,N_6707);
xnor U8592 (N_8592,N_6546,N_6062);
nor U8593 (N_8593,N_7009,N_7151);
or U8594 (N_8594,N_6164,N_7227);
nor U8595 (N_8595,N_7341,N_7279);
or U8596 (N_8596,N_7025,N_6314);
or U8597 (N_8597,N_7106,N_7016);
and U8598 (N_8598,N_7336,N_7252);
and U8599 (N_8599,N_6681,N_6442);
or U8600 (N_8600,N_6966,N_6497);
nand U8601 (N_8601,N_6027,N_6726);
and U8602 (N_8602,N_7337,N_6414);
xnor U8603 (N_8603,N_7465,N_7206);
nor U8604 (N_8604,N_6808,N_6175);
nor U8605 (N_8605,N_7270,N_6876);
and U8606 (N_8606,N_7199,N_6227);
nor U8607 (N_8607,N_6627,N_6874);
nand U8608 (N_8608,N_6844,N_7265);
or U8609 (N_8609,N_7007,N_6396);
nand U8610 (N_8610,N_6206,N_6016);
nand U8611 (N_8611,N_6747,N_6239);
or U8612 (N_8612,N_6613,N_6637);
and U8613 (N_8613,N_6599,N_6989);
and U8614 (N_8614,N_7137,N_7188);
or U8615 (N_8615,N_7003,N_6670);
nor U8616 (N_8616,N_6930,N_7283);
nand U8617 (N_8617,N_6958,N_6612);
nand U8618 (N_8618,N_6917,N_7035);
nand U8619 (N_8619,N_6084,N_7063);
nand U8620 (N_8620,N_7042,N_6425);
nand U8621 (N_8621,N_7215,N_7197);
or U8622 (N_8622,N_6870,N_6023);
and U8623 (N_8623,N_6588,N_6328);
or U8624 (N_8624,N_7436,N_6822);
xor U8625 (N_8625,N_6550,N_6567);
and U8626 (N_8626,N_6111,N_7183);
nand U8627 (N_8627,N_6220,N_7059);
nor U8628 (N_8628,N_6858,N_6374);
nor U8629 (N_8629,N_6967,N_6619);
or U8630 (N_8630,N_6814,N_6977);
and U8631 (N_8631,N_6783,N_6324);
and U8632 (N_8632,N_7327,N_6389);
nor U8633 (N_8633,N_6904,N_6759);
or U8634 (N_8634,N_6546,N_7070);
nor U8635 (N_8635,N_6798,N_6828);
nand U8636 (N_8636,N_6071,N_6941);
or U8637 (N_8637,N_6427,N_6634);
and U8638 (N_8638,N_6705,N_6684);
or U8639 (N_8639,N_6487,N_7483);
or U8640 (N_8640,N_6002,N_6702);
and U8641 (N_8641,N_7059,N_6457);
and U8642 (N_8642,N_6582,N_7367);
or U8643 (N_8643,N_6911,N_7126);
or U8644 (N_8644,N_6821,N_6163);
or U8645 (N_8645,N_6559,N_6316);
nor U8646 (N_8646,N_6847,N_7388);
nand U8647 (N_8647,N_7220,N_7293);
nand U8648 (N_8648,N_7239,N_7165);
or U8649 (N_8649,N_6074,N_7352);
or U8650 (N_8650,N_6875,N_6958);
nand U8651 (N_8651,N_6348,N_6196);
nand U8652 (N_8652,N_6374,N_6719);
and U8653 (N_8653,N_7471,N_7472);
nor U8654 (N_8654,N_7242,N_6370);
and U8655 (N_8655,N_6614,N_6346);
or U8656 (N_8656,N_7405,N_6776);
or U8657 (N_8657,N_6823,N_6004);
or U8658 (N_8658,N_6080,N_7334);
nor U8659 (N_8659,N_6986,N_6093);
or U8660 (N_8660,N_7069,N_7391);
nor U8661 (N_8661,N_7497,N_6057);
nand U8662 (N_8662,N_6600,N_6858);
nand U8663 (N_8663,N_6903,N_7001);
nand U8664 (N_8664,N_6130,N_7150);
nor U8665 (N_8665,N_6440,N_7485);
and U8666 (N_8666,N_6100,N_6314);
and U8667 (N_8667,N_6584,N_7012);
nor U8668 (N_8668,N_6460,N_6716);
or U8669 (N_8669,N_7312,N_6896);
or U8670 (N_8670,N_7138,N_6745);
and U8671 (N_8671,N_6939,N_6899);
nor U8672 (N_8672,N_7499,N_7294);
and U8673 (N_8673,N_6809,N_6011);
nand U8674 (N_8674,N_7261,N_6287);
and U8675 (N_8675,N_6656,N_6091);
and U8676 (N_8676,N_7137,N_6176);
nand U8677 (N_8677,N_6474,N_7310);
xnor U8678 (N_8678,N_7487,N_6382);
or U8679 (N_8679,N_7425,N_6500);
and U8680 (N_8680,N_7351,N_6369);
nor U8681 (N_8681,N_6194,N_6279);
nand U8682 (N_8682,N_6637,N_7208);
and U8683 (N_8683,N_6996,N_6849);
nand U8684 (N_8684,N_6829,N_6447);
and U8685 (N_8685,N_7426,N_6003);
or U8686 (N_8686,N_6388,N_6013);
or U8687 (N_8687,N_6592,N_6590);
nor U8688 (N_8688,N_6673,N_6309);
nor U8689 (N_8689,N_7228,N_6022);
or U8690 (N_8690,N_6541,N_7451);
or U8691 (N_8691,N_6901,N_6007);
nor U8692 (N_8692,N_7196,N_7316);
nor U8693 (N_8693,N_6817,N_6933);
or U8694 (N_8694,N_6986,N_6690);
nor U8695 (N_8695,N_6454,N_6516);
or U8696 (N_8696,N_6776,N_6962);
or U8697 (N_8697,N_6357,N_7423);
and U8698 (N_8698,N_7225,N_7059);
nor U8699 (N_8699,N_7395,N_6694);
nor U8700 (N_8700,N_6692,N_6277);
nor U8701 (N_8701,N_6902,N_6461);
and U8702 (N_8702,N_6685,N_6228);
or U8703 (N_8703,N_6941,N_6010);
nor U8704 (N_8704,N_7259,N_7063);
xor U8705 (N_8705,N_6636,N_6452);
nor U8706 (N_8706,N_7004,N_6524);
nand U8707 (N_8707,N_6264,N_7452);
or U8708 (N_8708,N_6639,N_6415);
nand U8709 (N_8709,N_7438,N_7082);
nand U8710 (N_8710,N_7466,N_6034);
nand U8711 (N_8711,N_6131,N_6884);
nor U8712 (N_8712,N_7061,N_7335);
or U8713 (N_8713,N_6628,N_6811);
nor U8714 (N_8714,N_6703,N_6627);
xor U8715 (N_8715,N_6749,N_6540);
or U8716 (N_8716,N_6612,N_7374);
nor U8717 (N_8717,N_6654,N_6668);
xnor U8718 (N_8718,N_7478,N_6759);
or U8719 (N_8719,N_7047,N_6608);
nand U8720 (N_8720,N_7272,N_6906);
nand U8721 (N_8721,N_7394,N_6799);
xnor U8722 (N_8722,N_6229,N_6347);
nor U8723 (N_8723,N_7157,N_7459);
and U8724 (N_8724,N_7017,N_6980);
or U8725 (N_8725,N_6419,N_7466);
xnor U8726 (N_8726,N_6223,N_6152);
nand U8727 (N_8727,N_7181,N_7376);
nor U8728 (N_8728,N_7387,N_6902);
nor U8729 (N_8729,N_6590,N_7223);
nand U8730 (N_8730,N_6792,N_6386);
nand U8731 (N_8731,N_7151,N_6083);
nor U8732 (N_8732,N_6483,N_7259);
or U8733 (N_8733,N_6005,N_6101);
or U8734 (N_8734,N_6774,N_7021);
xnor U8735 (N_8735,N_7232,N_6658);
nor U8736 (N_8736,N_6657,N_6968);
and U8737 (N_8737,N_6247,N_6858);
nor U8738 (N_8738,N_6647,N_6580);
nand U8739 (N_8739,N_6830,N_6088);
or U8740 (N_8740,N_7153,N_7032);
xnor U8741 (N_8741,N_7450,N_6711);
or U8742 (N_8742,N_6239,N_7132);
nor U8743 (N_8743,N_6923,N_7029);
nand U8744 (N_8744,N_7017,N_6872);
and U8745 (N_8745,N_6476,N_6281);
and U8746 (N_8746,N_6011,N_6371);
nor U8747 (N_8747,N_6166,N_6337);
nor U8748 (N_8748,N_6290,N_6168);
or U8749 (N_8749,N_7410,N_7092);
nor U8750 (N_8750,N_6861,N_7409);
or U8751 (N_8751,N_6781,N_6170);
nor U8752 (N_8752,N_6656,N_6786);
nand U8753 (N_8753,N_6157,N_7113);
and U8754 (N_8754,N_7096,N_6977);
or U8755 (N_8755,N_7138,N_7318);
and U8756 (N_8756,N_6961,N_6551);
nand U8757 (N_8757,N_6885,N_6386);
nand U8758 (N_8758,N_6689,N_6895);
and U8759 (N_8759,N_6458,N_6753);
nor U8760 (N_8760,N_7055,N_6812);
nand U8761 (N_8761,N_6100,N_7084);
or U8762 (N_8762,N_7031,N_6410);
and U8763 (N_8763,N_6852,N_6614);
nor U8764 (N_8764,N_7022,N_6350);
nand U8765 (N_8765,N_6474,N_6929);
nand U8766 (N_8766,N_6024,N_6013);
nand U8767 (N_8767,N_6158,N_6413);
or U8768 (N_8768,N_6404,N_6579);
and U8769 (N_8769,N_6739,N_6469);
nor U8770 (N_8770,N_6834,N_7274);
nor U8771 (N_8771,N_6086,N_7498);
nand U8772 (N_8772,N_6928,N_7391);
nand U8773 (N_8773,N_6316,N_6161);
and U8774 (N_8774,N_7314,N_7291);
nor U8775 (N_8775,N_6834,N_7147);
and U8776 (N_8776,N_6595,N_6618);
or U8777 (N_8777,N_6617,N_6707);
nor U8778 (N_8778,N_6380,N_7187);
or U8779 (N_8779,N_6342,N_6091);
nand U8780 (N_8780,N_6422,N_7332);
and U8781 (N_8781,N_7499,N_7485);
xnor U8782 (N_8782,N_7275,N_6427);
and U8783 (N_8783,N_6537,N_7490);
nor U8784 (N_8784,N_7140,N_6234);
and U8785 (N_8785,N_6103,N_6329);
nand U8786 (N_8786,N_6915,N_7064);
nand U8787 (N_8787,N_6807,N_7050);
xor U8788 (N_8788,N_7322,N_7429);
nand U8789 (N_8789,N_7425,N_7239);
xor U8790 (N_8790,N_6457,N_7499);
nor U8791 (N_8791,N_7321,N_7285);
nor U8792 (N_8792,N_6117,N_7315);
or U8793 (N_8793,N_7263,N_7180);
nor U8794 (N_8794,N_6112,N_6159);
nand U8795 (N_8795,N_7062,N_6499);
and U8796 (N_8796,N_6615,N_7069);
nor U8797 (N_8797,N_6033,N_6824);
and U8798 (N_8798,N_7019,N_6067);
nor U8799 (N_8799,N_6272,N_7175);
nand U8800 (N_8800,N_6155,N_7297);
xnor U8801 (N_8801,N_6120,N_7265);
or U8802 (N_8802,N_6657,N_6166);
xnor U8803 (N_8803,N_6272,N_7075);
nand U8804 (N_8804,N_6753,N_7396);
nor U8805 (N_8805,N_6184,N_7197);
and U8806 (N_8806,N_6129,N_6959);
and U8807 (N_8807,N_7402,N_7172);
nor U8808 (N_8808,N_7485,N_7234);
or U8809 (N_8809,N_6326,N_6840);
xor U8810 (N_8810,N_6997,N_7190);
nand U8811 (N_8811,N_7076,N_7201);
nor U8812 (N_8812,N_7337,N_6927);
nor U8813 (N_8813,N_6695,N_6843);
nor U8814 (N_8814,N_7136,N_6955);
nand U8815 (N_8815,N_6462,N_6432);
nand U8816 (N_8816,N_6893,N_7283);
or U8817 (N_8817,N_7217,N_7341);
or U8818 (N_8818,N_6908,N_6112);
or U8819 (N_8819,N_6382,N_6240);
and U8820 (N_8820,N_7282,N_7408);
or U8821 (N_8821,N_7351,N_6882);
and U8822 (N_8822,N_6278,N_6604);
or U8823 (N_8823,N_7374,N_6946);
nor U8824 (N_8824,N_6443,N_6724);
and U8825 (N_8825,N_6289,N_6539);
and U8826 (N_8826,N_6693,N_6730);
nor U8827 (N_8827,N_6307,N_7112);
nand U8828 (N_8828,N_6193,N_7376);
nand U8829 (N_8829,N_6811,N_6692);
nand U8830 (N_8830,N_7224,N_6693);
nor U8831 (N_8831,N_6941,N_6100);
and U8832 (N_8832,N_6796,N_6745);
and U8833 (N_8833,N_7072,N_7276);
or U8834 (N_8834,N_7313,N_6589);
nor U8835 (N_8835,N_7020,N_6039);
nand U8836 (N_8836,N_7013,N_6543);
or U8837 (N_8837,N_7335,N_7282);
nor U8838 (N_8838,N_6810,N_6597);
and U8839 (N_8839,N_6268,N_7382);
nand U8840 (N_8840,N_6242,N_7452);
or U8841 (N_8841,N_6856,N_6637);
nor U8842 (N_8842,N_6313,N_6334);
or U8843 (N_8843,N_6815,N_7322);
and U8844 (N_8844,N_6189,N_6895);
nand U8845 (N_8845,N_6285,N_6836);
nand U8846 (N_8846,N_6981,N_6111);
xnor U8847 (N_8847,N_7093,N_7051);
and U8848 (N_8848,N_7206,N_6161);
and U8849 (N_8849,N_6866,N_6967);
nand U8850 (N_8850,N_6844,N_7136);
and U8851 (N_8851,N_7370,N_6863);
xor U8852 (N_8852,N_7082,N_6762);
nand U8853 (N_8853,N_6712,N_6562);
or U8854 (N_8854,N_6041,N_6463);
nor U8855 (N_8855,N_6932,N_6683);
or U8856 (N_8856,N_6051,N_6819);
nand U8857 (N_8857,N_7055,N_6064);
and U8858 (N_8858,N_6160,N_6085);
nand U8859 (N_8859,N_6856,N_6844);
or U8860 (N_8860,N_6650,N_6503);
or U8861 (N_8861,N_7077,N_6088);
xnor U8862 (N_8862,N_6810,N_6957);
or U8863 (N_8863,N_6100,N_6460);
nand U8864 (N_8864,N_7331,N_6659);
and U8865 (N_8865,N_6154,N_6772);
nand U8866 (N_8866,N_6199,N_7127);
xnor U8867 (N_8867,N_6490,N_6746);
and U8868 (N_8868,N_7222,N_6391);
nor U8869 (N_8869,N_6182,N_6855);
and U8870 (N_8870,N_7125,N_6966);
and U8871 (N_8871,N_7062,N_6945);
nand U8872 (N_8872,N_6959,N_6404);
and U8873 (N_8873,N_7426,N_6676);
nand U8874 (N_8874,N_6270,N_6147);
nand U8875 (N_8875,N_7220,N_7246);
nor U8876 (N_8876,N_7269,N_7326);
xor U8877 (N_8877,N_7200,N_7113);
or U8878 (N_8878,N_6587,N_6908);
and U8879 (N_8879,N_7369,N_7406);
xnor U8880 (N_8880,N_7114,N_7000);
and U8881 (N_8881,N_7340,N_7120);
nor U8882 (N_8882,N_6298,N_6899);
xnor U8883 (N_8883,N_7219,N_7134);
or U8884 (N_8884,N_7276,N_7497);
nor U8885 (N_8885,N_6778,N_6155);
or U8886 (N_8886,N_6694,N_6447);
xor U8887 (N_8887,N_6089,N_6401);
nor U8888 (N_8888,N_6862,N_6133);
nand U8889 (N_8889,N_7419,N_6475);
nand U8890 (N_8890,N_6597,N_7028);
and U8891 (N_8891,N_6701,N_6261);
and U8892 (N_8892,N_7166,N_6616);
or U8893 (N_8893,N_6752,N_6521);
and U8894 (N_8894,N_7201,N_7294);
xnor U8895 (N_8895,N_6976,N_6702);
and U8896 (N_8896,N_7204,N_6223);
or U8897 (N_8897,N_7008,N_6016);
and U8898 (N_8898,N_7475,N_6676);
nand U8899 (N_8899,N_7282,N_7262);
nor U8900 (N_8900,N_6803,N_7354);
nand U8901 (N_8901,N_7048,N_6802);
or U8902 (N_8902,N_6148,N_6693);
nor U8903 (N_8903,N_7461,N_6123);
nand U8904 (N_8904,N_6811,N_6517);
nor U8905 (N_8905,N_6187,N_7486);
nor U8906 (N_8906,N_6135,N_6725);
and U8907 (N_8907,N_6638,N_7423);
xor U8908 (N_8908,N_7181,N_7138);
nor U8909 (N_8909,N_6697,N_6790);
and U8910 (N_8910,N_6334,N_6805);
nand U8911 (N_8911,N_6368,N_6931);
and U8912 (N_8912,N_6961,N_6752);
and U8913 (N_8913,N_7114,N_6146);
nand U8914 (N_8914,N_7401,N_6425);
nand U8915 (N_8915,N_7030,N_6346);
nor U8916 (N_8916,N_6882,N_6120);
nor U8917 (N_8917,N_7294,N_6644);
or U8918 (N_8918,N_6565,N_6188);
and U8919 (N_8919,N_6618,N_6312);
or U8920 (N_8920,N_6272,N_6344);
nor U8921 (N_8921,N_6150,N_6021);
or U8922 (N_8922,N_6910,N_6380);
or U8923 (N_8923,N_7212,N_6440);
nand U8924 (N_8924,N_6702,N_6567);
nand U8925 (N_8925,N_6331,N_6774);
and U8926 (N_8926,N_6392,N_6605);
nand U8927 (N_8927,N_7152,N_7267);
nand U8928 (N_8928,N_6649,N_7033);
xnor U8929 (N_8929,N_6710,N_6252);
nand U8930 (N_8930,N_6468,N_7229);
and U8931 (N_8931,N_7354,N_6559);
nor U8932 (N_8932,N_7033,N_6690);
xor U8933 (N_8933,N_6182,N_7113);
or U8934 (N_8934,N_6217,N_7489);
and U8935 (N_8935,N_6541,N_6987);
and U8936 (N_8936,N_6098,N_7273);
nor U8937 (N_8937,N_7011,N_6649);
xnor U8938 (N_8938,N_6320,N_7184);
nand U8939 (N_8939,N_7078,N_6848);
nor U8940 (N_8940,N_7040,N_6633);
and U8941 (N_8941,N_6520,N_7259);
nand U8942 (N_8942,N_6418,N_6746);
nand U8943 (N_8943,N_7134,N_6049);
and U8944 (N_8944,N_7413,N_6948);
xnor U8945 (N_8945,N_6054,N_6889);
and U8946 (N_8946,N_6897,N_7196);
nand U8947 (N_8947,N_6399,N_7478);
and U8948 (N_8948,N_6127,N_7138);
nor U8949 (N_8949,N_6098,N_7100);
nor U8950 (N_8950,N_6491,N_6089);
or U8951 (N_8951,N_6220,N_7068);
nor U8952 (N_8952,N_6566,N_6951);
nor U8953 (N_8953,N_7385,N_6127);
nor U8954 (N_8954,N_6847,N_7266);
nand U8955 (N_8955,N_6212,N_7246);
and U8956 (N_8956,N_7172,N_7367);
nor U8957 (N_8957,N_7091,N_6241);
and U8958 (N_8958,N_6468,N_6355);
nor U8959 (N_8959,N_6548,N_6068);
xor U8960 (N_8960,N_7054,N_6427);
or U8961 (N_8961,N_6042,N_6993);
xor U8962 (N_8962,N_6653,N_7462);
and U8963 (N_8963,N_6378,N_6994);
or U8964 (N_8964,N_6477,N_6655);
nor U8965 (N_8965,N_6037,N_6728);
nor U8966 (N_8966,N_6308,N_6754);
and U8967 (N_8967,N_6724,N_6256);
nor U8968 (N_8968,N_6457,N_6580);
nand U8969 (N_8969,N_7059,N_6187);
or U8970 (N_8970,N_6731,N_7485);
or U8971 (N_8971,N_7290,N_6078);
or U8972 (N_8972,N_6820,N_6989);
nand U8973 (N_8973,N_6199,N_6020);
nor U8974 (N_8974,N_7234,N_7336);
nor U8975 (N_8975,N_6398,N_6930);
and U8976 (N_8976,N_6756,N_7403);
nor U8977 (N_8977,N_7034,N_7400);
or U8978 (N_8978,N_6598,N_7100);
or U8979 (N_8979,N_6714,N_6030);
nor U8980 (N_8980,N_6931,N_7360);
nor U8981 (N_8981,N_7447,N_6653);
or U8982 (N_8982,N_7450,N_6392);
nand U8983 (N_8983,N_6336,N_6991);
nand U8984 (N_8984,N_7306,N_7004);
and U8985 (N_8985,N_6742,N_6287);
nor U8986 (N_8986,N_7020,N_6963);
nor U8987 (N_8987,N_6419,N_7312);
and U8988 (N_8988,N_7284,N_6240);
and U8989 (N_8989,N_6748,N_6155);
nand U8990 (N_8990,N_7479,N_6998);
or U8991 (N_8991,N_7125,N_6721);
and U8992 (N_8992,N_6069,N_6977);
or U8993 (N_8993,N_7433,N_6476);
and U8994 (N_8994,N_6539,N_7178);
or U8995 (N_8995,N_6294,N_7280);
xor U8996 (N_8996,N_6690,N_6778);
or U8997 (N_8997,N_6534,N_7428);
nand U8998 (N_8998,N_6271,N_7036);
nor U8999 (N_8999,N_6638,N_6993);
or U9000 (N_9000,N_8677,N_7978);
nand U9001 (N_9001,N_7989,N_8909);
xor U9002 (N_9002,N_8838,N_8679);
nand U9003 (N_9003,N_8334,N_8456);
or U9004 (N_9004,N_8697,N_7905);
or U9005 (N_9005,N_8702,N_7760);
xor U9006 (N_9006,N_7911,N_8524);
xor U9007 (N_9007,N_8671,N_8757);
or U9008 (N_9008,N_8703,N_8799);
or U9009 (N_9009,N_7998,N_8045);
nand U9010 (N_9010,N_7930,N_7832);
nand U9011 (N_9011,N_8234,N_7710);
nand U9012 (N_9012,N_8177,N_8607);
or U9013 (N_9013,N_7879,N_8304);
nand U9014 (N_9014,N_8988,N_8758);
nor U9015 (N_9015,N_8765,N_8180);
and U9016 (N_9016,N_8257,N_8565);
nand U9017 (N_9017,N_7561,N_7650);
or U9018 (N_9018,N_8483,N_8916);
and U9019 (N_9019,N_7637,N_8961);
and U9020 (N_9020,N_8638,N_7606);
or U9021 (N_9021,N_7762,N_8754);
nor U9022 (N_9022,N_8720,N_8984);
and U9023 (N_9023,N_8171,N_8642);
or U9024 (N_9024,N_8135,N_7822);
or U9025 (N_9025,N_8778,N_7805);
nor U9026 (N_9026,N_8481,N_8381);
or U9027 (N_9027,N_8212,N_8733);
or U9028 (N_9028,N_7546,N_8827);
nor U9029 (N_9029,N_7575,N_7607);
nor U9030 (N_9030,N_8943,N_8400);
nor U9031 (N_9031,N_8359,N_8536);
nand U9032 (N_9032,N_8709,N_8455);
nand U9033 (N_9033,N_8141,N_8725);
nand U9034 (N_9034,N_8941,N_7816);
nand U9035 (N_9035,N_8581,N_8611);
or U9036 (N_9036,N_7746,N_8477);
and U9037 (N_9037,N_8914,N_7984);
or U9038 (N_9038,N_7956,N_7541);
or U9039 (N_9039,N_8841,N_8219);
nor U9040 (N_9040,N_7712,N_8098);
nor U9041 (N_9041,N_8661,N_8705);
and U9042 (N_9042,N_8589,N_8884);
nor U9043 (N_9043,N_8734,N_8378);
nor U9044 (N_9044,N_7971,N_7960);
nand U9045 (N_9045,N_8223,N_7918);
xnor U9046 (N_9046,N_7671,N_8208);
nor U9047 (N_9047,N_8227,N_8615);
nor U9048 (N_9048,N_7661,N_7646);
and U9049 (N_9049,N_8279,N_7724);
and U9050 (N_9050,N_7864,N_8357);
xnor U9051 (N_9051,N_7522,N_8361);
or U9052 (N_9052,N_7949,N_7627);
and U9053 (N_9053,N_8463,N_8544);
and U9054 (N_9054,N_7632,N_8789);
or U9055 (N_9055,N_8881,N_8922);
nor U9056 (N_9056,N_8667,N_8094);
and U9057 (N_9057,N_7898,N_7631);
and U9058 (N_9058,N_8618,N_8830);
nor U9059 (N_9059,N_7991,N_8383);
nor U9060 (N_9060,N_8823,N_8440);
nand U9061 (N_9061,N_7969,N_8254);
nor U9062 (N_9062,N_8067,N_8639);
xor U9063 (N_9063,N_7741,N_8306);
nor U9064 (N_9064,N_8179,N_8230);
xnor U9065 (N_9065,N_8027,N_8132);
nand U9066 (N_9066,N_8151,N_7518);
or U9067 (N_9067,N_8103,N_7626);
xnor U9068 (N_9068,N_8111,N_8484);
or U9069 (N_9069,N_7686,N_8319);
nor U9070 (N_9070,N_7802,N_8023);
or U9071 (N_9071,N_8732,N_8728);
nand U9072 (N_9072,N_8547,N_8576);
or U9073 (N_9073,N_7828,N_7700);
nand U9074 (N_9074,N_8968,N_8727);
and U9075 (N_9075,N_7558,N_8805);
nand U9076 (N_9076,N_7769,N_8902);
or U9077 (N_9077,N_7945,N_7917);
or U9078 (N_9078,N_8039,N_7555);
and U9079 (N_9079,N_8476,N_8056);
nand U9080 (N_9080,N_7619,N_7734);
or U9081 (N_9081,N_7653,N_8253);
and U9082 (N_9082,N_8859,N_8942);
or U9083 (N_9083,N_8967,N_7564);
nand U9084 (N_9084,N_7778,N_8731);
nor U9085 (N_9085,N_7549,N_8612);
or U9086 (N_9086,N_7537,N_8165);
and U9087 (N_9087,N_8529,N_8152);
and U9088 (N_9088,N_7994,N_8118);
nand U9089 (N_9089,N_8566,N_8299);
and U9090 (N_9090,N_7657,N_8181);
and U9091 (N_9091,N_8489,N_8123);
or U9092 (N_9092,N_8788,N_8043);
and U9093 (N_9093,N_8211,N_8792);
nand U9094 (N_9094,N_7780,N_8974);
nand U9095 (N_9095,N_7885,N_7732);
nor U9096 (N_9096,N_8284,N_8164);
and U9097 (N_9097,N_7744,N_8995);
nand U9098 (N_9098,N_7841,N_7717);
xor U9099 (N_9099,N_8715,N_7967);
nand U9100 (N_9100,N_8794,N_8991);
nor U9101 (N_9101,N_8110,N_8289);
nor U9102 (N_9102,N_7526,N_8194);
nand U9103 (N_9103,N_8136,N_8882);
or U9104 (N_9104,N_8201,N_8466);
nor U9105 (N_9105,N_8250,N_7784);
nor U9106 (N_9106,N_7533,N_8911);
xnor U9107 (N_9107,N_8206,N_8633);
nor U9108 (N_9108,N_7892,N_7829);
nor U9109 (N_9109,N_8142,N_8224);
nand U9110 (N_9110,N_7603,N_7757);
nand U9111 (N_9111,N_7512,N_8225);
or U9112 (N_9112,N_7691,N_8480);
and U9113 (N_9113,N_8663,N_8447);
nand U9114 (N_9114,N_8325,N_8949);
nand U9115 (N_9115,N_7853,N_8444);
nand U9116 (N_9116,N_7635,N_7500);
xor U9117 (N_9117,N_8680,N_7781);
or U9118 (N_9118,N_8798,N_8915);
and U9119 (N_9119,N_7617,N_8760);
xnor U9120 (N_9120,N_7770,N_8590);
nand U9121 (N_9121,N_8519,N_8651);
nand U9122 (N_9122,N_7980,N_8600);
nor U9123 (N_9123,N_7662,N_8109);
xnor U9124 (N_9124,N_8232,N_8843);
nand U9125 (N_9125,N_8129,N_8150);
and U9126 (N_9126,N_7854,N_7654);
nor U9127 (N_9127,N_7753,N_8331);
nor U9128 (N_9128,N_8775,N_8835);
and U9129 (N_9129,N_8269,N_8005);
nor U9130 (N_9130,N_7915,N_8393);
or U9131 (N_9131,N_7525,N_7697);
nand U9132 (N_9132,N_8948,N_7756);
nand U9133 (N_9133,N_7752,N_8312);
nand U9134 (N_9134,N_8233,N_7833);
or U9135 (N_9135,N_7877,N_7842);
nor U9136 (N_9136,N_8527,N_8271);
and U9137 (N_9137,N_7993,N_7620);
nor U9138 (N_9138,N_8176,N_8928);
nand U9139 (N_9139,N_8428,N_8817);
nor U9140 (N_9140,N_8097,N_8953);
nor U9141 (N_9141,N_7723,N_7594);
nor U9142 (N_9142,N_8749,N_8903);
and U9143 (N_9143,N_8630,N_8218);
or U9144 (N_9144,N_7882,N_8356);
and U9145 (N_9145,N_7645,N_8351);
nor U9146 (N_9146,N_7502,N_8926);
xnor U9147 (N_9147,N_7869,N_8376);
and U9148 (N_9148,N_8912,N_8921);
and U9149 (N_9149,N_8239,N_8235);
nor U9150 (N_9150,N_8867,N_8753);
and U9151 (N_9151,N_8585,N_8837);
nand U9152 (N_9152,N_8657,N_7649);
or U9153 (N_9153,N_7665,N_8931);
nor U9154 (N_9154,N_8365,N_8090);
or U9155 (N_9155,N_8857,N_8530);
nor U9156 (N_9156,N_8982,N_7601);
or U9157 (N_9157,N_7644,N_8354);
and U9158 (N_9158,N_7939,N_7571);
and U9159 (N_9159,N_8310,N_8917);
and U9160 (N_9160,N_7677,N_8465);
and U9161 (N_9161,N_8115,N_8127);
or U9162 (N_9162,N_8736,N_8072);
or U9163 (N_9163,N_8836,N_7941);
nand U9164 (N_9164,N_8471,N_7559);
and U9165 (N_9165,N_8070,N_8300);
and U9166 (N_9166,N_8787,N_7944);
nor U9167 (N_9167,N_8012,N_7576);
nor U9168 (N_9168,N_7729,N_8384);
and U9169 (N_9169,N_8082,N_8971);
nand U9170 (N_9170,N_8845,N_7641);
nor U9171 (N_9171,N_8932,N_7593);
nor U9172 (N_9172,N_8852,N_8553);
or U9173 (N_9173,N_7718,N_8691);
nor U9174 (N_9174,N_8644,N_8617);
xnor U9175 (N_9175,N_8091,N_8445);
nand U9176 (N_9176,N_7706,N_8018);
or U9177 (N_9177,N_8498,N_8797);
nor U9178 (N_9178,N_8419,N_8486);
and U9179 (N_9179,N_8923,N_8874);
or U9180 (N_9180,N_7873,N_7777);
nand U9181 (N_9181,N_8375,N_8429);
nor U9182 (N_9182,N_8810,N_8640);
or U9183 (N_9183,N_7859,N_8598);
xnor U9184 (N_9184,N_8495,N_8759);
nor U9185 (N_9185,N_8369,N_8128);
or U9186 (N_9186,N_8636,N_8020);
and U9187 (N_9187,N_8997,N_7615);
nor U9188 (N_9188,N_7974,N_8762);
and U9189 (N_9189,N_7800,N_7690);
and U9190 (N_9190,N_8270,N_8950);
and U9191 (N_9191,N_7584,N_8050);
and U9192 (N_9192,N_8048,N_8105);
nor U9193 (N_9193,N_8267,N_8552);
and U9194 (N_9194,N_8689,N_7895);
or U9195 (N_9195,N_8578,N_8034);
or U9196 (N_9196,N_8113,N_7764);
and U9197 (N_9197,N_8341,N_8220);
nand U9198 (N_9198,N_8349,N_7912);
and U9199 (N_9199,N_7680,N_7768);
or U9200 (N_9200,N_7600,N_7733);
nor U9201 (N_9201,N_8302,N_7588);
xnor U9202 (N_9202,N_8674,N_8573);
and U9203 (N_9203,N_7609,N_8761);
or U9204 (N_9204,N_8947,N_8117);
and U9205 (N_9205,N_7742,N_8044);
or U9206 (N_9206,N_8277,N_8170);
and U9207 (N_9207,N_8739,N_7887);
or U9208 (N_9208,N_7605,N_8610);
and U9209 (N_9209,N_8907,N_8621);
nor U9210 (N_9210,N_8398,N_8275);
nand U9211 (N_9211,N_8643,N_7825);
xor U9212 (N_9212,N_7846,N_8575);
and U9213 (N_9213,N_7904,N_8894);
and U9214 (N_9214,N_8457,N_7596);
nand U9215 (N_9215,N_7808,N_8723);
nand U9216 (N_9216,N_7580,N_8266);
nor U9217 (N_9217,N_7738,N_8174);
nor U9218 (N_9218,N_7516,N_8764);
nand U9219 (N_9219,N_8983,N_8287);
or U9220 (N_9220,N_8930,N_8729);
nand U9221 (N_9221,N_8404,N_8475);
nor U9222 (N_9222,N_8200,N_8646);
or U9223 (N_9223,N_8685,N_8675);
nand U9224 (N_9224,N_8078,N_8352);
or U9225 (N_9225,N_8714,N_8972);
xor U9226 (N_9226,N_7625,N_8162);
or U9227 (N_9227,N_8293,N_8478);
and U9228 (N_9228,N_7783,N_8274);
nor U9229 (N_9229,N_8454,N_7501);
nor U9230 (N_9230,N_7914,N_8467);
nand U9231 (N_9231,N_8583,N_8358);
nor U9232 (N_9232,N_8395,N_8877);
or U9233 (N_9233,N_8379,N_8185);
or U9234 (N_9234,N_8172,N_8488);
nand U9235 (N_9235,N_8410,N_8425);
nand U9236 (N_9236,N_8790,N_8541);
nand U9237 (N_9237,N_8055,N_8169);
and U9238 (N_9238,N_8957,N_8460);
and U9239 (N_9239,N_8330,N_8413);
nor U9240 (N_9240,N_8965,N_8672);
nand U9241 (N_9241,N_8970,N_8847);
nor U9242 (N_9242,N_8084,N_8580);
xnor U9243 (N_9243,N_8920,N_7868);
and U9244 (N_9244,N_8592,N_8140);
and U9245 (N_9245,N_8493,N_8409);
and U9246 (N_9246,N_7581,N_7880);
nor U9247 (N_9247,N_8603,N_8442);
nor U9248 (N_9248,N_7557,N_8510);
and U9249 (N_9249,N_8695,N_8851);
xnor U9250 (N_9250,N_7683,N_8015);
nor U9251 (N_9251,N_8831,N_8624);
nand U9252 (N_9252,N_7623,N_7684);
nand U9253 (N_9253,N_7772,N_7527);
or U9254 (N_9254,N_7597,N_8614);
nor U9255 (N_9255,N_8872,N_7611);
nor U9256 (N_9256,N_8973,N_8936);
nor U9257 (N_9257,N_8106,N_8594);
and U9258 (N_9258,N_8768,N_8774);
or U9259 (N_9259,N_8255,N_7651);
or U9260 (N_9260,N_8060,N_8355);
nand U9261 (N_9261,N_8556,N_8243);
or U9262 (N_9262,N_8588,N_7672);
nor U9263 (N_9263,N_8286,N_7938);
xor U9264 (N_9264,N_8013,N_7867);
nand U9265 (N_9265,N_8153,N_8522);
nand U9266 (N_9266,N_8137,N_8245);
nor U9267 (N_9267,N_8101,N_8411);
and U9268 (N_9268,N_8335,N_7910);
xnor U9269 (N_9269,N_7679,N_8199);
nor U9270 (N_9270,N_8386,N_8030);
nor U9271 (N_9271,N_7595,N_8840);
xor U9272 (N_9272,N_8403,N_8708);
nand U9273 (N_9273,N_8508,N_8517);
and U9274 (N_9274,N_7883,N_8821);
and U9275 (N_9275,N_7586,N_7530);
nand U9276 (N_9276,N_8875,N_8721);
or U9277 (N_9277,N_8433,N_8571);
or U9278 (N_9278,N_7634,N_8904);
nand U9279 (N_9279,N_8858,N_8025);
nand U9280 (N_9280,N_8423,N_8616);
nor U9281 (N_9281,N_8550,N_7705);
nor U9282 (N_9282,N_8333,N_7639);
xnor U9283 (N_9283,N_8771,N_8999);
nand U9284 (N_9284,N_8315,N_8684);
or U9285 (N_9285,N_7692,N_8593);
or U9286 (N_9286,N_8626,N_8119);
nand U9287 (N_9287,N_7797,N_8564);
nor U9288 (N_9288,N_8345,N_8427);
or U9289 (N_9289,N_8148,N_8748);
and U9290 (N_9290,N_8237,N_8769);
and U9291 (N_9291,N_8276,N_7668);
and U9292 (N_9292,N_8570,N_8554);
and U9293 (N_9293,N_8742,N_7920);
and U9294 (N_9294,N_8869,N_8131);
or U9295 (N_9295,N_8855,N_7608);
nand U9296 (N_9296,N_7509,N_8264);
nor U9297 (N_9297,N_8766,N_8301);
nor U9298 (N_9298,N_8818,N_8149);
nor U9299 (N_9299,N_8421,N_8462);
or U9300 (N_9300,N_8184,N_8628);
xor U9301 (N_9301,N_8558,N_8813);
nand U9302 (N_9302,N_8374,N_7888);
or U9303 (N_9303,N_8139,N_8548);
nand U9304 (N_9304,N_8503,N_7714);
nor U9305 (N_9305,N_8856,N_8743);
xnor U9306 (N_9306,N_7795,N_7536);
or U9307 (N_9307,N_8625,N_8202);
and U9308 (N_9308,N_7973,N_8210);
xor U9309 (N_9309,N_8196,N_8978);
and U9310 (N_9310,N_8776,N_8168);
nor U9311 (N_9311,N_8897,N_8088);
and U9312 (N_9312,N_8468,N_8686);
or U9313 (N_9313,N_7618,N_8247);
and U9314 (N_9314,N_7730,N_8108);
nand U9315 (N_9315,N_8215,N_8938);
nor U9316 (N_9316,N_7809,N_8832);
nand U9317 (N_9317,N_8133,N_8125);
nor U9318 (N_9318,N_8735,N_8415);
and U9319 (N_9319,N_8124,N_8143);
and U9320 (N_9320,N_8022,N_7852);
nor U9321 (N_9321,N_8058,N_7936);
or U9322 (N_9322,N_8815,N_8826);
or U9323 (N_9323,N_8010,N_8291);
or U9324 (N_9324,N_7587,N_7702);
nand U9325 (N_9325,N_7970,N_7823);
nand U9326 (N_9326,N_7716,N_7804);
or U9327 (N_9327,N_7874,N_8883);
or U9328 (N_9328,N_7891,N_7897);
xnor U9329 (N_9329,N_8619,N_7819);
nand U9330 (N_9330,N_8112,N_8864);
and U9331 (N_9331,N_8298,N_8311);
nor U9332 (N_9332,N_8763,N_7574);
nor U9333 (N_9333,N_8041,N_7943);
xor U9334 (N_9334,N_8673,N_8586);
xnor U9335 (N_9335,N_8320,N_7789);
and U9336 (N_9336,N_8839,N_8795);
nand U9337 (N_9337,N_7827,N_8051);
xnor U9338 (N_9338,N_8996,N_8104);
and U9339 (N_9339,N_8648,N_8577);
xnor U9340 (N_9340,N_8525,N_8157);
nor U9341 (N_9341,N_7511,N_7831);
nand U9342 (N_9342,N_8652,N_8074);
nor U9343 (N_9343,N_8551,N_8087);
or U9344 (N_9344,N_8854,N_7708);
xor U9345 (N_9345,N_8371,N_8887);
nor U9346 (N_9346,N_7515,N_8649);
and U9347 (N_9347,N_7886,N_8669);
or U9348 (N_9348,N_8035,N_8077);
or U9349 (N_9349,N_8308,N_8102);
and U9350 (N_9350,N_8407,N_7624);
and U9351 (N_9351,N_8579,N_7834);
nor U9352 (N_9352,N_8891,N_8167);
nor U9353 (N_9353,N_8509,N_8756);
nand U9354 (N_9354,N_8863,N_7982);
and U9355 (N_9355,N_8500,N_7896);
nor U9356 (N_9356,N_8944,N_7929);
or U9357 (N_9357,N_8737,N_8523);
nand U9358 (N_9358,N_8173,N_8303);
nor U9359 (N_9359,N_7689,N_7591);
or U9360 (N_9360,N_8719,N_8231);
and U9361 (N_9361,N_7582,N_7547);
nor U9362 (N_9362,N_8008,N_7849);
or U9363 (N_9363,N_7957,N_8038);
nor U9364 (N_9364,N_8750,N_8712);
nor U9365 (N_9365,N_8353,N_8314);
and U9366 (N_9366,N_8449,N_8017);
or U9367 (N_9367,N_7871,N_8079);
and U9368 (N_9368,N_7847,N_8099);
nor U9369 (N_9369,N_8962,N_8402);
or U9370 (N_9370,N_8741,N_7721);
nand U9371 (N_9371,N_7745,N_7862);
xnor U9372 (N_9372,N_8326,N_7935);
nand U9373 (N_9373,N_8747,N_7775);
or U9374 (N_9374,N_8432,N_8392);
xnor U9375 (N_9375,N_8542,N_8681);
and U9376 (N_9376,N_7709,N_8031);
nor U9377 (N_9377,N_7932,N_8808);
nand U9378 (N_9378,N_8706,N_8704);
and U9379 (N_9379,N_7676,N_7545);
or U9380 (N_9380,N_7585,N_8226);
nand U9381 (N_9381,N_7556,N_7663);
or U9382 (N_9382,N_8693,N_7505);
nand U9383 (N_9383,N_8144,N_7563);
and U9384 (N_9384,N_7965,N_8929);
nand U9385 (N_9385,N_8338,N_7807);
or U9386 (N_9386,N_8512,N_7985);
and U9387 (N_9387,N_7630,N_8666);
or U9388 (N_9388,N_8898,N_8065);
nand U9389 (N_9389,N_8390,N_8385);
and U9390 (N_9390,N_7782,N_8587);
nor U9391 (N_9391,N_8406,N_7739);
and U9392 (N_9392,N_8388,N_8925);
or U9393 (N_9393,N_8986,N_8107);
nand U9394 (N_9394,N_8324,N_8698);
xnor U9395 (N_9395,N_8958,N_8849);
or U9396 (N_9396,N_8412,N_8183);
or U9397 (N_9397,N_8464,N_8985);
and U9398 (N_9398,N_8900,N_8833);
nand U9399 (N_9399,N_8420,N_7667);
nand U9400 (N_9400,N_7899,N_7798);
nor U9401 (N_9401,N_8062,N_7952);
or U9402 (N_9402,N_8182,N_7693);
or U9403 (N_9403,N_8258,N_7664);
nor U9404 (N_9404,N_8535,N_7785);
nand U9405 (N_9405,N_7513,N_8373);
nand U9406 (N_9406,N_8888,N_8871);
xor U9407 (N_9407,N_7790,N_7902);
nand U9408 (N_9408,N_7903,N_7979);
and U9409 (N_9409,N_7583,N_7726);
nand U9410 (N_9410,N_8155,N_8976);
or U9411 (N_9411,N_8595,N_7719);
and U9412 (N_9412,N_8811,N_8138);
nand U9413 (N_9413,N_7698,N_7817);
xnor U9414 (N_9414,N_7573,N_8809);
or U9415 (N_9415,N_7507,N_8453);
and U9416 (N_9416,N_7538,N_8539);
nor U9417 (N_9417,N_8297,N_7670);
nand U9418 (N_9418,N_7755,N_7843);
nor U9419 (N_9419,N_7673,N_8901);
or U9420 (N_9420,N_8309,N_8676);
nor U9421 (N_9421,N_8229,N_8052);
nand U9422 (N_9422,N_8417,N_8399);
nor U9423 (N_9423,N_8418,N_8337);
nor U9424 (N_9424,N_7577,N_8473);
or U9425 (N_9425,N_8664,N_8634);
xnor U9426 (N_9426,N_8853,N_7925);
nand U9427 (N_9427,N_8213,N_8092);
nor U9428 (N_9428,N_7514,N_8006);
xor U9429 (N_9429,N_7906,N_7751);
or U9430 (N_9430,N_7870,N_7953);
nand U9431 (N_9431,N_8204,N_8670);
nand U9432 (N_9432,N_8387,N_8033);
or U9433 (N_9433,N_7942,N_8631);
xor U9434 (N_9434,N_8273,N_8003);
and U9435 (N_9435,N_8846,N_7821);
or U9436 (N_9436,N_8609,N_8469);
nor U9437 (N_9437,N_8599,N_8307);
nand U9438 (N_9438,N_8613,N_8222);
xnor U9439 (N_9439,N_8694,N_8130);
nor U9440 (N_9440,N_8933,N_8120);
xor U9441 (N_9441,N_8975,N_8019);
nor U9442 (N_9442,N_8802,N_8401);
nor U9443 (N_9443,N_8977,N_7535);
nor U9444 (N_9444,N_8145,N_7848);
or U9445 (N_9445,N_8063,N_8574);
nand U9446 (N_9446,N_7928,N_7983);
xnor U9447 (N_9447,N_8037,N_8927);
and U9448 (N_9448,N_7612,N_7958);
or U9449 (N_9449,N_7565,N_8779);
or U9450 (N_9450,N_8288,N_8531);
nor U9451 (N_9451,N_8540,N_8193);
nand U9452 (N_9452,N_7579,N_7681);
and U9453 (N_9453,N_8740,N_8781);
nor U9454 (N_9454,N_7999,N_8414);
or U9455 (N_9455,N_7740,N_8436);
and U9456 (N_9456,N_8203,N_7523);
nor U9457 (N_9457,N_7722,N_7997);
nand U9458 (N_9458,N_8641,N_8394);
xnor U9459 (N_9459,N_8717,N_8683);
nor U9460 (N_9460,N_8545,N_8238);
and U9461 (N_9461,N_7539,N_8437);
xnor U9462 (N_9462,N_8040,N_8629);
xor U9463 (N_9463,N_7810,N_8435);
and U9464 (N_9464,N_8336,N_8434);
nand U9465 (N_9465,N_7976,N_7735);
nor U9466 (N_9466,N_7858,N_8175);
nand U9467 (N_9467,N_8268,N_7933);
nand U9468 (N_9468,N_8507,N_8492);
nor U9469 (N_9469,N_8520,N_8952);
or U9470 (N_9470,N_7963,N_8687);
or U9471 (N_9471,N_8259,N_7959);
xnor U9472 (N_9472,N_8602,N_8328);
nor U9473 (N_9473,N_7695,N_7647);
nor U9474 (N_9474,N_8147,N_8770);
nor U9475 (N_9475,N_7727,N_7946);
or U9476 (N_9476,N_8561,N_8458);
nor U9477 (N_9477,N_8793,N_7567);
nor U9478 (N_9478,N_7633,N_8688);
and U9479 (N_9479,N_8007,N_7961);
nand U9480 (N_9480,N_8662,N_8647);
nor U9481 (N_9481,N_7643,N_8391);
nand U9482 (N_9482,N_7658,N_7796);
or U9483 (N_9483,N_8004,N_8470);
xnor U9484 (N_9484,N_8890,N_8606);
and U9485 (N_9485,N_8236,N_7992);
xnor U9486 (N_9486,N_8377,N_8713);
nand U9487 (N_9487,N_7972,N_8597);
xnor U9488 (N_9488,N_8924,N_8046);
nor U9489 (N_9489,N_8880,N_8623);
and U9490 (N_9490,N_7884,N_8389);
or U9491 (N_9491,N_8446,N_8886);
nor U9492 (N_9492,N_8342,N_8514);
nor U9493 (N_9493,N_8896,N_7771);
nand U9494 (N_9494,N_8710,N_8755);
or U9495 (N_9495,N_7678,N_7687);
nor U9496 (N_9496,N_7720,N_8511);
nor U9497 (N_9497,N_7765,N_8494);
nor U9498 (N_9498,N_8521,N_7728);
or U9499 (N_9499,N_7750,N_7614);
nand U9500 (N_9500,N_8866,N_7642);
and U9501 (N_9501,N_8360,N_8159);
and U9502 (N_9502,N_8814,N_8262);
or U9503 (N_9503,N_7844,N_7531);
nand U9504 (N_9504,N_7551,N_7590);
nand U9505 (N_9505,N_8584,N_8772);
and U9506 (N_9506,N_8563,N_8682);
xnor U9507 (N_9507,N_8186,N_8317);
nor U9508 (N_9508,N_8622,N_8767);
nor U9509 (N_9509,N_7532,N_7799);
or U9510 (N_9510,N_8370,N_7866);
nand U9511 (N_9511,N_8828,N_7836);
and U9512 (N_9512,N_8207,N_8217);
nand U9513 (N_9513,N_7774,N_7995);
nor U9514 (N_9514,N_8026,N_7543);
xor U9515 (N_9515,N_7975,N_7826);
xnor U9516 (N_9516,N_7907,N_8878);
and U9517 (N_9517,N_8549,N_8653);
xor U9518 (N_9518,N_8246,N_7704);
or U9519 (N_9519,N_7703,N_7801);
and U9520 (N_9520,N_8295,N_8472);
or U9521 (N_9521,N_8850,N_7950);
and U9522 (N_9522,N_8513,N_8221);
nand U9523 (N_9523,N_8989,N_7747);
nand U9524 (N_9524,N_8028,N_7863);
or U9525 (N_9525,N_8533,N_7737);
or U9526 (N_9526,N_8959,N_8343);
nor U9527 (N_9527,N_7921,N_7812);
xnor U9528 (N_9528,N_8981,N_8656);
nor U9529 (N_9529,N_7968,N_8296);
and U9530 (N_9530,N_8501,N_8431);
nor U9531 (N_9531,N_7793,N_8195);
nand U9532 (N_9532,N_7763,N_7955);
and U9533 (N_9533,N_7659,N_8318);
nor U9534 (N_9534,N_8085,N_7715);
and U9535 (N_9535,N_8865,N_8568);
or U9536 (N_9536,N_8591,N_8908);
or U9537 (N_9537,N_8627,N_8724);
nor U9538 (N_9538,N_7566,N_7621);
or U9539 (N_9539,N_7894,N_8408);
nor U9540 (N_9540,N_8868,N_8348);
or U9541 (N_9541,N_7977,N_8879);
nor U9542 (N_9542,N_8860,N_8668);
nand U9543 (N_9543,N_8987,N_8745);
and U9544 (N_9544,N_8339,N_8001);
and U9545 (N_9545,N_8346,N_8047);
nor U9546 (N_9546,N_8479,N_8969);
nor U9547 (N_9547,N_7948,N_7916);
or U9548 (N_9548,N_8362,N_8448);
xor U9549 (N_9549,N_7856,N_8504);
nand U9550 (N_9550,N_8786,N_7688);
or U9551 (N_9551,N_8485,N_8963);
nand U9552 (N_9552,N_7540,N_8516);
nand U9553 (N_9553,N_8156,N_8939);
nand U9554 (N_9554,N_7508,N_8899);
and U9555 (N_9555,N_8780,N_7510);
and U9556 (N_9556,N_7924,N_7570);
or U9557 (N_9557,N_8819,N_8260);
nor U9558 (N_9558,N_7987,N_8178);
and U9559 (N_9559,N_8526,N_8885);
nor U9560 (N_9560,N_8282,N_8011);
nand U9561 (N_9561,N_7743,N_7875);
and U9562 (N_9562,N_7840,N_8491);
and U9563 (N_9563,N_7544,N_8800);
nor U9564 (N_9564,N_8146,N_8189);
nor U9565 (N_9565,N_8057,N_8773);
or U9566 (N_9566,N_8347,N_7830);
or U9567 (N_9567,N_7542,N_8042);
nor U9568 (N_9568,N_8073,N_8265);
nor U9569 (N_9569,N_7996,N_8608);
nand U9570 (N_9570,N_8187,N_7937);
xor U9571 (N_9571,N_7981,N_7922);
and U9572 (N_9572,N_8946,N_8848);
nand U9573 (N_9573,N_7675,N_8696);
nand U9574 (N_9574,N_7954,N_8744);
and U9575 (N_9575,N_8834,N_7813);
xnor U9576 (N_9576,N_7934,N_8816);
or U9577 (N_9577,N_8956,N_8114);
nor U9578 (N_9578,N_8659,N_7776);
and U9579 (N_9579,N_7865,N_8405);
or U9580 (N_9580,N_7749,N_8021);
xnor U9581 (N_9581,N_8126,N_8893);
nand U9582 (N_9582,N_8054,N_8474);
nand U9583 (N_9583,N_8241,N_7568);
nor U9584 (N_9584,N_8191,N_8784);
or U9585 (N_9585,N_8080,N_8380);
nor U9586 (N_9586,N_7638,N_7521);
and U9587 (N_9587,N_8650,N_8160);
nand U9588 (N_9588,N_8635,N_8283);
nor U9589 (N_9589,N_8016,N_8014);
nor U9590 (N_9590,N_8992,N_8998);
xor U9591 (N_9591,N_7725,N_7940);
nor U9592 (N_9592,N_8954,N_8482);
nand U9593 (N_9593,N_7900,N_7919);
nand U9594 (N_9594,N_8327,N_7589);
xor U9595 (N_9595,N_7855,N_8844);
xnor U9596 (N_9596,N_8332,N_8862);
nor U9597 (N_9597,N_7773,N_8081);
nor U9598 (N_9598,N_8935,N_8032);
nor U9599 (N_9599,N_7602,N_8572);
nor U9600 (N_9600,N_8198,N_7592);
nand U9601 (N_9601,N_8261,N_7820);
nand U9602 (N_9602,N_8555,N_7554);
and U9603 (N_9603,N_8502,N_7881);
xnor U9604 (N_9604,N_7947,N_8919);
or U9605 (N_9605,N_7660,N_8256);
nor U9606 (N_9606,N_8121,N_8278);
nand U9607 (N_9607,N_8543,N_7872);
nand U9608 (N_9608,N_8538,N_8228);
and U9609 (N_9609,N_8316,N_8945);
nor U9610 (N_9610,N_8979,N_7529);
or U9611 (N_9611,N_7966,N_8163);
nand U9612 (N_9612,N_8562,N_8518);
xor U9613 (N_9613,N_7767,N_8604);
nor U9614 (N_9614,N_7988,N_8892);
and U9615 (N_9615,N_8397,N_8461);
nand U9616 (N_9616,N_7748,N_7779);
nand U9617 (N_9617,N_8438,N_7517);
and U9618 (N_9618,N_8560,N_8738);
nand U9619 (N_9619,N_8000,N_7713);
and U9620 (N_9620,N_7598,N_7699);
xnor U9621 (N_9621,N_7908,N_8251);
nor U9622 (N_9622,N_8722,N_8582);
nand U9623 (N_9623,N_7791,N_8083);
nor U9624 (N_9624,N_7622,N_7964);
nor U9625 (N_9625,N_8918,N_8701);
nand U9626 (N_9626,N_7669,N_8870);
or U9627 (N_9627,N_7506,N_8829);
or U9628 (N_9628,N_8059,N_8645);
nor U9629 (N_9629,N_8824,N_8430);
or U9630 (N_9630,N_7562,N_8752);
nor U9631 (N_9631,N_8537,N_7550);
nand U9632 (N_9632,N_8158,N_8532);
or U9633 (N_9633,N_8340,N_8730);
and U9634 (N_9634,N_7835,N_8116);
and U9635 (N_9635,N_8329,N_8906);
nor U9636 (N_9636,N_8487,N_8692);
or U9637 (N_9637,N_8980,N_8188);
or U9638 (N_9638,N_8796,N_8096);
and U9639 (N_9639,N_8422,N_8053);
nor U9640 (N_9640,N_8093,N_7838);
nor U9641 (N_9641,N_8426,N_8654);
nand U9642 (N_9642,N_8166,N_8895);
or U9643 (N_9643,N_8305,N_8450);
nand U9644 (N_9644,N_8807,N_8690);
and U9645 (N_9645,N_8363,N_7803);
or U9646 (N_9646,N_8439,N_8069);
nor U9647 (N_9647,N_8825,N_8966);
or U9648 (N_9648,N_7837,N_8777);
nand U9649 (N_9649,N_8064,N_8658);
xor U9650 (N_9650,N_8049,N_7766);
and U9651 (N_9651,N_8751,N_8323);
nand U9652 (N_9652,N_8960,N_8424);
and U9653 (N_9653,N_7652,N_7857);
or U9654 (N_9654,N_7931,N_8746);
and U9655 (N_9655,N_7655,N_7569);
nand U9656 (N_9656,N_7504,N_8071);
or U9657 (N_9657,N_8528,N_8002);
or U9658 (N_9658,N_8076,N_7761);
or U9659 (N_9659,N_8249,N_7694);
and U9660 (N_9660,N_7850,N_8822);
xnor U9661 (N_9661,N_8964,N_8913);
and U9662 (N_9662,N_8322,N_7787);
and U9663 (N_9663,N_8451,N_8122);
or U9664 (N_9664,N_7528,N_8364);
nand U9665 (N_9665,N_8496,N_7736);
nand U9666 (N_9666,N_8655,N_8244);
or U9667 (N_9667,N_8061,N_8214);
or U9668 (N_9668,N_8459,N_7553);
nand U9669 (N_9669,N_7534,N_8716);
nor U9670 (N_9670,N_7927,N_8785);
nor U9671 (N_9671,N_8382,N_8567);
or U9672 (N_9672,N_8350,N_7674);
nor U9673 (N_9673,N_7786,N_7913);
and U9674 (N_9674,N_8910,N_7792);
xor U9675 (N_9675,N_7616,N_7851);
and U9676 (N_9676,N_8100,N_8842);
or U9677 (N_9677,N_7986,N_8791);
and U9678 (N_9678,N_8515,N_8368);
and U9679 (N_9679,N_7814,N_8095);
and U9680 (N_9680,N_7754,N_8699);
nand U9681 (N_9681,N_7656,N_8216);
nor U9682 (N_9682,N_7889,N_8861);
nand U9683 (N_9683,N_8372,N_8905);
or U9684 (N_9684,N_8443,N_8637);
xor U9685 (N_9685,N_8313,N_8205);
nor U9686 (N_9686,N_7845,N_7878);
and U9687 (N_9687,N_8873,N_8281);
and U9688 (N_9688,N_7711,N_8660);
or U9689 (N_9689,N_7640,N_7909);
and U9690 (N_9690,N_8280,N_8441);
xnor U9691 (N_9691,N_8024,N_7815);
nor U9692 (N_9692,N_8546,N_8190);
nand U9693 (N_9693,N_8569,N_8086);
or U9694 (N_9694,N_8366,N_8134);
nor U9695 (N_9695,N_7893,N_7636);
or U9696 (N_9696,N_8209,N_8605);
nor U9697 (N_9697,N_8726,N_7599);
or U9698 (N_9698,N_7682,N_7758);
nand U9699 (N_9699,N_8036,N_7548);
or U9700 (N_9700,N_7572,N_8596);
nor U9701 (N_9701,N_8711,N_8490);
nor U9702 (N_9702,N_7613,N_8990);
nor U9703 (N_9703,N_7818,N_8994);
xnor U9704 (N_9704,N_8940,N_8876);
or U9705 (N_9705,N_8248,N_7685);
or U9706 (N_9706,N_8506,N_7560);
and U9707 (N_9707,N_7788,N_8534);
or U9708 (N_9708,N_8272,N_7629);
and U9709 (N_9709,N_8285,N_7923);
xnor U9710 (N_9710,N_8242,N_7628);
or U9711 (N_9711,N_7876,N_8029);
nand U9712 (N_9712,N_7707,N_8559);
and U9713 (N_9713,N_7578,N_7926);
and U9714 (N_9714,N_8452,N_8601);
or U9715 (N_9715,N_8934,N_8089);
and U9716 (N_9716,N_8806,N_8557);
xor U9717 (N_9717,N_8396,N_8718);
and U9718 (N_9718,N_8497,N_7811);
xnor U9719 (N_9719,N_7696,N_7520);
or U9720 (N_9720,N_7552,N_8367);
or U9721 (N_9721,N_7806,N_8499);
nor U9722 (N_9722,N_7901,N_7524);
xnor U9723 (N_9723,N_8252,N_8707);
or U9724 (N_9724,N_7861,N_7951);
or U9725 (N_9725,N_8290,N_7890);
nand U9726 (N_9726,N_7701,N_8782);
and U9727 (N_9727,N_7519,N_8951);
nand U9728 (N_9728,N_8075,N_8263);
xor U9729 (N_9729,N_8820,N_7824);
and U9730 (N_9730,N_8620,N_8154);
nand U9731 (N_9731,N_8161,N_8009);
or U9732 (N_9732,N_7794,N_8993);
and U9733 (N_9733,N_8955,N_8632);
nand U9734 (N_9734,N_7759,N_8804);
xnor U9735 (N_9735,N_8240,N_8700);
nor U9736 (N_9736,N_8678,N_8889);
nand U9737 (N_9737,N_8321,N_8812);
nand U9738 (N_9738,N_7666,N_7503);
or U9739 (N_9739,N_7648,N_8505);
nor U9740 (N_9740,N_8783,N_7990);
nand U9741 (N_9741,N_8197,N_8803);
xnor U9742 (N_9742,N_8344,N_7962);
nand U9743 (N_9743,N_8292,N_8294);
or U9744 (N_9744,N_8937,N_7604);
nor U9745 (N_9745,N_7731,N_8192);
nor U9746 (N_9746,N_8801,N_8665);
nand U9747 (N_9747,N_7839,N_8068);
nor U9748 (N_9748,N_7860,N_8066);
nand U9749 (N_9749,N_8416,N_7610);
nor U9750 (N_9750,N_7656,N_8236);
nor U9751 (N_9751,N_7736,N_7709);
or U9752 (N_9752,N_7775,N_8487);
and U9753 (N_9753,N_8560,N_8948);
or U9754 (N_9754,N_8314,N_7958);
nand U9755 (N_9755,N_8153,N_7793);
or U9756 (N_9756,N_7515,N_7629);
and U9757 (N_9757,N_8551,N_7811);
nand U9758 (N_9758,N_8788,N_8348);
or U9759 (N_9759,N_8184,N_7912);
nand U9760 (N_9760,N_8551,N_8384);
xor U9761 (N_9761,N_8896,N_7833);
and U9762 (N_9762,N_8016,N_8994);
or U9763 (N_9763,N_7770,N_8862);
nand U9764 (N_9764,N_7906,N_7803);
xor U9765 (N_9765,N_8671,N_8380);
nand U9766 (N_9766,N_8372,N_7959);
nand U9767 (N_9767,N_7548,N_8214);
and U9768 (N_9768,N_7921,N_8760);
and U9769 (N_9769,N_7584,N_7738);
and U9770 (N_9770,N_8295,N_8225);
nand U9771 (N_9771,N_8472,N_8283);
xnor U9772 (N_9772,N_7945,N_8958);
nor U9773 (N_9773,N_7912,N_8332);
and U9774 (N_9774,N_8902,N_8176);
nand U9775 (N_9775,N_8675,N_7915);
nor U9776 (N_9776,N_8895,N_8505);
or U9777 (N_9777,N_8620,N_8915);
nor U9778 (N_9778,N_8936,N_7770);
and U9779 (N_9779,N_8840,N_8666);
nand U9780 (N_9780,N_8720,N_8633);
xnor U9781 (N_9781,N_7554,N_7951);
nand U9782 (N_9782,N_8416,N_8775);
and U9783 (N_9783,N_7840,N_8539);
and U9784 (N_9784,N_7578,N_7657);
and U9785 (N_9785,N_8395,N_8389);
nand U9786 (N_9786,N_8564,N_7567);
nor U9787 (N_9787,N_8489,N_8555);
or U9788 (N_9788,N_8178,N_8763);
nand U9789 (N_9789,N_8247,N_8376);
nor U9790 (N_9790,N_8470,N_7762);
xnor U9791 (N_9791,N_7664,N_8956);
nor U9792 (N_9792,N_8838,N_7927);
nor U9793 (N_9793,N_8911,N_8853);
and U9794 (N_9794,N_8739,N_7994);
or U9795 (N_9795,N_7670,N_8446);
xor U9796 (N_9796,N_8185,N_8860);
nand U9797 (N_9797,N_8439,N_8358);
nor U9798 (N_9798,N_8860,N_7981);
nor U9799 (N_9799,N_8704,N_7626);
and U9800 (N_9800,N_8875,N_8009);
or U9801 (N_9801,N_7704,N_8668);
or U9802 (N_9802,N_8667,N_7790);
nand U9803 (N_9803,N_7637,N_8109);
nand U9804 (N_9804,N_8870,N_8678);
or U9805 (N_9805,N_7872,N_8675);
nand U9806 (N_9806,N_8575,N_8636);
nor U9807 (N_9807,N_8449,N_8913);
and U9808 (N_9808,N_8878,N_8086);
nor U9809 (N_9809,N_8196,N_7993);
and U9810 (N_9810,N_8259,N_8961);
and U9811 (N_9811,N_8026,N_8555);
and U9812 (N_9812,N_7771,N_7878);
and U9813 (N_9813,N_8805,N_7676);
xor U9814 (N_9814,N_8335,N_8607);
or U9815 (N_9815,N_8924,N_8205);
or U9816 (N_9816,N_8900,N_7632);
or U9817 (N_9817,N_7769,N_8476);
and U9818 (N_9818,N_7777,N_7764);
and U9819 (N_9819,N_7883,N_8721);
xnor U9820 (N_9820,N_8091,N_8661);
nand U9821 (N_9821,N_8860,N_8350);
or U9822 (N_9822,N_7721,N_8827);
or U9823 (N_9823,N_7788,N_8346);
nor U9824 (N_9824,N_8809,N_8283);
nand U9825 (N_9825,N_8421,N_7958);
and U9826 (N_9826,N_8159,N_8496);
and U9827 (N_9827,N_8137,N_8952);
xnor U9828 (N_9828,N_7796,N_8479);
nor U9829 (N_9829,N_8651,N_8539);
nor U9830 (N_9830,N_8824,N_7540);
nand U9831 (N_9831,N_8122,N_8130);
or U9832 (N_9832,N_8343,N_8243);
nor U9833 (N_9833,N_8710,N_8875);
or U9834 (N_9834,N_8890,N_8989);
nor U9835 (N_9835,N_8979,N_7966);
nor U9836 (N_9836,N_8009,N_8137);
and U9837 (N_9837,N_8184,N_8663);
nand U9838 (N_9838,N_7835,N_7549);
and U9839 (N_9839,N_8122,N_8941);
nor U9840 (N_9840,N_7641,N_8132);
or U9841 (N_9841,N_8007,N_7874);
xor U9842 (N_9842,N_8957,N_8647);
nor U9843 (N_9843,N_8850,N_7737);
nor U9844 (N_9844,N_8828,N_8541);
xnor U9845 (N_9845,N_7501,N_7557);
and U9846 (N_9846,N_7934,N_8734);
nor U9847 (N_9847,N_8592,N_8551);
nand U9848 (N_9848,N_7567,N_8512);
nand U9849 (N_9849,N_8138,N_7641);
and U9850 (N_9850,N_7773,N_7717);
nand U9851 (N_9851,N_7935,N_8877);
xnor U9852 (N_9852,N_8533,N_8078);
nand U9853 (N_9853,N_8958,N_8156);
and U9854 (N_9854,N_8446,N_7569);
and U9855 (N_9855,N_7512,N_7911);
nand U9856 (N_9856,N_8731,N_7565);
nand U9857 (N_9857,N_8468,N_8249);
nor U9858 (N_9858,N_8416,N_7738);
xor U9859 (N_9859,N_7745,N_7698);
or U9860 (N_9860,N_7753,N_7592);
and U9861 (N_9861,N_8658,N_8641);
nand U9862 (N_9862,N_8373,N_8259);
or U9863 (N_9863,N_8966,N_7748);
nand U9864 (N_9864,N_8758,N_8628);
nor U9865 (N_9865,N_7711,N_7934);
and U9866 (N_9866,N_8843,N_8438);
nand U9867 (N_9867,N_8429,N_8484);
or U9868 (N_9868,N_8420,N_8253);
nor U9869 (N_9869,N_7678,N_7654);
nand U9870 (N_9870,N_8095,N_8497);
or U9871 (N_9871,N_7673,N_8135);
xnor U9872 (N_9872,N_8428,N_8526);
nand U9873 (N_9873,N_8049,N_8350);
xor U9874 (N_9874,N_8076,N_8862);
nand U9875 (N_9875,N_8041,N_8414);
or U9876 (N_9876,N_7529,N_7929);
or U9877 (N_9877,N_8816,N_8247);
nor U9878 (N_9878,N_8312,N_8580);
nand U9879 (N_9879,N_8158,N_8557);
nor U9880 (N_9880,N_8367,N_8154);
nor U9881 (N_9881,N_8458,N_8726);
nor U9882 (N_9882,N_7705,N_8985);
nor U9883 (N_9883,N_8541,N_7939);
or U9884 (N_9884,N_8859,N_8446);
nor U9885 (N_9885,N_8282,N_7829);
and U9886 (N_9886,N_7606,N_8624);
or U9887 (N_9887,N_8012,N_7547);
nand U9888 (N_9888,N_8321,N_8515);
and U9889 (N_9889,N_7768,N_8186);
nand U9890 (N_9890,N_7899,N_8054);
and U9891 (N_9891,N_7606,N_8650);
nor U9892 (N_9892,N_8053,N_8485);
nand U9893 (N_9893,N_7612,N_8998);
or U9894 (N_9894,N_8714,N_8264);
nor U9895 (N_9895,N_7638,N_7604);
or U9896 (N_9896,N_8653,N_7742);
or U9897 (N_9897,N_8989,N_8038);
nor U9898 (N_9898,N_8099,N_7892);
nand U9899 (N_9899,N_8266,N_8267);
nand U9900 (N_9900,N_7878,N_8963);
nand U9901 (N_9901,N_8736,N_7568);
nor U9902 (N_9902,N_7841,N_7608);
nand U9903 (N_9903,N_8735,N_8218);
nor U9904 (N_9904,N_7754,N_8925);
and U9905 (N_9905,N_7773,N_7952);
nor U9906 (N_9906,N_8848,N_8407);
or U9907 (N_9907,N_8774,N_8465);
xnor U9908 (N_9908,N_7666,N_8484);
nand U9909 (N_9909,N_8757,N_8257);
nand U9910 (N_9910,N_8857,N_7770);
or U9911 (N_9911,N_7720,N_8257);
nand U9912 (N_9912,N_8384,N_8602);
nor U9913 (N_9913,N_8592,N_8429);
nor U9914 (N_9914,N_7802,N_8149);
nand U9915 (N_9915,N_8996,N_7569);
xor U9916 (N_9916,N_7597,N_8455);
and U9917 (N_9917,N_7941,N_7617);
xnor U9918 (N_9918,N_7989,N_8871);
nor U9919 (N_9919,N_8255,N_8725);
or U9920 (N_9920,N_7959,N_7984);
nand U9921 (N_9921,N_7725,N_8644);
or U9922 (N_9922,N_7864,N_7721);
nor U9923 (N_9923,N_8647,N_8864);
and U9924 (N_9924,N_8557,N_8481);
or U9925 (N_9925,N_8251,N_8492);
or U9926 (N_9926,N_8380,N_8490);
and U9927 (N_9927,N_8652,N_7901);
xnor U9928 (N_9928,N_8891,N_8763);
xor U9929 (N_9929,N_7646,N_8758);
nor U9930 (N_9930,N_7977,N_8357);
xnor U9931 (N_9931,N_8090,N_8597);
nor U9932 (N_9932,N_8380,N_8208);
nor U9933 (N_9933,N_8938,N_8196);
xnor U9934 (N_9934,N_8522,N_8911);
and U9935 (N_9935,N_7587,N_8713);
and U9936 (N_9936,N_8378,N_7891);
nor U9937 (N_9937,N_7961,N_8532);
nor U9938 (N_9938,N_7501,N_8279);
nand U9939 (N_9939,N_8010,N_8208);
and U9940 (N_9940,N_8656,N_8865);
or U9941 (N_9941,N_7616,N_7768);
nor U9942 (N_9942,N_8942,N_7633);
nand U9943 (N_9943,N_8266,N_8086);
or U9944 (N_9944,N_8021,N_7979);
nand U9945 (N_9945,N_8652,N_8876);
nor U9946 (N_9946,N_8229,N_8817);
and U9947 (N_9947,N_8890,N_8778);
nand U9948 (N_9948,N_7734,N_7878);
nor U9949 (N_9949,N_8923,N_8327);
and U9950 (N_9950,N_8301,N_8476);
nor U9951 (N_9951,N_8324,N_7796);
and U9952 (N_9952,N_8379,N_7797);
nor U9953 (N_9953,N_7875,N_8668);
nand U9954 (N_9954,N_7534,N_8639);
nand U9955 (N_9955,N_8786,N_7523);
and U9956 (N_9956,N_7604,N_8517);
xor U9957 (N_9957,N_7771,N_8612);
nand U9958 (N_9958,N_8861,N_8489);
nand U9959 (N_9959,N_8704,N_7627);
nor U9960 (N_9960,N_8071,N_7555);
and U9961 (N_9961,N_7833,N_8475);
and U9962 (N_9962,N_8430,N_8569);
nand U9963 (N_9963,N_8293,N_8102);
nor U9964 (N_9964,N_7613,N_8164);
nand U9965 (N_9965,N_8753,N_8455);
xnor U9966 (N_9966,N_8284,N_8016);
and U9967 (N_9967,N_8351,N_7722);
nand U9968 (N_9968,N_8872,N_8115);
nor U9969 (N_9969,N_8943,N_7654);
or U9970 (N_9970,N_8149,N_8174);
nand U9971 (N_9971,N_7587,N_8556);
xor U9972 (N_9972,N_8813,N_7675);
or U9973 (N_9973,N_8206,N_8826);
nand U9974 (N_9974,N_8127,N_8752);
nand U9975 (N_9975,N_7681,N_8844);
xor U9976 (N_9976,N_7868,N_7949);
xnor U9977 (N_9977,N_7828,N_7713);
nand U9978 (N_9978,N_8376,N_7590);
nor U9979 (N_9979,N_8408,N_8489);
nor U9980 (N_9980,N_7687,N_8947);
nor U9981 (N_9981,N_8434,N_8031);
nand U9982 (N_9982,N_8239,N_8605);
and U9983 (N_9983,N_8978,N_8552);
xnor U9984 (N_9984,N_7912,N_7941);
or U9985 (N_9985,N_8914,N_7500);
or U9986 (N_9986,N_7504,N_7681);
nor U9987 (N_9987,N_7941,N_7656);
or U9988 (N_9988,N_7846,N_8370);
and U9989 (N_9989,N_7855,N_8880);
nand U9990 (N_9990,N_8240,N_8968);
and U9991 (N_9991,N_7844,N_8958);
xor U9992 (N_9992,N_8645,N_8572);
and U9993 (N_9993,N_8617,N_8951);
or U9994 (N_9994,N_8135,N_8186);
nand U9995 (N_9995,N_8636,N_8405);
and U9996 (N_9996,N_8653,N_7824);
and U9997 (N_9997,N_8245,N_8824);
xnor U9998 (N_9998,N_7857,N_8783);
nor U9999 (N_9999,N_7636,N_7683);
and U10000 (N_10000,N_8623,N_7528);
or U10001 (N_10001,N_7527,N_8386);
nor U10002 (N_10002,N_7775,N_8852);
nand U10003 (N_10003,N_8798,N_8633);
xnor U10004 (N_10004,N_7673,N_7720);
nor U10005 (N_10005,N_7765,N_8421);
and U10006 (N_10006,N_7508,N_8405);
nand U10007 (N_10007,N_7750,N_8943);
and U10008 (N_10008,N_8810,N_8611);
nand U10009 (N_10009,N_8592,N_7514);
nand U10010 (N_10010,N_7586,N_8873);
nand U10011 (N_10011,N_8735,N_8499);
or U10012 (N_10012,N_8736,N_7539);
and U10013 (N_10013,N_7948,N_8432);
and U10014 (N_10014,N_8495,N_8110);
or U10015 (N_10015,N_8553,N_8663);
nand U10016 (N_10016,N_8868,N_8122);
nand U10017 (N_10017,N_7584,N_8708);
or U10018 (N_10018,N_8461,N_7681);
and U10019 (N_10019,N_8916,N_8788);
and U10020 (N_10020,N_8175,N_7703);
xor U10021 (N_10021,N_8697,N_8147);
or U10022 (N_10022,N_8464,N_7797);
or U10023 (N_10023,N_8259,N_8731);
and U10024 (N_10024,N_8164,N_8876);
nor U10025 (N_10025,N_8557,N_7776);
and U10026 (N_10026,N_7891,N_8176);
or U10027 (N_10027,N_8272,N_7735);
and U10028 (N_10028,N_8686,N_8750);
nand U10029 (N_10029,N_8136,N_7926);
nand U10030 (N_10030,N_7638,N_8779);
nor U10031 (N_10031,N_7684,N_7845);
and U10032 (N_10032,N_8501,N_8576);
nand U10033 (N_10033,N_8197,N_8104);
nor U10034 (N_10034,N_7902,N_7695);
nor U10035 (N_10035,N_8572,N_8712);
or U10036 (N_10036,N_7877,N_8867);
nor U10037 (N_10037,N_7615,N_8400);
nand U10038 (N_10038,N_7617,N_8460);
xor U10039 (N_10039,N_8983,N_8830);
or U10040 (N_10040,N_8291,N_8884);
nand U10041 (N_10041,N_7933,N_8914);
nor U10042 (N_10042,N_8543,N_8805);
and U10043 (N_10043,N_8511,N_7769);
nand U10044 (N_10044,N_7725,N_8899);
nand U10045 (N_10045,N_7881,N_8313);
or U10046 (N_10046,N_7773,N_7970);
and U10047 (N_10047,N_8401,N_7844);
xor U10048 (N_10048,N_7576,N_8247);
nand U10049 (N_10049,N_7924,N_8907);
and U10050 (N_10050,N_7590,N_7869);
nand U10051 (N_10051,N_8753,N_8298);
and U10052 (N_10052,N_8049,N_7892);
or U10053 (N_10053,N_8661,N_8330);
and U10054 (N_10054,N_7907,N_8262);
or U10055 (N_10055,N_7900,N_8364);
nand U10056 (N_10056,N_7995,N_8555);
and U10057 (N_10057,N_7785,N_8901);
nor U10058 (N_10058,N_7885,N_7698);
and U10059 (N_10059,N_8140,N_7957);
nor U10060 (N_10060,N_8177,N_8356);
nor U10061 (N_10061,N_8352,N_8016);
nand U10062 (N_10062,N_7748,N_8529);
xnor U10063 (N_10063,N_7710,N_7766);
nor U10064 (N_10064,N_8697,N_7869);
and U10065 (N_10065,N_8327,N_7733);
and U10066 (N_10066,N_7784,N_8030);
and U10067 (N_10067,N_8304,N_8368);
nor U10068 (N_10068,N_8517,N_8515);
nand U10069 (N_10069,N_8864,N_8602);
or U10070 (N_10070,N_7974,N_8266);
xnor U10071 (N_10071,N_8359,N_8021);
or U10072 (N_10072,N_7969,N_8955);
xor U10073 (N_10073,N_7841,N_7620);
nor U10074 (N_10074,N_8828,N_8704);
xor U10075 (N_10075,N_8015,N_7853);
or U10076 (N_10076,N_8743,N_8860);
nor U10077 (N_10077,N_7558,N_8839);
or U10078 (N_10078,N_8753,N_8113);
nor U10079 (N_10079,N_7842,N_8480);
nand U10080 (N_10080,N_8416,N_7970);
or U10081 (N_10081,N_8675,N_7860);
nand U10082 (N_10082,N_8211,N_7767);
xnor U10083 (N_10083,N_8228,N_7928);
nor U10084 (N_10084,N_7998,N_7658);
nand U10085 (N_10085,N_8435,N_8140);
and U10086 (N_10086,N_8293,N_8516);
nand U10087 (N_10087,N_7552,N_7673);
nor U10088 (N_10088,N_8434,N_8754);
xnor U10089 (N_10089,N_8628,N_8424);
and U10090 (N_10090,N_8013,N_8638);
nor U10091 (N_10091,N_8463,N_8362);
nand U10092 (N_10092,N_8754,N_7817);
and U10093 (N_10093,N_7599,N_7677);
or U10094 (N_10094,N_8429,N_7763);
or U10095 (N_10095,N_8750,N_8708);
and U10096 (N_10096,N_7919,N_7937);
nor U10097 (N_10097,N_8411,N_8658);
and U10098 (N_10098,N_8063,N_8135);
or U10099 (N_10099,N_7567,N_8118);
xor U10100 (N_10100,N_8959,N_7822);
xor U10101 (N_10101,N_7933,N_8063);
nor U10102 (N_10102,N_8988,N_7607);
and U10103 (N_10103,N_8382,N_8312);
nor U10104 (N_10104,N_8910,N_8452);
or U10105 (N_10105,N_8841,N_7643);
or U10106 (N_10106,N_8089,N_8766);
and U10107 (N_10107,N_8135,N_8852);
nand U10108 (N_10108,N_8866,N_8242);
and U10109 (N_10109,N_8786,N_8412);
xor U10110 (N_10110,N_8269,N_7586);
nor U10111 (N_10111,N_8544,N_8394);
xor U10112 (N_10112,N_8010,N_8184);
and U10113 (N_10113,N_7605,N_8406);
xnor U10114 (N_10114,N_7635,N_8506);
nor U10115 (N_10115,N_8939,N_8695);
and U10116 (N_10116,N_8282,N_7733);
or U10117 (N_10117,N_8905,N_8898);
xnor U10118 (N_10118,N_8993,N_8610);
and U10119 (N_10119,N_8302,N_8767);
or U10120 (N_10120,N_7804,N_7637);
or U10121 (N_10121,N_8857,N_8326);
xnor U10122 (N_10122,N_8437,N_7771);
or U10123 (N_10123,N_8562,N_8998);
nand U10124 (N_10124,N_8695,N_8891);
or U10125 (N_10125,N_8542,N_8913);
or U10126 (N_10126,N_7683,N_8391);
and U10127 (N_10127,N_8340,N_7604);
or U10128 (N_10128,N_8527,N_8371);
and U10129 (N_10129,N_7941,N_8322);
or U10130 (N_10130,N_7680,N_8351);
or U10131 (N_10131,N_8680,N_7584);
and U10132 (N_10132,N_8779,N_7902);
nor U10133 (N_10133,N_8887,N_7677);
and U10134 (N_10134,N_7857,N_8152);
nor U10135 (N_10135,N_8073,N_8730);
or U10136 (N_10136,N_7802,N_7552);
xnor U10137 (N_10137,N_8029,N_7713);
xnor U10138 (N_10138,N_8833,N_8890);
and U10139 (N_10139,N_8299,N_7665);
or U10140 (N_10140,N_7991,N_8604);
or U10141 (N_10141,N_8629,N_8466);
and U10142 (N_10142,N_8709,N_8220);
and U10143 (N_10143,N_8000,N_8430);
nand U10144 (N_10144,N_8351,N_7652);
xnor U10145 (N_10145,N_8685,N_8585);
nor U10146 (N_10146,N_8385,N_7640);
or U10147 (N_10147,N_8795,N_7944);
nand U10148 (N_10148,N_8654,N_8558);
nand U10149 (N_10149,N_8362,N_8922);
nand U10150 (N_10150,N_8536,N_7692);
nand U10151 (N_10151,N_8171,N_7750);
or U10152 (N_10152,N_8887,N_8893);
nand U10153 (N_10153,N_8693,N_8282);
nand U10154 (N_10154,N_8988,N_8302);
xor U10155 (N_10155,N_8192,N_8270);
xor U10156 (N_10156,N_7548,N_7514);
nor U10157 (N_10157,N_8707,N_7993);
xor U10158 (N_10158,N_8160,N_8660);
nand U10159 (N_10159,N_8108,N_7924);
and U10160 (N_10160,N_7567,N_7950);
nor U10161 (N_10161,N_8217,N_7780);
or U10162 (N_10162,N_7963,N_8097);
nand U10163 (N_10163,N_8757,N_7639);
nand U10164 (N_10164,N_7569,N_7547);
nand U10165 (N_10165,N_7584,N_8087);
and U10166 (N_10166,N_8591,N_8834);
or U10167 (N_10167,N_7961,N_8675);
nand U10168 (N_10168,N_8291,N_8091);
or U10169 (N_10169,N_7716,N_7817);
nor U10170 (N_10170,N_8210,N_8537);
nand U10171 (N_10171,N_8970,N_8702);
and U10172 (N_10172,N_8341,N_8268);
nand U10173 (N_10173,N_7894,N_8096);
or U10174 (N_10174,N_8263,N_8480);
nand U10175 (N_10175,N_7999,N_8173);
and U10176 (N_10176,N_8728,N_7804);
or U10177 (N_10177,N_8824,N_8468);
or U10178 (N_10178,N_8761,N_8473);
xnor U10179 (N_10179,N_8702,N_7860);
xor U10180 (N_10180,N_8164,N_7838);
nand U10181 (N_10181,N_7918,N_7692);
or U10182 (N_10182,N_8138,N_7514);
xnor U10183 (N_10183,N_8955,N_8535);
xnor U10184 (N_10184,N_8037,N_8076);
nor U10185 (N_10185,N_7733,N_8858);
nand U10186 (N_10186,N_8326,N_8517);
and U10187 (N_10187,N_8184,N_8314);
or U10188 (N_10188,N_8661,N_8902);
or U10189 (N_10189,N_7741,N_8700);
or U10190 (N_10190,N_8517,N_8363);
and U10191 (N_10191,N_8370,N_8881);
nand U10192 (N_10192,N_8350,N_8035);
nor U10193 (N_10193,N_8808,N_8212);
or U10194 (N_10194,N_8476,N_7969);
and U10195 (N_10195,N_8975,N_7586);
and U10196 (N_10196,N_8723,N_7543);
or U10197 (N_10197,N_8441,N_8763);
or U10198 (N_10198,N_8988,N_8469);
or U10199 (N_10199,N_8167,N_7745);
and U10200 (N_10200,N_7788,N_8960);
and U10201 (N_10201,N_7931,N_7803);
and U10202 (N_10202,N_8435,N_7847);
or U10203 (N_10203,N_7746,N_8060);
and U10204 (N_10204,N_8109,N_7937);
and U10205 (N_10205,N_7893,N_8854);
and U10206 (N_10206,N_8833,N_8700);
nor U10207 (N_10207,N_8985,N_8404);
nor U10208 (N_10208,N_7749,N_8690);
nand U10209 (N_10209,N_7659,N_7861);
and U10210 (N_10210,N_8129,N_7628);
and U10211 (N_10211,N_8624,N_8117);
and U10212 (N_10212,N_8746,N_8684);
and U10213 (N_10213,N_8779,N_8439);
or U10214 (N_10214,N_8010,N_7561);
nand U10215 (N_10215,N_7768,N_7512);
xnor U10216 (N_10216,N_8089,N_8442);
nor U10217 (N_10217,N_8366,N_8075);
xnor U10218 (N_10218,N_7993,N_7630);
nor U10219 (N_10219,N_7755,N_8446);
nand U10220 (N_10220,N_7876,N_8995);
xnor U10221 (N_10221,N_8174,N_8934);
and U10222 (N_10222,N_7789,N_7766);
or U10223 (N_10223,N_7950,N_7746);
nand U10224 (N_10224,N_8380,N_8475);
or U10225 (N_10225,N_7808,N_7987);
or U10226 (N_10226,N_7885,N_7650);
nand U10227 (N_10227,N_8993,N_8128);
and U10228 (N_10228,N_8039,N_8227);
nand U10229 (N_10229,N_8843,N_8817);
nand U10230 (N_10230,N_8673,N_7640);
xnor U10231 (N_10231,N_8537,N_7725);
xor U10232 (N_10232,N_7569,N_7887);
nand U10233 (N_10233,N_7972,N_8274);
nor U10234 (N_10234,N_7517,N_8239);
nand U10235 (N_10235,N_7655,N_8281);
and U10236 (N_10236,N_8138,N_8930);
nor U10237 (N_10237,N_7743,N_7806);
or U10238 (N_10238,N_8116,N_7549);
or U10239 (N_10239,N_8467,N_8134);
nand U10240 (N_10240,N_7997,N_8619);
nand U10241 (N_10241,N_8388,N_7720);
or U10242 (N_10242,N_8923,N_8974);
xnor U10243 (N_10243,N_7534,N_8979);
nand U10244 (N_10244,N_8744,N_8748);
or U10245 (N_10245,N_8953,N_8323);
and U10246 (N_10246,N_8210,N_8772);
and U10247 (N_10247,N_8047,N_7563);
nand U10248 (N_10248,N_8716,N_8374);
nand U10249 (N_10249,N_8518,N_7632);
nor U10250 (N_10250,N_8247,N_8756);
and U10251 (N_10251,N_7638,N_7689);
and U10252 (N_10252,N_8500,N_8872);
and U10253 (N_10253,N_8460,N_8592);
and U10254 (N_10254,N_8147,N_7870);
xnor U10255 (N_10255,N_8747,N_8729);
xor U10256 (N_10256,N_8401,N_8704);
nor U10257 (N_10257,N_7709,N_8989);
nand U10258 (N_10258,N_7883,N_8802);
xor U10259 (N_10259,N_8678,N_8796);
and U10260 (N_10260,N_7606,N_8472);
nor U10261 (N_10261,N_8037,N_8649);
and U10262 (N_10262,N_8583,N_8298);
or U10263 (N_10263,N_8927,N_7822);
and U10264 (N_10264,N_8868,N_7685);
and U10265 (N_10265,N_8142,N_8046);
xnor U10266 (N_10266,N_8565,N_8860);
or U10267 (N_10267,N_8798,N_8461);
or U10268 (N_10268,N_8785,N_8879);
and U10269 (N_10269,N_8552,N_8777);
nor U10270 (N_10270,N_8017,N_8289);
or U10271 (N_10271,N_8513,N_8125);
nor U10272 (N_10272,N_8816,N_8932);
or U10273 (N_10273,N_7845,N_8332);
and U10274 (N_10274,N_8305,N_7784);
nor U10275 (N_10275,N_8704,N_8224);
nand U10276 (N_10276,N_8962,N_8541);
nor U10277 (N_10277,N_7992,N_8790);
and U10278 (N_10278,N_8750,N_8773);
nor U10279 (N_10279,N_8511,N_8847);
nand U10280 (N_10280,N_8843,N_7854);
or U10281 (N_10281,N_8092,N_8285);
or U10282 (N_10282,N_7718,N_8379);
nand U10283 (N_10283,N_8505,N_8452);
xor U10284 (N_10284,N_7882,N_7658);
and U10285 (N_10285,N_8559,N_7665);
nor U10286 (N_10286,N_8901,N_7598);
and U10287 (N_10287,N_7605,N_8535);
nand U10288 (N_10288,N_8631,N_7542);
or U10289 (N_10289,N_8046,N_8578);
nand U10290 (N_10290,N_7517,N_8997);
nor U10291 (N_10291,N_7665,N_7849);
nand U10292 (N_10292,N_8951,N_7734);
or U10293 (N_10293,N_7685,N_8009);
nand U10294 (N_10294,N_8616,N_7650);
nand U10295 (N_10295,N_7552,N_7583);
and U10296 (N_10296,N_8715,N_8706);
nor U10297 (N_10297,N_8441,N_8210);
and U10298 (N_10298,N_7744,N_7584);
xnor U10299 (N_10299,N_8908,N_7688);
nor U10300 (N_10300,N_8785,N_8145);
and U10301 (N_10301,N_8721,N_8902);
nand U10302 (N_10302,N_7691,N_7540);
xnor U10303 (N_10303,N_8989,N_8008);
nand U10304 (N_10304,N_7805,N_8566);
and U10305 (N_10305,N_8473,N_8853);
nor U10306 (N_10306,N_8841,N_7652);
nor U10307 (N_10307,N_8736,N_8753);
or U10308 (N_10308,N_7677,N_7853);
and U10309 (N_10309,N_8989,N_7617);
and U10310 (N_10310,N_8899,N_7596);
nand U10311 (N_10311,N_8449,N_8968);
nand U10312 (N_10312,N_7968,N_8161);
nor U10313 (N_10313,N_8777,N_8630);
nor U10314 (N_10314,N_8905,N_8602);
nand U10315 (N_10315,N_7697,N_7915);
or U10316 (N_10316,N_7701,N_8521);
or U10317 (N_10317,N_8078,N_7723);
or U10318 (N_10318,N_7679,N_8610);
nand U10319 (N_10319,N_8039,N_8127);
nor U10320 (N_10320,N_8561,N_8543);
nor U10321 (N_10321,N_7502,N_7550);
and U10322 (N_10322,N_7931,N_8236);
nand U10323 (N_10323,N_7840,N_8421);
nor U10324 (N_10324,N_7544,N_8711);
or U10325 (N_10325,N_8934,N_8422);
nor U10326 (N_10326,N_7990,N_8691);
nand U10327 (N_10327,N_8040,N_8025);
nor U10328 (N_10328,N_8632,N_7599);
nand U10329 (N_10329,N_8461,N_8762);
or U10330 (N_10330,N_7520,N_7512);
nand U10331 (N_10331,N_8700,N_8825);
and U10332 (N_10332,N_8761,N_7880);
nor U10333 (N_10333,N_8085,N_7739);
nand U10334 (N_10334,N_7718,N_8934);
or U10335 (N_10335,N_8657,N_8457);
nor U10336 (N_10336,N_7620,N_7680);
nor U10337 (N_10337,N_7933,N_8526);
xor U10338 (N_10338,N_8197,N_8106);
nand U10339 (N_10339,N_8284,N_8711);
nand U10340 (N_10340,N_7585,N_8581);
or U10341 (N_10341,N_7558,N_8862);
and U10342 (N_10342,N_8153,N_7654);
nand U10343 (N_10343,N_8426,N_7667);
nand U10344 (N_10344,N_8080,N_8533);
or U10345 (N_10345,N_8299,N_8308);
nand U10346 (N_10346,N_7864,N_8236);
xnor U10347 (N_10347,N_8085,N_7769);
nand U10348 (N_10348,N_8651,N_8124);
and U10349 (N_10349,N_8953,N_8801);
and U10350 (N_10350,N_8430,N_8873);
nor U10351 (N_10351,N_8827,N_8263);
nor U10352 (N_10352,N_8529,N_8202);
nor U10353 (N_10353,N_7739,N_8154);
or U10354 (N_10354,N_7696,N_7894);
and U10355 (N_10355,N_8764,N_7860);
or U10356 (N_10356,N_7756,N_7799);
or U10357 (N_10357,N_8866,N_8626);
nor U10358 (N_10358,N_8089,N_7559);
or U10359 (N_10359,N_8086,N_8591);
nor U10360 (N_10360,N_8302,N_8984);
nor U10361 (N_10361,N_8220,N_7565);
nand U10362 (N_10362,N_7734,N_7568);
nor U10363 (N_10363,N_8430,N_7594);
and U10364 (N_10364,N_8191,N_8545);
and U10365 (N_10365,N_8930,N_7961);
xnor U10366 (N_10366,N_7917,N_8373);
and U10367 (N_10367,N_8150,N_7507);
nand U10368 (N_10368,N_8204,N_8751);
xnor U10369 (N_10369,N_8980,N_8467);
nand U10370 (N_10370,N_8204,N_8589);
or U10371 (N_10371,N_8518,N_8616);
and U10372 (N_10372,N_8151,N_7877);
and U10373 (N_10373,N_8366,N_8182);
or U10374 (N_10374,N_8200,N_7851);
and U10375 (N_10375,N_8873,N_8343);
or U10376 (N_10376,N_8498,N_7868);
nor U10377 (N_10377,N_8035,N_8088);
or U10378 (N_10378,N_8848,N_7870);
nor U10379 (N_10379,N_8858,N_8316);
nor U10380 (N_10380,N_7537,N_7690);
xnor U10381 (N_10381,N_8968,N_8861);
nor U10382 (N_10382,N_8880,N_8768);
and U10383 (N_10383,N_7931,N_7659);
or U10384 (N_10384,N_8095,N_8703);
and U10385 (N_10385,N_8731,N_8206);
nand U10386 (N_10386,N_8893,N_7768);
and U10387 (N_10387,N_8338,N_8930);
xnor U10388 (N_10388,N_8771,N_8087);
nand U10389 (N_10389,N_8382,N_8807);
nand U10390 (N_10390,N_7604,N_7539);
nor U10391 (N_10391,N_8505,N_7651);
and U10392 (N_10392,N_7854,N_7659);
xor U10393 (N_10393,N_8070,N_7571);
and U10394 (N_10394,N_7557,N_8524);
xnor U10395 (N_10395,N_7724,N_7746);
and U10396 (N_10396,N_8643,N_7627);
and U10397 (N_10397,N_7760,N_7651);
or U10398 (N_10398,N_8362,N_8251);
nor U10399 (N_10399,N_8487,N_8115);
nor U10400 (N_10400,N_8274,N_7888);
xor U10401 (N_10401,N_7510,N_8812);
or U10402 (N_10402,N_8262,N_8459);
nor U10403 (N_10403,N_8208,N_7988);
xor U10404 (N_10404,N_7727,N_7759);
or U10405 (N_10405,N_7976,N_7736);
nor U10406 (N_10406,N_8660,N_8340);
and U10407 (N_10407,N_7908,N_8732);
nand U10408 (N_10408,N_7839,N_8945);
or U10409 (N_10409,N_7680,N_8562);
and U10410 (N_10410,N_7601,N_8486);
or U10411 (N_10411,N_7629,N_8032);
xnor U10412 (N_10412,N_8697,N_8878);
nand U10413 (N_10413,N_8446,N_8596);
or U10414 (N_10414,N_8606,N_8752);
nand U10415 (N_10415,N_8984,N_8877);
or U10416 (N_10416,N_8243,N_8607);
xnor U10417 (N_10417,N_8364,N_8155);
or U10418 (N_10418,N_7933,N_8310);
nand U10419 (N_10419,N_7836,N_7992);
nand U10420 (N_10420,N_8996,N_8342);
nand U10421 (N_10421,N_8640,N_8625);
or U10422 (N_10422,N_7828,N_8617);
or U10423 (N_10423,N_7683,N_7967);
nand U10424 (N_10424,N_8564,N_8254);
nor U10425 (N_10425,N_8466,N_8576);
and U10426 (N_10426,N_8676,N_7519);
xnor U10427 (N_10427,N_8802,N_8770);
xnor U10428 (N_10428,N_8186,N_8003);
nand U10429 (N_10429,N_8347,N_8339);
nand U10430 (N_10430,N_7943,N_8982);
or U10431 (N_10431,N_8179,N_8445);
and U10432 (N_10432,N_8298,N_7751);
nor U10433 (N_10433,N_8807,N_8799);
or U10434 (N_10434,N_8441,N_7669);
nand U10435 (N_10435,N_7637,N_8298);
nor U10436 (N_10436,N_8192,N_8085);
or U10437 (N_10437,N_8528,N_8893);
and U10438 (N_10438,N_8299,N_8706);
nor U10439 (N_10439,N_7931,N_8511);
nand U10440 (N_10440,N_8194,N_8849);
nand U10441 (N_10441,N_8654,N_8256);
and U10442 (N_10442,N_8919,N_7942);
nor U10443 (N_10443,N_8190,N_8246);
nor U10444 (N_10444,N_8842,N_7791);
nand U10445 (N_10445,N_8767,N_8113);
nor U10446 (N_10446,N_7814,N_8074);
or U10447 (N_10447,N_7822,N_7560);
and U10448 (N_10448,N_8075,N_8264);
nand U10449 (N_10449,N_8514,N_8494);
nand U10450 (N_10450,N_7763,N_8637);
xnor U10451 (N_10451,N_7753,N_8273);
nand U10452 (N_10452,N_8619,N_8296);
nand U10453 (N_10453,N_8018,N_8807);
nand U10454 (N_10454,N_8667,N_7574);
nor U10455 (N_10455,N_8556,N_8514);
nor U10456 (N_10456,N_8325,N_8279);
nor U10457 (N_10457,N_8659,N_8972);
nand U10458 (N_10458,N_8496,N_8977);
nand U10459 (N_10459,N_8761,N_7981);
or U10460 (N_10460,N_8266,N_8426);
and U10461 (N_10461,N_7786,N_8917);
xnor U10462 (N_10462,N_7900,N_8486);
nor U10463 (N_10463,N_8655,N_7814);
and U10464 (N_10464,N_8694,N_8426);
nand U10465 (N_10465,N_7739,N_7626);
nor U10466 (N_10466,N_7638,N_8087);
nand U10467 (N_10467,N_7635,N_8416);
xnor U10468 (N_10468,N_8642,N_8542);
nand U10469 (N_10469,N_7562,N_8238);
or U10470 (N_10470,N_8328,N_8210);
or U10471 (N_10471,N_8880,N_8956);
and U10472 (N_10472,N_8004,N_7751);
nand U10473 (N_10473,N_8590,N_7799);
nor U10474 (N_10474,N_8558,N_8589);
nand U10475 (N_10475,N_7983,N_8622);
or U10476 (N_10476,N_8506,N_8313);
or U10477 (N_10477,N_8511,N_8547);
or U10478 (N_10478,N_8878,N_8064);
or U10479 (N_10479,N_8304,N_8756);
nand U10480 (N_10480,N_7562,N_8216);
nand U10481 (N_10481,N_8778,N_7944);
xnor U10482 (N_10482,N_8605,N_8103);
xnor U10483 (N_10483,N_8770,N_8140);
or U10484 (N_10484,N_8475,N_7614);
nor U10485 (N_10485,N_8211,N_8275);
and U10486 (N_10486,N_8630,N_7666);
nand U10487 (N_10487,N_8518,N_8454);
or U10488 (N_10488,N_7871,N_8561);
nand U10489 (N_10489,N_8312,N_7830);
nand U10490 (N_10490,N_7757,N_8076);
nor U10491 (N_10491,N_7585,N_8980);
and U10492 (N_10492,N_8765,N_7858);
xnor U10493 (N_10493,N_8569,N_8642);
xnor U10494 (N_10494,N_7505,N_8876);
nand U10495 (N_10495,N_8118,N_8728);
nand U10496 (N_10496,N_8032,N_7859);
nor U10497 (N_10497,N_8682,N_7645);
xor U10498 (N_10498,N_7593,N_8063);
nor U10499 (N_10499,N_8354,N_8879);
nand U10500 (N_10500,N_10490,N_9433);
or U10501 (N_10501,N_9041,N_10450);
nor U10502 (N_10502,N_10259,N_9100);
nand U10503 (N_10503,N_9118,N_9925);
nand U10504 (N_10504,N_9023,N_10073);
nor U10505 (N_10505,N_10439,N_10030);
nor U10506 (N_10506,N_9368,N_10068);
or U10507 (N_10507,N_10369,N_10031);
or U10508 (N_10508,N_10447,N_9224);
nor U10509 (N_10509,N_9779,N_10260);
xor U10510 (N_10510,N_10434,N_9838);
nor U10511 (N_10511,N_9822,N_10164);
or U10512 (N_10512,N_9062,N_9871);
nand U10513 (N_10513,N_9374,N_9587);
xnor U10514 (N_10514,N_10291,N_9780);
nand U10515 (N_10515,N_10248,N_10322);
nor U10516 (N_10516,N_9198,N_9693);
xor U10517 (N_10517,N_10377,N_9643);
and U10518 (N_10518,N_9778,N_9622);
xor U10519 (N_10519,N_10430,N_10213);
xnor U10520 (N_10520,N_9088,N_10029);
nor U10521 (N_10521,N_10080,N_9133);
or U10522 (N_10522,N_10237,N_9534);
and U10523 (N_10523,N_9045,N_10192);
nand U10524 (N_10524,N_9136,N_9730);
and U10525 (N_10525,N_9801,N_9843);
nor U10526 (N_10526,N_10395,N_9781);
xnor U10527 (N_10527,N_10462,N_10421);
and U10528 (N_10528,N_9501,N_10306);
nand U10529 (N_10529,N_9272,N_9735);
nand U10530 (N_10530,N_10338,N_9457);
nand U10531 (N_10531,N_10140,N_9867);
and U10532 (N_10532,N_9628,N_9619);
and U10533 (N_10533,N_9896,N_9655);
or U10534 (N_10534,N_9018,N_10361);
nand U10535 (N_10535,N_9446,N_9279);
nand U10536 (N_10536,N_9346,N_9357);
nand U10537 (N_10537,N_9511,N_10319);
nor U10538 (N_10538,N_9836,N_9848);
nor U10539 (N_10539,N_9676,N_9505);
xnor U10540 (N_10540,N_9086,N_10337);
nor U10541 (N_10541,N_9303,N_9153);
nor U10542 (N_10542,N_9868,N_10046);
nor U10543 (N_10543,N_10116,N_10406);
or U10544 (N_10544,N_10044,N_10240);
nor U10545 (N_10545,N_9015,N_9466);
nor U10546 (N_10546,N_10011,N_10081);
and U10547 (N_10547,N_9448,N_9349);
or U10548 (N_10548,N_9365,N_10339);
or U10549 (N_10549,N_10124,N_9308);
nor U10550 (N_10550,N_9788,N_10346);
nand U10551 (N_10551,N_10372,N_9234);
and U10552 (N_10552,N_10344,N_9751);
xor U10553 (N_10553,N_9502,N_9179);
or U10554 (N_10554,N_10489,N_10302);
or U10555 (N_10555,N_9219,N_10463);
and U10556 (N_10556,N_9020,N_10300);
nand U10557 (N_10557,N_10008,N_10028);
or U10558 (N_10558,N_9954,N_9769);
nand U10559 (N_10559,N_9340,N_9356);
or U10560 (N_10560,N_9532,N_10095);
nor U10561 (N_10561,N_9116,N_9957);
and U10562 (N_10562,N_10254,N_9561);
and U10563 (N_10563,N_10429,N_10146);
xnor U10564 (N_10564,N_9296,N_9911);
or U10565 (N_10565,N_10403,N_9550);
xor U10566 (N_10566,N_9402,N_9996);
or U10567 (N_10567,N_10191,N_9053);
or U10568 (N_10568,N_10088,N_9207);
nor U10569 (N_10569,N_9940,N_9326);
nand U10570 (N_10570,N_10303,N_9991);
and U10571 (N_10571,N_10170,N_9266);
nand U10572 (N_10572,N_9560,N_10190);
nand U10573 (N_10573,N_10202,N_9385);
and U10574 (N_10574,N_9804,N_9396);
nor U10575 (N_10575,N_9264,N_9080);
nor U10576 (N_10576,N_9414,N_9943);
nand U10577 (N_10577,N_9454,N_9019);
and U10578 (N_10578,N_10482,N_10043);
or U10579 (N_10579,N_9339,N_9874);
xnor U10580 (N_10580,N_9003,N_9076);
nand U10581 (N_10581,N_9503,N_9802);
and U10582 (N_10582,N_10267,N_9885);
nor U10583 (N_10583,N_10304,N_9872);
nand U10584 (N_10584,N_9223,N_10492);
and U10585 (N_10585,N_9125,N_9001);
nand U10586 (N_10586,N_10065,N_10066);
nand U10587 (N_10587,N_10071,N_9586);
and U10588 (N_10588,N_9737,N_9172);
and U10589 (N_10589,N_9005,N_10126);
and U10590 (N_10590,N_10472,N_9343);
and U10591 (N_10591,N_9662,N_9312);
xor U10592 (N_10592,N_9409,N_9582);
nand U10593 (N_10593,N_10138,N_9362);
nor U10594 (N_10594,N_9825,N_10148);
nand U10595 (N_10595,N_9151,N_10469);
and U10596 (N_10596,N_10311,N_9858);
and U10597 (N_10597,N_9174,N_9170);
nand U10598 (N_10598,N_9820,N_10448);
nor U10599 (N_10599,N_9334,N_10210);
nor U10600 (N_10600,N_10105,N_10035);
and U10601 (N_10601,N_10166,N_9504);
and U10602 (N_10602,N_9932,N_9097);
nand U10603 (N_10603,N_10340,N_9766);
nand U10604 (N_10604,N_9623,N_10175);
xnor U10605 (N_10605,N_9635,N_10057);
nand U10606 (N_10606,N_10464,N_9739);
xnor U10607 (N_10607,N_10263,N_10015);
or U10608 (N_10608,N_9884,N_9301);
or U10609 (N_10609,N_9220,N_10324);
or U10610 (N_10610,N_9493,N_9875);
and U10611 (N_10611,N_9064,N_9255);
or U10612 (N_10612,N_9700,N_10039);
nor U10613 (N_10613,N_9948,N_10089);
nor U10614 (N_10614,N_9383,N_10010);
nor U10615 (N_10615,N_9541,N_9039);
nor U10616 (N_10616,N_9525,N_10180);
or U10617 (N_10617,N_10370,N_9682);
and U10618 (N_10618,N_9074,N_9661);
nor U10619 (N_10619,N_9947,N_10474);
and U10620 (N_10620,N_9554,N_9427);
nor U10621 (N_10621,N_10000,N_10273);
or U10622 (N_10622,N_9063,N_9258);
nor U10623 (N_10623,N_10204,N_10113);
nor U10624 (N_10624,N_9036,N_9920);
nand U10625 (N_10625,N_10173,N_9071);
nand U10626 (N_10626,N_9341,N_10280);
nand U10627 (N_10627,N_9621,N_9696);
nor U10628 (N_10628,N_9453,N_9973);
xnor U10629 (N_10629,N_9160,N_10085);
xor U10630 (N_10630,N_9579,N_9564);
or U10631 (N_10631,N_9854,N_9703);
nand U10632 (N_10632,N_9157,N_10145);
nand U10633 (N_10633,N_10378,N_9846);
xnor U10634 (N_10634,N_9906,N_9862);
and U10635 (N_10635,N_10309,N_9016);
nor U10636 (N_10636,N_9360,N_9028);
and U10637 (N_10637,N_10432,N_10056);
or U10638 (N_10638,N_9197,N_10392);
and U10639 (N_10639,N_9800,N_9611);
nand U10640 (N_10640,N_10215,N_9096);
nor U10641 (N_10641,N_9320,N_10161);
nand U10642 (N_10642,N_10257,N_9314);
nand U10643 (N_10643,N_10022,N_9189);
or U10644 (N_10644,N_10241,N_10147);
or U10645 (N_10645,N_10365,N_10315);
nor U10646 (N_10646,N_9990,N_10150);
nor U10647 (N_10647,N_9390,N_9165);
or U10648 (N_10648,N_9372,N_9995);
and U10649 (N_10649,N_9674,N_9119);
and U10650 (N_10650,N_10108,N_9070);
nand U10651 (N_10651,N_10208,N_10007);
nor U10652 (N_10652,N_9888,N_9715);
and U10653 (N_10653,N_9120,N_10364);
nand U10654 (N_10654,N_10314,N_9930);
and U10655 (N_10655,N_9772,N_9458);
nor U10656 (N_10656,N_10288,N_9997);
or U10657 (N_10657,N_9783,N_9926);
and U10658 (N_10658,N_9404,N_9900);
nand U10659 (N_10659,N_9608,N_10358);
nand U10660 (N_10660,N_9209,N_9759);
or U10661 (N_10661,N_10379,N_9529);
or U10662 (N_10662,N_9352,N_9006);
or U10663 (N_10663,N_10197,N_9573);
xor U10664 (N_10664,N_10373,N_10341);
nand U10665 (N_10665,N_9934,N_9842);
nor U10666 (N_10666,N_9426,N_9555);
and U10667 (N_10667,N_9306,N_10299);
nand U10668 (N_10668,N_9022,N_9317);
nor U10669 (N_10669,N_9513,N_10473);
nand U10670 (N_10670,N_9687,N_9978);
nor U10671 (N_10671,N_9413,N_10194);
and U10672 (N_10672,N_9826,N_9733);
nand U10673 (N_10673,N_9130,N_9147);
nand U10674 (N_10674,N_9060,N_10082);
or U10675 (N_10675,N_10078,N_10227);
and U10676 (N_10676,N_10075,N_9269);
nor U10677 (N_10677,N_9649,N_9091);
or U10678 (N_10678,N_9870,N_10312);
nand U10679 (N_10679,N_9175,N_10349);
nand U10680 (N_10680,N_10282,N_9112);
or U10681 (N_10681,N_9916,N_9734);
and U10682 (N_10682,N_9637,N_10343);
nor U10683 (N_10683,N_10268,N_10062);
nor U10684 (N_10684,N_9178,N_9110);
nand U10685 (N_10685,N_9650,N_9371);
and U10686 (N_10686,N_9468,N_9748);
or U10687 (N_10687,N_10021,N_9618);
nand U10688 (N_10688,N_10196,N_10048);
or U10689 (N_10689,N_9988,N_9857);
xor U10690 (N_10690,N_9976,N_9217);
nand U10691 (N_10691,N_9205,N_9845);
xnor U10692 (N_10692,N_9139,N_9704);
or U10693 (N_10693,N_9585,N_10331);
or U10694 (N_10694,N_9685,N_10053);
or U10695 (N_10695,N_10092,N_10086);
nand U10696 (N_10696,N_9447,N_9399);
and U10697 (N_10697,N_9889,N_9945);
nand U10698 (N_10698,N_10209,N_9031);
nor U10699 (N_10699,N_10396,N_9578);
nand U10700 (N_10700,N_9285,N_9672);
and U10701 (N_10701,N_10265,N_9725);
and U10702 (N_10702,N_9986,N_9809);
nor U10703 (N_10703,N_9192,N_9512);
or U10704 (N_10704,N_9380,N_9497);
xnor U10705 (N_10705,N_9606,N_9998);
nor U10706 (N_10706,N_9971,N_9850);
nand U10707 (N_10707,N_10249,N_10231);
nand U10708 (N_10708,N_10363,N_9090);
or U10709 (N_10709,N_10405,N_9210);
xor U10710 (N_10710,N_9008,N_9232);
xor U10711 (N_10711,N_10033,N_9955);
nor U10712 (N_10712,N_9571,N_10200);
nor U10713 (N_10713,N_9283,N_10497);
nand U10714 (N_10714,N_10245,N_9007);
nor U10715 (N_10715,N_9823,N_9524);
or U10716 (N_10716,N_9358,N_10366);
and U10717 (N_10717,N_9690,N_10342);
xor U10718 (N_10718,N_10367,N_10467);
nand U10719 (N_10719,N_9467,N_9882);
nor U10720 (N_10720,N_9811,N_10480);
or U10721 (N_10721,N_9345,N_9329);
nand U10722 (N_10722,N_9043,N_9040);
xor U10723 (N_10723,N_9794,N_10067);
xor U10724 (N_10724,N_9364,N_9068);
xor U10725 (N_10725,N_9065,N_10156);
nor U10726 (N_10726,N_10079,N_9231);
nor U10727 (N_10727,N_10454,N_10069);
and U10728 (N_10728,N_10328,N_9714);
and U10729 (N_10729,N_10375,N_9441);
nand U10730 (N_10730,N_9496,N_9247);
and U10731 (N_10731,N_9230,N_9167);
and U10732 (N_10732,N_10002,N_10440);
nand U10733 (N_10733,N_10335,N_9961);
xor U10734 (N_10734,N_9051,N_10123);
and U10735 (N_10735,N_10098,N_9559);
nand U10736 (N_10736,N_10054,N_9261);
and U10737 (N_10737,N_9083,N_9121);
nand U10738 (N_10738,N_10225,N_10049);
or U10739 (N_10739,N_9057,N_9200);
nor U10740 (N_10740,N_9239,N_9977);
nor U10741 (N_10741,N_10277,N_9631);
nor U10742 (N_10742,N_10136,N_9292);
xnor U10743 (N_10743,N_10368,N_9143);
and U10744 (N_10744,N_9675,N_10444);
and U10745 (N_10745,N_10040,N_10333);
nor U10746 (N_10746,N_10295,N_9324);
and U10747 (N_10747,N_10347,N_10435);
nand U10748 (N_10748,N_9092,N_10132);
and U10749 (N_10749,N_9475,N_10184);
nor U10750 (N_10750,N_9939,N_9913);
nor U10751 (N_10751,N_10470,N_9681);
or U10752 (N_10752,N_10034,N_9032);
nand U10753 (N_10753,N_9983,N_9046);
or U10754 (N_10754,N_9442,N_10386);
xor U10755 (N_10755,N_9054,N_9716);
nor U10756 (N_10756,N_9240,N_9771);
nor U10757 (N_10757,N_9227,N_9879);
or U10758 (N_10758,N_9342,N_9464);
nor U10759 (N_10759,N_9952,N_9294);
nand U10760 (N_10760,N_9514,N_9401);
and U10761 (N_10761,N_9812,N_9455);
nor U10762 (N_10762,N_9421,N_9833);
or U10763 (N_10763,N_9304,N_10313);
or U10764 (N_10764,N_9403,N_10220);
and U10765 (N_10765,N_9892,N_9411);
and U10766 (N_10766,N_9377,N_9485);
or U10767 (N_10767,N_9353,N_9979);
nor U10768 (N_10768,N_9536,N_9914);
nor U10769 (N_10769,N_10168,N_9705);
nor U10770 (N_10770,N_9894,N_9449);
and U10771 (N_10771,N_9904,N_9335);
and U10772 (N_10772,N_9658,N_9935);
nand U10773 (N_10773,N_9236,N_9840);
and U10774 (N_10774,N_9177,N_9336);
nand U10775 (N_10775,N_9969,N_9389);
nor U10776 (N_10776,N_10416,N_9545);
or U10777 (N_10777,N_10233,N_9465);
xnor U10778 (N_10778,N_10498,N_10045);
or U10779 (N_10779,N_9533,N_9395);
and U10780 (N_10780,N_9187,N_10238);
or U10781 (N_10781,N_9055,N_9479);
nand U10782 (N_10782,N_10228,N_9087);
nor U10783 (N_10783,N_9841,N_9203);
nor U10784 (N_10784,N_9262,N_10266);
nor U10785 (N_10785,N_10137,N_10388);
nand U10786 (N_10786,N_9653,N_9280);
xnor U10787 (N_10787,N_9012,N_9905);
or U10788 (N_10788,N_9756,N_9790);
nor U10789 (N_10789,N_9516,N_10475);
xor U10790 (N_10790,N_9010,N_10360);
or U10791 (N_10791,N_10001,N_9201);
or U10792 (N_10792,N_9689,N_9480);
and U10793 (N_10793,N_10422,N_10258);
or U10794 (N_10794,N_10070,N_9946);
xnor U10795 (N_10795,N_10418,N_9067);
or U10796 (N_10796,N_9056,N_9648);
or U10797 (N_10797,N_10409,N_9141);
nand U10798 (N_10798,N_9489,N_9860);
or U10799 (N_10799,N_9741,N_9123);
nor U10800 (N_10800,N_10326,N_10055);
and U10801 (N_10801,N_9697,N_9557);
xor U10802 (N_10802,N_10290,N_9819);
and U10803 (N_10803,N_9965,N_10401);
or U10804 (N_10804,N_10308,N_9162);
xnor U10805 (N_10805,N_9128,N_10399);
or U10806 (N_10806,N_9218,N_10102);
and U10807 (N_10807,N_9225,N_9770);
and U10808 (N_10808,N_10253,N_9106);
nand U10809 (N_10809,N_9615,N_9760);
and U10810 (N_10810,N_10461,N_10090);
nor U10811 (N_10811,N_9099,N_9712);
nor U10812 (N_10812,N_10143,N_10398);
or U10813 (N_10813,N_9058,N_10491);
nor U10814 (N_10814,N_9267,N_9994);
and U10815 (N_10815,N_9834,N_9439);
and U10816 (N_10816,N_10255,N_10296);
nand U10817 (N_10817,N_9936,N_10023);
nor U10818 (N_10818,N_9873,N_9597);
xor U10819 (N_10819,N_9035,N_9907);
and U10820 (N_10820,N_10376,N_9962);
nor U10821 (N_10821,N_9691,N_10169);
xnor U10822 (N_10822,N_9290,N_9764);
and U10823 (N_10823,N_9246,N_9482);
nor U10824 (N_10824,N_10016,N_9235);
and U10825 (N_10825,N_9720,N_10264);
and U10826 (N_10826,N_10094,N_9271);
or U10827 (N_10827,N_9678,N_9393);
nand U10828 (N_10828,N_9021,N_9103);
or U10829 (N_10829,N_10423,N_9355);
or U10830 (N_10830,N_9866,N_9749);
and U10831 (N_10831,N_9037,N_9366);
nand U10832 (N_10832,N_9755,N_9274);
nor U10833 (N_10833,N_9424,N_9050);
nand U10834 (N_10834,N_10061,N_9297);
or U10835 (N_10835,N_9107,N_9124);
or U10836 (N_10836,N_9437,N_9476);
and U10837 (N_10837,N_9922,N_10292);
and U10838 (N_10838,N_9249,N_9415);
nor U10839 (N_10839,N_9797,N_10445);
nand U10840 (N_10840,N_10077,N_9665);
nand U10841 (N_10841,N_9078,N_9315);
nand U10842 (N_10842,N_10256,N_9963);
nand U10843 (N_10843,N_9707,N_10214);
and U10844 (N_10844,N_10047,N_9757);
nand U10845 (N_10845,N_10018,N_10354);
nand U10846 (N_10846,N_10381,N_9698);
nand U10847 (N_10847,N_10400,N_9169);
or U10848 (N_10848,N_9150,N_9066);
and U10849 (N_10849,N_9478,N_9193);
nor U10850 (N_10850,N_10020,N_10019);
and U10851 (N_10851,N_10415,N_10076);
nor U10852 (N_10852,N_9252,N_9101);
nand U10853 (N_10853,N_9630,N_9422);
or U10854 (N_10854,N_10410,N_9669);
or U10855 (N_10855,N_9644,N_10483);
and U10856 (N_10856,N_10486,N_9602);
xor U10857 (N_10857,N_10443,N_9259);
xnor U10858 (N_10858,N_9499,N_9569);
nor U10859 (N_10859,N_9350,N_9565);
and U10860 (N_10860,N_9987,N_10003);
xor U10861 (N_10861,N_9593,N_9382);
or U10862 (N_10862,N_9488,N_10345);
and U10863 (N_10863,N_9386,N_9310);
nand U10864 (N_10864,N_10133,N_10305);
nor U10865 (N_10865,N_9543,N_9847);
or U10866 (N_10866,N_9982,N_10160);
and U10867 (N_10867,N_9347,N_9430);
nor U10868 (N_10868,N_10058,N_10437);
or U10869 (N_10869,N_9989,N_9639);
and U10870 (N_10870,N_9508,N_10350);
and U10871 (N_10871,N_9332,N_9617);
and U10872 (N_10872,N_10110,N_9853);
or U10873 (N_10873,N_9138,N_9281);
xnor U10874 (N_10874,N_9807,N_9243);
nor U10875 (N_10875,N_10281,N_10420);
and U10876 (N_10876,N_10247,N_10230);
and U10877 (N_10877,N_10004,N_9278);
xor U10878 (N_10878,N_9284,N_9042);
nand U10879 (N_10879,N_9902,N_9754);
or U10880 (N_10880,N_9298,N_10287);
nor U10881 (N_10881,N_10005,N_9709);
nor U10882 (N_10882,N_9864,N_9795);
nor U10883 (N_10883,N_9319,N_9625);
or U10884 (N_10884,N_10433,N_10074);
nor U10885 (N_10885,N_10427,N_9387);
nor U10886 (N_10886,N_9463,N_10407);
nor U10887 (N_10887,N_9890,N_9477);
nand U10888 (N_10888,N_9333,N_9338);
nor U10889 (N_10889,N_9898,N_10096);
nor U10890 (N_10890,N_9859,N_9061);
and U10891 (N_10891,N_10471,N_9721);
xor U10892 (N_10892,N_9108,N_9918);
or U10893 (N_10893,N_10224,N_9852);
or U10894 (N_10894,N_10374,N_9863);
and U10895 (N_10895,N_9491,N_9584);
xor U10896 (N_10896,N_9519,N_9311);
or U10897 (N_10897,N_9695,N_9282);
nand U10898 (N_10898,N_10325,N_10411);
and U10899 (N_10899,N_9713,N_9670);
and U10900 (N_10900,N_9701,N_10059);
nand U10901 (N_10901,N_9928,N_9406);
nor U10902 (N_10902,N_9923,N_9786);
and U10903 (N_10903,N_9487,N_10320);
nor U10904 (N_10904,N_9830,N_9581);
or U10905 (N_10905,N_9014,N_9710);
nand U10906 (N_10906,N_9002,N_9486);
and U10907 (N_10907,N_10103,N_10465);
or U10908 (N_10908,N_9694,N_10130);
and U10909 (N_10909,N_9024,N_9194);
nand U10910 (N_10910,N_9131,N_10212);
nand U10911 (N_10911,N_9026,N_9089);
or U10912 (N_10912,N_9627,N_9740);
nor U10913 (N_10913,N_9416,N_9079);
nor U10914 (N_10914,N_9048,N_9775);
and U10915 (N_10915,N_9429,N_9134);
nand U10916 (N_10916,N_9601,N_9363);
nor U10917 (N_10917,N_10431,N_10177);
and U10918 (N_10918,N_9075,N_10487);
nand U10919 (N_10919,N_9663,N_9588);
nand U10920 (N_10920,N_10185,N_9495);
nor U10921 (N_10921,N_9762,N_9527);
and U10922 (N_10922,N_10216,N_9484);
nor U10923 (N_10923,N_9299,N_10179);
and U10924 (N_10924,N_9213,N_9470);
nor U10925 (N_10925,N_9855,N_9277);
and U10926 (N_10926,N_9154,N_9168);
nand U10927 (N_10927,N_10207,N_9148);
or U10928 (N_10928,N_9105,N_9958);
or U10929 (N_10929,N_9069,N_9348);
or U10930 (N_10930,N_9456,N_9981);
or U10931 (N_10931,N_9185,N_9145);
nand U10932 (N_10932,N_9967,N_10457);
nor U10933 (N_10933,N_9507,N_9440);
or U10934 (N_10934,N_10222,N_9785);
nor U10935 (N_10935,N_9184,N_10413);
and U10936 (N_10936,N_10246,N_10332);
or U10937 (N_10937,N_10468,N_9419);
or U10938 (N_10938,N_9199,N_10390);
nand U10939 (N_10939,N_9238,N_10206);
nor U10940 (N_10940,N_10310,N_10459);
or U10941 (N_10941,N_10294,N_9082);
nor U10942 (N_10942,N_10244,N_10106);
and U10943 (N_10943,N_9196,N_9202);
xor U10944 (N_10944,N_9960,N_9736);
nand U10945 (N_10945,N_9104,N_9114);
nand U10946 (N_10946,N_9265,N_9450);
and U10947 (N_10947,N_9049,N_9975);
nand U10948 (N_10948,N_9251,N_9126);
nor U10949 (N_10949,N_9706,N_9717);
or U10950 (N_10950,N_9323,N_9328);
nand U10951 (N_10951,N_9221,N_9684);
or U10952 (N_10952,N_9761,N_10189);
xor U10953 (N_10953,N_10171,N_9592);
and U10954 (N_10954,N_10460,N_9330);
nor U10955 (N_10955,N_9500,N_10119);
nor U10956 (N_10956,N_9451,N_10493);
nand U10957 (N_10957,N_9526,N_10151);
or U10958 (N_10958,N_10234,N_9181);
nand U10959 (N_10959,N_10152,N_9275);
or U10960 (N_10960,N_9642,N_9999);
nor U10961 (N_10961,N_9445,N_9723);
or U10962 (N_10962,N_10174,N_9773);
and U10963 (N_10963,N_9244,N_10402);
nor U10964 (N_10964,N_9747,N_10201);
nand U10965 (N_10965,N_10316,N_9897);
nand U10966 (N_10966,N_9420,N_9191);
and U10967 (N_10967,N_9044,N_9728);
and U10968 (N_10968,N_9034,N_9899);
or U10969 (N_10969,N_9572,N_9915);
or U10970 (N_10970,N_9398,N_9951);
xor U10971 (N_10971,N_9077,N_9286);
nor U10972 (N_10972,N_9369,N_9129);
nand U10973 (N_10973,N_9752,N_10250);
nand U10974 (N_10974,N_10101,N_9208);
nand U10975 (N_10975,N_9742,N_10037);
and U10976 (N_10976,N_10301,N_9827);
and U10977 (N_10977,N_9798,N_10155);
xnor U10978 (N_10978,N_9745,N_10391);
nand U10979 (N_10979,N_9392,N_9547);
or U10980 (N_10980,N_10485,N_10356);
nand U10981 (N_10981,N_9492,N_9835);
nor U10982 (N_10982,N_10205,N_9763);
xor U10983 (N_10983,N_9553,N_9388);
and U10984 (N_10984,N_10478,N_10442);
nor U10985 (N_10985,N_10236,N_10451);
nand U10986 (N_10986,N_9816,N_9861);
or U10987 (N_10987,N_9241,N_9832);
or U10988 (N_10988,N_9654,N_9784);
and U10989 (N_10989,N_9291,N_9481);
and U10990 (N_10990,N_9711,N_9344);
and U10991 (N_10991,N_9521,N_10318);
nand U10992 (N_10992,N_9237,N_9367);
xor U10993 (N_10993,N_9188,N_10162);
nor U10994 (N_10994,N_10017,N_9460);
and U10995 (N_10995,N_9626,N_10229);
and U10996 (N_10996,N_10154,N_9746);
and U10997 (N_10997,N_10449,N_10336);
nand U10998 (N_10998,N_9796,N_9980);
and U10999 (N_10999,N_9410,N_9880);
and U11000 (N_11000,N_10084,N_9242);
nor U11001 (N_11001,N_9146,N_10144);
nand U11002 (N_11002,N_9562,N_9186);
or U11003 (N_11003,N_10120,N_9821);
nor U11004 (N_11004,N_9435,N_9538);
nor U11005 (N_11005,N_9966,N_10232);
and U11006 (N_11006,N_10012,N_9229);
nor U11007 (N_11007,N_10394,N_9612);
nand U11008 (N_11008,N_9614,N_10484);
or U11009 (N_11009,N_9959,N_9313);
nor U11010 (N_11010,N_9651,N_10285);
or U11011 (N_11011,N_9865,N_9473);
xnor U11012 (N_11012,N_9517,N_9814);
xor U11013 (N_11013,N_10109,N_9542);
or U11014 (N_11014,N_10278,N_10083);
nor U11015 (N_11015,N_9791,N_9636);
and U11016 (N_11016,N_10495,N_9590);
nand U11017 (N_11017,N_9808,N_10293);
xor U11018 (N_11018,N_10235,N_9144);
or U11019 (N_11019,N_9127,N_10226);
and U11020 (N_11020,N_9758,N_9029);
nand U11021 (N_11021,N_9418,N_9025);
nor U11022 (N_11022,N_9632,N_9589);
and U11023 (N_11023,N_10298,N_10149);
xnor U11024 (N_11024,N_9903,N_9474);
nor U11025 (N_11025,N_10359,N_9161);
nor U11026 (N_11026,N_10159,N_9309);
or U11027 (N_11027,N_9287,N_10382);
or U11028 (N_11028,N_9708,N_9204);
and U11029 (N_11029,N_9397,N_10383);
and U11030 (N_11030,N_10323,N_9599);
nor U11031 (N_11031,N_9577,N_9017);
and U11032 (N_11032,N_9909,N_9288);
or U11033 (N_11033,N_10252,N_10334);
nand U11034 (N_11034,N_9893,N_10283);
and U11035 (N_11035,N_9743,N_10052);
and U11036 (N_11036,N_9515,N_10217);
nor U11037 (N_11037,N_9596,N_10125);
nand U11038 (N_11038,N_9027,N_9753);
nand U11039 (N_11039,N_10389,N_9671);
xnor U11040 (N_11040,N_9595,N_9719);
nand U11041 (N_11041,N_9607,N_9680);
nor U11042 (N_11042,N_10072,N_10131);
nand U11043 (N_11043,N_10122,N_9917);
or U11044 (N_11044,N_9774,N_9895);
or U11045 (N_11045,N_10091,N_10157);
and U11046 (N_11046,N_9302,N_10186);
and U11047 (N_11047,N_10193,N_9093);
nor U11048 (N_11048,N_10438,N_9594);
nor U11049 (N_11049,N_9984,N_9767);
or U11050 (N_11050,N_10167,N_9953);
nor U11051 (N_11051,N_9140,N_10397);
and U11052 (N_11052,N_10165,N_9452);
or U11053 (N_11053,N_9539,N_9657);
and U11054 (N_11054,N_9052,N_9226);
or U11055 (N_11055,N_9974,N_10417);
and U11056 (N_11056,N_10188,N_10251);
xor U11057 (N_11057,N_10139,N_9552);
nor U11058 (N_11058,N_9647,N_9011);
nor U11059 (N_11059,N_9081,N_9732);
nand U11060 (N_11060,N_9095,N_9509);
and U11061 (N_11061,N_9993,N_9180);
nand U11062 (N_11062,N_10453,N_9233);
or U11063 (N_11063,N_9520,N_9222);
nand U11064 (N_11064,N_10387,N_9257);
nand U11065 (N_11065,N_9881,N_9793);
and U11066 (N_11066,N_10218,N_9985);
nand U11067 (N_11067,N_10223,N_9351);
nand U11068 (N_11068,N_9354,N_9883);
nor U11069 (N_11069,N_10353,N_10114);
and U11070 (N_11070,N_9423,N_9438);
nor U11071 (N_11071,N_9551,N_10441);
and U11072 (N_11072,N_9163,N_9668);
nand U11073 (N_11073,N_9459,N_9805);
nand U11074 (N_11074,N_9727,N_9295);
nand U11075 (N_11075,N_9724,N_10203);
or U11076 (N_11076,N_10118,N_10466);
nor U11077 (N_11077,N_9400,N_10499);
nor U11078 (N_11078,N_9535,N_9891);
nor U11079 (N_11079,N_9849,N_9765);
and U11080 (N_11080,N_10425,N_10211);
and U11081 (N_11081,N_10488,N_9634);
or U11082 (N_11082,N_10271,N_9444);
and U11083 (N_11083,N_10269,N_10496);
nor U11084 (N_11084,N_9245,N_9924);
xnor U11085 (N_11085,N_9789,N_9931);
or U11086 (N_11086,N_10426,N_10093);
nor U11087 (N_11087,N_9856,N_9667);
nor U11088 (N_11088,N_9558,N_9432);
nor U11089 (N_11089,N_9307,N_10198);
and U11090 (N_11090,N_9370,N_9293);
and U11091 (N_11091,N_10274,N_9603);
nand U11092 (N_11092,N_10307,N_9469);
nor U11093 (N_11093,N_9268,N_9498);
or U11094 (N_11094,N_9111,N_9575);
and U11095 (N_11095,N_9327,N_9098);
and U11096 (N_11096,N_9912,N_9009);
and U11097 (N_11097,N_10452,N_9152);
and U11098 (N_11098,N_9461,N_9276);
and U11099 (N_11099,N_9471,N_9378);
or U11100 (N_11100,N_9744,N_9531);
or U11101 (N_11101,N_9182,N_9806);
nand U11102 (N_11102,N_9731,N_9666);
nand U11103 (N_11103,N_10038,N_9776);
nor U11104 (N_11104,N_9702,N_10404);
nand U11105 (N_11105,N_9813,N_10371);
and U11106 (N_11106,N_9563,N_10087);
or U11107 (N_11107,N_10286,N_9250);
and U11108 (N_11108,N_9013,N_10172);
xnor U11109 (N_11109,N_9391,N_9877);
or U11110 (N_11110,N_9394,N_10408);
nor U11111 (N_11111,N_10127,N_9038);
or U11112 (N_11112,N_9428,N_10024);
nand U11113 (N_11113,N_9300,N_9950);
or U11114 (N_11114,N_10289,N_9620);
nand U11115 (N_11115,N_9817,N_9518);
nor U11116 (N_11116,N_10412,N_9659);
and U11117 (N_11117,N_10362,N_9686);
or U11118 (N_11118,N_10134,N_10221);
nor U11119 (N_11119,N_9164,N_9155);
and U11120 (N_11120,N_9699,N_10327);
nor U11121 (N_11121,N_9815,N_10330);
nor U11122 (N_11122,N_9692,N_9102);
or U11123 (N_11123,N_9331,N_9537);
nand U11124 (N_11124,N_9522,N_10041);
xnor U11125 (N_11125,N_9878,N_9640);
and U11126 (N_11126,N_9616,N_10476);
nand U11127 (N_11127,N_10297,N_9132);
and U11128 (N_11128,N_9528,N_10115);
nor U11129 (N_11129,N_9679,N_9901);
nor U11130 (N_11130,N_10393,N_10481);
nand U11131 (N_11131,N_9381,N_10097);
and U11132 (N_11132,N_10419,N_9254);
nor U11133 (N_11133,N_9777,N_10163);
nand U11134 (N_11134,N_9321,N_9949);
and U11135 (N_11135,N_9072,N_10270);
nand U11136 (N_11136,N_9570,N_10357);
or U11137 (N_11137,N_10195,N_10099);
or U11138 (N_11138,N_9270,N_9624);
or U11139 (N_11139,N_10181,N_10036);
nor U11140 (N_11140,N_10009,N_9887);
nand U11141 (N_11141,N_10479,N_10117);
xor U11142 (N_11142,N_9122,N_9583);
or U11143 (N_11143,N_9510,N_9156);
or U11144 (N_11144,N_9787,N_10284);
and U11145 (N_11145,N_9506,N_10128);
nand U11146 (N_11146,N_9260,N_9792);
nand U11147 (N_11147,N_9000,N_9316);
nor U11148 (N_11148,N_10063,N_9722);
nand U11149 (N_11149,N_9540,N_9115);
nor U11150 (N_11150,N_9253,N_10153);
nor U11151 (N_11151,N_10329,N_9117);
nor U11152 (N_11152,N_10385,N_9729);
and U11153 (N_11153,N_9738,N_9768);
or U11154 (N_11154,N_9084,N_9567);
or U11155 (N_11155,N_9109,N_10187);
or U11156 (N_11156,N_9972,N_9664);
nor U11157 (N_11157,N_9228,N_9803);
or U11158 (N_11158,N_10279,N_9673);
or U11159 (N_11159,N_10026,N_9384);
nor U11160 (N_11160,N_9113,N_9869);
nand U11161 (N_11161,N_10261,N_9556);
nand U11162 (N_11162,N_10494,N_9137);
and U11163 (N_11163,N_9273,N_9094);
nand U11164 (N_11164,N_9047,N_10428);
or U11165 (N_11165,N_9322,N_9910);
or U11166 (N_11166,N_9944,N_9831);
nor U11167 (N_11167,N_9652,N_9549);
and U11168 (N_11168,N_10352,N_9605);
xor U11169 (N_11169,N_9568,N_10112);
or U11170 (N_11170,N_9574,N_10060);
and U11171 (N_11171,N_9598,N_9576);
nor U11172 (N_11172,N_9824,N_9810);
nand U11173 (N_11173,N_9851,N_10348);
and U11174 (N_11174,N_9546,N_10042);
nor U11175 (N_11175,N_9206,N_9263);
or U11176 (N_11176,N_9173,N_10064);
and U11177 (N_11177,N_10199,N_10456);
nor U11178 (N_11178,N_9214,N_9927);
and U11179 (N_11179,N_9490,N_9135);
or U11180 (N_11180,N_10014,N_9600);
and U11181 (N_11181,N_10321,N_10182);
nand U11182 (N_11182,N_10414,N_9921);
and U11183 (N_11183,N_9190,N_10276);
and U11184 (N_11184,N_9142,N_9970);
or U11185 (N_11185,N_10446,N_10380);
and U11186 (N_11186,N_9376,N_9876);
or U11187 (N_11187,N_10384,N_9085);
and U11188 (N_11188,N_10051,N_9677);
or U11189 (N_11189,N_9472,N_9929);
xor U11190 (N_11190,N_9844,N_9530);
or U11191 (N_11191,N_9750,N_9494);
nor U11192 (N_11192,N_9443,N_10242);
nand U11193 (N_11193,N_9633,N_9938);
or U11194 (N_11194,N_9375,N_9158);
xor U11195 (N_11195,N_9610,N_10183);
nand U11196 (N_11196,N_9483,N_10272);
nand U11197 (N_11197,N_10006,N_10436);
or U11198 (N_11198,N_10013,N_9818);
and U11199 (N_11199,N_9629,N_9829);
and U11200 (N_11200,N_9171,N_9325);
xor U11201 (N_11201,N_9373,N_9645);
nor U11202 (N_11202,N_9417,N_9256);
xnor U11203 (N_11203,N_9030,N_9660);
or U11204 (N_11204,N_9782,N_10141);
nor U11205 (N_11205,N_9216,N_10104);
or U11206 (N_11206,N_9580,N_9613);
nor U11207 (N_11207,N_10032,N_9305);
and U11208 (N_11208,N_9523,N_10107);
and U11209 (N_11209,N_9361,N_10455);
nand U11210 (N_11210,N_9799,N_9964);
nor U11211 (N_11211,N_9641,N_10129);
nand U11212 (N_11212,N_9908,N_9638);
xor U11213 (N_11213,N_9425,N_10424);
or U11214 (N_11214,N_10477,N_9059);
nor U11215 (N_11215,N_10158,N_9408);
nand U11216 (N_11216,N_9215,N_9176);
xor U11217 (N_11217,N_9886,N_9289);
or U11218 (N_11218,N_9726,N_9548);
xor U11219 (N_11219,N_9609,N_9407);
nand U11220 (N_11220,N_9159,N_9166);
nand U11221 (N_11221,N_10176,N_9379);
nor U11222 (N_11222,N_10050,N_9604);
and U11223 (N_11223,N_10121,N_9591);
xor U11224 (N_11224,N_9183,N_10219);
xor U11225 (N_11225,N_10111,N_9718);
xor U11226 (N_11226,N_10355,N_9566);
nand U11227 (N_11227,N_9942,N_9828);
nand U11228 (N_11228,N_9837,N_10142);
nand U11229 (N_11229,N_9212,N_9211);
nand U11230 (N_11230,N_9004,N_9149);
or U11231 (N_11231,N_9919,N_10100);
xnor U11232 (N_11232,N_9688,N_9968);
nor U11233 (N_11233,N_9073,N_9359);
and U11234 (N_11234,N_10262,N_9248);
or U11235 (N_11235,N_9405,N_10317);
xor U11236 (N_11236,N_9933,N_9431);
or U11237 (N_11237,N_10025,N_9937);
nor U11238 (N_11238,N_9656,N_9992);
and U11239 (N_11239,N_9337,N_9412);
and U11240 (N_11240,N_10243,N_9033);
and U11241 (N_11241,N_10458,N_9646);
and U11242 (N_11242,N_10239,N_9544);
or U11243 (N_11243,N_9941,N_9956);
or U11244 (N_11244,N_9318,N_10351);
nand U11245 (N_11245,N_10027,N_9434);
nand U11246 (N_11246,N_9436,N_9839);
nor U11247 (N_11247,N_10178,N_10275);
and U11248 (N_11248,N_9683,N_9462);
and U11249 (N_11249,N_9195,N_10135);
nand U11250 (N_11250,N_9374,N_10254);
xor U11251 (N_11251,N_9423,N_9410);
xnor U11252 (N_11252,N_9118,N_10454);
and U11253 (N_11253,N_9707,N_9869);
nand U11254 (N_11254,N_10343,N_10217);
xnor U11255 (N_11255,N_9241,N_9316);
nor U11256 (N_11256,N_9459,N_9457);
xnor U11257 (N_11257,N_10435,N_10480);
xor U11258 (N_11258,N_10343,N_10423);
or U11259 (N_11259,N_10459,N_10016);
nand U11260 (N_11260,N_10409,N_10152);
and U11261 (N_11261,N_9429,N_9547);
nor U11262 (N_11262,N_10297,N_9416);
nor U11263 (N_11263,N_10304,N_9171);
or U11264 (N_11264,N_9152,N_9601);
and U11265 (N_11265,N_10456,N_10358);
or U11266 (N_11266,N_9021,N_9140);
or U11267 (N_11267,N_10416,N_9518);
nor U11268 (N_11268,N_10213,N_10278);
and U11269 (N_11269,N_10186,N_9403);
or U11270 (N_11270,N_9348,N_9771);
or U11271 (N_11271,N_10363,N_9470);
xnor U11272 (N_11272,N_9675,N_10295);
and U11273 (N_11273,N_9024,N_9013);
nor U11274 (N_11274,N_9252,N_10256);
nor U11275 (N_11275,N_9543,N_10346);
nor U11276 (N_11276,N_9969,N_10317);
nand U11277 (N_11277,N_9291,N_10311);
or U11278 (N_11278,N_9326,N_10182);
nand U11279 (N_11279,N_9994,N_9251);
nand U11280 (N_11280,N_9057,N_9721);
and U11281 (N_11281,N_9079,N_9828);
nor U11282 (N_11282,N_10143,N_10237);
xnor U11283 (N_11283,N_9478,N_10437);
or U11284 (N_11284,N_9818,N_10217);
nand U11285 (N_11285,N_10445,N_9783);
or U11286 (N_11286,N_9529,N_9627);
nand U11287 (N_11287,N_9709,N_10089);
and U11288 (N_11288,N_9621,N_10378);
nand U11289 (N_11289,N_9954,N_9090);
or U11290 (N_11290,N_9437,N_9267);
and U11291 (N_11291,N_10207,N_9348);
or U11292 (N_11292,N_9060,N_10218);
nand U11293 (N_11293,N_9988,N_9251);
nor U11294 (N_11294,N_9853,N_9915);
and U11295 (N_11295,N_9831,N_10101);
or U11296 (N_11296,N_9555,N_9148);
and U11297 (N_11297,N_9357,N_9680);
and U11298 (N_11298,N_10152,N_9726);
xor U11299 (N_11299,N_10432,N_10088);
nand U11300 (N_11300,N_9707,N_10226);
xor U11301 (N_11301,N_9206,N_9067);
nor U11302 (N_11302,N_9245,N_9197);
xor U11303 (N_11303,N_10439,N_9378);
xnor U11304 (N_11304,N_10170,N_9789);
nand U11305 (N_11305,N_9990,N_10278);
and U11306 (N_11306,N_9459,N_10004);
xor U11307 (N_11307,N_9136,N_10225);
nor U11308 (N_11308,N_10448,N_9841);
xor U11309 (N_11309,N_10188,N_10411);
nor U11310 (N_11310,N_10390,N_9464);
nand U11311 (N_11311,N_9379,N_9124);
nor U11312 (N_11312,N_10077,N_9944);
xor U11313 (N_11313,N_9915,N_9626);
nor U11314 (N_11314,N_9460,N_10399);
nand U11315 (N_11315,N_9451,N_9527);
or U11316 (N_11316,N_9674,N_10352);
and U11317 (N_11317,N_10271,N_10299);
nor U11318 (N_11318,N_9834,N_10150);
or U11319 (N_11319,N_10154,N_9904);
and U11320 (N_11320,N_9244,N_9972);
nor U11321 (N_11321,N_10498,N_9375);
and U11322 (N_11322,N_9724,N_9736);
xor U11323 (N_11323,N_9312,N_9096);
and U11324 (N_11324,N_9042,N_10364);
nor U11325 (N_11325,N_9387,N_9293);
and U11326 (N_11326,N_10061,N_9600);
nor U11327 (N_11327,N_9167,N_10100);
or U11328 (N_11328,N_9418,N_9904);
and U11329 (N_11329,N_9737,N_10318);
nor U11330 (N_11330,N_9050,N_9446);
nor U11331 (N_11331,N_10223,N_10166);
nor U11332 (N_11332,N_9941,N_9605);
and U11333 (N_11333,N_9143,N_9597);
xnor U11334 (N_11334,N_10386,N_9828);
or U11335 (N_11335,N_10045,N_10292);
nor U11336 (N_11336,N_10108,N_9918);
and U11337 (N_11337,N_9605,N_10397);
and U11338 (N_11338,N_9342,N_10385);
or U11339 (N_11339,N_9738,N_9312);
nand U11340 (N_11340,N_9839,N_9230);
and U11341 (N_11341,N_10282,N_9426);
nor U11342 (N_11342,N_10249,N_9936);
or U11343 (N_11343,N_9735,N_9224);
and U11344 (N_11344,N_10137,N_10432);
xor U11345 (N_11345,N_9371,N_9933);
nand U11346 (N_11346,N_9617,N_10246);
nor U11347 (N_11347,N_9030,N_9522);
xnor U11348 (N_11348,N_9728,N_10115);
nor U11349 (N_11349,N_10475,N_9696);
and U11350 (N_11350,N_10197,N_10102);
and U11351 (N_11351,N_10025,N_9054);
xor U11352 (N_11352,N_9028,N_9864);
nor U11353 (N_11353,N_9817,N_9891);
and U11354 (N_11354,N_10095,N_9816);
nand U11355 (N_11355,N_9306,N_10392);
or U11356 (N_11356,N_9174,N_10385);
nor U11357 (N_11357,N_9298,N_9511);
or U11358 (N_11358,N_9467,N_9440);
nand U11359 (N_11359,N_9304,N_10059);
nor U11360 (N_11360,N_9756,N_9356);
nand U11361 (N_11361,N_9065,N_9005);
nor U11362 (N_11362,N_9941,N_9426);
xnor U11363 (N_11363,N_9460,N_10241);
nor U11364 (N_11364,N_9475,N_10156);
and U11365 (N_11365,N_10240,N_9362);
nor U11366 (N_11366,N_10106,N_9016);
or U11367 (N_11367,N_9627,N_9572);
nand U11368 (N_11368,N_10392,N_10337);
nand U11369 (N_11369,N_9962,N_9475);
nand U11370 (N_11370,N_9045,N_10485);
xnor U11371 (N_11371,N_10249,N_10429);
and U11372 (N_11372,N_9309,N_9377);
nand U11373 (N_11373,N_10200,N_9071);
or U11374 (N_11374,N_9956,N_9085);
nand U11375 (N_11375,N_9728,N_10263);
nand U11376 (N_11376,N_9137,N_9296);
xnor U11377 (N_11377,N_9795,N_9432);
xnor U11378 (N_11378,N_9163,N_9952);
or U11379 (N_11379,N_9112,N_9094);
nor U11380 (N_11380,N_10249,N_9728);
or U11381 (N_11381,N_9857,N_9151);
or U11382 (N_11382,N_10342,N_10387);
or U11383 (N_11383,N_9266,N_10375);
and U11384 (N_11384,N_10494,N_10085);
nor U11385 (N_11385,N_9378,N_9327);
nor U11386 (N_11386,N_10381,N_10176);
nor U11387 (N_11387,N_9681,N_9934);
or U11388 (N_11388,N_9535,N_9214);
and U11389 (N_11389,N_10011,N_10170);
and U11390 (N_11390,N_9718,N_9745);
nand U11391 (N_11391,N_9765,N_9426);
and U11392 (N_11392,N_9228,N_9030);
nand U11393 (N_11393,N_9716,N_10478);
nor U11394 (N_11394,N_9273,N_9762);
nor U11395 (N_11395,N_9053,N_10174);
and U11396 (N_11396,N_9772,N_9730);
and U11397 (N_11397,N_9553,N_9711);
nand U11398 (N_11398,N_9631,N_9855);
or U11399 (N_11399,N_9703,N_9863);
nor U11400 (N_11400,N_10474,N_9115);
or U11401 (N_11401,N_9131,N_10148);
nor U11402 (N_11402,N_9065,N_9168);
or U11403 (N_11403,N_9248,N_9927);
nor U11404 (N_11404,N_9256,N_9840);
or U11405 (N_11405,N_10347,N_9188);
nand U11406 (N_11406,N_9121,N_9861);
nand U11407 (N_11407,N_9891,N_10370);
nor U11408 (N_11408,N_10480,N_9887);
nand U11409 (N_11409,N_9046,N_9050);
nor U11410 (N_11410,N_10003,N_9427);
or U11411 (N_11411,N_9350,N_9065);
nor U11412 (N_11412,N_9545,N_9527);
nor U11413 (N_11413,N_10022,N_9382);
nor U11414 (N_11414,N_10261,N_10266);
nor U11415 (N_11415,N_9391,N_10264);
nor U11416 (N_11416,N_10336,N_9501);
xnor U11417 (N_11417,N_9346,N_9180);
and U11418 (N_11418,N_9505,N_9947);
nor U11419 (N_11419,N_9851,N_10151);
and U11420 (N_11420,N_9841,N_9306);
nor U11421 (N_11421,N_9415,N_9235);
and U11422 (N_11422,N_9982,N_9979);
or U11423 (N_11423,N_9224,N_9937);
or U11424 (N_11424,N_9281,N_10016);
or U11425 (N_11425,N_9616,N_10083);
or U11426 (N_11426,N_10150,N_9732);
or U11427 (N_11427,N_10082,N_9205);
nand U11428 (N_11428,N_9170,N_10369);
nand U11429 (N_11429,N_9966,N_9218);
nand U11430 (N_11430,N_9912,N_10054);
and U11431 (N_11431,N_9525,N_9783);
xor U11432 (N_11432,N_9138,N_10381);
nor U11433 (N_11433,N_10493,N_10252);
or U11434 (N_11434,N_10291,N_9093);
nor U11435 (N_11435,N_10411,N_9275);
nor U11436 (N_11436,N_9542,N_9773);
nor U11437 (N_11437,N_9302,N_9480);
xnor U11438 (N_11438,N_9429,N_9856);
nand U11439 (N_11439,N_9090,N_9052);
xor U11440 (N_11440,N_10012,N_10345);
nand U11441 (N_11441,N_9591,N_10498);
nand U11442 (N_11442,N_9323,N_9994);
and U11443 (N_11443,N_9174,N_10294);
xor U11444 (N_11444,N_10054,N_9515);
xnor U11445 (N_11445,N_10349,N_9997);
nor U11446 (N_11446,N_9935,N_9533);
nand U11447 (N_11447,N_10054,N_10217);
or U11448 (N_11448,N_10362,N_9142);
or U11449 (N_11449,N_9425,N_10331);
or U11450 (N_11450,N_9494,N_10314);
or U11451 (N_11451,N_9686,N_9055);
or U11452 (N_11452,N_9393,N_9545);
or U11453 (N_11453,N_9156,N_10063);
nand U11454 (N_11454,N_10201,N_10092);
nand U11455 (N_11455,N_9040,N_10399);
nor U11456 (N_11456,N_9724,N_9322);
nand U11457 (N_11457,N_9433,N_10315);
nor U11458 (N_11458,N_10037,N_9639);
nor U11459 (N_11459,N_10351,N_10472);
nor U11460 (N_11460,N_10021,N_9939);
or U11461 (N_11461,N_9267,N_9495);
nor U11462 (N_11462,N_9938,N_9710);
and U11463 (N_11463,N_9726,N_9770);
nor U11464 (N_11464,N_10009,N_9674);
and U11465 (N_11465,N_9834,N_10426);
nor U11466 (N_11466,N_10299,N_9194);
and U11467 (N_11467,N_9226,N_10302);
or U11468 (N_11468,N_9894,N_9187);
nor U11469 (N_11469,N_9739,N_10107);
or U11470 (N_11470,N_9845,N_10140);
and U11471 (N_11471,N_10120,N_9303);
and U11472 (N_11472,N_10417,N_9556);
or U11473 (N_11473,N_9329,N_9692);
nor U11474 (N_11474,N_9879,N_9294);
nor U11475 (N_11475,N_10468,N_9505);
nor U11476 (N_11476,N_9479,N_10019);
nor U11477 (N_11477,N_9445,N_9424);
and U11478 (N_11478,N_9973,N_10298);
nand U11479 (N_11479,N_10204,N_9610);
or U11480 (N_11480,N_9706,N_10432);
and U11481 (N_11481,N_10155,N_9544);
xnor U11482 (N_11482,N_10449,N_10167);
or U11483 (N_11483,N_9755,N_9221);
nor U11484 (N_11484,N_9045,N_9512);
nand U11485 (N_11485,N_10240,N_9882);
nor U11486 (N_11486,N_9841,N_9240);
xor U11487 (N_11487,N_10025,N_10270);
and U11488 (N_11488,N_10113,N_9044);
nor U11489 (N_11489,N_9445,N_10067);
or U11490 (N_11490,N_9229,N_10159);
and U11491 (N_11491,N_10238,N_9614);
or U11492 (N_11492,N_9818,N_9878);
nor U11493 (N_11493,N_9232,N_10218);
nor U11494 (N_11494,N_9782,N_9596);
nand U11495 (N_11495,N_9112,N_9283);
nand U11496 (N_11496,N_10297,N_9640);
or U11497 (N_11497,N_10341,N_9728);
xor U11498 (N_11498,N_9875,N_9451);
and U11499 (N_11499,N_10262,N_9497);
and U11500 (N_11500,N_9438,N_10321);
and U11501 (N_11501,N_9216,N_10385);
nor U11502 (N_11502,N_9528,N_9320);
nand U11503 (N_11503,N_9871,N_10320);
nor U11504 (N_11504,N_9456,N_9750);
or U11505 (N_11505,N_9222,N_9509);
nor U11506 (N_11506,N_9087,N_9635);
nand U11507 (N_11507,N_9902,N_9445);
and U11508 (N_11508,N_10497,N_9415);
nor U11509 (N_11509,N_10235,N_9742);
or U11510 (N_11510,N_9151,N_9245);
nand U11511 (N_11511,N_10267,N_9596);
nor U11512 (N_11512,N_10370,N_9986);
nand U11513 (N_11513,N_9704,N_9500);
and U11514 (N_11514,N_9052,N_9404);
or U11515 (N_11515,N_10420,N_10383);
nand U11516 (N_11516,N_9107,N_9811);
xor U11517 (N_11517,N_9606,N_10069);
and U11518 (N_11518,N_10317,N_9248);
xor U11519 (N_11519,N_10288,N_10023);
or U11520 (N_11520,N_9385,N_9577);
xnor U11521 (N_11521,N_9007,N_9829);
xnor U11522 (N_11522,N_9394,N_9339);
xor U11523 (N_11523,N_10227,N_9902);
and U11524 (N_11524,N_10203,N_10349);
or U11525 (N_11525,N_9660,N_9384);
nand U11526 (N_11526,N_9448,N_10260);
and U11527 (N_11527,N_9880,N_10204);
or U11528 (N_11528,N_9190,N_9823);
nor U11529 (N_11529,N_9632,N_9358);
xor U11530 (N_11530,N_9721,N_10079);
xor U11531 (N_11531,N_10127,N_9557);
nor U11532 (N_11532,N_9434,N_10236);
and U11533 (N_11533,N_9186,N_9325);
nor U11534 (N_11534,N_9063,N_9835);
xnor U11535 (N_11535,N_9965,N_9613);
nand U11536 (N_11536,N_9331,N_9129);
xor U11537 (N_11537,N_9769,N_10246);
nand U11538 (N_11538,N_9385,N_9404);
and U11539 (N_11539,N_10010,N_9721);
nor U11540 (N_11540,N_9780,N_9988);
and U11541 (N_11541,N_9547,N_9344);
nand U11542 (N_11542,N_9710,N_9744);
nor U11543 (N_11543,N_9203,N_9446);
nor U11544 (N_11544,N_10186,N_10075);
nor U11545 (N_11545,N_10237,N_10387);
or U11546 (N_11546,N_10325,N_9432);
or U11547 (N_11547,N_9462,N_10235);
nand U11548 (N_11548,N_9220,N_9860);
nor U11549 (N_11549,N_9431,N_9963);
nand U11550 (N_11550,N_9116,N_9491);
and U11551 (N_11551,N_9715,N_9683);
nand U11552 (N_11552,N_9921,N_10499);
nand U11553 (N_11553,N_9747,N_9393);
nor U11554 (N_11554,N_10095,N_10098);
or U11555 (N_11555,N_9216,N_9648);
and U11556 (N_11556,N_10277,N_9899);
nand U11557 (N_11557,N_9296,N_9234);
or U11558 (N_11558,N_10465,N_10374);
or U11559 (N_11559,N_9994,N_10203);
nand U11560 (N_11560,N_9495,N_10269);
or U11561 (N_11561,N_9331,N_10183);
nor U11562 (N_11562,N_9422,N_10458);
nand U11563 (N_11563,N_9365,N_9800);
xor U11564 (N_11564,N_9245,N_9539);
nor U11565 (N_11565,N_10331,N_9929);
nor U11566 (N_11566,N_10184,N_9664);
nand U11567 (N_11567,N_10135,N_10283);
xnor U11568 (N_11568,N_9110,N_9479);
nor U11569 (N_11569,N_9058,N_10141);
nor U11570 (N_11570,N_10258,N_10244);
or U11571 (N_11571,N_9765,N_9766);
xor U11572 (N_11572,N_9847,N_10303);
nor U11573 (N_11573,N_9142,N_9107);
or U11574 (N_11574,N_9516,N_9858);
or U11575 (N_11575,N_9335,N_9438);
nand U11576 (N_11576,N_9539,N_9832);
nand U11577 (N_11577,N_9545,N_10108);
nor U11578 (N_11578,N_9905,N_10012);
nor U11579 (N_11579,N_9181,N_9856);
nand U11580 (N_11580,N_9103,N_9554);
nor U11581 (N_11581,N_10268,N_10463);
and U11582 (N_11582,N_9822,N_10498);
or U11583 (N_11583,N_10270,N_10481);
and U11584 (N_11584,N_9659,N_9406);
nand U11585 (N_11585,N_9652,N_10217);
or U11586 (N_11586,N_9923,N_9444);
nand U11587 (N_11587,N_10288,N_9357);
and U11588 (N_11588,N_9995,N_9257);
or U11589 (N_11589,N_9290,N_9496);
and U11590 (N_11590,N_9933,N_10330);
nand U11591 (N_11591,N_9041,N_9305);
nor U11592 (N_11592,N_10217,N_9111);
or U11593 (N_11593,N_9801,N_10292);
nand U11594 (N_11594,N_10209,N_9621);
and U11595 (N_11595,N_9479,N_10352);
nor U11596 (N_11596,N_9225,N_10258);
xor U11597 (N_11597,N_9490,N_9487);
and U11598 (N_11598,N_9451,N_9872);
and U11599 (N_11599,N_9061,N_9131);
xnor U11600 (N_11600,N_9346,N_10332);
or U11601 (N_11601,N_9696,N_9435);
nor U11602 (N_11602,N_10231,N_9216);
xnor U11603 (N_11603,N_9857,N_10109);
nand U11604 (N_11604,N_9092,N_10009);
nand U11605 (N_11605,N_10075,N_9764);
and U11606 (N_11606,N_10355,N_9666);
nand U11607 (N_11607,N_10172,N_9082);
or U11608 (N_11608,N_9249,N_10398);
and U11609 (N_11609,N_9668,N_10082);
xor U11610 (N_11610,N_9133,N_10232);
nor U11611 (N_11611,N_9008,N_9088);
and U11612 (N_11612,N_9002,N_10114);
nand U11613 (N_11613,N_9132,N_10121);
xor U11614 (N_11614,N_9154,N_9469);
and U11615 (N_11615,N_10210,N_9071);
nand U11616 (N_11616,N_9436,N_9064);
and U11617 (N_11617,N_9735,N_9603);
nand U11618 (N_11618,N_9868,N_10215);
xnor U11619 (N_11619,N_9347,N_10390);
nand U11620 (N_11620,N_10114,N_9886);
or U11621 (N_11621,N_9930,N_10468);
and U11622 (N_11622,N_10465,N_9459);
or U11623 (N_11623,N_10035,N_9737);
nand U11624 (N_11624,N_9348,N_9709);
or U11625 (N_11625,N_9963,N_10108);
or U11626 (N_11626,N_9691,N_9306);
nand U11627 (N_11627,N_9705,N_10165);
nand U11628 (N_11628,N_9387,N_9650);
or U11629 (N_11629,N_10254,N_10066);
nor U11630 (N_11630,N_9305,N_9960);
or U11631 (N_11631,N_10036,N_9777);
xor U11632 (N_11632,N_9780,N_9350);
nor U11633 (N_11633,N_9565,N_9962);
nor U11634 (N_11634,N_9689,N_9241);
nor U11635 (N_11635,N_9928,N_9439);
nand U11636 (N_11636,N_10136,N_10499);
or U11637 (N_11637,N_9659,N_10083);
nand U11638 (N_11638,N_9531,N_10148);
xor U11639 (N_11639,N_9301,N_9117);
xnor U11640 (N_11640,N_10026,N_9911);
and U11641 (N_11641,N_9857,N_9626);
xnor U11642 (N_11642,N_10005,N_9811);
and U11643 (N_11643,N_10192,N_10412);
or U11644 (N_11644,N_10410,N_10250);
nand U11645 (N_11645,N_9283,N_9306);
and U11646 (N_11646,N_9663,N_9658);
nor U11647 (N_11647,N_9883,N_9743);
nand U11648 (N_11648,N_9157,N_10210);
or U11649 (N_11649,N_10260,N_9318);
and U11650 (N_11650,N_10338,N_9089);
nor U11651 (N_11651,N_10317,N_9599);
nor U11652 (N_11652,N_10109,N_10412);
or U11653 (N_11653,N_10427,N_9571);
nor U11654 (N_11654,N_10104,N_9106);
nand U11655 (N_11655,N_10140,N_10292);
nor U11656 (N_11656,N_9583,N_9272);
or U11657 (N_11657,N_9457,N_9689);
and U11658 (N_11658,N_10486,N_10103);
or U11659 (N_11659,N_10166,N_9818);
nor U11660 (N_11660,N_10355,N_10267);
and U11661 (N_11661,N_9169,N_9520);
nor U11662 (N_11662,N_10110,N_10229);
nor U11663 (N_11663,N_9637,N_9093);
and U11664 (N_11664,N_9225,N_9255);
or U11665 (N_11665,N_9149,N_10001);
nor U11666 (N_11666,N_9067,N_9665);
and U11667 (N_11667,N_9319,N_10145);
nor U11668 (N_11668,N_10314,N_9548);
and U11669 (N_11669,N_10061,N_10287);
nor U11670 (N_11670,N_10278,N_9779);
nor U11671 (N_11671,N_9164,N_9972);
or U11672 (N_11672,N_9576,N_9975);
and U11673 (N_11673,N_9060,N_10413);
nand U11674 (N_11674,N_9359,N_9541);
nor U11675 (N_11675,N_9096,N_9826);
or U11676 (N_11676,N_9207,N_9244);
or U11677 (N_11677,N_10139,N_10469);
nor U11678 (N_11678,N_9468,N_9643);
nand U11679 (N_11679,N_9939,N_9416);
and U11680 (N_11680,N_10477,N_9100);
or U11681 (N_11681,N_10463,N_9028);
nand U11682 (N_11682,N_9826,N_10161);
xor U11683 (N_11683,N_9127,N_9126);
xnor U11684 (N_11684,N_9169,N_9663);
and U11685 (N_11685,N_10129,N_9483);
and U11686 (N_11686,N_9881,N_9942);
nor U11687 (N_11687,N_9484,N_9666);
nor U11688 (N_11688,N_9275,N_9704);
nand U11689 (N_11689,N_10427,N_9122);
and U11690 (N_11690,N_9681,N_9789);
or U11691 (N_11691,N_9812,N_9909);
nand U11692 (N_11692,N_9887,N_9633);
xor U11693 (N_11693,N_9541,N_9272);
and U11694 (N_11694,N_9848,N_9162);
nor U11695 (N_11695,N_10231,N_9818);
or U11696 (N_11696,N_9306,N_9751);
or U11697 (N_11697,N_10169,N_10151);
nand U11698 (N_11698,N_10003,N_9433);
or U11699 (N_11699,N_9362,N_9188);
and U11700 (N_11700,N_9331,N_9562);
and U11701 (N_11701,N_9429,N_9897);
nor U11702 (N_11702,N_10471,N_9398);
nand U11703 (N_11703,N_9366,N_9470);
and U11704 (N_11704,N_9558,N_9994);
nor U11705 (N_11705,N_10468,N_9569);
and U11706 (N_11706,N_9598,N_10249);
or U11707 (N_11707,N_10321,N_10052);
and U11708 (N_11708,N_10082,N_10155);
and U11709 (N_11709,N_9304,N_9285);
nand U11710 (N_11710,N_9126,N_10384);
and U11711 (N_11711,N_9424,N_9251);
nor U11712 (N_11712,N_9212,N_9291);
nand U11713 (N_11713,N_9462,N_9269);
and U11714 (N_11714,N_9582,N_10353);
and U11715 (N_11715,N_9456,N_9785);
nor U11716 (N_11716,N_9668,N_9374);
nand U11717 (N_11717,N_10180,N_9602);
nand U11718 (N_11718,N_10331,N_9600);
nor U11719 (N_11719,N_10036,N_9917);
nand U11720 (N_11720,N_9907,N_9368);
nor U11721 (N_11721,N_9150,N_9333);
nand U11722 (N_11722,N_9631,N_9100);
and U11723 (N_11723,N_10386,N_9232);
nor U11724 (N_11724,N_10172,N_10051);
or U11725 (N_11725,N_10079,N_10496);
and U11726 (N_11726,N_9664,N_9955);
nor U11727 (N_11727,N_9843,N_9148);
and U11728 (N_11728,N_9723,N_9178);
or U11729 (N_11729,N_9266,N_9288);
nor U11730 (N_11730,N_9204,N_10487);
and U11731 (N_11731,N_9124,N_9293);
nor U11732 (N_11732,N_10392,N_9419);
nor U11733 (N_11733,N_9874,N_10209);
nand U11734 (N_11734,N_10175,N_10080);
or U11735 (N_11735,N_9241,N_10368);
and U11736 (N_11736,N_9763,N_9723);
nand U11737 (N_11737,N_10073,N_9682);
and U11738 (N_11738,N_9314,N_9662);
nor U11739 (N_11739,N_9107,N_9890);
nand U11740 (N_11740,N_10279,N_9754);
nand U11741 (N_11741,N_9754,N_9672);
nor U11742 (N_11742,N_10445,N_9870);
or U11743 (N_11743,N_9486,N_10204);
or U11744 (N_11744,N_10267,N_9570);
or U11745 (N_11745,N_9794,N_10035);
xnor U11746 (N_11746,N_9174,N_9536);
nor U11747 (N_11747,N_9718,N_9026);
nand U11748 (N_11748,N_10226,N_9090);
nand U11749 (N_11749,N_9641,N_9070);
and U11750 (N_11750,N_10250,N_9501);
and U11751 (N_11751,N_9091,N_9201);
nand U11752 (N_11752,N_10327,N_9938);
nor U11753 (N_11753,N_9870,N_10413);
nor U11754 (N_11754,N_10411,N_9004);
nand U11755 (N_11755,N_9763,N_9998);
nand U11756 (N_11756,N_9312,N_9056);
nand U11757 (N_11757,N_9037,N_9182);
or U11758 (N_11758,N_9055,N_10350);
nor U11759 (N_11759,N_10134,N_9273);
nand U11760 (N_11760,N_9889,N_9351);
nor U11761 (N_11761,N_10161,N_10049);
xnor U11762 (N_11762,N_9172,N_10039);
or U11763 (N_11763,N_10167,N_10190);
xor U11764 (N_11764,N_9796,N_10477);
xor U11765 (N_11765,N_9233,N_9529);
or U11766 (N_11766,N_10453,N_10092);
or U11767 (N_11767,N_9617,N_9997);
or U11768 (N_11768,N_10119,N_9990);
xnor U11769 (N_11769,N_10281,N_9938);
or U11770 (N_11770,N_9171,N_9890);
nand U11771 (N_11771,N_9687,N_9626);
nor U11772 (N_11772,N_9860,N_10192);
and U11773 (N_11773,N_10425,N_9591);
nor U11774 (N_11774,N_9649,N_9285);
nor U11775 (N_11775,N_9367,N_9454);
and U11776 (N_11776,N_9959,N_9257);
nor U11777 (N_11777,N_10175,N_10137);
and U11778 (N_11778,N_9603,N_9785);
xor U11779 (N_11779,N_9583,N_9762);
nand U11780 (N_11780,N_9102,N_9476);
or U11781 (N_11781,N_9485,N_9702);
and U11782 (N_11782,N_9207,N_10025);
nand U11783 (N_11783,N_9085,N_9256);
and U11784 (N_11784,N_9987,N_9330);
xor U11785 (N_11785,N_9355,N_10469);
nand U11786 (N_11786,N_9182,N_9660);
and U11787 (N_11787,N_9615,N_9302);
and U11788 (N_11788,N_10290,N_10072);
nand U11789 (N_11789,N_9807,N_9074);
nor U11790 (N_11790,N_9096,N_9762);
nand U11791 (N_11791,N_10303,N_9237);
xnor U11792 (N_11792,N_9431,N_9029);
or U11793 (N_11793,N_9329,N_9065);
xor U11794 (N_11794,N_10124,N_9837);
nand U11795 (N_11795,N_10172,N_9220);
nor U11796 (N_11796,N_9885,N_9056);
and U11797 (N_11797,N_9510,N_10052);
nand U11798 (N_11798,N_9903,N_10404);
and U11799 (N_11799,N_9348,N_9027);
and U11800 (N_11800,N_10117,N_10317);
or U11801 (N_11801,N_9720,N_9179);
and U11802 (N_11802,N_10048,N_10051);
nand U11803 (N_11803,N_10317,N_9059);
nor U11804 (N_11804,N_10449,N_10350);
and U11805 (N_11805,N_9417,N_9046);
xor U11806 (N_11806,N_9942,N_10454);
nand U11807 (N_11807,N_9845,N_10260);
nand U11808 (N_11808,N_9102,N_9654);
xor U11809 (N_11809,N_10182,N_9715);
nor U11810 (N_11810,N_10073,N_10207);
and U11811 (N_11811,N_10061,N_9371);
nand U11812 (N_11812,N_10241,N_9089);
and U11813 (N_11813,N_9872,N_9578);
and U11814 (N_11814,N_10023,N_10124);
or U11815 (N_11815,N_9776,N_10273);
and U11816 (N_11816,N_9460,N_10069);
or U11817 (N_11817,N_10272,N_10386);
nor U11818 (N_11818,N_9840,N_9929);
or U11819 (N_11819,N_10451,N_9594);
or U11820 (N_11820,N_9534,N_10215);
nand U11821 (N_11821,N_10310,N_9801);
nor U11822 (N_11822,N_10021,N_9537);
nor U11823 (N_11823,N_10002,N_9327);
or U11824 (N_11824,N_9521,N_9409);
and U11825 (N_11825,N_10484,N_10287);
or U11826 (N_11826,N_9390,N_9892);
or U11827 (N_11827,N_10444,N_9707);
or U11828 (N_11828,N_9146,N_9565);
or U11829 (N_11829,N_9384,N_9017);
and U11830 (N_11830,N_10296,N_10217);
and U11831 (N_11831,N_9049,N_9835);
nor U11832 (N_11832,N_10338,N_10387);
xor U11833 (N_11833,N_10234,N_9404);
or U11834 (N_11834,N_9933,N_9076);
or U11835 (N_11835,N_9434,N_9166);
nor U11836 (N_11836,N_10332,N_9921);
nand U11837 (N_11837,N_9545,N_9690);
or U11838 (N_11838,N_10444,N_9911);
nor U11839 (N_11839,N_9169,N_9292);
xnor U11840 (N_11840,N_9297,N_9161);
nor U11841 (N_11841,N_9183,N_10151);
nor U11842 (N_11842,N_10421,N_9626);
or U11843 (N_11843,N_10479,N_10071);
or U11844 (N_11844,N_10459,N_9197);
nand U11845 (N_11845,N_9469,N_10357);
and U11846 (N_11846,N_9823,N_9059);
and U11847 (N_11847,N_10490,N_9422);
nand U11848 (N_11848,N_9241,N_9870);
xnor U11849 (N_11849,N_9288,N_9237);
or U11850 (N_11850,N_10212,N_9602);
nand U11851 (N_11851,N_9647,N_10067);
nor U11852 (N_11852,N_9856,N_10335);
or U11853 (N_11853,N_9068,N_10471);
and U11854 (N_11854,N_10364,N_9734);
nand U11855 (N_11855,N_9022,N_10137);
nand U11856 (N_11856,N_9738,N_9106);
nor U11857 (N_11857,N_9232,N_9571);
nor U11858 (N_11858,N_9965,N_9353);
or U11859 (N_11859,N_9258,N_9978);
or U11860 (N_11860,N_10170,N_10140);
and U11861 (N_11861,N_10226,N_9331);
nor U11862 (N_11862,N_10096,N_9026);
nand U11863 (N_11863,N_9163,N_9004);
nor U11864 (N_11864,N_9011,N_9152);
nand U11865 (N_11865,N_9026,N_9204);
or U11866 (N_11866,N_10350,N_9122);
nor U11867 (N_11867,N_9842,N_9254);
nand U11868 (N_11868,N_9642,N_9295);
or U11869 (N_11869,N_9073,N_9436);
nor U11870 (N_11870,N_9800,N_9461);
and U11871 (N_11871,N_10163,N_10101);
nor U11872 (N_11872,N_9101,N_9537);
nor U11873 (N_11873,N_9620,N_10267);
or U11874 (N_11874,N_9831,N_9596);
nor U11875 (N_11875,N_10470,N_10229);
and U11876 (N_11876,N_10280,N_9521);
nand U11877 (N_11877,N_9908,N_10306);
or U11878 (N_11878,N_9051,N_9699);
nand U11879 (N_11879,N_9728,N_9721);
nand U11880 (N_11880,N_9017,N_9449);
nand U11881 (N_11881,N_9048,N_9418);
nor U11882 (N_11882,N_9613,N_9649);
nand U11883 (N_11883,N_9065,N_9493);
and U11884 (N_11884,N_9339,N_10146);
nand U11885 (N_11885,N_10164,N_9068);
or U11886 (N_11886,N_9336,N_10106);
and U11887 (N_11887,N_9327,N_10348);
nor U11888 (N_11888,N_9386,N_9213);
or U11889 (N_11889,N_9936,N_10137);
and U11890 (N_11890,N_10460,N_9181);
and U11891 (N_11891,N_9521,N_9767);
nor U11892 (N_11892,N_10267,N_9754);
and U11893 (N_11893,N_10339,N_10490);
or U11894 (N_11894,N_9943,N_9352);
and U11895 (N_11895,N_10316,N_9792);
and U11896 (N_11896,N_9185,N_9997);
and U11897 (N_11897,N_9567,N_9200);
nand U11898 (N_11898,N_10306,N_9237);
or U11899 (N_11899,N_9422,N_10351);
and U11900 (N_11900,N_10374,N_9482);
nand U11901 (N_11901,N_9189,N_9738);
or U11902 (N_11902,N_10243,N_9275);
or U11903 (N_11903,N_10312,N_9339);
nor U11904 (N_11904,N_9361,N_9346);
or U11905 (N_11905,N_10347,N_10346);
nand U11906 (N_11906,N_10137,N_9136);
or U11907 (N_11907,N_9461,N_9984);
or U11908 (N_11908,N_10052,N_9762);
or U11909 (N_11909,N_9881,N_10110);
xnor U11910 (N_11910,N_9477,N_9585);
xor U11911 (N_11911,N_9954,N_9635);
and U11912 (N_11912,N_10319,N_9200);
and U11913 (N_11913,N_9355,N_9723);
nor U11914 (N_11914,N_9457,N_9909);
nor U11915 (N_11915,N_9202,N_9586);
nand U11916 (N_11916,N_9205,N_9149);
nand U11917 (N_11917,N_9601,N_9943);
nor U11918 (N_11918,N_9202,N_9432);
and U11919 (N_11919,N_9616,N_9600);
nor U11920 (N_11920,N_10287,N_10037);
xnor U11921 (N_11921,N_9189,N_10188);
xor U11922 (N_11922,N_10316,N_10140);
nor U11923 (N_11923,N_9162,N_10011);
nand U11924 (N_11924,N_9583,N_10224);
and U11925 (N_11925,N_10008,N_10417);
nand U11926 (N_11926,N_10113,N_9383);
nor U11927 (N_11927,N_9123,N_10028);
xnor U11928 (N_11928,N_9338,N_10359);
nand U11929 (N_11929,N_10345,N_9247);
nand U11930 (N_11930,N_10163,N_9372);
or U11931 (N_11931,N_9921,N_9429);
xor U11932 (N_11932,N_9613,N_10331);
nor U11933 (N_11933,N_10332,N_9759);
nor U11934 (N_11934,N_10474,N_9128);
xnor U11935 (N_11935,N_9515,N_10108);
or U11936 (N_11936,N_9437,N_9546);
nor U11937 (N_11937,N_9966,N_10425);
and U11938 (N_11938,N_9678,N_9441);
nand U11939 (N_11939,N_9658,N_10133);
nor U11940 (N_11940,N_10109,N_9049);
or U11941 (N_11941,N_10098,N_9315);
and U11942 (N_11942,N_10220,N_9715);
nor U11943 (N_11943,N_10280,N_9160);
nand U11944 (N_11944,N_9214,N_9488);
and U11945 (N_11945,N_9343,N_9166);
nand U11946 (N_11946,N_9434,N_9395);
nand U11947 (N_11947,N_9695,N_9453);
nor U11948 (N_11948,N_10213,N_9926);
or U11949 (N_11949,N_9360,N_10026);
nand U11950 (N_11950,N_9440,N_9907);
xnor U11951 (N_11951,N_9476,N_9055);
nor U11952 (N_11952,N_9583,N_9874);
nor U11953 (N_11953,N_10291,N_9250);
nor U11954 (N_11954,N_9410,N_9039);
nand U11955 (N_11955,N_10435,N_9345);
or U11956 (N_11956,N_9561,N_9134);
nand U11957 (N_11957,N_10322,N_9864);
nand U11958 (N_11958,N_10008,N_10140);
and U11959 (N_11959,N_9989,N_9408);
and U11960 (N_11960,N_9599,N_9077);
and U11961 (N_11961,N_10050,N_9036);
and U11962 (N_11962,N_9795,N_10047);
nor U11963 (N_11963,N_9582,N_9901);
or U11964 (N_11964,N_10359,N_10463);
nor U11965 (N_11965,N_9084,N_9963);
and U11966 (N_11966,N_9500,N_9855);
or U11967 (N_11967,N_10003,N_9515);
nand U11968 (N_11968,N_10014,N_9374);
and U11969 (N_11969,N_9171,N_10373);
xnor U11970 (N_11970,N_10124,N_9754);
and U11971 (N_11971,N_10101,N_9310);
or U11972 (N_11972,N_10052,N_10216);
nand U11973 (N_11973,N_10408,N_9326);
nor U11974 (N_11974,N_9819,N_9565);
nand U11975 (N_11975,N_9453,N_9098);
nand U11976 (N_11976,N_9981,N_9502);
xnor U11977 (N_11977,N_10003,N_9937);
nand U11978 (N_11978,N_9712,N_9575);
and U11979 (N_11979,N_10012,N_9314);
or U11980 (N_11980,N_9138,N_10491);
nor U11981 (N_11981,N_9818,N_9208);
nand U11982 (N_11982,N_10090,N_10319);
nand U11983 (N_11983,N_10186,N_9405);
nand U11984 (N_11984,N_10133,N_9344);
nor U11985 (N_11985,N_9396,N_9761);
or U11986 (N_11986,N_10256,N_10372);
and U11987 (N_11987,N_9964,N_9284);
or U11988 (N_11988,N_9713,N_9474);
or U11989 (N_11989,N_9243,N_9879);
or U11990 (N_11990,N_9769,N_10076);
and U11991 (N_11991,N_9421,N_9777);
or U11992 (N_11992,N_9503,N_9895);
xnor U11993 (N_11993,N_10356,N_9011);
nor U11994 (N_11994,N_10267,N_9269);
and U11995 (N_11995,N_10187,N_9917);
and U11996 (N_11996,N_10394,N_9182);
and U11997 (N_11997,N_9932,N_9076);
nor U11998 (N_11998,N_9661,N_9859);
xor U11999 (N_11999,N_9202,N_10037);
and U12000 (N_12000,N_11084,N_11906);
nand U12001 (N_12001,N_11104,N_10596);
nand U12002 (N_12002,N_11551,N_11735);
and U12003 (N_12003,N_11020,N_11648);
or U12004 (N_12004,N_11847,N_10698);
nor U12005 (N_12005,N_10713,N_10819);
nor U12006 (N_12006,N_11943,N_11527);
xor U12007 (N_12007,N_10738,N_11662);
and U12008 (N_12008,N_11297,N_11508);
nand U12009 (N_12009,N_10830,N_11808);
or U12010 (N_12010,N_11058,N_11122);
nand U12011 (N_12011,N_11180,N_10924);
nor U12012 (N_12012,N_10918,N_10817);
and U12013 (N_12013,N_11251,N_11628);
or U12014 (N_12014,N_11330,N_11468);
and U12015 (N_12015,N_10616,N_11756);
or U12016 (N_12016,N_11718,N_11770);
and U12017 (N_12017,N_11797,N_10591);
or U12018 (N_12018,N_11607,N_11392);
or U12019 (N_12019,N_11445,N_10753);
or U12020 (N_12020,N_11779,N_11912);
or U12021 (N_12021,N_10896,N_10768);
or U12022 (N_12022,N_11731,N_11097);
nand U12023 (N_12023,N_11929,N_11518);
nand U12024 (N_12024,N_11126,N_11444);
or U12025 (N_12025,N_11114,N_10856);
nand U12026 (N_12026,N_11576,N_11064);
or U12027 (N_12027,N_11321,N_11855);
nor U12028 (N_12028,N_11841,N_11402);
and U12029 (N_12029,N_10609,N_11510);
or U12030 (N_12030,N_11582,N_11303);
nor U12031 (N_12031,N_11981,N_11646);
and U12032 (N_12032,N_10561,N_10673);
and U12033 (N_12033,N_11758,N_10938);
or U12034 (N_12034,N_11430,N_10672);
nand U12035 (N_12035,N_11208,N_10993);
xor U12036 (N_12036,N_11577,N_10663);
xor U12037 (N_12037,N_10560,N_11734);
and U12038 (N_12038,N_10878,N_11903);
or U12039 (N_12039,N_11026,N_11546);
or U12040 (N_12040,N_10539,N_11827);
or U12041 (N_12041,N_10893,N_10718);
or U12042 (N_12042,N_11106,N_11947);
and U12043 (N_12043,N_11443,N_11952);
nor U12044 (N_12044,N_11421,N_10628);
or U12045 (N_12045,N_11678,N_10955);
nor U12046 (N_12046,N_11203,N_11766);
nand U12047 (N_12047,N_11506,N_11273);
or U12048 (N_12048,N_10797,N_11983);
nand U12049 (N_12049,N_10970,N_10829);
nand U12050 (N_12050,N_10890,N_10631);
and U12051 (N_12051,N_11659,N_11773);
or U12052 (N_12052,N_11636,N_11156);
nand U12053 (N_12053,N_11075,N_10909);
and U12054 (N_12054,N_11959,N_11798);
nand U12055 (N_12055,N_11617,N_11562);
nand U12056 (N_12056,N_11516,N_11459);
or U12057 (N_12057,N_10534,N_11138);
and U12058 (N_12058,N_10528,N_11883);
or U12059 (N_12059,N_11334,N_11489);
nor U12060 (N_12060,N_11067,N_10593);
and U12061 (N_12061,N_11751,N_11343);
xor U12062 (N_12062,N_11086,N_11614);
xnor U12063 (N_12063,N_11812,N_11805);
or U12064 (N_12064,N_10719,N_11483);
or U12065 (N_12065,N_10971,N_11570);
nand U12066 (N_12066,N_11829,N_10919);
or U12067 (N_12067,N_10681,N_10660);
and U12068 (N_12068,N_11736,N_10553);
nor U12069 (N_12069,N_10604,N_11140);
xnor U12070 (N_12070,N_11656,N_11099);
and U12071 (N_12071,N_10676,N_11495);
nor U12072 (N_12072,N_10857,N_11365);
nand U12073 (N_12073,N_10769,N_10658);
and U12074 (N_12074,N_10712,N_11622);
nand U12075 (N_12075,N_11085,N_11214);
or U12076 (N_12076,N_11804,N_11428);
nor U12077 (N_12077,N_11749,N_10607);
xor U12078 (N_12078,N_11187,N_11644);
nor U12079 (N_12079,N_11984,N_11029);
nand U12080 (N_12080,N_11174,N_11599);
and U12081 (N_12081,N_11282,N_11536);
and U12082 (N_12082,N_11532,N_11728);
xnor U12083 (N_12083,N_10739,N_10541);
or U12084 (N_12084,N_10965,N_11715);
xor U12085 (N_12085,N_11839,N_11675);
nand U12086 (N_12086,N_10980,N_10781);
or U12087 (N_12087,N_11200,N_11862);
and U12088 (N_12088,N_10869,N_10899);
or U12089 (N_12089,N_11836,N_10888);
and U12090 (N_12090,N_11207,N_11463);
or U12091 (N_12091,N_11711,N_10633);
nand U12092 (N_12092,N_10551,N_10538);
nor U12093 (N_12093,N_11264,N_11046);
or U12094 (N_12094,N_11466,N_10599);
nand U12095 (N_12095,N_11295,N_11485);
nand U12096 (N_12096,N_11131,N_11250);
or U12097 (N_12097,N_10707,N_11567);
or U12098 (N_12098,N_10515,N_11332);
and U12099 (N_12099,N_11048,N_10642);
or U12100 (N_12100,N_11143,N_11574);
nand U12101 (N_12101,N_10925,N_11815);
or U12102 (N_12102,N_10763,N_10917);
xor U12103 (N_12103,N_10977,N_11842);
and U12104 (N_12104,N_10812,N_11647);
nand U12105 (N_12105,N_11367,N_11157);
or U12106 (N_12106,N_11217,N_11604);
xnor U12107 (N_12107,N_10537,N_11349);
nand U12108 (N_12108,N_11949,N_11145);
or U12109 (N_12109,N_11277,N_11061);
and U12110 (N_12110,N_10847,N_11924);
nand U12111 (N_12111,N_11922,N_11871);
nor U12112 (N_12112,N_11181,N_11720);
nand U12113 (N_12113,N_11997,N_11471);
and U12114 (N_12114,N_11920,N_10838);
or U12115 (N_12115,N_11291,N_10685);
nor U12116 (N_12116,N_10851,N_11882);
nor U12117 (N_12117,N_11164,N_11917);
or U12118 (N_12118,N_11951,N_11202);
and U12119 (N_12119,N_11125,N_11654);
nand U12120 (N_12120,N_11939,N_10505);
or U12121 (N_12121,N_11918,N_11930);
nor U12122 (N_12122,N_11670,N_11358);
and U12123 (N_12123,N_10986,N_11826);
and U12124 (N_12124,N_11389,N_10766);
nor U12125 (N_12125,N_10737,N_11155);
xor U12126 (N_12126,N_10532,N_10506);
or U12127 (N_12127,N_11394,N_10735);
nor U12128 (N_12128,N_10686,N_11750);
or U12129 (N_12129,N_11287,N_11860);
nor U12130 (N_12130,N_11645,N_11962);
and U12131 (N_12131,N_10746,N_11854);
or U12132 (N_12132,N_10948,N_10972);
or U12133 (N_12133,N_10854,N_11103);
xnor U12134 (N_12134,N_11945,N_10529);
nor U12135 (N_12135,N_11256,N_11995);
or U12136 (N_12136,N_11973,N_11848);
nand U12137 (N_12137,N_10708,N_10826);
or U12138 (N_12138,N_11176,N_11938);
nor U12139 (N_12139,N_10855,N_11120);
nor U12140 (N_12140,N_10790,N_11726);
and U12141 (N_12141,N_11727,N_11721);
nor U12142 (N_12142,N_10870,N_10689);
nand U12143 (N_12143,N_10680,N_10555);
and U12144 (N_12144,N_10873,N_11034);
nand U12145 (N_12145,N_11741,N_10876);
nand U12146 (N_12146,N_11305,N_10587);
nand U12147 (N_12147,N_10935,N_11783);
or U12148 (N_12148,N_10942,N_11616);
nand U12149 (N_12149,N_11115,N_11626);
and U12150 (N_12150,N_11960,N_10511);
and U12151 (N_12151,N_11159,N_11012);
nand U12152 (N_12152,N_11436,N_11141);
xnor U12153 (N_12153,N_11209,N_11892);
nor U12154 (N_12154,N_11618,N_11692);
xnor U12155 (N_12155,N_11565,N_10879);
xor U12156 (N_12156,N_10862,N_11889);
nand U12157 (N_12157,N_11254,N_11031);
and U12158 (N_12158,N_11969,N_11878);
nand U12159 (N_12159,N_11395,N_10783);
nor U12160 (N_12160,N_10792,N_11080);
and U12161 (N_12161,N_10531,N_11792);
or U12162 (N_12162,N_11698,N_10754);
or U12163 (N_12163,N_10775,N_11425);
xnor U12164 (N_12164,N_11496,N_10585);
nor U12165 (N_12165,N_11350,N_11825);
nand U12166 (N_12166,N_10974,N_11042);
nand U12167 (N_12167,N_10747,N_11213);
nand U12168 (N_12168,N_11447,N_11375);
nand U12169 (N_12169,N_11399,N_11397);
nand U12170 (N_12170,N_11769,N_11413);
or U12171 (N_12171,N_11151,N_10844);
nor U12172 (N_12172,N_11589,N_11033);
nor U12173 (N_12173,N_11894,N_10600);
or U12174 (N_12174,N_10800,N_11925);
or U12175 (N_12175,N_10833,N_10540);
or U12176 (N_12176,N_11002,N_11270);
or U12177 (N_12177,N_11239,N_10982);
nand U12178 (N_12178,N_11807,N_11417);
nand U12179 (N_12179,N_10772,N_10821);
nor U12180 (N_12180,N_11879,N_11348);
xor U12181 (N_12181,N_11594,N_11474);
nand U12182 (N_12182,N_10882,N_11457);
nor U12183 (N_12183,N_10729,N_11638);
nor U12184 (N_12184,N_11927,N_11975);
nand U12185 (N_12185,N_11245,N_10858);
and U12186 (N_12186,N_11666,N_11027);
and U12187 (N_12187,N_10589,N_11429);
and U12188 (N_12188,N_10552,N_11269);
and U12189 (N_12189,N_11197,N_11488);
nor U12190 (N_12190,N_10776,N_10877);
or U12191 (N_12191,N_11241,N_11028);
nor U12192 (N_12192,N_10656,N_11540);
nand U12193 (N_12193,N_11105,N_11979);
and U12194 (N_12194,N_10693,N_11230);
or U12195 (N_12195,N_11021,N_11653);
nor U12196 (N_12196,N_11405,N_11262);
xor U12197 (N_12197,N_10923,N_11011);
or U12198 (N_12198,N_11461,N_11416);
nand U12199 (N_12199,N_11781,N_11094);
nand U12200 (N_12200,N_10978,N_11049);
xnor U12201 (N_12201,N_10611,N_11407);
xor U12202 (N_12202,N_11761,N_11539);
nor U12203 (N_12203,N_11658,N_11811);
xor U12204 (N_12204,N_10894,N_11828);
or U12205 (N_12205,N_10533,N_11767);
nor U12206 (N_12206,N_11581,N_11246);
or U12207 (N_12207,N_10704,N_10949);
nor U12208 (N_12208,N_11861,N_11363);
and U12209 (N_12209,N_10931,N_10613);
nor U12210 (N_12210,N_11738,N_11052);
nor U12211 (N_12211,N_11832,N_11837);
or U12212 (N_12212,N_10786,N_11001);
and U12213 (N_12213,N_11458,N_11494);
nor U12214 (N_12214,N_11146,N_11921);
and U12215 (N_12215,N_11383,N_10927);
nand U12216 (N_12216,N_10548,N_11677);
or U12217 (N_12217,N_11036,N_10654);
nor U12218 (N_12218,N_11130,N_10582);
nor U12219 (N_12219,N_11830,N_11555);
nand U12220 (N_12220,N_11948,N_11802);
and U12221 (N_12221,N_10827,N_11346);
nand U12222 (N_12222,N_10644,N_11603);
nor U12223 (N_12223,N_11584,N_11127);
and U12224 (N_12224,N_10760,N_10535);
or U12225 (N_12225,N_10887,N_11624);
and U12226 (N_12226,N_11822,N_11440);
and U12227 (N_12227,N_10588,N_11703);
or U12228 (N_12228,N_10848,N_10525);
and U12229 (N_12229,N_10653,N_10788);
or U12230 (N_12230,N_11956,N_11077);
or U12231 (N_12231,N_11598,N_10751);
or U12232 (N_12232,N_10731,N_11742);
or U12233 (N_12233,N_11409,N_11763);
and U12234 (N_12234,N_10922,N_10715);
and U12235 (N_12235,N_10850,N_11554);
nor U12236 (N_12236,N_11932,N_11989);
nand U12237 (N_12237,N_11896,N_11649);
nor U12238 (N_12238,N_11091,N_11667);
and U12239 (N_12239,N_11869,N_10522);
nor U12240 (N_12240,N_11326,N_11700);
nand U12241 (N_12241,N_11403,N_11840);
and U12242 (N_12242,N_10814,N_10661);
nor U12243 (N_12243,N_11774,N_11037);
or U12244 (N_12244,N_11154,N_11136);
nand U12245 (N_12245,N_11509,N_10774);
nand U12246 (N_12246,N_11212,N_11994);
and U12247 (N_12247,N_10655,N_11331);
and U12248 (N_12248,N_11401,N_11743);
nor U12249 (N_12249,N_11147,N_11398);
xor U12250 (N_12250,N_11740,N_11550);
xor U12251 (N_12251,N_11188,N_11490);
nor U12252 (N_12252,N_11323,N_10597);
or U12253 (N_12253,N_11071,N_10668);
nor U12254 (N_12254,N_10976,N_11857);
or U12255 (N_12255,N_10626,N_10682);
and U12256 (N_12256,N_10697,N_11404);
or U12257 (N_12257,N_11017,N_11193);
or U12258 (N_12258,N_10710,N_11933);
xor U12259 (N_12259,N_11322,N_11548);
nand U12260 (N_12260,N_10943,N_11427);
xor U12261 (N_12261,N_11814,N_11886);
nand U12262 (N_12262,N_11557,N_10665);
and U12263 (N_12263,N_11846,N_11915);
nor U12264 (N_12264,N_10892,N_10615);
and U12265 (N_12265,N_10578,N_10900);
xnor U12266 (N_12266,N_11911,N_11679);
nor U12267 (N_12267,N_11530,N_11306);
or U12268 (N_12268,N_11759,N_10975);
nor U12269 (N_12269,N_11613,N_11177);
or U12270 (N_12270,N_11222,N_10958);
nand U12271 (N_12271,N_11010,N_11953);
and U12272 (N_12272,N_10543,N_11856);
and U12273 (N_12273,N_11190,N_11660);
nor U12274 (N_12274,N_10650,N_10988);
and U12275 (N_12275,N_11928,N_11507);
nor U12276 (N_12276,N_10520,N_11873);
and U12277 (N_12277,N_11923,N_10999);
nand U12278 (N_12278,N_11591,N_10610);
and U12279 (N_12279,N_11133,N_11313);
or U12280 (N_12280,N_11347,N_11118);
or U12281 (N_12281,N_11266,N_10632);
or U12282 (N_12282,N_10785,N_11746);
or U12283 (N_12283,N_10816,N_11359);
nand U12284 (N_12284,N_10939,N_11587);
nand U12285 (N_12285,N_10671,N_11556);
nor U12286 (N_12286,N_10575,N_11940);
xnor U12287 (N_12287,N_11867,N_11535);
nor U12288 (N_12288,N_11423,N_11681);
and U12289 (N_12289,N_11639,N_10886);
nand U12290 (N_12290,N_11179,N_11484);
xnor U12291 (N_12291,N_10957,N_11876);
and U12292 (N_12292,N_10973,N_11795);
and U12293 (N_12293,N_11253,N_11621);
nor U12294 (N_12294,N_11237,N_10780);
or U12295 (N_12295,N_10852,N_11976);
nand U12296 (N_12296,N_10761,N_10963);
or U12297 (N_12297,N_11820,N_11119);
nor U12298 (N_12298,N_11035,N_11885);
nor U12299 (N_12299,N_11312,N_10512);
or U12300 (N_12300,N_11941,N_11259);
nor U12301 (N_12301,N_11890,N_11631);
nand U12302 (N_12302,N_10572,N_10871);
nand U12303 (N_12303,N_11970,N_10777);
and U12304 (N_12304,N_10700,N_11559);
nor U12305 (N_12305,N_10523,N_11116);
nand U12306 (N_12306,N_11102,N_10806);
nand U12307 (N_12307,N_11977,N_11452);
or U12308 (N_12308,N_11833,N_11476);
and U12309 (N_12309,N_10726,N_11632);
and U12310 (N_12310,N_10524,N_10803);
nor U12311 (N_12311,N_11112,N_10728);
and U12312 (N_12312,N_11480,N_10885);
nor U12313 (N_12313,N_10645,N_11782);
or U12314 (N_12314,N_10962,N_10836);
nor U12315 (N_12315,N_11324,N_11041);
and U12316 (N_12316,N_11198,N_11370);
xnor U12317 (N_12317,N_11082,N_11004);
nor U12318 (N_12318,N_11893,N_11030);
xnor U12319 (N_12319,N_10714,N_11661);
or U12320 (N_12320,N_11818,N_11898);
and U12321 (N_12321,N_11884,N_11081);
nor U12322 (N_12322,N_11806,N_11547);
and U12323 (N_12323,N_11688,N_10567);
and U12324 (N_12324,N_11784,N_11369);
or U12325 (N_12325,N_11128,N_10779);
or U12326 (N_12326,N_11498,N_10581);
nor U12327 (N_12327,N_10592,N_11655);
xor U12328 (N_12328,N_11289,N_11134);
or U12329 (N_12329,N_11673,N_11709);
or U12330 (N_12330,N_11233,N_11218);
xnor U12331 (N_12331,N_11714,N_11148);
and U12332 (N_12332,N_11610,N_11088);
and U12333 (N_12333,N_11877,N_11754);
or U12334 (N_12334,N_10880,N_11637);
and U12335 (N_12335,N_10901,N_11946);
nor U12336 (N_12336,N_11400,N_11328);
or U12337 (N_12337,N_11796,N_10995);
nor U12338 (N_12338,N_10601,N_11513);
nand U12339 (N_12339,N_11694,N_11909);
nand U12340 (N_12340,N_11479,N_10799);
or U12341 (N_12341,N_10989,N_11185);
nor U12342 (N_12342,N_11462,N_11998);
nand U12343 (N_12343,N_11290,N_11844);
nand U12344 (N_12344,N_11695,N_11006);
and U12345 (N_12345,N_10967,N_10569);
xnor U12346 (N_12346,N_11705,N_11593);
xor U12347 (N_12347,N_10510,N_10595);
and U12348 (N_12348,N_10690,N_10767);
nor U12349 (N_12349,N_11016,N_11578);
and U12350 (N_12350,N_10677,N_11384);
and U12351 (N_12351,N_11776,N_11283);
and U12352 (N_12352,N_11907,N_10577);
and U12353 (N_12353,N_11542,N_10913);
nor U12354 (N_12354,N_11596,N_11755);
nand U12355 (N_12355,N_11451,N_11132);
nand U12356 (N_12356,N_10960,N_11340);
or U12357 (N_12357,N_11449,N_11139);
or U12358 (N_12358,N_11764,N_11719);
or U12359 (N_12359,N_11066,N_11153);
and U12360 (N_12360,N_10787,N_11315);
and U12361 (N_12361,N_10868,N_11378);
nor U12362 (N_12362,N_10641,N_10621);
nand U12363 (N_12363,N_11433,N_11005);
nor U12364 (N_12364,N_10742,N_11791);
nor U12365 (N_12365,N_11038,N_11453);
xnor U12366 (N_12366,N_10831,N_11117);
nand U12367 (N_12367,N_10921,N_10750);
and U12368 (N_12368,N_11364,N_11482);
and U12369 (N_12369,N_10692,N_11520);
nor U12370 (N_12370,N_10932,N_11481);
or U12371 (N_12371,N_11657,N_11595);
nor U12372 (N_12372,N_11210,N_11108);
and U12373 (N_12373,N_10985,N_11868);
nor U12374 (N_12374,N_11329,N_10934);
nand U12375 (N_12375,N_11696,N_11579);
and U12376 (N_12376,N_11170,N_11572);
nor U12377 (N_12377,N_11651,N_10562);
nor U12378 (N_12378,N_11563,N_11205);
and U12379 (N_12379,N_11963,N_11414);
xor U12380 (N_12380,N_11730,N_10674);
nand U12381 (N_12381,N_10782,N_11276);
nand U12382 (N_12382,N_11044,N_10657);
nand U12383 (N_12383,N_11630,N_11487);
nor U12384 (N_12384,N_11702,N_11519);
nand U12385 (N_12385,N_11689,N_11432);
or U12386 (N_12386,N_11265,N_11672);
and U12387 (N_12387,N_10765,N_10834);
nand U12388 (N_12388,N_11183,N_10634);
and U12389 (N_12389,N_11286,N_11913);
or U12390 (N_12390,N_11107,N_10846);
nand U12391 (N_12391,N_11142,N_11110);
xnor U12392 (N_12392,N_11990,N_11093);
nor U12393 (N_12393,N_11000,N_10670);
nor U12394 (N_12394,N_11062,N_10773);
and U12395 (N_12395,N_10623,N_10791);
nor U12396 (N_12396,N_10516,N_10701);
and U12397 (N_12397,N_11993,N_10903);
and U12398 (N_12398,N_11240,N_11271);
nand U12399 (N_12399,N_11019,N_10815);
nand U12400 (N_12400,N_11902,N_11493);
or U12401 (N_12401,N_11460,N_10636);
nor U12402 (N_12402,N_10648,N_10669);
nor U12403 (N_12403,N_10678,N_10998);
and U12404 (N_12404,N_10839,N_11184);
nor U12405 (N_12405,N_10579,N_11100);
nand U12406 (N_12406,N_11664,N_10796);
or U12407 (N_12407,N_11683,N_11411);
nand U12408 (N_12408,N_11712,N_10504);
or U12409 (N_12409,N_11919,N_10527);
and U12410 (N_12410,N_10916,N_11492);
nor U12411 (N_12411,N_10627,N_11353);
nor U12412 (N_12412,N_11611,N_11853);
and U12413 (N_12413,N_11745,N_11788);
nor U12414 (N_12414,N_10643,N_11319);
nor U12415 (N_12415,N_10564,N_10810);
nand U12416 (N_12416,N_11777,N_10614);
or U12417 (N_12417,N_10915,N_10884);
nor U12418 (N_12418,N_11261,N_11528);
and U12419 (N_12419,N_10947,N_10576);
nor U12420 (N_12420,N_11671,N_11704);
nor U12421 (N_12421,N_11327,N_11526);
and U12422 (N_12422,N_11454,N_11302);
and U12423 (N_12423,N_11691,N_10959);
or U12424 (N_12424,N_10625,N_11961);
or U12425 (N_12425,N_11355,N_11248);
nand U12426 (N_12426,N_10667,N_10566);
and U12427 (N_12427,N_10554,N_10649);
or U12428 (N_12428,N_11865,N_10752);
and U12429 (N_12429,N_11794,N_11014);
xnor U12430 (N_12430,N_11982,N_11499);
nand U12431 (N_12431,N_10991,N_10571);
xor U12432 (N_12432,N_11529,N_11229);
nor U12433 (N_12433,N_11580,N_11249);
or U12434 (N_12434,N_11824,N_11819);
nand U12435 (N_12435,N_11024,N_10602);
nand U12436 (N_12436,N_11101,N_11866);
and U12437 (N_12437,N_10969,N_11195);
and U12438 (N_12438,N_11583,N_11521);
nand U12439 (N_12439,N_11393,N_10984);
or U12440 (N_12440,N_11450,N_11022);
xor U12441 (N_12441,N_11235,N_11859);
and U12442 (N_12442,N_10651,N_11723);
or U12443 (N_12443,N_10549,N_10598);
and U12444 (N_12444,N_10687,N_10647);
nor U12445 (N_12445,N_11388,N_10867);
and U12446 (N_12446,N_10853,N_10759);
and U12447 (N_12447,N_11175,N_11419);
and U12448 (N_12448,N_11965,N_11412);
nand U12449 (N_12449,N_11040,N_11025);
nor U12450 (N_12450,N_10914,N_11051);
or U12451 (N_12451,N_10736,N_11008);
nand U12452 (N_12452,N_11722,N_11298);
nand U12453 (N_12453,N_10825,N_10946);
nand U12454 (N_12454,N_11944,N_10526);
xnor U12455 (N_12455,N_11601,N_11431);
xnor U12456 (N_12456,N_11371,N_11511);
nand U12457 (N_12457,N_11219,N_11768);
nand U12458 (N_12458,N_11335,N_10911);
and U12459 (N_12459,N_11469,N_10794);
xor U12460 (N_12460,N_10717,N_11368);
xor U12461 (N_12461,N_10733,N_11843);
or U12462 (N_12462,N_11434,N_11252);
nor U12463 (N_12463,N_10500,N_11267);
or U12464 (N_12464,N_11422,N_10705);
xor U12465 (N_12465,N_11352,N_11633);
or U12466 (N_12466,N_11744,N_11910);
nand U12467 (N_12467,N_11465,N_11070);
nand U12468 (N_12468,N_11189,N_11477);
nand U12469 (N_12469,N_11408,N_11166);
nor U12470 (N_12470,N_11294,N_11958);
nand U12471 (N_12471,N_11299,N_10703);
nand U12472 (N_12472,N_11699,N_11713);
nor U12473 (N_12473,N_11231,N_11096);
nor U12474 (N_12474,N_10513,N_11455);
nand U12475 (N_12475,N_11676,N_11800);
or U12476 (N_12476,N_11390,N_11162);
nand U12477 (N_12477,N_11293,N_11056);
and U12478 (N_12478,N_11361,N_11003);
or U12479 (N_12479,N_10546,N_10820);
nand U12480 (N_12480,N_11663,N_11227);
nand U12481 (N_12481,N_11609,N_10620);
and U12482 (N_12482,N_11602,N_11045);
nand U12483 (N_12483,N_11972,N_10688);
or U12484 (N_12484,N_11351,N_11475);
and U12485 (N_12485,N_11385,N_11525);
nor U12486 (N_12486,N_11426,N_10709);
and U12487 (N_12487,N_10987,N_11054);
nor U12488 (N_12488,N_11809,N_11872);
nand U12489 (N_12489,N_11284,N_11575);
and U12490 (N_12490,N_10864,N_11171);
and U12491 (N_12491,N_11888,N_11372);
and U12492 (N_12492,N_10920,N_11074);
nand U12493 (N_12493,N_11870,N_11491);
xor U12494 (N_12494,N_11957,N_11605);
nand U12495 (N_12495,N_10906,N_10740);
nor U12496 (N_12496,N_10996,N_11382);
and U12497 (N_12497,N_11223,N_10683);
nand U12498 (N_12498,N_11534,N_10699);
nor U12499 (N_12499,N_11308,N_11897);
nor U12500 (N_12500,N_11123,N_10994);
xnor U12501 (N_12501,N_11379,N_11092);
nand U12502 (N_12502,N_11354,N_11083);
nand U12503 (N_12503,N_11733,N_10568);
nand U12504 (N_12504,N_11242,N_10940);
nand U12505 (N_12505,N_11448,N_11473);
nand U12506 (N_12506,N_11762,N_10702);
or U12507 (N_12507,N_11339,N_10928);
nor U12508 (N_12508,N_10813,N_11533);
nor U12509 (N_12509,N_11737,N_11055);
and U12510 (N_12510,N_11338,N_11172);
and U12511 (N_12511,N_11059,N_11640);
and U12512 (N_12512,N_10638,N_11564);
nand U12513 (N_12513,N_10696,N_10635);
and U12514 (N_12514,N_11748,N_11517);
or U12515 (N_12515,N_11849,N_10675);
nand U12516 (N_12516,N_11620,N_11191);
nand U12517 (N_12517,N_10630,N_11281);
and U12518 (N_12518,N_11851,N_11739);
and U12519 (N_12519,N_11072,N_11864);
nand U12520 (N_12520,N_10694,N_11775);
nand U12521 (N_12521,N_11936,N_10666);
and U12522 (N_12522,N_11801,N_11161);
or U12523 (N_12523,N_10964,N_11914);
xnor U12524 (N_12524,N_11221,N_10908);
nor U12525 (N_12525,N_10695,N_10824);
nor U12526 (N_12526,N_11568,N_11901);
or U12527 (N_12527,N_11226,N_10849);
and U12528 (N_12528,N_11505,N_11124);
and U12529 (N_12529,N_11007,N_10983);
nand U12530 (N_12530,N_11199,N_11366);
nand U12531 (N_12531,N_10603,N_11747);
xor U12532 (N_12532,N_10547,N_10594);
xnor U12533 (N_12533,N_11701,N_10981);
nor U12534 (N_12534,N_11360,N_11435);
nor U12535 (N_12535,N_10646,N_11874);
or U12536 (N_12536,N_11627,N_10570);
and U12537 (N_12537,N_10872,N_11109);
or U12538 (N_12538,N_11320,N_11336);
and U12539 (N_12539,N_10556,N_10612);
or U12540 (N_12540,N_11987,N_11023);
nand U12541 (N_12541,N_11895,N_11971);
nand U12542 (N_12542,N_11725,N_11467);
nand U12543 (N_12543,N_10992,N_10748);
xor U12544 (N_12544,N_11357,N_11192);
nor U12545 (N_12545,N_11087,N_10590);
xnor U12546 (N_12546,N_11258,N_11968);
nor U12547 (N_12547,N_11247,N_11438);
nor U12548 (N_12548,N_11376,N_11486);
xor U12549 (N_12549,N_11377,N_11950);
nand U12550 (N_12550,N_11524,N_11803);
or U12551 (N_12551,N_11863,N_11665);
nor U12552 (N_12552,N_11150,N_11716);
and U12553 (N_12553,N_11032,N_11149);
nor U12554 (N_12554,N_11135,N_10881);
nand U12555 (N_12555,N_10756,N_10823);
xor U12556 (N_12556,N_11121,N_11515);
or U12557 (N_12557,N_11345,N_10637);
nor U12558 (N_12558,N_11641,N_11502);
nand U12559 (N_12559,N_11643,N_11999);
and U12560 (N_12560,N_11342,N_11985);
and U12561 (N_12561,N_10842,N_11439);
or U12562 (N_12562,N_11380,N_10762);
nand U12563 (N_12563,N_10802,N_11634);
nand U12564 (N_12564,N_10749,N_10811);
or U12565 (N_12565,N_10904,N_11437);
or U12566 (N_12566,N_11793,N_10798);
xor U12567 (N_12567,N_10837,N_10950);
and U12568 (N_12568,N_11296,N_11472);
and U12569 (N_12569,N_10745,N_11615);
and U12570 (N_12570,N_11787,N_11687);
nor U12571 (N_12571,N_11707,N_11904);
nor U12572 (N_12572,N_10514,N_11018);
nand U12573 (N_12573,N_11224,N_10954);
and U12574 (N_12574,N_11612,N_11680);
or U12575 (N_12575,N_11813,N_10720);
or U12576 (N_12576,N_11178,N_11571);
and U12577 (N_12577,N_10617,N_11668);
nand U12578 (N_12578,N_11980,N_11076);
nand U12579 (N_12579,N_10912,N_10933);
and U12580 (N_12580,N_11160,N_11586);
nand U12581 (N_12581,N_11053,N_11771);
nand U12582 (N_12582,N_10559,N_11344);
nand U12583 (N_12583,N_11942,N_10727);
nor U12584 (N_12584,N_11690,N_11850);
nand U12585 (N_12585,N_10652,N_10778);
and U12586 (N_12586,N_10805,N_11015);
xor U12587 (N_12587,N_11543,N_11597);
and U12588 (N_12588,N_10711,N_11799);
xor U12589 (N_12589,N_11710,N_11625);
or U12590 (N_12590,N_10544,N_11724);
nor U12591 (N_12591,N_10889,N_10679);
and U12592 (N_12592,N_10910,N_11558);
nand U12593 (N_12593,N_11560,N_11541);
or U12594 (N_12594,N_11307,N_11934);
nor U12595 (N_12595,N_11186,N_11585);
or U12596 (N_12596,N_11373,N_11243);
xor U12597 (N_12597,N_11978,N_11301);
nor U12598 (N_12598,N_11238,N_11279);
nand U12599 (N_12599,N_11514,N_11522);
nor U12600 (N_12600,N_10907,N_10684);
nor U12601 (N_12601,N_10563,N_11039);
or U12602 (N_12602,N_11232,N_11954);
or U12603 (N_12603,N_11729,N_10956);
nand U12604 (N_12604,N_10606,N_11167);
and U12605 (N_12605,N_11905,N_10517);
nand U12606 (N_12606,N_10664,N_11986);
nor U12607 (N_12607,N_10691,N_10507);
nor U12608 (N_12608,N_10659,N_11955);
nand U12609 (N_12609,N_11706,N_10770);
and U12610 (N_12610,N_10926,N_11234);
and U12611 (N_12611,N_11966,N_11047);
nand U12612 (N_12612,N_11089,N_11717);
or U12613 (N_12613,N_10584,N_11789);
nor U12614 (N_12614,N_10758,N_11441);
and U12615 (N_12615,N_10861,N_11988);
and U12616 (N_12616,N_10979,N_11916);
nor U12617 (N_12617,N_11635,N_11823);
or U12618 (N_12618,N_10809,N_10997);
nor U12619 (N_12619,N_10895,N_11470);
or U12620 (N_12620,N_11974,N_10502);
or U12621 (N_12621,N_10764,N_10706);
or U12622 (N_12622,N_11442,N_11310);
and U12623 (N_12623,N_11553,N_11194);
nor U12624 (N_12624,N_11215,N_10757);
or U12625 (N_12625,N_11504,N_11387);
and U12626 (N_12626,N_11606,N_10818);
nor U12627 (N_12627,N_10716,N_11549);
nand U12628 (N_12628,N_11079,N_11785);
or U12629 (N_12629,N_11908,N_11073);
nor U12630 (N_12630,N_11216,N_11835);
xnor U12631 (N_12631,N_11497,N_11069);
and U12632 (N_12632,N_11652,N_11552);
nor U12633 (N_12633,N_11420,N_11317);
nor U12634 (N_12634,N_11292,N_10521);
or U12635 (N_12635,N_11569,N_10944);
nand U12636 (N_12636,N_10840,N_11418);
nor U12637 (N_12637,N_11790,N_11778);
nand U12638 (N_12638,N_11693,N_11752);
xnor U12639 (N_12639,N_11236,N_11182);
nor U12640 (N_12640,N_11501,N_11674);
nor U12641 (N_12641,N_10509,N_11137);
or U12642 (N_12642,N_10966,N_11887);
xnor U12643 (N_12643,N_10898,N_11891);
or U12644 (N_12644,N_10542,N_11845);
and U12645 (N_12645,N_10859,N_10937);
nor U12646 (N_12646,N_11900,N_11244);
and U12647 (N_12647,N_11446,N_10550);
nor U12648 (N_12648,N_11415,N_10929);
nor U12649 (N_12649,N_11255,N_11288);
nor U12650 (N_12650,N_11196,N_11685);
or U12651 (N_12651,N_10518,N_11057);
and U12652 (N_12652,N_10624,N_10744);
and U12653 (N_12653,N_11545,N_10734);
and U12654 (N_12654,N_10945,N_10503);
and U12655 (N_12655,N_11228,N_11318);
or U12656 (N_12656,N_11852,N_11588);
or U12657 (N_12657,N_11753,N_11899);
and U12658 (N_12658,N_10743,N_11478);
xor U12659 (N_12659,N_10557,N_10835);
and U12660 (N_12660,N_11537,N_11013);
nand U12661 (N_12661,N_10902,N_11406);
xnor U12662 (N_12662,N_10725,N_10860);
or U12663 (N_12663,N_11926,N_11992);
and U12664 (N_12664,N_10619,N_11316);
nand U12665 (N_12665,N_11078,N_11732);
and U12666 (N_12666,N_10640,N_11561);
nand U12667 (N_12667,N_11165,N_11931);
xnor U12668 (N_12668,N_11263,N_10722);
or U12669 (N_12669,N_11817,N_11362);
and U12670 (N_12670,N_11111,N_10583);
nor U12671 (N_12671,N_11875,N_11391);
and U12672 (N_12672,N_11386,N_11211);
nor U12673 (N_12673,N_11260,N_11765);
nor U12674 (N_12674,N_11341,N_10565);
or U12675 (N_12675,N_11374,N_10573);
xor U12676 (N_12676,N_11274,N_11996);
or U12677 (N_12677,N_10501,N_11566);
and U12678 (N_12678,N_10808,N_11821);
nand U12679 (N_12679,N_10639,N_10897);
nor U12680 (N_12680,N_11285,N_11600);
nand U12681 (N_12681,N_11337,N_11275);
or U12682 (N_12682,N_11512,N_11573);
nor U12683 (N_12683,N_11642,N_11098);
nor U12684 (N_12684,N_11786,N_10530);
nor U12685 (N_12685,N_11168,N_10941);
nand U12686 (N_12686,N_10723,N_10605);
nand U12687 (N_12687,N_10545,N_10863);
and U12688 (N_12688,N_10832,N_11592);
nand U12689 (N_12689,N_11590,N_11206);
or U12690 (N_12690,N_10558,N_11619);
and U12691 (N_12691,N_11881,N_11424);
and U12692 (N_12692,N_10662,N_10771);
or U12693 (N_12693,N_11757,N_10807);
nand U12694 (N_12694,N_11043,N_10586);
xnor U12695 (N_12695,N_10508,N_11531);
and U12696 (N_12696,N_10891,N_11257);
nor U12697 (N_12697,N_11204,N_10804);
nand U12698 (N_12698,N_10724,N_10828);
or U12699 (N_12699,N_10519,N_11009);
or U12700 (N_12700,N_11629,N_11225);
xor U12701 (N_12701,N_10574,N_11544);
nand U12702 (N_12702,N_10930,N_10793);
or U12703 (N_12703,N_11060,N_11816);
nand U12704 (N_12704,N_11456,N_10822);
nor U12705 (N_12705,N_11523,N_10953);
and U12706 (N_12706,N_10874,N_11158);
or U12707 (N_12707,N_11113,N_11500);
nor U12708 (N_12708,N_11858,N_11090);
or U12709 (N_12709,N_10961,N_11538);
nor U12710 (N_12710,N_11991,N_10618);
or U12711 (N_12711,N_11356,N_10875);
and U12712 (N_12712,N_11937,N_10841);
nor U12713 (N_12713,N_11964,N_10721);
nor U12714 (N_12714,N_11669,N_11068);
xnor U12715 (N_12715,N_11831,N_11144);
nor U12716 (N_12716,N_11268,N_10801);
or U12717 (N_12717,N_10730,N_11410);
and U12718 (N_12718,N_10905,N_11201);
or U12719 (N_12719,N_11300,N_11935);
xnor U12720 (N_12720,N_10755,N_11772);
nand U12721 (N_12721,N_10580,N_11129);
nand U12722 (N_12722,N_10865,N_11708);
xor U12723 (N_12723,N_11967,N_10990);
nor U12724 (N_12724,N_10608,N_11152);
nor U12725 (N_12725,N_11311,N_11220);
nand U12726 (N_12726,N_10732,N_11063);
or U12727 (N_12727,N_11304,N_11464);
nand U12728 (N_12728,N_11834,N_11333);
nor U12729 (N_12729,N_10936,N_11272);
nand U12730 (N_12730,N_10866,N_10536);
nor U12731 (N_12731,N_11280,N_11381);
nor U12732 (N_12732,N_11278,N_11623);
xor U12733 (N_12733,N_11163,N_11686);
nor U12734 (N_12734,N_11697,N_10883);
xnor U12735 (N_12735,N_11050,N_11760);
or U12736 (N_12736,N_10843,N_11608);
nand U12737 (N_12737,N_11682,N_10951);
xnor U12738 (N_12738,N_10741,N_11684);
nor U12739 (N_12739,N_11309,N_11780);
or U12740 (N_12740,N_11880,N_11314);
and U12741 (N_12741,N_11095,N_11325);
nor U12742 (N_12742,N_10795,N_10629);
or U12743 (N_12743,N_11169,N_11838);
or U12744 (N_12744,N_11650,N_11810);
nor U12745 (N_12745,N_10789,N_10622);
xnor U12746 (N_12746,N_10784,N_11065);
and U12747 (N_12747,N_10845,N_11396);
nand U12748 (N_12748,N_10968,N_10952);
and U12749 (N_12749,N_11173,N_11503);
nor U12750 (N_12750,N_10539,N_11407);
or U12751 (N_12751,N_10692,N_10586);
xnor U12752 (N_12752,N_10662,N_10862);
nor U12753 (N_12753,N_11375,N_11859);
nand U12754 (N_12754,N_11919,N_11291);
and U12755 (N_12755,N_11015,N_10848);
xnor U12756 (N_12756,N_11902,N_11720);
nand U12757 (N_12757,N_11434,N_11066);
nand U12758 (N_12758,N_10663,N_10706);
or U12759 (N_12759,N_10953,N_11591);
and U12760 (N_12760,N_11192,N_11218);
nand U12761 (N_12761,N_11100,N_10584);
or U12762 (N_12762,N_11607,N_11328);
nand U12763 (N_12763,N_11325,N_11747);
nor U12764 (N_12764,N_10871,N_11258);
nand U12765 (N_12765,N_11530,N_10903);
or U12766 (N_12766,N_10585,N_11406);
or U12767 (N_12767,N_11342,N_10960);
nor U12768 (N_12768,N_10648,N_11382);
or U12769 (N_12769,N_10665,N_11479);
or U12770 (N_12770,N_11983,N_11751);
nand U12771 (N_12771,N_11264,N_11030);
nor U12772 (N_12772,N_10916,N_11798);
or U12773 (N_12773,N_10642,N_11917);
or U12774 (N_12774,N_11669,N_10648);
nor U12775 (N_12775,N_11587,N_11970);
nand U12776 (N_12776,N_11578,N_11118);
or U12777 (N_12777,N_10781,N_10574);
nor U12778 (N_12778,N_11840,N_11499);
and U12779 (N_12779,N_11612,N_10979);
nor U12780 (N_12780,N_11803,N_10534);
and U12781 (N_12781,N_10566,N_11976);
nor U12782 (N_12782,N_11881,N_11125);
or U12783 (N_12783,N_11367,N_11529);
xnor U12784 (N_12784,N_11309,N_10710);
and U12785 (N_12785,N_11442,N_10920);
or U12786 (N_12786,N_10870,N_11478);
xor U12787 (N_12787,N_10755,N_11281);
or U12788 (N_12788,N_10826,N_11396);
and U12789 (N_12789,N_11616,N_11095);
or U12790 (N_12790,N_11871,N_11254);
and U12791 (N_12791,N_10551,N_11285);
or U12792 (N_12792,N_10886,N_10987);
or U12793 (N_12793,N_11638,N_11634);
nor U12794 (N_12794,N_10655,N_10962);
or U12795 (N_12795,N_10658,N_11491);
nand U12796 (N_12796,N_11714,N_10573);
nor U12797 (N_12797,N_10700,N_11986);
nand U12798 (N_12798,N_11119,N_11811);
nor U12799 (N_12799,N_11603,N_11103);
nor U12800 (N_12800,N_11481,N_10568);
nand U12801 (N_12801,N_11873,N_10553);
and U12802 (N_12802,N_11316,N_11443);
nor U12803 (N_12803,N_11989,N_10806);
nor U12804 (N_12804,N_10744,N_11384);
or U12805 (N_12805,N_10696,N_11584);
nand U12806 (N_12806,N_11472,N_10933);
or U12807 (N_12807,N_11152,N_11434);
nor U12808 (N_12808,N_10679,N_11363);
and U12809 (N_12809,N_11439,N_11477);
or U12810 (N_12810,N_11862,N_11682);
or U12811 (N_12811,N_11851,N_10822);
or U12812 (N_12812,N_11204,N_11645);
nand U12813 (N_12813,N_10665,N_10622);
nand U12814 (N_12814,N_11339,N_11068);
and U12815 (N_12815,N_11775,N_11028);
nand U12816 (N_12816,N_10881,N_11699);
and U12817 (N_12817,N_11202,N_11726);
nor U12818 (N_12818,N_10692,N_11293);
nand U12819 (N_12819,N_10882,N_11045);
or U12820 (N_12820,N_11147,N_10544);
and U12821 (N_12821,N_11079,N_11553);
and U12822 (N_12822,N_11914,N_11242);
nor U12823 (N_12823,N_11584,N_10632);
and U12824 (N_12824,N_11129,N_10750);
and U12825 (N_12825,N_11351,N_10560);
xnor U12826 (N_12826,N_10541,N_11153);
nand U12827 (N_12827,N_11790,N_11823);
or U12828 (N_12828,N_11599,N_11200);
xnor U12829 (N_12829,N_11668,N_10577);
or U12830 (N_12830,N_11766,N_10759);
xor U12831 (N_12831,N_11681,N_11052);
and U12832 (N_12832,N_10888,N_10589);
nand U12833 (N_12833,N_11829,N_10697);
or U12834 (N_12834,N_10530,N_11111);
nand U12835 (N_12835,N_11467,N_11980);
xnor U12836 (N_12836,N_10793,N_11022);
xor U12837 (N_12837,N_11036,N_11122);
xnor U12838 (N_12838,N_11452,N_10865);
or U12839 (N_12839,N_10655,N_10584);
nor U12840 (N_12840,N_10753,N_10502);
or U12841 (N_12841,N_11933,N_11418);
nor U12842 (N_12842,N_11869,N_11613);
nand U12843 (N_12843,N_11702,N_10897);
nand U12844 (N_12844,N_11115,N_11049);
and U12845 (N_12845,N_11934,N_10911);
or U12846 (N_12846,N_11841,N_11346);
or U12847 (N_12847,N_11348,N_11150);
or U12848 (N_12848,N_10877,N_11167);
nor U12849 (N_12849,N_11319,N_11129);
and U12850 (N_12850,N_11822,N_10558);
nand U12851 (N_12851,N_10843,N_11692);
nand U12852 (N_12852,N_10639,N_10772);
nand U12853 (N_12853,N_11597,N_10773);
and U12854 (N_12854,N_10941,N_10739);
or U12855 (N_12855,N_10740,N_11996);
and U12856 (N_12856,N_11280,N_11560);
nand U12857 (N_12857,N_11706,N_10608);
or U12858 (N_12858,N_11303,N_10981);
nor U12859 (N_12859,N_11727,N_11329);
nor U12860 (N_12860,N_11667,N_11712);
nand U12861 (N_12861,N_10577,N_11243);
xor U12862 (N_12862,N_11247,N_11889);
xor U12863 (N_12863,N_10694,N_11116);
and U12864 (N_12864,N_11894,N_11364);
or U12865 (N_12865,N_11801,N_11504);
and U12866 (N_12866,N_11943,N_11126);
or U12867 (N_12867,N_10651,N_10595);
and U12868 (N_12868,N_10621,N_11749);
nor U12869 (N_12869,N_10572,N_11181);
xor U12870 (N_12870,N_11952,N_11789);
nor U12871 (N_12871,N_10538,N_11321);
nor U12872 (N_12872,N_10984,N_10872);
or U12873 (N_12873,N_10948,N_10613);
nand U12874 (N_12874,N_11954,N_11744);
or U12875 (N_12875,N_11450,N_11162);
nor U12876 (N_12876,N_11742,N_11204);
xnor U12877 (N_12877,N_11519,N_11034);
nand U12878 (N_12878,N_11683,N_10858);
nor U12879 (N_12879,N_11132,N_10828);
xnor U12880 (N_12880,N_11321,N_11100);
or U12881 (N_12881,N_11333,N_10690);
and U12882 (N_12882,N_11777,N_10721);
nor U12883 (N_12883,N_10685,N_11319);
and U12884 (N_12884,N_10628,N_11902);
or U12885 (N_12885,N_11551,N_11619);
or U12886 (N_12886,N_11982,N_11219);
or U12887 (N_12887,N_11242,N_11588);
or U12888 (N_12888,N_11557,N_11642);
nand U12889 (N_12889,N_10851,N_11503);
nor U12890 (N_12890,N_11925,N_11323);
nand U12891 (N_12891,N_11036,N_11498);
xnor U12892 (N_12892,N_11279,N_11171);
xnor U12893 (N_12893,N_10675,N_11015);
nor U12894 (N_12894,N_10691,N_11780);
nor U12895 (N_12895,N_10892,N_11791);
nor U12896 (N_12896,N_11527,N_10660);
and U12897 (N_12897,N_10737,N_11747);
nor U12898 (N_12898,N_11687,N_10711);
and U12899 (N_12899,N_10832,N_10566);
or U12900 (N_12900,N_11978,N_11687);
or U12901 (N_12901,N_11169,N_11992);
or U12902 (N_12902,N_11765,N_11067);
or U12903 (N_12903,N_11355,N_11432);
nand U12904 (N_12904,N_11851,N_11649);
or U12905 (N_12905,N_11106,N_10993);
xor U12906 (N_12906,N_10756,N_11605);
nor U12907 (N_12907,N_10955,N_11292);
nor U12908 (N_12908,N_10756,N_10900);
nand U12909 (N_12909,N_11350,N_11345);
nor U12910 (N_12910,N_11453,N_11224);
and U12911 (N_12911,N_11362,N_10595);
nand U12912 (N_12912,N_11819,N_10800);
nand U12913 (N_12913,N_11071,N_11259);
or U12914 (N_12914,N_11405,N_11348);
xnor U12915 (N_12915,N_10808,N_10889);
nor U12916 (N_12916,N_11796,N_11148);
or U12917 (N_12917,N_11595,N_10945);
xnor U12918 (N_12918,N_11710,N_11276);
nor U12919 (N_12919,N_10579,N_11787);
or U12920 (N_12920,N_11652,N_11673);
nor U12921 (N_12921,N_11793,N_10595);
or U12922 (N_12922,N_11688,N_10935);
or U12923 (N_12923,N_11621,N_10780);
and U12924 (N_12924,N_11685,N_11711);
and U12925 (N_12925,N_11957,N_11207);
and U12926 (N_12926,N_11596,N_10846);
nor U12927 (N_12927,N_10845,N_11290);
nand U12928 (N_12928,N_11130,N_10940);
nand U12929 (N_12929,N_11237,N_11947);
or U12930 (N_12930,N_11635,N_11498);
or U12931 (N_12931,N_10970,N_11933);
nor U12932 (N_12932,N_10639,N_11734);
nor U12933 (N_12933,N_11992,N_11751);
nor U12934 (N_12934,N_11083,N_11782);
nand U12935 (N_12935,N_11200,N_11561);
nand U12936 (N_12936,N_11541,N_10573);
and U12937 (N_12937,N_11094,N_11024);
or U12938 (N_12938,N_11277,N_11180);
nor U12939 (N_12939,N_10715,N_11437);
nand U12940 (N_12940,N_11135,N_11065);
nor U12941 (N_12941,N_11479,N_11388);
or U12942 (N_12942,N_11622,N_11836);
nor U12943 (N_12943,N_10501,N_11320);
nand U12944 (N_12944,N_11562,N_10557);
nand U12945 (N_12945,N_11352,N_11429);
or U12946 (N_12946,N_10547,N_11939);
xnor U12947 (N_12947,N_11709,N_11501);
and U12948 (N_12948,N_11208,N_11051);
nor U12949 (N_12949,N_11021,N_10637);
nor U12950 (N_12950,N_11549,N_10634);
and U12951 (N_12951,N_10963,N_11281);
or U12952 (N_12952,N_11491,N_11215);
nand U12953 (N_12953,N_11170,N_11364);
or U12954 (N_12954,N_11232,N_10646);
xor U12955 (N_12955,N_10897,N_11106);
nand U12956 (N_12956,N_11924,N_11727);
nand U12957 (N_12957,N_11274,N_11886);
nand U12958 (N_12958,N_11795,N_11417);
or U12959 (N_12959,N_10616,N_10874);
nor U12960 (N_12960,N_11499,N_10973);
xnor U12961 (N_12961,N_11103,N_10894);
nor U12962 (N_12962,N_10549,N_11784);
or U12963 (N_12963,N_11003,N_11479);
nor U12964 (N_12964,N_10790,N_10956);
xnor U12965 (N_12965,N_11976,N_10741);
and U12966 (N_12966,N_11724,N_10632);
nand U12967 (N_12967,N_11572,N_11515);
xnor U12968 (N_12968,N_11535,N_10998);
and U12969 (N_12969,N_11018,N_11398);
and U12970 (N_12970,N_11175,N_11560);
and U12971 (N_12971,N_11353,N_10637);
or U12972 (N_12972,N_11746,N_11877);
and U12973 (N_12973,N_11582,N_10507);
nand U12974 (N_12974,N_11929,N_10761);
xnor U12975 (N_12975,N_11680,N_10710);
nor U12976 (N_12976,N_11967,N_10767);
nand U12977 (N_12977,N_10902,N_11906);
nand U12978 (N_12978,N_11813,N_11312);
nor U12979 (N_12979,N_11422,N_11138);
xor U12980 (N_12980,N_10737,N_11129);
nand U12981 (N_12981,N_11681,N_11682);
and U12982 (N_12982,N_10956,N_11299);
nor U12983 (N_12983,N_10748,N_11235);
nand U12984 (N_12984,N_11621,N_11247);
nor U12985 (N_12985,N_11505,N_10846);
and U12986 (N_12986,N_10557,N_11211);
nor U12987 (N_12987,N_10610,N_11614);
nand U12988 (N_12988,N_11899,N_11440);
and U12989 (N_12989,N_11764,N_11435);
and U12990 (N_12990,N_11746,N_11658);
or U12991 (N_12991,N_11274,N_11823);
or U12992 (N_12992,N_10679,N_11836);
nor U12993 (N_12993,N_11134,N_11584);
nor U12994 (N_12994,N_10924,N_10540);
and U12995 (N_12995,N_11879,N_11900);
or U12996 (N_12996,N_11918,N_11854);
xor U12997 (N_12997,N_10757,N_11709);
and U12998 (N_12998,N_10541,N_11368);
or U12999 (N_12999,N_10646,N_11205);
nor U13000 (N_13000,N_11507,N_11386);
or U13001 (N_13001,N_10944,N_11079);
nor U13002 (N_13002,N_11581,N_10932);
nor U13003 (N_13003,N_10914,N_10858);
or U13004 (N_13004,N_11912,N_11879);
or U13005 (N_13005,N_11440,N_11413);
or U13006 (N_13006,N_11490,N_11057);
nand U13007 (N_13007,N_11328,N_11839);
or U13008 (N_13008,N_11128,N_11710);
or U13009 (N_13009,N_11366,N_10962);
xnor U13010 (N_13010,N_11941,N_11356);
and U13011 (N_13011,N_11577,N_11146);
or U13012 (N_13012,N_11237,N_11444);
nor U13013 (N_13013,N_11328,N_11198);
or U13014 (N_13014,N_11720,N_10616);
and U13015 (N_13015,N_11043,N_10792);
nor U13016 (N_13016,N_10794,N_11492);
nand U13017 (N_13017,N_11011,N_11487);
and U13018 (N_13018,N_11329,N_11150);
nor U13019 (N_13019,N_11092,N_11457);
nand U13020 (N_13020,N_11105,N_11582);
nor U13021 (N_13021,N_11108,N_11705);
and U13022 (N_13022,N_10547,N_11253);
xor U13023 (N_13023,N_10748,N_10758);
and U13024 (N_13024,N_10904,N_11124);
nand U13025 (N_13025,N_11332,N_11352);
nor U13026 (N_13026,N_10700,N_11226);
and U13027 (N_13027,N_10580,N_11172);
and U13028 (N_13028,N_11998,N_11548);
nor U13029 (N_13029,N_10726,N_11850);
and U13030 (N_13030,N_11452,N_11605);
nor U13031 (N_13031,N_10822,N_11167);
nand U13032 (N_13032,N_10891,N_10690);
and U13033 (N_13033,N_10661,N_11237);
nor U13034 (N_13034,N_11091,N_10716);
nor U13035 (N_13035,N_10515,N_10850);
nor U13036 (N_13036,N_11745,N_11879);
nand U13037 (N_13037,N_10993,N_10567);
and U13038 (N_13038,N_11530,N_11455);
or U13039 (N_13039,N_11758,N_11771);
and U13040 (N_13040,N_11781,N_11153);
or U13041 (N_13041,N_10664,N_11638);
nor U13042 (N_13042,N_11634,N_11695);
or U13043 (N_13043,N_11842,N_11218);
nor U13044 (N_13044,N_11268,N_11044);
or U13045 (N_13045,N_11574,N_10905);
nor U13046 (N_13046,N_10517,N_11953);
nor U13047 (N_13047,N_10805,N_11660);
or U13048 (N_13048,N_10676,N_11427);
nand U13049 (N_13049,N_11930,N_11255);
nor U13050 (N_13050,N_11958,N_11477);
nor U13051 (N_13051,N_11165,N_11549);
nand U13052 (N_13052,N_11875,N_10978);
or U13053 (N_13053,N_11291,N_10555);
xnor U13054 (N_13054,N_11314,N_10898);
nand U13055 (N_13055,N_11432,N_11034);
xnor U13056 (N_13056,N_11629,N_11149);
or U13057 (N_13057,N_11865,N_11473);
nand U13058 (N_13058,N_11257,N_10943);
or U13059 (N_13059,N_10877,N_10547);
and U13060 (N_13060,N_11555,N_11514);
nand U13061 (N_13061,N_11035,N_10585);
nand U13062 (N_13062,N_11059,N_11172);
nand U13063 (N_13063,N_11841,N_10703);
or U13064 (N_13064,N_11189,N_11133);
and U13065 (N_13065,N_11528,N_11510);
or U13066 (N_13066,N_11931,N_11959);
or U13067 (N_13067,N_10823,N_10717);
nor U13068 (N_13068,N_10847,N_10564);
nor U13069 (N_13069,N_11709,N_11395);
nand U13070 (N_13070,N_11698,N_11666);
nor U13071 (N_13071,N_10919,N_11674);
nand U13072 (N_13072,N_10615,N_11150);
nor U13073 (N_13073,N_11063,N_11862);
or U13074 (N_13074,N_11425,N_11960);
nand U13075 (N_13075,N_10958,N_10956);
nor U13076 (N_13076,N_10822,N_11829);
and U13077 (N_13077,N_11253,N_11507);
nand U13078 (N_13078,N_11034,N_10648);
and U13079 (N_13079,N_11830,N_11793);
or U13080 (N_13080,N_11883,N_11471);
or U13081 (N_13081,N_10506,N_10765);
or U13082 (N_13082,N_10920,N_10899);
xor U13083 (N_13083,N_10501,N_11592);
and U13084 (N_13084,N_10707,N_11276);
nand U13085 (N_13085,N_10690,N_11946);
nor U13086 (N_13086,N_11448,N_10721);
xor U13087 (N_13087,N_10987,N_10915);
nand U13088 (N_13088,N_10726,N_10636);
nand U13089 (N_13089,N_11114,N_11725);
nor U13090 (N_13090,N_11521,N_10869);
and U13091 (N_13091,N_10634,N_10687);
or U13092 (N_13092,N_10664,N_11212);
and U13093 (N_13093,N_11319,N_11193);
and U13094 (N_13094,N_11073,N_11529);
nor U13095 (N_13095,N_11872,N_11869);
or U13096 (N_13096,N_11239,N_11580);
nor U13097 (N_13097,N_11464,N_10506);
or U13098 (N_13098,N_11662,N_11554);
nor U13099 (N_13099,N_10532,N_11759);
xor U13100 (N_13100,N_11212,N_11159);
nand U13101 (N_13101,N_11812,N_11294);
nor U13102 (N_13102,N_11501,N_11645);
nor U13103 (N_13103,N_11482,N_11536);
and U13104 (N_13104,N_11875,N_11756);
and U13105 (N_13105,N_11762,N_10824);
and U13106 (N_13106,N_11053,N_11211);
nand U13107 (N_13107,N_10658,N_11523);
xnor U13108 (N_13108,N_10502,N_11129);
or U13109 (N_13109,N_10504,N_11091);
or U13110 (N_13110,N_11392,N_11649);
or U13111 (N_13111,N_10992,N_10775);
nor U13112 (N_13112,N_11370,N_11630);
and U13113 (N_13113,N_11207,N_10574);
nand U13114 (N_13114,N_11424,N_11002);
nand U13115 (N_13115,N_10745,N_11336);
and U13116 (N_13116,N_11138,N_10533);
nor U13117 (N_13117,N_10533,N_10693);
nor U13118 (N_13118,N_10955,N_11842);
or U13119 (N_13119,N_11064,N_11656);
nor U13120 (N_13120,N_10564,N_10683);
or U13121 (N_13121,N_10974,N_11150);
nor U13122 (N_13122,N_11204,N_11057);
nor U13123 (N_13123,N_10782,N_11122);
or U13124 (N_13124,N_11480,N_10845);
or U13125 (N_13125,N_10784,N_11998);
nor U13126 (N_13126,N_10828,N_11649);
or U13127 (N_13127,N_11819,N_11899);
nand U13128 (N_13128,N_11071,N_11749);
and U13129 (N_13129,N_11978,N_11580);
and U13130 (N_13130,N_10774,N_11679);
nand U13131 (N_13131,N_11615,N_10911);
nor U13132 (N_13132,N_11670,N_10609);
nor U13133 (N_13133,N_11310,N_11326);
xnor U13134 (N_13134,N_11881,N_10751);
nand U13135 (N_13135,N_11582,N_10992);
and U13136 (N_13136,N_11973,N_11637);
nand U13137 (N_13137,N_11743,N_11742);
or U13138 (N_13138,N_10530,N_10871);
nand U13139 (N_13139,N_10565,N_11629);
nor U13140 (N_13140,N_11456,N_11131);
or U13141 (N_13141,N_11581,N_10668);
and U13142 (N_13142,N_11366,N_10566);
xnor U13143 (N_13143,N_11759,N_11940);
nor U13144 (N_13144,N_11999,N_10917);
nor U13145 (N_13145,N_11888,N_11821);
nor U13146 (N_13146,N_11529,N_11748);
and U13147 (N_13147,N_11360,N_11934);
or U13148 (N_13148,N_11140,N_11633);
and U13149 (N_13149,N_11952,N_11538);
nor U13150 (N_13150,N_11732,N_10671);
and U13151 (N_13151,N_10864,N_10659);
and U13152 (N_13152,N_11069,N_11701);
nor U13153 (N_13153,N_11785,N_11882);
and U13154 (N_13154,N_11330,N_11878);
xor U13155 (N_13155,N_11685,N_11402);
and U13156 (N_13156,N_10673,N_10806);
or U13157 (N_13157,N_10568,N_11430);
nor U13158 (N_13158,N_11734,N_10540);
nor U13159 (N_13159,N_11100,N_11783);
nor U13160 (N_13160,N_10766,N_10955);
nand U13161 (N_13161,N_11059,N_11440);
and U13162 (N_13162,N_10557,N_10896);
or U13163 (N_13163,N_10909,N_11440);
xor U13164 (N_13164,N_11117,N_10784);
or U13165 (N_13165,N_11206,N_10708);
nand U13166 (N_13166,N_11173,N_11796);
nand U13167 (N_13167,N_10737,N_10638);
and U13168 (N_13168,N_11899,N_10852);
nand U13169 (N_13169,N_11162,N_11435);
or U13170 (N_13170,N_11545,N_10784);
or U13171 (N_13171,N_11642,N_11843);
and U13172 (N_13172,N_11440,N_10670);
nor U13173 (N_13173,N_11332,N_11281);
nand U13174 (N_13174,N_11725,N_11480);
nand U13175 (N_13175,N_11008,N_11710);
or U13176 (N_13176,N_11353,N_11690);
nand U13177 (N_13177,N_11671,N_11722);
nor U13178 (N_13178,N_10583,N_10562);
nor U13179 (N_13179,N_10797,N_10614);
nor U13180 (N_13180,N_10998,N_10668);
and U13181 (N_13181,N_10589,N_11976);
xnor U13182 (N_13182,N_10930,N_10528);
or U13183 (N_13183,N_10753,N_11777);
and U13184 (N_13184,N_10937,N_11349);
xnor U13185 (N_13185,N_11577,N_11178);
and U13186 (N_13186,N_11468,N_11198);
nor U13187 (N_13187,N_11673,N_11171);
nand U13188 (N_13188,N_10507,N_11607);
nor U13189 (N_13189,N_11585,N_11194);
and U13190 (N_13190,N_11334,N_10579);
and U13191 (N_13191,N_11489,N_11720);
xnor U13192 (N_13192,N_11520,N_11768);
xnor U13193 (N_13193,N_11676,N_10999);
or U13194 (N_13194,N_11643,N_11259);
nor U13195 (N_13195,N_10613,N_10592);
nand U13196 (N_13196,N_11121,N_11266);
or U13197 (N_13197,N_11563,N_11447);
nor U13198 (N_13198,N_11901,N_11358);
or U13199 (N_13199,N_10805,N_11918);
and U13200 (N_13200,N_11537,N_10803);
or U13201 (N_13201,N_11382,N_11476);
nor U13202 (N_13202,N_11748,N_10802);
nor U13203 (N_13203,N_11359,N_11763);
nand U13204 (N_13204,N_11633,N_11537);
nor U13205 (N_13205,N_11640,N_11053);
nand U13206 (N_13206,N_10731,N_11714);
nor U13207 (N_13207,N_10538,N_11220);
or U13208 (N_13208,N_10793,N_10892);
nor U13209 (N_13209,N_10661,N_10935);
or U13210 (N_13210,N_11950,N_10525);
xor U13211 (N_13211,N_10706,N_10778);
nor U13212 (N_13212,N_11365,N_11572);
nor U13213 (N_13213,N_11981,N_11257);
and U13214 (N_13214,N_10578,N_11450);
xnor U13215 (N_13215,N_11497,N_11182);
xor U13216 (N_13216,N_10769,N_11181);
or U13217 (N_13217,N_11051,N_10698);
and U13218 (N_13218,N_11119,N_10660);
nand U13219 (N_13219,N_11178,N_10638);
nor U13220 (N_13220,N_11746,N_11151);
nand U13221 (N_13221,N_10633,N_11253);
nand U13222 (N_13222,N_11438,N_10855);
or U13223 (N_13223,N_11633,N_11094);
nand U13224 (N_13224,N_11382,N_10701);
or U13225 (N_13225,N_11873,N_10570);
nand U13226 (N_13226,N_10840,N_10810);
xnor U13227 (N_13227,N_10647,N_11567);
nor U13228 (N_13228,N_11240,N_11249);
or U13229 (N_13229,N_11750,N_11934);
and U13230 (N_13230,N_11702,N_11004);
nand U13231 (N_13231,N_10877,N_11325);
and U13232 (N_13232,N_11390,N_11527);
nand U13233 (N_13233,N_10743,N_11681);
nand U13234 (N_13234,N_10524,N_10937);
nand U13235 (N_13235,N_11728,N_10738);
xor U13236 (N_13236,N_10846,N_11438);
nor U13237 (N_13237,N_10919,N_11064);
nor U13238 (N_13238,N_11508,N_11458);
or U13239 (N_13239,N_11332,N_11685);
and U13240 (N_13240,N_11028,N_11056);
and U13241 (N_13241,N_11481,N_10627);
or U13242 (N_13242,N_11147,N_10615);
or U13243 (N_13243,N_11860,N_11597);
xnor U13244 (N_13244,N_11522,N_10507);
nand U13245 (N_13245,N_11673,N_11451);
or U13246 (N_13246,N_10985,N_11355);
nand U13247 (N_13247,N_11692,N_10749);
or U13248 (N_13248,N_11263,N_11664);
and U13249 (N_13249,N_11945,N_11242);
nor U13250 (N_13250,N_10729,N_11210);
nor U13251 (N_13251,N_11735,N_11374);
xor U13252 (N_13252,N_11276,N_11905);
xnor U13253 (N_13253,N_11489,N_11288);
and U13254 (N_13254,N_11473,N_11563);
or U13255 (N_13255,N_10700,N_11623);
and U13256 (N_13256,N_11252,N_10955);
and U13257 (N_13257,N_11419,N_11540);
and U13258 (N_13258,N_10946,N_11219);
and U13259 (N_13259,N_11041,N_11618);
and U13260 (N_13260,N_11268,N_11397);
and U13261 (N_13261,N_11397,N_10750);
nand U13262 (N_13262,N_11483,N_10778);
nand U13263 (N_13263,N_11597,N_11715);
and U13264 (N_13264,N_10609,N_11564);
and U13265 (N_13265,N_11664,N_10822);
or U13266 (N_13266,N_10953,N_10646);
nor U13267 (N_13267,N_11407,N_10774);
nor U13268 (N_13268,N_10701,N_10727);
nor U13269 (N_13269,N_10704,N_11246);
nand U13270 (N_13270,N_10643,N_10579);
nor U13271 (N_13271,N_11895,N_11606);
or U13272 (N_13272,N_11083,N_11837);
or U13273 (N_13273,N_11970,N_10929);
nand U13274 (N_13274,N_11572,N_10774);
and U13275 (N_13275,N_11523,N_11271);
nor U13276 (N_13276,N_10866,N_11170);
nor U13277 (N_13277,N_11430,N_11723);
nor U13278 (N_13278,N_10843,N_11241);
xnor U13279 (N_13279,N_11569,N_11669);
or U13280 (N_13280,N_11983,N_10714);
nor U13281 (N_13281,N_11926,N_11303);
and U13282 (N_13282,N_11982,N_10820);
nor U13283 (N_13283,N_10589,N_11629);
nand U13284 (N_13284,N_10675,N_11296);
nor U13285 (N_13285,N_10779,N_11166);
or U13286 (N_13286,N_11299,N_11768);
and U13287 (N_13287,N_11870,N_11958);
and U13288 (N_13288,N_10893,N_10994);
nand U13289 (N_13289,N_10815,N_11219);
and U13290 (N_13290,N_11605,N_10511);
or U13291 (N_13291,N_11737,N_11640);
nor U13292 (N_13292,N_11639,N_10830);
or U13293 (N_13293,N_10635,N_11842);
nand U13294 (N_13294,N_11362,N_11834);
nand U13295 (N_13295,N_10958,N_11518);
nand U13296 (N_13296,N_10675,N_10848);
or U13297 (N_13297,N_10787,N_11078);
xor U13298 (N_13298,N_11473,N_10767);
nand U13299 (N_13299,N_11877,N_10695);
nor U13300 (N_13300,N_11327,N_10580);
nand U13301 (N_13301,N_11947,N_11335);
and U13302 (N_13302,N_10690,N_10984);
xor U13303 (N_13303,N_10576,N_10995);
and U13304 (N_13304,N_10853,N_11344);
nor U13305 (N_13305,N_11979,N_11069);
or U13306 (N_13306,N_11604,N_11372);
or U13307 (N_13307,N_10632,N_10925);
or U13308 (N_13308,N_11045,N_11339);
nand U13309 (N_13309,N_11212,N_11890);
and U13310 (N_13310,N_11179,N_11360);
and U13311 (N_13311,N_11562,N_11624);
nand U13312 (N_13312,N_10774,N_11015);
nand U13313 (N_13313,N_11046,N_10626);
and U13314 (N_13314,N_11051,N_11716);
nand U13315 (N_13315,N_11784,N_10874);
or U13316 (N_13316,N_11642,N_11080);
and U13317 (N_13317,N_10809,N_11253);
or U13318 (N_13318,N_10779,N_11793);
or U13319 (N_13319,N_10976,N_11064);
xor U13320 (N_13320,N_10703,N_11878);
or U13321 (N_13321,N_10650,N_11580);
or U13322 (N_13322,N_10897,N_11599);
nor U13323 (N_13323,N_10652,N_11302);
xnor U13324 (N_13324,N_10806,N_10884);
xor U13325 (N_13325,N_11786,N_11533);
or U13326 (N_13326,N_11003,N_11362);
nor U13327 (N_13327,N_10647,N_11750);
and U13328 (N_13328,N_11352,N_11295);
nor U13329 (N_13329,N_11942,N_10555);
nand U13330 (N_13330,N_10921,N_11832);
or U13331 (N_13331,N_10657,N_10783);
or U13332 (N_13332,N_11824,N_11346);
xnor U13333 (N_13333,N_11419,N_10925);
nor U13334 (N_13334,N_10679,N_11820);
or U13335 (N_13335,N_11592,N_11280);
and U13336 (N_13336,N_11977,N_11481);
or U13337 (N_13337,N_10653,N_10814);
or U13338 (N_13338,N_11684,N_10974);
xnor U13339 (N_13339,N_11234,N_11955);
and U13340 (N_13340,N_11871,N_11011);
nand U13341 (N_13341,N_10985,N_10964);
nor U13342 (N_13342,N_11329,N_11696);
nor U13343 (N_13343,N_10688,N_11126);
nand U13344 (N_13344,N_11656,N_11466);
nand U13345 (N_13345,N_11320,N_11052);
xnor U13346 (N_13346,N_10927,N_11100);
xnor U13347 (N_13347,N_11496,N_11219);
xor U13348 (N_13348,N_11612,N_10864);
xnor U13349 (N_13349,N_10975,N_10506);
or U13350 (N_13350,N_10914,N_11015);
or U13351 (N_13351,N_10925,N_11853);
nor U13352 (N_13352,N_10577,N_10704);
or U13353 (N_13353,N_11424,N_10673);
and U13354 (N_13354,N_11415,N_11480);
or U13355 (N_13355,N_11828,N_11137);
nand U13356 (N_13356,N_10839,N_11033);
or U13357 (N_13357,N_11877,N_11677);
or U13358 (N_13358,N_11062,N_11046);
or U13359 (N_13359,N_11327,N_11582);
and U13360 (N_13360,N_11343,N_11783);
nand U13361 (N_13361,N_10617,N_11338);
nand U13362 (N_13362,N_10807,N_11430);
nor U13363 (N_13363,N_11111,N_11746);
xnor U13364 (N_13364,N_11961,N_11042);
or U13365 (N_13365,N_11980,N_10798);
nor U13366 (N_13366,N_11830,N_11787);
or U13367 (N_13367,N_10736,N_11513);
or U13368 (N_13368,N_11606,N_11562);
or U13369 (N_13369,N_11282,N_10544);
or U13370 (N_13370,N_11623,N_10846);
or U13371 (N_13371,N_10572,N_11099);
nor U13372 (N_13372,N_10766,N_11857);
and U13373 (N_13373,N_10616,N_11775);
or U13374 (N_13374,N_11497,N_11720);
or U13375 (N_13375,N_11375,N_11633);
nor U13376 (N_13376,N_11386,N_11707);
nand U13377 (N_13377,N_11593,N_11631);
or U13378 (N_13378,N_11085,N_11660);
nor U13379 (N_13379,N_10887,N_10825);
or U13380 (N_13380,N_11251,N_11924);
and U13381 (N_13381,N_11324,N_11056);
and U13382 (N_13382,N_11147,N_11347);
or U13383 (N_13383,N_10945,N_11120);
nand U13384 (N_13384,N_10754,N_10686);
or U13385 (N_13385,N_11659,N_10580);
nor U13386 (N_13386,N_11602,N_11792);
xnor U13387 (N_13387,N_11234,N_11018);
nand U13388 (N_13388,N_11174,N_10877);
and U13389 (N_13389,N_11188,N_10758);
nand U13390 (N_13390,N_11340,N_11206);
or U13391 (N_13391,N_11222,N_11472);
and U13392 (N_13392,N_11776,N_11417);
or U13393 (N_13393,N_10736,N_11751);
nor U13394 (N_13394,N_10996,N_11887);
and U13395 (N_13395,N_10755,N_10549);
nor U13396 (N_13396,N_11580,N_11075);
nand U13397 (N_13397,N_10808,N_11698);
or U13398 (N_13398,N_11760,N_11891);
or U13399 (N_13399,N_11822,N_11684);
and U13400 (N_13400,N_10505,N_11050);
nor U13401 (N_13401,N_11597,N_11594);
or U13402 (N_13402,N_10557,N_10598);
nand U13403 (N_13403,N_10556,N_11332);
xnor U13404 (N_13404,N_10860,N_11024);
or U13405 (N_13405,N_11615,N_11302);
and U13406 (N_13406,N_11682,N_10531);
nand U13407 (N_13407,N_11558,N_10623);
and U13408 (N_13408,N_10540,N_11533);
xor U13409 (N_13409,N_10955,N_11635);
nand U13410 (N_13410,N_10898,N_10686);
nand U13411 (N_13411,N_11931,N_10517);
nor U13412 (N_13412,N_11271,N_10644);
nor U13413 (N_13413,N_11223,N_10705);
or U13414 (N_13414,N_11720,N_11630);
nand U13415 (N_13415,N_11134,N_10810);
nor U13416 (N_13416,N_10936,N_11873);
xnor U13417 (N_13417,N_11447,N_11277);
or U13418 (N_13418,N_11696,N_10700);
nor U13419 (N_13419,N_11267,N_10618);
nand U13420 (N_13420,N_11571,N_11690);
nand U13421 (N_13421,N_11587,N_10790);
nand U13422 (N_13422,N_11830,N_10781);
nor U13423 (N_13423,N_10682,N_11746);
nand U13424 (N_13424,N_11630,N_10921);
or U13425 (N_13425,N_11241,N_10614);
nor U13426 (N_13426,N_10601,N_11325);
nand U13427 (N_13427,N_11379,N_11470);
xnor U13428 (N_13428,N_11112,N_10590);
and U13429 (N_13429,N_11069,N_11855);
nor U13430 (N_13430,N_10636,N_11897);
nor U13431 (N_13431,N_11987,N_10663);
nor U13432 (N_13432,N_11866,N_11456);
nor U13433 (N_13433,N_11339,N_11816);
or U13434 (N_13434,N_11009,N_11183);
nor U13435 (N_13435,N_11583,N_11231);
nor U13436 (N_13436,N_11274,N_10690);
xnor U13437 (N_13437,N_10769,N_11378);
or U13438 (N_13438,N_11941,N_10850);
and U13439 (N_13439,N_10676,N_11759);
nand U13440 (N_13440,N_11896,N_11476);
nor U13441 (N_13441,N_11642,N_11855);
and U13442 (N_13442,N_11269,N_10725);
or U13443 (N_13443,N_11830,N_11144);
xnor U13444 (N_13444,N_10751,N_11009);
nor U13445 (N_13445,N_11480,N_11523);
nor U13446 (N_13446,N_11823,N_10502);
or U13447 (N_13447,N_10884,N_11243);
and U13448 (N_13448,N_11842,N_10889);
nor U13449 (N_13449,N_11307,N_10767);
or U13450 (N_13450,N_11355,N_10914);
or U13451 (N_13451,N_11651,N_11725);
and U13452 (N_13452,N_11237,N_11736);
or U13453 (N_13453,N_11949,N_10503);
and U13454 (N_13454,N_10922,N_10993);
and U13455 (N_13455,N_10572,N_10732);
or U13456 (N_13456,N_11156,N_11207);
or U13457 (N_13457,N_10819,N_10725);
nand U13458 (N_13458,N_11429,N_11230);
and U13459 (N_13459,N_11387,N_10631);
and U13460 (N_13460,N_11238,N_11423);
or U13461 (N_13461,N_11558,N_10580);
nor U13462 (N_13462,N_11902,N_11510);
nand U13463 (N_13463,N_10915,N_11418);
nand U13464 (N_13464,N_10715,N_11284);
nand U13465 (N_13465,N_11073,N_11238);
nand U13466 (N_13466,N_11493,N_11000);
or U13467 (N_13467,N_11646,N_11889);
nor U13468 (N_13468,N_11208,N_11739);
nor U13469 (N_13469,N_11745,N_10716);
and U13470 (N_13470,N_11200,N_11060);
and U13471 (N_13471,N_11998,N_11207);
or U13472 (N_13472,N_11323,N_11316);
xnor U13473 (N_13473,N_11011,N_10770);
nand U13474 (N_13474,N_11108,N_11596);
nand U13475 (N_13475,N_11120,N_11805);
nand U13476 (N_13476,N_10779,N_11806);
and U13477 (N_13477,N_11544,N_10912);
and U13478 (N_13478,N_11407,N_10777);
or U13479 (N_13479,N_10817,N_11665);
and U13480 (N_13480,N_11870,N_11076);
or U13481 (N_13481,N_11105,N_11788);
xnor U13482 (N_13482,N_11162,N_10867);
nor U13483 (N_13483,N_11192,N_11583);
and U13484 (N_13484,N_10590,N_11177);
and U13485 (N_13485,N_11134,N_11233);
nor U13486 (N_13486,N_10870,N_11831);
xnor U13487 (N_13487,N_11651,N_10818);
nand U13488 (N_13488,N_10756,N_11001);
nor U13489 (N_13489,N_11231,N_11377);
nor U13490 (N_13490,N_11559,N_10606);
or U13491 (N_13491,N_11146,N_11794);
nand U13492 (N_13492,N_11151,N_11160);
nand U13493 (N_13493,N_11128,N_11517);
nand U13494 (N_13494,N_10791,N_11282);
nand U13495 (N_13495,N_10686,N_11500);
or U13496 (N_13496,N_10944,N_11052);
or U13497 (N_13497,N_11600,N_10592);
nand U13498 (N_13498,N_11539,N_11107);
xnor U13499 (N_13499,N_10680,N_11687);
and U13500 (N_13500,N_12087,N_12305);
nor U13501 (N_13501,N_12724,N_12747);
xor U13502 (N_13502,N_13069,N_12862);
nand U13503 (N_13503,N_12292,N_13177);
or U13504 (N_13504,N_12112,N_12390);
xnor U13505 (N_13505,N_12071,N_12459);
and U13506 (N_13506,N_12773,N_13371);
or U13507 (N_13507,N_12059,N_13007);
or U13508 (N_13508,N_13485,N_12757);
or U13509 (N_13509,N_12870,N_12565);
nand U13510 (N_13510,N_12246,N_12906);
and U13511 (N_13511,N_12682,N_12483);
xnor U13512 (N_13512,N_12657,N_13135);
nor U13513 (N_13513,N_12984,N_13363);
nand U13514 (N_13514,N_12489,N_12027);
nor U13515 (N_13515,N_12350,N_13006);
or U13516 (N_13516,N_13410,N_13498);
or U13517 (N_13517,N_12078,N_12431);
nor U13518 (N_13518,N_12049,N_12405);
and U13519 (N_13519,N_13041,N_12374);
and U13520 (N_13520,N_12041,N_12905);
and U13521 (N_13521,N_12329,N_13122);
nor U13522 (N_13522,N_13308,N_12191);
nand U13523 (N_13523,N_13241,N_13348);
nand U13524 (N_13524,N_12019,N_13150);
and U13525 (N_13525,N_13310,N_13434);
nor U13526 (N_13526,N_12395,N_12077);
xor U13527 (N_13527,N_12408,N_12977);
nand U13528 (N_13528,N_12931,N_12532);
or U13529 (N_13529,N_13147,N_12504);
or U13530 (N_13530,N_13196,N_12451);
and U13531 (N_13531,N_13430,N_13367);
nor U13532 (N_13532,N_12605,N_12606);
nand U13533 (N_13533,N_13089,N_12326);
and U13534 (N_13534,N_13412,N_12704);
nand U13535 (N_13535,N_12879,N_12323);
nand U13536 (N_13536,N_13409,N_13232);
and U13537 (N_13537,N_12138,N_12342);
and U13538 (N_13538,N_13009,N_13372);
or U13539 (N_13539,N_12722,N_12830);
and U13540 (N_13540,N_12893,N_12332);
and U13541 (N_13541,N_12015,N_13316);
or U13542 (N_13542,N_12693,N_12691);
or U13543 (N_13543,N_12750,N_12473);
and U13544 (N_13544,N_13258,N_12120);
and U13545 (N_13545,N_12387,N_12122);
and U13546 (N_13546,N_12330,N_12419);
and U13547 (N_13547,N_12070,N_12783);
nand U13548 (N_13548,N_12232,N_12877);
nor U13549 (N_13549,N_13262,N_12766);
and U13550 (N_13550,N_12797,N_12638);
nand U13551 (N_13551,N_12658,N_13081);
or U13552 (N_13552,N_13183,N_12131);
nand U13553 (N_13553,N_12426,N_12669);
and U13554 (N_13554,N_12924,N_12527);
nor U13555 (N_13555,N_12282,N_12925);
nor U13556 (N_13556,N_13299,N_13458);
nand U13557 (N_13557,N_13428,N_13050);
and U13558 (N_13558,N_12202,N_12367);
and U13559 (N_13559,N_13438,N_13192);
nand U13560 (N_13560,N_13277,N_13231);
and U13561 (N_13561,N_13109,N_12683);
nor U13562 (N_13562,N_13392,N_12585);
nor U13563 (N_13563,N_12948,N_12018);
and U13564 (N_13564,N_12200,N_13088);
and U13565 (N_13565,N_12343,N_12793);
and U13566 (N_13566,N_12099,N_13017);
or U13567 (N_13567,N_12561,N_13380);
nor U13568 (N_13568,N_12397,N_12423);
nand U13569 (N_13569,N_13186,N_12789);
or U13570 (N_13570,N_12867,N_13357);
nor U13571 (N_13571,N_13489,N_12480);
nor U13572 (N_13572,N_12719,N_13097);
xor U13573 (N_13573,N_12438,N_12441);
or U13574 (N_13574,N_13301,N_13187);
and U13575 (N_13575,N_12577,N_13155);
and U13576 (N_13576,N_12072,N_12898);
nor U13577 (N_13577,N_13180,N_13397);
xnor U13578 (N_13578,N_12066,N_13208);
nor U13579 (N_13579,N_12567,N_13341);
or U13580 (N_13580,N_12951,N_12209);
nand U13581 (N_13581,N_13087,N_13379);
and U13582 (N_13582,N_12180,N_13045);
or U13583 (N_13583,N_12255,N_12702);
xnor U13584 (N_13584,N_12574,N_13239);
nand U13585 (N_13585,N_12083,N_12252);
or U13586 (N_13586,N_13336,N_12622);
xnor U13587 (N_13587,N_12006,N_12234);
and U13588 (N_13588,N_12111,N_13191);
and U13589 (N_13589,N_12692,N_12034);
nor U13590 (N_13590,N_12975,N_13320);
or U13591 (N_13591,N_12152,N_12067);
and U13592 (N_13592,N_13214,N_12220);
and U13593 (N_13593,N_12420,N_13100);
nand U13594 (N_13594,N_13233,N_12703);
nand U13595 (N_13595,N_13407,N_12579);
or U13596 (N_13596,N_12032,N_12626);
or U13597 (N_13597,N_12915,N_13174);
or U13598 (N_13598,N_12989,N_12449);
nor U13599 (N_13599,N_12236,N_13125);
nor U13600 (N_13600,N_12920,N_12543);
nor U13601 (N_13601,N_13390,N_12562);
or U13602 (N_13602,N_12031,N_12604);
nand U13603 (N_13603,N_12859,N_12586);
or U13604 (N_13604,N_12760,N_12164);
xnor U13605 (N_13605,N_12713,N_12617);
or U13606 (N_13606,N_12629,N_12340);
nor U13607 (N_13607,N_12641,N_12009);
nor U13608 (N_13608,N_12555,N_13153);
or U13609 (N_13609,N_12590,N_13207);
nand U13610 (N_13610,N_12721,N_12221);
or U13611 (N_13611,N_12248,N_12970);
or U13612 (N_13612,N_12318,N_12346);
and U13613 (N_13613,N_12536,N_13220);
xor U13614 (N_13614,N_12507,N_13166);
nand U13615 (N_13615,N_12681,N_13427);
nor U13616 (N_13616,N_12124,N_12229);
nand U13617 (N_13617,N_12790,N_12801);
nand U13618 (N_13618,N_12718,N_12631);
and U13619 (N_13619,N_13229,N_12444);
or U13620 (N_13620,N_13413,N_12194);
nor U13621 (N_13621,N_12936,N_12108);
and U13622 (N_13622,N_13090,N_12623);
nand U13623 (N_13623,N_12883,N_12436);
nand U13624 (N_13624,N_12291,N_12050);
nand U13625 (N_13625,N_13142,N_13033);
or U13626 (N_13626,N_12744,N_12815);
nor U13627 (N_13627,N_13286,N_12857);
nand U13628 (N_13628,N_12644,N_12685);
or U13629 (N_13629,N_12345,N_12190);
and U13630 (N_13630,N_13016,N_12647);
and U13631 (N_13631,N_12767,N_12778);
nand U13632 (N_13632,N_13243,N_13113);
nand U13633 (N_13633,N_12654,N_12466);
nor U13634 (N_13634,N_12491,N_12690);
or U13635 (N_13635,N_12937,N_12878);
xor U13636 (N_13636,N_12799,N_12934);
and U13637 (N_13637,N_13038,N_12094);
nor U13638 (N_13638,N_12554,N_12570);
and U13639 (N_13639,N_13476,N_13462);
nand U13640 (N_13640,N_12772,N_12521);
and U13641 (N_13641,N_13030,N_12950);
xnor U13642 (N_13642,N_12082,N_12795);
and U13643 (N_13643,N_13487,N_12646);
or U13644 (N_13644,N_12884,N_12380);
nor U13645 (N_13645,N_13169,N_12714);
or U13646 (N_13646,N_12996,N_13225);
nand U13647 (N_13647,N_12127,N_13394);
or U13648 (N_13648,N_12633,N_12356);
xnor U13649 (N_13649,N_13093,N_12929);
nor U13650 (N_13650,N_12860,N_12822);
xnor U13651 (N_13651,N_12674,N_12520);
and U13652 (N_13652,N_12811,N_12594);
and U13653 (N_13653,N_13012,N_12734);
and U13654 (N_13654,N_13014,N_12837);
or U13655 (N_13655,N_12065,N_12197);
or U13656 (N_13656,N_12804,N_12393);
or U13657 (N_13657,N_12228,N_13139);
or U13658 (N_13658,N_13439,N_12826);
or U13659 (N_13659,N_13193,N_12339);
or U13660 (N_13660,N_12852,N_12053);
nand U13661 (N_13661,N_12678,N_13028);
or U13662 (N_13662,N_12283,N_13337);
and U13663 (N_13663,N_13274,N_12981);
xor U13664 (N_13664,N_12814,N_13276);
nand U13665 (N_13665,N_13361,N_12875);
nand U13666 (N_13666,N_13102,N_13280);
or U13667 (N_13667,N_12680,N_12351);
and U13668 (N_13668,N_12582,N_12409);
nand U13669 (N_13669,N_12360,N_13278);
or U13670 (N_13670,N_12514,N_12497);
and U13671 (N_13671,N_12866,N_13159);
and U13672 (N_13672,N_12500,N_12551);
and U13673 (N_13673,N_12481,N_13408);
or U13674 (N_13674,N_12474,N_13035);
and U13675 (N_13675,N_12159,N_12130);
xor U13676 (N_13676,N_12776,N_13029);
or U13677 (N_13677,N_13201,N_12705);
nor U13678 (N_13678,N_12239,N_12979);
xor U13679 (N_13679,N_12132,N_13424);
or U13680 (N_13680,N_12634,N_12533);
nand U13681 (N_13681,N_12173,N_12834);
and U13682 (N_13682,N_13279,N_12188);
or U13683 (N_13683,N_12835,N_13366);
and U13684 (N_13684,N_12470,N_13256);
or U13685 (N_13685,N_12069,N_12911);
nand U13686 (N_13686,N_13449,N_12366);
and U13687 (N_13687,N_13053,N_12731);
nand U13688 (N_13688,N_12089,N_13251);
nand U13689 (N_13689,N_12935,N_13324);
nand U13690 (N_13690,N_12556,N_12103);
nor U13691 (N_13691,N_13403,N_12101);
xnor U13692 (N_13692,N_13254,N_12944);
nand U13693 (N_13693,N_12712,N_13417);
and U13694 (N_13694,N_12774,N_13161);
or U13695 (N_13695,N_12183,N_12043);
nand U13696 (N_13696,N_12257,N_12597);
xor U13697 (N_13697,N_12649,N_12385);
or U13698 (N_13698,N_13391,N_12897);
or U13699 (N_13699,N_12552,N_13168);
and U13700 (N_13700,N_12525,N_12238);
xor U13701 (N_13701,N_12081,N_13217);
or U13702 (N_13702,N_13205,N_13179);
xor U13703 (N_13703,N_12251,N_13475);
xor U13704 (N_13704,N_13211,N_12512);
and U13705 (N_13705,N_12378,N_13094);
nor U13706 (N_13706,N_13027,N_12526);
nor U13707 (N_13707,N_13369,N_13325);
nand U13708 (N_13708,N_13204,N_13343);
nand U13709 (N_13709,N_12888,N_13350);
and U13710 (N_13710,N_12439,N_13206);
or U13711 (N_13711,N_12002,N_13194);
and U13712 (N_13712,N_12416,N_12528);
or U13713 (N_13713,N_12394,N_13440);
and U13714 (N_13714,N_13025,N_13011);
and U13715 (N_13715,N_13005,N_13282);
nand U13716 (N_13716,N_12289,N_13300);
and U13717 (N_13717,N_12758,N_12918);
nand U13718 (N_13718,N_12745,N_12729);
nor U13719 (N_13719,N_12560,N_13216);
nand U13720 (N_13720,N_12843,N_13451);
nor U13721 (N_13721,N_12107,N_12913);
nor U13722 (N_13722,N_12598,N_12088);
and U13723 (N_13723,N_12335,N_12461);
or U13724 (N_13724,N_12187,N_12494);
or U13725 (N_13725,N_12240,N_13144);
xor U13726 (N_13726,N_13157,N_12794);
and U13727 (N_13727,N_12324,N_12014);
nor U13728 (N_13728,N_12307,N_12538);
and U13729 (N_13729,N_13312,N_12608);
and U13730 (N_13730,N_13178,N_13134);
nor U13731 (N_13731,N_13057,N_13074);
or U13732 (N_13732,N_12546,N_12262);
nor U13733 (N_13733,N_12095,N_13062);
or U13734 (N_13734,N_12347,N_12872);
or U13735 (N_13735,N_13288,N_13046);
nand U13736 (N_13736,N_13163,N_12261);
xnor U13737 (N_13737,N_13383,N_12425);
xnor U13738 (N_13738,N_12961,N_13387);
or U13739 (N_13739,N_13095,N_13446);
xor U13740 (N_13740,N_12237,N_13457);
nor U13741 (N_13741,N_13221,N_13215);
nor U13742 (N_13742,N_12762,N_12612);
nor U13743 (N_13743,N_12997,N_12845);
nand U13744 (N_13744,N_12084,N_12464);
and U13745 (N_13745,N_12624,N_12972);
xor U13746 (N_13746,N_12779,N_12802);
nor U13747 (N_13747,N_12973,N_12125);
xnor U13748 (N_13748,N_12457,N_13143);
and U13749 (N_13749,N_12847,N_13123);
or U13750 (N_13750,N_13411,N_12004);
nor U13751 (N_13751,N_12912,N_12696);
and U13752 (N_13752,N_12406,N_12167);
and U13753 (N_13753,N_12479,N_13461);
and U13754 (N_13754,N_12885,N_13339);
nor U13755 (N_13755,N_12825,N_12856);
nand U13756 (N_13756,N_12008,N_12170);
xnor U13757 (N_13757,N_13431,N_12672);
nor U13758 (N_13758,N_12296,N_12717);
nor U13759 (N_13759,N_13466,N_12593);
nor U13760 (N_13760,N_12381,N_13322);
or U13761 (N_13761,N_12091,N_13450);
or U13762 (N_13762,N_12012,N_13309);
nand U13763 (N_13763,N_12463,N_13447);
nand U13764 (N_13764,N_12448,N_12708);
and U13765 (N_13765,N_12388,N_12133);
or U13766 (N_13766,N_12475,N_13064);
and U13767 (N_13767,N_12576,N_13483);
xnor U13768 (N_13768,N_13078,N_12891);
nand U13769 (N_13769,N_12215,N_12478);
and U13770 (N_13770,N_12792,N_12104);
nor U13771 (N_13771,N_13026,N_12278);
or U13772 (N_13772,N_13145,N_12136);
nand U13773 (N_13773,N_13152,N_12192);
xnor U13774 (N_13774,N_12171,N_12198);
xor U13775 (N_13775,N_12035,N_13425);
nand U13776 (N_13776,N_12730,N_12816);
or U13777 (N_13777,N_12651,N_12495);
and U13778 (N_13778,N_12506,N_12735);
or U13779 (N_13779,N_13013,N_13480);
nand U13780 (N_13780,N_12761,N_12178);
or U13781 (N_13781,N_13259,N_13156);
nand U13782 (N_13782,N_12196,N_12020);
and U13783 (N_13783,N_12045,N_12829);
nand U13784 (N_13784,N_12235,N_13244);
or U13785 (N_13785,N_12341,N_12331);
nand U13786 (N_13786,N_12889,N_13465);
and U13787 (N_13787,N_12189,N_12039);
nand U13788 (N_13788,N_12454,N_12614);
nor U13789 (N_13789,N_12384,N_12317);
or U13790 (N_13790,N_12848,N_12828);
or U13791 (N_13791,N_13059,N_12595);
nand U13792 (N_13792,N_12575,N_13031);
xnor U13793 (N_13793,N_12748,N_13362);
and U13794 (N_13794,N_12844,N_12434);
or U13795 (N_13795,N_12280,N_13065);
and U13796 (N_13796,N_13120,N_13400);
and U13797 (N_13797,N_12686,N_12572);
nor U13798 (N_13798,N_12119,N_12741);
or U13799 (N_13799,N_12599,N_13154);
nand U13800 (N_13800,N_12281,N_13242);
nand U13801 (N_13801,N_13101,N_13070);
nor U13802 (N_13802,N_12573,N_12899);
nand U13803 (N_13803,N_12645,N_12440);
and U13804 (N_13804,N_12578,N_12941);
nand U13805 (N_13805,N_12616,N_12781);
nor U13806 (N_13806,N_12386,N_12222);
nor U13807 (N_13807,N_12382,N_12530);
nor U13808 (N_13808,N_13323,N_12142);
and U13809 (N_13809,N_13353,N_13080);
or U13810 (N_13810,N_13141,N_12433);
nand U13811 (N_13811,N_13401,N_12864);
xnor U13812 (N_13812,N_12135,N_12510);
and U13813 (N_13813,N_12592,N_13073);
nand U13814 (N_13814,N_12306,N_12791);
xnor U13815 (N_13815,N_12271,N_13052);
nand U13816 (N_13816,N_12224,N_13110);
nor U13817 (N_13817,N_12253,N_12338);
nand U13818 (N_13818,N_12411,N_12022);
nand U13819 (N_13819,N_12117,N_13433);
nand U13820 (N_13820,N_12610,N_13003);
xor U13821 (N_13821,N_12587,N_12179);
nand U13822 (N_13822,N_12218,N_13473);
nand U13823 (N_13823,N_12275,N_12471);
nand U13824 (N_13824,N_12967,N_13295);
or U13825 (N_13825,N_13236,N_12770);
or U13826 (N_13826,N_13092,N_13460);
and U13827 (N_13827,N_13347,N_12964);
and U13828 (N_13828,N_12571,N_12165);
nor U13829 (N_13829,N_12653,N_12694);
nor U13830 (N_13830,N_12858,N_12359);
or U13831 (N_13831,N_12186,N_13039);
nor U13832 (N_13832,N_12824,N_12214);
nand U13833 (N_13833,N_13360,N_12149);
or U13834 (N_13834,N_12226,N_13126);
nor U13835 (N_13835,N_12732,N_12619);
nand U13836 (N_13836,N_13263,N_13137);
nand U13837 (N_13837,N_12455,N_12971);
nand U13838 (N_13838,N_12499,N_12755);
nor U13839 (N_13839,N_12017,N_13048);
or U13840 (N_13840,N_13189,N_13115);
xnor U13841 (N_13841,N_13140,N_12100);
nand U13842 (N_13842,N_12817,N_13344);
and U13843 (N_13843,N_12230,N_12060);
nor U13844 (N_13844,N_13068,N_12379);
or U13845 (N_13845,N_12258,N_12273);
or U13846 (N_13846,N_12957,N_13484);
or U13847 (N_13847,N_13124,N_13112);
and U13848 (N_13848,N_13148,N_13453);
or U13849 (N_13849,N_12516,N_13010);
xor U13850 (N_13850,N_13315,N_12073);
nor U13851 (N_13851,N_12290,N_12064);
xnor U13852 (N_13852,N_12667,N_12000);
xor U13853 (N_13853,N_12524,N_13338);
and U13854 (N_13854,N_12160,N_12940);
and U13855 (N_13855,N_12569,N_13162);
nor U13856 (N_13856,N_13149,N_12371);
or U13857 (N_13857,N_12168,N_13002);
and U13858 (N_13858,N_12942,N_12450);
xnor U13859 (N_13859,N_12947,N_12472);
xor U13860 (N_13860,N_13203,N_12299);
nand U13861 (N_13861,N_12277,N_12093);
or U13862 (N_13862,N_12630,N_12810);
or U13863 (N_13863,N_13296,N_12684);
nor U13864 (N_13864,N_12163,N_12583);
nand U13865 (N_13865,N_12184,N_12410);
or U13866 (N_13866,N_12075,N_12916);
nor U13867 (N_13867,N_12563,N_12820);
or U13868 (N_13868,N_13289,N_13389);
or U13869 (N_13869,N_12819,N_12836);
nor U13870 (N_13870,N_12298,N_13294);
nand U13871 (N_13871,N_12016,N_12121);
nand U13872 (N_13872,N_13146,N_13329);
or U13873 (N_13873,N_13000,N_12033);
xor U13874 (N_13874,N_13314,N_12833);
and U13875 (N_13875,N_12739,N_12320);
nor U13876 (N_13876,N_12584,N_12661);
xnor U13877 (N_13877,N_12939,N_12021);
or U13878 (N_13878,N_12302,N_12383);
xor U13879 (N_13879,N_13266,N_13164);
nor U13880 (N_13880,N_12780,N_13429);
and U13881 (N_13881,N_13129,N_12643);
xnor U13882 (N_13882,N_12412,N_13238);
and U13883 (N_13883,N_13436,N_12508);
nand U13884 (N_13884,N_12706,N_13345);
and U13885 (N_13885,N_12659,N_12403);
and U13886 (N_13886,N_12853,N_13464);
xor U13887 (N_13887,N_12140,N_12895);
nand U13888 (N_13888,N_12547,N_12304);
nand U13889 (N_13889,N_12328,N_13319);
nor U13890 (N_13890,N_12655,N_13318);
or U13891 (N_13891,N_13273,N_13373);
nor U13892 (N_13892,N_12276,N_13245);
and U13893 (N_13893,N_13267,N_13423);
or U13894 (N_13894,N_12079,N_13086);
or U13895 (N_13895,N_13385,N_12118);
nand U13896 (N_13896,N_12851,N_12492);
and U13897 (N_13897,N_12662,N_12720);
nor U13898 (N_13898,N_13237,N_12618);
or U13899 (N_13899,N_13051,N_12648);
or U13900 (N_13900,N_12548,N_12312);
xnor U13901 (N_13901,N_12689,N_12055);
and U13902 (N_13902,N_13188,N_13224);
xor U13903 (N_13903,N_13479,N_13250);
nor U13904 (N_13904,N_13418,N_12293);
nor U13905 (N_13905,N_13377,N_12109);
or U13906 (N_13906,N_12148,N_13099);
and U13907 (N_13907,N_13328,N_12363);
nor U13908 (N_13908,N_13474,N_12223);
nor U13909 (N_13909,N_12949,N_12334);
and U13910 (N_13910,N_12010,N_12798);
nand U13911 (N_13911,N_12966,N_12496);
nor U13912 (N_13912,N_12003,N_12922);
or U13913 (N_13913,N_12764,N_13072);
nand U13914 (N_13914,N_13285,N_13018);
xor U13915 (N_13915,N_12174,N_12529);
nand U13916 (N_13916,N_12986,N_12611);
or U13917 (N_13917,N_13354,N_12746);
nand U13918 (N_13918,N_12207,N_12726);
xor U13919 (N_13919,N_13202,N_12736);
or U13920 (N_13920,N_12225,N_12498);
nand U13921 (N_13921,N_12476,N_13228);
nor U13922 (N_13922,N_13234,N_13253);
and U13923 (N_13923,N_13055,N_12699);
or U13924 (N_13924,N_12890,N_12710);
nor U13925 (N_13925,N_13032,N_13333);
nand U13926 (N_13926,N_13107,N_12509);
nand U13927 (N_13927,N_12687,N_13477);
nor U13928 (N_13928,N_12670,N_13227);
nor U13929 (N_13929,N_13198,N_12056);
and U13930 (N_13930,N_12316,N_12752);
nand U13931 (N_13931,N_13375,N_12637);
nor U13932 (N_13932,N_12876,N_13042);
and U13933 (N_13933,N_13437,N_12519);
nand U13934 (N_13934,N_12777,N_13355);
or U13935 (N_13935,N_12679,N_12621);
nor U13936 (N_13936,N_12839,N_12418);
xor U13937 (N_13937,N_13441,N_13098);
nand U13938 (N_13938,N_12580,N_12627);
nor U13939 (N_13939,N_12953,N_12782);
nand U13940 (N_13940,N_12846,N_12902);
nand U13941 (N_13941,N_12771,N_12753);
xnor U13942 (N_13942,N_13486,N_13399);
nor U13943 (N_13943,N_12697,N_12155);
nor U13944 (N_13944,N_12169,N_13036);
xor U13945 (N_13945,N_12358,N_13298);
and U13946 (N_13946,N_12542,N_13158);
nand U13947 (N_13947,N_12775,N_13118);
nor U13948 (N_13948,N_12272,N_12952);
nand U13949 (N_13949,N_13426,N_12417);
nor U13950 (N_13950,N_12854,N_12468);
or U13951 (N_13951,N_13212,N_12313);
and U13952 (N_13952,N_12665,N_12769);
and U13953 (N_13953,N_12873,N_12596);
nor U13954 (N_13954,N_13335,N_12181);
nand U13955 (N_13955,N_12377,N_12153);
nand U13956 (N_13956,N_13365,N_12227);
nor U13957 (N_13957,N_12123,N_12256);
nand U13958 (N_13958,N_12177,N_13040);
xnor U13959 (N_13959,N_12297,N_12490);
or U13960 (N_13960,N_13396,N_12295);
nand U13961 (N_13961,N_12531,N_12806);
or U13962 (N_13962,N_12357,N_13175);
or U13963 (N_13963,N_12727,N_12933);
or U13964 (N_13964,N_12965,N_13132);
nor U13965 (N_13965,N_12096,N_12432);
xor U13966 (N_13966,N_13414,N_13247);
and U13967 (N_13967,N_12245,N_12058);
or U13968 (N_13968,N_12013,N_12086);
or U13969 (N_13969,N_12503,N_13066);
xnor U13970 (N_13970,N_12663,N_12219);
or U13971 (N_13971,N_12881,N_12725);
xor U13972 (N_13972,N_12268,N_13269);
or U13973 (N_13973,N_12803,N_12541);
nand U13974 (N_13974,N_12928,N_12040);
nor U13975 (N_13975,N_13108,N_13321);
and U13976 (N_13976,N_13359,N_12517);
xor U13977 (N_13977,N_12129,N_13378);
or U13978 (N_13978,N_12005,N_12823);
nor U13979 (N_13979,N_12549,N_12901);
or U13980 (N_13980,N_12908,N_12932);
or U13981 (N_13981,N_13260,N_12400);
and U13982 (N_13982,N_12264,N_12763);
nor U13983 (N_13983,N_12141,N_12963);
and U13984 (N_13984,N_13422,N_12270);
and U13985 (N_13985,N_13172,N_13096);
and U13986 (N_13986,N_12539,N_13185);
xor U13987 (N_13987,N_12827,N_13182);
xnor U13988 (N_13988,N_13416,N_13165);
nor U13989 (N_13989,N_12211,N_13398);
nand U13990 (N_13990,N_12698,N_12182);
xor U13991 (N_13991,N_13252,N_12518);
nand U13992 (N_13992,N_12636,N_13415);
or U13993 (N_13993,N_12467,N_12676);
and U13994 (N_13994,N_13061,N_12613);
or U13995 (N_13995,N_12715,N_12716);
and U13996 (N_13996,N_13334,N_12137);
and U13997 (N_13997,N_12427,N_13272);
or U13998 (N_13998,N_13496,N_12242);
nand U13999 (N_13999,N_12892,N_12150);
and U14000 (N_14000,N_13381,N_12250);
or U14001 (N_14001,N_12743,N_12628);
nor U14002 (N_14002,N_12375,N_13459);
or U14003 (N_14003,N_12301,N_13306);
and U14004 (N_14004,N_12352,N_12660);
or U14005 (N_14005,N_12210,N_12401);
and U14006 (N_14006,N_12652,N_13302);
and U14007 (N_14007,N_13076,N_13305);
or U14008 (N_14008,N_12151,N_12603);
or U14009 (N_14009,N_12786,N_12368);
or U14010 (N_14010,N_12147,N_12909);
or U14011 (N_14011,N_13435,N_12205);
xnor U14012 (N_14012,N_12076,N_12392);
nand U14013 (N_14013,N_13481,N_12958);
or U14014 (N_14014,N_13384,N_12115);
and U14015 (N_14015,N_12999,N_12917);
nand U14016 (N_14016,N_13240,N_12092);
nand U14017 (N_14017,N_12429,N_13270);
nor U14018 (N_14018,N_12213,N_12288);
nor U14019 (N_14019,N_13127,N_12269);
nor U14020 (N_14020,N_12044,N_12267);
and U14021 (N_14021,N_13303,N_13223);
or U14022 (N_14022,N_12545,N_12456);
xnor U14023 (N_14023,N_13420,N_12788);
and U14024 (N_14024,N_12110,N_13151);
nor U14025 (N_14025,N_12675,N_13103);
xor U14026 (N_14026,N_13049,N_12442);
nor U14027 (N_14027,N_12784,N_12046);
nand U14028 (N_14028,N_13283,N_12217);
nor U14029 (N_14029,N_12796,N_12113);
nand U14030 (N_14030,N_13376,N_12303);
nand U14031 (N_14031,N_12029,N_12982);
nand U14032 (N_14032,N_13019,N_12315);
or U14033 (N_14033,N_12927,N_12868);
and U14034 (N_14034,N_12344,N_13222);
nand U14035 (N_14035,N_12588,N_13370);
xnor U14036 (N_14036,N_12144,N_13317);
xnor U14037 (N_14037,N_12907,N_13488);
or U14038 (N_14038,N_12024,N_12607);
xor U14039 (N_14039,N_13468,N_13356);
nor U14040 (N_14040,N_12068,N_12052);
nor U14041 (N_14041,N_13275,N_13463);
nand U14042 (N_14042,N_13311,N_12201);
or U14043 (N_14043,N_12208,N_12759);
and U14044 (N_14044,N_12300,N_12850);
or U14045 (N_14045,N_12286,N_12487);
nor U14046 (N_14046,N_12011,N_12821);
xnor U14047 (N_14047,N_13210,N_12337);
nor U14048 (N_14048,N_12249,N_13364);
and U14049 (N_14049,N_12443,N_13402);
xor U14050 (N_14050,N_12749,N_13004);
xnor U14051 (N_14051,N_13111,N_12640);
nand U14052 (N_14052,N_12469,N_13063);
and U14053 (N_14053,N_12404,N_12910);
nor U14054 (N_14054,N_12311,N_12399);
xor U14055 (N_14055,N_13313,N_13056);
nand U14056 (N_14056,N_12601,N_12785);
nor U14057 (N_14057,N_12945,N_13091);
nand U14058 (N_14058,N_12370,N_12143);
nand U14059 (N_14059,N_12322,N_12946);
or U14060 (N_14060,N_12711,N_12695);
nor U14061 (N_14061,N_13257,N_12513);
nand U14062 (N_14062,N_12709,N_12985);
nor U14063 (N_14063,N_13448,N_12900);
nor U14064 (N_14064,N_12284,N_12978);
xnor U14065 (N_14065,N_12145,N_13472);
or U14066 (N_14066,N_12505,N_12314);
nand U14067 (N_14067,N_13342,N_12849);
nor U14068 (N_14068,N_12493,N_12098);
or U14069 (N_14069,N_13307,N_12838);
nand U14070 (N_14070,N_12023,N_12620);
nor U14071 (N_14071,N_12048,N_13492);
and U14072 (N_14072,N_13352,N_12355);
nand U14073 (N_14073,N_12244,N_12841);
nor U14074 (N_14074,N_12051,N_13442);
or U14075 (N_14075,N_12172,N_13482);
or U14076 (N_14076,N_13291,N_13368);
nand U14077 (N_14077,N_13218,N_12193);
nor U14078 (N_14078,N_13470,N_12671);
nor U14079 (N_14079,N_13200,N_12537);
nor U14080 (N_14080,N_13495,N_13170);
nor U14081 (N_14081,N_12581,N_12740);
nor U14082 (N_14082,N_12482,N_12625);
nor U14083 (N_14083,N_12166,N_13199);
and U14084 (N_14084,N_13071,N_12501);
nand U14085 (N_14085,N_13497,N_13173);
or U14086 (N_14086,N_12212,N_12840);
xor U14087 (N_14087,N_12650,N_12589);
nor U14088 (N_14088,N_13213,N_12116);
nor U14089 (N_14089,N_12874,N_12414);
nor U14090 (N_14090,N_13190,N_12199);
or U14091 (N_14091,N_12921,N_12376);
and U14092 (N_14092,N_12751,N_13271);
or U14093 (N_14093,N_13024,N_12396);
and U14094 (N_14094,N_12600,N_12157);
or U14095 (N_14095,N_13195,N_12632);
nor U14096 (N_14096,N_12036,N_13297);
nand U14097 (N_14097,N_12156,N_12484);
nor U14098 (N_14098,N_12146,N_12259);
and U14099 (N_14099,N_12842,N_12424);
nand U14100 (N_14100,N_12274,N_13284);
or U14101 (N_14101,N_12700,N_12983);
nor U14102 (N_14102,N_13265,N_12809);
or U14103 (N_14103,N_12591,N_13281);
nor U14104 (N_14104,N_12285,N_13374);
or U14105 (N_14105,N_12001,N_13444);
xnor U14106 (N_14106,N_13404,N_13293);
nor U14107 (N_14107,N_13287,N_12511);
nor U14108 (N_14108,N_12389,N_13471);
xor U14109 (N_14109,N_12544,N_13226);
and U14110 (N_14110,N_12139,N_13114);
nand U14111 (N_14111,N_13268,N_12319);
nor U14112 (N_14112,N_12805,N_13083);
nor U14113 (N_14113,N_13406,N_12991);
xor U14114 (N_14114,N_12664,N_12522);
or U14115 (N_14115,N_12085,N_12333);
nand U14116 (N_14116,N_12994,N_13119);
and U14117 (N_14117,N_12914,N_12038);
nor U14118 (N_14118,N_12407,N_12800);
and U14119 (N_14119,N_13246,N_13264);
xor U14120 (N_14120,N_12818,N_12327);
nand U14121 (N_14121,N_13349,N_12865);
or U14122 (N_14122,N_12241,N_12061);
nor U14123 (N_14123,N_13290,N_12447);
and U14124 (N_14124,N_12437,N_12161);
nand U14125 (N_14125,N_12677,N_12765);
and U14126 (N_14126,N_12807,N_12954);
nand U14127 (N_14127,N_12254,N_12904);
nand U14128 (N_14128,N_12422,N_13001);
nand U14129 (N_14129,N_13085,N_12105);
nor U14130 (N_14130,N_13133,N_12462);
and U14131 (N_14131,N_13249,N_13395);
nand U14132 (N_14132,N_12348,N_13346);
nor U14133 (N_14133,N_12354,N_12428);
xnor U14134 (N_14134,N_12279,N_12488);
nor U14135 (N_14135,N_12446,N_12062);
nand U14136 (N_14136,N_13075,N_12486);
xnor U14137 (N_14137,N_12959,N_13037);
xor U14138 (N_14138,N_12869,N_12028);
nor U14139 (N_14139,N_12106,N_12233);
and U14140 (N_14140,N_12943,N_12688);
and U14141 (N_14141,N_12903,N_12402);
nor U14142 (N_14142,N_12263,N_13058);
and U14143 (N_14143,N_12373,N_13358);
xor U14144 (N_14144,N_12568,N_12287);
nor U14145 (N_14145,N_12266,N_13015);
nor U14146 (N_14146,N_12523,N_13060);
or U14147 (N_14147,N_12185,N_12855);
nor U14148 (N_14148,N_12362,N_13248);
nand U14149 (N_14149,N_12861,N_12321);
or U14150 (N_14150,N_12956,N_13490);
nor U14151 (N_14151,N_12832,N_12882);
xor U14152 (N_14152,N_13082,N_12502);
nor U14153 (N_14153,N_13171,N_12162);
nor U14154 (N_14154,N_12353,N_12988);
nor U14155 (N_14155,N_12886,N_12639);
and U14156 (N_14156,N_12025,N_12063);
nor U14157 (N_14157,N_12968,N_12465);
or U14158 (N_14158,N_13043,N_12026);
xnor U14159 (N_14159,N_12260,N_12042);
and U14160 (N_14160,N_13235,N_12976);
or U14161 (N_14161,N_12728,N_12325);
or U14162 (N_14162,N_13054,N_12980);
nand U14163 (N_14163,N_13067,N_13021);
and U14164 (N_14164,N_12564,N_12995);
and U14165 (N_14165,N_12880,N_12391);
nand U14166 (N_14166,N_12231,N_13181);
or U14167 (N_14167,N_13079,N_12871);
nor U14168 (N_14168,N_13138,N_13445);
nor U14169 (N_14169,N_12294,N_13327);
nand U14170 (N_14170,N_13499,N_12673);
nand U14171 (N_14171,N_12756,N_12372);
or U14172 (N_14172,N_13478,N_12308);
or U14173 (N_14173,N_12668,N_12030);
and U14174 (N_14174,N_12247,N_12707);
nor U14175 (N_14175,N_13494,N_12102);
nand U14176 (N_14176,N_12007,N_13136);
and U14177 (N_14177,N_12458,N_12887);
nor U14178 (N_14178,N_12550,N_12310);
or U14179 (N_14179,N_13160,N_12097);
nand U14180 (N_14180,N_13326,N_13044);
nand U14181 (N_14181,N_12609,N_13452);
nand U14182 (N_14182,N_13332,N_12435);
or U14183 (N_14183,N_13104,N_12926);
and U14184 (N_14184,N_12485,N_12452);
xor U14185 (N_14185,N_12787,N_13456);
and U14186 (N_14186,N_13047,N_12265);
nand U14187 (N_14187,N_13117,N_13077);
xor U14188 (N_14188,N_12534,N_12057);
nor U14189 (N_14189,N_12754,N_12566);
nor U14190 (N_14190,N_12602,N_12074);
or U14191 (N_14191,N_12080,N_12558);
nand U14192 (N_14192,N_12701,N_12894);
and U14193 (N_14193,N_12938,N_12768);
nor U14194 (N_14194,N_13351,N_12666);
and U14195 (N_14195,N_12128,N_12553);
or U14196 (N_14196,N_12430,N_12206);
nand U14197 (N_14197,N_13034,N_12930);
nand U14198 (N_14198,N_12515,N_13022);
nand U14199 (N_14199,N_12919,N_12398);
and U14200 (N_14200,N_13388,N_13340);
and U14201 (N_14201,N_12738,N_12962);
and U14202 (N_14202,N_13131,N_12413);
nor U14203 (N_14203,N_12134,N_12415);
nand U14204 (N_14204,N_12369,N_13008);
nand U14205 (N_14205,N_12987,N_12336);
nand U14206 (N_14206,N_12993,N_12453);
nand U14207 (N_14207,N_13020,N_12175);
and U14208 (N_14208,N_12126,N_13261);
nand U14209 (N_14209,N_12365,N_12960);
and U14210 (N_14210,N_12990,N_12808);
or U14211 (N_14211,N_12176,N_13330);
nand U14212 (N_14212,N_13382,N_12195);
and U14213 (N_14213,N_13455,N_12203);
nor U14214 (N_14214,N_12737,N_12047);
nand U14215 (N_14215,N_12037,N_12243);
and U14216 (N_14216,N_12054,N_12733);
and U14217 (N_14217,N_12559,N_12923);
xnor U14218 (N_14218,N_12896,N_13493);
nand U14219 (N_14219,N_12540,N_12955);
or U14220 (N_14220,N_12969,N_13084);
or U14221 (N_14221,N_12812,N_12557);
nand U14222 (N_14222,N_13386,N_13304);
nor U14223 (N_14223,N_12204,N_13116);
xor U14224 (N_14224,N_13130,N_12216);
or U14225 (N_14225,N_12831,N_13023);
xnor U14226 (N_14226,N_12813,N_12635);
nand U14227 (N_14227,N_12114,N_12723);
and U14228 (N_14228,N_13128,N_12477);
and U14229 (N_14229,N_12309,N_13331);
nor U14230 (N_14230,N_13393,N_12154);
nand U14231 (N_14231,N_13255,N_13230);
nor U14232 (N_14232,N_12364,N_12361);
nor U14233 (N_14233,N_13432,N_12863);
nand U14234 (N_14234,N_12460,N_13292);
nand U14235 (N_14235,N_12445,N_13105);
nor U14236 (N_14236,N_13467,N_12421);
nand U14237 (N_14237,N_13197,N_13421);
and U14238 (N_14238,N_12656,N_12158);
nand U14239 (N_14239,N_12742,N_12974);
or U14240 (N_14240,N_12998,N_13469);
and U14241 (N_14241,N_13167,N_13176);
or U14242 (N_14242,N_12090,N_12535);
nand U14243 (N_14243,N_12642,N_12349);
nand U14244 (N_14244,N_13106,N_13405);
nand U14245 (N_14245,N_13209,N_13491);
nor U14246 (N_14246,N_12615,N_13219);
nand U14247 (N_14247,N_13443,N_13121);
and U14248 (N_14248,N_13419,N_13184);
or U14249 (N_14249,N_13454,N_12992);
nor U14250 (N_14250,N_13471,N_13098);
and U14251 (N_14251,N_13033,N_13017);
and U14252 (N_14252,N_13319,N_13354);
nand U14253 (N_14253,N_12044,N_12358);
nand U14254 (N_14254,N_12201,N_12717);
xnor U14255 (N_14255,N_12692,N_12659);
and U14256 (N_14256,N_12681,N_13387);
nand U14257 (N_14257,N_12242,N_12054);
and U14258 (N_14258,N_13200,N_12876);
nor U14259 (N_14259,N_12846,N_13170);
nand U14260 (N_14260,N_13015,N_12234);
nor U14261 (N_14261,N_12800,N_12375);
nand U14262 (N_14262,N_13434,N_13031);
nor U14263 (N_14263,N_12788,N_13153);
and U14264 (N_14264,N_13237,N_12901);
nand U14265 (N_14265,N_12979,N_13144);
nand U14266 (N_14266,N_12511,N_12350);
nand U14267 (N_14267,N_13411,N_12450);
xnor U14268 (N_14268,N_12144,N_12528);
or U14269 (N_14269,N_12052,N_13232);
and U14270 (N_14270,N_13323,N_13381);
nor U14271 (N_14271,N_13266,N_12517);
nor U14272 (N_14272,N_12162,N_13433);
xnor U14273 (N_14273,N_12974,N_12749);
nand U14274 (N_14274,N_12336,N_12470);
and U14275 (N_14275,N_13248,N_12254);
and U14276 (N_14276,N_12644,N_13114);
or U14277 (N_14277,N_12352,N_12954);
nand U14278 (N_14278,N_12935,N_13232);
or U14279 (N_14279,N_12254,N_12443);
or U14280 (N_14280,N_12125,N_12944);
nor U14281 (N_14281,N_13307,N_12567);
xor U14282 (N_14282,N_12741,N_12894);
nand U14283 (N_14283,N_12108,N_13274);
and U14284 (N_14284,N_12338,N_13328);
xnor U14285 (N_14285,N_12134,N_12489);
nand U14286 (N_14286,N_13176,N_12881);
nand U14287 (N_14287,N_12278,N_13403);
nor U14288 (N_14288,N_12504,N_12069);
and U14289 (N_14289,N_13253,N_12594);
and U14290 (N_14290,N_12448,N_13162);
nand U14291 (N_14291,N_13259,N_13237);
or U14292 (N_14292,N_12322,N_12452);
xnor U14293 (N_14293,N_13145,N_13336);
or U14294 (N_14294,N_13233,N_12096);
nor U14295 (N_14295,N_13062,N_13401);
nor U14296 (N_14296,N_12388,N_12356);
xnor U14297 (N_14297,N_13099,N_13398);
nor U14298 (N_14298,N_13329,N_12476);
nand U14299 (N_14299,N_12284,N_13096);
xnor U14300 (N_14300,N_12665,N_13043);
nor U14301 (N_14301,N_12728,N_13476);
nand U14302 (N_14302,N_13349,N_12164);
nand U14303 (N_14303,N_12831,N_12613);
or U14304 (N_14304,N_12462,N_13177);
and U14305 (N_14305,N_12801,N_13200);
and U14306 (N_14306,N_13139,N_12683);
and U14307 (N_14307,N_12043,N_12710);
nand U14308 (N_14308,N_12463,N_12555);
nand U14309 (N_14309,N_12840,N_12762);
nand U14310 (N_14310,N_13250,N_12459);
xnor U14311 (N_14311,N_13155,N_12695);
nand U14312 (N_14312,N_12406,N_12874);
and U14313 (N_14313,N_12579,N_13054);
nor U14314 (N_14314,N_12670,N_12421);
nand U14315 (N_14315,N_13380,N_12218);
nand U14316 (N_14316,N_12941,N_13038);
nor U14317 (N_14317,N_12620,N_12880);
nand U14318 (N_14318,N_13408,N_13454);
and U14319 (N_14319,N_12820,N_12708);
nand U14320 (N_14320,N_13425,N_12573);
and U14321 (N_14321,N_12389,N_13016);
or U14322 (N_14322,N_12477,N_13291);
nor U14323 (N_14323,N_13479,N_13243);
or U14324 (N_14324,N_13338,N_12428);
xor U14325 (N_14325,N_13032,N_13409);
or U14326 (N_14326,N_12802,N_12375);
or U14327 (N_14327,N_12336,N_13040);
and U14328 (N_14328,N_12471,N_13164);
nor U14329 (N_14329,N_12580,N_13087);
or U14330 (N_14330,N_13244,N_12658);
or U14331 (N_14331,N_12050,N_12062);
and U14332 (N_14332,N_12759,N_13254);
nor U14333 (N_14333,N_13492,N_12155);
or U14334 (N_14334,N_13458,N_12072);
nand U14335 (N_14335,N_12510,N_12264);
xnor U14336 (N_14336,N_13359,N_12369);
or U14337 (N_14337,N_12874,N_12117);
nor U14338 (N_14338,N_12833,N_12034);
nand U14339 (N_14339,N_13247,N_12977);
or U14340 (N_14340,N_12150,N_12271);
nor U14341 (N_14341,N_12454,N_13359);
or U14342 (N_14342,N_12493,N_13223);
xnor U14343 (N_14343,N_12507,N_12506);
and U14344 (N_14344,N_13370,N_13243);
or U14345 (N_14345,N_12514,N_13240);
and U14346 (N_14346,N_12931,N_12134);
xnor U14347 (N_14347,N_13147,N_12272);
and U14348 (N_14348,N_12747,N_13040);
xor U14349 (N_14349,N_12357,N_13300);
nand U14350 (N_14350,N_13478,N_13132);
and U14351 (N_14351,N_12136,N_13227);
nand U14352 (N_14352,N_13408,N_12315);
and U14353 (N_14353,N_12986,N_12796);
and U14354 (N_14354,N_12092,N_12235);
or U14355 (N_14355,N_12988,N_12865);
or U14356 (N_14356,N_12848,N_13423);
nor U14357 (N_14357,N_12550,N_13055);
or U14358 (N_14358,N_12767,N_12553);
nor U14359 (N_14359,N_12744,N_12399);
xor U14360 (N_14360,N_13443,N_12979);
nand U14361 (N_14361,N_12756,N_12702);
or U14362 (N_14362,N_13047,N_13422);
nor U14363 (N_14363,N_13099,N_13358);
nor U14364 (N_14364,N_12922,N_13253);
nand U14365 (N_14365,N_13186,N_13185);
or U14366 (N_14366,N_12621,N_12415);
or U14367 (N_14367,N_12488,N_13409);
nor U14368 (N_14368,N_12824,N_12576);
nor U14369 (N_14369,N_13252,N_12564);
nand U14370 (N_14370,N_12832,N_13428);
nor U14371 (N_14371,N_12840,N_13457);
xor U14372 (N_14372,N_12641,N_13304);
nand U14373 (N_14373,N_13346,N_12670);
nand U14374 (N_14374,N_12302,N_12626);
or U14375 (N_14375,N_13066,N_13325);
nor U14376 (N_14376,N_12442,N_13440);
or U14377 (N_14377,N_12101,N_12202);
and U14378 (N_14378,N_12247,N_13130);
and U14379 (N_14379,N_12960,N_13293);
and U14380 (N_14380,N_12364,N_12635);
or U14381 (N_14381,N_12592,N_12462);
and U14382 (N_14382,N_13418,N_13287);
and U14383 (N_14383,N_13333,N_12584);
nand U14384 (N_14384,N_13019,N_13297);
and U14385 (N_14385,N_13263,N_12289);
and U14386 (N_14386,N_12610,N_12811);
nand U14387 (N_14387,N_13063,N_12971);
and U14388 (N_14388,N_12102,N_13027);
and U14389 (N_14389,N_12369,N_13303);
and U14390 (N_14390,N_12344,N_12041);
nor U14391 (N_14391,N_12709,N_12088);
and U14392 (N_14392,N_13455,N_12266);
nor U14393 (N_14393,N_12961,N_13306);
xnor U14394 (N_14394,N_13016,N_13256);
nor U14395 (N_14395,N_12933,N_13486);
and U14396 (N_14396,N_12710,N_12177);
nand U14397 (N_14397,N_12638,N_12808);
and U14398 (N_14398,N_12004,N_12230);
or U14399 (N_14399,N_12600,N_13297);
xor U14400 (N_14400,N_13196,N_13034);
nor U14401 (N_14401,N_12328,N_12702);
nand U14402 (N_14402,N_12634,N_12556);
nand U14403 (N_14403,N_12683,N_12370);
nand U14404 (N_14404,N_12551,N_13059);
or U14405 (N_14405,N_12813,N_13134);
nand U14406 (N_14406,N_12908,N_13192);
xor U14407 (N_14407,N_12715,N_12445);
and U14408 (N_14408,N_12084,N_13148);
and U14409 (N_14409,N_12392,N_12798);
nand U14410 (N_14410,N_12261,N_12305);
or U14411 (N_14411,N_12872,N_12690);
nand U14412 (N_14412,N_12667,N_12814);
nor U14413 (N_14413,N_13152,N_12098);
and U14414 (N_14414,N_12455,N_12107);
or U14415 (N_14415,N_12585,N_13237);
or U14416 (N_14416,N_13081,N_12452);
nor U14417 (N_14417,N_12777,N_13151);
xor U14418 (N_14418,N_12001,N_13106);
and U14419 (N_14419,N_12307,N_13066);
or U14420 (N_14420,N_12570,N_13120);
nand U14421 (N_14421,N_13047,N_12130);
nor U14422 (N_14422,N_12014,N_12851);
nor U14423 (N_14423,N_12999,N_12491);
nand U14424 (N_14424,N_13119,N_12379);
or U14425 (N_14425,N_12965,N_12461);
nor U14426 (N_14426,N_12904,N_12227);
nor U14427 (N_14427,N_13483,N_12787);
nor U14428 (N_14428,N_13081,N_12546);
and U14429 (N_14429,N_12662,N_12105);
or U14430 (N_14430,N_12791,N_12293);
nor U14431 (N_14431,N_13005,N_12867);
or U14432 (N_14432,N_12955,N_13240);
nor U14433 (N_14433,N_12145,N_13009);
nor U14434 (N_14434,N_12064,N_12808);
or U14435 (N_14435,N_13374,N_12450);
and U14436 (N_14436,N_12917,N_12300);
nor U14437 (N_14437,N_13454,N_12461);
nor U14438 (N_14438,N_13466,N_13131);
or U14439 (N_14439,N_13216,N_12331);
nor U14440 (N_14440,N_12743,N_13063);
or U14441 (N_14441,N_12296,N_13284);
or U14442 (N_14442,N_12782,N_13422);
and U14443 (N_14443,N_13295,N_12914);
nand U14444 (N_14444,N_13380,N_12376);
nand U14445 (N_14445,N_13198,N_12644);
xnor U14446 (N_14446,N_12989,N_13195);
or U14447 (N_14447,N_12172,N_13485);
nand U14448 (N_14448,N_12844,N_12512);
or U14449 (N_14449,N_12944,N_12473);
xor U14450 (N_14450,N_12220,N_12324);
nor U14451 (N_14451,N_13252,N_12234);
or U14452 (N_14452,N_12258,N_13437);
and U14453 (N_14453,N_12888,N_12343);
and U14454 (N_14454,N_13354,N_12373);
nor U14455 (N_14455,N_12106,N_12379);
xnor U14456 (N_14456,N_12853,N_13321);
or U14457 (N_14457,N_13456,N_12945);
or U14458 (N_14458,N_13100,N_13276);
and U14459 (N_14459,N_12026,N_12167);
xor U14460 (N_14460,N_12875,N_12343);
nand U14461 (N_14461,N_12918,N_12677);
and U14462 (N_14462,N_12648,N_12127);
nor U14463 (N_14463,N_12515,N_12748);
nand U14464 (N_14464,N_12728,N_12523);
nor U14465 (N_14465,N_13109,N_13011);
nand U14466 (N_14466,N_13053,N_12111);
nand U14467 (N_14467,N_12479,N_12239);
nor U14468 (N_14468,N_13164,N_12829);
or U14469 (N_14469,N_12816,N_12359);
or U14470 (N_14470,N_13356,N_13299);
nor U14471 (N_14471,N_13117,N_12971);
or U14472 (N_14472,N_12523,N_12347);
nor U14473 (N_14473,N_12626,N_12050);
xor U14474 (N_14474,N_12958,N_13348);
nor U14475 (N_14475,N_13034,N_12174);
and U14476 (N_14476,N_12477,N_12910);
nand U14477 (N_14477,N_13177,N_12688);
and U14478 (N_14478,N_12844,N_12011);
nand U14479 (N_14479,N_12785,N_12989);
nand U14480 (N_14480,N_13356,N_12124);
nor U14481 (N_14481,N_12942,N_13363);
nand U14482 (N_14482,N_13253,N_12338);
nor U14483 (N_14483,N_12086,N_13048);
xor U14484 (N_14484,N_12674,N_12723);
nor U14485 (N_14485,N_12443,N_13188);
nand U14486 (N_14486,N_13422,N_12216);
or U14487 (N_14487,N_13047,N_12667);
or U14488 (N_14488,N_12671,N_13047);
nand U14489 (N_14489,N_12723,N_12380);
or U14490 (N_14490,N_12404,N_12420);
and U14491 (N_14491,N_13034,N_13036);
or U14492 (N_14492,N_12455,N_13446);
and U14493 (N_14493,N_12527,N_12069);
nor U14494 (N_14494,N_12161,N_12641);
or U14495 (N_14495,N_12865,N_12877);
and U14496 (N_14496,N_13286,N_12525);
and U14497 (N_14497,N_12251,N_13165);
nor U14498 (N_14498,N_13211,N_12008);
nand U14499 (N_14499,N_13470,N_12139);
or U14500 (N_14500,N_13040,N_13272);
and U14501 (N_14501,N_12160,N_12941);
or U14502 (N_14502,N_12156,N_12514);
or U14503 (N_14503,N_13455,N_13484);
nor U14504 (N_14504,N_13172,N_12414);
nand U14505 (N_14505,N_12286,N_12339);
nand U14506 (N_14506,N_13367,N_13353);
or U14507 (N_14507,N_12035,N_13439);
nor U14508 (N_14508,N_12565,N_12529);
nor U14509 (N_14509,N_13042,N_12183);
and U14510 (N_14510,N_13217,N_12438);
nand U14511 (N_14511,N_12494,N_12549);
nand U14512 (N_14512,N_12341,N_12641);
nor U14513 (N_14513,N_12047,N_13143);
nor U14514 (N_14514,N_12510,N_12893);
or U14515 (N_14515,N_12562,N_12159);
and U14516 (N_14516,N_13036,N_12381);
or U14517 (N_14517,N_12154,N_12353);
and U14518 (N_14518,N_12413,N_13487);
and U14519 (N_14519,N_13380,N_12791);
nor U14520 (N_14520,N_12747,N_13066);
nand U14521 (N_14521,N_12353,N_12824);
nor U14522 (N_14522,N_12281,N_13114);
and U14523 (N_14523,N_13466,N_12558);
nand U14524 (N_14524,N_12578,N_12789);
or U14525 (N_14525,N_13224,N_12592);
or U14526 (N_14526,N_12016,N_12935);
nand U14527 (N_14527,N_12246,N_12188);
or U14528 (N_14528,N_12300,N_12778);
nor U14529 (N_14529,N_13318,N_12698);
or U14530 (N_14530,N_12178,N_12894);
nor U14531 (N_14531,N_12457,N_12613);
nand U14532 (N_14532,N_12813,N_13235);
xnor U14533 (N_14533,N_13045,N_12932);
nor U14534 (N_14534,N_12893,N_13165);
nand U14535 (N_14535,N_12334,N_12494);
and U14536 (N_14536,N_12632,N_12255);
xor U14537 (N_14537,N_12682,N_12619);
and U14538 (N_14538,N_12621,N_12386);
or U14539 (N_14539,N_13235,N_12360);
nor U14540 (N_14540,N_12939,N_13064);
nor U14541 (N_14541,N_13088,N_12559);
and U14542 (N_14542,N_13287,N_13045);
nor U14543 (N_14543,N_12046,N_13271);
and U14544 (N_14544,N_12363,N_12142);
nor U14545 (N_14545,N_12259,N_12385);
nand U14546 (N_14546,N_12680,N_13095);
nor U14547 (N_14547,N_12388,N_12979);
xnor U14548 (N_14548,N_13020,N_12267);
nor U14549 (N_14549,N_12999,N_13341);
nor U14550 (N_14550,N_12368,N_12317);
nand U14551 (N_14551,N_12034,N_12397);
nor U14552 (N_14552,N_12476,N_12369);
and U14553 (N_14553,N_12161,N_12642);
nor U14554 (N_14554,N_13447,N_12151);
nor U14555 (N_14555,N_13273,N_13121);
or U14556 (N_14556,N_12388,N_13227);
xor U14557 (N_14557,N_12261,N_12489);
or U14558 (N_14558,N_13435,N_12952);
xor U14559 (N_14559,N_12906,N_12346);
nor U14560 (N_14560,N_12593,N_13327);
or U14561 (N_14561,N_13304,N_13132);
or U14562 (N_14562,N_12036,N_12820);
and U14563 (N_14563,N_13195,N_12574);
and U14564 (N_14564,N_13166,N_12629);
nand U14565 (N_14565,N_13160,N_13084);
and U14566 (N_14566,N_13103,N_12369);
nor U14567 (N_14567,N_12334,N_12987);
nor U14568 (N_14568,N_13307,N_12378);
nor U14569 (N_14569,N_13182,N_13243);
or U14570 (N_14570,N_12869,N_12066);
nand U14571 (N_14571,N_12195,N_13067);
nor U14572 (N_14572,N_12652,N_13012);
and U14573 (N_14573,N_12412,N_13208);
or U14574 (N_14574,N_13055,N_13169);
or U14575 (N_14575,N_12907,N_12897);
nand U14576 (N_14576,N_12082,N_13181);
and U14577 (N_14577,N_13307,N_13131);
nand U14578 (N_14578,N_12637,N_12813);
and U14579 (N_14579,N_13080,N_13149);
or U14580 (N_14580,N_12844,N_12359);
nand U14581 (N_14581,N_12880,N_12084);
and U14582 (N_14582,N_13120,N_13415);
nand U14583 (N_14583,N_12916,N_12935);
nor U14584 (N_14584,N_13494,N_12271);
and U14585 (N_14585,N_12289,N_12703);
nand U14586 (N_14586,N_12954,N_12265);
nand U14587 (N_14587,N_12843,N_12589);
nor U14588 (N_14588,N_12845,N_13265);
nand U14589 (N_14589,N_12183,N_12386);
nand U14590 (N_14590,N_13333,N_12835);
and U14591 (N_14591,N_12946,N_12177);
xor U14592 (N_14592,N_12534,N_12218);
nor U14593 (N_14593,N_13465,N_12446);
and U14594 (N_14594,N_12308,N_12156);
or U14595 (N_14595,N_12475,N_13117);
xnor U14596 (N_14596,N_12168,N_12623);
or U14597 (N_14597,N_13455,N_12783);
nor U14598 (N_14598,N_13101,N_13433);
nor U14599 (N_14599,N_13427,N_13489);
nand U14600 (N_14600,N_12564,N_13289);
or U14601 (N_14601,N_12940,N_12275);
and U14602 (N_14602,N_12259,N_12990);
nor U14603 (N_14603,N_13307,N_12968);
nand U14604 (N_14604,N_12619,N_13171);
nand U14605 (N_14605,N_13484,N_13122);
nor U14606 (N_14606,N_12481,N_12037);
nand U14607 (N_14607,N_13087,N_12982);
and U14608 (N_14608,N_12120,N_13328);
nor U14609 (N_14609,N_12356,N_12162);
nor U14610 (N_14610,N_13109,N_12198);
nor U14611 (N_14611,N_13343,N_12465);
and U14612 (N_14612,N_13402,N_12440);
nand U14613 (N_14613,N_12648,N_13361);
or U14614 (N_14614,N_12481,N_12528);
or U14615 (N_14615,N_12325,N_13409);
and U14616 (N_14616,N_12344,N_12629);
nor U14617 (N_14617,N_12922,N_12051);
or U14618 (N_14618,N_13448,N_12408);
and U14619 (N_14619,N_12749,N_12950);
nand U14620 (N_14620,N_13043,N_12971);
nand U14621 (N_14621,N_13399,N_13218);
and U14622 (N_14622,N_13172,N_12869);
and U14623 (N_14623,N_13159,N_12578);
nand U14624 (N_14624,N_13078,N_13356);
or U14625 (N_14625,N_12240,N_12183);
and U14626 (N_14626,N_13413,N_12869);
nand U14627 (N_14627,N_12303,N_13497);
xnor U14628 (N_14628,N_12989,N_13083);
nand U14629 (N_14629,N_12150,N_12062);
nor U14630 (N_14630,N_12656,N_13332);
and U14631 (N_14631,N_12745,N_12317);
nand U14632 (N_14632,N_12007,N_12543);
and U14633 (N_14633,N_12049,N_12637);
or U14634 (N_14634,N_12237,N_13456);
or U14635 (N_14635,N_13169,N_12971);
nand U14636 (N_14636,N_12299,N_13269);
xnor U14637 (N_14637,N_12660,N_12035);
or U14638 (N_14638,N_12626,N_12202);
nor U14639 (N_14639,N_12760,N_12303);
nor U14640 (N_14640,N_12008,N_12090);
or U14641 (N_14641,N_12562,N_12957);
and U14642 (N_14642,N_13376,N_12227);
nor U14643 (N_14643,N_12648,N_13192);
and U14644 (N_14644,N_12545,N_13110);
xor U14645 (N_14645,N_12100,N_12966);
nand U14646 (N_14646,N_12745,N_12917);
nor U14647 (N_14647,N_12272,N_13385);
or U14648 (N_14648,N_12901,N_12404);
or U14649 (N_14649,N_13463,N_12407);
xor U14650 (N_14650,N_12714,N_12003);
and U14651 (N_14651,N_12505,N_12106);
nor U14652 (N_14652,N_12323,N_13161);
and U14653 (N_14653,N_13116,N_12770);
and U14654 (N_14654,N_13180,N_12809);
nand U14655 (N_14655,N_13356,N_13118);
or U14656 (N_14656,N_13324,N_12368);
and U14657 (N_14657,N_12782,N_13084);
and U14658 (N_14658,N_13234,N_13100);
nor U14659 (N_14659,N_12073,N_13279);
nor U14660 (N_14660,N_13358,N_13211);
or U14661 (N_14661,N_13219,N_12595);
nand U14662 (N_14662,N_12837,N_12353);
or U14663 (N_14663,N_12023,N_12936);
xor U14664 (N_14664,N_12018,N_12078);
nor U14665 (N_14665,N_13105,N_13093);
nor U14666 (N_14666,N_12150,N_12468);
nand U14667 (N_14667,N_12259,N_13361);
or U14668 (N_14668,N_13466,N_13381);
and U14669 (N_14669,N_12935,N_13213);
and U14670 (N_14670,N_13461,N_13067);
or U14671 (N_14671,N_13444,N_12236);
or U14672 (N_14672,N_12523,N_12849);
or U14673 (N_14673,N_13122,N_12244);
and U14674 (N_14674,N_13308,N_12525);
and U14675 (N_14675,N_13167,N_13244);
nand U14676 (N_14676,N_12378,N_12263);
nand U14677 (N_14677,N_13425,N_12713);
or U14678 (N_14678,N_13155,N_13063);
and U14679 (N_14679,N_12297,N_13388);
and U14680 (N_14680,N_13467,N_12496);
nor U14681 (N_14681,N_12720,N_13319);
xor U14682 (N_14682,N_12723,N_12584);
and U14683 (N_14683,N_12071,N_12989);
nand U14684 (N_14684,N_13444,N_12736);
or U14685 (N_14685,N_12452,N_12075);
or U14686 (N_14686,N_12957,N_12113);
and U14687 (N_14687,N_13395,N_12896);
or U14688 (N_14688,N_12429,N_12054);
or U14689 (N_14689,N_12305,N_12054);
or U14690 (N_14690,N_12486,N_13389);
nor U14691 (N_14691,N_13284,N_12285);
xor U14692 (N_14692,N_12381,N_12814);
nand U14693 (N_14693,N_12516,N_13379);
and U14694 (N_14694,N_12804,N_12631);
nand U14695 (N_14695,N_13432,N_13201);
or U14696 (N_14696,N_13180,N_13312);
xnor U14697 (N_14697,N_12372,N_12132);
xnor U14698 (N_14698,N_13138,N_13018);
nor U14699 (N_14699,N_12040,N_13237);
or U14700 (N_14700,N_12636,N_13491);
nor U14701 (N_14701,N_12961,N_12175);
or U14702 (N_14702,N_13053,N_12620);
xnor U14703 (N_14703,N_12932,N_12361);
nor U14704 (N_14704,N_12823,N_13305);
or U14705 (N_14705,N_13154,N_12035);
or U14706 (N_14706,N_12599,N_13055);
or U14707 (N_14707,N_13374,N_12216);
nand U14708 (N_14708,N_12627,N_13335);
nand U14709 (N_14709,N_12371,N_12354);
and U14710 (N_14710,N_13233,N_13470);
nor U14711 (N_14711,N_12194,N_13443);
or U14712 (N_14712,N_12030,N_12334);
nor U14713 (N_14713,N_12477,N_12887);
nand U14714 (N_14714,N_12393,N_12202);
xnor U14715 (N_14715,N_12721,N_12376);
and U14716 (N_14716,N_12084,N_12373);
nor U14717 (N_14717,N_12351,N_12337);
and U14718 (N_14718,N_12913,N_12232);
nor U14719 (N_14719,N_12437,N_12218);
and U14720 (N_14720,N_12478,N_12396);
or U14721 (N_14721,N_13330,N_12556);
or U14722 (N_14722,N_13364,N_12785);
nor U14723 (N_14723,N_12544,N_12098);
and U14724 (N_14724,N_12534,N_12711);
nand U14725 (N_14725,N_13340,N_13224);
nor U14726 (N_14726,N_12544,N_12015);
or U14727 (N_14727,N_12166,N_12864);
nand U14728 (N_14728,N_13094,N_12073);
or U14729 (N_14729,N_12575,N_12594);
nor U14730 (N_14730,N_12705,N_12603);
and U14731 (N_14731,N_12249,N_12926);
and U14732 (N_14732,N_12376,N_13320);
and U14733 (N_14733,N_12746,N_12081);
and U14734 (N_14734,N_12797,N_12101);
xnor U14735 (N_14735,N_12802,N_13305);
nand U14736 (N_14736,N_13229,N_12586);
nor U14737 (N_14737,N_12715,N_12108);
xor U14738 (N_14738,N_12432,N_12104);
nor U14739 (N_14739,N_12787,N_12278);
or U14740 (N_14740,N_12425,N_13005);
and U14741 (N_14741,N_12533,N_12962);
and U14742 (N_14742,N_12978,N_13161);
or U14743 (N_14743,N_12296,N_12271);
nor U14744 (N_14744,N_12104,N_12498);
nor U14745 (N_14745,N_13497,N_12273);
nor U14746 (N_14746,N_12596,N_12166);
or U14747 (N_14747,N_13388,N_13409);
and U14748 (N_14748,N_12956,N_12905);
nand U14749 (N_14749,N_12451,N_13360);
nor U14750 (N_14750,N_12099,N_13349);
or U14751 (N_14751,N_13176,N_12124);
nor U14752 (N_14752,N_13072,N_12194);
and U14753 (N_14753,N_12111,N_13377);
nand U14754 (N_14754,N_12355,N_12792);
nand U14755 (N_14755,N_12332,N_12956);
and U14756 (N_14756,N_12539,N_12841);
and U14757 (N_14757,N_13346,N_13325);
nand U14758 (N_14758,N_12373,N_12695);
xor U14759 (N_14759,N_13079,N_12375);
nand U14760 (N_14760,N_12946,N_13012);
and U14761 (N_14761,N_12637,N_12932);
or U14762 (N_14762,N_12996,N_12648);
nand U14763 (N_14763,N_12060,N_12038);
nand U14764 (N_14764,N_13499,N_12540);
nand U14765 (N_14765,N_13279,N_13232);
or U14766 (N_14766,N_13051,N_13222);
nand U14767 (N_14767,N_12505,N_13187);
xor U14768 (N_14768,N_12867,N_13319);
nand U14769 (N_14769,N_12900,N_13318);
and U14770 (N_14770,N_13101,N_12386);
nor U14771 (N_14771,N_12360,N_12956);
or U14772 (N_14772,N_12516,N_12912);
nand U14773 (N_14773,N_12729,N_13172);
and U14774 (N_14774,N_12693,N_12091);
and U14775 (N_14775,N_12487,N_12412);
nor U14776 (N_14776,N_12783,N_13411);
nand U14777 (N_14777,N_13020,N_12634);
or U14778 (N_14778,N_12936,N_13290);
and U14779 (N_14779,N_12674,N_12230);
and U14780 (N_14780,N_13216,N_12888);
nand U14781 (N_14781,N_13023,N_13186);
nand U14782 (N_14782,N_12631,N_13481);
or U14783 (N_14783,N_13381,N_12553);
nor U14784 (N_14784,N_13206,N_12484);
and U14785 (N_14785,N_12413,N_13021);
nand U14786 (N_14786,N_12101,N_13275);
nor U14787 (N_14787,N_12169,N_12418);
and U14788 (N_14788,N_12701,N_12003);
and U14789 (N_14789,N_13201,N_12247);
xor U14790 (N_14790,N_13378,N_13016);
nor U14791 (N_14791,N_13256,N_12863);
or U14792 (N_14792,N_12261,N_12688);
and U14793 (N_14793,N_12387,N_12282);
and U14794 (N_14794,N_13173,N_12274);
and U14795 (N_14795,N_12556,N_12908);
and U14796 (N_14796,N_12100,N_12047);
xor U14797 (N_14797,N_12336,N_13349);
or U14798 (N_14798,N_12396,N_12033);
nor U14799 (N_14799,N_12196,N_12451);
nand U14800 (N_14800,N_12401,N_13388);
xnor U14801 (N_14801,N_12976,N_12429);
nand U14802 (N_14802,N_12324,N_13463);
and U14803 (N_14803,N_12015,N_12244);
xor U14804 (N_14804,N_12599,N_13037);
or U14805 (N_14805,N_13332,N_12437);
nand U14806 (N_14806,N_12541,N_13409);
nand U14807 (N_14807,N_12086,N_12554);
and U14808 (N_14808,N_12618,N_12426);
nand U14809 (N_14809,N_13357,N_13033);
nor U14810 (N_14810,N_12128,N_12616);
or U14811 (N_14811,N_12589,N_13037);
or U14812 (N_14812,N_12111,N_12987);
or U14813 (N_14813,N_13220,N_13237);
nand U14814 (N_14814,N_12776,N_12069);
xnor U14815 (N_14815,N_12198,N_12653);
or U14816 (N_14816,N_13073,N_12941);
nand U14817 (N_14817,N_12858,N_13270);
nand U14818 (N_14818,N_13181,N_12942);
or U14819 (N_14819,N_12967,N_12231);
or U14820 (N_14820,N_12947,N_12203);
and U14821 (N_14821,N_13225,N_12911);
nor U14822 (N_14822,N_13215,N_12864);
xor U14823 (N_14823,N_12670,N_12978);
nor U14824 (N_14824,N_12072,N_12791);
nor U14825 (N_14825,N_12225,N_12819);
nor U14826 (N_14826,N_12308,N_12526);
or U14827 (N_14827,N_13435,N_12472);
or U14828 (N_14828,N_13120,N_13411);
nor U14829 (N_14829,N_12416,N_13240);
and U14830 (N_14830,N_12088,N_13251);
nor U14831 (N_14831,N_12042,N_13366);
and U14832 (N_14832,N_12060,N_12796);
xnor U14833 (N_14833,N_13440,N_12686);
or U14834 (N_14834,N_13163,N_12723);
nor U14835 (N_14835,N_12256,N_12711);
nor U14836 (N_14836,N_12276,N_13036);
and U14837 (N_14837,N_13112,N_12046);
xnor U14838 (N_14838,N_12783,N_13110);
nand U14839 (N_14839,N_12491,N_12819);
nand U14840 (N_14840,N_12678,N_13381);
or U14841 (N_14841,N_12965,N_12738);
nor U14842 (N_14842,N_13148,N_12647);
and U14843 (N_14843,N_13004,N_12831);
nor U14844 (N_14844,N_12085,N_12097);
xnor U14845 (N_14845,N_12396,N_12646);
nand U14846 (N_14846,N_12240,N_12305);
or U14847 (N_14847,N_13093,N_12192);
and U14848 (N_14848,N_13032,N_13211);
or U14849 (N_14849,N_13240,N_13312);
nand U14850 (N_14850,N_12700,N_12938);
nand U14851 (N_14851,N_13250,N_12155);
nand U14852 (N_14852,N_12067,N_12314);
nor U14853 (N_14853,N_12598,N_12953);
nor U14854 (N_14854,N_12000,N_13397);
nand U14855 (N_14855,N_12250,N_12589);
nor U14856 (N_14856,N_12052,N_12299);
nor U14857 (N_14857,N_12548,N_12044);
and U14858 (N_14858,N_13168,N_12922);
or U14859 (N_14859,N_12489,N_12214);
nand U14860 (N_14860,N_13106,N_12035);
nor U14861 (N_14861,N_13076,N_13150);
and U14862 (N_14862,N_12790,N_13488);
nor U14863 (N_14863,N_13493,N_12840);
nand U14864 (N_14864,N_13355,N_13359);
nor U14865 (N_14865,N_12394,N_13027);
nand U14866 (N_14866,N_13370,N_13207);
nand U14867 (N_14867,N_13477,N_12932);
nor U14868 (N_14868,N_12730,N_12838);
and U14869 (N_14869,N_12276,N_12976);
or U14870 (N_14870,N_12867,N_12077);
nor U14871 (N_14871,N_12309,N_13239);
and U14872 (N_14872,N_12696,N_12637);
or U14873 (N_14873,N_13426,N_13337);
or U14874 (N_14874,N_12746,N_13327);
xor U14875 (N_14875,N_12454,N_12859);
xnor U14876 (N_14876,N_12141,N_12320);
nand U14877 (N_14877,N_13377,N_12677);
nand U14878 (N_14878,N_12005,N_12410);
nand U14879 (N_14879,N_12924,N_13218);
nor U14880 (N_14880,N_12770,N_13161);
and U14881 (N_14881,N_12101,N_12186);
and U14882 (N_14882,N_12284,N_13120);
nand U14883 (N_14883,N_12471,N_12317);
or U14884 (N_14884,N_13278,N_12235);
nor U14885 (N_14885,N_12773,N_12598);
or U14886 (N_14886,N_12208,N_12212);
nand U14887 (N_14887,N_12742,N_12606);
and U14888 (N_14888,N_13146,N_13087);
nor U14889 (N_14889,N_12707,N_12069);
and U14890 (N_14890,N_13448,N_13191);
or U14891 (N_14891,N_12084,N_12852);
and U14892 (N_14892,N_13221,N_12503);
or U14893 (N_14893,N_13220,N_12659);
nand U14894 (N_14894,N_12703,N_12534);
nand U14895 (N_14895,N_13483,N_12680);
or U14896 (N_14896,N_13426,N_12021);
and U14897 (N_14897,N_13422,N_12055);
or U14898 (N_14898,N_13137,N_13000);
xor U14899 (N_14899,N_12582,N_12643);
or U14900 (N_14900,N_13409,N_12517);
xor U14901 (N_14901,N_12286,N_12615);
nand U14902 (N_14902,N_13097,N_12899);
nor U14903 (N_14903,N_13234,N_12480);
or U14904 (N_14904,N_12937,N_12936);
nor U14905 (N_14905,N_13416,N_12597);
nor U14906 (N_14906,N_12822,N_12517);
nor U14907 (N_14907,N_12876,N_13180);
xor U14908 (N_14908,N_12722,N_12605);
nand U14909 (N_14909,N_12388,N_13241);
nand U14910 (N_14910,N_12900,N_12033);
and U14911 (N_14911,N_13356,N_12351);
nand U14912 (N_14912,N_12011,N_12225);
or U14913 (N_14913,N_12016,N_12727);
or U14914 (N_14914,N_12081,N_12801);
nand U14915 (N_14915,N_12707,N_12213);
and U14916 (N_14916,N_12207,N_13028);
and U14917 (N_14917,N_12508,N_13417);
and U14918 (N_14918,N_12076,N_12924);
or U14919 (N_14919,N_12254,N_13463);
or U14920 (N_14920,N_12663,N_13302);
nand U14921 (N_14921,N_13300,N_13233);
and U14922 (N_14922,N_13054,N_12380);
nor U14923 (N_14923,N_12712,N_13419);
or U14924 (N_14924,N_12977,N_12511);
and U14925 (N_14925,N_13350,N_12072);
and U14926 (N_14926,N_12779,N_12281);
nor U14927 (N_14927,N_13163,N_12040);
or U14928 (N_14928,N_12358,N_12682);
or U14929 (N_14929,N_13380,N_12934);
or U14930 (N_14930,N_13043,N_13187);
nand U14931 (N_14931,N_12774,N_12521);
nand U14932 (N_14932,N_13174,N_12261);
and U14933 (N_14933,N_13224,N_12583);
nand U14934 (N_14934,N_13381,N_12487);
or U14935 (N_14935,N_12236,N_13391);
xor U14936 (N_14936,N_12153,N_13002);
xor U14937 (N_14937,N_12540,N_12321);
nor U14938 (N_14938,N_13444,N_13360);
nand U14939 (N_14939,N_12444,N_12331);
and U14940 (N_14940,N_12558,N_12631);
nand U14941 (N_14941,N_12040,N_13194);
nand U14942 (N_14942,N_12964,N_13168);
nand U14943 (N_14943,N_13491,N_12699);
and U14944 (N_14944,N_12938,N_12730);
and U14945 (N_14945,N_12391,N_12615);
nand U14946 (N_14946,N_12910,N_12554);
nor U14947 (N_14947,N_12348,N_13151);
nand U14948 (N_14948,N_12962,N_12676);
nor U14949 (N_14949,N_13399,N_13439);
nand U14950 (N_14950,N_12509,N_13329);
or U14951 (N_14951,N_13480,N_12683);
nor U14952 (N_14952,N_13274,N_12775);
or U14953 (N_14953,N_12359,N_13312);
and U14954 (N_14954,N_13069,N_13337);
or U14955 (N_14955,N_12634,N_12604);
nand U14956 (N_14956,N_12591,N_12225);
and U14957 (N_14957,N_12630,N_12699);
nor U14958 (N_14958,N_13009,N_13307);
xor U14959 (N_14959,N_12928,N_13440);
or U14960 (N_14960,N_12517,N_12273);
or U14961 (N_14961,N_13187,N_12088);
or U14962 (N_14962,N_12741,N_12716);
nand U14963 (N_14963,N_12627,N_12155);
nand U14964 (N_14964,N_12096,N_12713);
nand U14965 (N_14965,N_12939,N_12303);
nor U14966 (N_14966,N_13435,N_12015);
and U14967 (N_14967,N_13137,N_12753);
nand U14968 (N_14968,N_13395,N_12453);
nand U14969 (N_14969,N_13202,N_12038);
or U14970 (N_14970,N_12443,N_13050);
or U14971 (N_14971,N_12389,N_12073);
and U14972 (N_14972,N_13157,N_12497);
nand U14973 (N_14973,N_12702,N_13280);
nand U14974 (N_14974,N_12730,N_13223);
nand U14975 (N_14975,N_12547,N_12886);
or U14976 (N_14976,N_12732,N_13378);
or U14977 (N_14977,N_12591,N_12577);
nand U14978 (N_14978,N_13103,N_12006);
and U14979 (N_14979,N_12873,N_12955);
nand U14980 (N_14980,N_12693,N_13493);
nand U14981 (N_14981,N_12296,N_12308);
nand U14982 (N_14982,N_12764,N_13088);
or U14983 (N_14983,N_12297,N_12407);
nor U14984 (N_14984,N_12167,N_12299);
or U14985 (N_14985,N_12440,N_13071);
and U14986 (N_14986,N_12379,N_12312);
xor U14987 (N_14987,N_12405,N_12369);
and U14988 (N_14988,N_13397,N_13347);
xnor U14989 (N_14989,N_12890,N_12177);
nor U14990 (N_14990,N_12135,N_12367);
nor U14991 (N_14991,N_12809,N_13263);
xor U14992 (N_14992,N_13415,N_12053);
or U14993 (N_14993,N_12459,N_13021);
nor U14994 (N_14994,N_12764,N_12112);
and U14995 (N_14995,N_13343,N_12486);
and U14996 (N_14996,N_13035,N_12813);
nand U14997 (N_14997,N_12591,N_12774);
and U14998 (N_14998,N_12662,N_12043);
nor U14999 (N_14999,N_12288,N_12825);
or UO_0 (O_0,N_14825,N_14178);
and UO_1 (O_1,N_14498,N_13829);
nand UO_2 (O_2,N_14628,N_14126);
and UO_3 (O_3,N_13718,N_13586);
nand UO_4 (O_4,N_13523,N_13562);
nor UO_5 (O_5,N_13871,N_14461);
or UO_6 (O_6,N_13954,N_14381);
nor UO_7 (O_7,N_14151,N_14236);
nand UO_8 (O_8,N_13765,N_13982);
nor UO_9 (O_9,N_14692,N_14273);
xnor UO_10 (O_10,N_14726,N_14690);
nor UO_11 (O_11,N_13889,N_14362);
xor UO_12 (O_12,N_14788,N_13722);
and UO_13 (O_13,N_14086,N_13866);
or UO_14 (O_14,N_13703,N_14958);
and UO_15 (O_15,N_13815,N_14587);
xor UO_16 (O_16,N_14199,N_14089);
or UO_17 (O_17,N_13814,N_14987);
or UO_18 (O_18,N_14931,N_14801);
nand UO_19 (O_19,N_14096,N_14002);
or UO_20 (O_20,N_14186,N_14053);
xor UO_21 (O_21,N_13976,N_13846);
xnor UO_22 (O_22,N_14838,N_14757);
or UO_23 (O_23,N_14889,N_13971);
or UO_24 (O_24,N_14897,N_13755);
or UO_25 (O_25,N_14261,N_14643);
xnor UO_26 (O_26,N_14839,N_13842);
nor UO_27 (O_27,N_13538,N_13816);
or UO_28 (O_28,N_14067,N_14539);
or UO_29 (O_29,N_14443,N_14976);
nor UO_30 (O_30,N_13974,N_14828);
nand UO_31 (O_31,N_14548,N_13885);
nor UO_32 (O_32,N_14970,N_14909);
or UO_33 (O_33,N_14581,N_14729);
or UO_34 (O_34,N_14100,N_14473);
xnor UO_35 (O_35,N_14625,N_14365);
or UO_36 (O_36,N_14398,N_14413);
or UO_37 (O_37,N_13770,N_14046);
nand UO_38 (O_38,N_14194,N_14162);
nand UO_39 (O_39,N_14906,N_14167);
and UO_40 (O_40,N_14589,N_13942);
and UO_41 (O_41,N_13507,N_14940);
nand UO_42 (O_42,N_14934,N_13744);
nand UO_43 (O_43,N_14749,N_13978);
and UO_44 (O_44,N_14588,N_14693);
and UO_45 (O_45,N_14289,N_14016);
nand UO_46 (O_46,N_14630,N_13513);
nand UO_47 (O_47,N_14375,N_13527);
nand UO_48 (O_48,N_14139,N_13572);
xor UO_49 (O_49,N_14437,N_13831);
and UO_50 (O_50,N_14451,N_13693);
nand UO_51 (O_51,N_14545,N_14569);
nand UO_52 (O_52,N_14209,N_14306);
nand UO_53 (O_53,N_13966,N_14620);
nand UO_54 (O_54,N_14425,N_13964);
or UO_55 (O_55,N_14579,N_14416);
nand UO_56 (O_56,N_13967,N_13568);
nor UO_57 (O_57,N_14773,N_13707);
or UO_58 (O_58,N_13930,N_14813);
and UO_59 (O_59,N_13729,N_14611);
and UO_60 (O_60,N_14562,N_13856);
nor UO_61 (O_61,N_14383,N_14395);
nand UO_62 (O_62,N_13570,N_14925);
or UO_63 (O_63,N_14242,N_13702);
or UO_64 (O_64,N_13806,N_14501);
or UO_65 (O_65,N_14856,N_14103);
nand UO_66 (O_66,N_13780,N_14846);
and UO_67 (O_67,N_13725,N_14857);
and UO_68 (O_68,N_14850,N_14021);
or UO_69 (O_69,N_13953,N_14268);
nand UO_70 (O_70,N_14922,N_14304);
nor UO_71 (O_71,N_14699,N_13809);
and UO_72 (O_72,N_13767,N_14893);
nor UO_73 (O_73,N_14663,N_14927);
nand UO_74 (O_74,N_14314,N_14979);
and UO_75 (O_75,N_13848,N_13960);
xor UO_76 (O_76,N_14344,N_14800);
nand UO_77 (O_77,N_13514,N_14576);
xnor UO_78 (O_78,N_14883,N_14397);
nor UO_79 (O_79,N_14707,N_13731);
nor UO_80 (O_80,N_14082,N_14658);
nand UO_81 (O_81,N_14332,N_14034);
xor UO_82 (O_82,N_14718,N_14446);
nand UO_83 (O_83,N_14253,N_14973);
nor UO_84 (O_84,N_14674,N_13593);
and UO_85 (O_85,N_14227,N_13641);
nor UO_86 (O_86,N_14706,N_14324);
and UO_87 (O_87,N_14269,N_14168);
nand UO_88 (O_88,N_14563,N_13617);
xnor UO_89 (O_89,N_14632,N_14792);
nand UO_90 (O_90,N_13534,N_14346);
or UO_91 (O_91,N_13697,N_13608);
nor UO_92 (O_92,N_14008,N_14966);
nand UO_93 (O_93,N_14983,N_14121);
nor UO_94 (O_94,N_14391,N_14213);
xor UO_95 (O_95,N_13726,N_14335);
nor UO_96 (O_96,N_14438,N_14617);
and UO_97 (O_97,N_14600,N_14226);
xnor UO_98 (O_98,N_14784,N_13577);
nor UO_99 (O_99,N_14502,N_14240);
xor UO_100 (O_100,N_14762,N_14219);
nor UO_101 (O_101,N_13841,N_14482);
and UO_102 (O_102,N_14255,N_14481);
and UO_103 (O_103,N_13630,N_14170);
nor UO_104 (O_104,N_13656,N_14001);
and UO_105 (O_105,N_13992,N_13713);
or UO_106 (O_106,N_13798,N_14516);
nor UO_107 (O_107,N_14185,N_13680);
and UO_108 (O_108,N_14894,N_14531);
xnor UO_109 (O_109,N_14766,N_14975);
and UO_110 (O_110,N_13502,N_14929);
and UO_111 (O_111,N_13640,N_14373);
or UO_112 (O_112,N_14330,N_14159);
nor UO_113 (O_113,N_14254,N_14315);
or UO_114 (O_114,N_14129,N_14452);
nand UO_115 (O_115,N_13631,N_14566);
and UO_116 (O_116,N_14519,N_13837);
and UO_117 (O_117,N_14791,N_13855);
xor UO_118 (O_118,N_14812,N_13988);
nand UO_119 (O_119,N_13921,N_14187);
nor UO_120 (O_120,N_14327,N_14147);
or UO_121 (O_121,N_14740,N_13579);
or UO_122 (O_122,N_14285,N_14527);
and UO_123 (O_123,N_14688,N_13875);
xor UO_124 (O_124,N_14951,N_14442);
or UO_125 (O_125,N_13677,N_14877);
nor UO_126 (O_126,N_13795,N_13532);
or UO_127 (O_127,N_14528,N_14997);
nor UO_128 (O_128,N_14284,N_13894);
nand UO_129 (O_129,N_14043,N_14577);
and UO_130 (O_130,N_14274,N_14241);
or UO_131 (O_131,N_13606,N_13673);
nand UO_132 (O_132,N_14650,N_14945);
or UO_133 (O_133,N_14013,N_13773);
nand UO_134 (O_134,N_13510,N_14673);
nor UO_135 (O_135,N_14025,N_13900);
nand UO_136 (O_136,N_13588,N_13610);
and UO_137 (O_137,N_13892,N_13627);
xor UO_138 (O_138,N_13936,N_14294);
nor UO_139 (O_139,N_14491,N_14939);
nand UO_140 (O_140,N_14305,N_14736);
or UO_141 (O_141,N_13754,N_14064);
xnor UO_142 (O_142,N_13763,N_13832);
nor UO_143 (O_143,N_14078,N_14610);
nand UO_144 (O_144,N_14680,N_14465);
nor UO_145 (O_145,N_14052,N_13556);
nor UO_146 (O_146,N_14637,N_13671);
nor UO_147 (O_147,N_14212,N_14503);
nand UO_148 (O_148,N_14861,N_14799);
nand UO_149 (O_149,N_14320,N_14286);
nand UO_150 (O_150,N_13989,N_13574);
or UO_151 (O_151,N_14120,N_14638);
nand UO_152 (O_152,N_13857,N_14145);
nor UO_153 (O_153,N_13602,N_14480);
nor UO_154 (O_154,N_14768,N_14629);
nor UO_155 (O_155,N_13839,N_13565);
xnor UO_156 (O_156,N_13817,N_13666);
or UO_157 (O_157,N_14295,N_13660);
nand UO_158 (O_158,N_14095,N_14288);
nand UO_159 (O_159,N_13541,N_14770);
and UO_160 (O_160,N_13724,N_14148);
nor UO_161 (O_161,N_13528,N_14192);
or UO_162 (O_162,N_14822,N_13632);
or UO_163 (O_163,N_14733,N_14439);
and UO_164 (O_164,N_13694,N_14155);
xor UO_165 (O_165,N_14250,N_14180);
xor UO_166 (O_166,N_13653,N_13547);
or UO_167 (O_167,N_13977,N_13849);
and UO_168 (O_168,N_14623,N_14598);
and UO_169 (O_169,N_14028,N_14963);
and UO_170 (O_170,N_14796,N_14456);
nor UO_171 (O_171,N_14664,N_14419);
xnor UO_172 (O_172,N_13927,N_14660);
or UO_173 (O_173,N_14018,N_13776);
or UO_174 (O_174,N_14105,N_14328);
nor UO_175 (O_175,N_13799,N_14805);
nor UO_176 (O_176,N_14470,N_13564);
and UO_177 (O_177,N_14485,N_14634);
and UO_178 (O_178,N_14666,N_14550);
nand UO_179 (O_179,N_13860,N_13730);
xor UO_180 (O_180,N_14984,N_14942);
and UO_181 (O_181,N_14303,N_14318);
nor UO_182 (O_182,N_14841,N_14875);
and UO_183 (O_183,N_14696,N_14441);
and UO_184 (O_184,N_14127,N_14207);
or UO_185 (O_185,N_14190,N_14322);
or UO_186 (O_186,N_13880,N_14952);
nand UO_187 (O_187,N_14845,N_14410);
nor UO_188 (O_188,N_13874,N_14203);
nand UO_189 (O_189,N_14154,N_13929);
and UO_190 (O_190,N_14636,N_13833);
nand UO_191 (O_191,N_14440,N_13786);
xor UO_192 (O_192,N_14427,N_14272);
xor UO_193 (O_193,N_14532,N_14293);
or UO_194 (O_194,N_13994,N_13681);
or UO_195 (O_195,N_13840,N_13634);
and UO_196 (O_196,N_14672,N_13511);
nand UO_197 (O_197,N_14949,N_13609);
nand UO_198 (O_198,N_13990,N_13879);
nor UO_199 (O_199,N_14866,N_13700);
and UO_200 (O_200,N_14031,N_14826);
nand UO_201 (O_201,N_13947,N_13699);
or UO_202 (O_202,N_14281,N_13530);
xor UO_203 (O_203,N_13581,N_14251);
nor UO_204 (O_204,N_13872,N_14038);
or UO_205 (O_205,N_13659,N_13811);
nor UO_206 (O_206,N_14323,N_14267);
and UO_207 (O_207,N_13993,N_14353);
xnor UO_208 (O_208,N_14510,N_14153);
nand UO_209 (O_209,N_13813,N_14591);
or UO_210 (O_210,N_13720,N_14795);
nor UO_211 (O_211,N_13985,N_14526);
and UO_212 (O_212,N_13529,N_14535);
nand UO_213 (O_213,N_13526,N_14118);
nor UO_214 (O_214,N_13648,N_13756);
and UO_215 (O_215,N_14171,N_14978);
and UO_216 (O_216,N_14947,N_13774);
nor UO_217 (O_217,N_14309,N_14552);
or UO_218 (O_218,N_14087,N_14898);
nand UO_219 (O_219,N_14357,N_13844);
nand UO_220 (O_220,N_14197,N_13850);
and UO_221 (O_221,N_14886,N_14640);
and UO_222 (O_222,N_14202,N_14758);
or UO_223 (O_223,N_14543,N_14379);
nand UO_224 (O_224,N_14032,N_14435);
nor UO_225 (O_225,N_13934,N_14928);
nor UO_226 (O_226,N_13711,N_14659);
or UO_227 (O_227,N_14243,N_14752);
or UO_228 (O_228,N_13959,N_14950);
nand UO_229 (O_229,N_13682,N_14326);
and UO_230 (O_230,N_14702,N_14338);
or UO_231 (O_231,N_14734,N_14776);
and UO_232 (O_232,N_14819,N_13536);
and UO_233 (O_233,N_14024,N_14106);
and UO_234 (O_234,N_14406,N_14989);
xnor UO_235 (O_235,N_14135,N_14910);
and UO_236 (O_236,N_14725,N_14492);
nand UO_237 (O_237,N_14551,N_14609);
nand UO_238 (O_238,N_14084,N_14604);
and UO_239 (O_239,N_13594,N_13549);
nand UO_240 (O_240,N_14206,N_14872);
and UO_241 (O_241,N_14142,N_14399);
nor UO_242 (O_242,N_14648,N_14390);
and UO_243 (O_243,N_13623,N_13836);
and UO_244 (O_244,N_13843,N_14962);
xor UO_245 (O_245,N_14712,N_14351);
and UO_246 (O_246,N_14654,N_14280);
xnor UO_247 (O_247,N_14401,N_14723);
nand UO_248 (O_248,N_14062,N_14041);
or UO_249 (O_249,N_14027,N_14436);
or UO_250 (O_250,N_14149,N_14050);
and UO_251 (O_251,N_14618,N_13787);
and UO_252 (O_252,N_13591,N_14635);
nor UO_253 (O_253,N_14182,N_14123);
nor UO_254 (O_254,N_13919,N_14574);
and UO_255 (O_255,N_14737,N_14714);
xor UO_256 (O_256,N_14361,N_14081);
and UO_257 (O_257,N_14376,N_14564);
xnor UO_258 (O_258,N_13638,N_13995);
nor UO_259 (O_259,N_14597,N_14593);
nand UO_260 (O_260,N_13950,N_14065);
nor UO_261 (O_261,N_14426,N_14895);
or UO_262 (O_262,N_13539,N_13557);
or UO_263 (O_263,N_14161,N_14512);
nor UO_264 (O_264,N_13788,N_14720);
nand UO_265 (O_265,N_14384,N_13597);
and UO_266 (O_266,N_14936,N_14964);
nand UO_267 (O_267,N_14460,N_14787);
xor UO_268 (O_268,N_14467,N_14665);
or UO_269 (O_269,N_14785,N_14003);
nor UO_270 (O_270,N_14462,N_13612);
nand UO_271 (O_271,N_13823,N_14504);
or UO_272 (O_272,N_14205,N_14751);
nor UO_273 (O_273,N_14697,N_13563);
or UO_274 (O_274,N_13975,N_14073);
and UO_275 (O_275,N_13757,N_14036);
nand UO_276 (O_276,N_14445,N_13521);
nand UO_277 (O_277,N_14468,N_14125);
xnor UO_278 (O_278,N_14724,N_13599);
xor UO_279 (O_279,N_14624,N_13624);
nor UO_280 (O_280,N_14370,N_13698);
nand UO_281 (O_281,N_13891,N_14809);
and UO_282 (O_282,N_14235,N_14099);
and UO_283 (O_283,N_14402,N_14112);
nand UO_284 (O_284,N_13550,N_14420);
and UO_285 (O_285,N_14619,N_13592);
and UO_286 (O_286,N_14108,N_14806);
and UO_287 (O_287,N_14228,N_14358);
nor UO_288 (O_288,N_14415,N_14642);
or UO_289 (O_289,N_13688,N_13812);
and UO_290 (O_290,N_13519,N_14133);
and UO_291 (O_291,N_13654,N_14216);
nand UO_292 (O_292,N_14360,N_14484);
xor UO_293 (O_293,N_13958,N_14891);
nor UO_294 (O_294,N_13636,N_14386);
nor UO_295 (O_295,N_13887,N_13674);
and UO_296 (O_296,N_14511,N_13893);
nor UO_297 (O_297,N_14308,N_13769);
xnor UO_298 (O_298,N_13969,N_13537);
or UO_299 (O_299,N_14310,N_13968);
and UO_300 (O_300,N_14810,N_13758);
nand UO_301 (O_301,N_14911,N_14888);
or UO_302 (O_302,N_14458,N_14592);
and UO_303 (O_303,N_14882,N_13973);
and UO_304 (O_304,N_14578,N_14144);
xnor UO_305 (O_305,N_14522,N_14546);
nand UO_306 (O_306,N_13999,N_14960);
nor UO_307 (O_307,N_13945,N_13622);
nand UO_308 (O_308,N_13895,N_13793);
xor UO_309 (O_309,N_14264,N_13943);
and UO_310 (O_310,N_13667,N_14899);
nand UO_311 (O_311,N_14716,N_14290);
and UO_312 (O_312,N_14671,N_13779);
or UO_313 (O_313,N_14183,N_14781);
nand UO_314 (O_314,N_14775,N_13917);
xor UO_315 (O_315,N_13932,N_13542);
and UO_316 (O_316,N_13664,N_14641);
or UO_317 (O_317,N_14450,N_13687);
and UO_318 (O_318,N_13749,N_13922);
nor UO_319 (O_319,N_13629,N_13512);
and UO_320 (O_320,N_14655,N_14488);
nand UO_321 (O_321,N_14074,N_14890);
nand UO_322 (O_322,N_14124,N_14292);
nand UO_323 (O_323,N_14573,N_14747);
and UO_324 (O_324,N_13672,N_14953);
nand UO_325 (O_325,N_14647,N_13984);
nor UO_326 (O_326,N_14605,N_14382);
nand UO_327 (O_327,N_13643,N_14990);
or UO_328 (O_328,N_14824,N_14019);
and UO_329 (O_329,N_14783,N_14266);
or UO_330 (O_330,N_14933,N_13826);
nand UO_331 (O_331,N_14150,N_13633);
nand UO_332 (O_332,N_13979,N_14196);
and UO_333 (O_333,N_13981,N_14333);
or UO_334 (O_334,N_14818,N_14163);
and UO_335 (O_335,N_13575,N_14683);
or UO_336 (O_336,N_13998,N_13918);
and UO_337 (O_337,N_14907,N_14372);
nor UO_338 (O_338,N_14862,N_14797);
or UO_339 (O_339,N_14107,N_14364);
or UO_340 (O_340,N_14859,N_14896);
and UO_341 (O_341,N_14471,N_14248);
xnor UO_342 (O_342,N_14014,N_13571);
nor UO_343 (O_343,N_14521,N_14307);
nor UO_344 (O_344,N_14012,N_14541);
or UO_345 (O_345,N_14529,N_13928);
and UO_346 (O_346,N_14430,N_13752);
nand UO_347 (O_347,N_13646,N_14919);
nand UO_348 (O_348,N_14662,N_14276);
nor UO_349 (O_349,N_13748,N_13775);
and UO_350 (O_350,N_13783,N_13583);
and UO_351 (O_351,N_13584,N_14408);
nand UO_352 (O_352,N_13506,N_14767);
and UO_353 (O_353,N_14750,N_14614);
or UO_354 (O_354,N_13941,N_14601);
nand UO_355 (O_355,N_14902,N_13870);
and UO_356 (O_356,N_14049,N_14411);
and UO_357 (O_357,N_13820,N_13873);
nand UO_358 (O_358,N_14653,N_14667);
nor UO_359 (O_359,N_13509,N_13746);
and UO_360 (O_360,N_13791,N_14299);
or UO_361 (O_361,N_14432,N_13690);
nand UO_362 (O_362,N_14230,N_14472);
nor UO_363 (O_363,N_13914,N_14011);
nand UO_364 (O_364,N_14130,N_14422);
and UO_365 (O_365,N_13605,N_14137);
and UO_366 (O_366,N_14853,N_14188);
and UO_367 (O_367,N_13926,N_14090);
or UO_368 (O_368,N_14337,N_14739);
nand UO_369 (O_369,N_13778,N_14218);
or UO_370 (O_370,N_14469,N_13937);
nand UO_371 (O_371,N_14677,N_14756);
nor UO_372 (O_372,N_13951,N_13576);
xor UO_373 (O_373,N_14753,N_14101);
nand UO_374 (O_374,N_14514,N_13626);
or UO_375 (O_375,N_14238,N_13695);
xnor UO_376 (O_376,N_14110,N_14967);
nor UO_377 (O_377,N_14802,N_14487);
nand UO_378 (O_378,N_14069,N_13683);
and UO_379 (O_379,N_13578,N_14463);
and UO_380 (O_380,N_13803,N_14263);
nand UO_381 (O_381,N_13500,N_13540);
nor UO_382 (O_382,N_13601,N_13807);
nor UO_383 (O_383,N_13533,N_13613);
xnor UO_384 (O_384,N_14369,N_13589);
nand UO_385 (O_385,N_14547,N_14079);
nor UO_386 (O_386,N_13719,N_14160);
and UO_387 (O_387,N_14444,N_14873);
nor UO_388 (O_388,N_13717,N_14232);
nand UO_389 (O_389,N_14394,N_14279);
or UO_390 (O_390,N_14705,N_13721);
nor UO_391 (O_391,N_13535,N_14039);
or UO_392 (O_392,N_14827,N_14955);
nor UO_393 (O_393,N_13804,N_13708);
or UO_394 (O_394,N_14275,N_14076);
nor UO_395 (O_395,N_14874,N_14136);
nand UO_396 (O_396,N_14257,N_14836);
and UO_397 (O_397,N_13789,N_14215);
or UO_398 (O_398,N_13925,N_14981);
or UO_399 (O_399,N_13531,N_14954);
or UO_400 (O_400,N_14143,N_14347);
nand UO_401 (O_401,N_13585,N_13706);
or UO_402 (O_402,N_14559,N_14865);
or UO_403 (O_403,N_14881,N_14044);
and UO_404 (O_404,N_13781,N_14917);
nand UO_405 (O_405,N_14520,N_14525);
nor UO_406 (O_406,N_13516,N_14026);
xor UO_407 (O_407,N_14533,N_14237);
nand UO_408 (O_408,N_14980,N_13980);
and UO_409 (O_409,N_14208,N_14695);
nand UO_410 (O_410,N_14412,N_14172);
and UO_411 (O_411,N_14554,N_13940);
xnor UO_412 (O_412,N_14138,N_13883);
nor UO_413 (O_413,N_14682,N_14530);
nand UO_414 (O_414,N_13662,N_13676);
or UO_415 (O_415,N_14270,N_14317);
and UO_416 (O_416,N_14908,N_13948);
and UO_417 (O_417,N_13761,N_13712);
nand UO_418 (O_418,N_13794,N_14374);
and UO_419 (O_419,N_14721,N_14176);
nand UO_420 (O_420,N_13963,N_14583);
or UO_421 (O_421,N_13741,N_14870);
xnor UO_422 (O_422,N_13735,N_14249);
nor UO_423 (O_423,N_14985,N_14259);
and UO_424 (O_424,N_14603,N_14098);
or UO_425 (O_425,N_13905,N_14884);
nor UO_426 (O_426,N_14177,N_13961);
nor UO_427 (O_427,N_14301,N_13675);
or UO_428 (O_428,N_14536,N_13825);
nor UO_429 (O_429,N_13637,N_14234);
nand UO_430 (O_430,N_13760,N_14345);
or UO_431 (O_431,N_14004,N_13595);
nor UO_432 (O_432,N_14164,N_14916);
or UO_433 (O_433,N_14823,N_14174);
nor UO_434 (O_434,N_14010,N_14992);
nand UO_435 (O_435,N_13603,N_14246);
nor UO_436 (O_436,N_14080,N_14282);
nand UO_437 (O_437,N_14509,N_14061);
nand UO_438 (O_438,N_14311,N_14479);
nand UO_439 (O_439,N_14007,N_13907);
or UO_440 (O_440,N_14225,N_14959);
xor UO_441 (O_441,N_14392,N_14670);
nand UO_442 (O_442,N_13649,N_13669);
or UO_443 (O_443,N_14029,N_14921);
and UO_444 (O_444,N_13915,N_13560);
nor UO_445 (O_445,N_14694,N_14602);
nor UO_446 (O_446,N_14972,N_14849);
nand UO_447 (O_447,N_14719,N_14811);
or UO_448 (O_448,N_14513,N_14222);
nor UO_449 (O_449,N_14599,N_14912);
or UO_450 (O_450,N_14804,N_14091);
xnor UO_451 (O_451,N_14855,N_14109);
or UO_452 (O_452,N_14341,N_14063);
and UO_453 (O_453,N_13518,N_14568);
nand UO_454 (O_454,N_14941,N_14005);
nor UO_455 (O_455,N_14200,N_14760);
nand UO_456 (O_456,N_14405,N_13580);
and UO_457 (O_457,N_13614,N_14497);
xor UO_458 (O_458,N_14956,N_14193);
nand UO_459 (O_459,N_13566,N_14146);
and UO_460 (O_460,N_13504,N_13802);
nand UO_461 (O_461,N_14239,N_14047);
nor UO_462 (O_462,N_14017,N_14937);
nand UO_463 (O_463,N_14378,N_14821);
nor UO_464 (O_464,N_14296,N_13587);
and UO_465 (O_465,N_14418,N_13670);
xor UO_466 (O_466,N_14639,N_13986);
nor UO_467 (O_467,N_14717,N_14119);
or UO_468 (O_468,N_14085,N_14627);
nor UO_469 (O_469,N_14020,N_13658);
and UO_470 (O_470,N_14913,N_14999);
nor UO_471 (O_471,N_14340,N_14500);
nand UO_472 (O_472,N_13827,N_14582);
and UO_473 (O_473,N_14901,N_14777);
nor UO_474 (O_474,N_14507,N_14924);
nor UO_475 (O_475,N_14343,N_14595);
or UO_476 (O_476,N_14971,N_14794);
nor UO_477 (O_477,N_13596,N_14957);
nand UO_478 (O_478,N_14741,N_14542);
or UO_479 (O_479,N_13704,N_13663);
nor UO_480 (O_480,N_14229,N_14414);
nor UO_481 (O_481,N_14555,N_14231);
xor UO_482 (O_482,N_13818,N_14388);
nor UO_483 (O_483,N_14403,N_13805);
or UO_484 (O_484,N_13935,N_14656);
xor UO_485 (O_485,N_14769,N_13904);
xnor UO_486 (O_486,N_13909,N_14968);
nand UO_487 (O_487,N_14868,N_13896);
or UO_488 (O_488,N_14015,N_14843);
and UO_489 (O_489,N_13946,N_14455);
and UO_490 (O_490,N_13657,N_14389);
nor UO_491 (O_491,N_14515,N_13692);
nand UO_492 (O_492,N_13644,N_14336);
or UO_493 (O_493,N_14057,N_14359);
nor UO_494 (O_494,N_14835,N_14490);
and UO_495 (O_495,N_14657,N_13972);
or UO_496 (O_496,N_14860,N_14914);
and UO_497 (O_497,N_13916,N_14903);
nor UO_498 (O_498,N_14068,N_14042);
and UO_499 (O_499,N_14499,N_13736);
nand UO_500 (O_500,N_13931,N_14974);
nor UO_501 (O_501,N_14366,N_14265);
nand UO_502 (O_502,N_14745,N_14128);
and UO_503 (O_503,N_14534,N_14058);
and UO_504 (O_504,N_13955,N_14549);
nand UO_505 (O_505,N_14056,N_14092);
or UO_506 (O_506,N_14687,N_13600);
and UO_507 (O_507,N_14429,N_14223);
nor UO_508 (O_508,N_14887,N_14506);
nand UO_509 (O_509,N_13742,N_14204);
nor UO_510 (O_510,N_13505,N_14363);
and UO_511 (O_511,N_13508,N_13835);
nor UO_512 (O_512,N_14173,N_14932);
nor UO_513 (O_513,N_13555,N_14114);
nor UO_514 (O_514,N_13517,N_13854);
xnor UO_515 (O_515,N_14115,N_14586);
or UO_516 (O_516,N_13903,N_14400);
xor UO_517 (O_517,N_14851,N_14453);
or UO_518 (O_518,N_13616,N_14368);
or UO_519 (O_519,N_14478,N_14575);
nand UO_520 (O_520,N_14508,N_14466);
and UO_521 (O_521,N_14840,N_14616);
nand UO_522 (O_522,N_14876,N_14037);
and UO_523 (O_523,N_14691,N_13908);
and UO_524 (O_524,N_13970,N_14764);
or UO_525 (O_525,N_14915,N_14704);
nand UO_526 (O_526,N_13762,N_14312);
nor UO_527 (O_527,N_13867,N_14496);
and UO_528 (O_528,N_13590,N_14580);
or UO_529 (O_529,N_13598,N_14111);
or UO_530 (O_530,N_14943,N_14329);
and UO_531 (O_531,N_14748,N_14354);
nor UO_532 (O_532,N_14077,N_14848);
nor UO_533 (O_533,N_13544,N_14867);
xor UO_534 (O_534,N_14698,N_14998);
and UO_535 (O_535,N_13714,N_13525);
nand UO_536 (O_536,N_14961,N_13750);
and UO_537 (O_537,N_14102,N_14083);
or UO_538 (O_538,N_13920,N_13877);
nand UO_539 (O_539,N_14104,N_13777);
or UO_540 (O_540,N_14048,N_14476);
xor UO_541 (O_541,N_14169,N_14367);
nor UO_542 (O_542,N_13652,N_13524);
and UO_543 (O_543,N_14755,N_14433);
nand UO_544 (O_544,N_14540,N_14612);
and UO_545 (O_545,N_13861,N_14727);
nor UO_546 (O_546,N_14715,N_14730);
nor UO_547 (O_547,N_14701,N_14782);
nor UO_548 (O_548,N_13738,N_14878);
and UO_549 (O_549,N_13751,N_14560);
and UO_550 (O_550,N_14558,N_14256);
nor UO_551 (O_551,N_14262,N_13766);
nand UO_552 (O_552,N_13834,N_14986);
or UO_553 (O_553,N_13933,N_14571);
or UO_554 (O_554,N_14651,N_14728);
and UO_555 (O_555,N_14457,N_14505);
nor UO_556 (O_556,N_14387,N_14675);
nand UO_557 (O_557,N_14608,N_14596);
and UO_558 (O_558,N_14926,N_14224);
or UO_559 (O_559,N_14407,N_14594);
xnor UO_560 (O_560,N_14424,N_14652);
and UO_561 (O_561,N_14352,N_14615);
or UO_562 (O_562,N_14217,N_14517);
nor UO_563 (O_563,N_14621,N_13902);
or UO_564 (O_564,N_14313,N_13882);
or UO_565 (O_565,N_13987,N_14761);
and UO_566 (O_566,N_13620,N_14556);
xnor UO_567 (O_567,N_14054,N_14731);
or UO_568 (O_568,N_14871,N_14244);
nor UO_569 (O_569,N_14117,N_13685);
or UO_570 (O_570,N_14334,N_13647);
or UO_571 (O_571,N_14661,N_14030);
or UO_572 (O_572,N_14071,N_14464);
nand UO_573 (O_573,N_14743,N_13790);
nor UO_574 (O_574,N_14132,N_14996);
and UO_575 (O_575,N_13701,N_14165);
or UO_576 (O_576,N_13991,N_14759);
or UO_577 (O_577,N_13678,N_14214);
or UO_578 (O_578,N_14681,N_14900);
nor UO_579 (O_579,N_14475,N_14994);
nor UO_580 (O_580,N_13665,N_14572);
nand UO_581 (O_581,N_14220,N_14093);
xor UO_582 (O_582,N_14565,N_13628);
and UO_583 (O_583,N_14544,N_14350);
and UO_584 (O_584,N_14287,N_14316);
nor UO_585 (O_585,N_13551,N_14072);
nor UO_586 (O_586,N_13661,N_14918);
nand UO_587 (O_587,N_14700,N_14669);
xor UO_588 (O_588,N_14709,N_14584);
and UO_589 (O_589,N_14746,N_13567);
nor UO_590 (O_590,N_14993,N_14489);
nand UO_591 (O_591,N_14302,N_14339);
and UO_592 (O_592,N_13983,N_14247);
and UO_593 (O_593,N_13822,N_14880);
nor UO_594 (O_594,N_13604,N_14676);
nor UO_595 (O_595,N_13864,N_13642);
nor UO_596 (O_596,N_14348,N_13621);
and UO_597 (O_597,N_14210,N_14803);
or UO_598 (O_598,N_13619,N_14935);
or UO_599 (O_599,N_14157,N_14885);
or UO_600 (O_600,N_14965,N_13553);
or UO_601 (O_601,N_14991,N_13747);
nor UO_602 (O_602,N_14837,N_14454);
and UO_603 (O_603,N_13944,N_14494);
nand UO_604 (O_604,N_13819,N_14607);
nor UO_605 (O_605,N_14606,N_13764);
nand UO_606 (O_606,N_14613,N_14537);
nor UO_607 (O_607,N_14070,N_14495);
nand UO_608 (O_608,N_13522,N_14181);
nor UO_609 (O_609,N_13759,N_13554);
nor UO_610 (O_610,N_14847,N_14832);
nand UO_611 (O_611,N_14703,N_13582);
nor UO_612 (O_612,N_14946,N_13847);
nor UO_613 (O_613,N_13863,N_13888);
or UO_614 (O_614,N_13723,N_13828);
and UO_615 (O_615,N_13625,N_14355);
xor UO_616 (O_616,N_14833,N_14448);
or UO_617 (O_617,N_13897,N_14944);
nor UO_618 (O_618,N_13865,N_14184);
nor UO_619 (O_619,N_13852,N_14152);
nand UO_620 (O_620,N_13545,N_14732);
and UO_621 (O_621,N_14431,N_14685);
xor UO_622 (O_622,N_14858,N_14793);
nand UO_623 (O_623,N_14221,N_14300);
and UO_624 (O_624,N_14116,N_14055);
or UO_625 (O_625,N_13739,N_13569);
and UO_626 (O_626,N_13797,N_14075);
or UO_627 (O_627,N_14982,N_13956);
and UO_628 (O_628,N_13784,N_14798);
nand UO_629 (O_629,N_13997,N_13876);
nand UO_630 (O_630,N_13886,N_14816);
xnor UO_631 (O_631,N_13772,N_14829);
nor UO_632 (O_632,N_13655,N_14158);
or UO_633 (O_633,N_14678,N_13558);
nand UO_634 (O_634,N_14423,N_14022);
xor UO_635 (O_635,N_14000,N_14892);
nand UO_636 (O_636,N_13645,N_14977);
or UO_637 (O_637,N_13884,N_13573);
or UO_638 (O_638,N_14060,N_14371);
and UO_639 (O_639,N_14122,N_14879);
nand UO_640 (O_640,N_14708,N_14772);
and UO_641 (O_641,N_14040,N_14820);
nand UO_642 (O_642,N_14141,N_14342);
xnor UO_643 (O_643,N_13996,N_14260);
nor UO_644 (O_644,N_13503,N_14742);
xnor UO_645 (O_645,N_14023,N_14417);
or UO_646 (O_646,N_14277,N_14166);
nor UO_647 (O_647,N_13686,N_13901);
or UO_648 (O_648,N_14252,N_13923);
nor UO_649 (O_649,N_13862,N_14258);
nand UO_650 (O_650,N_14864,N_14298);
xor UO_651 (O_651,N_14493,N_14006);
or UO_652 (O_652,N_13650,N_14771);
and UO_653 (O_653,N_14486,N_14088);
nand UO_654 (O_654,N_14140,N_14869);
and UO_655 (O_655,N_13845,N_14686);
or UO_656 (O_656,N_14283,N_14807);
nor UO_657 (O_657,N_13824,N_14518);
or UO_658 (O_658,N_13838,N_14814);
nand UO_659 (O_659,N_14668,N_13796);
nor UO_660 (O_660,N_14325,N_13821);
nand UO_661 (O_661,N_14684,N_13716);
nand UO_662 (O_662,N_14201,N_14134);
nor UO_663 (O_663,N_14830,N_14428);
nor UO_664 (O_664,N_13684,N_13710);
or UO_665 (O_665,N_14988,N_13501);
nor UO_666 (O_666,N_13728,N_13520);
nand UO_667 (O_667,N_13853,N_14175);
or UO_668 (O_668,N_13607,N_14195);
or UO_669 (O_669,N_13543,N_13952);
nand UO_670 (O_670,N_14538,N_14059);
nor UO_671 (O_671,N_14561,N_13691);
nand UO_672 (O_672,N_14646,N_13771);
or UO_673 (O_673,N_14995,N_14711);
or UO_674 (O_674,N_14245,N_13548);
nand UO_675 (O_675,N_14844,N_14590);
and UO_676 (O_676,N_14765,N_14297);
or UO_677 (O_677,N_13792,N_14808);
nand UO_678 (O_678,N_13912,N_14409);
and UO_679 (O_679,N_13515,N_13830);
and UO_680 (O_680,N_14524,N_13939);
nor UO_681 (O_681,N_14396,N_14191);
nor UO_682 (O_682,N_14854,N_13651);
nor UO_683 (O_683,N_14633,N_13740);
nand UO_684 (O_684,N_13869,N_13801);
nand UO_685 (O_685,N_13858,N_14905);
nor UO_686 (O_686,N_13851,N_13910);
or UO_687 (O_687,N_14377,N_14923);
nand UO_688 (O_688,N_13615,N_14904);
or UO_689 (O_689,N_14198,N_13906);
nand UO_690 (O_690,N_13611,N_13639);
and UO_691 (O_691,N_13810,N_13635);
nand UO_692 (O_692,N_14585,N_14626);
nand UO_693 (O_693,N_13808,N_14066);
or UO_694 (O_694,N_14722,N_14331);
or UO_695 (O_695,N_14385,N_13679);
or UO_696 (O_696,N_14278,N_14033);
xnor UO_697 (O_697,N_13668,N_13785);
nand UO_698 (O_698,N_13881,N_14094);
and UO_699 (O_699,N_13949,N_14557);
nand UO_700 (O_700,N_13899,N_14713);
or UO_701 (O_701,N_14817,N_13689);
or UO_702 (O_702,N_14447,N_14421);
nand UO_703 (O_703,N_14930,N_13957);
or UO_704 (O_704,N_13938,N_14009);
xor UO_705 (O_705,N_14321,N_14477);
nor UO_706 (O_706,N_13559,N_13727);
nand UO_707 (O_707,N_14774,N_13859);
nand UO_708 (O_708,N_14045,N_13733);
nand UO_709 (O_709,N_14051,N_14831);
nand UO_710 (O_710,N_14763,N_13913);
nand UO_711 (O_711,N_13890,N_14567);
or UO_712 (O_712,N_14710,N_13705);
nand UO_713 (O_713,N_14644,N_14380);
xor UO_714 (O_714,N_14938,N_14449);
xor UO_715 (O_715,N_14156,N_13737);
nor UO_716 (O_716,N_14754,N_14735);
and UO_717 (O_717,N_14744,N_14815);
or UO_718 (O_718,N_13696,N_13753);
nor UO_719 (O_719,N_13618,N_14113);
nor UO_720 (O_720,N_14553,N_13734);
and UO_721 (O_721,N_14474,N_14790);
nand UO_722 (O_722,N_13800,N_14649);
nand UO_723 (O_723,N_14778,N_14645);
xor UO_724 (O_724,N_14233,N_14483);
or UO_725 (O_725,N_13911,N_13743);
xnor UO_726 (O_726,N_14570,N_14434);
and UO_727 (O_727,N_14786,N_13768);
or UO_728 (O_728,N_14319,N_14179);
nor UO_729 (O_729,N_14920,N_14679);
or UO_730 (O_730,N_14689,N_14271);
nand UO_731 (O_731,N_14852,N_13561);
nor UO_732 (O_732,N_14035,N_13898);
nor UO_733 (O_733,N_14779,N_14459);
or UO_734 (O_734,N_13709,N_14842);
nor UO_735 (O_735,N_14863,N_14834);
nand UO_736 (O_736,N_13965,N_14097);
nor UO_737 (O_737,N_14404,N_13715);
nor UO_738 (O_738,N_14631,N_14131);
xor UO_739 (O_739,N_14356,N_14738);
nor UO_740 (O_740,N_14349,N_13782);
nand UO_741 (O_741,N_14523,N_13552);
or UO_742 (O_742,N_14211,N_14969);
and UO_743 (O_743,N_13745,N_14789);
nand UO_744 (O_744,N_14189,N_14393);
or UO_745 (O_745,N_14622,N_13878);
or UO_746 (O_746,N_13732,N_14291);
xor UO_747 (O_747,N_13924,N_13868);
or UO_748 (O_748,N_14780,N_14948);
and UO_749 (O_749,N_13546,N_13962);
nor UO_750 (O_750,N_14707,N_14053);
and UO_751 (O_751,N_14323,N_13507);
or UO_752 (O_752,N_14982,N_14844);
and UO_753 (O_753,N_14735,N_13895);
nand UO_754 (O_754,N_14512,N_14517);
nand UO_755 (O_755,N_14217,N_14717);
nor UO_756 (O_756,N_14211,N_14841);
xnor UO_757 (O_757,N_14391,N_14643);
or UO_758 (O_758,N_14847,N_14015);
and UO_759 (O_759,N_14224,N_14162);
nand UO_760 (O_760,N_13887,N_14629);
xnor UO_761 (O_761,N_13609,N_13687);
nor UO_762 (O_762,N_14293,N_14793);
nand UO_763 (O_763,N_13899,N_13931);
or UO_764 (O_764,N_14537,N_14936);
or UO_765 (O_765,N_14130,N_14860);
and UO_766 (O_766,N_13610,N_14651);
or UO_767 (O_767,N_13599,N_14156);
nor UO_768 (O_768,N_14127,N_14806);
nor UO_769 (O_769,N_14034,N_14912);
or UO_770 (O_770,N_14300,N_14421);
xnor UO_771 (O_771,N_14133,N_14496);
nor UO_772 (O_772,N_14386,N_14071);
and UO_773 (O_773,N_14115,N_14574);
or UO_774 (O_774,N_14729,N_13942);
or UO_775 (O_775,N_13608,N_14159);
nor UO_776 (O_776,N_13528,N_14469);
nor UO_777 (O_777,N_13677,N_13550);
or UO_778 (O_778,N_14700,N_13560);
nand UO_779 (O_779,N_14678,N_13548);
xnor UO_780 (O_780,N_14915,N_14867);
xnor UO_781 (O_781,N_13616,N_14151);
or UO_782 (O_782,N_13714,N_13870);
nand UO_783 (O_783,N_14872,N_13949);
or UO_784 (O_784,N_14435,N_14120);
nor UO_785 (O_785,N_13552,N_14296);
and UO_786 (O_786,N_13988,N_14957);
or UO_787 (O_787,N_14399,N_14700);
nand UO_788 (O_788,N_13904,N_14643);
or UO_789 (O_789,N_14366,N_13874);
nor UO_790 (O_790,N_14429,N_14707);
or UO_791 (O_791,N_13680,N_13848);
and UO_792 (O_792,N_14784,N_13846);
and UO_793 (O_793,N_14778,N_14769);
nand UO_794 (O_794,N_14885,N_14425);
nor UO_795 (O_795,N_13780,N_14066);
or UO_796 (O_796,N_13842,N_13534);
nor UO_797 (O_797,N_14231,N_14489);
and UO_798 (O_798,N_13515,N_14275);
or UO_799 (O_799,N_14592,N_13677);
xor UO_800 (O_800,N_14631,N_13552);
or UO_801 (O_801,N_14311,N_14307);
xor UO_802 (O_802,N_14943,N_14355);
and UO_803 (O_803,N_13914,N_13866);
and UO_804 (O_804,N_14879,N_14317);
and UO_805 (O_805,N_13720,N_14169);
nor UO_806 (O_806,N_13579,N_13793);
nand UO_807 (O_807,N_14910,N_13818);
nand UO_808 (O_808,N_14552,N_13697);
nor UO_809 (O_809,N_14864,N_14317);
nor UO_810 (O_810,N_14259,N_14735);
or UO_811 (O_811,N_14476,N_13521);
and UO_812 (O_812,N_14572,N_14788);
and UO_813 (O_813,N_13504,N_13763);
xnor UO_814 (O_814,N_14736,N_14724);
and UO_815 (O_815,N_14631,N_14039);
or UO_816 (O_816,N_14444,N_13729);
xor UO_817 (O_817,N_14682,N_14975);
nor UO_818 (O_818,N_14320,N_13914);
or UO_819 (O_819,N_14957,N_14526);
nor UO_820 (O_820,N_14625,N_13824);
and UO_821 (O_821,N_14371,N_14648);
xor UO_822 (O_822,N_13969,N_14863);
and UO_823 (O_823,N_14634,N_14973);
or UO_824 (O_824,N_14376,N_14633);
and UO_825 (O_825,N_13835,N_14088);
nor UO_826 (O_826,N_14493,N_14514);
or UO_827 (O_827,N_14402,N_14427);
and UO_828 (O_828,N_14220,N_14158);
and UO_829 (O_829,N_13535,N_13826);
xnor UO_830 (O_830,N_13899,N_14108);
nand UO_831 (O_831,N_13658,N_14034);
or UO_832 (O_832,N_13553,N_14531);
or UO_833 (O_833,N_13567,N_13598);
nand UO_834 (O_834,N_14467,N_14196);
nor UO_835 (O_835,N_14464,N_14427);
nand UO_836 (O_836,N_14724,N_14645);
nor UO_837 (O_837,N_13626,N_14896);
nor UO_838 (O_838,N_14022,N_14397);
xor UO_839 (O_839,N_13616,N_14632);
and UO_840 (O_840,N_13750,N_14219);
or UO_841 (O_841,N_14548,N_14742);
and UO_842 (O_842,N_13855,N_14470);
nor UO_843 (O_843,N_14020,N_14337);
nor UO_844 (O_844,N_14821,N_13645);
nand UO_845 (O_845,N_14395,N_14146);
nor UO_846 (O_846,N_14703,N_14722);
or UO_847 (O_847,N_14305,N_13727);
xor UO_848 (O_848,N_14455,N_13800);
or UO_849 (O_849,N_14798,N_14759);
and UO_850 (O_850,N_13835,N_14217);
nand UO_851 (O_851,N_14654,N_14248);
nand UO_852 (O_852,N_13709,N_14719);
or UO_853 (O_853,N_14055,N_14397);
nor UO_854 (O_854,N_14759,N_14584);
and UO_855 (O_855,N_13754,N_14581);
or UO_856 (O_856,N_14084,N_13805);
xnor UO_857 (O_857,N_14604,N_13933);
nand UO_858 (O_858,N_14685,N_14167);
or UO_859 (O_859,N_14704,N_14903);
nor UO_860 (O_860,N_14735,N_13553);
nand UO_861 (O_861,N_13546,N_14937);
xor UO_862 (O_862,N_14165,N_14396);
nor UO_863 (O_863,N_13506,N_14958);
xnor UO_864 (O_864,N_14413,N_14479);
or UO_865 (O_865,N_14992,N_13528);
nand UO_866 (O_866,N_13734,N_13592);
or UO_867 (O_867,N_14708,N_13721);
and UO_868 (O_868,N_14864,N_13565);
nor UO_869 (O_869,N_14117,N_13665);
nor UO_870 (O_870,N_14428,N_14717);
or UO_871 (O_871,N_14583,N_14549);
and UO_872 (O_872,N_13634,N_14065);
xnor UO_873 (O_873,N_13678,N_13721);
or UO_874 (O_874,N_13925,N_13865);
and UO_875 (O_875,N_14995,N_13790);
or UO_876 (O_876,N_14202,N_14715);
and UO_877 (O_877,N_13961,N_14571);
xor UO_878 (O_878,N_14868,N_14776);
nand UO_879 (O_879,N_14047,N_14052);
or UO_880 (O_880,N_14459,N_13603);
nor UO_881 (O_881,N_14778,N_14118);
nand UO_882 (O_882,N_14579,N_14710);
or UO_883 (O_883,N_13807,N_14416);
and UO_884 (O_884,N_13567,N_14524);
xor UO_885 (O_885,N_14371,N_14777);
or UO_886 (O_886,N_14335,N_14109);
or UO_887 (O_887,N_14577,N_13504);
or UO_888 (O_888,N_14986,N_14203);
nor UO_889 (O_889,N_14922,N_13708);
nor UO_890 (O_890,N_14931,N_14062);
and UO_891 (O_891,N_14526,N_14320);
nand UO_892 (O_892,N_14931,N_14054);
and UO_893 (O_893,N_14043,N_14600);
nand UO_894 (O_894,N_13983,N_14654);
nor UO_895 (O_895,N_14046,N_14374);
nand UO_896 (O_896,N_14987,N_14277);
nand UO_897 (O_897,N_14095,N_13531);
or UO_898 (O_898,N_14054,N_14637);
nand UO_899 (O_899,N_14813,N_14556);
nand UO_900 (O_900,N_14189,N_14008);
nand UO_901 (O_901,N_13979,N_13754);
nand UO_902 (O_902,N_13618,N_13597);
or UO_903 (O_903,N_14935,N_13774);
nor UO_904 (O_904,N_14927,N_14973);
nor UO_905 (O_905,N_14246,N_14638);
or UO_906 (O_906,N_14819,N_14255);
and UO_907 (O_907,N_13600,N_14178);
or UO_908 (O_908,N_14257,N_14035);
nand UO_909 (O_909,N_14865,N_14195);
nor UO_910 (O_910,N_14030,N_13979);
or UO_911 (O_911,N_14590,N_13932);
nor UO_912 (O_912,N_14516,N_13545);
nand UO_913 (O_913,N_14765,N_13936);
nor UO_914 (O_914,N_14995,N_13844);
nand UO_915 (O_915,N_14910,N_13999);
and UO_916 (O_916,N_14884,N_13668);
nand UO_917 (O_917,N_14471,N_14705);
nand UO_918 (O_918,N_14087,N_14346);
nor UO_919 (O_919,N_14433,N_14056);
nand UO_920 (O_920,N_14628,N_14559);
nor UO_921 (O_921,N_13944,N_14836);
nor UO_922 (O_922,N_13511,N_13964);
or UO_923 (O_923,N_14747,N_13898);
nand UO_924 (O_924,N_13664,N_14364);
nand UO_925 (O_925,N_14174,N_13597);
and UO_926 (O_926,N_14538,N_13991);
and UO_927 (O_927,N_14781,N_14398);
or UO_928 (O_928,N_14085,N_14112);
nor UO_929 (O_929,N_13710,N_14393);
nor UO_930 (O_930,N_14874,N_14373);
and UO_931 (O_931,N_13606,N_14726);
nand UO_932 (O_932,N_13936,N_14834);
or UO_933 (O_933,N_14883,N_14148);
or UO_934 (O_934,N_14334,N_14199);
or UO_935 (O_935,N_13975,N_14652);
nor UO_936 (O_936,N_14451,N_14691);
and UO_937 (O_937,N_14090,N_13796);
or UO_938 (O_938,N_14385,N_13887);
and UO_939 (O_939,N_14787,N_14503);
nand UO_940 (O_940,N_13568,N_14974);
or UO_941 (O_941,N_14453,N_14380);
nor UO_942 (O_942,N_14448,N_13701);
nor UO_943 (O_943,N_14002,N_14566);
and UO_944 (O_944,N_13987,N_13805);
and UO_945 (O_945,N_13938,N_13841);
xor UO_946 (O_946,N_14723,N_14668);
and UO_947 (O_947,N_14458,N_14812);
and UO_948 (O_948,N_14921,N_13966);
and UO_949 (O_949,N_14951,N_14883);
nor UO_950 (O_950,N_14827,N_14106);
and UO_951 (O_951,N_13645,N_13919);
and UO_952 (O_952,N_14399,N_13931);
nor UO_953 (O_953,N_14023,N_13654);
or UO_954 (O_954,N_14904,N_14953);
nand UO_955 (O_955,N_14532,N_14338);
and UO_956 (O_956,N_13748,N_14063);
or UO_957 (O_957,N_14126,N_14316);
nor UO_958 (O_958,N_14797,N_14687);
and UO_959 (O_959,N_13925,N_13720);
nor UO_960 (O_960,N_13964,N_14762);
nand UO_961 (O_961,N_14472,N_14204);
nor UO_962 (O_962,N_13699,N_14061);
nor UO_963 (O_963,N_14644,N_14701);
nor UO_964 (O_964,N_14323,N_13878);
nand UO_965 (O_965,N_14313,N_14283);
or UO_966 (O_966,N_14624,N_14633);
nand UO_967 (O_967,N_14794,N_14907);
and UO_968 (O_968,N_13780,N_14200);
nand UO_969 (O_969,N_13988,N_14565);
nand UO_970 (O_970,N_13582,N_13828);
and UO_971 (O_971,N_14325,N_14363);
or UO_972 (O_972,N_14501,N_13988);
and UO_973 (O_973,N_14148,N_13513);
or UO_974 (O_974,N_13796,N_14884);
and UO_975 (O_975,N_13857,N_14937);
nor UO_976 (O_976,N_14260,N_13706);
nand UO_977 (O_977,N_13629,N_14053);
and UO_978 (O_978,N_14744,N_14870);
and UO_979 (O_979,N_14867,N_14455);
or UO_980 (O_980,N_14216,N_14087);
or UO_981 (O_981,N_14336,N_13690);
nor UO_982 (O_982,N_14976,N_13761);
nand UO_983 (O_983,N_14343,N_13597);
or UO_984 (O_984,N_14666,N_14356);
or UO_985 (O_985,N_13795,N_14688);
or UO_986 (O_986,N_13791,N_13832);
or UO_987 (O_987,N_14029,N_14796);
nand UO_988 (O_988,N_14710,N_14918);
and UO_989 (O_989,N_13834,N_14092);
nor UO_990 (O_990,N_14477,N_13861);
nand UO_991 (O_991,N_14130,N_13680);
xor UO_992 (O_992,N_14170,N_14348);
and UO_993 (O_993,N_14912,N_14352);
or UO_994 (O_994,N_14375,N_14490);
and UO_995 (O_995,N_13686,N_13833);
or UO_996 (O_996,N_13660,N_14654);
nand UO_997 (O_997,N_13980,N_14089);
nand UO_998 (O_998,N_14705,N_14567);
or UO_999 (O_999,N_14684,N_14830);
nand UO_1000 (O_1000,N_14719,N_14140);
xor UO_1001 (O_1001,N_14968,N_13671);
or UO_1002 (O_1002,N_14475,N_13753);
and UO_1003 (O_1003,N_14471,N_13592);
nand UO_1004 (O_1004,N_14071,N_14131);
and UO_1005 (O_1005,N_14831,N_13589);
or UO_1006 (O_1006,N_14045,N_13652);
or UO_1007 (O_1007,N_14785,N_14901);
nand UO_1008 (O_1008,N_13801,N_14378);
or UO_1009 (O_1009,N_13530,N_14589);
nor UO_1010 (O_1010,N_14661,N_14846);
nand UO_1011 (O_1011,N_14159,N_14872);
nor UO_1012 (O_1012,N_14299,N_14720);
nor UO_1013 (O_1013,N_14534,N_14925);
nor UO_1014 (O_1014,N_14177,N_14270);
xnor UO_1015 (O_1015,N_13980,N_14535);
or UO_1016 (O_1016,N_14387,N_14428);
nor UO_1017 (O_1017,N_13872,N_14423);
or UO_1018 (O_1018,N_14123,N_14890);
nand UO_1019 (O_1019,N_14462,N_14005);
nand UO_1020 (O_1020,N_13991,N_14295);
or UO_1021 (O_1021,N_14077,N_14316);
xnor UO_1022 (O_1022,N_14280,N_14514);
and UO_1023 (O_1023,N_14263,N_14793);
or UO_1024 (O_1024,N_13990,N_14531);
xor UO_1025 (O_1025,N_13686,N_14098);
nor UO_1026 (O_1026,N_13749,N_13619);
nor UO_1027 (O_1027,N_14971,N_14203);
nor UO_1028 (O_1028,N_14984,N_13631);
and UO_1029 (O_1029,N_14410,N_13666);
nor UO_1030 (O_1030,N_14695,N_13505);
and UO_1031 (O_1031,N_14891,N_14909);
nand UO_1032 (O_1032,N_13910,N_14899);
nor UO_1033 (O_1033,N_14408,N_13783);
or UO_1034 (O_1034,N_14406,N_14592);
nor UO_1035 (O_1035,N_14296,N_14916);
nor UO_1036 (O_1036,N_13705,N_14637);
xor UO_1037 (O_1037,N_14587,N_14710);
nor UO_1038 (O_1038,N_14718,N_14605);
nor UO_1039 (O_1039,N_13936,N_14011);
or UO_1040 (O_1040,N_14352,N_14983);
nand UO_1041 (O_1041,N_14168,N_13821);
or UO_1042 (O_1042,N_14908,N_14816);
nor UO_1043 (O_1043,N_14197,N_13974);
nand UO_1044 (O_1044,N_14219,N_13541);
or UO_1045 (O_1045,N_14537,N_14281);
xnor UO_1046 (O_1046,N_13697,N_13822);
nand UO_1047 (O_1047,N_14042,N_14495);
nand UO_1048 (O_1048,N_14970,N_14263);
and UO_1049 (O_1049,N_14770,N_13523);
or UO_1050 (O_1050,N_14839,N_13971);
nor UO_1051 (O_1051,N_14416,N_13893);
xnor UO_1052 (O_1052,N_13635,N_14259);
and UO_1053 (O_1053,N_14688,N_14485);
nor UO_1054 (O_1054,N_13779,N_14387);
nor UO_1055 (O_1055,N_13921,N_13753);
nor UO_1056 (O_1056,N_14258,N_14462);
xnor UO_1057 (O_1057,N_14135,N_13565);
xor UO_1058 (O_1058,N_13991,N_14096);
nor UO_1059 (O_1059,N_14772,N_14631);
and UO_1060 (O_1060,N_14242,N_13970);
or UO_1061 (O_1061,N_13887,N_14128);
and UO_1062 (O_1062,N_14914,N_14441);
nand UO_1063 (O_1063,N_13687,N_14612);
and UO_1064 (O_1064,N_14524,N_13663);
and UO_1065 (O_1065,N_14970,N_13934);
and UO_1066 (O_1066,N_13650,N_13976);
xnor UO_1067 (O_1067,N_14573,N_13890);
nand UO_1068 (O_1068,N_13920,N_13514);
and UO_1069 (O_1069,N_13805,N_14232);
nand UO_1070 (O_1070,N_13550,N_14224);
nor UO_1071 (O_1071,N_13891,N_13732);
or UO_1072 (O_1072,N_14813,N_13859);
or UO_1073 (O_1073,N_14136,N_13974);
nor UO_1074 (O_1074,N_13730,N_14676);
and UO_1075 (O_1075,N_14217,N_14393);
xor UO_1076 (O_1076,N_14022,N_14866);
nor UO_1077 (O_1077,N_14217,N_14789);
and UO_1078 (O_1078,N_14581,N_14178);
nor UO_1079 (O_1079,N_13810,N_14219);
nand UO_1080 (O_1080,N_14638,N_13975);
nor UO_1081 (O_1081,N_14063,N_14396);
and UO_1082 (O_1082,N_13763,N_14944);
xnor UO_1083 (O_1083,N_13553,N_14098);
nor UO_1084 (O_1084,N_14517,N_14547);
xnor UO_1085 (O_1085,N_13562,N_13559);
xnor UO_1086 (O_1086,N_14217,N_13935);
or UO_1087 (O_1087,N_14752,N_14483);
nor UO_1088 (O_1088,N_14059,N_14550);
or UO_1089 (O_1089,N_14114,N_13687);
nor UO_1090 (O_1090,N_13920,N_13660);
nor UO_1091 (O_1091,N_14273,N_14470);
nand UO_1092 (O_1092,N_14610,N_14359);
nor UO_1093 (O_1093,N_14323,N_14818);
or UO_1094 (O_1094,N_13528,N_14348);
nor UO_1095 (O_1095,N_14014,N_13601);
or UO_1096 (O_1096,N_14476,N_14305);
xnor UO_1097 (O_1097,N_14810,N_14236);
nand UO_1098 (O_1098,N_14927,N_14961);
nand UO_1099 (O_1099,N_14845,N_14942);
nor UO_1100 (O_1100,N_13810,N_13712);
nor UO_1101 (O_1101,N_13901,N_14910);
nand UO_1102 (O_1102,N_14990,N_14333);
and UO_1103 (O_1103,N_13799,N_14149);
or UO_1104 (O_1104,N_13921,N_13853);
nand UO_1105 (O_1105,N_13714,N_13865);
xnor UO_1106 (O_1106,N_13857,N_14601);
or UO_1107 (O_1107,N_13915,N_14392);
nor UO_1108 (O_1108,N_14823,N_14273);
or UO_1109 (O_1109,N_13980,N_13576);
or UO_1110 (O_1110,N_14570,N_14903);
nand UO_1111 (O_1111,N_14454,N_13972);
nand UO_1112 (O_1112,N_13514,N_14784);
and UO_1113 (O_1113,N_14082,N_14224);
or UO_1114 (O_1114,N_13981,N_13644);
and UO_1115 (O_1115,N_14698,N_13568);
nor UO_1116 (O_1116,N_14574,N_14486);
and UO_1117 (O_1117,N_14882,N_14945);
or UO_1118 (O_1118,N_14316,N_13816);
or UO_1119 (O_1119,N_14764,N_14743);
and UO_1120 (O_1120,N_14299,N_14482);
or UO_1121 (O_1121,N_14281,N_14050);
and UO_1122 (O_1122,N_13880,N_13517);
nand UO_1123 (O_1123,N_14076,N_14883);
nor UO_1124 (O_1124,N_14116,N_14414);
nand UO_1125 (O_1125,N_14661,N_14490);
nand UO_1126 (O_1126,N_14938,N_14563);
or UO_1127 (O_1127,N_14126,N_13888);
nand UO_1128 (O_1128,N_14006,N_14214);
nand UO_1129 (O_1129,N_14946,N_14126);
and UO_1130 (O_1130,N_13906,N_14139);
nor UO_1131 (O_1131,N_13972,N_14494);
or UO_1132 (O_1132,N_14801,N_13559);
and UO_1133 (O_1133,N_13905,N_14356);
nand UO_1134 (O_1134,N_14410,N_14116);
and UO_1135 (O_1135,N_14057,N_13884);
and UO_1136 (O_1136,N_14340,N_13687);
nor UO_1137 (O_1137,N_14877,N_14892);
nor UO_1138 (O_1138,N_14768,N_13927);
nand UO_1139 (O_1139,N_13637,N_14167);
and UO_1140 (O_1140,N_13978,N_14704);
and UO_1141 (O_1141,N_13828,N_13649);
xnor UO_1142 (O_1142,N_14186,N_14772);
nor UO_1143 (O_1143,N_14819,N_14850);
nand UO_1144 (O_1144,N_13781,N_14356);
and UO_1145 (O_1145,N_14828,N_13612);
nand UO_1146 (O_1146,N_14635,N_14297);
nand UO_1147 (O_1147,N_14594,N_14246);
nand UO_1148 (O_1148,N_14399,N_14011);
and UO_1149 (O_1149,N_13618,N_14579);
nor UO_1150 (O_1150,N_14949,N_13810);
or UO_1151 (O_1151,N_13545,N_13692);
nand UO_1152 (O_1152,N_13930,N_14269);
or UO_1153 (O_1153,N_13632,N_14134);
nor UO_1154 (O_1154,N_13621,N_14063);
or UO_1155 (O_1155,N_13785,N_14696);
or UO_1156 (O_1156,N_13902,N_14748);
nand UO_1157 (O_1157,N_14673,N_14958);
xor UO_1158 (O_1158,N_14412,N_14822);
or UO_1159 (O_1159,N_14041,N_14113);
or UO_1160 (O_1160,N_13563,N_13524);
xnor UO_1161 (O_1161,N_14720,N_14441);
nor UO_1162 (O_1162,N_14150,N_14443);
or UO_1163 (O_1163,N_13758,N_14142);
nor UO_1164 (O_1164,N_13630,N_14653);
xnor UO_1165 (O_1165,N_14550,N_14171);
nand UO_1166 (O_1166,N_14705,N_14694);
or UO_1167 (O_1167,N_13538,N_14322);
and UO_1168 (O_1168,N_14103,N_14823);
and UO_1169 (O_1169,N_14761,N_14660);
xor UO_1170 (O_1170,N_14350,N_14427);
or UO_1171 (O_1171,N_13747,N_14775);
nand UO_1172 (O_1172,N_14127,N_14858);
nor UO_1173 (O_1173,N_14006,N_14485);
xor UO_1174 (O_1174,N_13513,N_14860);
or UO_1175 (O_1175,N_14072,N_13628);
and UO_1176 (O_1176,N_14975,N_14888);
and UO_1177 (O_1177,N_14832,N_13914);
or UO_1178 (O_1178,N_14200,N_14303);
nor UO_1179 (O_1179,N_13511,N_14114);
xnor UO_1180 (O_1180,N_14488,N_14593);
nand UO_1181 (O_1181,N_14216,N_14176);
nand UO_1182 (O_1182,N_13928,N_13638);
and UO_1183 (O_1183,N_13992,N_14282);
nor UO_1184 (O_1184,N_14201,N_14070);
and UO_1185 (O_1185,N_14576,N_14521);
or UO_1186 (O_1186,N_14441,N_13946);
nor UO_1187 (O_1187,N_13782,N_14691);
nor UO_1188 (O_1188,N_14409,N_14198);
nor UO_1189 (O_1189,N_13887,N_14666);
and UO_1190 (O_1190,N_14672,N_14394);
nand UO_1191 (O_1191,N_13618,N_14355);
nand UO_1192 (O_1192,N_14207,N_14171);
or UO_1193 (O_1193,N_14141,N_14485);
and UO_1194 (O_1194,N_14855,N_13966);
and UO_1195 (O_1195,N_14676,N_14644);
nand UO_1196 (O_1196,N_14479,N_14142);
xnor UO_1197 (O_1197,N_14295,N_14833);
or UO_1198 (O_1198,N_14976,N_14449);
and UO_1199 (O_1199,N_14932,N_13799);
or UO_1200 (O_1200,N_14853,N_14583);
nor UO_1201 (O_1201,N_14100,N_14589);
nand UO_1202 (O_1202,N_14699,N_13700);
nor UO_1203 (O_1203,N_14292,N_13518);
xor UO_1204 (O_1204,N_14443,N_14497);
nand UO_1205 (O_1205,N_14283,N_13750);
or UO_1206 (O_1206,N_13831,N_14400);
nor UO_1207 (O_1207,N_14986,N_14294);
or UO_1208 (O_1208,N_13609,N_14343);
nor UO_1209 (O_1209,N_14904,N_14604);
or UO_1210 (O_1210,N_14802,N_14740);
nor UO_1211 (O_1211,N_14336,N_13529);
or UO_1212 (O_1212,N_13846,N_13516);
and UO_1213 (O_1213,N_13963,N_14174);
or UO_1214 (O_1214,N_13564,N_14370);
and UO_1215 (O_1215,N_14312,N_13994);
xnor UO_1216 (O_1216,N_14285,N_14872);
or UO_1217 (O_1217,N_14650,N_14396);
or UO_1218 (O_1218,N_13810,N_14100);
nor UO_1219 (O_1219,N_14458,N_14316);
nand UO_1220 (O_1220,N_13983,N_14669);
nor UO_1221 (O_1221,N_14716,N_13896);
or UO_1222 (O_1222,N_13759,N_13786);
and UO_1223 (O_1223,N_13688,N_14805);
and UO_1224 (O_1224,N_13675,N_14972);
nor UO_1225 (O_1225,N_14854,N_14681);
and UO_1226 (O_1226,N_14167,N_14347);
nor UO_1227 (O_1227,N_14884,N_14131);
nor UO_1228 (O_1228,N_14082,N_13590);
nor UO_1229 (O_1229,N_13522,N_14513);
xor UO_1230 (O_1230,N_13854,N_14390);
nor UO_1231 (O_1231,N_14510,N_14427);
or UO_1232 (O_1232,N_13940,N_14969);
nand UO_1233 (O_1233,N_14157,N_13668);
and UO_1234 (O_1234,N_13676,N_14357);
xor UO_1235 (O_1235,N_13568,N_13837);
nor UO_1236 (O_1236,N_13759,N_14193);
or UO_1237 (O_1237,N_13775,N_14292);
or UO_1238 (O_1238,N_14161,N_14755);
nand UO_1239 (O_1239,N_14635,N_13670);
nand UO_1240 (O_1240,N_13609,N_14315);
nor UO_1241 (O_1241,N_14553,N_14481);
nor UO_1242 (O_1242,N_13804,N_13571);
and UO_1243 (O_1243,N_14757,N_13976);
nand UO_1244 (O_1244,N_14307,N_14059);
nor UO_1245 (O_1245,N_13980,N_13699);
and UO_1246 (O_1246,N_14166,N_14612);
xnor UO_1247 (O_1247,N_14278,N_14271);
or UO_1248 (O_1248,N_14009,N_14015);
nand UO_1249 (O_1249,N_13595,N_14341);
or UO_1250 (O_1250,N_14869,N_14052);
and UO_1251 (O_1251,N_13668,N_14058);
nor UO_1252 (O_1252,N_13608,N_13533);
and UO_1253 (O_1253,N_13575,N_14066);
nand UO_1254 (O_1254,N_14389,N_14236);
nand UO_1255 (O_1255,N_14451,N_13810);
or UO_1256 (O_1256,N_14581,N_14467);
nand UO_1257 (O_1257,N_14604,N_14535);
and UO_1258 (O_1258,N_14743,N_14619);
xnor UO_1259 (O_1259,N_14897,N_14472);
and UO_1260 (O_1260,N_13591,N_14593);
or UO_1261 (O_1261,N_14320,N_14537);
or UO_1262 (O_1262,N_14018,N_14319);
nand UO_1263 (O_1263,N_14792,N_14837);
nor UO_1264 (O_1264,N_14753,N_14917);
nor UO_1265 (O_1265,N_13713,N_13833);
or UO_1266 (O_1266,N_14921,N_13656);
nor UO_1267 (O_1267,N_14552,N_14360);
and UO_1268 (O_1268,N_14816,N_14755);
or UO_1269 (O_1269,N_14366,N_14983);
nand UO_1270 (O_1270,N_14482,N_13947);
nand UO_1271 (O_1271,N_14384,N_13841);
nand UO_1272 (O_1272,N_14537,N_14999);
nand UO_1273 (O_1273,N_14713,N_14072);
nand UO_1274 (O_1274,N_13903,N_14432);
and UO_1275 (O_1275,N_13550,N_13525);
or UO_1276 (O_1276,N_13529,N_14795);
and UO_1277 (O_1277,N_13510,N_14443);
nor UO_1278 (O_1278,N_14447,N_14257);
or UO_1279 (O_1279,N_14110,N_14234);
nand UO_1280 (O_1280,N_14458,N_14143);
or UO_1281 (O_1281,N_13718,N_14390);
xnor UO_1282 (O_1282,N_14467,N_14395);
xor UO_1283 (O_1283,N_14244,N_13891);
or UO_1284 (O_1284,N_13874,N_13535);
and UO_1285 (O_1285,N_14096,N_13670);
nor UO_1286 (O_1286,N_14580,N_14503);
nor UO_1287 (O_1287,N_14919,N_13880);
nor UO_1288 (O_1288,N_13966,N_14089);
and UO_1289 (O_1289,N_14099,N_14667);
and UO_1290 (O_1290,N_14384,N_14142);
nor UO_1291 (O_1291,N_14554,N_14915);
nor UO_1292 (O_1292,N_13568,N_14013);
and UO_1293 (O_1293,N_13631,N_13985);
and UO_1294 (O_1294,N_14372,N_13945);
nand UO_1295 (O_1295,N_14005,N_14080);
nor UO_1296 (O_1296,N_13707,N_14646);
or UO_1297 (O_1297,N_14869,N_14233);
or UO_1298 (O_1298,N_14292,N_13523);
or UO_1299 (O_1299,N_14998,N_14470);
nor UO_1300 (O_1300,N_14976,N_14436);
nand UO_1301 (O_1301,N_13690,N_14711);
or UO_1302 (O_1302,N_13508,N_13571);
nand UO_1303 (O_1303,N_13860,N_14325);
nor UO_1304 (O_1304,N_14496,N_14766);
and UO_1305 (O_1305,N_13911,N_14924);
xor UO_1306 (O_1306,N_13791,N_14239);
and UO_1307 (O_1307,N_13856,N_14810);
nand UO_1308 (O_1308,N_14773,N_13947);
or UO_1309 (O_1309,N_14655,N_13938);
and UO_1310 (O_1310,N_13617,N_13808);
nor UO_1311 (O_1311,N_14798,N_13665);
nor UO_1312 (O_1312,N_14232,N_14815);
or UO_1313 (O_1313,N_14308,N_14445);
nor UO_1314 (O_1314,N_14098,N_13565);
and UO_1315 (O_1315,N_14813,N_13718);
or UO_1316 (O_1316,N_13814,N_13999);
or UO_1317 (O_1317,N_13834,N_14665);
or UO_1318 (O_1318,N_14760,N_14386);
or UO_1319 (O_1319,N_13523,N_13833);
or UO_1320 (O_1320,N_14325,N_13983);
nand UO_1321 (O_1321,N_14229,N_14006);
nand UO_1322 (O_1322,N_14049,N_13611);
nor UO_1323 (O_1323,N_14808,N_14897);
nor UO_1324 (O_1324,N_14993,N_14846);
nand UO_1325 (O_1325,N_14329,N_14693);
or UO_1326 (O_1326,N_13562,N_13947);
nand UO_1327 (O_1327,N_14399,N_13713);
nor UO_1328 (O_1328,N_14315,N_13674);
or UO_1329 (O_1329,N_13757,N_14280);
nor UO_1330 (O_1330,N_13760,N_13971);
and UO_1331 (O_1331,N_14524,N_14837);
or UO_1332 (O_1332,N_13846,N_14786);
or UO_1333 (O_1333,N_13621,N_14818);
and UO_1334 (O_1334,N_14387,N_14749);
nor UO_1335 (O_1335,N_14636,N_14742);
nand UO_1336 (O_1336,N_13672,N_14467);
or UO_1337 (O_1337,N_14669,N_14273);
and UO_1338 (O_1338,N_13567,N_13994);
nand UO_1339 (O_1339,N_14637,N_14719);
and UO_1340 (O_1340,N_14060,N_14032);
and UO_1341 (O_1341,N_14633,N_14890);
nand UO_1342 (O_1342,N_14092,N_14609);
nor UO_1343 (O_1343,N_13842,N_14831);
or UO_1344 (O_1344,N_14067,N_14516);
nor UO_1345 (O_1345,N_13709,N_14681);
xnor UO_1346 (O_1346,N_13570,N_14858);
and UO_1347 (O_1347,N_13996,N_14709);
and UO_1348 (O_1348,N_13595,N_14448);
or UO_1349 (O_1349,N_14061,N_14613);
nor UO_1350 (O_1350,N_13805,N_14432);
and UO_1351 (O_1351,N_14615,N_13808);
and UO_1352 (O_1352,N_14858,N_14135);
or UO_1353 (O_1353,N_14907,N_14367);
xnor UO_1354 (O_1354,N_14545,N_14596);
or UO_1355 (O_1355,N_14052,N_14578);
or UO_1356 (O_1356,N_14173,N_13660);
nand UO_1357 (O_1357,N_13576,N_13517);
nor UO_1358 (O_1358,N_14028,N_14428);
nand UO_1359 (O_1359,N_14995,N_14783);
nor UO_1360 (O_1360,N_14564,N_13722);
nor UO_1361 (O_1361,N_14748,N_14280);
nor UO_1362 (O_1362,N_13926,N_14104);
nand UO_1363 (O_1363,N_14792,N_14773);
nand UO_1364 (O_1364,N_13748,N_13715);
and UO_1365 (O_1365,N_14305,N_14052);
xnor UO_1366 (O_1366,N_13542,N_14449);
nand UO_1367 (O_1367,N_14400,N_14071);
and UO_1368 (O_1368,N_14533,N_14435);
nand UO_1369 (O_1369,N_14557,N_14637);
nand UO_1370 (O_1370,N_14188,N_14520);
and UO_1371 (O_1371,N_14485,N_14375);
nor UO_1372 (O_1372,N_14905,N_14811);
nand UO_1373 (O_1373,N_14551,N_14321);
xnor UO_1374 (O_1374,N_13726,N_14808);
and UO_1375 (O_1375,N_13852,N_14059);
and UO_1376 (O_1376,N_14257,N_14875);
nand UO_1377 (O_1377,N_14957,N_14616);
and UO_1378 (O_1378,N_14364,N_14401);
and UO_1379 (O_1379,N_14729,N_14485);
and UO_1380 (O_1380,N_14639,N_14827);
xor UO_1381 (O_1381,N_13631,N_14250);
nand UO_1382 (O_1382,N_14961,N_14017);
nor UO_1383 (O_1383,N_14950,N_13866);
nor UO_1384 (O_1384,N_14421,N_14141);
xnor UO_1385 (O_1385,N_14445,N_14742);
and UO_1386 (O_1386,N_14502,N_14040);
nor UO_1387 (O_1387,N_13712,N_14376);
or UO_1388 (O_1388,N_14117,N_13913);
nor UO_1389 (O_1389,N_14774,N_13880);
or UO_1390 (O_1390,N_14136,N_14002);
nor UO_1391 (O_1391,N_14980,N_14994);
nand UO_1392 (O_1392,N_14856,N_13686);
and UO_1393 (O_1393,N_13710,N_13810);
and UO_1394 (O_1394,N_13774,N_14816);
nand UO_1395 (O_1395,N_14293,N_14146);
nand UO_1396 (O_1396,N_14774,N_14124);
nor UO_1397 (O_1397,N_13871,N_13865);
nor UO_1398 (O_1398,N_13875,N_14880);
nand UO_1399 (O_1399,N_14511,N_14956);
and UO_1400 (O_1400,N_14673,N_13701);
and UO_1401 (O_1401,N_13686,N_14408);
nand UO_1402 (O_1402,N_13571,N_14572);
xor UO_1403 (O_1403,N_14062,N_14051);
nor UO_1404 (O_1404,N_14426,N_14632);
and UO_1405 (O_1405,N_14210,N_14729);
xnor UO_1406 (O_1406,N_14676,N_14767);
nor UO_1407 (O_1407,N_14401,N_14200);
nor UO_1408 (O_1408,N_14758,N_14479);
or UO_1409 (O_1409,N_14812,N_14378);
and UO_1410 (O_1410,N_14815,N_14550);
xnor UO_1411 (O_1411,N_14245,N_14436);
xor UO_1412 (O_1412,N_13935,N_13739);
and UO_1413 (O_1413,N_13626,N_14090);
or UO_1414 (O_1414,N_14892,N_13777);
and UO_1415 (O_1415,N_14266,N_14554);
and UO_1416 (O_1416,N_14634,N_13622);
nor UO_1417 (O_1417,N_14008,N_14033);
and UO_1418 (O_1418,N_14174,N_14189);
nor UO_1419 (O_1419,N_14477,N_14045);
and UO_1420 (O_1420,N_13506,N_14626);
or UO_1421 (O_1421,N_14344,N_14692);
and UO_1422 (O_1422,N_14351,N_14490);
and UO_1423 (O_1423,N_14013,N_14131);
nand UO_1424 (O_1424,N_14691,N_13646);
nor UO_1425 (O_1425,N_14152,N_14180);
nor UO_1426 (O_1426,N_14187,N_13871);
nand UO_1427 (O_1427,N_13786,N_13803);
xor UO_1428 (O_1428,N_13522,N_14496);
xor UO_1429 (O_1429,N_14562,N_13889);
nor UO_1430 (O_1430,N_14345,N_13526);
or UO_1431 (O_1431,N_14141,N_13988);
or UO_1432 (O_1432,N_14053,N_13964);
nand UO_1433 (O_1433,N_14624,N_14362);
nor UO_1434 (O_1434,N_14141,N_14700);
nor UO_1435 (O_1435,N_13802,N_14405);
nor UO_1436 (O_1436,N_14805,N_14484);
and UO_1437 (O_1437,N_14378,N_14141);
and UO_1438 (O_1438,N_14929,N_13509);
or UO_1439 (O_1439,N_14602,N_14863);
xnor UO_1440 (O_1440,N_14720,N_14148);
and UO_1441 (O_1441,N_13838,N_13947);
nand UO_1442 (O_1442,N_14786,N_13570);
nor UO_1443 (O_1443,N_13942,N_14796);
and UO_1444 (O_1444,N_13558,N_14355);
xor UO_1445 (O_1445,N_13668,N_13557);
nand UO_1446 (O_1446,N_14997,N_14219);
nor UO_1447 (O_1447,N_13688,N_14892);
nand UO_1448 (O_1448,N_14928,N_14987);
xnor UO_1449 (O_1449,N_14270,N_14471);
or UO_1450 (O_1450,N_13626,N_14836);
nor UO_1451 (O_1451,N_13552,N_14832);
or UO_1452 (O_1452,N_14283,N_13868);
nor UO_1453 (O_1453,N_14177,N_14565);
xor UO_1454 (O_1454,N_14381,N_14394);
and UO_1455 (O_1455,N_14981,N_13956);
and UO_1456 (O_1456,N_13502,N_13650);
nor UO_1457 (O_1457,N_14542,N_13653);
nand UO_1458 (O_1458,N_13772,N_14503);
xnor UO_1459 (O_1459,N_13900,N_13620);
nor UO_1460 (O_1460,N_14228,N_14244);
nor UO_1461 (O_1461,N_14997,N_14232);
or UO_1462 (O_1462,N_13995,N_14263);
nand UO_1463 (O_1463,N_14170,N_13784);
nor UO_1464 (O_1464,N_14895,N_14335);
and UO_1465 (O_1465,N_14611,N_13878);
nand UO_1466 (O_1466,N_14351,N_14519);
nor UO_1467 (O_1467,N_14737,N_14003);
nor UO_1468 (O_1468,N_14743,N_13543);
or UO_1469 (O_1469,N_13920,N_14421);
nor UO_1470 (O_1470,N_14196,N_13769);
nand UO_1471 (O_1471,N_13826,N_14088);
or UO_1472 (O_1472,N_13639,N_14532);
nand UO_1473 (O_1473,N_14818,N_14173);
nand UO_1474 (O_1474,N_14564,N_14784);
and UO_1475 (O_1475,N_14598,N_14475);
and UO_1476 (O_1476,N_14976,N_13524);
xnor UO_1477 (O_1477,N_14664,N_13795);
or UO_1478 (O_1478,N_13891,N_13799);
nand UO_1479 (O_1479,N_13627,N_14090);
or UO_1480 (O_1480,N_14334,N_14383);
and UO_1481 (O_1481,N_14923,N_14554);
and UO_1482 (O_1482,N_14545,N_14494);
xor UO_1483 (O_1483,N_14057,N_13679);
nand UO_1484 (O_1484,N_13925,N_14245);
and UO_1485 (O_1485,N_13705,N_13914);
nor UO_1486 (O_1486,N_14535,N_13984);
nand UO_1487 (O_1487,N_13635,N_14280);
nor UO_1488 (O_1488,N_14685,N_13864);
nor UO_1489 (O_1489,N_13741,N_14376);
nor UO_1490 (O_1490,N_14068,N_14771);
nor UO_1491 (O_1491,N_13935,N_13815);
or UO_1492 (O_1492,N_13978,N_13995);
or UO_1493 (O_1493,N_14315,N_14243);
nor UO_1494 (O_1494,N_14342,N_14806);
nor UO_1495 (O_1495,N_14241,N_14403);
or UO_1496 (O_1496,N_13528,N_14815);
nand UO_1497 (O_1497,N_14397,N_14145);
nand UO_1498 (O_1498,N_13773,N_13950);
and UO_1499 (O_1499,N_14455,N_14469);
nand UO_1500 (O_1500,N_14725,N_14575);
or UO_1501 (O_1501,N_14536,N_14551);
and UO_1502 (O_1502,N_14123,N_14290);
and UO_1503 (O_1503,N_14333,N_14551);
or UO_1504 (O_1504,N_14070,N_14982);
or UO_1505 (O_1505,N_13723,N_13727);
or UO_1506 (O_1506,N_13909,N_14620);
or UO_1507 (O_1507,N_13565,N_13682);
or UO_1508 (O_1508,N_13543,N_14883);
nand UO_1509 (O_1509,N_14046,N_13608);
xnor UO_1510 (O_1510,N_14258,N_14979);
nor UO_1511 (O_1511,N_13982,N_13966);
and UO_1512 (O_1512,N_14348,N_14886);
or UO_1513 (O_1513,N_14392,N_14361);
or UO_1514 (O_1514,N_14001,N_14084);
nand UO_1515 (O_1515,N_14130,N_14110);
or UO_1516 (O_1516,N_14704,N_14471);
and UO_1517 (O_1517,N_14384,N_13924);
nor UO_1518 (O_1518,N_14214,N_14102);
nand UO_1519 (O_1519,N_14960,N_14207);
or UO_1520 (O_1520,N_13809,N_13767);
nor UO_1521 (O_1521,N_13642,N_14779);
nor UO_1522 (O_1522,N_14304,N_13528);
nand UO_1523 (O_1523,N_14230,N_13560);
nor UO_1524 (O_1524,N_13963,N_14104);
nand UO_1525 (O_1525,N_14940,N_14648);
or UO_1526 (O_1526,N_14248,N_14237);
or UO_1527 (O_1527,N_14219,N_13947);
nor UO_1528 (O_1528,N_14580,N_13992);
and UO_1529 (O_1529,N_14357,N_14933);
and UO_1530 (O_1530,N_13990,N_14280);
and UO_1531 (O_1531,N_14874,N_14519);
nor UO_1532 (O_1532,N_13781,N_13766);
nor UO_1533 (O_1533,N_13552,N_13764);
nand UO_1534 (O_1534,N_14796,N_14126);
nand UO_1535 (O_1535,N_14951,N_13647);
nor UO_1536 (O_1536,N_13720,N_14027);
nor UO_1537 (O_1537,N_14369,N_13814);
and UO_1538 (O_1538,N_14283,N_13671);
nand UO_1539 (O_1539,N_13571,N_14370);
nand UO_1540 (O_1540,N_14280,N_14893);
or UO_1541 (O_1541,N_14723,N_13750);
and UO_1542 (O_1542,N_13794,N_14805);
xnor UO_1543 (O_1543,N_14155,N_13832);
and UO_1544 (O_1544,N_14905,N_14575);
or UO_1545 (O_1545,N_13513,N_13540);
or UO_1546 (O_1546,N_14393,N_14380);
or UO_1547 (O_1547,N_13633,N_14081);
nor UO_1548 (O_1548,N_14390,N_14704);
nor UO_1549 (O_1549,N_14403,N_14676);
xor UO_1550 (O_1550,N_14313,N_14429);
nand UO_1551 (O_1551,N_14836,N_13675);
nor UO_1552 (O_1552,N_14801,N_13898);
and UO_1553 (O_1553,N_14177,N_14187);
nor UO_1554 (O_1554,N_13908,N_13599);
nor UO_1555 (O_1555,N_14922,N_13693);
nor UO_1556 (O_1556,N_13787,N_14866);
nand UO_1557 (O_1557,N_14607,N_14090);
or UO_1558 (O_1558,N_14139,N_13824);
nand UO_1559 (O_1559,N_14379,N_14053);
nand UO_1560 (O_1560,N_14082,N_14997);
or UO_1561 (O_1561,N_14189,N_13959);
xor UO_1562 (O_1562,N_14568,N_14890);
nor UO_1563 (O_1563,N_14731,N_14457);
or UO_1564 (O_1564,N_13733,N_14972);
or UO_1565 (O_1565,N_14745,N_14632);
and UO_1566 (O_1566,N_14611,N_14804);
and UO_1567 (O_1567,N_14574,N_14490);
and UO_1568 (O_1568,N_13574,N_13781);
or UO_1569 (O_1569,N_14543,N_14069);
or UO_1570 (O_1570,N_14580,N_14779);
nand UO_1571 (O_1571,N_13934,N_14640);
nor UO_1572 (O_1572,N_14640,N_14112);
nor UO_1573 (O_1573,N_14861,N_14887);
or UO_1574 (O_1574,N_14056,N_14885);
and UO_1575 (O_1575,N_13666,N_13632);
and UO_1576 (O_1576,N_14584,N_14135);
nor UO_1577 (O_1577,N_13556,N_14353);
nand UO_1578 (O_1578,N_13951,N_14462);
and UO_1579 (O_1579,N_13688,N_14551);
or UO_1580 (O_1580,N_13567,N_14949);
and UO_1581 (O_1581,N_14903,N_13959);
and UO_1582 (O_1582,N_13929,N_14207);
xor UO_1583 (O_1583,N_14895,N_14153);
nand UO_1584 (O_1584,N_14993,N_14093);
nor UO_1585 (O_1585,N_14475,N_14643);
and UO_1586 (O_1586,N_13759,N_14595);
or UO_1587 (O_1587,N_14977,N_14320);
or UO_1588 (O_1588,N_14072,N_13845);
xnor UO_1589 (O_1589,N_14400,N_14930);
nor UO_1590 (O_1590,N_14970,N_14870);
or UO_1591 (O_1591,N_14819,N_13739);
xnor UO_1592 (O_1592,N_14821,N_13867);
xor UO_1593 (O_1593,N_14322,N_14384);
or UO_1594 (O_1594,N_14971,N_14969);
or UO_1595 (O_1595,N_14489,N_14118);
nand UO_1596 (O_1596,N_14315,N_14000);
xor UO_1597 (O_1597,N_13958,N_14219);
nor UO_1598 (O_1598,N_13863,N_14780);
nor UO_1599 (O_1599,N_13552,N_13683);
nand UO_1600 (O_1600,N_13627,N_14984);
and UO_1601 (O_1601,N_13659,N_14048);
xnor UO_1602 (O_1602,N_13998,N_14173);
nand UO_1603 (O_1603,N_14241,N_14171);
nand UO_1604 (O_1604,N_13520,N_14274);
nand UO_1605 (O_1605,N_14877,N_14256);
or UO_1606 (O_1606,N_14709,N_13916);
nand UO_1607 (O_1607,N_13568,N_14923);
or UO_1608 (O_1608,N_14068,N_13626);
nor UO_1609 (O_1609,N_14349,N_13500);
nor UO_1610 (O_1610,N_13672,N_14451);
nor UO_1611 (O_1611,N_14410,N_13669);
xor UO_1612 (O_1612,N_14393,N_13727);
or UO_1613 (O_1613,N_13639,N_14653);
nand UO_1614 (O_1614,N_14468,N_13534);
xor UO_1615 (O_1615,N_14764,N_14487);
and UO_1616 (O_1616,N_14666,N_14683);
nor UO_1617 (O_1617,N_13587,N_14558);
nand UO_1618 (O_1618,N_13745,N_14548);
and UO_1619 (O_1619,N_14113,N_14557);
nand UO_1620 (O_1620,N_14513,N_14199);
nor UO_1621 (O_1621,N_13622,N_14278);
nor UO_1622 (O_1622,N_13609,N_14053);
nor UO_1623 (O_1623,N_14706,N_14740);
and UO_1624 (O_1624,N_13645,N_13766);
nor UO_1625 (O_1625,N_14746,N_14007);
and UO_1626 (O_1626,N_14577,N_13655);
or UO_1627 (O_1627,N_14608,N_14181);
xnor UO_1628 (O_1628,N_14435,N_14863);
and UO_1629 (O_1629,N_14517,N_13753);
nor UO_1630 (O_1630,N_13898,N_14140);
nor UO_1631 (O_1631,N_14104,N_14954);
nor UO_1632 (O_1632,N_14524,N_14951);
and UO_1633 (O_1633,N_14690,N_13501);
nor UO_1634 (O_1634,N_13891,N_13560);
nor UO_1635 (O_1635,N_14879,N_14094);
or UO_1636 (O_1636,N_13913,N_14186);
and UO_1637 (O_1637,N_14931,N_14557);
or UO_1638 (O_1638,N_14152,N_14472);
nor UO_1639 (O_1639,N_14000,N_14527);
and UO_1640 (O_1640,N_13697,N_14867);
nor UO_1641 (O_1641,N_13912,N_13867);
or UO_1642 (O_1642,N_13917,N_14652);
nor UO_1643 (O_1643,N_13678,N_14079);
or UO_1644 (O_1644,N_13590,N_14243);
and UO_1645 (O_1645,N_13901,N_14815);
xnor UO_1646 (O_1646,N_14625,N_14233);
nor UO_1647 (O_1647,N_14520,N_13591);
xnor UO_1648 (O_1648,N_14259,N_13857);
or UO_1649 (O_1649,N_14621,N_14687);
and UO_1650 (O_1650,N_14456,N_14093);
and UO_1651 (O_1651,N_13721,N_14107);
nand UO_1652 (O_1652,N_14595,N_14126);
nor UO_1653 (O_1653,N_14096,N_14746);
or UO_1654 (O_1654,N_14480,N_13530);
and UO_1655 (O_1655,N_14931,N_14610);
nor UO_1656 (O_1656,N_14942,N_13697);
nand UO_1657 (O_1657,N_14552,N_14084);
and UO_1658 (O_1658,N_14997,N_13871);
nor UO_1659 (O_1659,N_13601,N_14547);
nand UO_1660 (O_1660,N_14102,N_14126);
nand UO_1661 (O_1661,N_14425,N_14141);
and UO_1662 (O_1662,N_13661,N_13894);
nor UO_1663 (O_1663,N_14881,N_14875);
or UO_1664 (O_1664,N_13640,N_13900);
nand UO_1665 (O_1665,N_14902,N_14998);
nor UO_1666 (O_1666,N_13737,N_14018);
nand UO_1667 (O_1667,N_14358,N_14590);
nand UO_1668 (O_1668,N_13566,N_13683);
xor UO_1669 (O_1669,N_13868,N_13933);
or UO_1670 (O_1670,N_13888,N_13855);
or UO_1671 (O_1671,N_14212,N_13591);
xor UO_1672 (O_1672,N_13818,N_14933);
or UO_1673 (O_1673,N_14020,N_13778);
nor UO_1674 (O_1674,N_14714,N_14861);
and UO_1675 (O_1675,N_14925,N_14438);
xor UO_1676 (O_1676,N_14152,N_13806);
and UO_1677 (O_1677,N_14937,N_14252);
nand UO_1678 (O_1678,N_13918,N_13555);
nand UO_1679 (O_1679,N_14003,N_14919);
nand UO_1680 (O_1680,N_13675,N_14022);
or UO_1681 (O_1681,N_14298,N_14910);
nand UO_1682 (O_1682,N_14197,N_14884);
nand UO_1683 (O_1683,N_13769,N_13972);
or UO_1684 (O_1684,N_14192,N_14919);
nand UO_1685 (O_1685,N_13728,N_14604);
and UO_1686 (O_1686,N_13922,N_13521);
and UO_1687 (O_1687,N_14807,N_14250);
nor UO_1688 (O_1688,N_13883,N_14355);
or UO_1689 (O_1689,N_14243,N_14560);
nor UO_1690 (O_1690,N_13841,N_14750);
or UO_1691 (O_1691,N_13873,N_14447);
nand UO_1692 (O_1692,N_14707,N_14670);
xnor UO_1693 (O_1693,N_14474,N_13864);
and UO_1694 (O_1694,N_14416,N_13603);
nand UO_1695 (O_1695,N_14270,N_14326);
xnor UO_1696 (O_1696,N_14863,N_13956);
xnor UO_1697 (O_1697,N_13902,N_14360);
nor UO_1698 (O_1698,N_14006,N_14906);
and UO_1699 (O_1699,N_13809,N_13638);
and UO_1700 (O_1700,N_14032,N_14110);
nor UO_1701 (O_1701,N_13753,N_14426);
and UO_1702 (O_1702,N_14809,N_14679);
xnor UO_1703 (O_1703,N_14209,N_14002);
nor UO_1704 (O_1704,N_13956,N_13549);
nor UO_1705 (O_1705,N_14802,N_14852);
nor UO_1706 (O_1706,N_13509,N_13810);
and UO_1707 (O_1707,N_14644,N_14614);
and UO_1708 (O_1708,N_13684,N_14044);
and UO_1709 (O_1709,N_13664,N_13570);
nor UO_1710 (O_1710,N_14407,N_14905);
and UO_1711 (O_1711,N_13508,N_14660);
xnor UO_1712 (O_1712,N_14761,N_14481);
xnor UO_1713 (O_1713,N_13691,N_14158);
xnor UO_1714 (O_1714,N_14564,N_14270);
and UO_1715 (O_1715,N_13707,N_13678);
and UO_1716 (O_1716,N_13717,N_14150);
nor UO_1717 (O_1717,N_14056,N_13869);
nor UO_1718 (O_1718,N_14958,N_14990);
nand UO_1719 (O_1719,N_13795,N_14506);
or UO_1720 (O_1720,N_13579,N_13612);
or UO_1721 (O_1721,N_14400,N_14063);
xor UO_1722 (O_1722,N_14360,N_14096);
nand UO_1723 (O_1723,N_13524,N_14651);
xnor UO_1724 (O_1724,N_13520,N_14783);
nand UO_1725 (O_1725,N_14953,N_14276);
nor UO_1726 (O_1726,N_13829,N_14675);
and UO_1727 (O_1727,N_13925,N_13759);
nor UO_1728 (O_1728,N_13819,N_14250);
nor UO_1729 (O_1729,N_14481,N_14473);
and UO_1730 (O_1730,N_14895,N_14766);
or UO_1731 (O_1731,N_14624,N_13794);
or UO_1732 (O_1732,N_14193,N_14018);
xnor UO_1733 (O_1733,N_14631,N_14909);
nand UO_1734 (O_1734,N_13682,N_14268);
and UO_1735 (O_1735,N_14688,N_13673);
xor UO_1736 (O_1736,N_14953,N_13714);
nor UO_1737 (O_1737,N_13556,N_14557);
or UO_1738 (O_1738,N_14820,N_14708);
and UO_1739 (O_1739,N_13944,N_14910);
xor UO_1740 (O_1740,N_13567,N_14115);
and UO_1741 (O_1741,N_14199,N_14843);
nor UO_1742 (O_1742,N_14707,N_14691);
and UO_1743 (O_1743,N_14835,N_13829);
nor UO_1744 (O_1744,N_14972,N_14385);
and UO_1745 (O_1745,N_14607,N_14310);
or UO_1746 (O_1746,N_14232,N_13760);
nor UO_1747 (O_1747,N_14928,N_13608);
and UO_1748 (O_1748,N_13873,N_14720);
nand UO_1749 (O_1749,N_14867,N_13676);
xor UO_1750 (O_1750,N_13600,N_14730);
nor UO_1751 (O_1751,N_14050,N_14476);
or UO_1752 (O_1752,N_14413,N_13608);
and UO_1753 (O_1753,N_14056,N_14554);
or UO_1754 (O_1754,N_14668,N_14696);
and UO_1755 (O_1755,N_14629,N_14440);
nor UO_1756 (O_1756,N_14252,N_13840);
xnor UO_1757 (O_1757,N_13644,N_14844);
and UO_1758 (O_1758,N_13541,N_13873);
or UO_1759 (O_1759,N_14669,N_13693);
nand UO_1760 (O_1760,N_13697,N_14295);
and UO_1761 (O_1761,N_14967,N_14604);
and UO_1762 (O_1762,N_14376,N_13955);
nor UO_1763 (O_1763,N_14678,N_14452);
or UO_1764 (O_1764,N_14508,N_14046);
or UO_1765 (O_1765,N_14863,N_14434);
xor UO_1766 (O_1766,N_13922,N_14596);
and UO_1767 (O_1767,N_14315,N_14638);
xor UO_1768 (O_1768,N_14619,N_14549);
nor UO_1769 (O_1769,N_14148,N_14343);
and UO_1770 (O_1770,N_14901,N_13998);
and UO_1771 (O_1771,N_14101,N_14328);
nand UO_1772 (O_1772,N_14247,N_14138);
xor UO_1773 (O_1773,N_14722,N_14501);
nand UO_1774 (O_1774,N_13885,N_14109);
and UO_1775 (O_1775,N_14109,N_13700);
and UO_1776 (O_1776,N_14153,N_14397);
nand UO_1777 (O_1777,N_13932,N_13778);
nand UO_1778 (O_1778,N_14461,N_14218);
and UO_1779 (O_1779,N_14044,N_14745);
nand UO_1780 (O_1780,N_13990,N_14981);
nand UO_1781 (O_1781,N_14253,N_14508);
nand UO_1782 (O_1782,N_13934,N_14082);
xor UO_1783 (O_1783,N_13653,N_13817);
and UO_1784 (O_1784,N_14079,N_14525);
nor UO_1785 (O_1785,N_14576,N_14490);
nor UO_1786 (O_1786,N_14329,N_14023);
xor UO_1787 (O_1787,N_13916,N_14622);
or UO_1788 (O_1788,N_13570,N_14547);
nand UO_1789 (O_1789,N_14177,N_13990);
or UO_1790 (O_1790,N_13532,N_14159);
nor UO_1791 (O_1791,N_13736,N_13971);
and UO_1792 (O_1792,N_14150,N_14598);
xnor UO_1793 (O_1793,N_14212,N_14440);
or UO_1794 (O_1794,N_14870,N_14840);
nor UO_1795 (O_1795,N_13648,N_14765);
and UO_1796 (O_1796,N_14609,N_14814);
nor UO_1797 (O_1797,N_13606,N_14012);
nor UO_1798 (O_1798,N_14483,N_14234);
or UO_1799 (O_1799,N_13559,N_14862);
and UO_1800 (O_1800,N_14495,N_14470);
nor UO_1801 (O_1801,N_13519,N_14256);
nor UO_1802 (O_1802,N_14539,N_14798);
nor UO_1803 (O_1803,N_14260,N_13783);
nand UO_1804 (O_1804,N_13562,N_14126);
nor UO_1805 (O_1805,N_14997,N_14220);
and UO_1806 (O_1806,N_13871,N_14838);
xnor UO_1807 (O_1807,N_14706,N_14310);
and UO_1808 (O_1808,N_14666,N_13689);
xnor UO_1809 (O_1809,N_14321,N_14909);
nor UO_1810 (O_1810,N_14573,N_14308);
and UO_1811 (O_1811,N_14382,N_14410);
xor UO_1812 (O_1812,N_14755,N_13731);
nor UO_1813 (O_1813,N_14452,N_14826);
nand UO_1814 (O_1814,N_13913,N_13767);
nor UO_1815 (O_1815,N_14902,N_14495);
nand UO_1816 (O_1816,N_14852,N_14097);
and UO_1817 (O_1817,N_13560,N_13859);
or UO_1818 (O_1818,N_14403,N_14533);
and UO_1819 (O_1819,N_14447,N_14734);
or UO_1820 (O_1820,N_13902,N_14366);
nor UO_1821 (O_1821,N_14647,N_14968);
xor UO_1822 (O_1822,N_13792,N_14113);
nor UO_1823 (O_1823,N_13656,N_14392);
xnor UO_1824 (O_1824,N_14962,N_14364);
and UO_1825 (O_1825,N_14195,N_13962);
xor UO_1826 (O_1826,N_13710,N_14309);
nor UO_1827 (O_1827,N_14003,N_14558);
nor UO_1828 (O_1828,N_14678,N_13810);
nor UO_1829 (O_1829,N_13577,N_14188);
nand UO_1830 (O_1830,N_14122,N_14522);
and UO_1831 (O_1831,N_14732,N_14437);
nor UO_1832 (O_1832,N_14154,N_14875);
nand UO_1833 (O_1833,N_13508,N_14076);
nand UO_1834 (O_1834,N_14791,N_13836);
nor UO_1835 (O_1835,N_14264,N_14978);
and UO_1836 (O_1836,N_14775,N_14357);
nand UO_1837 (O_1837,N_14615,N_13790);
nor UO_1838 (O_1838,N_14985,N_13876);
and UO_1839 (O_1839,N_14342,N_13944);
xnor UO_1840 (O_1840,N_13808,N_14802);
nor UO_1841 (O_1841,N_13971,N_14761);
nand UO_1842 (O_1842,N_14297,N_14717);
xor UO_1843 (O_1843,N_14564,N_14869);
and UO_1844 (O_1844,N_14822,N_14485);
nand UO_1845 (O_1845,N_13686,N_14312);
nand UO_1846 (O_1846,N_14914,N_14644);
or UO_1847 (O_1847,N_14951,N_14285);
and UO_1848 (O_1848,N_14392,N_13996);
xor UO_1849 (O_1849,N_14324,N_14756);
or UO_1850 (O_1850,N_13534,N_14378);
nor UO_1851 (O_1851,N_14041,N_14565);
nor UO_1852 (O_1852,N_14380,N_14576);
nor UO_1853 (O_1853,N_14026,N_14556);
xnor UO_1854 (O_1854,N_14622,N_13569);
and UO_1855 (O_1855,N_14489,N_14902);
and UO_1856 (O_1856,N_14943,N_14008);
and UO_1857 (O_1857,N_13801,N_14318);
nand UO_1858 (O_1858,N_14821,N_14220);
nor UO_1859 (O_1859,N_14510,N_14450);
nor UO_1860 (O_1860,N_14754,N_13969);
nand UO_1861 (O_1861,N_14740,N_14690);
and UO_1862 (O_1862,N_14855,N_14798);
or UO_1863 (O_1863,N_14578,N_14908);
or UO_1864 (O_1864,N_14921,N_14179);
xnor UO_1865 (O_1865,N_13906,N_13841);
or UO_1866 (O_1866,N_14399,N_13793);
or UO_1867 (O_1867,N_14395,N_13638);
or UO_1868 (O_1868,N_14446,N_14338);
nor UO_1869 (O_1869,N_14736,N_14677);
and UO_1870 (O_1870,N_14608,N_14251);
or UO_1871 (O_1871,N_14089,N_14404);
nor UO_1872 (O_1872,N_14380,N_14274);
nor UO_1873 (O_1873,N_13610,N_13927);
nand UO_1874 (O_1874,N_13572,N_13755);
or UO_1875 (O_1875,N_14282,N_13793);
nor UO_1876 (O_1876,N_14625,N_14051);
or UO_1877 (O_1877,N_13746,N_13735);
nor UO_1878 (O_1878,N_14889,N_13952);
or UO_1879 (O_1879,N_14193,N_13607);
and UO_1880 (O_1880,N_14454,N_13892);
and UO_1881 (O_1881,N_14146,N_14761);
nor UO_1882 (O_1882,N_14270,N_14580);
nand UO_1883 (O_1883,N_14740,N_14043);
xor UO_1884 (O_1884,N_13522,N_14180);
xnor UO_1885 (O_1885,N_13712,N_14367);
or UO_1886 (O_1886,N_14369,N_13920);
nand UO_1887 (O_1887,N_13939,N_14311);
and UO_1888 (O_1888,N_14497,N_14837);
nand UO_1889 (O_1889,N_13865,N_14618);
or UO_1890 (O_1890,N_14123,N_13625);
and UO_1891 (O_1891,N_14535,N_14408);
nor UO_1892 (O_1892,N_14063,N_13797);
nor UO_1893 (O_1893,N_14446,N_14727);
or UO_1894 (O_1894,N_13653,N_14910);
xnor UO_1895 (O_1895,N_14607,N_14247);
and UO_1896 (O_1896,N_14695,N_13526);
nand UO_1897 (O_1897,N_14098,N_14078);
and UO_1898 (O_1898,N_14314,N_14578);
or UO_1899 (O_1899,N_14835,N_13650);
nand UO_1900 (O_1900,N_14026,N_14517);
and UO_1901 (O_1901,N_14217,N_13818);
or UO_1902 (O_1902,N_14719,N_13568);
or UO_1903 (O_1903,N_14561,N_14255);
xnor UO_1904 (O_1904,N_14727,N_13813);
or UO_1905 (O_1905,N_13948,N_14975);
nor UO_1906 (O_1906,N_14215,N_14091);
or UO_1907 (O_1907,N_14977,N_13911);
or UO_1908 (O_1908,N_14418,N_14871);
nor UO_1909 (O_1909,N_14443,N_14872);
or UO_1910 (O_1910,N_14765,N_14905);
nor UO_1911 (O_1911,N_14716,N_14293);
xor UO_1912 (O_1912,N_14230,N_14319);
and UO_1913 (O_1913,N_13658,N_13800);
nor UO_1914 (O_1914,N_14492,N_14092);
or UO_1915 (O_1915,N_14067,N_14154);
nor UO_1916 (O_1916,N_14171,N_14549);
or UO_1917 (O_1917,N_13958,N_13605);
nor UO_1918 (O_1918,N_13585,N_14383);
nor UO_1919 (O_1919,N_14612,N_14635);
and UO_1920 (O_1920,N_13751,N_13937);
xor UO_1921 (O_1921,N_13509,N_14013);
and UO_1922 (O_1922,N_14331,N_14646);
or UO_1923 (O_1923,N_14699,N_14883);
and UO_1924 (O_1924,N_14500,N_14622);
and UO_1925 (O_1925,N_13686,N_14332);
and UO_1926 (O_1926,N_14335,N_14354);
nand UO_1927 (O_1927,N_13603,N_13568);
nor UO_1928 (O_1928,N_13558,N_14950);
nor UO_1929 (O_1929,N_14356,N_13680);
or UO_1930 (O_1930,N_14922,N_13798);
or UO_1931 (O_1931,N_13917,N_14037);
and UO_1932 (O_1932,N_13741,N_13617);
and UO_1933 (O_1933,N_13560,N_14801);
nand UO_1934 (O_1934,N_13710,N_14866);
xnor UO_1935 (O_1935,N_14520,N_14146);
nand UO_1936 (O_1936,N_14687,N_14587);
nor UO_1937 (O_1937,N_13841,N_13756);
or UO_1938 (O_1938,N_14262,N_14147);
or UO_1939 (O_1939,N_14001,N_14868);
or UO_1940 (O_1940,N_14595,N_13916);
xor UO_1941 (O_1941,N_14873,N_14309);
nor UO_1942 (O_1942,N_14384,N_14223);
nand UO_1943 (O_1943,N_14652,N_14062);
or UO_1944 (O_1944,N_14290,N_14182);
nor UO_1945 (O_1945,N_13748,N_14321);
nand UO_1946 (O_1946,N_14534,N_14687);
nor UO_1947 (O_1947,N_14579,N_14519);
or UO_1948 (O_1948,N_14371,N_14664);
and UO_1949 (O_1949,N_14223,N_14659);
and UO_1950 (O_1950,N_13715,N_14227);
and UO_1951 (O_1951,N_13918,N_13698);
xnor UO_1952 (O_1952,N_14863,N_14465);
and UO_1953 (O_1953,N_14543,N_14580);
xor UO_1954 (O_1954,N_14158,N_14659);
and UO_1955 (O_1955,N_13670,N_14485);
and UO_1956 (O_1956,N_13974,N_13525);
nand UO_1957 (O_1957,N_14493,N_14168);
and UO_1958 (O_1958,N_14216,N_13588);
xor UO_1959 (O_1959,N_14345,N_14080);
or UO_1960 (O_1960,N_14643,N_14913);
and UO_1961 (O_1961,N_14795,N_13513);
and UO_1962 (O_1962,N_14816,N_14738);
nand UO_1963 (O_1963,N_13655,N_13952);
and UO_1964 (O_1964,N_14607,N_14891);
or UO_1965 (O_1965,N_13533,N_14795);
and UO_1966 (O_1966,N_13729,N_13831);
or UO_1967 (O_1967,N_14136,N_14164);
nor UO_1968 (O_1968,N_14071,N_14936);
and UO_1969 (O_1969,N_13696,N_14666);
nor UO_1970 (O_1970,N_14343,N_13730);
or UO_1971 (O_1971,N_13520,N_14374);
nand UO_1972 (O_1972,N_14800,N_14946);
and UO_1973 (O_1973,N_14242,N_13552);
nand UO_1974 (O_1974,N_14134,N_13864);
nand UO_1975 (O_1975,N_14786,N_13682);
xnor UO_1976 (O_1976,N_14658,N_13898);
nand UO_1977 (O_1977,N_14795,N_14549);
or UO_1978 (O_1978,N_14000,N_13804);
xor UO_1979 (O_1979,N_13756,N_14817);
and UO_1980 (O_1980,N_14277,N_14982);
and UO_1981 (O_1981,N_14330,N_13999);
nor UO_1982 (O_1982,N_13863,N_13547);
nor UO_1983 (O_1983,N_13581,N_14041);
nor UO_1984 (O_1984,N_14908,N_14646);
nand UO_1985 (O_1985,N_13738,N_14151);
nor UO_1986 (O_1986,N_14465,N_14757);
xnor UO_1987 (O_1987,N_14183,N_13507);
nor UO_1988 (O_1988,N_13781,N_14770);
and UO_1989 (O_1989,N_13830,N_13843);
nor UO_1990 (O_1990,N_14772,N_14368);
or UO_1991 (O_1991,N_14825,N_14638);
nor UO_1992 (O_1992,N_14526,N_14884);
and UO_1993 (O_1993,N_14778,N_14791);
and UO_1994 (O_1994,N_14257,N_13553);
or UO_1995 (O_1995,N_14441,N_14202);
nor UO_1996 (O_1996,N_13766,N_14738);
or UO_1997 (O_1997,N_13874,N_14312);
and UO_1998 (O_1998,N_13941,N_13642);
nand UO_1999 (O_1999,N_14101,N_13557);
endmodule