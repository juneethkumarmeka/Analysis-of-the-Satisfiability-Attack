module basic_1000_10000_1500_10_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_617,In_344);
nor U1 (N_1,In_878,In_749);
nand U2 (N_2,In_108,In_971);
and U3 (N_3,In_133,In_355);
xnor U4 (N_4,In_451,In_301);
and U5 (N_5,In_574,In_171);
nand U6 (N_6,In_713,In_42);
nand U7 (N_7,In_558,In_189);
nand U8 (N_8,In_82,In_769);
and U9 (N_9,In_507,In_478);
nand U10 (N_10,In_13,In_907);
nor U11 (N_11,In_41,In_914);
or U12 (N_12,In_76,In_899);
or U13 (N_13,In_231,In_519);
and U14 (N_14,In_191,In_837);
nor U15 (N_15,In_604,In_658);
nand U16 (N_16,In_819,In_846);
nor U17 (N_17,In_710,In_93);
nand U18 (N_18,In_951,In_363);
nand U19 (N_19,In_619,In_47);
or U20 (N_20,In_159,In_849);
and U21 (N_21,In_14,In_320);
and U22 (N_22,In_77,In_917);
or U23 (N_23,In_804,In_556);
or U24 (N_24,In_15,In_938);
or U25 (N_25,In_341,In_591);
or U26 (N_26,In_516,In_226);
or U27 (N_27,In_957,In_889);
nor U28 (N_28,In_857,In_921);
nand U29 (N_29,In_902,In_598);
and U30 (N_30,In_655,In_873);
nand U31 (N_31,In_445,In_594);
nand U32 (N_32,In_151,In_186);
or U33 (N_33,In_496,In_648);
or U34 (N_34,In_979,In_221);
nand U35 (N_35,In_161,In_188);
and U36 (N_36,In_386,In_409);
nor U37 (N_37,In_7,In_261);
nor U38 (N_38,In_799,In_306);
and U39 (N_39,In_152,In_179);
nand U40 (N_40,In_909,In_501);
nor U41 (N_41,In_420,In_297);
or U42 (N_42,In_962,In_414);
or U43 (N_43,In_187,In_667);
or U44 (N_44,In_475,In_61);
or U45 (N_45,In_162,In_986);
and U46 (N_46,In_455,In_130);
nor U47 (N_47,In_148,In_612);
nand U48 (N_48,In_240,In_531);
and U49 (N_49,In_563,In_838);
and U50 (N_50,In_375,In_610);
nor U51 (N_51,In_722,In_416);
nand U52 (N_52,In_51,In_310);
nand U53 (N_53,In_721,In_298);
or U54 (N_54,In_2,In_918);
nor U55 (N_55,In_779,In_442);
and U56 (N_56,In_953,In_806);
nand U57 (N_57,In_506,In_967);
or U58 (N_58,In_803,In_318);
nand U59 (N_59,In_104,In_437);
nand U60 (N_60,In_754,In_374);
nand U61 (N_61,In_266,In_607);
nand U62 (N_62,In_595,In_239);
nand U63 (N_63,In_224,In_113);
nand U64 (N_64,In_941,In_787);
or U65 (N_65,In_812,In_650);
nor U66 (N_66,In_402,In_8);
nand U67 (N_67,In_985,In_517);
or U68 (N_68,In_639,In_682);
and U69 (N_69,In_342,In_925);
nand U70 (N_70,In_237,In_55);
or U71 (N_71,In_23,In_248);
nor U72 (N_72,In_465,In_331);
nor U73 (N_73,In_174,In_584);
nor U74 (N_74,In_391,In_602);
or U75 (N_75,In_348,In_369);
or U76 (N_76,In_949,In_980);
and U77 (N_77,In_141,In_659);
and U78 (N_78,In_50,In_101);
and U79 (N_79,In_305,In_218);
nand U80 (N_80,In_114,In_353);
nor U81 (N_81,In_945,In_714);
nor U82 (N_82,In_800,In_277);
and U83 (N_83,In_774,In_268);
and U84 (N_84,In_377,In_145);
nand U85 (N_85,In_974,In_820);
nor U86 (N_86,In_6,In_647);
nor U87 (N_87,In_815,In_698);
nand U88 (N_88,In_695,In_184);
nand U89 (N_89,In_760,In_903);
and U90 (N_90,In_782,In_222);
nand U91 (N_91,In_735,In_382);
and U92 (N_92,In_431,In_276);
nor U93 (N_93,In_468,In_768);
or U94 (N_94,In_410,In_669);
and U95 (N_95,In_615,In_250);
nor U96 (N_96,In_989,In_923);
nand U97 (N_97,In_272,In_347);
and U98 (N_98,In_705,In_508);
nor U99 (N_99,In_366,In_89);
or U100 (N_100,In_270,In_643);
and U101 (N_101,In_195,In_279);
and U102 (N_102,In_258,In_756);
nand U103 (N_103,In_396,In_349);
or U104 (N_104,In_38,In_217);
or U105 (N_105,In_614,In_958);
nand U106 (N_106,In_214,In_673);
nor U107 (N_107,In_327,In_16);
nor U108 (N_108,In_500,In_624);
or U109 (N_109,In_379,In_0);
and U110 (N_110,In_99,In_110);
nand U111 (N_111,In_841,In_361);
or U112 (N_112,In_888,In_523);
and U113 (N_113,In_733,In_763);
or U114 (N_114,In_213,In_160);
or U115 (N_115,In_510,In_84);
or U116 (N_116,In_177,In_470);
nor U117 (N_117,In_893,In_628);
nor U118 (N_118,In_4,In_679);
nor U119 (N_119,In_170,In_824);
nor U120 (N_120,In_915,In_392);
nand U121 (N_121,In_245,In_515);
nor U122 (N_122,In_227,In_703);
nor U123 (N_123,In_626,In_3);
or U124 (N_124,In_540,In_687);
or U125 (N_125,In_309,In_863);
and U126 (N_126,In_27,In_541);
nand U127 (N_127,In_371,In_532);
or U128 (N_128,In_886,In_326);
nor U129 (N_129,In_993,In_924);
or U130 (N_130,In_220,In_460);
nor U131 (N_131,In_429,In_536);
and U132 (N_132,In_172,In_976);
or U133 (N_133,In_632,In_75);
nand U134 (N_134,In_577,In_637);
and U135 (N_135,In_216,In_546);
nor U136 (N_136,In_573,In_645);
or U137 (N_137,In_977,In_491);
and U138 (N_138,In_587,In_872);
and U139 (N_139,In_209,In_193);
and U140 (N_140,In_895,In_393);
nand U141 (N_141,In_499,In_201);
nor U142 (N_142,In_406,In_64);
nor U143 (N_143,In_9,In_596);
or U144 (N_144,In_404,In_773);
nand U145 (N_145,In_477,In_850);
or U146 (N_146,In_818,In_96);
or U147 (N_147,In_57,In_443);
nor U148 (N_148,In_204,In_996);
and U149 (N_149,In_770,In_137);
or U150 (N_150,In_997,In_205);
or U151 (N_151,In_35,In_275);
nand U152 (N_152,In_808,In_85);
and U153 (N_153,In_131,In_879);
or U154 (N_154,In_944,In_107);
nor U155 (N_155,In_880,In_704);
nor U156 (N_156,In_388,In_700);
and U157 (N_157,In_946,In_814);
or U158 (N_158,In_593,In_807);
nand U159 (N_159,In_729,In_559);
nor U160 (N_160,In_555,In_701);
or U161 (N_161,In_330,In_94);
nand U162 (N_162,In_109,In_581);
and U163 (N_163,In_882,In_926);
nor U164 (N_164,In_63,In_464);
nor U165 (N_165,In_656,In_970);
and U166 (N_166,In_817,In_712);
or U167 (N_167,In_219,In_691);
or U168 (N_168,In_702,In_871);
and U169 (N_169,In_92,In_461);
and U170 (N_170,In_97,In_19);
and U171 (N_171,In_998,In_920);
nor U172 (N_172,In_434,In_79);
or U173 (N_173,In_585,In_982);
nand U174 (N_174,In_328,In_654);
nand U175 (N_175,In_795,In_288);
nor U176 (N_176,In_829,In_865);
and U177 (N_177,In_447,In_618);
nor U178 (N_178,In_883,In_296);
nand U179 (N_179,In_322,In_823);
or U180 (N_180,In_621,In_335);
and U181 (N_181,In_454,In_672);
nor U182 (N_182,In_132,In_480);
nand U183 (N_183,In_358,In_805);
and U184 (N_184,In_10,In_529);
and U185 (N_185,In_425,In_723);
nand U186 (N_186,In_436,In_955);
or U187 (N_187,In_395,In_70);
nor U188 (N_188,In_731,In_605);
nor U189 (N_189,In_860,In_357);
or U190 (N_190,In_183,In_987);
or U191 (N_191,In_198,In_332);
nor U192 (N_192,In_725,In_611);
xnor U193 (N_193,In_972,In_518);
xor U194 (N_194,In_586,In_257);
and U195 (N_195,In_33,In_26);
nor U196 (N_196,In_539,In_727);
and U197 (N_197,In_965,In_307);
and U198 (N_198,In_848,In_742);
or U199 (N_199,In_684,In_764);
and U200 (N_200,In_25,In_345);
or U201 (N_201,In_281,In_928);
and U202 (N_202,In_87,In_671);
nand U203 (N_203,In_947,In_367);
or U204 (N_204,In_831,In_329);
nor U205 (N_205,In_24,In_780);
or U206 (N_206,In_960,In_744);
or U207 (N_207,In_211,In_564);
nor U208 (N_208,In_285,In_324);
and U209 (N_209,In_155,In_467);
xor U210 (N_210,In_572,In_481);
or U211 (N_211,In_430,In_210);
and U212 (N_212,In_856,In_200);
nand U213 (N_213,In_686,In_469);
or U214 (N_214,In_642,In_796);
and U215 (N_215,In_11,In_992);
or U216 (N_216,In_571,In_271);
and U217 (N_217,In_147,In_816);
and U218 (N_218,In_407,In_234);
nand U219 (N_219,In_690,In_771);
and U220 (N_220,In_724,In_579);
and U221 (N_221,In_935,In_842);
or U222 (N_222,In_444,In_767);
nor U223 (N_223,In_606,In_827);
and U224 (N_224,In_149,In_590);
and U225 (N_225,In_492,In_427);
nand U226 (N_226,In_273,In_456);
and U227 (N_227,In_589,In_299);
and U228 (N_228,In_283,In_450);
or U229 (N_229,In_397,In_458);
nand U230 (N_230,In_192,In_543);
or U231 (N_231,In_660,In_566);
and U232 (N_232,In_575,In_653);
nand U233 (N_233,In_81,In_256);
nor U234 (N_234,In_157,In_663);
nand U235 (N_235,In_286,In_784);
nand U236 (N_236,In_153,In_280);
and U237 (N_237,In_711,In_565);
and U238 (N_238,In_674,In_498);
nand U239 (N_239,In_844,In_254);
nand U240 (N_240,In_116,In_384);
nand U241 (N_241,In_389,In_128);
and U242 (N_242,In_551,In_238);
or U243 (N_243,In_569,In_354);
nand U244 (N_244,In_828,In_534);
or U245 (N_245,In_576,In_822);
nor U246 (N_246,In_894,In_228);
xnor U247 (N_247,In_560,In_759);
xnor U248 (N_248,In_372,In_821);
xnor U249 (N_249,In_898,In_127);
and U250 (N_250,In_139,In_726);
and U251 (N_251,In_463,In_975);
or U252 (N_252,In_739,In_622);
and U253 (N_253,In_144,In_875);
or U254 (N_254,In_419,In_777);
or U255 (N_255,In_466,In_855);
or U256 (N_256,In_870,In_623);
nor U257 (N_257,In_826,In_930);
or U258 (N_258,In_683,In_428);
and U259 (N_259,In_994,In_412);
or U260 (N_260,In_740,In_265);
and U261 (N_261,In_236,In_916);
nor U262 (N_262,In_439,In_670);
nand U263 (N_263,In_325,In_750);
nand U264 (N_264,In_786,In_504);
or U265 (N_265,In_40,In_745);
nand U266 (N_266,In_202,In_190);
nand U267 (N_267,In_616,In_884);
or U268 (N_268,In_142,In_978);
and U269 (N_269,In_840,In_634);
nor U270 (N_270,In_956,In_44);
or U271 (N_271,In_524,In_422);
nand U272 (N_272,In_718,In_433);
and U273 (N_273,In_919,In_129);
or U274 (N_274,In_864,In_490);
nand U275 (N_275,In_49,In_343);
nand U276 (N_276,In_737,In_112);
and U277 (N_277,In_904,In_715);
or U278 (N_278,In_748,In_885);
or U279 (N_279,In_719,In_244);
nor U280 (N_280,In_680,In_462);
nor U281 (N_281,In_263,In_52);
and U282 (N_282,In_549,In_229);
or U283 (N_283,In_948,In_241);
nor U284 (N_284,In_675,In_115);
nor U285 (N_285,In_792,In_68);
nor U286 (N_286,In_599,In_43);
nand U287 (N_287,In_892,In_251);
and U288 (N_288,In_262,In_791);
and U289 (N_289,In_126,In_887);
nand U290 (N_290,In_494,In_746);
nor U291 (N_291,In_294,In_802);
and U292 (N_292,In_561,In_730);
or U293 (N_293,In_963,In_95);
nor U294 (N_294,In_772,In_991);
or U295 (N_295,In_853,In_897);
nor U296 (N_296,In_627,In_891);
and U297 (N_297,In_973,In_913);
and U298 (N_298,In_896,In_300);
nand U299 (N_299,In_39,In_922);
nand U300 (N_300,In_762,In_12);
or U301 (N_301,In_438,In_755);
and U302 (N_302,In_282,In_368);
or U303 (N_303,In_608,In_408);
nor U304 (N_304,In_253,In_693);
nand U305 (N_305,In_48,In_743);
or U306 (N_306,In_785,In_505);
and U307 (N_307,In_482,In_644);
nor U308 (N_308,In_689,In_212);
or U309 (N_309,In_381,In_53);
xnor U310 (N_310,In_527,In_988);
nand U311 (N_311,In_484,In_140);
nor U312 (N_312,In_448,In_485);
nor U313 (N_313,In_537,In_255);
and U314 (N_314,In_509,In_311);
nor U315 (N_315,In_990,In_36);
and U316 (N_316,In_497,In_609);
nor U317 (N_317,In_376,In_881);
nor U318 (N_318,In_495,In_338);
nand U319 (N_319,In_111,In_230);
and U320 (N_320,In_592,In_511);
or U321 (N_321,In_758,In_62);
nor U322 (N_322,In_810,In_578);
or U323 (N_323,In_521,In_514);
nand U324 (N_324,In_117,In_535);
nand U325 (N_325,In_45,In_432);
nor U326 (N_326,In_603,In_20);
and U327 (N_327,In_797,In_668);
nor U328 (N_328,In_175,In_910);
nor U329 (N_329,In_633,In_203);
nor U330 (N_330,In_168,In_512);
nand U331 (N_331,In_138,In_405);
nor U332 (N_332,In_440,In_665);
or U333 (N_333,In_765,In_208);
or U334 (N_334,In_29,In_751);
nor U335 (N_335,In_291,In_30);
nand U336 (N_336,In_287,In_474);
and U337 (N_337,In_636,In_123);
and U338 (N_338,In_34,In_493);
and U339 (N_339,In_403,In_657);
nor U340 (N_340,In_207,In_365);
and U341 (N_341,In_685,In_999);
nor U342 (N_342,In_119,In_781);
and U343 (N_343,In_666,In_638);
nand U344 (N_344,In_413,In_249);
nor U345 (N_345,In_252,In_798);
and U346 (N_346,In_259,In_264);
nand U347 (N_347,In_678,In_426);
nand U348 (N_348,In_314,In_315);
nand U349 (N_349,In_418,In_845);
or U350 (N_350,In_90,In_567);
and U351 (N_351,In_757,In_851);
nor U352 (N_352,In_37,In_316);
nand U353 (N_353,In_649,In_380);
and U354 (N_354,In_292,In_302);
or U355 (N_355,In_952,In_362);
or U356 (N_356,In_890,In_866);
nand U357 (N_357,In_105,In_950);
nand U358 (N_358,In_830,In_435);
nand U359 (N_359,In_295,In_934);
or U360 (N_360,In_242,In_677);
nand U361 (N_361,In_776,In_766);
nor U362 (N_362,In_232,In_525);
or U363 (N_363,In_940,In_370);
nor U364 (N_364,In_73,In_120);
and U365 (N_365,In_732,In_385);
nand U366 (N_366,In_290,In_630);
and U367 (N_367,In_334,In_778);
or U368 (N_368,In_71,In_199);
or U369 (N_369,In_847,In_908);
or U370 (N_370,In_854,In_267);
nor U371 (N_371,In_862,In_197);
nor U372 (N_372,In_303,In_900);
xor U373 (N_373,In_983,In_313);
xnor U374 (N_374,In_601,In_304);
and U375 (N_375,In_526,In_360);
and U376 (N_376,In_74,In_124);
nand U377 (N_377,In_629,In_323);
nand U378 (N_378,In_18,In_877);
or U379 (N_379,In_387,In_284);
nand U380 (N_380,In_28,In_86);
nor U381 (N_381,In_156,In_5);
nor U382 (N_382,In_350,In_471);
and U383 (N_383,In_134,In_869);
nand U384 (N_384,In_449,In_308);
nor U385 (N_385,In_457,In_932);
nor U386 (N_386,In_597,In_635);
nor U387 (N_387,In_570,In_196);
nand U388 (N_388,In_154,In_78);
or U389 (N_389,In_473,In_417);
xnor U390 (N_390,In_545,In_943);
and U391 (N_391,In_707,In_22);
or U392 (N_392,In_54,In_790);
and U393 (N_393,In_761,In_553);
nand U394 (N_394,In_734,In_233);
xnor U395 (N_395,In_60,In_708);
nand U396 (N_396,In_88,In_538);
or U397 (N_397,In_411,In_832);
or U398 (N_398,In_520,In_833);
nand U399 (N_399,In_662,In_479);
nor U400 (N_400,In_835,In_453);
nand U401 (N_401,In_118,In_364);
and U402 (N_402,In_911,In_483);
and U403 (N_403,In_582,In_813);
nand U404 (N_404,In_180,In_352);
and U405 (N_405,In_173,In_933);
nor U406 (N_406,In_83,In_927);
nor U407 (N_407,In_340,In_472);
or U408 (N_408,In_867,In_503);
or U409 (N_409,In_839,In_359);
and U410 (N_410,In_373,In_620);
xor U411 (N_411,In_640,In_699);
nand U412 (N_412,In_80,In_274);
nand U413 (N_413,In_122,In_278);
and U414 (N_414,In_641,In_931);
and U415 (N_415,In_905,In_929);
and U416 (N_416,In_194,In_65);
nand U417 (N_417,In_66,In_136);
and U418 (N_418,In_125,In_215);
or U419 (N_419,In_843,In_568);
nor U420 (N_420,In_775,In_452);
and U421 (N_421,In_46,In_809);
nand U422 (N_422,In_728,In_446);
nand U423 (N_423,In_459,In_696);
nand U424 (N_424,In_859,In_961);
nand U425 (N_425,In_158,In_178);
nor U426 (N_426,In_652,In_31);
and U427 (N_427,In_424,In_289);
and U428 (N_428,In_121,In_400);
and U429 (N_429,In_415,In_874);
and U430 (N_430,In_522,In_664);
nor U431 (N_431,In_176,In_789);
nor U432 (N_432,In_793,In_906);
nand U433 (N_433,In_401,In_981);
nor U434 (N_434,In_398,In_378);
nand U435 (N_435,In_681,In_544);
nor U436 (N_436,In_339,In_488);
nand U437 (N_437,In_530,In_557);
nand U438 (N_438,In_688,In_554);
nor U439 (N_439,In_717,In_390);
nand U440 (N_440,In_651,In_995);
nand U441 (N_441,In_293,In_801);
and U442 (N_442,In_336,In_346);
nor U443 (N_443,In_513,In_486);
nand U444 (N_444,In_394,In_1);
or U445 (N_445,In_260,In_588);
and U446 (N_446,In_32,In_548);
and U447 (N_447,In_72,In_333);
nand U448 (N_448,In_825,In_984);
nand U449 (N_449,In_312,In_321);
nor U450 (N_450,In_834,In_351);
nor U451 (N_451,In_646,In_337);
nor U452 (N_452,In_223,In_164);
nand U453 (N_453,In_163,In_716);
and U454 (N_454,In_959,In_692);
nor U455 (N_455,In_861,In_181);
and U456 (N_456,In_942,In_91);
and U457 (N_457,In_552,In_969);
nand U458 (N_458,In_69,In_966);
and U459 (N_459,In_489,In_736);
or U460 (N_460,In_939,In_166);
or U461 (N_461,In_487,In_17);
nand U462 (N_462,In_146,In_441);
and U463 (N_463,In_613,In_811);
nor U464 (N_464,In_528,In_21);
nand U465 (N_465,In_676,In_580);
nand U466 (N_466,In_858,In_135);
nor U467 (N_467,In_901,In_661);
nor U468 (N_468,In_150,In_269);
nand U469 (N_469,In_100,In_476);
nand U470 (N_470,In_182,In_56);
nand U471 (N_471,In_968,In_246);
and U472 (N_472,In_423,In_937);
or U473 (N_473,In_720,In_631);
xor U474 (N_474,In_243,In_876);
xor U475 (N_475,In_868,In_562);
or U476 (N_476,In_706,In_697);
nand U477 (N_477,In_59,In_356);
and U478 (N_478,In_852,In_936);
and U479 (N_479,In_225,In_788);
nor U480 (N_480,In_709,In_169);
and U481 (N_481,In_143,In_964);
and U482 (N_482,In_67,In_738);
and U483 (N_483,In_550,In_58);
nand U484 (N_484,In_421,In_98);
nor U485 (N_485,In_103,In_533);
or U486 (N_486,In_502,In_625);
and U487 (N_487,In_206,In_542);
nand U488 (N_488,In_747,In_165);
nor U489 (N_489,In_752,In_836);
and U490 (N_490,In_235,In_106);
and U491 (N_491,In_912,In_741);
or U492 (N_492,In_247,In_167);
nor U493 (N_493,In_600,In_694);
and U494 (N_494,In_185,In_583);
nor U495 (N_495,In_783,In_794);
nand U496 (N_496,In_399,In_317);
nor U497 (N_497,In_954,In_102);
and U498 (N_498,In_547,In_383);
and U499 (N_499,In_753,In_319);
nand U500 (N_500,In_554,In_379);
and U501 (N_501,In_873,In_333);
or U502 (N_502,In_841,In_684);
nand U503 (N_503,In_294,In_343);
or U504 (N_504,In_538,In_350);
nand U505 (N_505,In_802,In_198);
and U506 (N_506,In_922,In_245);
or U507 (N_507,In_922,In_13);
nor U508 (N_508,In_571,In_281);
nor U509 (N_509,In_162,In_911);
and U510 (N_510,In_525,In_145);
or U511 (N_511,In_916,In_154);
nor U512 (N_512,In_391,In_32);
nand U513 (N_513,In_11,In_786);
or U514 (N_514,In_274,In_590);
nand U515 (N_515,In_450,In_356);
nor U516 (N_516,In_361,In_571);
or U517 (N_517,In_371,In_662);
or U518 (N_518,In_776,In_626);
nand U519 (N_519,In_614,In_328);
or U520 (N_520,In_924,In_745);
nor U521 (N_521,In_590,In_176);
or U522 (N_522,In_283,In_95);
or U523 (N_523,In_656,In_772);
nor U524 (N_524,In_998,In_762);
nand U525 (N_525,In_503,In_210);
nor U526 (N_526,In_386,In_972);
or U527 (N_527,In_546,In_21);
or U528 (N_528,In_498,In_244);
nand U529 (N_529,In_272,In_494);
and U530 (N_530,In_977,In_48);
and U531 (N_531,In_336,In_677);
or U532 (N_532,In_640,In_886);
and U533 (N_533,In_784,In_727);
or U534 (N_534,In_302,In_512);
or U535 (N_535,In_209,In_98);
and U536 (N_536,In_581,In_130);
or U537 (N_537,In_771,In_391);
and U538 (N_538,In_909,In_145);
nand U539 (N_539,In_123,In_946);
nor U540 (N_540,In_675,In_742);
and U541 (N_541,In_940,In_177);
and U542 (N_542,In_568,In_892);
or U543 (N_543,In_178,In_254);
or U544 (N_544,In_266,In_20);
or U545 (N_545,In_699,In_322);
or U546 (N_546,In_783,In_27);
nor U547 (N_547,In_278,In_631);
nand U548 (N_548,In_727,In_329);
nand U549 (N_549,In_358,In_334);
nand U550 (N_550,In_488,In_709);
and U551 (N_551,In_733,In_0);
nand U552 (N_552,In_688,In_221);
and U553 (N_553,In_967,In_483);
nand U554 (N_554,In_186,In_522);
nand U555 (N_555,In_211,In_938);
nor U556 (N_556,In_597,In_850);
nand U557 (N_557,In_950,In_349);
xnor U558 (N_558,In_567,In_929);
nand U559 (N_559,In_889,In_904);
or U560 (N_560,In_630,In_591);
nor U561 (N_561,In_978,In_371);
and U562 (N_562,In_238,In_924);
nor U563 (N_563,In_994,In_713);
nor U564 (N_564,In_3,In_370);
and U565 (N_565,In_262,In_448);
or U566 (N_566,In_367,In_360);
and U567 (N_567,In_655,In_704);
nand U568 (N_568,In_496,In_9);
nand U569 (N_569,In_139,In_955);
nor U570 (N_570,In_409,In_547);
nand U571 (N_571,In_127,In_684);
nor U572 (N_572,In_260,In_783);
and U573 (N_573,In_861,In_870);
nor U574 (N_574,In_160,In_366);
nand U575 (N_575,In_718,In_985);
or U576 (N_576,In_585,In_398);
and U577 (N_577,In_639,In_883);
nor U578 (N_578,In_93,In_177);
or U579 (N_579,In_145,In_316);
or U580 (N_580,In_405,In_949);
and U581 (N_581,In_708,In_746);
nand U582 (N_582,In_448,In_466);
nor U583 (N_583,In_274,In_440);
or U584 (N_584,In_417,In_436);
or U585 (N_585,In_92,In_445);
nor U586 (N_586,In_914,In_616);
nor U587 (N_587,In_361,In_950);
nand U588 (N_588,In_376,In_925);
nor U589 (N_589,In_663,In_891);
and U590 (N_590,In_829,In_702);
and U591 (N_591,In_254,In_684);
and U592 (N_592,In_984,In_319);
nand U593 (N_593,In_764,In_761);
nand U594 (N_594,In_535,In_600);
or U595 (N_595,In_277,In_770);
and U596 (N_596,In_994,In_460);
nor U597 (N_597,In_366,In_655);
nand U598 (N_598,In_894,In_377);
or U599 (N_599,In_639,In_557);
and U600 (N_600,In_494,In_45);
or U601 (N_601,In_619,In_662);
nor U602 (N_602,In_805,In_612);
or U603 (N_603,In_643,In_599);
or U604 (N_604,In_119,In_670);
nand U605 (N_605,In_9,In_897);
and U606 (N_606,In_276,In_312);
or U607 (N_607,In_952,In_995);
nor U608 (N_608,In_971,In_452);
nand U609 (N_609,In_689,In_274);
nor U610 (N_610,In_35,In_527);
nand U611 (N_611,In_764,In_865);
nor U612 (N_612,In_619,In_759);
nor U613 (N_613,In_238,In_158);
or U614 (N_614,In_389,In_293);
nand U615 (N_615,In_94,In_502);
or U616 (N_616,In_6,In_278);
or U617 (N_617,In_247,In_275);
nor U618 (N_618,In_205,In_588);
and U619 (N_619,In_819,In_48);
and U620 (N_620,In_956,In_439);
and U621 (N_621,In_843,In_897);
nand U622 (N_622,In_947,In_555);
or U623 (N_623,In_601,In_553);
nor U624 (N_624,In_150,In_54);
or U625 (N_625,In_878,In_161);
xnor U626 (N_626,In_272,In_835);
nor U627 (N_627,In_218,In_941);
nor U628 (N_628,In_589,In_341);
nand U629 (N_629,In_894,In_154);
or U630 (N_630,In_511,In_622);
nor U631 (N_631,In_679,In_328);
or U632 (N_632,In_337,In_548);
or U633 (N_633,In_305,In_329);
nor U634 (N_634,In_40,In_1);
or U635 (N_635,In_448,In_856);
or U636 (N_636,In_272,In_405);
and U637 (N_637,In_132,In_978);
or U638 (N_638,In_406,In_500);
or U639 (N_639,In_855,In_569);
nand U640 (N_640,In_64,In_418);
nor U641 (N_641,In_110,In_769);
or U642 (N_642,In_574,In_494);
or U643 (N_643,In_495,In_75);
nor U644 (N_644,In_755,In_450);
and U645 (N_645,In_628,In_643);
nand U646 (N_646,In_560,In_720);
nand U647 (N_647,In_812,In_344);
and U648 (N_648,In_224,In_515);
and U649 (N_649,In_334,In_747);
nor U650 (N_650,In_653,In_460);
nor U651 (N_651,In_981,In_194);
nor U652 (N_652,In_702,In_821);
nand U653 (N_653,In_104,In_771);
nor U654 (N_654,In_181,In_980);
nor U655 (N_655,In_693,In_870);
nand U656 (N_656,In_302,In_140);
nor U657 (N_657,In_126,In_46);
nand U658 (N_658,In_643,In_610);
nand U659 (N_659,In_231,In_720);
nor U660 (N_660,In_143,In_278);
nor U661 (N_661,In_110,In_825);
nor U662 (N_662,In_884,In_757);
or U663 (N_663,In_39,In_174);
nor U664 (N_664,In_895,In_545);
or U665 (N_665,In_842,In_194);
and U666 (N_666,In_576,In_535);
and U667 (N_667,In_553,In_830);
nor U668 (N_668,In_327,In_228);
nor U669 (N_669,In_33,In_71);
nand U670 (N_670,In_648,In_843);
or U671 (N_671,In_108,In_209);
and U672 (N_672,In_600,In_494);
nand U673 (N_673,In_641,In_469);
nor U674 (N_674,In_274,In_677);
nand U675 (N_675,In_46,In_928);
nor U676 (N_676,In_424,In_881);
and U677 (N_677,In_24,In_611);
xor U678 (N_678,In_158,In_943);
and U679 (N_679,In_422,In_989);
nand U680 (N_680,In_126,In_43);
or U681 (N_681,In_55,In_799);
or U682 (N_682,In_672,In_898);
nand U683 (N_683,In_160,In_522);
xor U684 (N_684,In_160,In_531);
nor U685 (N_685,In_579,In_525);
or U686 (N_686,In_502,In_197);
or U687 (N_687,In_618,In_545);
or U688 (N_688,In_554,In_102);
nand U689 (N_689,In_940,In_776);
and U690 (N_690,In_124,In_176);
and U691 (N_691,In_698,In_909);
and U692 (N_692,In_561,In_56);
or U693 (N_693,In_170,In_37);
nand U694 (N_694,In_996,In_562);
nand U695 (N_695,In_523,In_487);
and U696 (N_696,In_690,In_185);
or U697 (N_697,In_714,In_709);
or U698 (N_698,In_384,In_79);
nand U699 (N_699,In_392,In_327);
nand U700 (N_700,In_921,In_266);
xnor U701 (N_701,In_944,In_425);
or U702 (N_702,In_936,In_402);
and U703 (N_703,In_415,In_171);
or U704 (N_704,In_750,In_435);
nor U705 (N_705,In_182,In_198);
or U706 (N_706,In_865,In_105);
nand U707 (N_707,In_95,In_409);
and U708 (N_708,In_78,In_722);
nor U709 (N_709,In_748,In_201);
nor U710 (N_710,In_553,In_863);
or U711 (N_711,In_2,In_875);
nor U712 (N_712,In_541,In_327);
and U713 (N_713,In_215,In_831);
or U714 (N_714,In_768,In_761);
and U715 (N_715,In_84,In_302);
and U716 (N_716,In_395,In_713);
or U717 (N_717,In_395,In_303);
or U718 (N_718,In_195,In_604);
nand U719 (N_719,In_15,In_338);
nor U720 (N_720,In_93,In_448);
nor U721 (N_721,In_540,In_156);
nor U722 (N_722,In_695,In_894);
or U723 (N_723,In_407,In_277);
nand U724 (N_724,In_797,In_552);
and U725 (N_725,In_188,In_971);
and U726 (N_726,In_185,In_773);
nor U727 (N_727,In_664,In_595);
and U728 (N_728,In_825,In_556);
nor U729 (N_729,In_956,In_831);
nand U730 (N_730,In_980,In_196);
nand U731 (N_731,In_252,In_51);
and U732 (N_732,In_121,In_861);
or U733 (N_733,In_483,In_265);
and U734 (N_734,In_37,In_280);
nand U735 (N_735,In_872,In_171);
nor U736 (N_736,In_221,In_655);
and U737 (N_737,In_862,In_107);
or U738 (N_738,In_92,In_208);
nor U739 (N_739,In_500,In_20);
or U740 (N_740,In_155,In_121);
and U741 (N_741,In_233,In_898);
or U742 (N_742,In_543,In_571);
and U743 (N_743,In_947,In_303);
nand U744 (N_744,In_674,In_172);
or U745 (N_745,In_280,In_904);
nand U746 (N_746,In_1,In_780);
or U747 (N_747,In_528,In_84);
or U748 (N_748,In_841,In_168);
or U749 (N_749,In_726,In_721);
nand U750 (N_750,In_341,In_70);
or U751 (N_751,In_437,In_681);
or U752 (N_752,In_809,In_440);
nor U753 (N_753,In_804,In_406);
or U754 (N_754,In_374,In_64);
nor U755 (N_755,In_874,In_69);
nor U756 (N_756,In_667,In_91);
or U757 (N_757,In_231,In_841);
and U758 (N_758,In_426,In_481);
nand U759 (N_759,In_316,In_374);
nor U760 (N_760,In_458,In_441);
nand U761 (N_761,In_372,In_123);
or U762 (N_762,In_817,In_399);
nand U763 (N_763,In_526,In_563);
and U764 (N_764,In_515,In_514);
or U765 (N_765,In_24,In_160);
nor U766 (N_766,In_866,In_429);
and U767 (N_767,In_460,In_896);
nor U768 (N_768,In_958,In_181);
and U769 (N_769,In_266,In_884);
nor U770 (N_770,In_784,In_765);
nor U771 (N_771,In_369,In_303);
or U772 (N_772,In_286,In_527);
nand U773 (N_773,In_393,In_741);
and U774 (N_774,In_939,In_5);
nand U775 (N_775,In_940,In_427);
or U776 (N_776,In_118,In_695);
or U777 (N_777,In_816,In_963);
nor U778 (N_778,In_54,In_182);
nand U779 (N_779,In_905,In_78);
or U780 (N_780,In_157,In_260);
and U781 (N_781,In_85,In_860);
nand U782 (N_782,In_305,In_776);
nand U783 (N_783,In_28,In_503);
and U784 (N_784,In_210,In_984);
nor U785 (N_785,In_146,In_771);
or U786 (N_786,In_310,In_798);
nand U787 (N_787,In_789,In_267);
or U788 (N_788,In_976,In_327);
nor U789 (N_789,In_883,In_217);
nor U790 (N_790,In_931,In_654);
or U791 (N_791,In_320,In_180);
nand U792 (N_792,In_763,In_301);
nand U793 (N_793,In_658,In_655);
nand U794 (N_794,In_553,In_488);
nor U795 (N_795,In_211,In_101);
or U796 (N_796,In_434,In_235);
and U797 (N_797,In_950,In_967);
nand U798 (N_798,In_781,In_108);
nand U799 (N_799,In_462,In_316);
or U800 (N_800,In_105,In_389);
nor U801 (N_801,In_601,In_556);
or U802 (N_802,In_950,In_273);
nor U803 (N_803,In_836,In_453);
nand U804 (N_804,In_742,In_884);
nand U805 (N_805,In_975,In_519);
and U806 (N_806,In_955,In_409);
and U807 (N_807,In_366,In_437);
and U808 (N_808,In_877,In_291);
nand U809 (N_809,In_279,In_894);
nor U810 (N_810,In_264,In_101);
nor U811 (N_811,In_667,In_440);
nand U812 (N_812,In_130,In_778);
nand U813 (N_813,In_90,In_304);
nand U814 (N_814,In_839,In_903);
or U815 (N_815,In_108,In_605);
nor U816 (N_816,In_181,In_216);
or U817 (N_817,In_802,In_947);
nor U818 (N_818,In_344,In_578);
nor U819 (N_819,In_730,In_396);
nor U820 (N_820,In_821,In_80);
nor U821 (N_821,In_198,In_880);
and U822 (N_822,In_122,In_372);
and U823 (N_823,In_569,In_460);
or U824 (N_824,In_762,In_323);
nor U825 (N_825,In_39,In_342);
nand U826 (N_826,In_146,In_750);
or U827 (N_827,In_464,In_713);
nand U828 (N_828,In_209,In_656);
nand U829 (N_829,In_258,In_530);
or U830 (N_830,In_684,In_405);
nand U831 (N_831,In_838,In_771);
nand U832 (N_832,In_405,In_831);
nand U833 (N_833,In_520,In_561);
and U834 (N_834,In_696,In_510);
nand U835 (N_835,In_196,In_566);
and U836 (N_836,In_481,In_347);
nor U837 (N_837,In_273,In_583);
or U838 (N_838,In_946,In_965);
or U839 (N_839,In_570,In_632);
nor U840 (N_840,In_756,In_402);
or U841 (N_841,In_267,In_371);
and U842 (N_842,In_391,In_348);
or U843 (N_843,In_794,In_909);
and U844 (N_844,In_752,In_391);
nor U845 (N_845,In_148,In_540);
or U846 (N_846,In_493,In_18);
nor U847 (N_847,In_6,In_920);
or U848 (N_848,In_658,In_507);
and U849 (N_849,In_140,In_817);
xnor U850 (N_850,In_855,In_317);
nand U851 (N_851,In_916,In_680);
and U852 (N_852,In_442,In_40);
nor U853 (N_853,In_427,In_985);
nand U854 (N_854,In_19,In_289);
nor U855 (N_855,In_237,In_61);
and U856 (N_856,In_851,In_959);
nor U857 (N_857,In_239,In_110);
nor U858 (N_858,In_981,In_466);
or U859 (N_859,In_658,In_306);
nor U860 (N_860,In_679,In_464);
nor U861 (N_861,In_226,In_74);
nand U862 (N_862,In_55,In_575);
nor U863 (N_863,In_811,In_5);
or U864 (N_864,In_997,In_118);
and U865 (N_865,In_270,In_849);
and U866 (N_866,In_741,In_943);
or U867 (N_867,In_277,In_185);
nor U868 (N_868,In_900,In_454);
nand U869 (N_869,In_86,In_737);
or U870 (N_870,In_165,In_926);
or U871 (N_871,In_321,In_6);
or U872 (N_872,In_82,In_89);
or U873 (N_873,In_321,In_884);
or U874 (N_874,In_919,In_720);
nor U875 (N_875,In_298,In_829);
nor U876 (N_876,In_770,In_371);
and U877 (N_877,In_609,In_30);
nor U878 (N_878,In_399,In_99);
nor U879 (N_879,In_697,In_781);
or U880 (N_880,In_579,In_388);
nand U881 (N_881,In_48,In_194);
and U882 (N_882,In_221,In_302);
or U883 (N_883,In_873,In_169);
nand U884 (N_884,In_963,In_256);
and U885 (N_885,In_175,In_234);
and U886 (N_886,In_419,In_820);
nor U887 (N_887,In_975,In_191);
or U888 (N_888,In_950,In_397);
or U889 (N_889,In_628,In_315);
nor U890 (N_890,In_390,In_96);
or U891 (N_891,In_349,In_895);
or U892 (N_892,In_263,In_723);
nand U893 (N_893,In_83,In_436);
nand U894 (N_894,In_529,In_977);
nand U895 (N_895,In_171,In_957);
and U896 (N_896,In_894,In_216);
nand U897 (N_897,In_558,In_480);
xor U898 (N_898,In_498,In_200);
nand U899 (N_899,In_334,In_679);
and U900 (N_900,In_949,In_679);
nor U901 (N_901,In_64,In_595);
nand U902 (N_902,In_684,In_92);
nor U903 (N_903,In_53,In_90);
nand U904 (N_904,In_441,In_361);
nor U905 (N_905,In_155,In_58);
nand U906 (N_906,In_371,In_184);
xor U907 (N_907,In_58,In_715);
nand U908 (N_908,In_919,In_39);
nand U909 (N_909,In_485,In_47);
and U910 (N_910,In_523,In_558);
or U911 (N_911,In_707,In_631);
or U912 (N_912,In_46,In_244);
nor U913 (N_913,In_184,In_203);
nor U914 (N_914,In_881,In_667);
and U915 (N_915,In_268,In_963);
and U916 (N_916,In_168,In_181);
and U917 (N_917,In_587,In_753);
xor U918 (N_918,In_403,In_451);
and U919 (N_919,In_936,In_124);
nor U920 (N_920,In_107,In_857);
and U921 (N_921,In_776,In_750);
and U922 (N_922,In_700,In_647);
nor U923 (N_923,In_636,In_659);
nor U924 (N_924,In_392,In_616);
nor U925 (N_925,In_864,In_604);
nand U926 (N_926,In_38,In_835);
nand U927 (N_927,In_102,In_281);
nor U928 (N_928,In_752,In_600);
and U929 (N_929,In_6,In_887);
nor U930 (N_930,In_23,In_382);
or U931 (N_931,In_972,In_704);
or U932 (N_932,In_322,In_409);
nor U933 (N_933,In_315,In_495);
or U934 (N_934,In_862,In_224);
nand U935 (N_935,In_22,In_393);
nor U936 (N_936,In_64,In_834);
nand U937 (N_937,In_754,In_174);
nand U938 (N_938,In_31,In_490);
and U939 (N_939,In_276,In_381);
and U940 (N_940,In_302,In_458);
and U941 (N_941,In_77,In_731);
and U942 (N_942,In_453,In_623);
and U943 (N_943,In_207,In_626);
or U944 (N_944,In_226,In_60);
nand U945 (N_945,In_451,In_443);
nor U946 (N_946,In_475,In_160);
and U947 (N_947,In_907,In_468);
or U948 (N_948,In_487,In_622);
or U949 (N_949,In_695,In_382);
nor U950 (N_950,In_376,In_654);
and U951 (N_951,In_317,In_639);
or U952 (N_952,In_293,In_891);
and U953 (N_953,In_527,In_324);
nor U954 (N_954,In_632,In_57);
nor U955 (N_955,In_880,In_255);
xnor U956 (N_956,In_978,In_955);
nand U957 (N_957,In_344,In_424);
nand U958 (N_958,In_261,In_330);
nor U959 (N_959,In_4,In_721);
nand U960 (N_960,In_21,In_581);
nand U961 (N_961,In_15,In_154);
nor U962 (N_962,In_300,In_441);
or U963 (N_963,In_992,In_122);
nor U964 (N_964,In_88,In_589);
nor U965 (N_965,In_978,In_31);
or U966 (N_966,In_142,In_746);
nor U967 (N_967,In_942,In_252);
nand U968 (N_968,In_778,In_518);
and U969 (N_969,In_276,In_9);
nand U970 (N_970,In_639,In_394);
and U971 (N_971,In_805,In_695);
nor U972 (N_972,In_324,In_345);
nor U973 (N_973,In_41,In_714);
or U974 (N_974,In_612,In_273);
nor U975 (N_975,In_610,In_815);
nor U976 (N_976,In_766,In_484);
nor U977 (N_977,In_78,In_298);
nand U978 (N_978,In_52,In_959);
and U979 (N_979,In_642,In_41);
nand U980 (N_980,In_480,In_821);
nand U981 (N_981,In_561,In_804);
nand U982 (N_982,In_51,In_139);
nor U983 (N_983,In_801,In_121);
and U984 (N_984,In_400,In_770);
or U985 (N_985,In_470,In_130);
nor U986 (N_986,In_980,In_430);
nand U987 (N_987,In_70,In_692);
nor U988 (N_988,In_200,In_795);
and U989 (N_989,In_295,In_355);
or U990 (N_990,In_439,In_995);
or U991 (N_991,In_462,In_434);
nand U992 (N_992,In_582,In_817);
and U993 (N_993,In_659,In_391);
or U994 (N_994,In_377,In_225);
nor U995 (N_995,In_490,In_875);
or U996 (N_996,In_835,In_957);
nand U997 (N_997,In_791,In_200);
nand U998 (N_998,In_652,In_88);
xnor U999 (N_999,In_826,In_909);
nand U1000 (N_1000,N_628,N_39);
nand U1001 (N_1001,N_639,N_836);
nor U1002 (N_1002,N_11,N_833);
nor U1003 (N_1003,N_436,N_122);
nand U1004 (N_1004,N_502,N_379);
nor U1005 (N_1005,N_848,N_160);
nor U1006 (N_1006,N_205,N_685);
nand U1007 (N_1007,N_821,N_13);
or U1008 (N_1008,N_906,N_267);
nor U1009 (N_1009,N_559,N_66);
nor U1010 (N_1010,N_359,N_940);
nor U1011 (N_1011,N_9,N_18);
nand U1012 (N_1012,N_979,N_963);
or U1013 (N_1013,N_869,N_218);
nand U1014 (N_1014,N_786,N_925);
and U1015 (N_1015,N_670,N_966);
nand U1016 (N_1016,N_686,N_866);
nor U1017 (N_1017,N_677,N_634);
nor U1018 (N_1018,N_624,N_131);
nand U1019 (N_1019,N_315,N_666);
or U1020 (N_1020,N_765,N_934);
or U1021 (N_1021,N_88,N_95);
nand U1022 (N_1022,N_87,N_727);
nor U1023 (N_1023,N_290,N_286);
or U1024 (N_1024,N_907,N_215);
or U1025 (N_1025,N_923,N_976);
nor U1026 (N_1026,N_690,N_544);
and U1027 (N_1027,N_945,N_737);
and U1028 (N_1028,N_785,N_431);
and U1029 (N_1029,N_904,N_266);
nor U1030 (N_1030,N_611,N_667);
nor U1031 (N_1031,N_949,N_76);
nor U1032 (N_1032,N_481,N_213);
or U1033 (N_1033,N_437,N_256);
and U1034 (N_1034,N_485,N_679);
and U1035 (N_1035,N_107,N_752);
nand U1036 (N_1036,N_393,N_135);
nand U1037 (N_1037,N_284,N_23);
and U1038 (N_1038,N_239,N_441);
or U1039 (N_1039,N_159,N_440);
nand U1040 (N_1040,N_568,N_506);
or U1041 (N_1041,N_369,N_692);
or U1042 (N_1042,N_96,N_19);
nand U1043 (N_1043,N_10,N_226);
nand U1044 (N_1044,N_45,N_199);
or U1045 (N_1045,N_178,N_227);
or U1046 (N_1046,N_989,N_987);
nor U1047 (N_1047,N_109,N_551);
nor U1048 (N_1048,N_442,N_162);
nor U1049 (N_1049,N_116,N_521);
nand U1050 (N_1050,N_416,N_926);
or U1051 (N_1051,N_224,N_15);
and U1052 (N_1052,N_222,N_274);
nand U1053 (N_1053,N_420,N_554);
nor U1054 (N_1054,N_905,N_853);
nand U1055 (N_1055,N_860,N_563);
or U1056 (N_1056,N_54,N_422);
and U1057 (N_1057,N_151,N_826);
and U1058 (N_1058,N_655,N_358);
or U1059 (N_1059,N_599,N_172);
nand U1060 (N_1060,N_457,N_443);
nand U1061 (N_1061,N_731,N_129);
nor U1062 (N_1062,N_922,N_936);
or U1063 (N_1063,N_540,N_591);
nor U1064 (N_1064,N_982,N_852);
and U1065 (N_1065,N_248,N_47);
and U1066 (N_1066,N_154,N_220);
nand U1067 (N_1067,N_492,N_360);
xnor U1068 (N_1068,N_748,N_813);
and U1069 (N_1069,N_430,N_627);
nand U1070 (N_1070,N_103,N_769);
or U1071 (N_1071,N_944,N_721);
or U1072 (N_1072,N_807,N_478);
nand U1073 (N_1073,N_29,N_38);
and U1074 (N_1074,N_520,N_604);
nor U1075 (N_1075,N_217,N_295);
nand U1076 (N_1076,N_503,N_687);
nand U1077 (N_1077,N_317,N_337);
nor U1078 (N_1078,N_75,N_454);
nor U1079 (N_1079,N_307,N_48);
and U1080 (N_1080,N_703,N_52);
nand U1081 (N_1081,N_78,N_288);
and U1082 (N_1082,N_528,N_743);
nand U1083 (N_1083,N_375,N_212);
and U1084 (N_1084,N_602,N_228);
or U1085 (N_1085,N_125,N_55);
and U1086 (N_1086,N_313,N_241);
nand U1087 (N_1087,N_827,N_582);
and U1088 (N_1088,N_882,N_383);
nor U1089 (N_1089,N_726,N_872);
or U1090 (N_1090,N_581,N_754);
nor U1091 (N_1091,N_879,N_252);
nor U1092 (N_1092,N_365,N_497);
or U1093 (N_1093,N_179,N_428);
nand U1094 (N_1094,N_838,N_883);
nand U1095 (N_1095,N_928,N_354);
nor U1096 (N_1096,N_186,N_58);
or U1097 (N_1097,N_712,N_778);
or U1098 (N_1098,N_631,N_353);
nor U1099 (N_1099,N_406,N_722);
nand U1100 (N_1100,N_641,N_49);
xnor U1101 (N_1101,N_493,N_7);
or U1102 (N_1102,N_347,N_930);
and U1103 (N_1103,N_865,N_501);
and U1104 (N_1104,N_148,N_128);
nor U1105 (N_1105,N_387,N_522);
or U1106 (N_1106,N_255,N_298);
and U1107 (N_1107,N_272,N_411);
nor U1108 (N_1108,N_847,N_401);
or U1109 (N_1109,N_204,N_601);
and U1110 (N_1110,N_890,N_291);
and U1111 (N_1111,N_843,N_849);
nor U1112 (N_1112,N_856,N_410);
nand U1113 (N_1113,N_665,N_450);
or U1114 (N_1114,N_216,N_796);
nand U1115 (N_1115,N_706,N_757);
and U1116 (N_1116,N_888,N_499);
or U1117 (N_1117,N_157,N_874);
nor U1118 (N_1118,N_962,N_133);
and U1119 (N_1119,N_746,N_57);
nor U1120 (N_1120,N_293,N_759);
nor U1121 (N_1121,N_788,N_278);
nor U1122 (N_1122,N_978,N_306);
nand U1123 (N_1123,N_142,N_418);
nor U1124 (N_1124,N_181,N_814);
nand U1125 (N_1125,N_645,N_539);
nor U1126 (N_1126,N_183,N_445);
nand U1127 (N_1127,N_483,N_768);
nand U1128 (N_1128,N_237,N_577);
nor U1129 (N_1129,N_793,N_408);
and U1130 (N_1130,N_767,N_968);
and U1131 (N_1131,N_834,N_913);
or U1132 (N_1132,N_388,N_439);
or U1133 (N_1133,N_973,N_123);
and U1134 (N_1134,N_89,N_893);
and U1135 (N_1135,N_891,N_651);
or U1136 (N_1136,N_514,N_211);
nor U1137 (N_1137,N_894,N_117);
or U1138 (N_1138,N_189,N_854);
and U1139 (N_1139,N_952,N_857);
or U1140 (N_1140,N_247,N_878);
nor U1141 (N_1141,N_36,N_802);
nand U1142 (N_1142,N_429,N_876);
or U1143 (N_1143,N_158,N_363);
nand U1144 (N_1144,N_772,N_305);
nor U1145 (N_1145,N_828,N_386);
or U1146 (N_1146,N_127,N_482);
and U1147 (N_1147,N_791,N_592);
nand U1148 (N_1148,N_68,N_467);
nand U1149 (N_1149,N_194,N_578);
nand U1150 (N_1150,N_661,N_993);
or U1151 (N_1151,N_161,N_565);
nand U1152 (N_1152,N_287,N_709);
or U1153 (N_1153,N_112,N_281);
or U1154 (N_1154,N_632,N_794);
nor U1155 (N_1155,N_986,N_996);
and U1156 (N_1156,N_822,N_955);
nand U1157 (N_1157,N_877,N_115);
or U1158 (N_1158,N_536,N_322);
or U1159 (N_1159,N_53,N_658);
nand U1160 (N_1160,N_362,N_176);
nand U1161 (N_1161,N_63,N_673);
nor U1162 (N_1162,N_533,N_170);
nand U1163 (N_1163,N_951,N_150);
nor U1164 (N_1164,N_417,N_953);
or U1165 (N_1165,N_817,N_323);
and U1166 (N_1166,N_21,N_165);
nor U1167 (N_1167,N_163,N_110);
and U1168 (N_1168,N_310,N_924);
or U1169 (N_1169,N_719,N_855);
and U1170 (N_1170,N_72,N_447);
or U1171 (N_1171,N_702,N_262);
or U1172 (N_1172,N_377,N_808);
or U1173 (N_1173,N_803,N_552);
nand U1174 (N_1174,N_105,N_798);
nor U1175 (N_1175,N_22,N_421);
nand U1176 (N_1176,N_839,N_525);
or U1177 (N_1177,N_534,N_662);
nand U1178 (N_1178,N_321,N_766);
nand U1179 (N_1179,N_398,N_120);
nor U1180 (N_1180,N_397,N_261);
and U1181 (N_1181,N_1,N_456);
nand U1182 (N_1182,N_395,N_143);
nor U1183 (N_1183,N_932,N_371);
and U1184 (N_1184,N_473,N_268);
nor U1185 (N_1185,N_498,N_177);
or U1186 (N_1186,N_711,N_509);
nand U1187 (N_1187,N_364,N_476);
and U1188 (N_1188,N_167,N_964);
nand U1189 (N_1189,N_625,N_590);
nand U1190 (N_1190,N_954,N_688);
nand U1191 (N_1191,N_648,N_235);
or U1192 (N_1192,N_607,N_931);
nor U1193 (N_1193,N_713,N_106);
nand U1194 (N_1194,N_546,N_74);
or U1195 (N_1195,N_541,N_258);
or U1196 (N_1196,N_474,N_487);
and U1197 (N_1197,N_361,N_881);
nor U1198 (N_1198,N_250,N_100);
xnor U1199 (N_1199,N_640,N_196);
and U1200 (N_1200,N_804,N_663);
nand U1201 (N_1201,N_781,N_198);
or U1202 (N_1202,N_265,N_101);
and U1203 (N_1203,N_192,N_399);
nand U1204 (N_1204,N_618,N_895);
nor U1205 (N_1205,N_385,N_596);
nand U1206 (N_1206,N_468,N_407);
nand U1207 (N_1207,N_489,N_214);
or U1208 (N_1208,N_391,N_419);
nor U1209 (N_1209,N_914,N_779);
and U1210 (N_1210,N_466,N_553);
or U1211 (N_1211,N_620,N_776);
and U1212 (N_1212,N_728,N_336);
nand U1213 (N_1213,N_260,N_531);
and U1214 (N_1214,N_27,N_367);
nor U1215 (N_1215,N_392,N_691);
or U1216 (N_1216,N_998,N_919);
nor U1217 (N_1217,N_34,N_118);
nand U1218 (N_1218,N_294,N_619);
or U1219 (N_1219,N_571,N_969);
and U1220 (N_1220,N_654,N_980);
nor U1221 (N_1221,N_515,N_114);
nand U1222 (N_1222,N_630,N_696);
nor U1223 (N_1223,N_200,N_168);
nand U1224 (N_1224,N_755,N_909);
and U1225 (N_1225,N_974,N_508);
and U1226 (N_1226,N_787,N_332);
or U1227 (N_1227,N_842,N_585);
nor U1228 (N_1228,N_345,N_720);
or U1229 (N_1229,N_800,N_912);
or U1230 (N_1230,N_69,N_862);
nor U1231 (N_1231,N_961,N_868);
nand U1232 (N_1232,N_950,N_762);
nor U1233 (N_1233,N_734,N_432);
or U1234 (N_1234,N_622,N_761);
and U1235 (N_1235,N_887,N_609);
nor U1236 (N_1236,N_583,N_471);
and U1237 (N_1237,N_635,N_144);
or U1238 (N_1238,N_263,N_911);
nor U1239 (N_1239,N_579,N_257);
nand U1240 (N_1240,N_17,N_901);
or U1241 (N_1241,N_999,N_242);
and U1242 (N_1242,N_378,N_269);
and U1243 (N_1243,N_309,N_613);
nand U1244 (N_1244,N_270,N_46);
and U1245 (N_1245,N_108,N_749);
or U1246 (N_1246,N_435,N_863);
and U1247 (N_1247,N_104,N_524);
nand U1248 (N_1248,N_513,N_0);
nor U1249 (N_1249,N_773,N_575);
or U1250 (N_1250,N_134,N_403);
or U1251 (N_1251,N_285,N_636);
nor U1252 (N_1252,N_234,N_169);
and U1253 (N_1253,N_606,N_516);
or U1254 (N_1254,N_138,N_277);
nor U1255 (N_1255,N_97,N_561);
nand U1256 (N_1256,N_861,N_898);
nand U1257 (N_1257,N_699,N_615);
nor U1258 (N_1258,N_85,N_542);
and U1259 (N_1259,N_355,N_126);
nand U1260 (N_1260,N_529,N_320);
and U1261 (N_1261,N_94,N_844);
nand U1262 (N_1262,N_614,N_790);
nor U1263 (N_1263,N_535,N_245);
nand U1264 (N_1264,N_598,N_740);
or U1265 (N_1265,N_548,N_545);
or U1266 (N_1266,N_623,N_396);
or U1267 (N_1267,N_308,N_490);
and U1268 (N_1268,N_219,N_517);
nor U1269 (N_1269,N_929,N_136);
and U1270 (N_1270,N_652,N_899);
nand U1271 (N_1271,N_958,N_707);
or U1272 (N_1272,N_801,N_564);
nand U1273 (N_1273,N_405,N_26);
and U1274 (N_1274,N_916,N_736);
or U1275 (N_1275,N_992,N_956);
and U1276 (N_1276,N_25,N_747);
or U1277 (N_1277,N_62,N_983);
and U1278 (N_1278,N_694,N_433);
nor U1279 (N_1279,N_723,N_90);
or U1280 (N_1280,N_684,N_210);
nand U1281 (N_1281,N_562,N_130);
nand U1282 (N_1282,N_465,N_352);
nand U1283 (N_1283,N_608,N_689);
nor U1284 (N_1284,N_760,N_672);
nor U1285 (N_1285,N_209,N_185);
nand U1286 (N_1286,N_900,N_811);
nand U1287 (N_1287,N_995,N_59);
or U1288 (N_1288,N_98,N_469);
nor U1289 (N_1289,N_795,N_244);
or U1290 (N_1290,N_413,N_35);
nand U1291 (N_1291,N_593,N_453);
or U1292 (N_1292,N_264,N_920);
or U1293 (N_1293,N_381,N_557);
or U1294 (N_1294,N_682,N_4);
nand U1295 (N_1295,N_147,N_784);
or U1296 (N_1296,N_67,N_586);
nand U1297 (N_1297,N_589,N_460);
or U1298 (N_1298,N_570,N_427);
and U1299 (N_1299,N_948,N_424);
or U1300 (N_1300,N_897,N_572);
and U1301 (N_1301,N_50,N_946);
or U1302 (N_1302,N_400,N_240);
nor U1303 (N_1303,N_343,N_547);
and U1304 (N_1304,N_935,N_943);
and U1305 (N_1305,N_191,N_43);
nand U1306 (N_1306,N_941,N_942);
nand U1307 (N_1307,N_384,N_331);
or U1308 (N_1308,N_937,N_600);
or U1309 (N_1309,N_902,N_461);
nor U1310 (N_1310,N_65,N_864);
or U1311 (N_1311,N_567,N_455);
or U1312 (N_1312,N_915,N_296);
nor U1313 (N_1313,N_197,N_5);
nor U1314 (N_1314,N_149,N_64);
nand U1315 (N_1315,N_574,N_806);
nor U1316 (N_1316,N_201,N_647);
nand U1317 (N_1317,N_612,N_140);
and U1318 (N_1318,N_644,N_873);
and U1319 (N_1319,N_238,N_959);
or U1320 (N_1320,N_903,N_875);
and U1321 (N_1321,N_809,N_31);
and U1322 (N_1322,N_30,N_870);
nor U1323 (N_1323,N_289,N_605);
nor U1324 (N_1324,N_111,N_818);
nand U1325 (N_1325,N_51,N_965);
nand U1326 (N_1326,N_668,N_452);
nand U1327 (N_1327,N_921,N_304);
and U1328 (N_1328,N_820,N_300);
nor U1329 (N_1329,N_484,N_470);
nand U1330 (N_1330,N_349,N_616);
nor U1331 (N_1331,N_412,N_86);
nor U1332 (N_1332,N_374,N_346);
nand U1333 (N_1333,N_710,N_40);
or U1334 (N_1334,N_939,N_44);
nor U1335 (N_1335,N_664,N_629);
nor U1336 (N_1336,N_174,N_896);
or U1337 (N_1337,N_254,N_797);
nand U1338 (N_1338,N_947,N_376);
nand U1339 (N_1339,N_695,N_171);
nand U1340 (N_1340,N_889,N_576);
and U1341 (N_1341,N_549,N_423);
or U1342 (N_1342,N_84,N_325);
nor U1343 (N_1343,N_141,N_495);
nand U1344 (N_1344,N_560,N_193);
and U1345 (N_1345,N_253,N_225);
nand U1346 (N_1346,N_472,N_16);
nand U1347 (N_1347,N_782,N_146);
and U1348 (N_1348,N_338,N_425);
and U1349 (N_1349,N_693,N_988);
nand U1350 (N_1350,N_751,N_328);
nand U1351 (N_1351,N_326,N_595);
or U1352 (N_1352,N_569,N_649);
nor U1353 (N_1353,N_477,N_507);
nand U1354 (N_1354,N_372,N_741);
and U1355 (N_1355,N_80,N_273);
and U1356 (N_1356,N_335,N_550);
nor U1357 (N_1357,N_637,N_164);
and U1358 (N_1358,N_56,N_770);
nand U1359 (N_1359,N_137,N_166);
nor U1360 (N_1360,N_446,N_918);
nand U1361 (N_1361,N_566,N_28);
nand U1362 (N_1362,N_223,N_312);
or U1363 (N_1363,N_858,N_957);
nor U1364 (N_1364,N_348,N_230);
nor U1365 (N_1365,N_229,N_573);
nand U1366 (N_1366,N_275,N_207);
nand U1367 (N_1367,N_537,N_527);
nor U1368 (N_1368,N_837,N_971);
nand U1369 (N_1369,N_459,N_738);
and U1370 (N_1370,N_885,N_488);
nand U1371 (N_1371,N_173,N_587);
nor U1372 (N_1372,N_697,N_314);
or U1373 (N_1373,N_742,N_175);
nand U1374 (N_1374,N_886,N_208);
and U1375 (N_1375,N_816,N_825);
or U1376 (N_1376,N_610,N_633);
or U1377 (N_1377,N_333,N_319);
nand U1378 (N_1378,N_236,N_449);
or U1379 (N_1379,N_32,N_880);
nor U1380 (N_1380,N_835,N_145);
or U1381 (N_1381,N_132,N_917);
nand U1382 (N_1382,N_70,N_580);
or U1383 (N_1383,N_202,N_671);
and U1384 (N_1384,N_638,N_496);
nand U1385 (N_1385,N_14,N_511);
and U1386 (N_1386,N_783,N_71);
nor U1387 (N_1387,N_42,N_280);
and U1388 (N_1388,N_701,N_938);
nand U1389 (N_1389,N_404,N_927);
nand U1390 (N_1390,N_475,N_434);
or U1391 (N_1391,N_933,N_61);
nor U1392 (N_1392,N_715,N_500);
or U1393 (N_1393,N_735,N_93);
nor U1394 (N_1394,N_316,N_990);
nor U1395 (N_1395,N_342,N_233);
xnor U1396 (N_1396,N_845,N_155);
and U1397 (N_1397,N_780,N_908);
and U1398 (N_1398,N_152,N_538);
nand U1399 (N_1399,N_739,N_92);
or U1400 (N_1400,N_37,N_119);
and U1401 (N_1401,N_805,N_243);
or U1402 (N_1402,N_351,N_678);
and U1403 (N_1403,N_829,N_182);
or U1404 (N_1404,N_232,N_716);
and U1405 (N_1405,N_819,N_777);
nand U1406 (N_1406,N_674,N_732);
nand U1407 (N_1407,N_910,N_504);
nand U1408 (N_1408,N_657,N_659);
nor U1409 (N_1409,N_479,N_124);
or U1410 (N_1410,N_246,N_994);
or U1411 (N_1411,N_279,N_523);
and U1412 (N_1412,N_350,N_184);
or U1413 (N_1413,N_683,N_301);
and U1414 (N_1414,N_729,N_60);
or U1415 (N_1415,N_656,N_714);
nand U1416 (N_1416,N_486,N_518);
nor U1417 (N_1417,N_3,N_370);
or U1418 (N_1418,N_12,N_815);
nand U1419 (N_1419,N_775,N_390);
and U1420 (N_1420,N_444,N_789);
or U1421 (N_1421,N_708,N_519);
nand U1422 (N_1422,N_283,N_660);
and U1423 (N_1423,N_594,N_597);
or U1424 (N_1424,N_382,N_6);
nor U1425 (N_1425,N_967,N_646);
nor U1426 (N_1426,N_438,N_366);
or U1427 (N_1427,N_700,N_823);
or U1428 (N_1428,N_763,N_451);
nand U1429 (N_1429,N_356,N_249);
nor U1430 (N_1430,N_299,N_680);
and U1431 (N_1431,N_681,N_705);
or U1432 (N_1432,N_730,N_82);
nand U1433 (N_1433,N_330,N_841);
and U1434 (N_1434,N_532,N_512);
and U1435 (N_1435,N_744,N_415);
nand U1436 (N_1436,N_774,N_409);
nand U1437 (N_1437,N_745,N_324);
nor U1438 (N_1438,N_970,N_650);
and U1439 (N_1439,N_318,N_41);
nand U1440 (N_1440,N_840,N_792);
or U1441 (N_1441,N_458,N_389);
and U1442 (N_1442,N_303,N_311);
and U1443 (N_1443,N_448,N_846);
and U1444 (N_1444,N_764,N_187);
or U1445 (N_1445,N_33,N_394);
nor U1446 (N_1446,N_758,N_603);
nor U1447 (N_1447,N_676,N_892);
and U1448 (N_1448,N_530,N_83);
or U1449 (N_1449,N_505,N_251);
and U1450 (N_1450,N_156,N_344);
or U1451 (N_1451,N_81,N_724);
nand U1452 (N_1452,N_341,N_77);
nand U1453 (N_1453,N_494,N_91);
nor U1454 (N_1454,N_556,N_79);
and U1455 (N_1455,N_99,N_960);
nor U1456 (N_1456,N_491,N_981);
nor U1457 (N_1457,N_733,N_717);
nand U1458 (N_1458,N_972,N_113);
and U1459 (N_1459,N_139,N_368);
or U1460 (N_1460,N_334,N_188);
and U1461 (N_1461,N_675,N_510);
and U1462 (N_1462,N_884,N_753);
and U1463 (N_1463,N_850,N_831);
or U1464 (N_1464,N_339,N_292);
or U1465 (N_1465,N_121,N_297);
and U1466 (N_1466,N_463,N_756);
nor U1467 (N_1467,N_799,N_329);
or U1468 (N_1468,N_357,N_8);
nor U1469 (N_1469,N_867,N_812);
xnor U1470 (N_1470,N_543,N_203);
and U1471 (N_1471,N_669,N_621);
and U1472 (N_1472,N_997,N_584);
or U1473 (N_1473,N_975,N_871);
and U1474 (N_1474,N_373,N_588);
nor U1475 (N_1475,N_626,N_984);
nand U1476 (N_1476,N_327,N_985);
and U1477 (N_1477,N_259,N_221);
or U1478 (N_1478,N_698,N_771);
nor U1479 (N_1479,N_526,N_282);
nand U1480 (N_1480,N_653,N_750);
or U1481 (N_1481,N_73,N_231);
nor U1482 (N_1482,N_462,N_340);
or U1483 (N_1483,N_704,N_642);
xor U1484 (N_1484,N_276,N_830);
xor U1485 (N_1485,N_617,N_977);
or U1486 (N_1486,N_480,N_426);
and U1487 (N_1487,N_206,N_153);
and U1488 (N_1488,N_832,N_414);
or U1489 (N_1489,N_180,N_195);
nand U1490 (N_1490,N_810,N_555);
nor U1491 (N_1491,N_190,N_991);
and U1492 (N_1492,N_2,N_725);
nand U1493 (N_1493,N_718,N_24);
or U1494 (N_1494,N_380,N_102);
or U1495 (N_1495,N_558,N_824);
nand U1496 (N_1496,N_271,N_20);
nand U1497 (N_1497,N_464,N_643);
nand U1498 (N_1498,N_302,N_402);
and U1499 (N_1499,N_851,N_859);
nand U1500 (N_1500,N_251,N_376);
nand U1501 (N_1501,N_633,N_338);
nor U1502 (N_1502,N_264,N_624);
nand U1503 (N_1503,N_106,N_46);
nand U1504 (N_1504,N_453,N_134);
nor U1505 (N_1505,N_90,N_901);
and U1506 (N_1506,N_799,N_999);
and U1507 (N_1507,N_392,N_770);
and U1508 (N_1508,N_228,N_727);
and U1509 (N_1509,N_268,N_185);
or U1510 (N_1510,N_157,N_556);
nand U1511 (N_1511,N_555,N_612);
nor U1512 (N_1512,N_180,N_237);
or U1513 (N_1513,N_192,N_61);
and U1514 (N_1514,N_200,N_529);
and U1515 (N_1515,N_128,N_593);
nand U1516 (N_1516,N_263,N_497);
nor U1517 (N_1517,N_499,N_964);
or U1518 (N_1518,N_343,N_749);
nor U1519 (N_1519,N_204,N_281);
nor U1520 (N_1520,N_189,N_579);
and U1521 (N_1521,N_105,N_206);
nand U1522 (N_1522,N_919,N_159);
nand U1523 (N_1523,N_200,N_86);
nand U1524 (N_1524,N_282,N_385);
or U1525 (N_1525,N_198,N_525);
or U1526 (N_1526,N_945,N_125);
and U1527 (N_1527,N_310,N_926);
and U1528 (N_1528,N_799,N_770);
or U1529 (N_1529,N_138,N_912);
nor U1530 (N_1530,N_61,N_891);
nor U1531 (N_1531,N_762,N_640);
nand U1532 (N_1532,N_749,N_940);
and U1533 (N_1533,N_31,N_414);
nand U1534 (N_1534,N_565,N_417);
nand U1535 (N_1535,N_286,N_952);
xnor U1536 (N_1536,N_398,N_21);
or U1537 (N_1537,N_507,N_367);
and U1538 (N_1538,N_972,N_24);
or U1539 (N_1539,N_690,N_181);
nor U1540 (N_1540,N_749,N_413);
nor U1541 (N_1541,N_559,N_548);
nand U1542 (N_1542,N_288,N_625);
and U1543 (N_1543,N_456,N_264);
or U1544 (N_1544,N_386,N_955);
or U1545 (N_1545,N_782,N_585);
or U1546 (N_1546,N_291,N_748);
xnor U1547 (N_1547,N_381,N_422);
and U1548 (N_1548,N_735,N_238);
nand U1549 (N_1549,N_999,N_738);
nand U1550 (N_1550,N_107,N_437);
or U1551 (N_1551,N_508,N_925);
nand U1552 (N_1552,N_937,N_609);
nand U1553 (N_1553,N_866,N_580);
or U1554 (N_1554,N_141,N_937);
or U1555 (N_1555,N_230,N_370);
and U1556 (N_1556,N_789,N_373);
nor U1557 (N_1557,N_458,N_541);
nor U1558 (N_1558,N_472,N_603);
or U1559 (N_1559,N_112,N_441);
xnor U1560 (N_1560,N_127,N_564);
or U1561 (N_1561,N_875,N_538);
nor U1562 (N_1562,N_764,N_252);
nor U1563 (N_1563,N_194,N_493);
nand U1564 (N_1564,N_19,N_436);
and U1565 (N_1565,N_279,N_188);
or U1566 (N_1566,N_697,N_866);
or U1567 (N_1567,N_321,N_17);
nand U1568 (N_1568,N_998,N_394);
or U1569 (N_1569,N_827,N_194);
nor U1570 (N_1570,N_379,N_812);
nand U1571 (N_1571,N_715,N_294);
and U1572 (N_1572,N_854,N_847);
and U1573 (N_1573,N_100,N_710);
xnor U1574 (N_1574,N_630,N_546);
nand U1575 (N_1575,N_50,N_262);
or U1576 (N_1576,N_65,N_389);
nor U1577 (N_1577,N_991,N_328);
and U1578 (N_1578,N_933,N_164);
and U1579 (N_1579,N_460,N_452);
or U1580 (N_1580,N_51,N_129);
or U1581 (N_1581,N_294,N_585);
nand U1582 (N_1582,N_190,N_918);
nor U1583 (N_1583,N_828,N_448);
and U1584 (N_1584,N_67,N_574);
and U1585 (N_1585,N_196,N_239);
nor U1586 (N_1586,N_640,N_349);
and U1587 (N_1587,N_532,N_547);
or U1588 (N_1588,N_668,N_630);
xor U1589 (N_1589,N_229,N_305);
or U1590 (N_1590,N_770,N_339);
or U1591 (N_1591,N_933,N_350);
nand U1592 (N_1592,N_266,N_980);
nand U1593 (N_1593,N_924,N_159);
nor U1594 (N_1594,N_868,N_170);
or U1595 (N_1595,N_92,N_223);
or U1596 (N_1596,N_125,N_90);
and U1597 (N_1597,N_903,N_49);
or U1598 (N_1598,N_89,N_82);
and U1599 (N_1599,N_753,N_137);
nor U1600 (N_1600,N_268,N_137);
nand U1601 (N_1601,N_33,N_414);
nor U1602 (N_1602,N_790,N_92);
nor U1603 (N_1603,N_620,N_742);
nand U1604 (N_1604,N_651,N_358);
nand U1605 (N_1605,N_216,N_248);
or U1606 (N_1606,N_291,N_895);
and U1607 (N_1607,N_480,N_219);
nor U1608 (N_1608,N_668,N_369);
and U1609 (N_1609,N_926,N_971);
and U1610 (N_1610,N_92,N_163);
xor U1611 (N_1611,N_781,N_41);
or U1612 (N_1612,N_152,N_236);
nor U1613 (N_1613,N_681,N_143);
and U1614 (N_1614,N_80,N_402);
nor U1615 (N_1615,N_382,N_934);
nor U1616 (N_1616,N_114,N_557);
and U1617 (N_1617,N_921,N_268);
nor U1618 (N_1618,N_998,N_920);
nor U1619 (N_1619,N_258,N_622);
nor U1620 (N_1620,N_374,N_352);
and U1621 (N_1621,N_74,N_540);
and U1622 (N_1622,N_503,N_500);
or U1623 (N_1623,N_562,N_55);
or U1624 (N_1624,N_972,N_274);
nor U1625 (N_1625,N_380,N_410);
nand U1626 (N_1626,N_638,N_797);
nor U1627 (N_1627,N_431,N_79);
nor U1628 (N_1628,N_553,N_874);
and U1629 (N_1629,N_86,N_227);
nand U1630 (N_1630,N_138,N_862);
nand U1631 (N_1631,N_380,N_470);
or U1632 (N_1632,N_302,N_389);
or U1633 (N_1633,N_19,N_183);
and U1634 (N_1634,N_92,N_960);
xor U1635 (N_1635,N_873,N_428);
nor U1636 (N_1636,N_308,N_126);
nor U1637 (N_1637,N_619,N_775);
or U1638 (N_1638,N_559,N_494);
or U1639 (N_1639,N_23,N_154);
nor U1640 (N_1640,N_8,N_643);
nor U1641 (N_1641,N_860,N_794);
or U1642 (N_1642,N_350,N_295);
nor U1643 (N_1643,N_441,N_152);
nor U1644 (N_1644,N_832,N_979);
nand U1645 (N_1645,N_235,N_316);
nor U1646 (N_1646,N_462,N_81);
or U1647 (N_1647,N_121,N_102);
and U1648 (N_1648,N_577,N_224);
or U1649 (N_1649,N_180,N_46);
nor U1650 (N_1650,N_324,N_380);
or U1651 (N_1651,N_128,N_251);
and U1652 (N_1652,N_427,N_633);
and U1653 (N_1653,N_312,N_199);
and U1654 (N_1654,N_642,N_79);
and U1655 (N_1655,N_126,N_864);
nand U1656 (N_1656,N_392,N_283);
nand U1657 (N_1657,N_699,N_766);
nor U1658 (N_1658,N_783,N_482);
or U1659 (N_1659,N_445,N_151);
and U1660 (N_1660,N_23,N_814);
nor U1661 (N_1661,N_957,N_703);
or U1662 (N_1662,N_565,N_200);
or U1663 (N_1663,N_749,N_407);
or U1664 (N_1664,N_713,N_479);
xor U1665 (N_1665,N_954,N_793);
or U1666 (N_1666,N_776,N_423);
nand U1667 (N_1667,N_169,N_104);
nand U1668 (N_1668,N_677,N_200);
nor U1669 (N_1669,N_109,N_940);
nand U1670 (N_1670,N_610,N_776);
nor U1671 (N_1671,N_149,N_210);
nand U1672 (N_1672,N_606,N_696);
and U1673 (N_1673,N_434,N_993);
nand U1674 (N_1674,N_811,N_873);
nand U1675 (N_1675,N_928,N_967);
nor U1676 (N_1676,N_709,N_405);
or U1677 (N_1677,N_105,N_557);
or U1678 (N_1678,N_541,N_14);
nor U1679 (N_1679,N_540,N_660);
nand U1680 (N_1680,N_842,N_404);
nand U1681 (N_1681,N_356,N_31);
and U1682 (N_1682,N_33,N_295);
or U1683 (N_1683,N_649,N_226);
and U1684 (N_1684,N_832,N_639);
nand U1685 (N_1685,N_287,N_994);
nor U1686 (N_1686,N_802,N_997);
nand U1687 (N_1687,N_328,N_503);
nand U1688 (N_1688,N_552,N_113);
nor U1689 (N_1689,N_976,N_968);
nand U1690 (N_1690,N_444,N_839);
or U1691 (N_1691,N_422,N_59);
nand U1692 (N_1692,N_38,N_27);
nor U1693 (N_1693,N_998,N_240);
and U1694 (N_1694,N_483,N_293);
or U1695 (N_1695,N_459,N_69);
or U1696 (N_1696,N_104,N_493);
nand U1697 (N_1697,N_496,N_375);
nand U1698 (N_1698,N_420,N_294);
nand U1699 (N_1699,N_70,N_562);
nand U1700 (N_1700,N_686,N_393);
or U1701 (N_1701,N_426,N_206);
and U1702 (N_1702,N_268,N_594);
nand U1703 (N_1703,N_445,N_932);
nand U1704 (N_1704,N_289,N_478);
nor U1705 (N_1705,N_737,N_987);
nor U1706 (N_1706,N_287,N_688);
nand U1707 (N_1707,N_805,N_490);
nand U1708 (N_1708,N_628,N_629);
or U1709 (N_1709,N_668,N_521);
nand U1710 (N_1710,N_61,N_243);
or U1711 (N_1711,N_682,N_392);
and U1712 (N_1712,N_784,N_696);
and U1713 (N_1713,N_556,N_906);
nand U1714 (N_1714,N_600,N_705);
or U1715 (N_1715,N_117,N_602);
and U1716 (N_1716,N_975,N_146);
nand U1717 (N_1717,N_510,N_18);
nor U1718 (N_1718,N_588,N_298);
nor U1719 (N_1719,N_31,N_908);
nor U1720 (N_1720,N_265,N_290);
and U1721 (N_1721,N_772,N_459);
or U1722 (N_1722,N_223,N_460);
nand U1723 (N_1723,N_627,N_781);
and U1724 (N_1724,N_558,N_728);
and U1725 (N_1725,N_273,N_228);
nor U1726 (N_1726,N_529,N_790);
and U1727 (N_1727,N_103,N_941);
or U1728 (N_1728,N_337,N_225);
nand U1729 (N_1729,N_2,N_996);
or U1730 (N_1730,N_937,N_567);
and U1731 (N_1731,N_931,N_311);
nor U1732 (N_1732,N_915,N_497);
nor U1733 (N_1733,N_15,N_721);
or U1734 (N_1734,N_446,N_397);
nand U1735 (N_1735,N_326,N_618);
and U1736 (N_1736,N_45,N_582);
nand U1737 (N_1737,N_579,N_629);
or U1738 (N_1738,N_412,N_410);
and U1739 (N_1739,N_329,N_668);
or U1740 (N_1740,N_511,N_257);
nor U1741 (N_1741,N_974,N_30);
nand U1742 (N_1742,N_989,N_144);
nor U1743 (N_1743,N_281,N_82);
nor U1744 (N_1744,N_898,N_401);
nor U1745 (N_1745,N_258,N_399);
nand U1746 (N_1746,N_921,N_154);
or U1747 (N_1747,N_11,N_571);
nand U1748 (N_1748,N_16,N_718);
nand U1749 (N_1749,N_988,N_321);
or U1750 (N_1750,N_259,N_535);
nand U1751 (N_1751,N_549,N_869);
or U1752 (N_1752,N_610,N_654);
nand U1753 (N_1753,N_62,N_24);
or U1754 (N_1754,N_482,N_765);
nor U1755 (N_1755,N_262,N_457);
and U1756 (N_1756,N_353,N_916);
or U1757 (N_1757,N_516,N_957);
nand U1758 (N_1758,N_33,N_718);
nand U1759 (N_1759,N_37,N_660);
or U1760 (N_1760,N_748,N_333);
or U1761 (N_1761,N_420,N_719);
nand U1762 (N_1762,N_718,N_947);
nor U1763 (N_1763,N_349,N_952);
or U1764 (N_1764,N_775,N_893);
and U1765 (N_1765,N_865,N_145);
and U1766 (N_1766,N_120,N_947);
nand U1767 (N_1767,N_586,N_648);
and U1768 (N_1768,N_437,N_860);
nor U1769 (N_1769,N_211,N_885);
nand U1770 (N_1770,N_980,N_850);
or U1771 (N_1771,N_746,N_766);
and U1772 (N_1772,N_220,N_347);
nor U1773 (N_1773,N_539,N_40);
and U1774 (N_1774,N_771,N_252);
nor U1775 (N_1775,N_994,N_521);
xor U1776 (N_1776,N_872,N_533);
or U1777 (N_1777,N_917,N_935);
and U1778 (N_1778,N_578,N_633);
and U1779 (N_1779,N_593,N_477);
nor U1780 (N_1780,N_563,N_252);
or U1781 (N_1781,N_873,N_67);
nand U1782 (N_1782,N_636,N_217);
and U1783 (N_1783,N_685,N_365);
nor U1784 (N_1784,N_387,N_14);
nor U1785 (N_1785,N_201,N_726);
and U1786 (N_1786,N_622,N_582);
nor U1787 (N_1787,N_697,N_788);
nor U1788 (N_1788,N_530,N_346);
nand U1789 (N_1789,N_356,N_665);
or U1790 (N_1790,N_875,N_77);
nor U1791 (N_1791,N_907,N_397);
nand U1792 (N_1792,N_456,N_409);
nand U1793 (N_1793,N_295,N_601);
nand U1794 (N_1794,N_538,N_695);
nor U1795 (N_1795,N_223,N_479);
and U1796 (N_1796,N_748,N_833);
nor U1797 (N_1797,N_867,N_281);
nor U1798 (N_1798,N_503,N_974);
xnor U1799 (N_1799,N_3,N_990);
or U1800 (N_1800,N_873,N_292);
nor U1801 (N_1801,N_916,N_232);
or U1802 (N_1802,N_699,N_394);
or U1803 (N_1803,N_128,N_248);
and U1804 (N_1804,N_961,N_21);
nor U1805 (N_1805,N_232,N_934);
nor U1806 (N_1806,N_29,N_151);
xor U1807 (N_1807,N_428,N_221);
or U1808 (N_1808,N_354,N_579);
or U1809 (N_1809,N_834,N_100);
xor U1810 (N_1810,N_549,N_614);
nor U1811 (N_1811,N_329,N_821);
and U1812 (N_1812,N_539,N_960);
and U1813 (N_1813,N_327,N_938);
nand U1814 (N_1814,N_493,N_70);
and U1815 (N_1815,N_640,N_105);
nand U1816 (N_1816,N_342,N_614);
or U1817 (N_1817,N_635,N_555);
or U1818 (N_1818,N_589,N_500);
or U1819 (N_1819,N_671,N_668);
nand U1820 (N_1820,N_960,N_193);
and U1821 (N_1821,N_427,N_903);
or U1822 (N_1822,N_126,N_215);
or U1823 (N_1823,N_534,N_332);
nand U1824 (N_1824,N_903,N_62);
and U1825 (N_1825,N_693,N_863);
nand U1826 (N_1826,N_939,N_898);
or U1827 (N_1827,N_764,N_592);
or U1828 (N_1828,N_587,N_856);
nor U1829 (N_1829,N_200,N_525);
nand U1830 (N_1830,N_788,N_926);
xor U1831 (N_1831,N_875,N_807);
and U1832 (N_1832,N_100,N_380);
nor U1833 (N_1833,N_295,N_35);
nand U1834 (N_1834,N_698,N_375);
or U1835 (N_1835,N_403,N_40);
and U1836 (N_1836,N_64,N_812);
nor U1837 (N_1837,N_941,N_247);
nand U1838 (N_1838,N_346,N_524);
nand U1839 (N_1839,N_498,N_740);
or U1840 (N_1840,N_728,N_229);
and U1841 (N_1841,N_737,N_776);
and U1842 (N_1842,N_639,N_84);
nor U1843 (N_1843,N_731,N_591);
or U1844 (N_1844,N_589,N_212);
and U1845 (N_1845,N_893,N_60);
or U1846 (N_1846,N_726,N_735);
nand U1847 (N_1847,N_799,N_750);
and U1848 (N_1848,N_42,N_616);
nor U1849 (N_1849,N_358,N_685);
or U1850 (N_1850,N_435,N_382);
or U1851 (N_1851,N_748,N_375);
nand U1852 (N_1852,N_884,N_678);
or U1853 (N_1853,N_532,N_856);
nand U1854 (N_1854,N_165,N_915);
nor U1855 (N_1855,N_190,N_558);
nor U1856 (N_1856,N_330,N_274);
nand U1857 (N_1857,N_324,N_59);
nor U1858 (N_1858,N_135,N_945);
and U1859 (N_1859,N_51,N_300);
nor U1860 (N_1860,N_646,N_485);
xor U1861 (N_1861,N_762,N_425);
or U1862 (N_1862,N_722,N_879);
or U1863 (N_1863,N_426,N_761);
nor U1864 (N_1864,N_574,N_116);
and U1865 (N_1865,N_130,N_943);
nor U1866 (N_1866,N_532,N_506);
xnor U1867 (N_1867,N_606,N_727);
or U1868 (N_1868,N_979,N_857);
or U1869 (N_1869,N_387,N_731);
and U1870 (N_1870,N_57,N_107);
or U1871 (N_1871,N_919,N_13);
nor U1872 (N_1872,N_218,N_349);
or U1873 (N_1873,N_9,N_891);
nor U1874 (N_1874,N_3,N_238);
nand U1875 (N_1875,N_7,N_411);
and U1876 (N_1876,N_678,N_261);
nor U1877 (N_1877,N_331,N_401);
and U1878 (N_1878,N_687,N_602);
or U1879 (N_1879,N_754,N_361);
or U1880 (N_1880,N_554,N_847);
and U1881 (N_1881,N_85,N_503);
or U1882 (N_1882,N_677,N_760);
or U1883 (N_1883,N_627,N_815);
nand U1884 (N_1884,N_527,N_971);
and U1885 (N_1885,N_754,N_416);
nor U1886 (N_1886,N_544,N_959);
nor U1887 (N_1887,N_883,N_415);
nand U1888 (N_1888,N_674,N_735);
xor U1889 (N_1889,N_715,N_501);
and U1890 (N_1890,N_863,N_898);
or U1891 (N_1891,N_89,N_874);
nand U1892 (N_1892,N_818,N_649);
and U1893 (N_1893,N_925,N_803);
or U1894 (N_1894,N_33,N_522);
nand U1895 (N_1895,N_490,N_286);
and U1896 (N_1896,N_327,N_280);
nand U1897 (N_1897,N_394,N_860);
or U1898 (N_1898,N_408,N_784);
nand U1899 (N_1899,N_908,N_210);
nor U1900 (N_1900,N_600,N_109);
nand U1901 (N_1901,N_971,N_207);
or U1902 (N_1902,N_596,N_707);
nand U1903 (N_1903,N_618,N_405);
nor U1904 (N_1904,N_958,N_966);
and U1905 (N_1905,N_665,N_927);
or U1906 (N_1906,N_37,N_147);
nand U1907 (N_1907,N_762,N_162);
or U1908 (N_1908,N_343,N_646);
and U1909 (N_1909,N_671,N_368);
or U1910 (N_1910,N_628,N_127);
and U1911 (N_1911,N_811,N_844);
or U1912 (N_1912,N_816,N_676);
nor U1913 (N_1913,N_836,N_898);
nor U1914 (N_1914,N_273,N_551);
and U1915 (N_1915,N_458,N_598);
nand U1916 (N_1916,N_957,N_124);
nor U1917 (N_1917,N_49,N_673);
nand U1918 (N_1918,N_137,N_779);
and U1919 (N_1919,N_998,N_132);
nand U1920 (N_1920,N_949,N_512);
nor U1921 (N_1921,N_714,N_608);
and U1922 (N_1922,N_995,N_860);
nand U1923 (N_1923,N_736,N_425);
and U1924 (N_1924,N_835,N_734);
nor U1925 (N_1925,N_426,N_32);
nor U1926 (N_1926,N_405,N_154);
or U1927 (N_1927,N_173,N_743);
or U1928 (N_1928,N_642,N_826);
or U1929 (N_1929,N_401,N_534);
and U1930 (N_1930,N_444,N_815);
and U1931 (N_1931,N_149,N_69);
nand U1932 (N_1932,N_290,N_82);
nor U1933 (N_1933,N_414,N_495);
nor U1934 (N_1934,N_428,N_245);
nor U1935 (N_1935,N_329,N_527);
or U1936 (N_1936,N_197,N_114);
or U1937 (N_1937,N_923,N_241);
nand U1938 (N_1938,N_27,N_152);
nor U1939 (N_1939,N_687,N_990);
nand U1940 (N_1940,N_693,N_666);
or U1941 (N_1941,N_580,N_432);
or U1942 (N_1942,N_120,N_187);
nand U1943 (N_1943,N_57,N_367);
nand U1944 (N_1944,N_308,N_596);
or U1945 (N_1945,N_100,N_27);
nor U1946 (N_1946,N_899,N_235);
nor U1947 (N_1947,N_121,N_514);
or U1948 (N_1948,N_23,N_679);
nor U1949 (N_1949,N_481,N_415);
nand U1950 (N_1950,N_695,N_340);
nor U1951 (N_1951,N_921,N_474);
and U1952 (N_1952,N_82,N_609);
nand U1953 (N_1953,N_690,N_790);
nor U1954 (N_1954,N_541,N_312);
nand U1955 (N_1955,N_98,N_148);
nand U1956 (N_1956,N_467,N_891);
nor U1957 (N_1957,N_389,N_396);
nand U1958 (N_1958,N_13,N_664);
and U1959 (N_1959,N_37,N_875);
or U1960 (N_1960,N_941,N_240);
or U1961 (N_1961,N_965,N_213);
nand U1962 (N_1962,N_535,N_574);
or U1963 (N_1963,N_846,N_851);
nor U1964 (N_1964,N_844,N_622);
or U1965 (N_1965,N_91,N_102);
or U1966 (N_1966,N_655,N_674);
nand U1967 (N_1967,N_251,N_345);
nor U1968 (N_1968,N_516,N_262);
nor U1969 (N_1969,N_585,N_313);
and U1970 (N_1970,N_470,N_116);
xor U1971 (N_1971,N_898,N_662);
and U1972 (N_1972,N_877,N_750);
nand U1973 (N_1973,N_285,N_985);
nor U1974 (N_1974,N_917,N_85);
and U1975 (N_1975,N_305,N_875);
nor U1976 (N_1976,N_103,N_693);
or U1977 (N_1977,N_947,N_181);
or U1978 (N_1978,N_225,N_930);
nand U1979 (N_1979,N_780,N_264);
nor U1980 (N_1980,N_657,N_136);
nand U1981 (N_1981,N_381,N_318);
nor U1982 (N_1982,N_354,N_273);
and U1983 (N_1983,N_869,N_937);
or U1984 (N_1984,N_642,N_695);
and U1985 (N_1985,N_406,N_437);
nand U1986 (N_1986,N_379,N_433);
or U1987 (N_1987,N_488,N_772);
or U1988 (N_1988,N_582,N_248);
and U1989 (N_1989,N_8,N_802);
nand U1990 (N_1990,N_602,N_212);
nor U1991 (N_1991,N_6,N_660);
nand U1992 (N_1992,N_618,N_855);
nor U1993 (N_1993,N_961,N_541);
or U1994 (N_1994,N_403,N_945);
nor U1995 (N_1995,N_508,N_760);
or U1996 (N_1996,N_981,N_927);
nand U1997 (N_1997,N_125,N_754);
nand U1998 (N_1998,N_726,N_712);
or U1999 (N_1999,N_610,N_566);
nor U2000 (N_2000,N_1837,N_1954);
and U2001 (N_2001,N_1951,N_1306);
or U2002 (N_2002,N_1680,N_1710);
nand U2003 (N_2003,N_1629,N_1350);
nor U2004 (N_2004,N_1151,N_1188);
and U2005 (N_2005,N_1155,N_1196);
and U2006 (N_2006,N_1846,N_1296);
or U2007 (N_2007,N_1735,N_1496);
nand U2008 (N_2008,N_1687,N_1560);
nand U2009 (N_2009,N_1011,N_1286);
nor U2010 (N_2010,N_1477,N_1912);
nor U2011 (N_2011,N_1720,N_1375);
nand U2012 (N_2012,N_1161,N_1473);
nand U2013 (N_2013,N_1441,N_1044);
and U2014 (N_2014,N_1120,N_1398);
nor U2015 (N_2015,N_1232,N_1952);
nor U2016 (N_2016,N_1834,N_1715);
nand U2017 (N_2017,N_1076,N_1499);
or U2018 (N_2018,N_1130,N_1182);
nor U2019 (N_2019,N_1276,N_1908);
or U2020 (N_2020,N_1364,N_1734);
nor U2021 (N_2021,N_1992,N_1063);
or U2022 (N_2022,N_1737,N_1452);
or U2023 (N_2023,N_1503,N_1465);
nand U2024 (N_2024,N_1858,N_1935);
nor U2025 (N_2025,N_1037,N_1875);
nor U2026 (N_2026,N_1368,N_1742);
and U2027 (N_2027,N_1913,N_1923);
nand U2028 (N_2028,N_1110,N_1684);
and U2029 (N_2029,N_1870,N_1975);
or U2030 (N_2030,N_1934,N_1245);
nand U2031 (N_2031,N_1509,N_1861);
or U2032 (N_2032,N_1024,N_1365);
nor U2033 (N_2033,N_1847,N_1816);
nand U2034 (N_2034,N_1936,N_1616);
xnor U2035 (N_2035,N_1813,N_1493);
and U2036 (N_2036,N_1279,N_1795);
nor U2037 (N_2037,N_1086,N_1422);
or U2038 (N_2038,N_1012,N_1964);
nor U2039 (N_2039,N_1378,N_1740);
and U2040 (N_2040,N_1454,N_1756);
nor U2041 (N_2041,N_1432,N_1318);
or U2042 (N_2042,N_1057,N_1209);
nor U2043 (N_2043,N_1307,N_1402);
or U2044 (N_2044,N_1755,N_1450);
or U2045 (N_2045,N_1361,N_1546);
and U2046 (N_2046,N_1930,N_1412);
and U2047 (N_2047,N_1494,N_1914);
nor U2048 (N_2048,N_1036,N_1367);
xor U2049 (N_2049,N_1303,N_1071);
nand U2050 (N_2050,N_1202,N_1143);
and U2051 (N_2051,N_1711,N_1467);
nor U2052 (N_2052,N_1114,N_1418);
nand U2053 (N_2053,N_1449,N_1396);
nand U2054 (N_2054,N_1772,N_1758);
nand U2055 (N_2055,N_1652,N_1280);
nand U2056 (N_2056,N_1391,N_1619);
and U2057 (N_2057,N_1163,N_1270);
and U2058 (N_2058,N_1134,N_1938);
nand U2059 (N_2059,N_1683,N_1943);
and U2060 (N_2060,N_1371,N_1738);
nor U2061 (N_2061,N_1713,N_1087);
nand U2062 (N_2062,N_1671,N_1215);
and U2063 (N_2063,N_1984,N_1828);
nand U2064 (N_2064,N_1133,N_1246);
and U2065 (N_2065,N_1067,N_1996);
and U2066 (N_2066,N_1778,N_1191);
nand U2067 (N_2067,N_1424,N_1453);
and U2068 (N_2068,N_1567,N_1839);
and U2069 (N_2069,N_1591,N_1323);
or U2070 (N_2070,N_1681,N_1405);
or U2071 (N_2071,N_1404,N_1670);
nor U2072 (N_2072,N_1920,N_1489);
nand U2073 (N_2073,N_1005,N_1138);
and U2074 (N_2074,N_1370,N_1458);
nand U2075 (N_2075,N_1158,N_1252);
or U2076 (N_2076,N_1115,N_1564);
nor U2077 (N_2077,N_1794,N_1127);
or U2078 (N_2078,N_1249,N_1132);
nor U2079 (N_2079,N_1113,N_1519);
and U2080 (N_2080,N_1430,N_1879);
or U2081 (N_2081,N_1167,N_1919);
and U2082 (N_2082,N_1853,N_1857);
or U2083 (N_2083,N_1198,N_1128);
nand U2084 (N_2084,N_1907,N_1312);
nor U2085 (N_2085,N_1906,N_1599);
nor U2086 (N_2086,N_1070,N_1866);
and U2087 (N_2087,N_1725,N_1208);
and U2088 (N_2088,N_1739,N_1317);
nand U2089 (N_2089,N_1692,N_1490);
nand U2090 (N_2090,N_1171,N_1457);
and U2091 (N_2091,N_1829,N_1135);
nor U2092 (N_2092,N_1123,N_1415);
or U2093 (N_2093,N_1041,N_1596);
nor U2094 (N_2094,N_1470,N_1302);
or U2095 (N_2095,N_1403,N_1408);
and U2096 (N_2096,N_1407,N_1886);
nand U2097 (N_2097,N_1379,N_1767);
and U2098 (N_2098,N_1807,N_1820);
nor U2099 (N_2099,N_1573,N_1961);
nor U2100 (N_2100,N_1637,N_1304);
or U2101 (N_2101,N_1508,N_1235);
or U2102 (N_2102,N_1401,N_1189);
nor U2103 (N_2103,N_1497,N_1145);
and U2104 (N_2104,N_1831,N_1360);
nor U2105 (N_2105,N_1417,N_1889);
or U2106 (N_2106,N_1008,N_1109);
nand U2107 (N_2107,N_1491,N_1200);
nor U2108 (N_2108,N_1221,N_1848);
and U2109 (N_2109,N_1763,N_1691);
or U2110 (N_2110,N_1605,N_1771);
nor U2111 (N_2111,N_1634,N_1849);
and U2112 (N_2112,N_1630,N_1594);
nand U2113 (N_2113,N_1881,N_1411);
nand U2114 (N_2114,N_1768,N_1156);
nand U2115 (N_2115,N_1278,N_1621);
and U2116 (N_2116,N_1520,N_1542);
and U2117 (N_2117,N_1856,N_1827);
nand U2118 (N_2118,N_1724,N_1141);
or U2119 (N_2119,N_1815,N_1655);
nor U2120 (N_2120,N_1474,N_1607);
nand U2121 (N_2121,N_1501,N_1841);
nor U2122 (N_2122,N_1150,N_1911);
nor U2123 (N_2123,N_1420,N_1259);
nand U2124 (N_2124,N_1268,N_1233);
and U2125 (N_2125,N_1618,N_1550);
or U2126 (N_2126,N_1210,N_1356);
nor U2127 (N_2127,N_1372,N_1170);
nor U2128 (N_2128,N_1104,N_1628);
nand U2129 (N_2129,N_1103,N_1184);
or U2130 (N_2130,N_1265,N_1043);
nor U2131 (N_2131,N_1970,N_1862);
or U2132 (N_2132,N_1531,N_1642);
or U2133 (N_2133,N_1603,N_1898);
and U2134 (N_2134,N_1785,N_1892);
nand U2135 (N_2135,N_1944,N_1777);
and U2136 (N_2136,N_1100,N_1878);
nand U2137 (N_2137,N_1525,N_1425);
and U2138 (N_2138,N_1002,N_1064);
nand U2139 (N_2139,N_1125,N_1993);
nor U2140 (N_2140,N_1787,N_1098);
and U2141 (N_2141,N_1714,N_1243);
nand U2142 (N_2142,N_1555,N_1721);
and U2143 (N_2143,N_1903,N_1038);
nor U2144 (N_2144,N_1685,N_1874);
and U2145 (N_2145,N_1593,N_1034);
nor U2146 (N_2146,N_1320,N_1447);
or U2147 (N_2147,N_1112,N_1102);
nand U2148 (N_2148,N_1662,N_1639);
xnor U2149 (N_2149,N_1595,N_1551);
or U2150 (N_2150,N_1389,N_1598);
and U2151 (N_2151,N_1495,N_1948);
nor U2152 (N_2152,N_1949,N_1747);
and U2153 (N_2153,N_1661,N_1040);
nand U2154 (N_2154,N_1337,N_1225);
nand U2155 (N_2155,N_1623,N_1230);
nor U2156 (N_2156,N_1958,N_1077);
nor U2157 (N_2157,N_1451,N_1313);
nor U2158 (N_2158,N_1987,N_1884);
nand U2159 (N_2159,N_1479,N_1448);
and U2160 (N_2160,N_1089,N_1678);
nor U2161 (N_2161,N_1674,N_1187);
nor U2162 (N_2162,N_1440,N_1237);
and U2163 (N_2163,N_1843,N_1563);
xnor U2164 (N_2164,N_1533,N_1649);
nor U2165 (N_2165,N_1290,N_1093);
nor U2166 (N_2166,N_1427,N_1705);
and U2167 (N_2167,N_1030,N_1169);
or U2168 (N_2168,N_1835,N_1255);
and U2169 (N_2169,N_1083,N_1275);
and U2170 (N_2170,N_1443,N_1055);
and U2171 (N_2171,N_1224,N_1324);
and U2172 (N_2172,N_1909,N_1969);
nor U2173 (N_2173,N_1695,N_1781);
nor U2174 (N_2174,N_1028,N_1314);
or U2175 (N_2175,N_1539,N_1585);
and U2176 (N_2176,N_1985,N_1199);
and U2177 (N_2177,N_1386,N_1216);
or U2178 (N_2178,N_1332,N_1883);
nand U2179 (N_2179,N_1601,N_1515);
or U2180 (N_2180,N_1696,N_1126);
nor U2181 (N_2181,N_1700,N_1543);
or U2182 (N_2182,N_1462,N_1287);
or U2183 (N_2183,N_1741,N_1111);
or U2184 (N_2184,N_1565,N_1090);
nor U2185 (N_2185,N_1343,N_1728);
and U2186 (N_2186,N_1798,N_1446);
nor U2187 (N_2187,N_1894,N_1885);
nand U2188 (N_2188,N_1393,N_1376);
or U2189 (N_2189,N_1284,N_1006);
or U2190 (N_2190,N_1385,N_1638);
nor U2191 (N_2191,N_1541,N_1010);
and U2192 (N_2192,N_1048,N_1776);
and U2193 (N_2193,N_1792,N_1810);
and U2194 (N_2194,N_1963,N_1693);
nor U2195 (N_2195,N_1609,N_1748);
nand U2196 (N_2196,N_1223,N_1622);
nand U2197 (N_2197,N_1485,N_1344);
nand U2198 (N_2198,N_1434,N_1097);
nor U2199 (N_2199,N_1178,N_1397);
nand U2200 (N_2200,N_1806,N_1081);
and U2201 (N_2201,N_1261,N_1234);
or U2202 (N_2202,N_1633,N_1207);
nand U2203 (N_2203,N_1289,N_1394);
nor U2204 (N_2204,N_1164,N_1995);
and U2205 (N_2205,N_1066,N_1990);
or U2206 (N_2206,N_1799,N_1088);
nand U2207 (N_2207,N_1615,N_1339);
and U2208 (N_2208,N_1780,N_1545);
nor U2209 (N_2209,N_1392,N_1084);
and U2210 (N_2210,N_1775,N_1877);
and U2211 (N_2211,N_1309,N_1597);
nand U2212 (N_2212,N_1193,N_1413);
and U2213 (N_2213,N_1698,N_1410);
and U2214 (N_2214,N_1973,N_1762);
nor U2215 (N_2215,N_1764,N_1487);
and U2216 (N_2216,N_1706,N_1718);
nand U2217 (N_2217,N_1014,N_1626);
or U2218 (N_2218,N_1352,N_1957);
and U2219 (N_2219,N_1635,N_1229);
nor U2220 (N_2220,N_1569,N_1068);
or U2221 (N_2221,N_1647,N_1850);
and U2222 (N_2222,N_1211,N_1459);
nand U2223 (N_2223,N_1643,N_1183);
or U2224 (N_2224,N_1940,N_1978);
and U2225 (N_2225,N_1802,N_1033);
nor U2226 (N_2226,N_1845,N_1997);
or U2227 (N_2227,N_1197,N_1466);
nor U2228 (N_2228,N_1521,N_1712);
and U2229 (N_2229,N_1013,N_1264);
and U2230 (N_2230,N_1315,N_1653);
and U2231 (N_2231,N_1836,N_1868);
nand U2232 (N_2232,N_1026,N_1108);
nand U2233 (N_2233,N_1650,N_1099);
and U2234 (N_2234,N_1004,N_1366);
nor U2235 (N_2235,N_1166,N_1950);
or U2236 (N_2236,N_1553,N_1932);
nor U2237 (N_2237,N_1482,N_1744);
nand U2238 (N_2238,N_1359,N_1173);
or U2239 (N_2239,N_1253,N_1241);
or U2240 (N_2240,N_1568,N_1078);
nand U2241 (N_2241,N_1056,N_1388);
nand U2242 (N_2242,N_1399,N_1617);
nand U2243 (N_2243,N_1025,N_1865);
or U2244 (N_2244,N_1334,N_1308);
nor U2245 (N_2245,N_1258,N_1727);
nor U2246 (N_2246,N_1291,N_1240);
nand U2247 (N_2247,N_1325,N_1073);
nand U2248 (N_2248,N_1460,N_1636);
and U2249 (N_2249,N_1904,N_1900);
nand U2250 (N_2250,N_1946,N_1227);
nand U2251 (N_2251,N_1974,N_1512);
nor U2252 (N_2252,N_1577,N_1529);
nor U2253 (N_2253,N_1212,N_1864);
or U2254 (N_2254,N_1994,N_1419);
nand U2255 (N_2255,N_1817,N_1916);
nand U2256 (N_2256,N_1119,N_1185);
or U2257 (N_2257,N_1065,N_1942);
and U2258 (N_2258,N_1625,N_1562);
nand U2259 (N_2259,N_1069,N_1266);
or U2260 (N_2260,N_1977,N_1690);
or U2261 (N_2261,N_1719,N_1540);
nand U2262 (N_2262,N_1971,N_1753);
or U2263 (N_2263,N_1558,N_1890);
or U2264 (N_2264,N_1377,N_1921);
or U2265 (N_2265,N_1736,N_1382);
or U2266 (N_2266,N_1707,N_1096);
nor U2267 (N_2267,N_1709,N_1080);
or U2268 (N_2268,N_1431,N_1075);
and U2269 (N_2269,N_1400,N_1165);
and U2270 (N_2270,N_1181,N_1094);
or U2271 (N_2271,N_1888,N_1613);
and U2272 (N_2272,N_1019,N_1640);
nand U2273 (N_2273,N_1283,N_1941);
xor U2274 (N_2274,N_1537,N_1154);
nand U2275 (N_2275,N_1136,N_1045);
nand U2276 (N_2276,N_1582,N_1106);
and U2277 (N_2277,N_1085,N_1373);
nand U2278 (N_2278,N_1395,N_1580);
and U2279 (N_2279,N_1242,N_1267);
or U2280 (N_2280,N_1105,N_1572);
nor U2281 (N_2281,N_1982,N_1179);
and U2282 (N_2282,N_1416,N_1142);
or U2283 (N_2283,N_1924,N_1821);
nand U2284 (N_2284,N_1620,N_1789);
and U2285 (N_2285,N_1757,N_1042);
and U2286 (N_2286,N_1631,N_1228);
and U2287 (N_2287,N_1770,N_1140);
nor U2288 (N_2288,N_1860,N_1483);
nor U2289 (N_2289,N_1654,N_1321);
nor U2290 (N_2290,N_1575,N_1688);
xnor U2291 (N_2291,N_1809,N_1147);
nand U2292 (N_2292,N_1513,N_1480);
or U2293 (N_2293,N_1192,N_1122);
or U2294 (N_2294,N_1651,N_1007);
or U2295 (N_2295,N_1020,N_1387);
nor U2296 (N_2296,N_1988,N_1703);
nand U2297 (N_2297,N_1863,N_1749);
or U2298 (N_2298,N_1701,N_1759);
nor U2299 (N_2299,N_1058,N_1316);
and U2300 (N_2300,N_1967,N_1524);
and U2301 (N_2301,N_1262,N_1476);
or U2302 (N_2302,N_1062,N_1588);
nor U2303 (N_2303,N_1047,N_1552);
nand U2304 (N_2304,N_1955,N_1137);
or U2305 (N_2305,N_1348,N_1330);
nand U2306 (N_2306,N_1897,N_1676);
or U2307 (N_2307,N_1390,N_1409);
or U2308 (N_2308,N_1061,N_1003);
and U2309 (N_2309,N_1902,N_1804);
or U2310 (N_2310,N_1426,N_1729);
nor U2311 (N_2311,N_1101,N_1292);
and U2312 (N_2312,N_1472,N_1733);
and U2313 (N_2313,N_1731,N_1374);
nand U2314 (N_2314,N_1338,N_1231);
or U2315 (N_2315,N_1664,N_1910);
and U2316 (N_2316,N_1561,N_1566);
nand U2317 (N_2317,N_1803,N_1819);
nor U2318 (N_2318,N_1592,N_1218);
nand U2319 (N_2319,N_1668,N_1646);
or U2320 (N_2320,N_1146,N_1851);
and U2321 (N_2321,N_1293,N_1027);
and U2322 (N_2322,N_1423,N_1722);
nand U2323 (N_2323,N_1752,N_1611);
or U2324 (N_2324,N_1554,N_1095);
or U2325 (N_2325,N_1523,N_1009);
nand U2326 (N_2326,N_1021,N_1018);
and U2327 (N_2327,N_1586,N_1257);
or U2328 (N_2328,N_1281,N_1659);
and U2329 (N_2329,N_1665,N_1072);
nand U2330 (N_2330,N_1331,N_1251);
nor U2331 (N_2331,N_1129,N_1250);
or U2332 (N_2332,N_1966,N_1438);
or U2333 (N_2333,N_1406,N_1478);
and U2334 (N_2334,N_1991,N_1750);
and U2335 (N_2335,N_1505,N_1269);
or U2336 (N_2336,N_1979,N_1172);
and U2337 (N_2337,N_1384,N_1148);
or U2338 (N_2338,N_1838,N_1301);
or U2339 (N_2339,N_1504,N_1825);
nand U2340 (N_2340,N_1644,N_1937);
nand U2341 (N_2341,N_1723,N_1669);
nor U2342 (N_2342,N_1786,N_1205);
and U2343 (N_2343,N_1213,N_1031);
or U2344 (N_2344,N_1627,N_1353);
and U2345 (N_2345,N_1514,N_1699);
or U2346 (N_2346,N_1238,N_1782);
or U2347 (N_2347,N_1354,N_1180);
or U2348 (N_2348,N_1867,N_1000);
nor U2349 (N_2349,N_1274,N_1805);
nor U2350 (N_2350,N_1830,N_1358);
or U2351 (N_2351,N_1282,N_1972);
and U2352 (N_2352,N_1689,N_1814);
or U2353 (N_2353,N_1190,N_1355);
nor U2354 (N_2354,N_1498,N_1606);
nand U2355 (N_2355,N_1023,N_1502);
nand U2356 (N_2356,N_1175,N_1186);
or U2357 (N_2357,N_1139,N_1437);
nand U2358 (N_2358,N_1931,N_1507);
and U2359 (N_2359,N_1801,N_1896);
and U2360 (N_2360,N_1357,N_1428);
or U2361 (N_2361,N_1796,N_1176);
and U2362 (N_2362,N_1162,N_1658);
nor U2363 (N_2363,N_1899,N_1107);
or U2364 (N_2364,N_1677,N_1947);
nand U2365 (N_2365,N_1694,N_1288);
nor U2366 (N_2366,N_1516,N_1578);
nand U2367 (N_2367,N_1918,N_1882);
and U2368 (N_2368,N_1029,N_1528);
or U2369 (N_2369,N_1570,N_1471);
xor U2370 (N_2370,N_1672,N_1660);
nand U2371 (N_2371,N_1214,N_1091);
and U2372 (N_2372,N_1832,N_1854);
nand U2373 (N_2373,N_1116,N_1206);
nand U2374 (N_2374,N_1239,N_1797);
nor U2375 (N_2375,N_1632,N_1435);
nor U2376 (N_2376,N_1362,N_1340);
or U2377 (N_2377,N_1160,N_1124);
nand U2378 (N_2378,N_1518,N_1842);
or U2379 (N_2379,N_1455,N_1702);
nor U2380 (N_2380,N_1981,N_1587);
nand U2381 (N_2381,N_1421,N_1880);
or U2382 (N_2382,N_1152,N_1998);
or U2383 (N_2383,N_1774,N_1891);
and U2384 (N_2384,N_1032,N_1769);
nor U2385 (N_2385,N_1745,N_1204);
and U2386 (N_2386,N_1244,N_1579);
and U2387 (N_2387,N_1201,N_1442);
and U2388 (N_2388,N_1547,N_1492);
or U2389 (N_2389,N_1926,N_1784);
or U2390 (N_2390,N_1534,N_1263);
nor U2391 (N_2391,N_1645,N_1793);
nor U2392 (N_2392,N_1035,N_1788);
nor U2393 (N_2393,N_1743,N_1463);
xnor U2394 (N_2394,N_1559,N_1818);
and U2395 (N_2395,N_1260,N_1117);
nor U2396 (N_2396,N_1351,N_1526);
xor U2397 (N_2397,N_1791,N_1604);
nor U2398 (N_2398,N_1581,N_1549);
nor U2399 (N_2399,N_1716,N_1369);
nand U2400 (N_2400,N_1544,N_1956);
nand U2401 (N_2401,N_1761,N_1965);
and U2402 (N_2402,N_1824,N_1663);
or U2403 (N_2403,N_1548,N_1329);
nor U2404 (N_2404,N_1667,N_1247);
nand U2405 (N_2405,N_1826,N_1294);
and U2406 (N_2406,N_1256,N_1049);
or U2407 (N_2407,N_1194,N_1174);
nor U2408 (N_2408,N_1469,N_1177);
or U2409 (N_2409,N_1871,N_1925);
or U2410 (N_2410,N_1149,N_1766);
nor U2411 (N_2411,N_1059,N_1872);
nor U2412 (N_2412,N_1050,N_1319);
and U2413 (N_2413,N_1046,N_1751);
or U2414 (N_2414,N_1574,N_1960);
nor U2415 (N_2415,N_1641,N_1989);
or U2416 (N_2416,N_1697,N_1530);
nand U2417 (N_2417,N_1612,N_1833);
nor U2418 (N_2418,N_1052,N_1610);
and U2419 (N_2419,N_1939,N_1682);
xnor U2420 (N_2420,N_1429,N_1708);
or U2421 (N_2421,N_1506,N_1273);
and U2422 (N_2422,N_1444,N_1962);
and U2423 (N_2423,N_1336,N_1905);
nand U2424 (N_2424,N_1051,N_1322);
nor U2425 (N_2425,N_1812,N_1657);
nor U2426 (N_2426,N_1779,N_1298);
or U2427 (N_2427,N_1153,N_1295);
nand U2428 (N_2428,N_1532,N_1060);
or U2429 (N_2429,N_1583,N_1760);
nor U2430 (N_2430,N_1203,N_1168);
nor U2431 (N_2431,N_1159,N_1349);
or U2432 (N_2432,N_1383,N_1277);
nand U2433 (N_2433,N_1873,N_1053);
nand U2434 (N_2434,N_1535,N_1517);
nand U2435 (N_2435,N_1922,N_1484);
nor U2436 (N_2436,N_1876,N_1686);
or U2437 (N_2437,N_1968,N_1345);
and U2438 (N_2438,N_1118,N_1039);
nor U2439 (N_2439,N_1976,N_1959);
nor U2440 (N_2440,N_1016,N_1488);
nand U2441 (N_2441,N_1022,N_1538);
nand U2442 (N_2442,N_1986,N_1980);
nor U2443 (N_2443,N_1486,N_1840);
nor U2444 (N_2444,N_1220,N_1576);
nand U2445 (N_2445,N_1363,N_1859);
nor U2446 (N_2446,N_1679,N_1335);
or U2447 (N_2447,N_1436,N_1226);
or U2448 (N_2448,N_1953,N_1844);
and U2449 (N_2449,N_1927,N_1675);
or U2450 (N_2450,N_1380,N_1217);
and U2451 (N_2451,N_1333,N_1614);
or U2452 (N_2452,N_1285,N_1726);
or U2453 (N_2453,N_1144,N_1999);
xor U2454 (N_2454,N_1536,N_1092);
nand U2455 (N_2455,N_1765,N_1461);
and U2456 (N_2456,N_1328,N_1717);
xor U2457 (N_2457,N_1254,N_1300);
and U2458 (N_2458,N_1666,N_1500);
or U2459 (N_2459,N_1624,N_1901);
nand U2460 (N_2460,N_1928,N_1945);
nand U2461 (N_2461,N_1915,N_1656);
or U2462 (N_2462,N_1602,N_1584);
nor U2463 (N_2463,N_1571,N_1790);
and U2464 (N_2464,N_1773,N_1445);
or U2465 (N_2465,N_1600,N_1248);
nand U2466 (N_2466,N_1887,N_1327);
and U2467 (N_2467,N_1299,N_1852);
and U2468 (N_2468,N_1310,N_1730);
nand U2469 (N_2469,N_1933,N_1855);
nor U2470 (N_2470,N_1608,N_1673);
nor U2471 (N_2471,N_1811,N_1917);
or U2472 (N_2472,N_1481,N_1510);
nor U2473 (N_2473,N_1131,N_1311);
and U2474 (N_2474,N_1305,N_1589);
nand U2475 (N_2475,N_1895,N_1381);
nor U2476 (N_2476,N_1556,N_1195);
or U2477 (N_2477,N_1522,N_1590);
nor U2478 (N_2478,N_1079,N_1464);
nand U2479 (N_2479,N_1704,N_1468);
or U2480 (N_2480,N_1475,N_1414);
and U2481 (N_2481,N_1869,N_1929);
nand U2482 (N_2482,N_1823,N_1732);
or U2483 (N_2483,N_1222,N_1219);
nand U2484 (N_2484,N_1326,N_1456);
nand U2485 (N_2485,N_1342,N_1433);
or U2486 (N_2486,N_1783,N_1236);
nor U2487 (N_2487,N_1297,N_1082);
nand U2488 (N_2488,N_1341,N_1054);
nand U2489 (N_2489,N_1800,N_1648);
nor U2490 (N_2490,N_1015,N_1983);
nand U2491 (N_2491,N_1746,N_1346);
nor U2492 (N_2492,N_1808,N_1439);
and U2493 (N_2493,N_1121,N_1347);
or U2494 (N_2494,N_1272,N_1557);
or U2495 (N_2495,N_1893,N_1271);
nor U2496 (N_2496,N_1017,N_1527);
nand U2497 (N_2497,N_1754,N_1157);
and U2498 (N_2498,N_1001,N_1511);
and U2499 (N_2499,N_1074,N_1822);
or U2500 (N_2500,N_1984,N_1506);
or U2501 (N_2501,N_1971,N_1287);
or U2502 (N_2502,N_1038,N_1229);
or U2503 (N_2503,N_1637,N_1680);
and U2504 (N_2504,N_1196,N_1388);
or U2505 (N_2505,N_1866,N_1158);
nand U2506 (N_2506,N_1437,N_1645);
or U2507 (N_2507,N_1996,N_1945);
nor U2508 (N_2508,N_1974,N_1389);
nor U2509 (N_2509,N_1149,N_1947);
nand U2510 (N_2510,N_1595,N_1587);
and U2511 (N_2511,N_1459,N_1756);
and U2512 (N_2512,N_1167,N_1624);
and U2513 (N_2513,N_1781,N_1043);
nor U2514 (N_2514,N_1731,N_1717);
nand U2515 (N_2515,N_1581,N_1331);
and U2516 (N_2516,N_1709,N_1812);
nand U2517 (N_2517,N_1593,N_1234);
nor U2518 (N_2518,N_1712,N_1848);
or U2519 (N_2519,N_1626,N_1782);
nor U2520 (N_2520,N_1106,N_1832);
or U2521 (N_2521,N_1134,N_1982);
nand U2522 (N_2522,N_1634,N_1546);
or U2523 (N_2523,N_1892,N_1277);
nand U2524 (N_2524,N_1984,N_1205);
nand U2525 (N_2525,N_1075,N_1544);
or U2526 (N_2526,N_1801,N_1601);
nor U2527 (N_2527,N_1438,N_1508);
and U2528 (N_2528,N_1616,N_1626);
nand U2529 (N_2529,N_1857,N_1395);
nand U2530 (N_2530,N_1797,N_1858);
and U2531 (N_2531,N_1079,N_1439);
nand U2532 (N_2532,N_1017,N_1993);
and U2533 (N_2533,N_1097,N_1096);
nand U2534 (N_2534,N_1949,N_1191);
nor U2535 (N_2535,N_1106,N_1618);
or U2536 (N_2536,N_1878,N_1359);
or U2537 (N_2537,N_1405,N_1960);
nand U2538 (N_2538,N_1680,N_1196);
nand U2539 (N_2539,N_1767,N_1226);
nor U2540 (N_2540,N_1225,N_1179);
or U2541 (N_2541,N_1708,N_1501);
and U2542 (N_2542,N_1867,N_1727);
or U2543 (N_2543,N_1117,N_1470);
nor U2544 (N_2544,N_1095,N_1992);
nor U2545 (N_2545,N_1710,N_1347);
nor U2546 (N_2546,N_1043,N_1364);
or U2547 (N_2547,N_1241,N_1666);
nand U2548 (N_2548,N_1112,N_1992);
and U2549 (N_2549,N_1707,N_1049);
nor U2550 (N_2550,N_1946,N_1852);
xor U2551 (N_2551,N_1525,N_1457);
and U2552 (N_2552,N_1642,N_1179);
nand U2553 (N_2553,N_1311,N_1929);
nor U2554 (N_2554,N_1717,N_1217);
nor U2555 (N_2555,N_1220,N_1426);
nor U2556 (N_2556,N_1519,N_1795);
and U2557 (N_2557,N_1378,N_1230);
and U2558 (N_2558,N_1268,N_1291);
or U2559 (N_2559,N_1953,N_1081);
nor U2560 (N_2560,N_1646,N_1803);
nor U2561 (N_2561,N_1429,N_1103);
nor U2562 (N_2562,N_1813,N_1716);
nand U2563 (N_2563,N_1955,N_1426);
nor U2564 (N_2564,N_1545,N_1439);
nor U2565 (N_2565,N_1123,N_1108);
and U2566 (N_2566,N_1901,N_1785);
or U2567 (N_2567,N_1962,N_1491);
or U2568 (N_2568,N_1213,N_1626);
and U2569 (N_2569,N_1521,N_1155);
nor U2570 (N_2570,N_1072,N_1818);
nor U2571 (N_2571,N_1557,N_1968);
or U2572 (N_2572,N_1326,N_1586);
or U2573 (N_2573,N_1726,N_1580);
nand U2574 (N_2574,N_1783,N_1563);
and U2575 (N_2575,N_1755,N_1207);
nor U2576 (N_2576,N_1683,N_1218);
nor U2577 (N_2577,N_1793,N_1220);
or U2578 (N_2578,N_1781,N_1465);
and U2579 (N_2579,N_1422,N_1837);
nand U2580 (N_2580,N_1980,N_1104);
and U2581 (N_2581,N_1775,N_1463);
or U2582 (N_2582,N_1781,N_1266);
and U2583 (N_2583,N_1849,N_1671);
nand U2584 (N_2584,N_1671,N_1443);
nand U2585 (N_2585,N_1765,N_1970);
or U2586 (N_2586,N_1245,N_1061);
nand U2587 (N_2587,N_1331,N_1977);
or U2588 (N_2588,N_1316,N_1875);
nand U2589 (N_2589,N_1347,N_1250);
nor U2590 (N_2590,N_1252,N_1987);
nand U2591 (N_2591,N_1457,N_1147);
or U2592 (N_2592,N_1855,N_1002);
and U2593 (N_2593,N_1905,N_1298);
nand U2594 (N_2594,N_1872,N_1788);
and U2595 (N_2595,N_1906,N_1238);
or U2596 (N_2596,N_1238,N_1000);
nor U2597 (N_2597,N_1841,N_1709);
and U2598 (N_2598,N_1313,N_1382);
or U2599 (N_2599,N_1122,N_1654);
nor U2600 (N_2600,N_1741,N_1496);
and U2601 (N_2601,N_1187,N_1607);
nand U2602 (N_2602,N_1240,N_1208);
or U2603 (N_2603,N_1445,N_1552);
and U2604 (N_2604,N_1302,N_1194);
nand U2605 (N_2605,N_1808,N_1345);
nand U2606 (N_2606,N_1261,N_1337);
and U2607 (N_2607,N_1587,N_1805);
nand U2608 (N_2608,N_1629,N_1087);
or U2609 (N_2609,N_1880,N_1098);
and U2610 (N_2610,N_1813,N_1536);
nand U2611 (N_2611,N_1157,N_1819);
or U2612 (N_2612,N_1733,N_1670);
and U2613 (N_2613,N_1398,N_1339);
or U2614 (N_2614,N_1396,N_1760);
and U2615 (N_2615,N_1720,N_1059);
nand U2616 (N_2616,N_1725,N_1424);
or U2617 (N_2617,N_1902,N_1387);
nor U2618 (N_2618,N_1343,N_1593);
nand U2619 (N_2619,N_1854,N_1999);
nor U2620 (N_2620,N_1564,N_1851);
or U2621 (N_2621,N_1334,N_1526);
or U2622 (N_2622,N_1520,N_1349);
nor U2623 (N_2623,N_1448,N_1179);
or U2624 (N_2624,N_1874,N_1766);
nor U2625 (N_2625,N_1323,N_1396);
nor U2626 (N_2626,N_1280,N_1672);
nor U2627 (N_2627,N_1570,N_1394);
and U2628 (N_2628,N_1872,N_1439);
nand U2629 (N_2629,N_1271,N_1626);
nor U2630 (N_2630,N_1027,N_1328);
nand U2631 (N_2631,N_1136,N_1618);
or U2632 (N_2632,N_1975,N_1042);
and U2633 (N_2633,N_1945,N_1717);
and U2634 (N_2634,N_1072,N_1832);
nand U2635 (N_2635,N_1026,N_1107);
nor U2636 (N_2636,N_1511,N_1052);
nor U2637 (N_2637,N_1593,N_1307);
and U2638 (N_2638,N_1614,N_1026);
nand U2639 (N_2639,N_1533,N_1124);
nor U2640 (N_2640,N_1158,N_1435);
nand U2641 (N_2641,N_1656,N_1693);
and U2642 (N_2642,N_1827,N_1797);
or U2643 (N_2643,N_1949,N_1008);
nand U2644 (N_2644,N_1055,N_1729);
and U2645 (N_2645,N_1692,N_1107);
or U2646 (N_2646,N_1649,N_1014);
nand U2647 (N_2647,N_1010,N_1285);
or U2648 (N_2648,N_1803,N_1130);
nand U2649 (N_2649,N_1819,N_1970);
nor U2650 (N_2650,N_1842,N_1453);
and U2651 (N_2651,N_1602,N_1525);
nor U2652 (N_2652,N_1647,N_1670);
or U2653 (N_2653,N_1752,N_1950);
nor U2654 (N_2654,N_1242,N_1421);
nand U2655 (N_2655,N_1791,N_1027);
nand U2656 (N_2656,N_1305,N_1521);
nand U2657 (N_2657,N_1421,N_1938);
nand U2658 (N_2658,N_1395,N_1563);
nor U2659 (N_2659,N_1418,N_1716);
nor U2660 (N_2660,N_1492,N_1135);
nor U2661 (N_2661,N_1775,N_1711);
nor U2662 (N_2662,N_1484,N_1827);
xor U2663 (N_2663,N_1497,N_1660);
or U2664 (N_2664,N_1257,N_1676);
nand U2665 (N_2665,N_1537,N_1799);
nand U2666 (N_2666,N_1993,N_1007);
or U2667 (N_2667,N_1404,N_1019);
nand U2668 (N_2668,N_1945,N_1321);
nor U2669 (N_2669,N_1236,N_1603);
nor U2670 (N_2670,N_1526,N_1235);
nor U2671 (N_2671,N_1601,N_1704);
and U2672 (N_2672,N_1870,N_1286);
nor U2673 (N_2673,N_1253,N_1166);
nor U2674 (N_2674,N_1324,N_1562);
nor U2675 (N_2675,N_1440,N_1755);
nand U2676 (N_2676,N_1437,N_1438);
and U2677 (N_2677,N_1061,N_1006);
or U2678 (N_2678,N_1852,N_1036);
nor U2679 (N_2679,N_1916,N_1690);
and U2680 (N_2680,N_1614,N_1520);
nor U2681 (N_2681,N_1263,N_1370);
and U2682 (N_2682,N_1183,N_1508);
and U2683 (N_2683,N_1636,N_1588);
nor U2684 (N_2684,N_1309,N_1228);
nor U2685 (N_2685,N_1506,N_1619);
nand U2686 (N_2686,N_1242,N_1826);
or U2687 (N_2687,N_1784,N_1007);
nand U2688 (N_2688,N_1178,N_1770);
and U2689 (N_2689,N_1771,N_1053);
and U2690 (N_2690,N_1171,N_1674);
and U2691 (N_2691,N_1119,N_1491);
nor U2692 (N_2692,N_1461,N_1816);
nor U2693 (N_2693,N_1256,N_1925);
nand U2694 (N_2694,N_1625,N_1767);
xnor U2695 (N_2695,N_1285,N_1971);
and U2696 (N_2696,N_1460,N_1044);
nor U2697 (N_2697,N_1656,N_1660);
or U2698 (N_2698,N_1570,N_1908);
nor U2699 (N_2699,N_1803,N_1879);
nor U2700 (N_2700,N_1169,N_1355);
and U2701 (N_2701,N_1646,N_1120);
nand U2702 (N_2702,N_1699,N_1452);
xnor U2703 (N_2703,N_1960,N_1584);
nor U2704 (N_2704,N_1689,N_1992);
or U2705 (N_2705,N_1252,N_1844);
or U2706 (N_2706,N_1989,N_1108);
and U2707 (N_2707,N_1084,N_1367);
nand U2708 (N_2708,N_1821,N_1720);
or U2709 (N_2709,N_1503,N_1604);
or U2710 (N_2710,N_1173,N_1852);
nand U2711 (N_2711,N_1137,N_1590);
nand U2712 (N_2712,N_1828,N_1090);
nand U2713 (N_2713,N_1788,N_1571);
nor U2714 (N_2714,N_1252,N_1667);
nor U2715 (N_2715,N_1317,N_1110);
and U2716 (N_2716,N_1334,N_1668);
nor U2717 (N_2717,N_1517,N_1626);
nor U2718 (N_2718,N_1251,N_1711);
nor U2719 (N_2719,N_1294,N_1427);
or U2720 (N_2720,N_1543,N_1473);
or U2721 (N_2721,N_1121,N_1042);
and U2722 (N_2722,N_1498,N_1800);
or U2723 (N_2723,N_1585,N_1697);
and U2724 (N_2724,N_1528,N_1082);
or U2725 (N_2725,N_1053,N_1135);
nor U2726 (N_2726,N_1144,N_1633);
or U2727 (N_2727,N_1911,N_1204);
or U2728 (N_2728,N_1257,N_1601);
nand U2729 (N_2729,N_1916,N_1412);
or U2730 (N_2730,N_1428,N_1549);
nand U2731 (N_2731,N_1248,N_1791);
nor U2732 (N_2732,N_1645,N_1598);
or U2733 (N_2733,N_1350,N_1695);
and U2734 (N_2734,N_1482,N_1967);
nor U2735 (N_2735,N_1310,N_1511);
nand U2736 (N_2736,N_1226,N_1608);
and U2737 (N_2737,N_1073,N_1077);
nor U2738 (N_2738,N_1277,N_1054);
nor U2739 (N_2739,N_1421,N_1263);
nand U2740 (N_2740,N_1203,N_1141);
nand U2741 (N_2741,N_1759,N_1632);
nor U2742 (N_2742,N_1736,N_1546);
or U2743 (N_2743,N_1417,N_1038);
nor U2744 (N_2744,N_1427,N_1531);
and U2745 (N_2745,N_1214,N_1189);
nor U2746 (N_2746,N_1787,N_1550);
nand U2747 (N_2747,N_1988,N_1808);
and U2748 (N_2748,N_1755,N_1146);
nor U2749 (N_2749,N_1556,N_1019);
or U2750 (N_2750,N_1899,N_1447);
nand U2751 (N_2751,N_1195,N_1859);
and U2752 (N_2752,N_1478,N_1719);
and U2753 (N_2753,N_1372,N_1567);
or U2754 (N_2754,N_1560,N_1599);
nand U2755 (N_2755,N_1643,N_1763);
or U2756 (N_2756,N_1922,N_1904);
and U2757 (N_2757,N_1805,N_1007);
nor U2758 (N_2758,N_1230,N_1281);
nand U2759 (N_2759,N_1259,N_1882);
and U2760 (N_2760,N_1791,N_1058);
or U2761 (N_2761,N_1099,N_1795);
and U2762 (N_2762,N_1588,N_1779);
nand U2763 (N_2763,N_1445,N_1182);
and U2764 (N_2764,N_1446,N_1322);
or U2765 (N_2765,N_1724,N_1284);
and U2766 (N_2766,N_1212,N_1646);
and U2767 (N_2767,N_1491,N_1079);
nor U2768 (N_2768,N_1622,N_1281);
and U2769 (N_2769,N_1443,N_1367);
nor U2770 (N_2770,N_1849,N_1384);
and U2771 (N_2771,N_1914,N_1493);
nor U2772 (N_2772,N_1568,N_1868);
nor U2773 (N_2773,N_1904,N_1263);
or U2774 (N_2774,N_1961,N_1819);
nand U2775 (N_2775,N_1646,N_1326);
xnor U2776 (N_2776,N_1938,N_1600);
or U2777 (N_2777,N_1642,N_1602);
and U2778 (N_2778,N_1995,N_1362);
nor U2779 (N_2779,N_1277,N_1426);
nand U2780 (N_2780,N_1297,N_1100);
nor U2781 (N_2781,N_1759,N_1018);
nand U2782 (N_2782,N_1728,N_1575);
xnor U2783 (N_2783,N_1152,N_1627);
nor U2784 (N_2784,N_1774,N_1554);
or U2785 (N_2785,N_1485,N_1321);
and U2786 (N_2786,N_1930,N_1899);
xnor U2787 (N_2787,N_1317,N_1569);
nand U2788 (N_2788,N_1932,N_1196);
nand U2789 (N_2789,N_1555,N_1235);
nor U2790 (N_2790,N_1176,N_1797);
nor U2791 (N_2791,N_1884,N_1787);
or U2792 (N_2792,N_1952,N_1556);
nor U2793 (N_2793,N_1409,N_1341);
or U2794 (N_2794,N_1571,N_1594);
nor U2795 (N_2795,N_1827,N_1263);
and U2796 (N_2796,N_1875,N_1850);
nand U2797 (N_2797,N_1363,N_1170);
and U2798 (N_2798,N_1160,N_1197);
nor U2799 (N_2799,N_1734,N_1259);
or U2800 (N_2800,N_1105,N_1319);
xnor U2801 (N_2801,N_1448,N_1630);
or U2802 (N_2802,N_1247,N_1920);
nor U2803 (N_2803,N_1849,N_1861);
and U2804 (N_2804,N_1889,N_1061);
nor U2805 (N_2805,N_1026,N_1774);
or U2806 (N_2806,N_1868,N_1438);
or U2807 (N_2807,N_1615,N_1453);
or U2808 (N_2808,N_1151,N_1106);
or U2809 (N_2809,N_1463,N_1886);
and U2810 (N_2810,N_1734,N_1412);
nor U2811 (N_2811,N_1847,N_1392);
or U2812 (N_2812,N_1411,N_1885);
or U2813 (N_2813,N_1171,N_1979);
and U2814 (N_2814,N_1220,N_1212);
nor U2815 (N_2815,N_1016,N_1417);
or U2816 (N_2816,N_1071,N_1446);
or U2817 (N_2817,N_1398,N_1793);
nor U2818 (N_2818,N_1342,N_1038);
nor U2819 (N_2819,N_1702,N_1840);
and U2820 (N_2820,N_1819,N_1031);
nor U2821 (N_2821,N_1751,N_1406);
or U2822 (N_2822,N_1109,N_1386);
nand U2823 (N_2823,N_1771,N_1427);
or U2824 (N_2824,N_1971,N_1678);
or U2825 (N_2825,N_1493,N_1528);
or U2826 (N_2826,N_1634,N_1749);
nand U2827 (N_2827,N_1766,N_1322);
nor U2828 (N_2828,N_1964,N_1552);
nor U2829 (N_2829,N_1491,N_1442);
nor U2830 (N_2830,N_1657,N_1507);
nand U2831 (N_2831,N_1625,N_1760);
nor U2832 (N_2832,N_1520,N_1480);
nor U2833 (N_2833,N_1206,N_1375);
or U2834 (N_2834,N_1685,N_1875);
or U2835 (N_2835,N_1332,N_1075);
nor U2836 (N_2836,N_1448,N_1875);
or U2837 (N_2837,N_1882,N_1713);
and U2838 (N_2838,N_1332,N_1435);
nor U2839 (N_2839,N_1762,N_1112);
nand U2840 (N_2840,N_1660,N_1045);
and U2841 (N_2841,N_1413,N_1593);
or U2842 (N_2842,N_1027,N_1195);
nand U2843 (N_2843,N_1307,N_1484);
nand U2844 (N_2844,N_1682,N_1533);
and U2845 (N_2845,N_1189,N_1670);
or U2846 (N_2846,N_1341,N_1806);
nor U2847 (N_2847,N_1214,N_1367);
or U2848 (N_2848,N_1652,N_1409);
nor U2849 (N_2849,N_1335,N_1095);
or U2850 (N_2850,N_1488,N_1380);
nor U2851 (N_2851,N_1348,N_1805);
nor U2852 (N_2852,N_1387,N_1094);
nand U2853 (N_2853,N_1860,N_1931);
and U2854 (N_2854,N_1706,N_1268);
or U2855 (N_2855,N_1311,N_1284);
or U2856 (N_2856,N_1911,N_1957);
nor U2857 (N_2857,N_1670,N_1088);
nand U2858 (N_2858,N_1388,N_1067);
nor U2859 (N_2859,N_1764,N_1181);
nor U2860 (N_2860,N_1287,N_1106);
nor U2861 (N_2861,N_1948,N_1896);
and U2862 (N_2862,N_1166,N_1186);
nor U2863 (N_2863,N_1506,N_1557);
or U2864 (N_2864,N_1092,N_1992);
nor U2865 (N_2865,N_1163,N_1199);
nand U2866 (N_2866,N_1210,N_1528);
or U2867 (N_2867,N_1343,N_1238);
nor U2868 (N_2868,N_1326,N_1012);
nor U2869 (N_2869,N_1072,N_1602);
nor U2870 (N_2870,N_1083,N_1534);
or U2871 (N_2871,N_1086,N_1867);
nor U2872 (N_2872,N_1420,N_1430);
nor U2873 (N_2873,N_1398,N_1528);
nand U2874 (N_2874,N_1800,N_1255);
nand U2875 (N_2875,N_1651,N_1905);
or U2876 (N_2876,N_1434,N_1518);
and U2877 (N_2877,N_1286,N_1989);
nor U2878 (N_2878,N_1478,N_1807);
nand U2879 (N_2879,N_1529,N_1769);
and U2880 (N_2880,N_1021,N_1906);
and U2881 (N_2881,N_1235,N_1583);
and U2882 (N_2882,N_1585,N_1140);
or U2883 (N_2883,N_1679,N_1379);
and U2884 (N_2884,N_1881,N_1612);
nand U2885 (N_2885,N_1706,N_1424);
nand U2886 (N_2886,N_1890,N_1009);
and U2887 (N_2887,N_1251,N_1223);
or U2888 (N_2888,N_1663,N_1405);
or U2889 (N_2889,N_1085,N_1890);
nor U2890 (N_2890,N_1259,N_1191);
or U2891 (N_2891,N_1862,N_1414);
and U2892 (N_2892,N_1509,N_1083);
nor U2893 (N_2893,N_1829,N_1775);
nor U2894 (N_2894,N_1250,N_1280);
and U2895 (N_2895,N_1903,N_1935);
nor U2896 (N_2896,N_1631,N_1404);
nor U2897 (N_2897,N_1164,N_1074);
or U2898 (N_2898,N_1765,N_1020);
nand U2899 (N_2899,N_1935,N_1566);
or U2900 (N_2900,N_1450,N_1580);
nor U2901 (N_2901,N_1351,N_1504);
or U2902 (N_2902,N_1112,N_1592);
and U2903 (N_2903,N_1471,N_1688);
and U2904 (N_2904,N_1572,N_1821);
and U2905 (N_2905,N_1468,N_1770);
or U2906 (N_2906,N_1556,N_1502);
nor U2907 (N_2907,N_1752,N_1993);
xnor U2908 (N_2908,N_1877,N_1113);
nand U2909 (N_2909,N_1141,N_1974);
or U2910 (N_2910,N_1485,N_1198);
or U2911 (N_2911,N_1360,N_1176);
nor U2912 (N_2912,N_1996,N_1567);
and U2913 (N_2913,N_1513,N_1335);
or U2914 (N_2914,N_1088,N_1153);
nor U2915 (N_2915,N_1346,N_1476);
nor U2916 (N_2916,N_1358,N_1153);
or U2917 (N_2917,N_1157,N_1123);
nor U2918 (N_2918,N_1502,N_1352);
and U2919 (N_2919,N_1747,N_1109);
or U2920 (N_2920,N_1857,N_1262);
nor U2921 (N_2921,N_1151,N_1294);
nand U2922 (N_2922,N_1770,N_1092);
nor U2923 (N_2923,N_1975,N_1709);
nand U2924 (N_2924,N_1570,N_1835);
and U2925 (N_2925,N_1791,N_1040);
or U2926 (N_2926,N_1079,N_1259);
and U2927 (N_2927,N_1150,N_1098);
or U2928 (N_2928,N_1876,N_1860);
or U2929 (N_2929,N_1862,N_1686);
and U2930 (N_2930,N_1709,N_1531);
or U2931 (N_2931,N_1390,N_1983);
nor U2932 (N_2932,N_1919,N_1922);
nand U2933 (N_2933,N_1891,N_1838);
nor U2934 (N_2934,N_1559,N_1767);
nor U2935 (N_2935,N_1414,N_1306);
nand U2936 (N_2936,N_1583,N_1154);
and U2937 (N_2937,N_1152,N_1827);
nand U2938 (N_2938,N_1914,N_1570);
and U2939 (N_2939,N_1571,N_1378);
or U2940 (N_2940,N_1795,N_1033);
nor U2941 (N_2941,N_1513,N_1751);
nor U2942 (N_2942,N_1274,N_1421);
nor U2943 (N_2943,N_1894,N_1547);
or U2944 (N_2944,N_1958,N_1530);
nor U2945 (N_2945,N_1240,N_1003);
nor U2946 (N_2946,N_1656,N_1024);
or U2947 (N_2947,N_1314,N_1249);
or U2948 (N_2948,N_1509,N_1882);
or U2949 (N_2949,N_1918,N_1322);
nand U2950 (N_2950,N_1634,N_1710);
nor U2951 (N_2951,N_1476,N_1511);
and U2952 (N_2952,N_1703,N_1588);
nand U2953 (N_2953,N_1057,N_1595);
and U2954 (N_2954,N_1173,N_1218);
and U2955 (N_2955,N_1453,N_1647);
nor U2956 (N_2956,N_1129,N_1615);
nor U2957 (N_2957,N_1599,N_1569);
or U2958 (N_2958,N_1004,N_1118);
and U2959 (N_2959,N_1543,N_1313);
nor U2960 (N_2960,N_1079,N_1410);
and U2961 (N_2961,N_1650,N_1293);
or U2962 (N_2962,N_1953,N_1494);
or U2963 (N_2963,N_1285,N_1129);
nor U2964 (N_2964,N_1305,N_1484);
nor U2965 (N_2965,N_1853,N_1672);
or U2966 (N_2966,N_1955,N_1960);
or U2967 (N_2967,N_1406,N_1377);
or U2968 (N_2968,N_1589,N_1998);
nand U2969 (N_2969,N_1259,N_1589);
nor U2970 (N_2970,N_1236,N_1628);
or U2971 (N_2971,N_1942,N_1861);
nand U2972 (N_2972,N_1581,N_1863);
nor U2973 (N_2973,N_1936,N_1878);
nor U2974 (N_2974,N_1373,N_1061);
nor U2975 (N_2975,N_1145,N_1886);
nand U2976 (N_2976,N_1680,N_1664);
and U2977 (N_2977,N_1622,N_1681);
nor U2978 (N_2978,N_1463,N_1451);
nand U2979 (N_2979,N_1609,N_1400);
nand U2980 (N_2980,N_1209,N_1575);
nor U2981 (N_2981,N_1849,N_1092);
nor U2982 (N_2982,N_1105,N_1128);
or U2983 (N_2983,N_1177,N_1050);
and U2984 (N_2984,N_1013,N_1918);
nand U2985 (N_2985,N_1336,N_1919);
or U2986 (N_2986,N_1145,N_1624);
nor U2987 (N_2987,N_1470,N_1105);
nor U2988 (N_2988,N_1012,N_1318);
or U2989 (N_2989,N_1603,N_1086);
and U2990 (N_2990,N_1768,N_1993);
and U2991 (N_2991,N_1320,N_1048);
or U2992 (N_2992,N_1564,N_1979);
or U2993 (N_2993,N_1039,N_1565);
nand U2994 (N_2994,N_1480,N_1139);
and U2995 (N_2995,N_1868,N_1891);
or U2996 (N_2996,N_1325,N_1012);
and U2997 (N_2997,N_1055,N_1169);
nor U2998 (N_2998,N_1289,N_1462);
or U2999 (N_2999,N_1928,N_1064);
nand U3000 (N_3000,N_2766,N_2932);
nand U3001 (N_3001,N_2794,N_2456);
or U3002 (N_3002,N_2300,N_2645);
nand U3003 (N_3003,N_2542,N_2966);
nor U3004 (N_3004,N_2102,N_2910);
and U3005 (N_3005,N_2942,N_2013);
and U3006 (N_3006,N_2527,N_2577);
or U3007 (N_3007,N_2959,N_2851);
and U3008 (N_3008,N_2051,N_2607);
nor U3009 (N_3009,N_2280,N_2676);
nand U3010 (N_3010,N_2134,N_2435);
nand U3011 (N_3011,N_2546,N_2222);
nand U3012 (N_3012,N_2889,N_2681);
nor U3013 (N_3013,N_2077,N_2457);
nor U3014 (N_3014,N_2193,N_2253);
or U3015 (N_3015,N_2376,N_2005);
nand U3016 (N_3016,N_2985,N_2621);
nor U3017 (N_3017,N_2083,N_2793);
nor U3018 (N_3018,N_2273,N_2266);
or U3019 (N_3019,N_2707,N_2170);
and U3020 (N_3020,N_2229,N_2437);
nor U3021 (N_3021,N_2143,N_2439);
and U3022 (N_3022,N_2117,N_2241);
or U3023 (N_3023,N_2238,N_2227);
nor U3024 (N_3024,N_2294,N_2570);
and U3025 (N_3025,N_2832,N_2425);
or U3026 (N_3026,N_2200,N_2423);
and U3027 (N_3027,N_2606,N_2781);
and U3028 (N_3028,N_2902,N_2798);
nor U3029 (N_3029,N_2130,N_2509);
nor U3030 (N_3030,N_2878,N_2993);
nand U3031 (N_3031,N_2672,N_2937);
and U3032 (N_3032,N_2328,N_2353);
or U3033 (N_3033,N_2112,N_2689);
and U3034 (N_3034,N_2311,N_2014);
nor U3035 (N_3035,N_2345,N_2086);
and U3036 (N_3036,N_2740,N_2520);
xor U3037 (N_3037,N_2825,N_2669);
or U3038 (N_3038,N_2374,N_2250);
nor U3039 (N_3039,N_2749,N_2033);
or U3040 (N_3040,N_2135,N_2743);
nand U3041 (N_3041,N_2898,N_2507);
or U3042 (N_3042,N_2493,N_2792);
or U3043 (N_3043,N_2692,N_2747);
or U3044 (N_3044,N_2020,N_2009);
and U3045 (N_3045,N_2583,N_2189);
nor U3046 (N_3046,N_2239,N_2429);
and U3047 (N_3047,N_2268,N_2956);
nand U3048 (N_3048,N_2442,N_2325);
nand U3049 (N_3049,N_2615,N_2305);
or U3050 (N_3050,N_2110,N_2525);
nor U3051 (N_3051,N_2221,N_2500);
nand U3052 (N_3052,N_2824,N_2141);
nand U3053 (N_3053,N_2834,N_2626);
or U3054 (N_3054,N_2962,N_2999);
or U3055 (N_3055,N_2058,N_2516);
nand U3056 (N_3056,N_2714,N_2183);
nor U3057 (N_3057,N_2697,N_2225);
nand U3058 (N_3058,N_2984,N_2533);
and U3059 (N_3059,N_2441,N_2719);
and U3060 (N_3060,N_2981,N_2003);
and U3061 (N_3061,N_2177,N_2124);
or U3062 (N_3062,N_2201,N_2826);
nor U3063 (N_3063,N_2796,N_2675);
and U3064 (N_3064,N_2769,N_2330);
or U3065 (N_3065,N_2031,N_2436);
nand U3066 (N_3066,N_2819,N_2145);
nand U3067 (N_3067,N_2568,N_2945);
or U3068 (N_3068,N_2599,N_2363);
nor U3069 (N_3069,N_2257,N_2059);
nand U3070 (N_3070,N_2006,N_2562);
or U3071 (N_3071,N_2677,N_2730);
nor U3072 (N_3072,N_2858,N_2590);
nand U3073 (N_3073,N_2987,N_2641);
nand U3074 (N_3074,N_2162,N_2139);
nand U3075 (N_3075,N_2592,N_2256);
or U3076 (N_3076,N_2195,N_2775);
and U3077 (N_3077,N_2099,N_2665);
nor U3078 (N_3078,N_2404,N_2365);
or U3079 (N_3079,N_2283,N_2630);
nand U3080 (N_3080,N_2119,N_2847);
and U3081 (N_3081,N_2960,N_2165);
and U3082 (N_3082,N_2089,N_2354);
and U3083 (N_3083,N_2440,N_2887);
and U3084 (N_3084,N_2382,N_2424);
nor U3085 (N_3085,N_2232,N_2275);
nand U3086 (N_3086,N_2093,N_2398);
or U3087 (N_3087,N_2657,N_2973);
and U3088 (N_3088,N_2835,N_2136);
nand U3089 (N_3089,N_2282,N_2808);
nand U3090 (N_3090,N_2073,N_2394);
nor U3091 (N_3091,N_2434,N_2510);
nor U3092 (N_3092,N_2048,N_2385);
nor U3093 (N_3093,N_2062,N_2197);
nand U3094 (N_3094,N_2748,N_2968);
or U3095 (N_3095,N_2652,N_2414);
or U3096 (N_3096,N_2355,N_2701);
nor U3097 (N_3097,N_2067,N_2741);
and U3098 (N_3098,N_2478,N_2762);
nand U3099 (N_3099,N_2420,N_2705);
and U3100 (N_3100,N_2421,N_2632);
nor U3101 (N_3101,N_2074,N_2184);
or U3102 (N_3102,N_2799,N_2380);
and U3103 (N_3103,N_2773,N_2674);
nor U3104 (N_3104,N_2446,N_2349);
nor U3105 (N_3105,N_2377,N_2765);
and U3106 (N_3106,N_2471,N_2894);
or U3107 (N_3107,N_2584,N_2848);
and U3108 (N_3108,N_2347,N_2767);
and U3109 (N_3109,N_2597,N_2078);
nand U3110 (N_3110,N_2501,N_2123);
or U3111 (N_3111,N_2523,N_2503);
or U3112 (N_3112,N_2179,N_2742);
or U3113 (N_3113,N_2274,N_2155);
and U3114 (N_3114,N_2933,N_2928);
nor U3115 (N_3115,N_2053,N_2426);
nand U3116 (N_3116,N_2302,N_2369);
nor U3117 (N_3117,N_2589,N_2978);
or U3118 (N_3118,N_2109,N_2696);
and U3119 (N_3119,N_2821,N_2567);
nand U3120 (N_3120,N_2277,N_2852);
or U3121 (N_3121,N_2843,N_2718);
nor U3122 (N_3122,N_2327,N_2759);
nor U3123 (N_3123,N_2097,N_2656);
and U3124 (N_3124,N_2463,N_2983);
nor U3125 (N_3125,N_2359,N_2151);
nand U3126 (N_3126,N_2941,N_2194);
nor U3127 (N_3127,N_2254,N_2484);
nand U3128 (N_3128,N_2921,N_2288);
nand U3129 (N_3129,N_2367,N_2691);
nand U3130 (N_3130,N_2737,N_2116);
and U3131 (N_3131,N_2559,N_2723);
or U3132 (N_3132,N_2512,N_2764);
and U3133 (N_3133,N_2337,N_2455);
nand U3134 (N_3134,N_2829,N_2498);
nor U3135 (N_3135,N_2133,N_2447);
nand U3136 (N_3136,N_2923,N_2903);
or U3137 (N_3137,N_2344,N_2042);
nand U3138 (N_3138,N_2017,N_2870);
nor U3139 (N_3139,N_2223,N_2160);
nand U3140 (N_3140,N_2506,N_2205);
nand U3141 (N_3141,N_2602,N_2536);
or U3142 (N_3142,N_2244,N_2866);
nand U3143 (N_3143,N_2298,N_2057);
and U3144 (N_3144,N_2336,N_2880);
or U3145 (N_3145,N_2443,N_2988);
and U3146 (N_3146,N_2087,N_2040);
nand U3147 (N_3147,N_2576,N_2678);
nand U3148 (N_3148,N_2948,N_2936);
nor U3149 (N_3149,N_2018,N_2303);
or U3150 (N_3150,N_2855,N_2432);
and U3151 (N_3151,N_2026,N_2373);
nor U3152 (N_3152,N_2248,N_2638);
and U3153 (N_3153,N_2085,N_2531);
nand U3154 (N_3154,N_2998,N_2056);
and U3155 (N_3155,N_2156,N_2857);
or U3156 (N_3156,N_2909,N_2381);
nor U3157 (N_3157,N_2846,N_2322);
nand U3158 (N_3158,N_2296,N_2472);
and U3159 (N_3159,N_2905,N_2636);
nand U3160 (N_3160,N_2529,N_2515);
nand U3161 (N_3161,N_2012,N_2395);
or U3162 (N_3162,N_2480,N_2571);
or U3163 (N_3163,N_2594,N_2845);
nand U3164 (N_3164,N_2668,N_2886);
nand U3165 (N_3165,N_2551,N_2240);
nor U3166 (N_3166,N_2650,N_2262);
and U3167 (N_3167,N_2947,N_2617);
nand U3168 (N_3168,N_2735,N_2708);
and U3169 (N_3169,N_2098,N_2154);
and U3170 (N_3170,N_2348,N_2791);
or U3171 (N_3171,N_2451,N_2784);
nor U3172 (N_3172,N_2153,N_2895);
nor U3173 (N_3173,N_2408,N_2137);
nor U3174 (N_3174,N_2548,N_2150);
or U3175 (N_3175,N_2315,N_2532);
and U3176 (N_3176,N_2164,N_2586);
nand U3177 (N_3177,N_2623,N_2655);
or U3178 (N_3178,N_2545,N_2561);
nor U3179 (N_3179,N_2182,N_2579);
nor U3180 (N_3180,N_2263,N_2445);
nor U3181 (N_3181,N_2514,N_2259);
or U3182 (N_3182,N_2483,N_2982);
or U3183 (N_3183,N_2663,N_2739);
or U3184 (N_3184,N_2490,N_2949);
or U3185 (N_3185,N_2543,N_2030);
and U3186 (N_3186,N_2768,N_2476);
nor U3187 (N_3187,N_2756,N_2528);
and U3188 (N_3188,N_2066,N_2706);
nand U3189 (N_3189,N_2482,N_2412);
nor U3190 (N_3190,N_2774,N_2831);
and U3191 (N_3191,N_2535,N_2169);
nand U3192 (N_3192,N_2861,N_2486);
nor U3193 (N_3193,N_2777,N_2856);
or U3194 (N_3194,N_2470,N_2897);
and U3195 (N_3195,N_2564,N_2350);
nand U3196 (N_3196,N_2011,N_2815);
and U3197 (N_3197,N_2913,N_2438);
and U3198 (N_3198,N_2301,N_2876);
and U3199 (N_3199,N_2402,N_2753);
and U3200 (N_3200,N_2967,N_2215);
nand U3201 (N_3201,N_2297,N_2310);
nor U3202 (N_3202,N_2635,N_2497);
or U3203 (N_3203,N_2024,N_2260);
nor U3204 (N_3204,N_2771,N_2530);
nand U3205 (N_3205,N_2547,N_2001);
nand U3206 (N_3206,N_2969,N_2991);
nor U3207 (N_3207,N_2734,N_2392);
nand U3208 (N_3208,N_2499,N_2433);
nor U3209 (N_3209,N_2877,N_2035);
nand U3210 (N_3210,N_2292,N_2218);
nor U3211 (N_3211,N_2469,N_2495);
and U3212 (N_3212,N_2849,N_2859);
and U3213 (N_3213,N_2752,N_2906);
nor U3214 (N_3214,N_2710,N_2055);
nor U3215 (N_3215,N_2795,N_2744);
and U3216 (N_3216,N_2673,N_2558);
or U3217 (N_3217,N_2658,N_2252);
and U3218 (N_3218,N_2027,N_2128);
nand U3219 (N_3219,N_2574,N_2619);
or U3220 (N_3220,N_2094,N_2299);
nand U3221 (N_3221,N_2122,N_2401);
nor U3222 (N_3222,N_2549,N_2780);
or U3223 (N_3223,N_2521,N_2820);
nand U3224 (N_3224,N_2192,N_2582);
or U3225 (N_3225,N_2428,N_2125);
or U3226 (N_3226,N_2068,N_2025);
nor U3227 (N_3227,N_2918,N_2351);
or U3228 (N_3228,N_2338,N_2202);
or U3229 (N_3229,N_2578,N_2550);
or U3230 (N_3230,N_2680,N_2173);
nand U3231 (N_3231,N_2092,N_2639);
nand U3232 (N_3232,N_2148,N_2272);
nand U3233 (N_3233,N_2776,N_2721);
or U3234 (N_3234,N_2651,N_2333);
nor U3235 (N_3235,N_2464,N_2335);
nand U3236 (N_3236,N_2778,N_2237);
nand U3237 (N_3237,N_2452,N_2188);
nand U3238 (N_3238,N_2587,N_2511);
and U3239 (N_3239,N_2904,N_2920);
or U3240 (N_3240,N_2841,N_2113);
nand U3241 (N_3241,N_2378,N_2649);
nor U3242 (N_3242,N_2806,N_2801);
or U3243 (N_3243,N_2317,N_2008);
or U3244 (N_3244,N_2994,N_2285);
and U3245 (N_3245,N_2817,N_2647);
or U3246 (N_3246,N_2684,N_2618);
nor U3247 (N_3247,N_2196,N_2295);
nor U3248 (N_3248,N_2611,N_2726);
nor U3249 (N_3249,N_2996,N_2409);
nor U3250 (N_3250,N_2002,N_2209);
nor U3251 (N_3251,N_2612,N_2388);
or U3252 (N_3252,N_2290,N_2271);
or U3253 (N_3253,N_2037,N_2213);
nor U3254 (N_3254,N_2888,N_2308);
and U3255 (N_3255,N_2935,N_2076);
nor U3256 (N_3256,N_2938,N_2236);
or U3257 (N_3257,N_2247,N_2468);
nor U3258 (N_3258,N_2811,N_2211);
or U3259 (N_3259,N_2450,N_2419);
nor U3260 (N_3260,N_2276,N_2961);
nor U3261 (N_3261,N_2041,N_2802);
and U3262 (N_3262,N_2823,N_2867);
and U3263 (N_3263,N_2724,N_2390);
nand U3264 (N_3264,N_2810,N_2807);
nand U3265 (N_3265,N_2812,N_2990);
nand U3266 (N_3266,N_2770,N_2624);
nand U3267 (N_3267,N_2838,N_2963);
nor U3268 (N_3268,N_2896,N_2270);
or U3269 (N_3269,N_2608,N_2943);
nand U3270 (N_3270,N_2517,N_2627);
nand U3271 (N_3271,N_2716,N_2406);
or U3272 (N_3272,N_2258,N_2603);
xnor U3273 (N_3273,N_2403,N_2324);
and U3274 (N_3274,N_2953,N_2036);
or U3275 (N_3275,N_2459,N_2204);
or U3276 (N_3276,N_2473,N_2703);
nor U3277 (N_3277,N_2871,N_2717);
nor U3278 (N_3278,N_2108,N_2989);
nand U3279 (N_3279,N_2465,N_2900);
nand U3280 (N_3280,N_2107,N_2699);
or U3281 (N_3281,N_2163,N_2595);
and U3282 (N_3282,N_2518,N_2600);
nand U3283 (N_3283,N_2954,N_2126);
or U3284 (N_3284,N_2371,N_2788);
nor U3285 (N_3285,N_2720,N_2032);
or U3286 (N_3286,N_2782,N_2090);
nand U3287 (N_3287,N_2760,N_2581);
and U3288 (N_3288,N_2569,N_2418);
and U3289 (N_3289,N_2563,N_2265);
and U3290 (N_3290,N_2732,N_2103);
and U3291 (N_3291,N_2049,N_2477);
nand U3292 (N_3292,N_2422,N_2683);
and U3293 (N_3293,N_2178,N_2946);
and U3294 (N_3294,N_2513,N_2269);
and U3295 (N_3295,N_2833,N_2341);
and U3296 (N_3296,N_2079,N_2131);
nor U3297 (N_3297,N_2844,N_2364);
nand U3298 (N_3298,N_2757,N_2411);
and U3299 (N_3299,N_2198,N_2924);
and U3300 (N_3300,N_2487,N_2475);
nor U3301 (N_3301,N_2679,N_2115);
nor U3302 (N_3302,N_2565,N_2659);
nor U3303 (N_3303,N_2485,N_2105);
nand U3304 (N_3304,N_2264,N_2454);
nor U3305 (N_3305,N_2181,N_2000);
or U3306 (N_3306,N_2316,N_2736);
nor U3307 (N_3307,N_2940,N_2916);
nand U3308 (N_3308,N_2572,N_2854);
nand U3309 (N_3309,N_2023,N_2755);
and U3310 (N_3310,N_2648,N_2286);
and U3311 (N_3311,N_2687,N_2929);
or U3312 (N_3312,N_2144,N_2199);
and U3313 (N_3313,N_2063,N_2029);
and U3314 (N_3314,N_2491,N_2343);
nor U3315 (N_3315,N_2702,N_2357);
nand U3316 (N_3316,N_2539,N_2502);
nor U3317 (N_3317,N_2214,N_2800);
and U3318 (N_3318,N_2964,N_2553);
nor U3319 (N_3319,N_2329,N_2175);
or U3320 (N_3320,N_2167,N_2901);
nand U3321 (N_3321,N_2671,N_2604);
nor U3322 (N_3322,N_2114,N_2111);
and U3323 (N_3323,N_2952,N_2187);
nand U3324 (N_3324,N_2084,N_2761);
nand U3325 (N_3325,N_2206,N_2789);
and U3326 (N_3326,N_2415,N_2082);
nor U3327 (N_3327,N_2142,N_2171);
and U3328 (N_3328,N_2389,N_2120);
nor U3329 (N_3329,N_2416,N_2152);
nor U3330 (N_3330,N_2230,N_2400);
nand U3331 (N_3331,N_2462,N_2289);
nand U3332 (N_3332,N_2267,N_2814);
and U3333 (N_3333,N_2556,N_2862);
or U3334 (N_3334,N_2346,N_2284);
and U3335 (N_3335,N_2786,N_2908);
or U3336 (N_3336,N_2631,N_2869);
or U3337 (N_3337,N_2883,N_2479);
nand U3338 (N_3338,N_2207,N_2190);
nor U3339 (N_3339,N_2809,N_2830);
and U3340 (N_3340,N_2922,N_2874);
xnor U3341 (N_3341,N_2541,N_2504);
and U3342 (N_3342,N_2427,N_2226);
and U3343 (N_3343,N_2596,N_2186);
nor U3344 (N_3344,N_2593,N_2004);
and U3345 (N_3345,N_2321,N_2772);
nor U3346 (N_3346,N_2712,N_2925);
nand U3347 (N_3347,N_2879,N_2839);
and U3348 (N_3348,N_2616,N_2505);
nand U3349 (N_3349,N_2104,N_2914);
nand U3350 (N_3350,N_2287,N_2955);
nand U3351 (N_3351,N_2816,N_2080);
or U3352 (N_3352,N_2050,N_2931);
nor U3353 (N_3353,N_2965,N_2368);
nor U3354 (N_3354,N_2733,N_2711);
nor U3355 (N_3355,N_2233,N_2361);
or U3356 (N_3356,N_2970,N_2243);
nor U3357 (N_3357,N_2166,N_2660);
nor U3358 (N_3358,N_2637,N_2410);
or U3359 (N_3359,N_2557,N_2646);
and U3360 (N_3360,N_2091,N_2172);
and U3361 (N_3361,N_2304,N_2065);
nand U3362 (N_3362,N_2613,N_2944);
nand U3363 (N_3363,N_2822,N_2850);
nand U3364 (N_3364,N_2872,N_2670);
nor U3365 (N_3365,N_2804,N_2890);
nor U3366 (N_3366,N_2360,N_2974);
or U3367 (N_3367,N_2106,N_2088);
nand U3368 (N_3368,N_2912,N_2957);
nand U3369 (N_3369,N_2458,N_2149);
nor U3370 (N_3370,N_2038,N_2314);
nand U3371 (N_3371,N_2666,N_2661);
and U3372 (N_3372,N_2161,N_2339);
and U3373 (N_3373,N_2185,N_2016);
and U3374 (N_3374,N_2840,N_2580);
nand U3375 (N_3375,N_2245,N_2951);
nand U3376 (N_3376,N_2694,N_2598);
or U3377 (N_3377,N_2309,N_2601);
nor U3378 (N_3378,N_2234,N_2555);
nor U3379 (N_3379,N_2803,N_2654);
nand U3380 (N_3380,N_2827,N_2045);
or U3381 (N_3381,N_2728,N_2047);
or U3382 (N_3382,N_2007,N_2892);
nand U3383 (N_3383,N_2386,N_2640);
nor U3384 (N_3384,N_2837,N_2407);
nand U3385 (N_3385,N_2704,N_2934);
and U3386 (N_3386,N_2629,N_2853);
and U3387 (N_3387,N_2882,N_2828);
or U3388 (N_3388,N_2453,N_2358);
nor U3389 (N_3389,N_2127,N_2307);
or U3390 (N_3390,N_2174,N_2069);
or U3391 (N_3391,N_2919,N_2979);
nor U3392 (N_3392,N_2644,N_2915);
or U3393 (N_3393,N_2319,N_2064);
and U3394 (N_3394,N_2071,N_2779);
nand U3395 (N_3395,N_2039,N_2129);
or U3396 (N_3396,N_2818,N_2146);
nor U3397 (N_3397,N_2693,N_2318);
or U3398 (N_3398,N_2334,N_2836);
or U3399 (N_3399,N_2095,N_2231);
and U3400 (N_3400,N_2216,N_2217);
nor U3401 (N_3401,N_2642,N_2034);
nor U3402 (N_3402,N_2397,N_2391);
and U3403 (N_3403,N_2375,N_2797);
and U3404 (N_3404,N_2980,N_2323);
or U3405 (N_3405,N_2538,N_2573);
nand U3406 (N_3406,N_2010,N_2488);
and U3407 (N_3407,N_2413,N_2588);
nor U3408 (N_3408,N_2384,N_2695);
nand U3409 (N_3409,N_2917,N_2713);
nand U3410 (N_3410,N_2899,N_2725);
and U3411 (N_3411,N_2977,N_2868);
nand U3412 (N_3412,N_2246,N_2044);
nand U3413 (N_3413,N_2727,N_2585);
or U3414 (N_3414,N_2790,N_2249);
xor U3415 (N_3415,N_2643,N_2159);
and U3416 (N_3416,N_2865,N_2686);
nor U3417 (N_3417,N_2489,N_2291);
nor U3418 (N_3418,N_2101,N_2927);
and U3419 (N_3419,N_2046,N_2813);
nor U3420 (N_3420,N_2763,N_2634);
and U3421 (N_3421,N_2688,N_2224);
or U3422 (N_3422,N_2907,N_2492);
nand U3423 (N_3423,N_2787,N_2332);
nand U3424 (N_3424,N_2754,N_2387);
nand U3425 (N_3425,N_2995,N_2591);
nor U3426 (N_3426,N_2842,N_2986);
and U3427 (N_3427,N_2210,N_2628);
or U3428 (N_3428,N_2312,N_2015);
and U3429 (N_3429,N_2072,N_2622);
nor U3430 (N_3430,N_2242,N_2605);
nand U3431 (N_3431,N_2208,N_2158);
or U3432 (N_3432,N_2860,N_2331);
nand U3433 (N_3433,N_2560,N_2805);
and U3434 (N_3434,N_2235,N_2519);
nor U3435 (N_3435,N_2203,N_2138);
nand U3436 (N_3436,N_2633,N_2751);
nand U3437 (N_3437,N_2715,N_2522);
nor U3438 (N_3438,N_2132,N_2320);
or U3439 (N_3439,N_2019,N_2971);
nand U3440 (N_3440,N_2534,N_2180);
nor U3441 (N_3441,N_2620,N_2052);
and U3442 (N_3442,N_2746,N_2610);
and U3443 (N_3443,N_2021,N_2460);
and U3444 (N_3444,N_2544,N_2992);
and U3445 (N_3445,N_2372,N_2864);
and U3446 (N_3446,N_2157,N_2625);
nand U3447 (N_3447,N_2251,N_2043);
and U3448 (N_3448,N_2885,N_2494);
and U3449 (N_3449,N_2745,N_2061);
or U3450 (N_3450,N_2508,N_2313);
and U3451 (N_3451,N_2911,N_2191);
or U3452 (N_3452,N_2939,N_2212);
and U3453 (N_3453,N_2340,N_2664);
and U3454 (N_3454,N_2653,N_2405);
nor U3455 (N_3455,N_2417,N_2891);
and U3456 (N_3456,N_2444,N_2575);
or U3457 (N_3457,N_2682,N_2366);
nand U3458 (N_3458,N_2396,N_2958);
nand U3459 (N_3459,N_2750,N_2893);
and U3460 (N_3460,N_2709,N_2100);
and U3461 (N_3461,N_2028,N_2281);
nor U3462 (N_3462,N_2875,N_2700);
and U3463 (N_3463,N_2731,N_2540);
or U3464 (N_3464,N_2698,N_2379);
or U3465 (N_3465,N_2261,N_2976);
or U3466 (N_3466,N_2526,N_2685);
or U3467 (N_3467,N_2609,N_2147);
nand U3468 (N_3468,N_2926,N_2975);
and U3469 (N_3469,N_2884,N_2255);
nor U3470 (N_3470,N_2449,N_2219);
nor U3471 (N_3471,N_2293,N_2118);
nand U3472 (N_3472,N_2554,N_2729);
and U3473 (N_3473,N_2863,N_2552);
and U3474 (N_3474,N_2722,N_2614);
nand U3475 (N_3475,N_2662,N_2326);
nand U3476 (N_3476,N_2758,N_2690);
and U3477 (N_3477,N_2356,N_2431);
nor U3478 (N_3478,N_2467,N_2461);
or U3479 (N_3479,N_2496,N_2474);
or U3480 (N_3480,N_2972,N_2370);
nand U3481 (N_3481,N_2667,N_2352);
nor U3482 (N_3482,N_2054,N_2081);
nand U3483 (N_3483,N_2783,N_2220);
nand U3484 (N_3484,N_2466,N_2448);
and U3485 (N_3485,N_2881,N_2785);
or U3486 (N_3486,N_2430,N_2096);
or U3487 (N_3487,N_2930,N_2873);
nor U3488 (N_3488,N_2228,N_2278);
and U3489 (N_3489,N_2950,N_2075);
nor U3490 (N_3490,N_2524,N_2121);
nand U3491 (N_3491,N_2342,N_2566);
nor U3492 (N_3492,N_2140,N_2362);
or U3493 (N_3493,N_2537,N_2393);
or U3494 (N_3494,N_2383,N_2399);
and U3495 (N_3495,N_2168,N_2022);
nor U3496 (N_3496,N_2306,N_2176);
nor U3497 (N_3497,N_2070,N_2738);
nand U3498 (N_3498,N_2060,N_2481);
or U3499 (N_3499,N_2279,N_2997);
nor U3500 (N_3500,N_2507,N_2257);
nand U3501 (N_3501,N_2064,N_2142);
or U3502 (N_3502,N_2834,N_2379);
and U3503 (N_3503,N_2579,N_2218);
nand U3504 (N_3504,N_2816,N_2801);
nand U3505 (N_3505,N_2441,N_2616);
nand U3506 (N_3506,N_2031,N_2145);
and U3507 (N_3507,N_2065,N_2054);
nand U3508 (N_3508,N_2797,N_2037);
nand U3509 (N_3509,N_2068,N_2550);
and U3510 (N_3510,N_2858,N_2925);
or U3511 (N_3511,N_2210,N_2626);
nor U3512 (N_3512,N_2738,N_2487);
nor U3513 (N_3513,N_2013,N_2782);
and U3514 (N_3514,N_2593,N_2184);
nor U3515 (N_3515,N_2542,N_2765);
or U3516 (N_3516,N_2556,N_2545);
and U3517 (N_3517,N_2617,N_2175);
nor U3518 (N_3518,N_2157,N_2104);
and U3519 (N_3519,N_2249,N_2832);
and U3520 (N_3520,N_2818,N_2796);
or U3521 (N_3521,N_2799,N_2301);
nor U3522 (N_3522,N_2811,N_2869);
nand U3523 (N_3523,N_2662,N_2978);
or U3524 (N_3524,N_2615,N_2966);
or U3525 (N_3525,N_2631,N_2574);
nand U3526 (N_3526,N_2514,N_2022);
or U3527 (N_3527,N_2115,N_2964);
nor U3528 (N_3528,N_2536,N_2369);
and U3529 (N_3529,N_2448,N_2648);
and U3530 (N_3530,N_2060,N_2631);
nand U3531 (N_3531,N_2630,N_2382);
nor U3532 (N_3532,N_2370,N_2460);
or U3533 (N_3533,N_2444,N_2514);
or U3534 (N_3534,N_2664,N_2149);
nand U3535 (N_3535,N_2757,N_2334);
or U3536 (N_3536,N_2879,N_2492);
or U3537 (N_3537,N_2581,N_2793);
nor U3538 (N_3538,N_2955,N_2379);
or U3539 (N_3539,N_2038,N_2418);
and U3540 (N_3540,N_2115,N_2981);
or U3541 (N_3541,N_2285,N_2613);
or U3542 (N_3542,N_2752,N_2389);
nand U3543 (N_3543,N_2286,N_2341);
and U3544 (N_3544,N_2431,N_2381);
and U3545 (N_3545,N_2377,N_2166);
or U3546 (N_3546,N_2562,N_2418);
nor U3547 (N_3547,N_2899,N_2053);
or U3548 (N_3548,N_2413,N_2142);
and U3549 (N_3549,N_2270,N_2287);
and U3550 (N_3550,N_2636,N_2722);
nor U3551 (N_3551,N_2204,N_2906);
or U3552 (N_3552,N_2492,N_2036);
nor U3553 (N_3553,N_2861,N_2359);
xnor U3554 (N_3554,N_2291,N_2127);
nand U3555 (N_3555,N_2384,N_2699);
nand U3556 (N_3556,N_2772,N_2841);
or U3557 (N_3557,N_2480,N_2137);
or U3558 (N_3558,N_2076,N_2989);
nand U3559 (N_3559,N_2337,N_2507);
and U3560 (N_3560,N_2993,N_2576);
and U3561 (N_3561,N_2723,N_2946);
and U3562 (N_3562,N_2753,N_2258);
or U3563 (N_3563,N_2061,N_2208);
and U3564 (N_3564,N_2508,N_2401);
nor U3565 (N_3565,N_2934,N_2886);
nand U3566 (N_3566,N_2689,N_2692);
nand U3567 (N_3567,N_2443,N_2087);
and U3568 (N_3568,N_2534,N_2004);
and U3569 (N_3569,N_2120,N_2733);
nand U3570 (N_3570,N_2995,N_2846);
xor U3571 (N_3571,N_2548,N_2401);
nor U3572 (N_3572,N_2625,N_2595);
and U3573 (N_3573,N_2386,N_2477);
nor U3574 (N_3574,N_2479,N_2553);
or U3575 (N_3575,N_2181,N_2667);
or U3576 (N_3576,N_2522,N_2396);
and U3577 (N_3577,N_2758,N_2679);
nand U3578 (N_3578,N_2358,N_2670);
nand U3579 (N_3579,N_2338,N_2400);
nand U3580 (N_3580,N_2889,N_2267);
nand U3581 (N_3581,N_2937,N_2412);
and U3582 (N_3582,N_2216,N_2545);
and U3583 (N_3583,N_2811,N_2305);
or U3584 (N_3584,N_2541,N_2494);
nand U3585 (N_3585,N_2486,N_2435);
nand U3586 (N_3586,N_2459,N_2986);
nor U3587 (N_3587,N_2402,N_2028);
nor U3588 (N_3588,N_2049,N_2196);
and U3589 (N_3589,N_2897,N_2700);
or U3590 (N_3590,N_2631,N_2101);
nor U3591 (N_3591,N_2886,N_2805);
or U3592 (N_3592,N_2111,N_2542);
nand U3593 (N_3593,N_2506,N_2027);
and U3594 (N_3594,N_2799,N_2239);
or U3595 (N_3595,N_2576,N_2823);
nand U3596 (N_3596,N_2480,N_2182);
nor U3597 (N_3597,N_2770,N_2901);
nor U3598 (N_3598,N_2467,N_2965);
nand U3599 (N_3599,N_2988,N_2664);
and U3600 (N_3600,N_2687,N_2257);
nand U3601 (N_3601,N_2818,N_2401);
nand U3602 (N_3602,N_2417,N_2086);
or U3603 (N_3603,N_2951,N_2081);
nor U3604 (N_3604,N_2700,N_2997);
and U3605 (N_3605,N_2322,N_2913);
nand U3606 (N_3606,N_2099,N_2446);
and U3607 (N_3607,N_2384,N_2757);
nor U3608 (N_3608,N_2788,N_2864);
nor U3609 (N_3609,N_2690,N_2766);
nor U3610 (N_3610,N_2511,N_2906);
nand U3611 (N_3611,N_2295,N_2979);
or U3612 (N_3612,N_2632,N_2219);
nand U3613 (N_3613,N_2696,N_2434);
or U3614 (N_3614,N_2044,N_2353);
nor U3615 (N_3615,N_2063,N_2561);
nor U3616 (N_3616,N_2108,N_2080);
xor U3617 (N_3617,N_2372,N_2064);
nor U3618 (N_3618,N_2069,N_2994);
or U3619 (N_3619,N_2862,N_2674);
nand U3620 (N_3620,N_2607,N_2669);
and U3621 (N_3621,N_2136,N_2768);
and U3622 (N_3622,N_2291,N_2372);
nor U3623 (N_3623,N_2021,N_2424);
and U3624 (N_3624,N_2266,N_2584);
and U3625 (N_3625,N_2226,N_2689);
and U3626 (N_3626,N_2227,N_2437);
nand U3627 (N_3627,N_2733,N_2663);
or U3628 (N_3628,N_2331,N_2594);
and U3629 (N_3629,N_2444,N_2038);
and U3630 (N_3630,N_2151,N_2288);
and U3631 (N_3631,N_2136,N_2057);
nor U3632 (N_3632,N_2972,N_2708);
or U3633 (N_3633,N_2828,N_2175);
and U3634 (N_3634,N_2193,N_2229);
nor U3635 (N_3635,N_2189,N_2926);
nor U3636 (N_3636,N_2526,N_2141);
nand U3637 (N_3637,N_2247,N_2018);
nor U3638 (N_3638,N_2060,N_2391);
and U3639 (N_3639,N_2397,N_2283);
or U3640 (N_3640,N_2827,N_2325);
or U3641 (N_3641,N_2730,N_2477);
nand U3642 (N_3642,N_2252,N_2423);
and U3643 (N_3643,N_2449,N_2477);
nand U3644 (N_3644,N_2451,N_2717);
nor U3645 (N_3645,N_2997,N_2652);
nor U3646 (N_3646,N_2856,N_2013);
or U3647 (N_3647,N_2924,N_2391);
nand U3648 (N_3648,N_2141,N_2542);
nand U3649 (N_3649,N_2455,N_2368);
and U3650 (N_3650,N_2173,N_2103);
nor U3651 (N_3651,N_2569,N_2386);
or U3652 (N_3652,N_2537,N_2307);
or U3653 (N_3653,N_2646,N_2392);
and U3654 (N_3654,N_2338,N_2108);
xnor U3655 (N_3655,N_2732,N_2587);
or U3656 (N_3656,N_2603,N_2373);
and U3657 (N_3657,N_2729,N_2335);
or U3658 (N_3658,N_2856,N_2347);
and U3659 (N_3659,N_2633,N_2176);
or U3660 (N_3660,N_2331,N_2387);
nand U3661 (N_3661,N_2260,N_2097);
nand U3662 (N_3662,N_2391,N_2913);
and U3663 (N_3663,N_2155,N_2908);
and U3664 (N_3664,N_2899,N_2101);
nor U3665 (N_3665,N_2995,N_2835);
nand U3666 (N_3666,N_2872,N_2452);
and U3667 (N_3667,N_2978,N_2257);
and U3668 (N_3668,N_2844,N_2703);
or U3669 (N_3669,N_2219,N_2759);
and U3670 (N_3670,N_2719,N_2009);
nor U3671 (N_3671,N_2608,N_2400);
nand U3672 (N_3672,N_2705,N_2258);
nand U3673 (N_3673,N_2552,N_2403);
and U3674 (N_3674,N_2175,N_2433);
and U3675 (N_3675,N_2777,N_2628);
nor U3676 (N_3676,N_2890,N_2976);
and U3677 (N_3677,N_2274,N_2629);
nor U3678 (N_3678,N_2072,N_2976);
and U3679 (N_3679,N_2946,N_2292);
nor U3680 (N_3680,N_2559,N_2428);
nand U3681 (N_3681,N_2301,N_2607);
nand U3682 (N_3682,N_2349,N_2635);
nor U3683 (N_3683,N_2314,N_2686);
nor U3684 (N_3684,N_2681,N_2513);
or U3685 (N_3685,N_2184,N_2316);
nor U3686 (N_3686,N_2476,N_2694);
or U3687 (N_3687,N_2085,N_2783);
and U3688 (N_3688,N_2245,N_2183);
nand U3689 (N_3689,N_2432,N_2960);
nand U3690 (N_3690,N_2396,N_2428);
or U3691 (N_3691,N_2945,N_2261);
and U3692 (N_3692,N_2006,N_2174);
and U3693 (N_3693,N_2196,N_2197);
xor U3694 (N_3694,N_2715,N_2518);
nor U3695 (N_3695,N_2109,N_2120);
and U3696 (N_3696,N_2080,N_2369);
or U3697 (N_3697,N_2402,N_2879);
or U3698 (N_3698,N_2940,N_2286);
or U3699 (N_3699,N_2215,N_2936);
or U3700 (N_3700,N_2695,N_2920);
and U3701 (N_3701,N_2154,N_2374);
and U3702 (N_3702,N_2155,N_2516);
nand U3703 (N_3703,N_2151,N_2835);
nand U3704 (N_3704,N_2988,N_2653);
nand U3705 (N_3705,N_2781,N_2423);
nand U3706 (N_3706,N_2612,N_2939);
and U3707 (N_3707,N_2759,N_2606);
nor U3708 (N_3708,N_2200,N_2166);
nand U3709 (N_3709,N_2325,N_2731);
nor U3710 (N_3710,N_2195,N_2826);
or U3711 (N_3711,N_2378,N_2950);
and U3712 (N_3712,N_2058,N_2396);
or U3713 (N_3713,N_2801,N_2674);
nand U3714 (N_3714,N_2698,N_2389);
or U3715 (N_3715,N_2441,N_2422);
nand U3716 (N_3716,N_2847,N_2284);
or U3717 (N_3717,N_2204,N_2015);
xor U3718 (N_3718,N_2354,N_2954);
and U3719 (N_3719,N_2925,N_2391);
and U3720 (N_3720,N_2285,N_2009);
or U3721 (N_3721,N_2543,N_2756);
and U3722 (N_3722,N_2507,N_2549);
and U3723 (N_3723,N_2611,N_2017);
and U3724 (N_3724,N_2816,N_2776);
nor U3725 (N_3725,N_2822,N_2578);
nand U3726 (N_3726,N_2725,N_2549);
and U3727 (N_3727,N_2732,N_2083);
nand U3728 (N_3728,N_2104,N_2079);
nand U3729 (N_3729,N_2030,N_2059);
nor U3730 (N_3730,N_2433,N_2651);
or U3731 (N_3731,N_2039,N_2730);
nor U3732 (N_3732,N_2944,N_2949);
or U3733 (N_3733,N_2417,N_2555);
nand U3734 (N_3734,N_2636,N_2509);
nand U3735 (N_3735,N_2493,N_2820);
or U3736 (N_3736,N_2540,N_2845);
and U3737 (N_3737,N_2836,N_2546);
nor U3738 (N_3738,N_2968,N_2901);
and U3739 (N_3739,N_2967,N_2936);
nand U3740 (N_3740,N_2927,N_2973);
nor U3741 (N_3741,N_2340,N_2283);
or U3742 (N_3742,N_2557,N_2913);
nor U3743 (N_3743,N_2309,N_2319);
and U3744 (N_3744,N_2758,N_2484);
nand U3745 (N_3745,N_2892,N_2403);
xor U3746 (N_3746,N_2626,N_2984);
and U3747 (N_3747,N_2120,N_2845);
and U3748 (N_3748,N_2062,N_2894);
or U3749 (N_3749,N_2826,N_2228);
nand U3750 (N_3750,N_2776,N_2131);
nor U3751 (N_3751,N_2048,N_2886);
and U3752 (N_3752,N_2111,N_2108);
nor U3753 (N_3753,N_2932,N_2020);
or U3754 (N_3754,N_2093,N_2255);
nand U3755 (N_3755,N_2054,N_2770);
or U3756 (N_3756,N_2564,N_2674);
nand U3757 (N_3757,N_2570,N_2591);
nand U3758 (N_3758,N_2080,N_2649);
or U3759 (N_3759,N_2312,N_2155);
and U3760 (N_3760,N_2173,N_2653);
or U3761 (N_3761,N_2859,N_2839);
and U3762 (N_3762,N_2792,N_2647);
and U3763 (N_3763,N_2083,N_2213);
or U3764 (N_3764,N_2562,N_2383);
nand U3765 (N_3765,N_2393,N_2368);
nor U3766 (N_3766,N_2060,N_2814);
nand U3767 (N_3767,N_2093,N_2376);
nor U3768 (N_3768,N_2309,N_2934);
nor U3769 (N_3769,N_2246,N_2399);
or U3770 (N_3770,N_2062,N_2989);
nand U3771 (N_3771,N_2653,N_2480);
or U3772 (N_3772,N_2827,N_2088);
nor U3773 (N_3773,N_2584,N_2930);
and U3774 (N_3774,N_2071,N_2230);
and U3775 (N_3775,N_2484,N_2445);
and U3776 (N_3776,N_2025,N_2675);
or U3777 (N_3777,N_2334,N_2264);
or U3778 (N_3778,N_2356,N_2337);
nor U3779 (N_3779,N_2466,N_2810);
or U3780 (N_3780,N_2117,N_2649);
and U3781 (N_3781,N_2260,N_2479);
and U3782 (N_3782,N_2568,N_2730);
nand U3783 (N_3783,N_2445,N_2521);
or U3784 (N_3784,N_2123,N_2499);
nor U3785 (N_3785,N_2097,N_2686);
nor U3786 (N_3786,N_2482,N_2358);
or U3787 (N_3787,N_2137,N_2154);
or U3788 (N_3788,N_2746,N_2658);
nand U3789 (N_3789,N_2107,N_2054);
nand U3790 (N_3790,N_2485,N_2550);
nand U3791 (N_3791,N_2106,N_2353);
nor U3792 (N_3792,N_2707,N_2144);
and U3793 (N_3793,N_2965,N_2967);
or U3794 (N_3794,N_2564,N_2608);
nand U3795 (N_3795,N_2623,N_2058);
nand U3796 (N_3796,N_2867,N_2805);
or U3797 (N_3797,N_2137,N_2558);
or U3798 (N_3798,N_2356,N_2406);
nor U3799 (N_3799,N_2230,N_2733);
and U3800 (N_3800,N_2953,N_2623);
nor U3801 (N_3801,N_2792,N_2197);
nor U3802 (N_3802,N_2070,N_2890);
nand U3803 (N_3803,N_2728,N_2813);
nor U3804 (N_3804,N_2054,N_2705);
nand U3805 (N_3805,N_2634,N_2171);
nor U3806 (N_3806,N_2392,N_2543);
or U3807 (N_3807,N_2178,N_2849);
nand U3808 (N_3808,N_2930,N_2469);
and U3809 (N_3809,N_2034,N_2194);
and U3810 (N_3810,N_2819,N_2101);
or U3811 (N_3811,N_2463,N_2102);
or U3812 (N_3812,N_2878,N_2066);
nand U3813 (N_3813,N_2091,N_2935);
nand U3814 (N_3814,N_2698,N_2496);
nand U3815 (N_3815,N_2256,N_2723);
or U3816 (N_3816,N_2763,N_2743);
and U3817 (N_3817,N_2381,N_2027);
or U3818 (N_3818,N_2633,N_2600);
and U3819 (N_3819,N_2957,N_2333);
nand U3820 (N_3820,N_2720,N_2328);
or U3821 (N_3821,N_2631,N_2859);
and U3822 (N_3822,N_2992,N_2492);
and U3823 (N_3823,N_2156,N_2898);
nor U3824 (N_3824,N_2236,N_2451);
nor U3825 (N_3825,N_2311,N_2580);
nor U3826 (N_3826,N_2644,N_2936);
and U3827 (N_3827,N_2556,N_2108);
nand U3828 (N_3828,N_2818,N_2105);
nor U3829 (N_3829,N_2301,N_2858);
nor U3830 (N_3830,N_2843,N_2087);
nor U3831 (N_3831,N_2325,N_2386);
and U3832 (N_3832,N_2694,N_2744);
nor U3833 (N_3833,N_2349,N_2754);
nor U3834 (N_3834,N_2684,N_2895);
or U3835 (N_3835,N_2641,N_2721);
or U3836 (N_3836,N_2004,N_2924);
or U3837 (N_3837,N_2707,N_2019);
nand U3838 (N_3838,N_2036,N_2234);
nor U3839 (N_3839,N_2217,N_2812);
and U3840 (N_3840,N_2283,N_2595);
nand U3841 (N_3841,N_2775,N_2716);
and U3842 (N_3842,N_2831,N_2263);
and U3843 (N_3843,N_2979,N_2966);
nand U3844 (N_3844,N_2681,N_2096);
nor U3845 (N_3845,N_2901,N_2661);
or U3846 (N_3846,N_2007,N_2912);
nand U3847 (N_3847,N_2214,N_2749);
nand U3848 (N_3848,N_2748,N_2695);
nor U3849 (N_3849,N_2814,N_2717);
and U3850 (N_3850,N_2040,N_2685);
nand U3851 (N_3851,N_2826,N_2861);
or U3852 (N_3852,N_2356,N_2229);
nor U3853 (N_3853,N_2210,N_2257);
nand U3854 (N_3854,N_2733,N_2482);
or U3855 (N_3855,N_2414,N_2666);
and U3856 (N_3856,N_2912,N_2907);
nand U3857 (N_3857,N_2029,N_2165);
or U3858 (N_3858,N_2101,N_2447);
or U3859 (N_3859,N_2005,N_2427);
nor U3860 (N_3860,N_2181,N_2847);
and U3861 (N_3861,N_2221,N_2439);
nor U3862 (N_3862,N_2484,N_2045);
or U3863 (N_3863,N_2855,N_2538);
nor U3864 (N_3864,N_2999,N_2129);
nand U3865 (N_3865,N_2348,N_2932);
nor U3866 (N_3866,N_2685,N_2940);
nand U3867 (N_3867,N_2714,N_2124);
and U3868 (N_3868,N_2962,N_2498);
and U3869 (N_3869,N_2338,N_2614);
or U3870 (N_3870,N_2572,N_2271);
and U3871 (N_3871,N_2530,N_2940);
and U3872 (N_3872,N_2498,N_2041);
nand U3873 (N_3873,N_2300,N_2241);
nor U3874 (N_3874,N_2540,N_2473);
and U3875 (N_3875,N_2963,N_2324);
and U3876 (N_3876,N_2120,N_2242);
or U3877 (N_3877,N_2883,N_2714);
nor U3878 (N_3878,N_2682,N_2725);
nor U3879 (N_3879,N_2370,N_2396);
nor U3880 (N_3880,N_2392,N_2528);
nor U3881 (N_3881,N_2347,N_2926);
nor U3882 (N_3882,N_2972,N_2081);
nor U3883 (N_3883,N_2249,N_2883);
nand U3884 (N_3884,N_2960,N_2090);
nand U3885 (N_3885,N_2858,N_2979);
and U3886 (N_3886,N_2033,N_2639);
nand U3887 (N_3887,N_2418,N_2034);
nand U3888 (N_3888,N_2787,N_2735);
and U3889 (N_3889,N_2915,N_2094);
nand U3890 (N_3890,N_2011,N_2599);
or U3891 (N_3891,N_2252,N_2853);
or U3892 (N_3892,N_2652,N_2550);
and U3893 (N_3893,N_2721,N_2522);
or U3894 (N_3894,N_2882,N_2016);
or U3895 (N_3895,N_2337,N_2414);
nor U3896 (N_3896,N_2053,N_2960);
nor U3897 (N_3897,N_2034,N_2065);
nand U3898 (N_3898,N_2016,N_2712);
nand U3899 (N_3899,N_2199,N_2277);
nand U3900 (N_3900,N_2192,N_2710);
or U3901 (N_3901,N_2976,N_2236);
or U3902 (N_3902,N_2896,N_2849);
and U3903 (N_3903,N_2737,N_2281);
nand U3904 (N_3904,N_2992,N_2010);
and U3905 (N_3905,N_2756,N_2675);
nor U3906 (N_3906,N_2889,N_2860);
or U3907 (N_3907,N_2421,N_2916);
nand U3908 (N_3908,N_2338,N_2873);
and U3909 (N_3909,N_2422,N_2514);
or U3910 (N_3910,N_2151,N_2275);
and U3911 (N_3911,N_2812,N_2561);
nand U3912 (N_3912,N_2306,N_2542);
nor U3913 (N_3913,N_2351,N_2155);
xnor U3914 (N_3914,N_2854,N_2233);
and U3915 (N_3915,N_2546,N_2995);
and U3916 (N_3916,N_2705,N_2029);
and U3917 (N_3917,N_2301,N_2358);
nand U3918 (N_3918,N_2859,N_2971);
nor U3919 (N_3919,N_2153,N_2168);
or U3920 (N_3920,N_2705,N_2042);
nand U3921 (N_3921,N_2572,N_2609);
or U3922 (N_3922,N_2192,N_2458);
and U3923 (N_3923,N_2782,N_2435);
nor U3924 (N_3924,N_2404,N_2790);
nor U3925 (N_3925,N_2861,N_2705);
nand U3926 (N_3926,N_2183,N_2641);
nand U3927 (N_3927,N_2950,N_2983);
or U3928 (N_3928,N_2791,N_2536);
nor U3929 (N_3929,N_2682,N_2460);
and U3930 (N_3930,N_2755,N_2054);
and U3931 (N_3931,N_2989,N_2866);
nor U3932 (N_3932,N_2092,N_2017);
nor U3933 (N_3933,N_2894,N_2337);
and U3934 (N_3934,N_2015,N_2442);
nor U3935 (N_3935,N_2307,N_2882);
nand U3936 (N_3936,N_2199,N_2377);
nor U3937 (N_3937,N_2337,N_2442);
nand U3938 (N_3938,N_2633,N_2303);
nor U3939 (N_3939,N_2873,N_2989);
or U3940 (N_3940,N_2968,N_2846);
nand U3941 (N_3941,N_2652,N_2804);
nand U3942 (N_3942,N_2982,N_2320);
and U3943 (N_3943,N_2488,N_2261);
or U3944 (N_3944,N_2418,N_2962);
nor U3945 (N_3945,N_2718,N_2192);
nor U3946 (N_3946,N_2504,N_2902);
nor U3947 (N_3947,N_2971,N_2786);
nor U3948 (N_3948,N_2199,N_2585);
nor U3949 (N_3949,N_2658,N_2897);
and U3950 (N_3950,N_2800,N_2544);
nand U3951 (N_3951,N_2033,N_2984);
nor U3952 (N_3952,N_2266,N_2158);
and U3953 (N_3953,N_2029,N_2709);
nand U3954 (N_3954,N_2321,N_2481);
and U3955 (N_3955,N_2011,N_2857);
nor U3956 (N_3956,N_2354,N_2345);
and U3957 (N_3957,N_2670,N_2132);
nor U3958 (N_3958,N_2603,N_2702);
and U3959 (N_3959,N_2995,N_2764);
nor U3960 (N_3960,N_2049,N_2654);
nand U3961 (N_3961,N_2611,N_2825);
and U3962 (N_3962,N_2790,N_2206);
nand U3963 (N_3963,N_2711,N_2447);
or U3964 (N_3964,N_2389,N_2098);
and U3965 (N_3965,N_2160,N_2481);
and U3966 (N_3966,N_2254,N_2315);
and U3967 (N_3967,N_2042,N_2771);
nand U3968 (N_3968,N_2733,N_2112);
or U3969 (N_3969,N_2697,N_2091);
or U3970 (N_3970,N_2276,N_2928);
or U3971 (N_3971,N_2606,N_2343);
nand U3972 (N_3972,N_2652,N_2200);
or U3973 (N_3973,N_2007,N_2001);
and U3974 (N_3974,N_2763,N_2685);
or U3975 (N_3975,N_2933,N_2168);
nor U3976 (N_3976,N_2106,N_2494);
or U3977 (N_3977,N_2828,N_2587);
or U3978 (N_3978,N_2433,N_2598);
nor U3979 (N_3979,N_2631,N_2976);
nor U3980 (N_3980,N_2384,N_2394);
or U3981 (N_3981,N_2764,N_2915);
nand U3982 (N_3982,N_2498,N_2261);
nor U3983 (N_3983,N_2480,N_2943);
nor U3984 (N_3984,N_2746,N_2009);
and U3985 (N_3985,N_2375,N_2144);
nand U3986 (N_3986,N_2619,N_2729);
nand U3987 (N_3987,N_2977,N_2711);
nand U3988 (N_3988,N_2183,N_2405);
nand U3989 (N_3989,N_2534,N_2424);
nor U3990 (N_3990,N_2858,N_2273);
nand U3991 (N_3991,N_2499,N_2801);
nor U3992 (N_3992,N_2548,N_2462);
or U3993 (N_3993,N_2634,N_2467);
and U3994 (N_3994,N_2655,N_2819);
or U3995 (N_3995,N_2640,N_2145);
nor U3996 (N_3996,N_2017,N_2123);
and U3997 (N_3997,N_2910,N_2509);
or U3998 (N_3998,N_2769,N_2961);
nand U3999 (N_3999,N_2540,N_2718);
nor U4000 (N_4000,N_3637,N_3880);
nor U4001 (N_4001,N_3118,N_3583);
nand U4002 (N_4002,N_3343,N_3531);
and U4003 (N_4003,N_3937,N_3138);
or U4004 (N_4004,N_3823,N_3845);
and U4005 (N_4005,N_3542,N_3368);
xor U4006 (N_4006,N_3490,N_3738);
nand U4007 (N_4007,N_3928,N_3509);
and U4008 (N_4008,N_3636,N_3361);
and U4009 (N_4009,N_3161,N_3305);
or U4010 (N_4010,N_3570,N_3471);
nand U4011 (N_4011,N_3914,N_3489);
nor U4012 (N_4012,N_3781,N_3815);
or U4013 (N_4013,N_3959,N_3847);
or U4014 (N_4014,N_3609,N_3960);
or U4015 (N_4015,N_3818,N_3034);
or U4016 (N_4016,N_3836,N_3094);
and U4017 (N_4017,N_3271,N_3200);
nor U4018 (N_4018,N_3719,N_3619);
and U4019 (N_4019,N_3463,N_3771);
and U4020 (N_4020,N_3042,N_3301);
or U4021 (N_4021,N_3546,N_3026);
and U4022 (N_4022,N_3057,N_3088);
and U4023 (N_4023,N_3076,N_3616);
or U4024 (N_4024,N_3576,N_3601);
and U4025 (N_4025,N_3188,N_3434);
and U4026 (N_4026,N_3505,N_3851);
or U4027 (N_4027,N_3220,N_3497);
nand U4028 (N_4028,N_3116,N_3491);
or U4029 (N_4029,N_3268,N_3354);
nand U4030 (N_4030,N_3260,N_3371);
nand U4031 (N_4031,N_3930,N_3902);
nand U4032 (N_4032,N_3174,N_3833);
or U4033 (N_4033,N_3310,N_3538);
and U4034 (N_4034,N_3723,N_3429);
and U4035 (N_4035,N_3108,N_3910);
nor U4036 (N_4036,N_3496,N_3228);
nor U4037 (N_4037,N_3341,N_3025);
and U4038 (N_4038,N_3993,N_3473);
nor U4039 (N_4039,N_3573,N_3911);
and U4040 (N_4040,N_3657,N_3886);
nand U4041 (N_4041,N_3877,N_3926);
or U4042 (N_4042,N_3043,N_3058);
xnor U4043 (N_4043,N_3452,N_3824);
nor U4044 (N_4044,N_3762,N_3387);
and U4045 (N_4045,N_3949,N_3905);
and U4046 (N_4046,N_3101,N_3339);
and U4047 (N_4047,N_3769,N_3376);
or U4048 (N_4048,N_3250,N_3385);
and U4049 (N_4049,N_3751,N_3224);
or U4050 (N_4050,N_3875,N_3501);
nor U4051 (N_4051,N_3523,N_3077);
or U4052 (N_4052,N_3715,N_3780);
nor U4053 (N_4053,N_3622,N_3592);
or U4054 (N_4054,N_3205,N_3537);
nand U4055 (N_4055,N_3165,N_3030);
and U4056 (N_4056,N_3774,N_3962);
nand U4057 (N_4057,N_3667,N_3915);
nor U4058 (N_4058,N_3721,N_3210);
nor U4059 (N_4059,N_3010,N_3096);
nor U4060 (N_4060,N_3488,N_3425);
nor U4061 (N_4061,N_3122,N_3628);
nand U4062 (N_4062,N_3690,N_3579);
and U4063 (N_4063,N_3702,N_3175);
nor U4064 (N_4064,N_3014,N_3194);
nor U4065 (N_4065,N_3066,N_3532);
or U4066 (N_4066,N_3044,N_3166);
nand U4067 (N_4067,N_3016,N_3292);
nor U4068 (N_4068,N_3209,N_3445);
or U4069 (N_4069,N_3347,N_3067);
or U4070 (N_4070,N_3262,N_3747);
nand U4071 (N_4071,N_3394,N_3896);
nor U4072 (N_4072,N_3689,N_3775);
nor U4073 (N_4073,N_3396,N_3989);
or U4074 (N_4074,N_3104,N_3925);
nand U4075 (N_4075,N_3516,N_3481);
nor U4076 (N_4076,N_3085,N_3696);
nor U4077 (N_4077,N_3363,N_3897);
and U4078 (N_4078,N_3778,N_3627);
nand U4079 (N_4079,N_3403,N_3678);
and U4080 (N_4080,N_3587,N_3199);
and U4081 (N_4081,N_3257,N_3229);
nand U4082 (N_4082,N_3817,N_3267);
or U4083 (N_4083,N_3097,N_3519);
and U4084 (N_4084,N_3961,N_3699);
nor U4085 (N_4085,N_3284,N_3470);
nand U4086 (N_4086,N_3838,N_3536);
nand U4087 (N_4087,N_3631,N_3350);
nor U4088 (N_4088,N_3040,N_3236);
nand U4089 (N_4089,N_3302,N_3029);
or U4090 (N_4090,N_3648,N_3211);
or U4091 (N_4091,N_3712,N_3948);
nor U4092 (N_4092,N_3317,N_3547);
or U4093 (N_4093,N_3173,N_3287);
nand U4094 (N_4094,N_3869,N_3770);
nor U4095 (N_4095,N_3759,N_3072);
or U4096 (N_4096,N_3863,N_3594);
nor U4097 (N_4097,N_3180,N_3308);
nor U4098 (N_4098,N_3968,N_3632);
nor U4099 (N_4099,N_3714,N_3840);
nor U4100 (N_4100,N_3599,N_3704);
nor U4101 (N_4101,N_3453,N_3127);
or U4102 (N_4102,N_3917,N_3716);
nand U4103 (N_4103,N_3359,N_3617);
nand U4104 (N_4104,N_3272,N_3410);
or U4105 (N_4105,N_3419,N_3381);
nor U4106 (N_4106,N_3316,N_3144);
nor U4107 (N_4107,N_3682,N_3395);
or U4108 (N_4108,N_3612,N_3325);
and U4109 (N_4109,N_3136,N_3084);
or U4110 (N_4110,N_3100,N_3558);
or U4111 (N_4111,N_3859,N_3055);
and U4112 (N_4112,N_3729,N_3764);
and U4113 (N_4113,N_3052,N_3462);
nor U4114 (N_4114,N_3391,N_3977);
nand U4115 (N_4115,N_3692,N_3335);
nor U4116 (N_4116,N_3294,N_3171);
and U4117 (N_4117,N_3665,N_3786);
or U4118 (N_4118,N_3157,N_3743);
nor U4119 (N_4119,N_3620,N_3373);
and U4120 (N_4120,N_3214,N_3023);
and U4121 (N_4121,N_3821,N_3276);
or U4122 (N_4122,N_3768,N_3345);
and U4123 (N_4123,N_3513,N_3584);
and U4124 (N_4124,N_3980,N_3849);
nor U4125 (N_4125,N_3602,N_3883);
or U4126 (N_4126,N_3295,N_3389);
nor U4127 (N_4127,N_3881,N_3867);
nor U4128 (N_4128,N_3447,N_3801);
nand U4129 (N_4129,N_3564,N_3603);
and U4130 (N_4130,N_3830,N_3724);
or U4131 (N_4131,N_3132,N_3553);
and U4132 (N_4132,N_3595,N_3870);
or U4133 (N_4133,N_3380,N_3983);
nand U4134 (N_4134,N_3423,N_3472);
nor U4135 (N_4135,N_3237,N_3701);
or U4136 (N_4136,N_3435,N_3195);
nor U4137 (N_4137,N_3009,N_3650);
nor U4138 (N_4138,N_3231,N_3258);
or U4139 (N_4139,N_3324,N_3777);
or U4140 (N_4140,N_3129,N_3071);
nor U4141 (N_4141,N_3252,N_3124);
and U4142 (N_4142,N_3069,N_3145);
nor U4143 (N_4143,N_3213,N_3502);
nor U4144 (N_4144,N_3179,N_3464);
or U4145 (N_4145,N_3854,N_3659);
nand U4146 (N_4146,N_3107,N_3326);
or U4147 (N_4147,N_3728,N_3251);
and U4148 (N_4148,N_3369,N_3556);
and U4149 (N_4149,N_3186,N_3827);
or U4150 (N_4150,N_3559,N_3647);
nor U4151 (N_4151,N_3498,N_3311);
or U4152 (N_4152,N_3282,N_3053);
nand U4153 (N_4153,N_3624,N_3934);
or U4154 (N_4154,N_3374,N_3586);
or U4155 (N_4155,N_3427,N_3901);
or U4156 (N_4156,N_3154,N_3791);
nor U4157 (N_4157,N_3451,N_3545);
and U4158 (N_4158,N_3718,N_3608);
or U4159 (N_4159,N_3405,N_3795);
xnor U4160 (N_4160,N_3691,N_3318);
and U4161 (N_4161,N_3408,N_3543);
nor U4162 (N_4162,N_3921,N_3709);
nand U4163 (N_4163,N_3889,N_3710);
or U4164 (N_4164,N_3215,N_3755);
or U4165 (N_4165,N_3190,N_3511);
nand U4166 (N_4166,N_3806,N_3858);
nor U4167 (N_4167,N_3874,N_3286);
and U4168 (N_4168,N_3758,N_3614);
nor U4169 (N_4169,N_3019,N_3035);
or U4170 (N_4170,N_3856,N_3500);
nor U4171 (N_4171,N_3388,N_3593);
and U4172 (N_4172,N_3951,N_3015);
xor U4173 (N_4173,N_3688,N_3540);
nand U4174 (N_4174,N_3499,N_3244);
nand U4175 (N_4175,N_3207,N_3800);
or U4176 (N_4176,N_3033,N_3274);
or U4177 (N_4177,N_3431,N_3909);
and U4178 (N_4178,N_3455,N_3525);
and U4179 (N_4179,N_3613,N_3012);
and U4180 (N_4180,N_3242,N_3984);
nor U4181 (N_4181,N_3280,N_3739);
or U4182 (N_4182,N_3591,N_3046);
and U4183 (N_4183,N_3837,N_3168);
nor U4184 (N_4184,N_3259,N_3932);
nand U4185 (N_4185,N_3152,N_3086);
nor U4186 (N_4186,N_3985,N_3080);
nor U4187 (N_4187,N_3634,N_3328);
nor U4188 (N_4188,N_3146,N_3254);
nor U4189 (N_4189,N_3810,N_3045);
nand U4190 (N_4190,N_3417,N_3649);
nand U4191 (N_4191,N_3933,N_3130);
or U4192 (N_4192,N_3176,N_3398);
nor U4193 (N_4193,N_3296,N_3298);
or U4194 (N_4194,N_3117,N_3623);
nor U4195 (N_4195,N_3020,N_3275);
nor U4196 (N_4196,N_3248,N_3039);
and U4197 (N_4197,N_3799,N_3589);
or U4198 (N_4198,N_3652,N_3796);
or U4199 (N_4199,N_3742,N_3448);
nor U4200 (N_4200,N_3309,N_3585);
or U4201 (N_4201,N_3633,N_3013);
or U4202 (N_4202,N_3203,N_3736);
nand U4203 (N_4203,N_3572,N_3312);
and U4204 (N_4204,N_3606,N_3588);
nand U4205 (N_4205,N_3748,N_3997);
or U4206 (N_4206,N_3114,N_3457);
or U4207 (N_4207,N_3115,N_3342);
nor U4208 (N_4208,N_3041,N_3565);
or U4209 (N_4209,N_3264,N_3575);
and U4210 (N_4210,N_3008,N_3773);
or U4211 (N_4211,N_3574,N_3642);
or U4212 (N_4212,N_3185,N_3333);
nand U4213 (N_4213,N_3518,N_3646);
and U4214 (N_4214,N_3021,N_3459);
and U4215 (N_4215,N_3611,N_3697);
or U4216 (N_4216,N_3234,N_3153);
and U4217 (N_4217,N_3323,N_3803);
nand U4218 (N_4218,N_3994,N_3437);
nand U4219 (N_4219,N_3375,N_3393);
nor U4220 (N_4220,N_3163,N_3842);
nor U4221 (N_4221,N_3814,N_3879);
and U4222 (N_4222,N_3358,N_3050);
nor U4223 (N_4223,N_3285,N_3444);
and U4224 (N_4224,N_3861,N_3202);
nor U4225 (N_4225,N_3112,N_3119);
nand U4226 (N_4226,N_3607,N_3390);
nor U4227 (N_4227,N_3037,N_3899);
and U4228 (N_4228,N_3635,N_3562);
nand U4229 (N_4229,N_3032,N_3197);
xnor U4230 (N_4230,N_3300,N_3142);
and U4231 (N_4231,N_3973,N_3544);
and U4232 (N_4232,N_3283,N_3629);
and U4233 (N_4233,N_3279,N_3420);
or U4234 (N_4234,N_3507,N_3018);
or U4235 (N_4235,N_3740,N_3675);
nor U4236 (N_4236,N_3281,N_3133);
nand U4237 (N_4237,N_3788,N_3663);
nand U4238 (N_4238,N_3766,N_3478);
and U4239 (N_4239,N_3508,N_3192);
and U4240 (N_4240,N_3946,N_3201);
or U4241 (N_4241,N_3965,N_3098);
nor U4242 (N_4242,N_3327,N_3123);
nand U4243 (N_4243,N_3936,N_3204);
or U4244 (N_4244,N_3454,N_3772);
nor U4245 (N_4245,N_3426,N_3226);
nand U4246 (N_4246,N_3089,N_3844);
and U4247 (N_4247,N_3289,N_3139);
or U4248 (N_4248,N_3348,N_3539);
nor U4249 (N_4249,N_3535,N_3843);
nor U4250 (N_4250,N_3137,N_3477);
nor U4251 (N_4251,N_3126,N_3450);
nand U4252 (N_4252,N_3517,N_3666);
nand U4253 (N_4253,N_3456,N_3352);
nor U4254 (N_4254,N_3480,N_3460);
nand U4255 (N_4255,N_3293,N_3940);
nand U4256 (N_4256,N_3950,N_3876);
nand U4257 (N_4257,N_3693,N_3338);
nor U4258 (N_4258,N_3908,N_3804);
nand U4259 (N_4259,N_3277,N_3007);
nand U4260 (N_4260,N_3991,N_3256);
nand U4261 (N_4261,N_3597,N_3064);
nand U4262 (N_4262,N_3253,N_3418);
nor U4263 (N_4263,N_3038,N_3669);
nor U4264 (N_4264,N_3906,N_3964);
nand U4265 (N_4265,N_3563,N_3241);
and U4266 (N_4266,N_3193,N_3075);
or U4267 (N_4267,N_3436,N_3664);
or U4268 (N_4268,N_3492,N_3852);
and U4269 (N_4269,N_3087,N_3346);
or U4270 (N_4270,N_3430,N_3763);
and U4271 (N_4271,N_3812,N_3494);
nand U4272 (N_4272,N_3534,N_3217);
and U4273 (N_4273,N_3982,N_3105);
nand U4274 (N_4274,N_3571,N_3885);
nor U4275 (N_4275,N_3732,N_3320);
nand U4276 (N_4276,N_3734,N_3110);
and U4277 (N_4277,N_3578,N_3245);
nor U4278 (N_4278,N_3722,N_3401);
nand U4279 (N_4279,N_3760,N_3467);
and U4280 (N_4280,N_3641,N_3998);
or U4281 (N_4281,N_3036,N_3073);
nand U4282 (N_4282,N_3337,N_3522);
nand U4283 (N_4283,N_3953,N_3947);
nand U4284 (N_4284,N_3265,N_3249);
nand U4285 (N_4285,N_3683,N_3125);
or U4286 (N_4286,N_3752,N_3240);
xor U4287 (N_4287,N_3626,N_3465);
or U4288 (N_4288,N_3733,N_3860);
nand U4289 (N_4289,N_3735,N_3416);
nor U4290 (N_4290,N_3924,N_3695);
nor U4291 (N_4291,N_3191,N_3196);
nor U4292 (N_4292,N_3676,N_3938);
and U4293 (N_4293,N_3708,N_3750);
nand U4294 (N_4294,N_3159,N_3412);
or U4295 (N_4295,N_3894,N_3783);
nor U4296 (N_4296,N_3744,N_3898);
or U4297 (N_4297,N_3336,N_3206);
or U4298 (N_4298,N_3767,N_3261);
nor U4299 (N_4299,N_3307,N_3485);
and U4300 (N_4300,N_3530,N_3364);
nor U4301 (N_4301,N_3484,N_3099);
xnor U4302 (N_4302,N_3379,N_3230);
nand U4303 (N_4303,N_3003,N_3313);
nand U4304 (N_4304,N_3344,N_3990);
and U4305 (N_4305,N_3872,N_3081);
or U4306 (N_4306,N_3263,N_3919);
or U4307 (N_4307,N_3551,N_3967);
nor U4308 (N_4308,N_3978,N_3474);
or U4309 (N_4309,N_3935,N_3510);
and U4310 (N_4310,N_3141,N_3068);
nand U4311 (N_4311,N_3255,N_3172);
nand U4312 (N_4312,N_3785,N_3221);
nand U4313 (N_4313,N_3944,N_3103);
and U4314 (N_4314,N_3560,N_3140);
or U4315 (N_4315,N_3605,N_3864);
nor U4316 (N_4316,N_3054,N_3314);
nor U4317 (N_4317,N_3923,N_3566);
nand U4318 (N_4318,N_3349,N_3550);
and U4319 (N_4319,N_3903,N_3671);
or U4320 (N_4320,N_3147,N_3273);
nor U4321 (N_4321,N_3807,N_3218);
nor U4322 (N_4322,N_3422,N_3793);
nand U4323 (N_4323,N_3731,N_3841);
nor U4324 (N_4324,N_3332,N_3670);
nand U4325 (N_4325,N_3329,N_3970);
nor U4326 (N_4326,N_3061,N_3406);
and U4327 (N_4327,N_3432,N_3362);
nand U4328 (N_4328,N_3177,N_3868);
or U4329 (N_4329,N_3981,N_3850);
nor U4330 (N_4330,N_3839,N_3331);
or U4331 (N_4331,N_3674,N_3643);
nor U4332 (N_4332,N_3878,N_3005);
and U4333 (N_4333,N_3918,N_3972);
or U4334 (N_4334,N_3668,N_3561);
nor U4335 (N_4335,N_3567,N_3825);
and U4336 (N_4336,N_3737,N_3568);
or U4337 (N_4337,N_3533,N_3384);
or U4338 (N_4338,N_3999,N_3645);
or U4339 (N_4339,N_3904,N_3183);
and U4340 (N_4340,N_3835,N_3805);
nand U4341 (N_4341,N_3527,N_3216);
or U4342 (N_4342,N_3006,N_3581);
nor U4343 (N_4343,N_3580,N_3548);
or U4344 (N_4344,N_3654,N_3826);
and U4345 (N_4345,N_3979,N_3920);
nand U4346 (N_4346,N_3392,N_3618);
nor U4347 (N_4347,N_3212,N_3976);
nand U4348 (N_4348,N_3662,N_3091);
nor U4349 (N_4349,N_3169,N_3707);
nor U4350 (N_4350,N_3776,N_3787);
and U4351 (N_4351,N_3297,N_3658);
nand U4352 (N_4352,N_3079,N_3644);
nand U4353 (N_4353,N_3988,N_3577);
and U4354 (N_4354,N_3278,N_3414);
or U4355 (N_4355,N_3761,N_3882);
and U4356 (N_4356,N_3383,N_3059);
nand U4357 (N_4357,N_3782,N_3167);
nand U4358 (N_4358,N_3809,N_3070);
nor U4359 (N_4359,N_3655,N_3653);
and U4360 (N_4360,N_3916,N_3090);
and U4361 (N_4361,N_3621,N_3515);
nor U4362 (N_4362,N_3969,N_3065);
nand U4363 (N_4363,N_3834,N_3873);
or U4364 (N_4364,N_3987,N_3208);
nor U4365 (N_4365,N_3357,N_3402);
nor U4366 (N_4366,N_3756,N_3640);
nand U4367 (N_4367,N_3330,N_3468);
nor U4368 (N_4368,N_3887,N_3952);
or U4369 (N_4369,N_3865,N_3002);
and U4370 (N_4370,N_3706,N_3466);
nor U4371 (N_4371,N_3554,N_3757);
and U4372 (N_4372,N_3082,N_3028);
and U4373 (N_4373,N_3912,N_3615);
or U4374 (N_4374,N_3794,N_3943);
and U4375 (N_4375,N_3219,N_3945);
nand U4376 (N_4376,N_3048,N_3529);
nor U4377 (N_4377,N_3672,N_3789);
or U4378 (N_4378,N_3479,N_3150);
and U4379 (N_4379,N_3027,N_3004);
or U4380 (N_4380,N_3093,N_3487);
nor U4381 (N_4381,N_3512,N_3441);
nand U4382 (N_4382,N_3074,N_3247);
nor U4383 (N_4383,N_3685,N_3319);
or U4384 (N_4384,N_3893,N_3971);
or U4385 (N_4385,N_3049,N_3700);
and U4386 (N_4386,N_3922,N_3975);
nand U4387 (N_4387,N_3954,N_3409);
nor U4388 (N_4388,N_3846,N_3684);
nor U4389 (N_4389,N_3372,N_3017);
nand U4390 (N_4390,N_3360,N_3439);
nand U4391 (N_4391,N_3433,N_3895);
nor U4392 (N_4392,N_3596,N_3131);
and U4393 (N_4393,N_3504,N_3822);
or U4394 (N_4394,N_3890,N_3449);
nor U4395 (N_4395,N_3638,N_3829);
or U4396 (N_4396,N_3891,N_3941);
nand U4397 (N_4397,N_3000,N_3270);
nor U4398 (N_4398,N_3446,N_3677);
and U4399 (N_4399,N_3149,N_3322);
nand U4400 (N_4400,N_3400,N_3503);
nand U4401 (N_4401,N_3816,N_3939);
nand U4402 (N_4402,N_3811,N_3604);
nor U4403 (N_4403,N_3120,N_3482);
nand U4404 (N_4404,N_3957,N_3113);
xor U4405 (N_4405,N_3746,N_3582);
nand U4406 (N_4406,N_3155,N_3399);
nand U4407 (N_4407,N_3528,N_3820);
xnor U4408 (N_4408,N_3158,N_3428);
nand U4409 (N_4409,N_3966,N_3694);
and U4410 (N_4410,N_3625,N_3754);
or U4411 (N_4411,N_3730,N_3156);
or U4412 (N_4412,N_3725,N_3095);
nand U4413 (N_4413,N_3741,N_3862);
or U4414 (N_4414,N_3238,N_3639);
nor U4415 (N_4415,N_3661,N_3711);
nand U4416 (N_4416,N_3340,N_3239);
or U4417 (N_4417,N_3024,N_3178);
nand U4418 (N_4418,N_3942,N_3673);
and U4419 (N_4419,N_3727,N_3288);
or U4420 (N_4420,N_3365,N_3424);
nor U4421 (N_4421,N_3521,N_3442);
and U4422 (N_4422,N_3458,N_3148);
or U4423 (N_4423,N_3857,N_3808);
and U4424 (N_4424,N_3557,N_3181);
nor U4425 (N_4425,N_3001,N_3143);
nand U4426 (N_4426,N_3060,N_3051);
or U4427 (N_4427,N_3411,N_3382);
or U4428 (N_4428,N_3266,N_3370);
nor U4429 (N_4429,N_3386,N_3520);
or U4430 (N_4430,N_3995,N_3083);
nor U4431 (N_4431,N_3269,N_3109);
nand U4432 (N_4432,N_3321,N_3160);
nor U4433 (N_4433,N_3223,N_3486);
and U4434 (N_4434,N_3900,N_3929);
and U4435 (N_4435,N_3407,N_3871);
nor U4436 (N_4436,N_3855,N_3598);
or U4437 (N_4437,N_3182,N_3687);
nor U4438 (N_4438,N_3726,N_3656);
nor U4439 (N_4439,N_3866,N_3170);
nor U4440 (N_4440,N_3290,N_3549);
and U4441 (N_4441,N_3334,N_3506);
nand U4442 (N_4442,N_3956,N_3749);
nor U4443 (N_4443,N_3415,N_3047);
or U4444 (N_4444,N_3106,N_3630);
nand U4445 (N_4445,N_3443,N_3128);
and U4446 (N_4446,N_3600,N_3686);
or U4447 (N_4447,N_3713,N_3790);
nor U4448 (N_4448,N_3660,N_3151);
or U4449 (N_4449,N_3848,N_3888);
nor U4450 (N_4450,N_3495,N_3135);
nand U4451 (N_4451,N_3121,N_3377);
or U4452 (N_4452,N_3189,N_3681);
and U4453 (N_4453,N_3679,N_3802);
nand U4454 (N_4454,N_3355,N_3698);
nand U4455 (N_4455,N_3552,N_3031);
nor U4456 (N_4456,N_3222,N_3303);
nand U4457 (N_4457,N_3555,N_3792);
or U4458 (N_4458,N_3541,N_3819);
nor U4459 (N_4459,N_3366,N_3720);
nor U4460 (N_4460,N_3963,N_3056);
or U4461 (N_4461,N_3476,N_3892);
and U4462 (N_4462,N_3356,N_3353);
nor U4463 (N_4463,N_3651,N_3705);
nand U4464 (N_4464,N_3421,N_3765);
nor U4465 (N_4465,N_3514,N_3986);
and U4466 (N_4466,N_3913,N_3590);
nand U4467 (N_4467,N_3828,N_3062);
or U4468 (N_4468,N_3974,N_3187);
and U4469 (N_4469,N_3797,N_3299);
nand U4470 (N_4470,N_3102,N_3092);
nor U4471 (N_4471,N_3232,N_3469);
nand U4472 (N_4472,N_3784,N_3996);
and U4473 (N_4473,N_3198,N_3483);
nand U4474 (N_4474,N_3955,N_3745);
xnor U4475 (N_4475,N_3703,N_3798);
or U4476 (N_4476,N_3884,N_3227);
or U4477 (N_4477,N_3404,N_3461);
nand U4478 (N_4478,N_3304,N_3853);
nor U4479 (N_4479,N_3717,N_3958);
and U4480 (N_4480,N_3291,N_3832);
nor U4481 (N_4481,N_3351,N_3526);
nor U4482 (N_4482,N_3931,N_3367);
or U4483 (N_4483,N_3235,N_3680);
nor U4484 (N_4484,N_3306,N_3022);
nand U4485 (N_4485,N_3413,N_3992);
nand U4486 (N_4486,N_3011,N_3164);
or U4487 (N_4487,N_3907,N_3440);
or U4488 (N_4488,N_3315,N_3078);
or U4489 (N_4489,N_3233,N_3225);
or U4490 (N_4490,N_3753,N_3610);
and U4491 (N_4491,N_3813,N_3111);
or U4492 (N_4492,N_3493,N_3243);
nand U4493 (N_4493,N_3831,N_3524);
nor U4494 (N_4494,N_3378,N_3162);
nor U4495 (N_4495,N_3475,N_3184);
nor U4496 (N_4496,N_3063,N_3397);
nor U4497 (N_4497,N_3569,N_3927);
or U4498 (N_4498,N_3134,N_3779);
or U4499 (N_4499,N_3438,N_3246);
and U4500 (N_4500,N_3679,N_3955);
and U4501 (N_4501,N_3145,N_3257);
nand U4502 (N_4502,N_3045,N_3975);
and U4503 (N_4503,N_3150,N_3555);
or U4504 (N_4504,N_3218,N_3889);
nor U4505 (N_4505,N_3696,N_3325);
nand U4506 (N_4506,N_3036,N_3444);
and U4507 (N_4507,N_3221,N_3399);
nand U4508 (N_4508,N_3029,N_3404);
xor U4509 (N_4509,N_3950,N_3735);
nor U4510 (N_4510,N_3316,N_3091);
and U4511 (N_4511,N_3038,N_3542);
nand U4512 (N_4512,N_3934,N_3177);
nor U4513 (N_4513,N_3653,N_3360);
nand U4514 (N_4514,N_3412,N_3390);
or U4515 (N_4515,N_3979,N_3394);
nand U4516 (N_4516,N_3944,N_3986);
nor U4517 (N_4517,N_3232,N_3009);
and U4518 (N_4518,N_3776,N_3403);
or U4519 (N_4519,N_3040,N_3514);
and U4520 (N_4520,N_3107,N_3866);
nor U4521 (N_4521,N_3372,N_3543);
or U4522 (N_4522,N_3325,N_3473);
and U4523 (N_4523,N_3974,N_3139);
and U4524 (N_4524,N_3725,N_3122);
or U4525 (N_4525,N_3874,N_3796);
or U4526 (N_4526,N_3561,N_3601);
nor U4527 (N_4527,N_3747,N_3955);
nor U4528 (N_4528,N_3680,N_3662);
nor U4529 (N_4529,N_3951,N_3272);
and U4530 (N_4530,N_3989,N_3395);
nand U4531 (N_4531,N_3785,N_3916);
nor U4532 (N_4532,N_3961,N_3838);
and U4533 (N_4533,N_3230,N_3833);
nand U4534 (N_4534,N_3385,N_3338);
and U4535 (N_4535,N_3805,N_3424);
or U4536 (N_4536,N_3623,N_3854);
nor U4537 (N_4537,N_3186,N_3115);
or U4538 (N_4538,N_3963,N_3980);
nor U4539 (N_4539,N_3283,N_3598);
nor U4540 (N_4540,N_3045,N_3276);
or U4541 (N_4541,N_3582,N_3913);
and U4542 (N_4542,N_3603,N_3076);
nor U4543 (N_4543,N_3689,N_3351);
nor U4544 (N_4544,N_3224,N_3146);
nand U4545 (N_4545,N_3070,N_3335);
nor U4546 (N_4546,N_3733,N_3601);
and U4547 (N_4547,N_3259,N_3890);
nor U4548 (N_4548,N_3279,N_3465);
nand U4549 (N_4549,N_3137,N_3798);
nor U4550 (N_4550,N_3644,N_3994);
nor U4551 (N_4551,N_3039,N_3988);
nand U4552 (N_4552,N_3203,N_3182);
and U4553 (N_4553,N_3592,N_3429);
or U4554 (N_4554,N_3685,N_3772);
nand U4555 (N_4555,N_3165,N_3997);
nand U4556 (N_4556,N_3675,N_3940);
nand U4557 (N_4557,N_3669,N_3944);
or U4558 (N_4558,N_3976,N_3757);
nand U4559 (N_4559,N_3481,N_3373);
nand U4560 (N_4560,N_3641,N_3620);
xor U4561 (N_4561,N_3963,N_3537);
nor U4562 (N_4562,N_3752,N_3315);
nor U4563 (N_4563,N_3314,N_3883);
and U4564 (N_4564,N_3570,N_3168);
and U4565 (N_4565,N_3021,N_3332);
nor U4566 (N_4566,N_3052,N_3439);
nor U4567 (N_4567,N_3260,N_3745);
xor U4568 (N_4568,N_3250,N_3854);
nand U4569 (N_4569,N_3529,N_3350);
and U4570 (N_4570,N_3583,N_3641);
or U4571 (N_4571,N_3426,N_3401);
and U4572 (N_4572,N_3600,N_3021);
and U4573 (N_4573,N_3910,N_3299);
nand U4574 (N_4574,N_3001,N_3081);
nand U4575 (N_4575,N_3077,N_3175);
nand U4576 (N_4576,N_3030,N_3979);
nor U4577 (N_4577,N_3703,N_3811);
and U4578 (N_4578,N_3482,N_3534);
nand U4579 (N_4579,N_3022,N_3044);
nor U4580 (N_4580,N_3326,N_3720);
nand U4581 (N_4581,N_3031,N_3431);
nand U4582 (N_4582,N_3169,N_3087);
nand U4583 (N_4583,N_3912,N_3450);
and U4584 (N_4584,N_3840,N_3606);
nand U4585 (N_4585,N_3311,N_3910);
nand U4586 (N_4586,N_3566,N_3103);
and U4587 (N_4587,N_3418,N_3348);
and U4588 (N_4588,N_3207,N_3740);
and U4589 (N_4589,N_3203,N_3353);
and U4590 (N_4590,N_3926,N_3502);
nand U4591 (N_4591,N_3295,N_3984);
or U4592 (N_4592,N_3994,N_3178);
nor U4593 (N_4593,N_3246,N_3503);
and U4594 (N_4594,N_3561,N_3929);
nand U4595 (N_4595,N_3107,N_3454);
nand U4596 (N_4596,N_3556,N_3184);
nand U4597 (N_4597,N_3916,N_3981);
nand U4598 (N_4598,N_3153,N_3402);
or U4599 (N_4599,N_3637,N_3525);
nand U4600 (N_4600,N_3553,N_3871);
or U4601 (N_4601,N_3852,N_3403);
or U4602 (N_4602,N_3931,N_3855);
and U4603 (N_4603,N_3412,N_3764);
and U4604 (N_4604,N_3501,N_3970);
nor U4605 (N_4605,N_3395,N_3553);
or U4606 (N_4606,N_3651,N_3328);
or U4607 (N_4607,N_3953,N_3294);
nand U4608 (N_4608,N_3866,N_3359);
nand U4609 (N_4609,N_3854,N_3651);
nor U4610 (N_4610,N_3088,N_3205);
and U4611 (N_4611,N_3730,N_3593);
or U4612 (N_4612,N_3296,N_3875);
nor U4613 (N_4613,N_3306,N_3094);
nand U4614 (N_4614,N_3142,N_3222);
nand U4615 (N_4615,N_3422,N_3982);
or U4616 (N_4616,N_3823,N_3637);
nor U4617 (N_4617,N_3725,N_3774);
or U4618 (N_4618,N_3476,N_3523);
nand U4619 (N_4619,N_3047,N_3610);
nand U4620 (N_4620,N_3164,N_3316);
and U4621 (N_4621,N_3241,N_3036);
or U4622 (N_4622,N_3897,N_3856);
nand U4623 (N_4623,N_3445,N_3629);
or U4624 (N_4624,N_3676,N_3359);
or U4625 (N_4625,N_3204,N_3655);
or U4626 (N_4626,N_3469,N_3873);
and U4627 (N_4627,N_3970,N_3572);
and U4628 (N_4628,N_3007,N_3293);
or U4629 (N_4629,N_3854,N_3598);
nand U4630 (N_4630,N_3055,N_3815);
and U4631 (N_4631,N_3094,N_3881);
or U4632 (N_4632,N_3770,N_3126);
and U4633 (N_4633,N_3468,N_3284);
nor U4634 (N_4634,N_3007,N_3903);
or U4635 (N_4635,N_3804,N_3654);
and U4636 (N_4636,N_3087,N_3725);
and U4637 (N_4637,N_3974,N_3151);
nand U4638 (N_4638,N_3617,N_3541);
nor U4639 (N_4639,N_3378,N_3660);
and U4640 (N_4640,N_3657,N_3606);
nand U4641 (N_4641,N_3567,N_3053);
nor U4642 (N_4642,N_3499,N_3968);
and U4643 (N_4643,N_3434,N_3640);
nand U4644 (N_4644,N_3433,N_3779);
nand U4645 (N_4645,N_3786,N_3388);
and U4646 (N_4646,N_3880,N_3894);
xnor U4647 (N_4647,N_3455,N_3754);
nor U4648 (N_4648,N_3027,N_3150);
and U4649 (N_4649,N_3230,N_3255);
and U4650 (N_4650,N_3236,N_3741);
nor U4651 (N_4651,N_3829,N_3818);
nand U4652 (N_4652,N_3472,N_3572);
nor U4653 (N_4653,N_3721,N_3661);
or U4654 (N_4654,N_3474,N_3063);
nand U4655 (N_4655,N_3973,N_3268);
or U4656 (N_4656,N_3527,N_3203);
or U4657 (N_4657,N_3730,N_3114);
nand U4658 (N_4658,N_3773,N_3496);
nor U4659 (N_4659,N_3751,N_3133);
or U4660 (N_4660,N_3951,N_3036);
nand U4661 (N_4661,N_3159,N_3471);
nand U4662 (N_4662,N_3545,N_3859);
nor U4663 (N_4663,N_3142,N_3934);
or U4664 (N_4664,N_3811,N_3118);
nand U4665 (N_4665,N_3192,N_3382);
and U4666 (N_4666,N_3200,N_3615);
and U4667 (N_4667,N_3791,N_3958);
nor U4668 (N_4668,N_3668,N_3705);
and U4669 (N_4669,N_3616,N_3402);
or U4670 (N_4670,N_3326,N_3304);
nand U4671 (N_4671,N_3590,N_3736);
and U4672 (N_4672,N_3120,N_3295);
nor U4673 (N_4673,N_3618,N_3400);
or U4674 (N_4674,N_3893,N_3941);
nand U4675 (N_4675,N_3899,N_3159);
nor U4676 (N_4676,N_3134,N_3578);
and U4677 (N_4677,N_3219,N_3601);
or U4678 (N_4678,N_3170,N_3741);
nor U4679 (N_4679,N_3708,N_3215);
or U4680 (N_4680,N_3418,N_3735);
nor U4681 (N_4681,N_3913,N_3647);
or U4682 (N_4682,N_3627,N_3272);
or U4683 (N_4683,N_3292,N_3329);
nand U4684 (N_4684,N_3607,N_3901);
or U4685 (N_4685,N_3836,N_3924);
and U4686 (N_4686,N_3987,N_3633);
nand U4687 (N_4687,N_3393,N_3239);
and U4688 (N_4688,N_3776,N_3352);
nor U4689 (N_4689,N_3688,N_3064);
nor U4690 (N_4690,N_3314,N_3262);
nor U4691 (N_4691,N_3494,N_3258);
nand U4692 (N_4692,N_3263,N_3223);
or U4693 (N_4693,N_3169,N_3725);
nor U4694 (N_4694,N_3903,N_3918);
nor U4695 (N_4695,N_3863,N_3787);
nor U4696 (N_4696,N_3059,N_3467);
and U4697 (N_4697,N_3274,N_3989);
and U4698 (N_4698,N_3202,N_3064);
nand U4699 (N_4699,N_3965,N_3948);
or U4700 (N_4700,N_3833,N_3466);
or U4701 (N_4701,N_3420,N_3276);
or U4702 (N_4702,N_3355,N_3389);
or U4703 (N_4703,N_3631,N_3371);
or U4704 (N_4704,N_3329,N_3405);
nand U4705 (N_4705,N_3084,N_3882);
or U4706 (N_4706,N_3375,N_3197);
nand U4707 (N_4707,N_3363,N_3623);
and U4708 (N_4708,N_3584,N_3685);
nand U4709 (N_4709,N_3915,N_3676);
nand U4710 (N_4710,N_3638,N_3846);
nand U4711 (N_4711,N_3083,N_3161);
nor U4712 (N_4712,N_3057,N_3094);
nor U4713 (N_4713,N_3911,N_3153);
nor U4714 (N_4714,N_3131,N_3284);
nor U4715 (N_4715,N_3776,N_3089);
and U4716 (N_4716,N_3569,N_3537);
nand U4717 (N_4717,N_3991,N_3070);
and U4718 (N_4718,N_3066,N_3171);
and U4719 (N_4719,N_3530,N_3515);
nor U4720 (N_4720,N_3683,N_3950);
nor U4721 (N_4721,N_3608,N_3975);
or U4722 (N_4722,N_3192,N_3096);
or U4723 (N_4723,N_3163,N_3493);
or U4724 (N_4724,N_3196,N_3430);
and U4725 (N_4725,N_3220,N_3288);
or U4726 (N_4726,N_3244,N_3355);
nand U4727 (N_4727,N_3710,N_3212);
nor U4728 (N_4728,N_3346,N_3676);
nand U4729 (N_4729,N_3587,N_3481);
nand U4730 (N_4730,N_3525,N_3017);
nand U4731 (N_4731,N_3042,N_3632);
nor U4732 (N_4732,N_3756,N_3308);
nor U4733 (N_4733,N_3438,N_3124);
nand U4734 (N_4734,N_3831,N_3336);
nor U4735 (N_4735,N_3321,N_3809);
nand U4736 (N_4736,N_3738,N_3633);
or U4737 (N_4737,N_3060,N_3127);
or U4738 (N_4738,N_3147,N_3107);
or U4739 (N_4739,N_3147,N_3771);
or U4740 (N_4740,N_3179,N_3459);
nand U4741 (N_4741,N_3573,N_3152);
and U4742 (N_4742,N_3198,N_3630);
and U4743 (N_4743,N_3136,N_3685);
nand U4744 (N_4744,N_3321,N_3102);
xnor U4745 (N_4745,N_3736,N_3259);
or U4746 (N_4746,N_3752,N_3478);
or U4747 (N_4747,N_3042,N_3712);
nand U4748 (N_4748,N_3567,N_3638);
nor U4749 (N_4749,N_3000,N_3794);
nor U4750 (N_4750,N_3454,N_3987);
nand U4751 (N_4751,N_3836,N_3940);
nand U4752 (N_4752,N_3930,N_3268);
nor U4753 (N_4753,N_3057,N_3159);
nand U4754 (N_4754,N_3014,N_3957);
nand U4755 (N_4755,N_3011,N_3840);
and U4756 (N_4756,N_3606,N_3669);
nand U4757 (N_4757,N_3687,N_3231);
and U4758 (N_4758,N_3050,N_3023);
nand U4759 (N_4759,N_3804,N_3306);
nand U4760 (N_4760,N_3370,N_3879);
nor U4761 (N_4761,N_3486,N_3360);
and U4762 (N_4762,N_3475,N_3804);
nor U4763 (N_4763,N_3461,N_3325);
or U4764 (N_4764,N_3635,N_3369);
nor U4765 (N_4765,N_3161,N_3009);
nand U4766 (N_4766,N_3677,N_3508);
nor U4767 (N_4767,N_3555,N_3382);
nor U4768 (N_4768,N_3551,N_3103);
nor U4769 (N_4769,N_3394,N_3982);
nor U4770 (N_4770,N_3826,N_3082);
nand U4771 (N_4771,N_3041,N_3780);
nand U4772 (N_4772,N_3171,N_3581);
xor U4773 (N_4773,N_3869,N_3226);
and U4774 (N_4774,N_3683,N_3385);
nand U4775 (N_4775,N_3692,N_3289);
nor U4776 (N_4776,N_3583,N_3846);
nand U4777 (N_4777,N_3955,N_3463);
nand U4778 (N_4778,N_3157,N_3152);
and U4779 (N_4779,N_3523,N_3313);
nor U4780 (N_4780,N_3390,N_3799);
and U4781 (N_4781,N_3508,N_3572);
nor U4782 (N_4782,N_3540,N_3572);
nand U4783 (N_4783,N_3328,N_3932);
nor U4784 (N_4784,N_3565,N_3354);
or U4785 (N_4785,N_3822,N_3538);
or U4786 (N_4786,N_3592,N_3813);
or U4787 (N_4787,N_3021,N_3503);
or U4788 (N_4788,N_3456,N_3137);
nor U4789 (N_4789,N_3958,N_3831);
and U4790 (N_4790,N_3405,N_3719);
or U4791 (N_4791,N_3954,N_3627);
nor U4792 (N_4792,N_3189,N_3013);
nor U4793 (N_4793,N_3237,N_3823);
or U4794 (N_4794,N_3877,N_3398);
xnor U4795 (N_4795,N_3364,N_3086);
nand U4796 (N_4796,N_3965,N_3073);
nand U4797 (N_4797,N_3590,N_3893);
nand U4798 (N_4798,N_3778,N_3624);
or U4799 (N_4799,N_3409,N_3382);
nor U4800 (N_4800,N_3572,N_3632);
and U4801 (N_4801,N_3129,N_3238);
nand U4802 (N_4802,N_3590,N_3081);
nand U4803 (N_4803,N_3768,N_3906);
xor U4804 (N_4804,N_3188,N_3435);
nor U4805 (N_4805,N_3207,N_3590);
nor U4806 (N_4806,N_3145,N_3123);
and U4807 (N_4807,N_3669,N_3819);
nor U4808 (N_4808,N_3408,N_3959);
nor U4809 (N_4809,N_3688,N_3632);
nor U4810 (N_4810,N_3768,N_3252);
or U4811 (N_4811,N_3781,N_3791);
or U4812 (N_4812,N_3781,N_3930);
or U4813 (N_4813,N_3109,N_3988);
and U4814 (N_4814,N_3460,N_3696);
or U4815 (N_4815,N_3880,N_3521);
or U4816 (N_4816,N_3900,N_3804);
and U4817 (N_4817,N_3342,N_3544);
or U4818 (N_4818,N_3231,N_3715);
nor U4819 (N_4819,N_3267,N_3621);
nor U4820 (N_4820,N_3341,N_3463);
nand U4821 (N_4821,N_3994,N_3542);
nor U4822 (N_4822,N_3804,N_3399);
or U4823 (N_4823,N_3920,N_3958);
or U4824 (N_4824,N_3724,N_3605);
nor U4825 (N_4825,N_3771,N_3217);
nor U4826 (N_4826,N_3886,N_3219);
and U4827 (N_4827,N_3193,N_3038);
and U4828 (N_4828,N_3415,N_3398);
or U4829 (N_4829,N_3894,N_3278);
and U4830 (N_4830,N_3021,N_3980);
nand U4831 (N_4831,N_3751,N_3956);
nand U4832 (N_4832,N_3242,N_3176);
nand U4833 (N_4833,N_3661,N_3413);
nor U4834 (N_4834,N_3602,N_3487);
and U4835 (N_4835,N_3514,N_3135);
nand U4836 (N_4836,N_3156,N_3776);
nand U4837 (N_4837,N_3816,N_3561);
nand U4838 (N_4838,N_3975,N_3484);
nor U4839 (N_4839,N_3262,N_3162);
nand U4840 (N_4840,N_3654,N_3022);
nand U4841 (N_4841,N_3142,N_3824);
or U4842 (N_4842,N_3422,N_3264);
and U4843 (N_4843,N_3562,N_3953);
or U4844 (N_4844,N_3687,N_3272);
nand U4845 (N_4845,N_3740,N_3209);
nor U4846 (N_4846,N_3183,N_3394);
and U4847 (N_4847,N_3433,N_3888);
and U4848 (N_4848,N_3890,N_3891);
and U4849 (N_4849,N_3033,N_3671);
and U4850 (N_4850,N_3324,N_3988);
or U4851 (N_4851,N_3013,N_3073);
nand U4852 (N_4852,N_3571,N_3144);
or U4853 (N_4853,N_3656,N_3847);
and U4854 (N_4854,N_3342,N_3517);
nand U4855 (N_4855,N_3780,N_3530);
or U4856 (N_4856,N_3216,N_3072);
and U4857 (N_4857,N_3386,N_3361);
or U4858 (N_4858,N_3063,N_3975);
nor U4859 (N_4859,N_3638,N_3956);
or U4860 (N_4860,N_3784,N_3117);
nor U4861 (N_4861,N_3417,N_3463);
or U4862 (N_4862,N_3156,N_3941);
nand U4863 (N_4863,N_3923,N_3885);
or U4864 (N_4864,N_3920,N_3929);
or U4865 (N_4865,N_3402,N_3230);
nor U4866 (N_4866,N_3923,N_3916);
or U4867 (N_4867,N_3655,N_3954);
nand U4868 (N_4868,N_3424,N_3130);
and U4869 (N_4869,N_3339,N_3409);
or U4870 (N_4870,N_3424,N_3046);
or U4871 (N_4871,N_3788,N_3146);
nor U4872 (N_4872,N_3282,N_3137);
nand U4873 (N_4873,N_3088,N_3243);
nand U4874 (N_4874,N_3052,N_3303);
or U4875 (N_4875,N_3320,N_3345);
nor U4876 (N_4876,N_3112,N_3323);
nand U4877 (N_4877,N_3269,N_3193);
nand U4878 (N_4878,N_3698,N_3670);
nor U4879 (N_4879,N_3874,N_3691);
or U4880 (N_4880,N_3391,N_3327);
and U4881 (N_4881,N_3347,N_3235);
nor U4882 (N_4882,N_3905,N_3501);
nor U4883 (N_4883,N_3083,N_3400);
nand U4884 (N_4884,N_3022,N_3650);
nor U4885 (N_4885,N_3269,N_3948);
and U4886 (N_4886,N_3524,N_3693);
nor U4887 (N_4887,N_3126,N_3552);
and U4888 (N_4888,N_3579,N_3566);
nor U4889 (N_4889,N_3989,N_3929);
nand U4890 (N_4890,N_3281,N_3174);
or U4891 (N_4891,N_3832,N_3398);
nor U4892 (N_4892,N_3247,N_3713);
nand U4893 (N_4893,N_3957,N_3394);
nor U4894 (N_4894,N_3794,N_3054);
nand U4895 (N_4895,N_3467,N_3386);
or U4896 (N_4896,N_3439,N_3010);
or U4897 (N_4897,N_3601,N_3899);
and U4898 (N_4898,N_3781,N_3315);
nor U4899 (N_4899,N_3675,N_3029);
or U4900 (N_4900,N_3961,N_3567);
or U4901 (N_4901,N_3837,N_3510);
and U4902 (N_4902,N_3535,N_3258);
nand U4903 (N_4903,N_3261,N_3581);
or U4904 (N_4904,N_3849,N_3619);
and U4905 (N_4905,N_3349,N_3529);
or U4906 (N_4906,N_3666,N_3098);
nor U4907 (N_4907,N_3055,N_3188);
or U4908 (N_4908,N_3533,N_3210);
nand U4909 (N_4909,N_3317,N_3891);
and U4910 (N_4910,N_3708,N_3205);
and U4911 (N_4911,N_3142,N_3642);
nand U4912 (N_4912,N_3151,N_3798);
and U4913 (N_4913,N_3982,N_3330);
or U4914 (N_4914,N_3598,N_3634);
and U4915 (N_4915,N_3628,N_3431);
nand U4916 (N_4916,N_3895,N_3234);
nor U4917 (N_4917,N_3170,N_3370);
or U4918 (N_4918,N_3076,N_3895);
and U4919 (N_4919,N_3499,N_3703);
and U4920 (N_4920,N_3799,N_3463);
and U4921 (N_4921,N_3194,N_3070);
nor U4922 (N_4922,N_3183,N_3295);
nand U4923 (N_4923,N_3551,N_3323);
or U4924 (N_4924,N_3384,N_3435);
nand U4925 (N_4925,N_3358,N_3130);
nand U4926 (N_4926,N_3272,N_3760);
or U4927 (N_4927,N_3433,N_3657);
nand U4928 (N_4928,N_3536,N_3173);
nand U4929 (N_4929,N_3980,N_3233);
or U4930 (N_4930,N_3588,N_3930);
nor U4931 (N_4931,N_3304,N_3225);
and U4932 (N_4932,N_3549,N_3345);
or U4933 (N_4933,N_3866,N_3531);
nand U4934 (N_4934,N_3687,N_3512);
nand U4935 (N_4935,N_3148,N_3093);
nor U4936 (N_4936,N_3129,N_3170);
nand U4937 (N_4937,N_3561,N_3759);
nor U4938 (N_4938,N_3376,N_3477);
and U4939 (N_4939,N_3458,N_3096);
and U4940 (N_4940,N_3531,N_3070);
or U4941 (N_4941,N_3333,N_3104);
and U4942 (N_4942,N_3460,N_3931);
or U4943 (N_4943,N_3459,N_3029);
nor U4944 (N_4944,N_3088,N_3937);
and U4945 (N_4945,N_3010,N_3691);
nor U4946 (N_4946,N_3680,N_3330);
nor U4947 (N_4947,N_3031,N_3523);
and U4948 (N_4948,N_3786,N_3992);
nand U4949 (N_4949,N_3318,N_3433);
nor U4950 (N_4950,N_3803,N_3990);
nor U4951 (N_4951,N_3143,N_3537);
nand U4952 (N_4952,N_3705,N_3129);
and U4953 (N_4953,N_3717,N_3527);
and U4954 (N_4954,N_3033,N_3272);
nand U4955 (N_4955,N_3966,N_3062);
or U4956 (N_4956,N_3351,N_3243);
or U4957 (N_4957,N_3754,N_3503);
and U4958 (N_4958,N_3994,N_3951);
or U4959 (N_4959,N_3933,N_3458);
nand U4960 (N_4960,N_3956,N_3458);
nor U4961 (N_4961,N_3635,N_3504);
or U4962 (N_4962,N_3937,N_3126);
or U4963 (N_4963,N_3934,N_3915);
nor U4964 (N_4964,N_3401,N_3502);
or U4965 (N_4965,N_3120,N_3490);
nor U4966 (N_4966,N_3776,N_3529);
or U4967 (N_4967,N_3450,N_3978);
nor U4968 (N_4968,N_3981,N_3448);
or U4969 (N_4969,N_3831,N_3935);
nand U4970 (N_4970,N_3287,N_3176);
nor U4971 (N_4971,N_3516,N_3815);
nand U4972 (N_4972,N_3610,N_3160);
nor U4973 (N_4973,N_3981,N_3089);
or U4974 (N_4974,N_3333,N_3875);
and U4975 (N_4975,N_3398,N_3103);
nand U4976 (N_4976,N_3398,N_3710);
or U4977 (N_4977,N_3358,N_3896);
nand U4978 (N_4978,N_3787,N_3620);
nand U4979 (N_4979,N_3277,N_3564);
and U4980 (N_4980,N_3943,N_3634);
nor U4981 (N_4981,N_3819,N_3832);
and U4982 (N_4982,N_3392,N_3736);
nand U4983 (N_4983,N_3287,N_3964);
nand U4984 (N_4984,N_3888,N_3699);
nand U4985 (N_4985,N_3202,N_3518);
nand U4986 (N_4986,N_3734,N_3221);
and U4987 (N_4987,N_3072,N_3340);
nor U4988 (N_4988,N_3955,N_3749);
or U4989 (N_4989,N_3054,N_3863);
nand U4990 (N_4990,N_3942,N_3046);
and U4991 (N_4991,N_3693,N_3684);
nor U4992 (N_4992,N_3886,N_3796);
and U4993 (N_4993,N_3865,N_3544);
or U4994 (N_4994,N_3469,N_3713);
and U4995 (N_4995,N_3010,N_3094);
nand U4996 (N_4996,N_3351,N_3824);
nand U4997 (N_4997,N_3217,N_3461);
nor U4998 (N_4998,N_3057,N_3800);
or U4999 (N_4999,N_3419,N_3908);
nand U5000 (N_5000,N_4715,N_4159);
nand U5001 (N_5001,N_4095,N_4708);
or U5002 (N_5002,N_4440,N_4416);
nand U5003 (N_5003,N_4814,N_4300);
nand U5004 (N_5004,N_4997,N_4446);
nor U5005 (N_5005,N_4077,N_4692);
or U5006 (N_5006,N_4928,N_4459);
or U5007 (N_5007,N_4114,N_4398);
nand U5008 (N_5008,N_4029,N_4962);
and U5009 (N_5009,N_4554,N_4979);
or U5010 (N_5010,N_4295,N_4000);
and U5011 (N_5011,N_4031,N_4690);
nor U5012 (N_5012,N_4966,N_4901);
or U5013 (N_5013,N_4863,N_4004);
nor U5014 (N_5014,N_4206,N_4591);
and U5015 (N_5015,N_4856,N_4162);
nand U5016 (N_5016,N_4353,N_4054);
or U5017 (N_5017,N_4084,N_4164);
nor U5018 (N_5018,N_4977,N_4243);
nor U5019 (N_5019,N_4713,N_4804);
and U5020 (N_5020,N_4303,N_4677);
nor U5021 (N_5021,N_4891,N_4697);
nand U5022 (N_5022,N_4800,N_4781);
and U5023 (N_5023,N_4465,N_4755);
nand U5024 (N_5024,N_4847,N_4887);
and U5025 (N_5025,N_4382,N_4080);
nor U5026 (N_5026,N_4128,N_4870);
or U5027 (N_5027,N_4504,N_4925);
and U5028 (N_5028,N_4920,N_4195);
or U5029 (N_5029,N_4593,N_4457);
nand U5030 (N_5030,N_4628,N_4638);
nand U5031 (N_5031,N_4896,N_4409);
or U5032 (N_5032,N_4245,N_4536);
or U5033 (N_5033,N_4744,N_4189);
nand U5034 (N_5034,N_4970,N_4795);
or U5035 (N_5035,N_4914,N_4170);
nor U5036 (N_5036,N_4100,N_4249);
nand U5037 (N_5037,N_4130,N_4293);
nor U5038 (N_5038,N_4540,N_4579);
nand U5039 (N_5039,N_4949,N_4855);
nand U5040 (N_5040,N_4771,N_4493);
nand U5041 (N_5041,N_4684,N_4965);
and U5042 (N_5042,N_4972,N_4786);
or U5043 (N_5043,N_4803,N_4263);
nand U5044 (N_5044,N_4287,N_4065);
and U5045 (N_5045,N_4611,N_4655);
and U5046 (N_5046,N_4422,N_4840);
nor U5047 (N_5047,N_4028,N_4710);
nor U5048 (N_5048,N_4144,N_4559);
nor U5049 (N_5049,N_4044,N_4235);
nand U5050 (N_5050,N_4403,N_4799);
nand U5051 (N_5051,N_4435,N_4318);
or U5052 (N_5052,N_4760,N_4305);
and U5053 (N_5053,N_4034,N_4228);
nand U5054 (N_5054,N_4212,N_4889);
nand U5055 (N_5055,N_4820,N_4074);
or U5056 (N_5056,N_4464,N_4735);
or U5057 (N_5057,N_4973,N_4311);
nand U5058 (N_5058,N_4665,N_4830);
or U5059 (N_5059,N_4660,N_4132);
and U5060 (N_5060,N_4227,N_4268);
and U5061 (N_5061,N_4201,N_4815);
nor U5062 (N_5062,N_4340,N_4753);
and U5063 (N_5063,N_4556,N_4161);
and U5064 (N_5064,N_4401,N_4989);
and U5065 (N_5065,N_4772,N_4936);
nor U5066 (N_5066,N_4653,N_4298);
nor U5067 (N_5067,N_4903,N_4023);
nor U5068 (N_5068,N_4750,N_4853);
nand U5069 (N_5069,N_4687,N_4876);
nor U5070 (N_5070,N_4109,N_4939);
nand U5071 (N_5071,N_4551,N_4354);
nor U5072 (N_5072,N_4886,N_4788);
nor U5073 (N_5073,N_4127,N_4385);
and U5074 (N_5074,N_4614,N_4154);
nand U5075 (N_5075,N_4501,N_4766);
and U5076 (N_5076,N_4905,N_4499);
nor U5077 (N_5077,N_4240,N_4476);
nand U5078 (N_5078,N_4296,N_4995);
or U5079 (N_5079,N_4012,N_4445);
nor U5080 (N_5080,N_4884,N_4819);
and U5081 (N_5081,N_4858,N_4583);
and U5082 (N_5082,N_4654,N_4711);
and U5083 (N_5083,N_4328,N_4125);
or U5084 (N_5084,N_4273,N_4014);
nor U5085 (N_5085,N_4265,N_4165);
or U5086 (N_5086,N_4941,N_4810);
nor U5087 (N_5087,N_4112,N_4906);
nor U5088 (N_5088,N_4651,N_4289);
or U5089 (N_5089,N_4529,N_4010);
nand U5090 (N_5090,N_4907,N_4141);
nand U5091 (N_5091,N_4242,N_4473);
and U5092 (N_5092,N_4344,N_4573);
and U5093 (N_5093,N_4734,N_4616);
or U5094 (N_5094,N_4151,N_4454);
nand U5095 (N_5095,N_4836,N_4937);
nand U5096 (N_5096,N_4261,N_4759);
xor U5097 (N_5097,N_4661,N_4738);
nor U5098 (N_5098,N_4775,N_4236);
nand U5099 (N_5099,N_4520,N_4498);
nand U5100 (N_5100,N_4363,N_4866);
and U5101 (N_5101,N_4740,N_4873);
nor U5102 (N_5102,N_4862,N_4481);
or U5103 (N_5103,N_4003,N_4105);
nor U5104 (N_5104,N_4073,N_4177);
and U5105 (N_5105,N_4592,N_4066);
nand U5106 (N_5106,N_4299,N_4883);
and U5107 (N_5107,N_4586,N_4680);
nand U5108 (N_5108,N_4857,N_4461);
nand U5109 (N_5109,N_4221,N_4868);
nor U5110 (N_5110,N_4895,N_4676);
and U5111 (N_5111,N_4247,N_4779);
and U5112 (N_5112,N_4533,N_4269);
or U5113 (N_5113,N_4013,N_4005);
nand U5114 (N_5114,N_4349,N_4570);
nor U5115 (N_5115,N_4069,N_4279);
nand U5116 (N_5116,N_4686,N_4731);
nor U5117 (N_5117,N_4399,N_4094);
and U5118 (N_5118,N_4267,N_4754);
nand U5119 (N_5119,N_4329,N_4657);
or U5120 (N_5120,N_4537,N_4530);
xnor U5121 (N_5121,N_4612,N_4444);
nor U5122 (N_5122,N_4449,N_4341);
and U5123 (N_5123,N_4531,N_4514);
or U5124 (N_5124,N_4769,N_4669);
or U5125 (N_5125,N_4270,N_4811);
and U5126 (N_5126,N_4333,N_4765);
and U5127 (N_5127,N_4429,N_4027);
and U5128 (N_5128,N_4550,N_4637);
or U5129 (N_5129,N_4641,N_4081);
and U5130 (N_5130,N_4926,N_4699);
and U5131 (N_5131,N_4487,N_4496);
nor U5132 (N_5132,N_4679,N_4575);
nor U5133 (N_5133,N_4272,N_4251);
nand U5134 (N_5134,N_4248,N_4780);
nand U5135 (N_5135,N_4945,N_4695);
and U5136 (N_5136,N_4275,N_4597);
and U5137 (N_5137,N_4698,N_4336);
nor U5138 (N_5138,N_4745,N_4996);
nor U5139 (N_5139,N_4670,N_4683);
nor U5140 (N_5140,N_4075,N_4838);
nand U5141 (N_5141,N_4601,N_4813);
nand U5142 (N_5142,N_4549,N_4246);
or U5143 (N_5143,N_4384,N_4584);
nand U5144 (N_5144,N_4721,N_4992);
and U5145 (N_5145,N_4229,N_4867);
and U5146 (N_5146,N_4430,N_4707);
nor U5147 (N_5147,N_4960,N_4264);
or U5148 (N_5148,N_4046,N_4747);
or U5149 (N_5149,N_4358,N_4291);
and U5150 (N_5150,N_4739,N_4136);
and U5151 (N_5151,N_4033,N_4523);
nor U5152 (N_5152,N_4223,N_4567);
xor U5153 (N_5153,N_4436,N_4041);
nor U5154 (N_5154,N_4338,N_4681);
nor U5155 (N_5155,N_4178,N_4304);
nand U5156 (N_5156,N_4527,N_4039);
nor U5157 (N_5157,N_4600,N_4950);
nand U5158 (N_5158,N_4122,N_4623);
nor U5159 (N_5159,N_4281,N_4405);
nand U5160 (N_5160,N_4426,N_4659);
and U5161 (N_5161,N_4630,N_4629);
nand U5162 (N_5162,N_4667,N_4673);
or U5163 (N_5163,N_4088,N_4411);
nand U5164 (N_5164,N_4434,N_4480);
nand U5165 (N_5165,N_4139,N_4598);
or U5166 (N_5166,N_4952,N_4194);
nand U5167 (N_5167,N_4390,N_4563);
and U5168 (N_5168,N_4233,N_4326);
and U5169 (N_5169,N_4448,N_4288);
nand U5170 (N_5170,N_4809,N_4343);
or U5171 (N_5171,N_4850,N_4851);
or U5172 (N_5172,N_4622,N_4124);
xnor U5173 (N_5173,N_4045,N_4050);
or U5174 (N_5174,N_4726,N_4322);
nand U5175 (N_5175,N_4463,N_4730);
nand U5176 (N_5176,N_4736,N_4576);
nor U5177 (N_5177,N_4916,N_4404);
nor U5178 (N_5178,N_4208,N_4179);
and U5179 (N_5179,N_4560,N_4143);
and U5180 (N_5180,N_4763,N_4828);
nor U5181 (N_5181,N_4947,N_4668);
nor U5182 (N_5182,N_4967,N_4256);
and U5183 (N_5183,N_4852,N_4181);
nor U5184 (N_5184,N_4990,N_4596);
and U5185 (N_5185,N_4935,N_4986);
or U5186 (N_5186,N_4368,N_4595);
or U5187 (N_5187,N_4059,N_4477);
nor U5188 (N_5188,N_4488,N_4145);
or U5189 (N_5189,N_4762,N_4585);
or U5190 (N_5190,N_4790,N_4716);
or U5191 (N_5191,N_4571,N_4787);
or U5192 (N_5192,N_4024,N_4047);
and U5193 (N_5193,N_4331,N_4861);
and U5194 (N_5194,N_4521,N_4522);
or U5195 (N_5195,N_4006,N_4097);
nand U5196 (N_5196,N_4717,N_4250);
nand U5197 (N_5197,N_4147,N_4020);
or U5198 (N_5198,N_4335,N_4696);
nand U5199 (N_5199,N_4196,N_4016);
or U5200 (N_5200,N_4266,N_4361);
nor U5201 (N_5201,N_4482,N_4175);
nand U5202 (N_5202,N_4455,N_4961);
nor U5203 (N_5203,N_4371,N_4207);
or U5204 (N_5204,N_4627,N_4718);
or U5205 (N_5205,N_4366,N_4152);
nor U5206 (N_5206,N_4509,N_4462);
nand U5207 (N_5207,N_4802,N_4241);
nand U5208 (N_5208,N_4479,N_4214);
nand U5209 (N_5209,N_4982,N_4816);
or U5210 (N_5210,N_4484,N_4342);
nor U5211 (N_5211,N_4534,N_4607);
nor U5212 (N_5212,N_4259,N_4749);
and U5213 (N_5213,N_4829,N_4632);
nor U5214 (N_5214,N_4388,N_4032);
and U5215 (N_5215,N_4980,N_4347);
nand U5216 (N_5216,N_4098,N_4915);
nand U5217 (N_5217,N_4994,N_4352);
nand U5218 (N_5218,N_4211,N_4386);
nor U5219 (N_5219,N_4225,N_4116);
and U5220 (N_5220,N_4458,N_4346);
or U5221 (N_5221,N_4126,N_4515);
nand U5222 (N_5222,N_4091,N_4923);
and U5223 (N_5223,N_4337,N_4513);
and U5224 (N_5224,N_4378,N_4674);
nand U5225 (N_5225,N_4869,N_4035);
or U5226 (N_5226,N_4778,N_4555);
or U5227 (N_5227,N_4334,N_4140);
nand U5228 (N_5228,N_4313,N_4257);
nor U5229 (N_5229,N_4693,N_4090);
nor U5230 (N_5230,N_4737,N_4437);
and U5231 (N_5231,N_4700,N_4002);
and U5232 (N_5232,N_4543,N_4215);
or U5233 (N_5233,N_4443,N_4969);
and U5234 (N_5234,N_4118,N_4723);
and U5235 (N_5235,N_4425,N_4541);
or U5236 (N_5236,N_4193,N_4805);
or U5237 (N_5237,N_4649,N_4774);
nor U5238 (N_5238,N_4691,N_4625);
or U5239 (N_5239,N_4226,N_4061);
xnor U5240 (N_5240,N_4017,N_4834);
nor U5241 (N_5241,N_4260,N_4874);
or U5242 (N_5242,N_4198,N_4049);
or U5243 (N_5243,N_4284,N_4581);
or U5244 (N_5244,N_4183,N_4909);
and U5245 (N_5245,N_4042,N_4030);
or U5246 (N_5246,N_4146,N_4733);
and U5247 (N_5247,N_4350,N_4213);
or U5248 (N_5248,N_4782,N_4741);
nor U5249 (N_5249,N_4978,N_4964);
nor U5250 (N_5250,N_4546,N_4647);
or U5251 (N_5251,N_4101,N_4040);
and U5252 (N_5252,N_4392,N_4312);
and U5253 (N_5253,N_4357,N_4930);
or U5254 (N_5254,N_4468,N_4639);
or U5255 (N_5255,N_4872,N_4106);
and U5256 (N_5256,N_4943,N_4704);
nor U5257 (N_5257,N_4899,N_4929);
and U5258 (N_5258,N_4824,N_4566);
nand U5259 (N_5259,N_4156,N_4238);
nor U5260 (N_5260,N_4325,N_4957);
nor U5261 (N_5261,N_4441,N_4784);
nand U5262 (N_5262,N_4577,N_4280);
nand U5263 (N_5263,N_4910,N_4317);
or U5264 (N_5264,N_4432,N_4569);
nor U5265 (N_5265,N_4383,N_4806);
nand U5266 (N_5266,N_4672,N_4609);
nand U5267 (N_5267,N_4283,N_4688);
or U5268 (N_5268,N_4330,N_4316);
nor U5269 (N_5269,N_4424,N_4190);
nor U5270 (N_5270,N_4773,N_4018);
nand U5271 (N_5271,N_4702,N_4083);
nand U5272 (N_5272,N_4643,N_4666);
or U5273 (N_5273,N_4051,N_4324);
or U5274 (N_5274,N_4135,N_4934);
or U5275 (N_5275,N_4808,N_4348);
or U5276 (N_5276,N_4599,N_4525);
or U5277 (N_5277,N_4290,N_4558);
nand U5278 (N_5278,N_4848,N_4489);
and U5279 (N_5279,N_4645,N_4955);
nor U5280 (N_5280,N_4068,N_4492);
and U5281 (N_5281,N_4608,N_4714);
nor U5282 (N_5282,N_4648,N_4319);
nor U5283 (N_5283,N_4203,N_4142);
nand U5284 (N_5284,N_4842,N_4911);
or U5285 (N_5285,N_4987,N_4535);
or U5286 (N_5286,N_4332,N_4174);
nor U5287 (N_5287,N_4991,N_4797);
nor U5288 (N_5288,N_4373,N_4603);
nor U5289 (N_5289,N_4913,N_4633);
or U5290 (N_5290,N_4224,N_4621);
and U5291 (N_5291,N_4274,N_4355);
nand U5292 (N_5292,N_4940,N_4552);
nand U5293 (N_5293,N_4180,N_4137);
nand U5294 (N_5294,N_4709,N_4120);
nor U5295 (N_5295,N_4456,N_4210);
nor U5296 (N_5296,N_4825,N_4428);
nand U5297 (N_5297,N_4956,N_4902);
nor U5298 (N_5298,N_4652,N_4860);
and U5299 (N_5299,N_4176,N_4412);
nor U5300 (N_5300,N_4199,N_4219);
and U5301 (N_5301,N_4471,N_4239);
nor U5302 (N_5302,N_4580,N_4427);
and U5303 (N_5303,N_4822,N_4921);
nand U5304 (N_5304,N_4064,N_4182);
or U5305 (N_5305,N_4244,N_4933);
and U5306 (N_5306,N_4237,N_4516);
or U5307 (N_5307,N_4380,N_4590);
nand U5308 (N_5308,N_4589,N_4231);
nand U5309 (N_5309,N_4547,N_4230);
nor U5310 (N_5310,N_4841,N_4093);
nand U5311 (N_5311,N_4308,N_4983);
nand U5312 (N_5312,N_4924,N_4396);
or U5313 (N_5313,N_4993,N_4833);
nand U5314 (N_5314,N_4108,N_4505);
nand U5315 (N_5315,N_4631,N_4297);
nand U5316 (N_5316,N_4104,N_4582);
nor U5317 (N_5317,N_4209,N_4192);
and U5318 (N_5318,N_4685,N_4369);
nand U5319 (N_5319,N_4837,N_4134);
nand U5320 (N_5320,N_4467,N_4561);
nand U5321 (N_5321,N_4092,N_4019);
nand U5322 (N_5322,N_4286,N_4604);
nor U5323 (N_5323,N_4785,N_4999);
nand U5324 (N_5324,N_4150,N_4306);
nor U5325 (N_5325,N_4732,N_4783);
or U5326 (N_5326,N_4946,N_4483);
and U5327 (N_5327,N_4491,N_4402);
nor U5328 (N_5328,N_4663,N_4832);
or U5329 (N_5329,N_4932,N_4121);
or U5330 (N_5330,N_4526,N_4725);
nand U5331 (N_5331,N_4807,N_4954);
nand U5332 (N_5332,N_4938,N_4919);
and U5333 (N_5333,N_4878,N_4419);
nand U5334 (N_5334,N_4724,N_4205);
or U5335 (N_5335,N_4705,N_4951);
and U5336 (N_5336,N_4115,N_4278);
nand U5337 (N_5337,N_4890,N_4370);
or U5338 (N_5338,N_4984,N_4880);
and U5339 (N_5339,N_4460,N_4694);
nand U5340 (N_5340,N_4400,N_4442);
nor U5341 (N_5341,N_4974,N_4107);
or U5342 (N_5342,N_4276,N_4397);
or U5343 (N_5343,N_4367,N_4624);
nor U5344 (N_5344,N_4727,N_4610);
nand U5345 (N_5345,N_4506,N_4985);
or U5346 (N_5346,N_4218,N_4301);
nor U5347 (N_5347,N_4539,N_4067);
and U5348 (N_5348,N_4008,N_4752);
nor U5349 (N_5349,N_4187,N_4321);
nor U5350 (N_5350,N_4968,N_4011);
nor U5351 (N_5351,N_4391,N_4153);
nand U5352 (N_5352,N_4758,N_4234);
nand U5353 (N_5353,N_4757,N_4475);
nor U5354 (N_5354,N_4078,N_4009);
nor U5355 (N_5355,N_4021,N_4431);
or U5356 (N_5356,N_4712,N_4931);
or U5357 (N_5357,N_4057,N_4053);
and U5358 (N_5358,N_4789,N_4172);
nand U5359 (N_5359,N_4155,N_4485);
nand U5360 (N_5360,N_4001,N_4944);
or U5361 (N_5361,N_4310,N_4022);
nor U5362 (N_5362,N_4418,N_4232);
and U5363 (N_5363,N_4015,N_4365);
nor U5364 (N_5364,N_4096,N_4038);
nor U5365 (N_5365,N_4486,N_4254);
and U5366 (N_5366,N_4617,N_4133);
or U5367 (N_5367,N_4678,N_4846);
nor U5368 (N_5368,N_4085,N_4528);
nand U5369 (N_5369,N_4618,N_4323);
nor U5370 (N_5370,N_4048,N_4553);
nand U5371 (N_5371,N_4262,N_4719);
or U5372 (N_5372,N_4613,N_4768);
nand U5373 (N_5373,N_4087,N_4538);
nand U5374 (N_5374,N_4518,N_4844);
nor U5375 (N_5375,N_4387,N_4292);
xor U5376 (N_5376,N_4588,N_4395);
nand U5377 (N_5377,N_4071,N_4729);
or U5378 (N_5378,N_4507,N_4315);
and U5379 (N_5379,N_4908,N_4043);
or U5380 (N_5380,N_4113,N_4052);
nand U5381 (N_5381,N_4157,N_4200);
and U5382 (N_5382,N_4831,N_4407);
nand U5383 (N_5383,N_4423,N_4548);
nor U5384 (N_5384,N_4892,N_4394);
xnor U5385 (N_5385,N_4217,N_4345);
nand U5386 (N_5386,N_4339,N_4417);
nor U5387 (N_5387,N_4309,N_4512);
nand U5388 (N_5388,N_4942,N_4843);
or U5389 (N_5389,N_4258,N_4511);
nand U5390 (N_5390,N_4376,N_4742);
or U5391 (N_5391,N_4882,N_4893);
or U5392 (N_5392,N_4314,N_4362);
or U5393 (N_5393,N_4060,N_4058);
and U5394 (N_5394,N_4149,N_4578);
or U5395 (N_5395,N_4202,N_4379);
nor U5396 (N_5396,N_4171,N_4220);
and U5397 (N_5397,N_4953,N_4801);
or U5398 (N_5398,N_4099,N_4671);
nor U5399 (N_5399,N_4377,N_4619);
nand U5400 (N_5400,N_4393,N_4037);
nor U5401 (N_5401,N_4359,N_4111);
and U5402 (N_5402,N_4307,N_4503);
and U5403 (N_5403,N_4917,N_4451);
nor U5404 (N_5404,N_4703,N_4900);
and U5405 (N_5405,N_4079,N_4615);
and U5406 (N_5406,N_4988,N_4545);
or U5407 (N_5407,N_4277,N_4253);
nor U5408 (N_5408,N_4510,N_4500);
or U5409 (N_5409,N_4381,N_4565);
and U5410 (N_5410,N_4129,N_4374);
nor U5411 (N_5411,N_4433,N_4414);
nor U5412 (N_5412,N_4662,N_4894);
nand U5413 (N_5413,N_4594,N_4644);
nand U5414 (N_5414,N_4865,N_4497);
nor U5415 (N_5415,N_4776,N_4364);
and U5416 (N_5416,N_4327,N_4474);
and U5417 (N_5417,N_4119,N_4117);
or U5418 (N_5418,N_4036,N_4452);
xor U5419 (N_5419,N_4375,N_4821);
and U5420 (N_5420,N_4185,N_4706);
or U5421 (N_5421,N_4971,N_4796);
nor U5422 (N_5422,N_4495,N_4854);
nand U5423 (N_5423,N_4186,N_4602);
nand U5424 (N_5424,N_4490,N_4767);
nor U5425 (N_5425,N_4439,N_4421);
nand U5426 (N_5426,N_4728,N_4191);
and U5427 (N_5427,N_4360,N_4568);
nand U5428 (N_5428,N_4798,N_4372);
or U5429 (N_5429,N_4131,N_4466);
nor U5430 (N_5430,N_4875,N_4871);
or U5431 (N_5431,N_4204,N_4222);
nor U5432 (N_5432,N_4879,N_4720);
or U5433 (N_5433,N_4658,N_4794);
and U5434 (N_5434,N_4701,N_4640);
nor U5435 (N_5435,N_4826,N_4845);
or U5436 (N_5436,N_4062,N_4963);
nor U5437 (N_5437,N_4897,N_4351);
and U5438 (N_5438,N_4642,N_4904);
nand U5439 (N_5439,N_4302,N_4415);
and U5440 (N_5440,N_4881,N_4410);
and U5441 (N_5441,N_4646,N_4123);
nor U5442 (N_5442,N_4959,N_4025);
or U5443 (N_5443,N_4148,N_4166);
nand U5444 (N_5444,N_4158,N_4722);
or U5445 (N_5445,N_4605,N_4469);
or U5446 (N_5446,N_4682,N_4564);
or U5447 (N_5447,N_4502,N_4517);
nor U5448 (N_5448,N_4777,N_4070);
or U5449 (N_5449,N_4519,N_4587);
nand U5450 (N_5450,N_4761,N_4948);
or U5451 (N_5451,N_4793,N_4076);
nor U5452 (N_5452,N_4770,N_4635);
and U5453 (N_5453,N_4656,N_4285);
or U5454 (N_5454,N_4792,N_4160);
nor U5455 (N_5455,N_4818,N_4748);
or U5456 (N_5456,N_4524,N_4138);
nor U5457 (N_5457,N_4173,N_4557);
nand U5458 (N_5458,N_4542,N_4184);
or U5459 (N_5459,N_4089,N_4626);
nor U5460 (N_5460,N_4252,N_4664);
and U5461 (N_5461,N_4976,N_4827);
and U5462 (N_5462,N_4636,N_4574);
and U5463 (N_5463,N_4072,N_4055);
xnor U5464 (N_5464,N_4438,N_4885);
or U5465 (N_5465,N_4216,N_4898);
or U5466 (N_5466,N_4197,N_4188);
or U5467 (N_5467,N_4888,N_4026);
or U5468 (N_5468,N_4453,N_4918);
or U5469 (N_5469,N_4413,N_4791);
and U5470 (N_5470,N_4606,N_4746);
nand U5471 (N_5471,N_4102,N_4927);
or U5472 (N_5472,N_4167,N_4420);
nor U5473 (N_5473,N_4082,N_4532);
and U5474 (N_5474,N_4572,N_4007);
nor U5475 (N_5475,N_4056,N_4447);
and U5476 (N_5476,N_4255,N_4958);
or U5477 (N_5477,N_4751,N_4472);
and U5478 (N_5478,N_4168,N_4998);
or U5479 (N_5479,N_4294,N_4922);
nand U5480 (N_5480,N_4086,N_4389);
and U5481 (N_5481,N_4450,N_4823);
nand U5482 (N_5482,N_4764,N_4163);
nand U5483 (N_5483,N_4864,N_4877);
or U5484 (N_5484,N_4817,N_4063);
and U5485 (N_5485,N_4620,N_4650);
or U5486 (N_5486,N_4408,N_4494);
and U5487 (N_5487,N_4634,N_4912);
nor U5488 (N_5488,N_4103,N_4839);
nor U5489 (N_5489,N_4169,N_4282);
nor U5490 (N_5490,N_4508,N_4320);
xnor U5491 (N_5491,N_4562,N_4743);
nand U5492 (N_5492,N_4478,N_4975);
or U5493 (N_5493,N_4406,N_4689);
nor U5494 (N_5494,N_4110,N_4271);
nor U5495 (N_5495,N_4470,N_4812);
nor U5496 (N_5496,N_4849,N_4859);
or U5497 (N_5497,N_4981,N_4544);
or U5498 (N_5498,N_4356,N_4756);
nor U5499 (N_5499,N_4835,N_4675);
and U5500 (N_5500,N_4296,N_4795);
or U5501 (N_5501,N_4554,N_4286);
nand U5502 (N_5502,N_4676,N_4440);
and U5503 (N_5503,N_4548,N_4592);
nand U5504 (N_5504,N_4440,N_4871);
and U5505 (N_5505,N_4171,N_4531);
nand U5506 (N_5506,N_4464,N_4003);
nor U5507 (N_5507,N_4912,N_4647);
nand U5508 (N_5508,N_4967,N_4519);
nand U5509 (N_5509,N_4053,N_4244);
or U5510 (N_5510,N_4643,N_4576);
and U5511 (N_5511,N_4483,N_4570);
and U5512 (N_5512,N_4557,N_4071);
or U5513 (N_5513,N_4852,N_4998);
nand U5514 (N_5514,N_4826,N_4706);
or U5515 (N_5515,N_4983,N_4685);
and U5516 (N_5516,N_4338,N_4346);
nand U5517 (N_5517,N_4109,N_4211);
nand U5518 (N_5518,N_4915,N_4224);
nand U5519 (N_5519,N_4171,N_4281);
and U5520 (N_5520,N_4902,N_4060);
nand U5521 (N_5521,N_4504,N_4949);
nand U5522 (N_5522,N_4722,N_4032);
nor U5523 (N_5523,N_4417,N_4509);
nand U5524 (N_5524,N_4676,N_4633);
nor U5525 (N_5525,N_4563,N_4735);
nand U5526 (N_5526,N_4576,N_4502);
nor U5527 (N_5527,N_4786,N_4286);
nor U5528 (N_5528,N_4020,N_4743);
nor U5529 (N_5529,N_4861,N_4609);
nor U5530 (N_5530,N_4754,N_4625);
nor U5531 (N_5531,N_4663,N_4208);
nor U5532 (N_5532,N_4349,N_4695);
xor U5533 (N_5533,N_4747,N_4622);
nor U5534 (N_5534,N_4435,N_4303);
nand U5535 (N_5535,N_4980,N_4555);
or U5536 (N_5536,N_4207,N_4178);
nor U5537 (N_5537,N_4402,N_4692);
nor U5538 (N_5538,N_4424,N_4705);
xor U5539 (N_5539,N_4090,N_4064);
and U5540 (N_5540,N_4936,N_4729);
nand U5541 (N_5541,N_4709,N_4188);
or U5542 (N_5542,N_4409,N_4367);
and U5543 (N_5543,N_4170,N_4502);
nor U5544 (N_5544,N_4972,N_4577);
nand U5545 (N_5545,N_4963,N_4878);
and U5546 (N_5546,N_4452,N_4845);
or U5547 (N_5547,N_4103,N_4699);
or U5548 (N_5548,N_4638,N_4448);
nand U5549 (N_5549,N_4131,N_4005);
nand U5550 (N_5550,N_4087,N_4777);
nor U5551 (N_5551,N_4165,N_4127);
and U5552 (N_5552,N_4334,N_4039);
or U5553 (N_5553,N_4700,N_4481);
nor U5554 (N_5554,N_4555,N_4801);
nor U5555 (N_5555,N_4543,N_4773);
or U5556 (N_5556,N_4415,N_4082);
and U5557 (N_5557,N_4128,N_4534);
or U5558 (N_5558,N_4646,N_4199);
nand U5559 (N_5559,N_4312,N_4160);
and U5560 (N_5560,N_4864,N_4384);
or U5561 (N_5561,N_4463,N_4320);
nor U5562 (N_5562,N_4108,N_4423);
nand U5563 (N_5563,N_4249,N_4453);
nand U5564 (N_5564,N_4430,N_4103);
and U5565 (N_5565,N_4529,N_4113);
and U5566 (N_5566,N_4467,N_4672);
and U5567 (N_5567,N_4922,N_4843);
nand U5568 (N_5568,N_4831,N_4413);
and U5569 (N_5569,N_4325,N_4973);
nand U5570 (N_5570,N_4940,N_4890);
nand U5571 (N_5571,N_4203,N_4276);
nand U5572 (N_5572,N_4602,N_4446);
and U5573 (N_5573,N_4187,N_4603);
or U5574 (N_5574,N_4495,N_4974);
and U5575 (N_5575,N_4099,N_4387);
xnor U5576 (N_5576,N_4187,N_4954);
and U5577 (N_5577,N_4127,N_4465);
nor U5578 (N_5578,N_4026,N_4917);
nand U5579 (N_5579,N_4695,N_4363);
or U5580 (N_5580,N_4503,N_4572);
nand U5581 (N_5581,N_4796,N_4738);
nor U5582 (N_5582,N_4315,N_4465);
xor U5583 (N_5583,N_4379,N_4041);
nor U5584 (N_5584,N_4756,N_4777);
nand U5585 (N_5585,N_4478,N_4706);
nand U5586 (N_5586,N_4412,N_4046);
and U5587 (N_5587,N_4210,N_4375);
nor U5588 (N_5588,N_4890,N_4257);
nand U5589 (N_5589,N_4667,N_4138);
and U5590 (N_5590,N_4114,N_4250);
nand U5591 (N_5591,N_4254,N_4627);
nand U5592 (N_5592,N_4585,N_4738);
nor U5593 (N_5593,N_4309,N_4794);
or U5594 (N_5594,N_4907,N_4657);
and U5595 (N_5595,N_4012,N_4892);
and U5596 (N_5596,N_4893,N_4045);
or U5597 (N_5597,N_4642,N_4707);
nor U5598 (N_5598,N_4392,N_4218);
and U5599 (N_5599,N_4453,N_4783);
or U5600 (N_5600,N_4516,N_4578);
or U5601 (N_5601,N_4508,N_4866);
nand U5602 (N_5602,N_4672,N_4420);
or U5603 (N_5603,N_4601,N_4588);
nor U5604 (N_5604,N_4261,N_4763);
and U5605 (N_5605,N_4923,N_4437);
or U5606 (N_5606,N_4508,N_4755);
nor U5607 (N_5607,N_4966,N_4511);
or U5608 (N_5608,N_4606,N_4602);
and U5609 (N_5609,N_4563,N_4656);
nor U5610 (N_5610,N_4739,N_4800);
or U5611 (N_5611,N_4036,N_4908);
or U5612 (N_5612,N_4261,N_4206);
and U5613 (N_5613,N_4344,N_4558);
nor U5614 (N_5614,N_4614,N_4104);
and U5615 (N_5615,N_4842,N_4555);
nor U5616 (N_5616,N_4208,N_4558);
nand U5617 (N_5617,N_4393,N_4294);
nor U5618 (N_5618,N_4269,N_4042);
nand U5619 (N_5619,N_4022,N_4552);
and U5620 (N_5620,N_4781,N_4196);
and U5621 (N_5621,N_4108,N_4486);
nor U5622 (N_5622,N_4367,N_4557);
or U5623 (N_5623,N_4919,N_4490);
nor U5624 (N_5624,N_4369,N_4482);
nor U5625 (N_5625,N_4698,N_4826);
and U5626 (N_5626,N_4567,N_4353);
nand U5627 (N_5627,N_4521,N_4861);
nor U5628 (N_5628,N_4597,N_4766);
or U5629 (N_5629,N_4921,N_4878);
and U5630 (N_5630,N_4648,N_4523);
or U5631 (N_5631,N_4827,N_4178);
nor U5632 (N_5632,N_4962,N_4498);
and U5633 (N_5633,N_4415,N_4057);
or U5634 (N_5634,N_4166,N_4180);
nor U5635 (N_5635,N_4774,N_4988);
and U5636 (N_5636,N_4547,N_4813);
or U5637 (N_5637,N_4752,N_4445);
nand U5638 (N_5638,N_4787,N_4564);
and U5639 (N_5639,N_4211,N_4765);
or U5640 (N_5640,N_4831,N_4972);
xnor U5641 (N_5641,N_4192,N_4831);
nand U5642 (N_5642,N_4326,N_4108);
or U5643 (N_5643,N_4677,N_4647);
or U5644 (N_5644,N_4959,N_4143);
nor U5645 (N_5645,N_4172,N_4683);
nor U5646 (N_5646,N_4802,N_4851);
and U5647 (N_5647,N_4141,N_4230);
or U5648 (N_5648,N_4258,N_4177);
nor U5649 (N_5649,N_4583,N_4113);
nor U5650 (N_5650,N_4745,N_4924);
and U5651 (N_5651,N_4219,N_4419);
or U5652 (N_5652,N_4969,N_4840);
and U5653 (N_5653,N_4928,N_4647);
and U5654 (N_5654,N_4070,N_4521);
nand U5655 (N_5655,N_4642,N_4150);
and U5656 (N_5656,N_4596,N_4549);
and U5657 (N_5657,N_4992,N_4840);
or U5658 (N_5658,N_4966,N_4903);
or U5659 (N_5659,N_4377,N_4086);
nand U5660 (N_5660,N_4771,N_4594);
nand U5661 (N_5661,N_4966,N_4420);
or U5662 (N_5662,N_4544,N_4731);
nor U5663 (N_5663,N_4423,N_4709);
nand U5664 (N_5664,N_4631,N_4273);
and U5665 (N_5665,N_4237,N_4762);
or U5666 (N_5666,N_4500,N_4923);
or U5667 (N_5667,N_4058,N_4975);
and U5668 (N_5668,N_4297,N_4250);
nor U5669 (N_5669,N_4100,N_4185);
nand U5670 (N_5670,N_4658,N_4292);
or U5671 (N_5671,N_4808,N_4459);
or U5672 (N_5672,N_4614,N_4966);
nor U5673 (N_5673,N_4352,N_4550);
or U5674 (N_5674,N_4706,N_4722);
nor U5675 (N_5675,N_4641,N_4983);
nand U5676 (N_5676,N_4990,N_4348);
or U5677 (N_5677,N_4824,N_4506);
nor U5678 (N_5678,N_4538,N_4129);
nand U5679 (N_5679,N_4667,N_4832);
and U5680 (N_5680,N_4980,N_4234);
nand U5681 (N_5681,N_4125,N_4839);
nand U5682 (N_5682,N_4296,N_4124);
nand U5683 (N_5683,N_4517,N_4060);
nand U5684 (N_5684,N_4086,N_4935);
and U5685 (N_5685,N_4257,N_4983);
xnor U5686 (N_5686,N_4789,N_4553);
nor U5687 (N_5687,N_4181,N_4927);
nor U5688 (N_5688,N_4068,N_4921);
or U5689 (N_5689,N_4891,N_4769);
or U5690 (N_5690,N_4544,N_4267);
nand U5691 (N_5691,N_4992,N_4741);
nor U5692 (N_5692,N_4581,N_4217);
or U5693 (N_5693,N_4172,N_4294);
and U5694 (N_5694,N_4896,N_4349);
or U5695 (N_5695,N_4458,N_4687);
nand U5696 (N_5696,N_4407,N_4122);
nand U5697 (N_5697,N_4778,N_4176);
or U5698 (N_5698,N_4817,N_4013);
or U5699 (N_5699,N_4606,N_4642);
or U5700 (N_5700,N_4120,N_4473);
and U5701 (N_5701,N_4054,N_4656);
or U5702 (N_5702,N_4987,N_4274);
nand U5703 (N_5703,N_4106,N_4050);
nand U5704 (N_5704,N_4387,N_4261);
or U5705 (N_5705,N_4104,N_4434);
or U5706 (N_5706,N_4044,N_4257);
or U5707 (N_5707,N_4248,N_4425);
nand U5708 (N_5708,N_4006,N_4840);
nor U5709 (N_5709,N_4857,N_4221);
nand U5710 (N_5710,N_4727,N_4261);
nor U5711 (N_5711,N_4000,N_4437);
or U5712 (N_5712,N_4086,N_4100);
and U5713 (N_5713,N_4761,N_4774);
nor U5714 (N_5714,N_4963,N_4234);
nor U5715 (N_5715,N_4108,N_4475);
nor U5716 (N_5716,N_4453,N_4923);
nand U5717 (N_5717,N_4691,N_4217);
nor U5718 (N_5718,N_4694,N_4353);
nand U5719 (N_5719,N_4675,N_4580);
nor U5720 (N_5720,N_4187,N_4791);
and U5721 (N_5721,N_4114,N_4157);
or U5722 (N_5722,N_4702,N_4384);
or U5723 (N_5723,N_4283,N_4618);
nor U5724 (N_5724,N_4725,N_4603);
nand U5725 (N_5725,N_4381,N_4733);
or U5726 (N_5726,N_4710,N_4890);
nand U5727 (N_5727,N_4269,N_4884);
and U5728 (N_5728,N_4319,N_4860);
or U5729 (N_5729,N_4686,N_4409);
and U5730 (N_5730,N_4176,N_4720);
and U5731 (N_5731,N_4991,N_4662);
nand U5732 (N_5732,N_4559,N_4192);
and U5733 (N_5733,N_4367,N_4075);
and U5734 (N_5734,N_4692,N_4897);
and U5735 (N_5735,N_4743,N_4454);
and U5736 (N_5736,N_4944,N_4278);
or U5737 (N_5737,N_4478,N_4851);
nor U5738 (N_5738,N_4758,N_4221);
or U5739 (N_5739,N_4864,N_4953);
nor U5740 (N_5740,N_4987,N_4167);
and U5741 (N_5741,N_4511,N_4093);
or U5742 (N_5742,N_4522,N_4111);
nor U5743 (N_5743,N_4849,N_4722);
nor U5744 (N_5744,N_4646,N_4826);
nor U5745 (N_5745,N_4650,N_4420);
nand U5746 (N_5746,N_4309,N_4361);
or U5747 (N_5747,N_4169,N_4291);
or U5748 (N_5748,N_4252,N_4374);
or U5749 (N_5749,N_4500,N_4005);
nor U5750 (N_5750,N_4442,N_4882);
nand U5751 (N_5751,N_4177,N_4712);
or U5752 (N_5752,N_4493,N_4085);
or U5753 (N_5753,N_4899,N_4544);
and U5754 (N_5754,N_4489,N_4622);
nand U5755 (N_5755,N_4466,N_4092);
and U5756 (N_5756,N_4544,N_4790);
nor U5757 (N_5757,N_4398,N_4505);
or U5758 (N_5758,N_4358,N_4356);
nand U5759 (N_5759,N_4800,N_4514);
or U5760 (N_5760,N_4039,N_4923);
or U5761 (N_5761,N_4409,N_4378);
and U5762 (N_5762,N_4486,N_4034);
and U5763 (N_5763,N_4476,N_4654);
nor U5764 (N_5764,N_4144,N_4959);
nand U5765 (N_5765,N_4542,N_4894);
nand U5766 (N_5766,N_4656,N_4730);
nand U5767 (N_5767,N_4686,N_4933);
or U5768 (N_5768,N_4417,N_4066);
nand U5769 (N_5769,N_4027,N_4582);
and U5770 (N_5770,N_4343,N_4518);
nand U5771 (N_5771,N_4180,N_4834);
nor U5772 (N_5772,N_4189,N_4631);
and U5773 (N_5773,N_4064,N_4660);
nor U5774 (N_5774,N_4302,N_4372);
or U5775 (N_5775,N_4909,N_4690);
nand U5776 (N_5776,N_4563,N_4655);
or U5777 (N_5777,N_4347,N_4536);
nor U5778 (N_5778,N_4100,N_4289);
nand U5779 (N_5779,N_4677,N_4891);
and U5780 (N_5780,N_4999,N_4680);
and U5781 (N_5781,N_4199,N_4084);
and U5782 (N_5782,N_4201,N_4681);
and U5783 (N_5783,N_4644,N_4077);
and U5784 (N_5784,N_4254,N_4313);
and U5785 (N_5785,N_4068,N_4976);
and U5786 (N_5786,N_4067,N_4208);
nor U5787 (N_5787,N_4635,N_4605);
nand U5788 (N_5788,N_4313,N_4781);
nand U5789 (N_5789,N_4705,N_4316);
and U5790 (N_5790,N_4415,N_4996);
nor U5791 (N_5791,N_4549,N_4947);
or U5792 (N_5792,N_4810,N_4851);
and U5793 (N_5793,N_4083,N_4672);
or U5794 (N_5794,N_4990,N_4708);
nand U5795 (N_5795,N_4729,N_4031);
and U5796 (N_5796,N_4900,N_4447);
nor U5797 (N_5797,N_4430,N_4931);
or U5798 (N_5798,N_4223,N_4452);
nor U5799 (N_5799,N_4008,N_4634);
or U5800 (N_5800,N_4650,N_4802);
or U5801 (N_5801,N_4917,N_4123);
xnor U5802 (N_5802,N_4259,N_4458);
nand U5803 (N_5803,N_4538,N_4165);
nor U5804 (N_5804,N_4413,N_4368);
nor U5805 (N_5805,N_4389,N_4026);
nor U5806 (N_5806,N_4892,N_4601);
or U5807 (N_5807,N_4800,N_4505);
nand U5808 (N_5808,N_4960,N_4845);
and U5809 (N_5809,N_4592,N_4237);
nand U5810 (N_5810,N_4291,N_4621);
and U5811 (N_5811,N_4037,N_4099);
nand U5812 (N_5812,N_4431,N_4964);
and U5813 (N_5813,N_4354,N_4127);
nor U5814 (N_5814,N_4899,N_4342);
nor U5815 (N_5815,N_4485,N_4255);
or U5816 (N_5816,N_4352,N_4072);
and U5817 (N_5817,N_4088,N_4355);
and U5818 (N_5818,N_4307,N_4538);
and U5819 (N_5819,N_4608,N_4801);
or U5820 (N_5820,N_4366,N_4748);
nor U5821 (N_5821,N_4138,N_4367);
or U5822 (N_5822,N_4586,N_4839);
or U5823 (N_5823,N_4126,N_4152);
or U5824 (N_5824,N_4290,N_4818);
or U5825 (N_5825,N_4854,N_4983);
and U5826 (N_5826,N_4492,N_4691);
and U5827 (N_5827,N_4273,N_4025);
nor U5828 (N_5828,N_4647,N_4558);
nor U5829 (N_5829,N_4948,N_4705);
or U5830 (N_5830,N_4010,N_4219);
or U5831 (N_5831,N_4633,N_4700);
or U5832 (N_5832,N_4442,N_4137);
nand U5833 (N_5833,N_4292,N_4319);
nand U5834 (N_5834,N_4715,N_4619);
xor U5835 (N_5835,N_4199,N_4800);
nor U5836 (N_5836,N_4291,N_4753);
nor U5837 (N_5837,N_4735,N_4276);
and U5838 (N_5838,N_4599,N_4735);
nor U5839 (N_5839,N_4355,N_4705);
nand U5840 (N_5840,N_4676,N_4981);
nor U5841 (N_5841,N_4755,N_4765);
and U5842 (N_5842,N_4723,N_4525);
or U5843 (N_5843,N_4670,N_4624);
xor U5844 (N_5844,N_4378,N_4281);
and U5845 (N_5845,N_4577,N_4824);
nor U5846 (N_5846,N_4246,N_4860);
nand U5847 (N_5847,N_4095,N_4106);
nor U5848 (N_5848,N_4740,N_4839);
or U5849 (N_5849,N_4433,N_4131);
or U5850 (N_5850,N_4734,N_4916);
or U5851 (N_5851,N_4982,N_4762);
and U5852 (N_5852,N_4165,N_4734);
nand U5853 (N_5853,N_4564,N_4099);
nand U5854 (N_5854,N_4430,N_4615);
or U5855 (N_5855,N_4312,N_4148);
nor U5856 (N_5856,N_4225,N_4204);
and U5857 (N_5857,N_4923,N_4166);
nor U5858 (N_5858,N_4041,N_4735);
and U5859 (N_5859,N_4084,N_4119);
nand U5860 (N_5860,N_4696,N_4391);
nand U5861 (N_5861,N_4243,N_4918);
nor U5862 (N_5862,N_4396,N_4691);
or U5863 (N_5863,N_4209,N_4563);
nor U5864 (N_5864,N_4520,N_4020);
nand U5865 (N_5865,N_4315,N_4250);
or U5866 (N_5866,N_4699,N_4812);
or U5867 (N_5867,N_4470,N_4492);
and U5868 (N_5868,N_4130,N_4398);
nand U5869 (N_5869,N_4619,N_4456);
or U5870 (N_5870,N_4322,N_4918);
nor U5871 (N_5871,N_4928,N_4618);
or U5872 (N_5872,N_4690,N_4973);
nand U5873 (N_5873,N_4686,N_4763);
nand U5874 (N_5874,N_4458,N_4497);
nand U5875 (N_5875,N_4692,N_4258);
xor U5876 (N_5876,N_4171,N_4427);
and U5877 (N_5877,N_4690,N_4376);
or U5878 (N_5878,N_4689,N_4988);
nor U5879 (N_5879,N_4345,N_4105);
nand U5880 (N_5880,N_4772,N_4577);
nor U5881 (N_5881,N_4427,N_4918);
nor U5882 (N_5882,N_4940,N_4041);
nor U5883 (N_5883,N_4442,N_4033);
or U5884 (N_5884,N_4139,N_4748);
nor U5885 (N_5885,N_4142,N_4948);
or U5886 (N_5886,N_4416,N_4411);
nor U5887 (N_5887,N_4932,N_4815);
or U5888 (N_5888,N_4874,N_4248);
nor U5889 (N_5889,N_4091,N_4967);
nand U5890 (N_5890,N_4290,N_4130);
and U5891 (N_5891,N_4304,N_4565);
and U5892 (N_5892,N_4412,N_4818);
or U5893 (N_5893,N_4955,N_4333);
nand U5894 (N_5894,N_4669,N_4541);
xnor U5895 (N_5895,N_4696,N_4331);
nand U5896 (N_5896,N_4283,N_4030);
or U5897 (N_5897,N_4918,N_4966);
xor U5898 (N_5898,N_4535,N_4515);
nand U5899 (N_5899,N_4705,N_4695);
and U5900 (N_5900,N_4343,N_4407);
nor U5901 (N_5901,N_4559,N_4137);
and U5902 (N_5902,N_4557,N_4616);
and U5903 (N_5903,N_4865,N_4092);
nor U5904 (N_5904,N_4507,N_4461);
nand U5905 (N_5905,N_4082,N_4203);
nor U5906 (N_5906,N_4479,N_4725);
and U5907 (N_5907,N_4704,N_4138);
and U5908 (N_5908,N_4877,N_4569);
and U5909 (N_5909,N_4146,N_4002);
or U5910 (N_5910,N_4559,N_4873);
nor U5911 (N_5911,N_4080,N_4154);
and U5912 (N_5912,N_4922,N_4551);
nor U5913 (N_5913,N_4505,N_4328);
or U5914 (N_5914,N_4839,N_4811);
and U5915 (N_5915,N_4575,N_4834);
nand U5916 (N_5916,N_4953,N_4193);
nand U5917 (N_5917,N_4281,N_4804);
nor U5918 (N_5918,N_4165,N_4272);
nand U5919 (N_5919,N_4015,N_4076);
and U5920 (N_5920,N_4006,N_4808);
or U5921 (N_5921,N_4689,N_4938);
nor U5922 (N_5922,N_4003,N_4173);
and U5923 (N_5923,N_4089,N_4198);
and U5924 (N_5924,N_4468,N_4576);
nand U5925 (N_5925,N_4712,N_4885);
and U5926 (N_5926,N_4388,N_4835);
nand U5927 (N_5927,N_4293,N_4117);
and U5928 (N_5928,N_4045,N_4317);
or U5929 (N_5929,N_4918,N_4003);
and U5930 (N_5930,N_4100,N_4283);
or U5931 (N_5931,N_4455,N_4745);
or U5932 (N_5932,N_4572,N_4462);
or U5933 (N_5933,N_4435,N_4515);
nand U5934 (N_5934,N_4851,N_4593);
or U5935 (N_5935,N_4071,N_4849);
nand U5936 (N_5936,N_4751,N_4256);
nor U5937 (N_5937,N_4703,N_4638);
and U5938 (N_5938,N_4579,N_4174);
and U5939 (N_5939,N_4784,N_4380);
or U5940 (N_5940,N_4410,N_4087);
and U5941 (N_5941,N_4373,N_4009);
xor U5942 (N_5942,N_4020,N_4425);
and U5943 (N_5943,N_4020,N_4490);
nand U5944 (N_5944,N_4017,N_4361);
or U5945 (N_5945,N_4006,N_4559);
nand U5946 (N_5946,N_4395,N_4753);
nor U5947 (N_5947,N_4859,N_4963);
or U5948 (N_5948,N_4944,N_4581);
nor U5949 (N_5949,N_4065,N_4230);
nor U5950 (N_5950,N_4106,N_4962);
nor U5951 (N_5951,N_4729,N_4233);
nor U5952 (N_5952,N_4211,N_4700);
nor U5953 (N_5953,N_4251,N_4022);
nor U5954 (N_5954,N_4554,N_4173);
or U5955 (N_5955,N_4797,N_4883);
nor U5956 (N_5956,N_4059,N_4886);
and U5957 (N_5957,N_4512,N_4838);
or U5958 (N_5958,N_4785,N_4290);
nand U5959 (N_5959,N_4141,N_4972);
and U5960 (N_5960,N_4439,N_4332);
nand U5961 (N_5961,N_4189,N_4456);
and U5962 (N_5962,N_4060,N_4003);
nand U5963 (N_5963,N_4712,N_4799);
or U5964 (N_5964,N_4061,N_4128);
nor U5965 (N_5965,N_4988,N_4328);
nor U5966 (N_5966,N_4832,N_4868);
and U5967 (N_5967,N_4897,N_4903);
nor U5968 (N_5968,N_4797,N_4300);
and U5969 (N_5969,N_4444,N_4234);
or U5970 (N_5970,N_4442,N_4046);
and U5971 (N_5971,N_4541,N_4312);
nand U5972 (N_5972,N_4227,N_4511);
and U5973 (N_5973,N_4162,N_4460);
and U5974 (N_5974,N_4667,N_4562);
nand U5975 (N_5975,N_4962,N_4006);
nand U5976 (N_5976,N_4097,N_4162);
nand U5977 (N_5977,N_4981,N_4872);
or U5978 (N_5978,N_4999,N_4282);
and U5979 (N_5979,N_4913,N_4886);
nor U5980 (N_5980,N_4054,N_4017);
nand U5981 (N_5981,N_4427,N_4114);
nand U5982 (N_5982,N_4390,N_4500);
nor U5983 (N_5983,N_4820,N_4883);
and U5984 (N_5984,N_4829,N_4615);
nor U5985 (N_5985,N_4227,N_4005);
nand U5986 (N_5986,N_4244,N_4361);
or U5987 (N_5987,N_4231,N_4338);
nand U5988 (N_5988,N_4639,N_4237);
nor U5989 (N_5989,N_4398,N_4965);
nor U5990 (N_5990,N_4118,N_4833);
nor U5991 (N_5991,N_4892,N_4757);
or U5992 (N_5992,N_4235,N_4056);
nand U5993 (N_5993,N_4068,N_4430);
nand U5994 (N_5994,N_4096,N_4567);
nand U5995 (N_5995,N_4904,N_4546);
nor U5996 (N_5996,N_4200,N_4775);
or U5997 (N_5997,N_4993,N_4161);
nand U5998 (N_5998,N_4059,N_4265);
xnor U5999 (N_5999,N_4956,N_4769);
and U6000 (N_6000,N_5231,N_5697);
nand U6001 (N_6001,N_5308,N_5781);
and U6002 (N_6002,N_5803,N_5069);
nand U6003 (N_6003,N_5336,N_5515);
nand U6004 (N_6004,N_5162,N_5153);
and U6005 (N_6005,N_5199,N_5679);
nand U6006 (N_6006,N_5943,N_5648);
or U6007 (N_6007,N_5433,N_5120);
nor U6008 (N_6008,N_5259,N_5823);
nand U6009 (N_6009,N_5414,N_5819);
nand U6010 (N_6010,N_5317,N_5569);
nor U6011 (N_6011,N_5953,N_5845);
nand U6012 (N_6012,N_5022,N_5482);
nor U6013 (N_6013,N_5493,N_5264);
or U6014 (N_6014,N_5738,N_5502);
and U6015 (N_6015,N_5028,N_5649);
or U6016 (N_6016,N_5665,N_5533);
or U6017 (N_6017,N_5034,N_5172);
and U6018 (N_6018,N_5391,N_5088);
nor U6019 (N_6019,N_5454,N_5423);
nor U6020 (N_6020,N_5689,N_5480);
or U6021 (N_6021,N_5239,N_5927);
and U6022 (N_6022,N_5990,N_5353);
or U6023 (N_6023,N_5019,N_5381);
and U6024 (N_6024,N_5211,N_5776);
nand U6025 (N_6025,N_5835,N_5914);
nand U6026 (N_6026,N_5384,N_5411);
nand U6027 (N_6027,N_5624,N_5327);
nand U6028 (N_6028,N_5002,N_5179);
nand U6029 (N_6029,N_5437,N_5464);
nor U6030 (N_6030,N_5106,N_5169);
and U6031 (N_6031,N_5071,N_5006);
or U6032 (N_6032,N_5673,N_5097);
or U6033 (N_6033,N_5770,N_5060);
or U6034 (N_6034,N_5444,N_5431);
or U6035 (N_6035,N_5969,N_5559);
or U6036 (N_6036,N_5813,N_5677);
nor U6037 (N_6037,N_5042,N_5198);
nor U6038 (N_6038,N_5050,N_5903);
nor U6039 (N_6039,N_5175,N_5012);
or U6040 (N_6040,N_5495,N_5562);
nand U6041 (N_6041,N_5950,N_5589);
nand U6042 (N_6042,N_5843,N_5100);
and U6043 (N_6043,N_5426,N_5832);
or U6044 (N_6044,N_5152,N_5430);
or U6045 (N_6045,N_5500,N_5509);
or U6046 (N_6046,N_5385,N_5070);
nand U6047 (N_6047,N_5834,N_5200);
nand U6048 (N_6048,N_5185,N_5829);
nor U6049 (N_6049,N_5349,N_5514);
nand U6050 (N_6050,N_5955,N_5506);
and U6051 (N_6051,N_5429,N_5145);
and U6052 (N_6052,N_5268,N_5292);
nand U6053 (N_6053,N_5314,N_5485);
nor U6054 (N_6054,N_5432,N_5084);
nand U6055 (N_6055,N_5147,N_5761);
or U6056 (N_6056,N_5475,N_5144);
nand U6057 (N_6057,N_5379,N_5068);
nor U6058 (N_6058,N_5644,N_5357);
nand U6059 (N_6059,N_5702,N_5688);
or U6060 (N_6060,N_5610,N_5261);
or U6061 (N_6061,N_5396,N_5399);
or U6062 (N_6062,N_5092,N_5960);
and U6063 (N_6063,N_5858,N_5743);
or U6064 (N_6064,N_5039,N_5057);
nor U6065 (N_6065,N_5089,N_5224);
and U6066 (N_6066,N_5365,N_5300);
nand U6067 (N_6067,N_5944,N_5220);
nand U6068 (N_6068,N_5635,N_5575);
nand U6069 (N_6069,N_5170,N_5346);
and U6070 (N_6070,N_5664,N_5730);
nor U6071 (N_6071,N_5894,N_5510);
nand U6072 (N_6072,N_5877,N_5310);
or U6073 (N_6073,N_5904,N_5208);
or U6074 (N_6074,N_5983,N_5612);
nor U6075 (N_6075,N_5301,N_5272);
and U6076 (N_6076,N_5837,N_5724);
nor U6077 (N_6077,N_5529,N_5866);
nand U6078 (N_6078,N_5109,N_5230);
or U6079 (N_6079,N_5585,N_5735);
nand U6080 (N_6080,N_5271,N_5187);
nor U6081 (N_6081,N_5893,N_5979);
nand U6082 (N_6082,N_5263,N_5658);
nor U6083 (N_6083,N_5755,N_5104);
xor U6084 (N_6084,N_5784,N_5795);
and U6085 (N_6085,N_5322,N_5691);
nor U6086 (N_6086,N_5283,N_5001);
nor U6087 (N_6087,N_5815,N_5099);
nand U6088 (N_6088,N_5958,N_5841);
nand U6089 (N_6089,N_5974,N_5872);
nand U6090 (N_6090,N_5094,N_5407);
xnor U6091 (N_6091,N_5328,N_5519);
nor U6092 (N_6092,N_5377,N_5151);
nor U6093 (N_6093,N_5478,N_5672);
and U6094 (N_6094,N_5465,N_5289);
or U6095 (N_6095,N_5463,N_5551);
nor U6096 (N_6096,N_5363,N_5132);
and U6097 (N_6097,N_5698,N_5476);
and U6098 (N_6098,N_5256,N_5458);
nor U6099 (N_6099,N_5507,N_5687);
nor U6100 (N_6100,N_5825,N_5809);
nand U6101 (N_6101,N_5098,N_5274);
and U6102 (N_6102,N_5532,N_5371);
and U6103 (N_6103,N_5078,N_5453);
nand U6104 (N_6104,N_5930,N_5362);
nand U6105 (N_6105,N_5382,N_5055);
or U6106 (N_6106,N_5622,N_5018);
and U6107 (N_6107,N_5721,N_5748);
and U6108 (N_6108,N_5949,N_5330);
and U6109 (N_6109,N_5269,N_5184);
nor U6110 (N_6110,N_5709,N_5549);
nand U6111 (N_6111,N_5294,N_5650);
or U6112 (N_6112,N_5400,N_5545);
nand U6113 (N_6113,N_5621,N_5202);
and U6114 (N_6114,N_5758,N_5354);
xnor U6115 (N_6115,N_5530,N_5600);
or U6116 (N_6116,N_5626,N_5150);
and U6117 (N_6117,N_5970,N_5544);
and U6118 (N_6118,N_5847,N_5339);
nand U6119 (N_6119,N_5865,N_5981);
or U6120 (N_6120,N_5752,N_5686);
and U6121 (N_6121,N_5293,N_5277);
and U6122 (N_6122,N_5867,N_5996);
nand U6123 (N_6123,N_5547,N_5871);
and U6124 (N_6124,N_5217,N_5262);
nor U6125 (N_6125,N_5237,N_5690);
nor U6126 (N_6126,N_5766,N_5616);
or U6127 (N_6127,N_5275,N_5338);
and U6128 (N_6128,N_5810,N_5772);
and U6129 (N_6129,N_5410,N_5557);
nand U6130 (N_6130,N_5991,N_5986);
nand U6131 (N_6131,N_5728,N_5309);
and U6132 (N_6132,N_5555,N_5014);
nand U6133 (N_6133,N_5731,N_5820);
nor U6134 (N_6134,N_5675,N_5049);
or U6135 (N_6135,N_5483,N_5613);
nand U6136 (N_6136,N_5773,N_5148);
nor U6137 (N_6137,N_5488,N_5937);
or U6138 (N_6138,N_5251,N_5787);
and U6139 (N_6139,N_5074,N_5938);
and U6140 (N_6140,N_5403,N_5143);
and U6141 (N_6141,N_5062,N_5242);
or U6142 (N_6142,N_5606,N_5802);
xnor U6143 (N_6143,N_5503,N_5248);
nand U6144 (N_6144,N_5467,N_5750);
nand U6145 (N_6145,N_5628,N_5064);
nor U6146 (N_6146,N_5358,N_5707);
or U6147 (N_6147,N_5124,N_5838);
nor U6148 (N_6148,N_5901,N_5887);
and U6149 (N_6149,N_5594,N_5494);
nor U6150 (N_6150,N_5121,N_5449);
and U6151 (N_6151,N_5025,N_5692);
and U6152 (N_6152,N_5597,N_5405);
nand U6153 (N_6153,N_5003,N_5421);
and U6154 (N_6154,N_5550,N_5997);
and U6155 (N_6155,N_5527,N_5189);
nand U6156 (N_6156,N_5993,N_5971);
nand U6157 (N_6157,N_5722,N_5817);
or U6158 (N_6158,N_5246,N_5674);
nand U6159 (N_6159,N_5980,N_5469);
and U6160 (N_6160,N_5737,N_5190);
or U6161 (N_6161,N_5791,N_5627);
and U6162 (N_6162,N_5222,N_5374);
nor U6163 (N_6163,N_5701,N_5215);
or U6164 (N_6164,N_5020,N_5900);
or U6165 (N_6165,N_5554,N_5592);
xnor U6166 (N_6166,N_5298,N_5048);
and U6167 (N_6167,N_5576,N_5040);
and U6168 (N_6168,N_5563,N_5956);
or U6169 (N_6169,N_5951,N_5361);
nor U6170 (N_6170,N_5178,N_5862);
and U6171 (N_6171,N_5741,N_5140);
and U6172 (N_6172,N_5704,N_5523);
or U6173 (N_6173,N_5061,N_5171);
nand U6174 (N_6174,N_5219,N_5366);
or U6175 (N_6175,N_5149,N_5636);
nand U6176 (N_6176,N_5933,N_5499);
and U6177 (N_6177,N_5378,N_5605);
and U6178 (N_6178,N_5935,N_5114);
nor U6179 (N_6179,N_5204,N_5305);
or U6180 (N_6180,N_5270,N_5964);
nor U6181 (N_6181,N_5646,N_5236);
and U6182 (N_6182,N_5513,N_5888);
or U6183 (N_6183,N_5553,N_5343);
nor U6184 (N_6184,N_5266,N_5528);
or U6185 (N_6185,N_5718,N_5978);
and U6186 (N_6186,N_5440,N_5004);
and U6187 (N_6187,N_5032,N_5645);
or U6188 (N_6188,N_5824,N_5041);
and U6189 (N_6189,N_5418,N_5870);
and U6190 (N_6190,N_5534,N_5136);
nor U6191 (N_6191,N_5319,N_5678);
and U6192 (N_6192,N_5988,N_5214);
and U6193 (N_6193,N_5356,N_5355);
nand U6194 (N_6194,N_5233,N_5693);
nor U6195 (N_6195,N_5936,N_5180);
nand U6196 (N_6196,N_5046,N_5586);
nor U6197 (N_6197,N_5985,N_5801);
or U6198 (N_6198,N_5110,N_5921);
nor U6199 (N_6199,N_5695,N_5827);
nand U6200 (N_6200,N_5183,N_5769);
and U6201 (N_6201,N_5130,N_5705);
nand U6202 (N_6202,N_5525,N_5762);
nor U6203 (N_6203,N_5267,N_5734);
nor U6204 (N_6204,N_5751,N_5116);
nor U6205 (N_6205,N_5158,N_5299);
nor U6206 (N_6206,N_5924,N_5987);
and U6207 (N_6207,N_5512,N_5736);
nand U6208 (N_6208,N_5670,N_5347);
nor U6209 (N_6209,N_5367,N_5254);
or U6210 (N_6210,N_5497,N_5915);
nor U6211 (N_6211,N_5380,N_5203);
nand U6212 (N_6212,N_5853,N_5614);
nand U6213 (N_6213,N_5588,N_5386);
and U6214 (N_6214,N_5126,N_5455);
xor U6215 (N_6215,N_5010,N_5470);
or U6216 (N_6216,N_5417,N_5369);
and U6217 (N_6217,N_5492,N_5727);
or U6218 (N_6218,N_5290,N_5443);
or U6219 (N_6219,N_5947,N_5511);
nor U6220 (N_6220,N_5015,N_5923);
and U6221 (N_6221,N_5794,N_5427);
nor U6222 (N_6222,N_5481,N_5931);
and U6223 (N_6223,N_5973,N_5804);
nand U6224 (N_6224,N_5344,N_5812);
and U6225 (N_6225,N_5552,N_5854);
nand U6226 (N_6226,N_5072,N_5591);
and U6227 (N_6227,N_5388,N_5196);
and U6228 (N_6228,N_5182,N_5580);
or U6229 (N_6229,N_5874,N_5681);
or U6230 (N_6230,N_5311,N_5850);
and U6231 (N_6231,N_5643,N_5942);
nand U6232 (N_6232,N_5630,N_5756);
and U6233 (N_6233,N_5397,N_5083);
and U6234 (N_6234,N_5067,N_5508);
nand U6235 (N_6235,N_5581,N_5123);
nor U6236 (N_6236,N_5902,N_5296);
and U6237 (N_6237,N_5886,N_5725);
or U6238 (N_6238,N_5565,N_5840);
and U6239 (N_6239,N_5146,N_5714);
or U6240 (N_6240,N_5875,N_5333);
nor U6241 (N_6241,N_5491,N_5007);
and U6242 (N_6242,N_5360,N_5700);
and U6243 (N_6243,N_5653,N_5176);
nand U6244 (N_6244,N_5561,N_5873);
and U6245 (N_6245,N_5177,N_5404);
and U6246 (N_6246,N_5047,N_5717);
or U6247 (N_6247,N_5839,N_5876);
nor U6248 (N_6248,N_5913,N_5051);
or U6249 (N_6249,N_5764,N_5726);
or U6250 (N_6250,N_5186,N_5059);
and U6251 (N_6251,N_5640,N_5450);
nor U6252 (N_6252,N_5157,N_5436);
and U6253 (N_6253,N_5424,N_5984);
and U6254 (N_6254,N_5212,N_5790);
nor U6255 (N_6255,N_5058,N_5779);
or U6256 (N_6256,N_5265,N_5638);
nand U6257 (N_6257,N_5889,N_5760);
nor U6258 (N_6258,N_5484,N_5155);
or U6259 (N_6259,N_5389,N_5660);
xnor U6260 (N_6260,N_5584,N_5422);
and U6261 (N_6261,N_5940,N_5966);
and U6262 (N_6262,N_5744,N_5168);
nand U6263 (N_6263,N_5863,N_5568);
and U6264 (N_6264,N_5468,N_5461);
and U6265 (N_6265,N_5774,N_5593);
or U6266 (N_6266,N_5253,N_5836);
nand U6267 (N_6267,N_5320,N_5244);
nand U6268 (N_6268,N_5948,N_5685);
nand U6269 (N_6269,N_5789,N_5415);
nor U6270 (N_6270,N_5021,N_5273);
or U6271 (N_6271,N_5163,N_5788);
nor U6272 (N_6272,N_5572,N_5107);
nor U6273 (N_6273,N_5079,N_5370);
and U6274 (N_6274,N_5255,N_5516);
nor U6275 (N_6275,N_5757,N_5666);
nand U6276 (N_6276,N_5448,N_5976);
and U6277 (N_6277,N_5390,N_5297);
or U6278 (N_6278,N_5054,N_5570);
nand U6279 (N_6279,N_5925,N_5206);
and U6280 (N_6280,N_5316,N_5395);
nor U6281 (N_6281,N_5831,N_5579);
and U6282 (N_6282,N_5618,N_5279);
or U6283 (N_6283,N_5035,N_5192);
or U6284 (N_6284,N_5908,N_5864);
and U6285 (N_6285,N_5911,N_5241);
or U6286 (N_6286,N_5611,N_5425);
nand U6287 (N_6287,N_5138,N_5031);
or U6288 (N_6288,N_5442,N_5232);
nand U6289 (N_6289,N_5745,N_5890);
nor U6290 (N_6290,N_5669,N_5807);
and U6291 (N_6291,N_5141,N_5387);
and U6292 (N_6292,N_5504,N_5671);
nor U6293 (N_6293,N_5383,N_5181);
nor U6294 (N_6294,N_5209,N_5142);
nor U6295 (N_6295,N_5663,N_5892);
and U6296 (N_6296,N_5771,N_5538);
nand U6297 (N_6297,N_5856,N_5195);
nand U6298 (N_6298,N_5647,N_5221);
or U6299 (N_6299,N_5945,N_5216);
or U6300 (N_6300,N_5982,N_5754);
and U6301 (N_6301,N_5975,N_5992);
nor U6302 (N_6302,N_5303,N_5998);
nor U6303 (N_6303,N_5030,N_5617);
xnor U6304 (N_6304,N_5783,N_5699);
and U6305 (N_6305,N_5194,N_5043);
nor U6306 (N_6306,N_5117,N_5201);
or U6307 (N_6307,N_5822,N_5934);
or U6308 (N_6308,N_5451,N_5742);
nand U6309 (N_6309,N_5218,N_5315);
nor U6310 (N_6310,N_5521,N_5590);
nand U6311 (N_6311,N_5364,N_5599);
nor U6312 (N_6312,N_5323,N_5103);
and U6313 (N_6313,N_5193,N_5307);
nand U6314 (N_6314,N_5490,N_5537);
or U6315 (N_6315,N_5166,N_5406);
and U6316 (N_6316,N_5814,N_5119);
or U6317 (N_6317,N_5898,N_5720);
and U6318 (N_6318,N_5753,N_5466);
nand U6319 (N_6319,N_5286,N_5325);
or U6320 (N_6320,N_5623,N_5287);
and U6321 (N_6321,N_5578,N_5118);
and U6322 (N_6322,N_5487,N_5564);
nor U6323 (N_6323,N_5247,N_5747);
nand U6324 (N_6324,N_5260,N_5416);
nor U6325 (N_6325,N_5474,N_5879);
nor U6326 (N_6326,N_5306,N_5026);
and U6327 (N_6327,N_5932,N_5235);
nand U6328 (N_6328,N_5501,N_5160);
nor U6329 (N_6329,N_5716,N_5438);
and U6330 (N_6330,N_5816,N_5526);
nor U6331 (N_6331,N_5703,N_5479);
or U6332 (N_6332,N_5066,N_5111);
nand U6333 (N_6333,N_5250,N_5226);
and U6334 (N_6334,N_5368,N_5135);
nand U6335 (N_6335,N_5556,N_5321);
nor U6336 (N_6336,N_5602,N_5348);
nand U6337 (N_6337,N_5447,N_5792);
nand U6338 (N_6338,N_5740,N_5460);
or U6339 (N_6339,N_5191,N_5928);
nor U6340 (N_6340,N_5238,N_5905);
nand U6341 (N_6341,N_5571,N_5329);
nor U6342 (N_6342,N_5826,N_5133);
or U6343 (N_6343,N_5024,N_5412);
nor U6344 (N_6344,N_5651,N_5918);
or U6345 (N_6345,N_5324,N_5633);
nand U6346 (N_6346,N_5625,N_5828);
nor U6347 (N_6347,N_5435,N_5880);
and U6348 (N_6348,N_5715,N_5278);
nor U6349 (N_6349,N_5090,N_5401);
or U6350 (N_6350,N_5805,N_5659);
and U6351 (N_6351,N_5486,N_5821);
nand U6352 (N_6352,N_5723,N_5245);
nand U6353 (N_6353,N_5775,N_5077);
nand U6354 (N_6354,N_5619,N_5326);
nor U6355 (N_6355,N_5962,N_5567);
nand U6356 (N_6356,N_5536,N_5352);
and U6357 (N_6357,N_5159,N_5027);
nor U6358 (N_6358,N_5281,N_5456);
and U6359 (N_6359,N_5113,N_5080);
xor U6360 (N_6360,N_5818,N_5258);
and U6361 (N_6361,N_5086,N_5065);
or U6362 (N_6362,N_5808,N_5335);
nand U6363 (N_6363,N_5188,N_5855);
nand U6364 (N_6364,N_5786,N_5896);
and U6365 (N_6365,N_5676,N_5517);
or U6366 (N_6366,N_5075,N_5161);
and U6367 (N_6367,N_5852,N_5295);
and U6368 (N_6368,N_5989,N_5799);
nor U6369 (N_6369,N_5139,N_5225);
and U6370 (N_6370,N_5712,N_5505);
or U6371 (N_6371,N_5023,N_5878);
or U6372 (N_6372,N_5739,N_5869);
and U6373 (N_6373,N_5013,N_5341);
or U6374 (N_6374,N_5881,N_5000);
or U6375 (N_6375,N_5037,N_5861);
or U6376 (N_6376,N_5398,N_5137);
or U6377 (N_6377,N_5304,N_5073);
nand U6378 (N_6378,N_5234,N_5345);
or U6379 (N_6379,N_5005,N_5654);
nor U6380 (N_6380,N_5767,N_5667);
nand U6381 (N_6381,N_5972,N_5342);
and U6382 (N_6382,N_5402,N_5782);
and U6383 (N_6383,N_5009,N_5531);
nand U6384 (N_6384,N_5359,N_5288);
and U6385 (N_6385,N_5052,N_5229);
nor U6386 (N_6386,N_5796,N_5639);
nand U6387 (N_6387,N_5105,N_5632);
or U6388 (N_6388,N_5409,N_5008);
and U6389 (N_6389,N_5965,N_5708);
nor U6390 (N_6390,N_5207,N_5457);
nor U6391 (N_6391,N_5115,N_5473);
nand U6392 (N_6392,N_5729,N_5939);
and U6393 (N_6393,N_5608,N_5539);
nand U6394 (N_6394,N_5318,N_5434);
nand U6395 (N_6395,N_5164,N_5285);
nand U6396 (N_6396,N_5350,N_5909);
or U6397 (N_6397,N_5102,N_5785);
and U6398 (N_6398,N_5768,N_5372);
or U6399 (N_6399,N_5641,N_5541);
nor U6400 (N_6400,N_5101,N_5087);
nand U6401 (N_6401,N_5252,N_5128);
or U6402 (N_6402,N_5011,N_5952);
nor U6403 (N_6403,N_5332,N_5276);
nor U6404 (N_6404,N_5376,N_5213);
and U6405 (N_6405,N_5800,N_5941);
nand U6406 (N_6406,N_5240,N_5249);
nor U6407 (N_6407,N_5312,N_5848);
nor U6408 (N_6408,N_5849,N_5857);
nand U6409 (N_6409,N_5711,N_5780);
or U6410 (N_6410,N_5710,N_5620);
nand U6411 (N_6411,N_5842,N_5680);
nand U6412 (N_6412,N_5408,N_5897);
and U6413 (N_6413,N_5154,N_5907);
and U6414 (N_6414,N_5540,N_5922);
nand U6415 (N_6415,N_5895,N_5122);
nor U6416 (N_6416,N_5652,N_5033);
nand U6417 (N_6417,N_5657,N_5582);
nor U6418 (N_6418,N_5899,N_5916);
nand U6419 (N_6419,N_5134,N_5587);
or U6420 (N_6420,N_5156,N_5609);
nand U6421 (N_6421,N_5733,N_5542);
or U6422 (N_6422,N_5096,N_5053);
and U6423 (N_6423,N_5777,N_5125);
or U6424 (N_6424,N_5518,N_5957);
or U6425 (N_6425,N_5496,N_5637);
nand U6426 (N_6426,N_5603,N_5656);
nor U6427 (N_6427,N_5706,N_5167);
nand U6428 (N_6428,N_5477,N_5056);
nand U6429 (N_6429,N_5954,N_5520);
nand U6430 (N_6430,N_5929,N_5489);
and U6431 (N_6431,N_5683,N_5601);
nand U6432 (N_6432,N_5860,N_5883);
nand U6433 (N_6433,N_5995,N_5573);
nor U6434 (N_6434,N_5732,N_5446);
or U6435 (N_6435,N_5375,N_5441);
or U6436 (N_6436,N_5661,N_5351);
nand U6437 (N_6437,N_5713,N_5917);
nor U6438 (N_6438,N_5227,N_5558);
and U6439 (N_6439,N_5910,N_5472);
nand U6440 (N_6440,N_5413,N_5577);
nor U6441 (N_6441,N_5793,N_5977);
or U6442 (N_6442,N_5108,N_5548);
and U6443 (N_6443,N_5129,N_5165);
nand U6444 (N_6444,N_5811,N_5604);
nand U6445 (N_6445,N_5082,N_5459);
nor U6446 (N_6446,N_5566,N_5394);
and U6447 (N_6447,N_5598,N_5868);
nor U6448 (N_6448,N_5174,N_5968);
nor U6449 (N_6449,N_5017,N_5631);
xnor U6450 (N_6450,N_5280,N_5302);
nor U6451 (N_6451,N_5498,N_5445);
nand U6452 (N_6452,N_5471,N_5629);
or U6453 (N_6453,N_5085,N_5830);
nand U6454 (N_6454,N_5334,N_5282);
or U6455 (N_6455,N_5419,N_5546);
and U6456 (N_6456,N_5615,N_5036);
nand U6457 (N_6457,N_5337,N_5919);
and U6458 (N_6458,N_5420,N_5806);
nor U6459 (N_6459,N_5462,N_5127);
nand U6460 (N_6460,N_5763,N_5223);
nor U6461 (N_6461,N_5076,N_5885);
xnor U6462 (N_6462,N_5044,N_5778);
nor U6463 (N_6463,N_5063,N_5243);
and U6464 (N_6464,N_5798,N_5291);
and U6465 (N_6465,N_5642,N_5655);
or U6466 (N_6466,N_5891,N_5844);
nor U6467 (N_6467,N_5393,N_5882);
nand U6468 (N_6468,N_5016,N_5920);
and U6469 (N_6469,N_5906,N_5859);
nor U6470 (N_6470,N_5884,N_5682);
or U6471 (N_6471,N_5331,N_5963);
nand U6472 (N_6472,N_5340,N_5257);
or U6473 (N_6473,N_5091,N_5392);
and U6474 (N_6474,N_5197,N_5583);
and U6475 (N_6475,N_5765,N_5524);
nand U6476 (N_6476,N_5205,N_5946);
and U6477 (N_6477,N_5093,N_5719);
or U6478 (N_6478,N_5959,N_5694);
or U6479 (N_6479,N_5284,N_5313);
or U6480 (N_6480,N_5595,N_5535);
nor U6481 (N_6481,N_5574,N_5668);
nand U6482 (N_6482,N_5846,N_5112);
nor U6483 (N_6483,N_5045,N_5029);
and U6484 (N_6484,N_5696,N_5038);
nor U6485 (N_6485,N_5759,N_5228);
nor U6486 (N_6486,N_5749,N_5428);
nand U6487 (N_6487,N_5095,N_5662);
or U6488 (N_6488,N_5994,N_5684);
and U6489 (N_6489,N_5961,N_5797);
or U6490 (N_6490,N_5131,N_5746);
and U6491 (N_6491,N_5926,N_5543);
and U6492 (N_6492,N_5210,N_5833);
and U6493 (N_6493,N_5596,N_5522);
and U6494 (N_6494,N_5560,N_5439);
nor U6495 (N_6495,N_5373,N_5173);
and U6496 (N_6496,N_5999,N_5967);
nor U6497 (N_6497,N_5912,N_5851);
and U6498 (N_6498,N_5634,N_5081);
or U6499 (N_6499,N_5607,N_5452);
nor U6500 (N_6500,N_5290,N_5511);
or U6501 (N_6501,N_5463,N_5299);
nand U6502 (N_6502,N_5184,N_5915);
nor U6503 (N_6503,N_5342,N_5842);
nor U6504 (N_6504,N_5974,N_5379);
or U6505 (N_6505,N_5704,N_5821);
nor U6506 (N_6506,N_5745,N_5265);
nor U6507 (N_6507,N_5024,N_5582);
and U6508 (N_6508,N_5458,N_5798);
nand U6509 (N_6509,N_5612,N_5794);
and U6510 (N_6510,N_5458,N_5552);
nand U6511 (N_6511,N_5297,N_5593);
and U6512 (N_6512,N_5290,N_5669);
nor U6513 (N_6513,N_5233,N_5125);
nor U6514 (N_6514,N_5759,N_5139);
and U6515 (N_6515,N_5323,N_5910);
or U6516 (N_6516,N_5121,N_5581);
or U6517 (N_6517,N_5255,N_5004);
nor U6518 (N_6518,N_5976,N_5856);
and U6519 (N_6519,N_5163,N_5576);
or U6520 (N_6520,N_5681,N_5629);
and U6521 (N_6521,N_5236,N_5479);
nand U6522 (N_6522,N_5792,N_5366);
or U6523 (N_6523,N_5432,N_5668);
nor U6524 (N_6524,N_5303,N_5171);
nor U6525 (N_6525,N_5073,N_5576);
and U6526 (N_6526,N_5880,N_5199);
nor U6527 (N_6527,N_5531,N_5582);
and U6528 (N_6528,N_5082,N_5407);
nor U6529 (N_6529,N_5429,N_5428);
nor U6530 (N_6530,N_5140,N_5380);
nand U6531 (N_6531,N_5088,N_5181);
or U6532 (N_6532,N_5461,N_5469);
nor U6533 (N_6533,N_5903,N_5708);
or U6534 (N_6534,N_5609,N_5864);
and U6535 (N_6535,N_5315,N_5777);
nand U6536 (N_6536,N_5375,N_5943);
or U6537 (N_6537,N_5172,N_5256);
or U6538 (N_6538,N_5551,N_5544);
nor U6539 (N_6539,N_5395,N_5045);
nor U6540 (N_6540,N_5162,N_5013);
or U6541 (N_6541,N_5685,N_5777);
and U6542 (N_6542,N_5954,N_5722);
nor U6543 (N_6543,N_5632,N_5329);
or U6544 (N_6544,N_5301,N_5665);
nor U6545 (N_6545,N_5166,N_5963);
nor U6546 (N_6546,N_5710,N_5314);
nand U6547 (N_6547,N_5673,N_5714);
nand U6548 (N_6548,N_5148,N_5200);
or U6549 (N_6549,N_5593,N_5989);
and U6550 (N_6550,N_5047,N_5129);
nand U6551 (N_6551,N_5173,N_5804);
nor U6552 (N_6552,N_5490,N_5644);
nor U6553 (N_6553,N_5157,N_5815);
nor U6554 (N_6554,N_5576,N_5616);
nand U6555 (N_6555,N_5450,N_5136);
nor U6556 (N_6556,N_5433,N_5474);
nor U6557 (N_6557,N_5944,N_5262);
or U6558 (N_6558,N_5700,N_5031);
nor U6559 (N_6559,N_5109,N_5990);
nand U6560 (N_6560,N_5565,N_5556);
xor U6561 (N_6561,N_5518,N_5140);
and U6562 (N_6562,N_5605,N_5451);
nand U6563 (N_6563,N_5969,N_5048);
or U6564 (N_6564,N_5762,N_5799);
nor U6565 (N_6565,N_5221,N_5340);
nand U6566 (N_6566,N_5798,N_5832);
or U6567 (N_6567,N_5269,N_5060);
and U6568 (N_6568,N_5195,N_5640);
and U6569 (N_6569,N_5169,N_5746);
nor U6570 (N_6570,N_5854,N_5344);
nor U6571 (N_6571,N_5381,N_5687);
or U6572 (N_6572,N_5160,N_5092);
nor U6573 (N_6573,N_5946,N_5520);
nand U6574 (N_6574,N_5077,N_5539);
nor U6575 (N_6575,N_5082,N_5587);
nand U6576 (N_6576,N_5208,N_5505);
nand U6577 (N_6577,N_5445,N_5974);
nand U6578 (N_6578,N_5631,N_5346);
nor U6579 (N_6579,N_5051,N_5488);
or U6580 (N_6580,N_5792,N_5190);
nand U6581 (N_6581,N_5000,N_5396);
and U6582 (N_6582,N_5375,N_5201);
nor U6583 (N_6583,N_5384,N_5232);
or U6584 (N_6584,N_5457,N_5981);
or U6585 (N_6585,N_5467,N_5799);
or U6586 (N_6586,N_5030,N_5864);
nand U6587 (N_6587,N_5415,N_5112);
nor U6588 (N_6588,N_5184,N_5831);
or U6589 (N_6589,N_5676,N_5329);
nand U6590 (N_6590,N_5430,N_5732);
nand U6591 (N_6591,N_5221,N_5673);
or U6592 (N_6592,N_5239,N_5802);
nor U6593 (N_6593,N_5707,N_5679);
nand U6594 (N_6594,N_5798,N_5587);
and U6595 (N_6595,N_5523,N_5792);
nor U6596 (N_6596,N_5156,N_5406);
nor U6597 (N_6597,N_5771,N_5117);
or U6598 (N_6598,N_5323,N_5486);
or U6599 (N_6599,N_5509,N_5153);
or U6600 (N_6600,N_5675,N_5798);
and U6601 (N_6601,N_5279,N_5806);
nand U6602 (N_6602,N_5636,N_5450);
or U6603 (N_6603,N_5799,N_5671);
nand U6604 (N_6604,N_5465,N_5040);
nor U6605 (N_6605,N_5126,N_5058);
or U6606 (N_6606,N_5048,N_5268);
nor U6607 (N_6607,N_5812,N_5835);
or U6608 (N_6608,N_5892,N_5515);
or U6609 (N_6609,N_5449,N_5623);
and U6610 (N_6610,N_5798,N_5258);
nand U6611 (N_6611,N_5374,N_5092);
and U6612 (N_6612,N_5974,N_5666);
and U6613 (N_6613,N_5498,N_5063);
or U6614 (N_6614,N_5729,N_5950);
nor U6615 (N_6615,N_5319,N_5030);
nor U6616 (N_6616,N_5789,N_5391);
and U6617 (N_6617,N_5267,N_5276);
nand U6618 (N_6618,N_5174,N_5412);
and U6619 (N_6619,N_5610,N_5127);
nand U6620 (N_6620,N_5667,N_5716);
and U6621 (N_6621,N_5240,N_5309);
and U6622 (N_6622,N_5767,N_5508);
nand U6623 (N_6623,N_5353,N_5966);
and U6624 (N_6624,N_5194,N_5291);
or U6625 (N_6625,N_5323,N_5935);
nand U6626 (N_6626,N_5052,N_5838);
nor U6627 (N_6627,N_5124,N_5229);
or U6628 (N_6628,N_5197,N_5631);
nor U6629 (N_6629,N_5530,N_5196);
or U6630 (N_6630,N_5523,N_5559);
nand U6631 (N_6631,N_5490,N_5088);
and U6632 (N_6632,N_5315,N_5133);
or U6633 (N_6633,N_5481,N_5627);
nor U6634 (N_6634,N_5974,N_5423);
nand U6635 (N_6635,N_5495,N_5961);
nand U6636 (N_6636,N_5316,N_5712);
nor U6637 (N_6637,N_5787,N_5913);
nand U6638 (N_6638,N_5774,N_5847);
and U6639 (N_6639,N_5585,N_5278);
nand U6640 (N_6640,N_5314,N_5305);
and U6641 (N_6641,N_5122,N_5662);
xnor U6642 (N_6642,N_5845,N_5240);
nand U6643 (N_6643,N_5515,N_5885);
nand U6644 (N_6644,N_5206,N_5504);
nand U6645 (N_6645,N_5386,N_5912);
and U6646 (N_6646,N_5577,N_5343);
or U6647 (N_6647,N_5832,N_5117);
nand U6648 (N_6648,N_5914,N_5246);
nor U6649 (N_6649,N_5747,N_5917);
nand U6650 (N_6650,N_5969,N_5582);
nand U6651 (N_6651,N_5875,N_5115);
or U6652 (N_6652,N_5828,N_5251);
and U6653 (N_6653,N_5358,N_5809);
and U6654 (N_6654,N_5227,N_5291);
or U6655 (N_6655,N_5311,N_5159);
nor U6656 (N_6656,N_5146,N_5776);
nand U6657 (N_6657,N_5222,N_5749);
and U6658 (N_6658,N_5930,N_5284);
nor U6659 (N_6659,N_5236,N_5834);
nand U6660 (N_6660,N_5643,N_5632);
nor U6661 (N_6661,N_5876,N_5731);
nor U6662 (N_6662,N_5545,N_5960);
nor U6663 (N_6663,N_5993,N_5567);
nand U6664 (N_6664,N_5906,N_5235);
nor U6665 (N_6665,N_5528,N_5296);
nor U6666 (N_6666,N_5545,N_5640);
and U6667 (N_6667,N_5092,N_5675);
nand U6668 (N_6668,N_5841,N_5253);
and U6669 (N_6669,N_5595,N_5202);
and U6670 (N_6670,N_5902,N_5380);
xnor U6671 (N_6671,N_5462,N_5731);
or U6672 (N_6672,N_5506,N_5531);
nor U6673 (N_6673,N_5341,N_5547);
nor U6674 (N_6674,N_5181,N_5218);
nor U6675 (N_6675,N_5993,N_5918);
and U6676 (N_6676,N_5574,N_5441);
nor U6677 (N_6677,N_5017,N_5964);
nor U6678 (N_6678,N_5488,N_5817);
or U6679 (N_6679,N_5684,N_5878);
nand U6680 (N_6680,N_5954,N_5658);
nor U6681 (N_6681,N_5213,N_5267);
nor U6682 (N_6682,N_5171,N_5181);
nor U6683 (N_6683,N_5797,N_5918);
nand U6684 (N_6684,N_5070,N_5748);
nand U6685 (N_6685,N_5542,N_5750);
or U6686 (N_6686,N_5900,N_5232);
or U6687 (N_6687,N_5301,N_5587);
nor U6688 (N_6688,N_5316,N_5541);
nand U6689 (N_6689,N_5856,N_5565);
and U6690 (N_6690,N_5610,N_5667);
and U6691 (N_6691,N_5041,N_5863);
nor U6692 (N_6692,N_5297,N_5817);
and U6693 (N_6693,N_5647,N_5476);
and U6694 (N_6694,N_5261,N_5962);
nor U6695 (N_6695,N_5728,N_5621);
or U6696 (N_6696,N_5585,N_5896);
nor U6697 (N_6697,N_5113,N_5445);
nand U6698 (N_6698,N_5100,N_5592);
nor U6699 (N_6699,N_5327,N_5312);
or U6700 (N_6700,N_5441,N_5150);
or U6701 (N_6701,N_5815,N_5509);
nand U6702 (N_6702,N_5942,N_5892);
and U6703 (N_6703,N_5153,N_5983);
or U6704 (N_6704,N_5638,N_5523);
nand U6705 (N_6705,N_5079,N_5479);
nand U6706 (N_6706,N_5410,N_5018);
and U6707 (N_6707,N_5154,N_5943);
nor U6708 (N_6708,N_5906,N_5111);
nand U6709 (N_6709,N_5082,N_5365);
nor U6710 (N_6710,N_5997,N_5897);
nor U6711 (N_6711,N_5692,N_5619);
nor U6712 (N_6712,N_5305,N_5736);
nand U6713 (N_6713,N_5005,N_5629);
nor U6714 (N_6714,N_5064,N_5354);
nand U6715 (N_6715,N_5238,N_5712);
and U6716 (N_6716,N_5123,N_5890);
and U6717 (N_6717,N_5193,N_5597);
or U6718 (N_6718,N_5281,N_5201);
nor U6719 (N_6719,N_5589,N_5159);
nor U6720 (N_6720,N_5473,N_5583);
nand U6721 (N_6721,N_5464,N_5160);
and U6722 (N_6722,N_5540,N_5995);
nor U6723 (N_6723,N_5830,N_5043);
nand U6724 (N_6724,N_5563,N_5500);
and U6725 (N_6725,N_5921,N_5977);
nor U6726 (N_6726,N_5389,N_5990);
or U6727 (N_6727,N_5026,N_5935);
or U6728 (N_6728,N_5240,N_5375);
or U6729 (N_6729,N_5014,N_5892);
and U6730 (N_6730,N_5590,N_5090);
nand U6731 (N_6731,N_5271,N_5837);
and U6732 (N_6732,N_5267,N_5682);
nand U6733 (N_6733,N_5603,N_5408);
nand U6734 (N_6734,N_5346,N_5556);
nor U6735 (N_6735,N_5035,N_5172);
or U6736 (N_6736,N_5379,N_5838);
and U6737 (N_6737,N_5983,N_5055);
nor U6738 (N_6738,N_5123,N_5190);
nand U6739 (N_6739,N_5498,N_5330);
nand U6740 (N_6740,N_5813,N_5319);
or U6741 (N_6741,N_5611,N_5487);
nor U6742 (N_6742,N_5771,N_5232);
and U6743 (N_6743,N_5829,N_5264);
and U6744 (N_6744,N_5970,N_5326);
and U6745 (N_6745,N_5662,N_5067);
and U6746 (N_6746,N_5062,N_5740);
and U6747 (N_6747,N_5467,N_5049);
or U6748 (N_6748,N_5510,N_5005);
nand U6749 (N_6749,N_5729,N_5887);
or U6750 (N_6750,N_5011,N_5057);
nor U6751 (N_6751,N_5927,N_5339);
and U6752 (N_6752,N_5665,N_5408);
and U6753 (N_6753,N_5189,N_5827);
nand U6754 (N_6754,N_5904,N_5184);
nor U6755 (N_6755,N_5543,N_5669);
or U6756 (N_6756,N_5649,N_5658);
or U6757 (N_6757,N_5413,N_5359);
and U6758 (N_6758,N_5554,N_5238);
nand U6759 (N_6759,N_5167,N_5348);
or U6760 (N_6760,N_5992,N_5000);
nor U6761 (N_6761,N_5450,N_5040);
and U6762 (N_6762,N_5056,N_5384);
and U6763 (N_6763,N_5602,N_5547);
nor U6764 (N_6764,N_5911,N_5105);
nor U6765 (N_6765,N_5398,N_5546);
nor U6766 (N_6766,N_5348,N_5783);
nand U6767 (N_6767,N_5820,N_5802);
or U6768 (N_6768,N_5461,N_5623);
nand U6769 (N_6769,N_5522,N_5224);
and U6770 (N_6770,N_5878,N_5356);
nor U6771 (N_6771,N_5756,N_5376);
xnor U6772 (N_6772,N_5836,N_5587);
nor U6773 (N_6773,N_5781,N_5716);
and U6774 (N_6774,N_5874,N_5401);
or U6775 (N_6775,N_5039,N_5267);
nor U6776 (N_6776,N_5186,N_5404);
nor U6777 (N_6777,N_5091,N_5989);
nand U6778 (N_6778,N_5754,N_5082);
and U6779 (N_6779,N_5903,N_5920);
and U6780 (N_6780,N_5667,N_5018);
or U6781 (N_6781,N_5186,N_5181);
nand U6782 (N_6782,N_5600,N_5346);
nor U6783 (N_6783,N_5766,N_5296);
nand U6784 (N_6784,N_5499,N_5081);
or U6785 (N_6785,N_5809,N_5886);
and U6786 (N_6786,N_5616,N_5710);
nor U6787 (N_6787,N_5652,N_5108);
or U6788 (N_6788,N_5238,N_5683);
or U6789 (N_6789,N_5803,N_5088);
nor U6790 (N_6790,N_5436,N_5971);
nor U6791 (N_6791,N_5904,N_5830);
nand U6792 (N_6792,N_5041,N_5604);
and U6793 (N_6793,N_5376,N_5332);
or U6794 (N_6794,N_5045,N_5504);
or U6795 (N_6795,N_5729,N_5811);
nor U6796 (N_6796,N_5420,N_5530);
nor U6797 (N_6797,N_5818,N_5904);
nand U6798 (N_6798,N_5937,N_5869);
nand U6799 (N_6799,N_5934,N_5870);
and U6800 (N_6800,N_5097,N_5322);
and U6801 (N_6801,N_5997,N_5128);
and U6802 (N_6802,N_5727,N_5417);
nand U6803 (N_6803,N_5246,N_5327);
nand U6804 (N_6804,N_5173,N_5688);
nor U6805 (N_6805,N_5108,N_5859);
nor U6806 (N_6806,N_5440,N_5738);
nor U6807 (N_6807,N_5843,N_5625);
and U6808 (N_6808,N_5400,N_5156);
and U6809 (N_6809,N_5980,N_5472);
nand U6810 (N_6810,N_5974,N_5132);
nand U6811 (N_6811,N_5246,N_5927);
nor U6812 (N_6812,N_5768,N_5848);
or U6813 (N_6813,N_5547,N_5256);
nor U6814 (N_6814,N_5492,N_5368);
and U6815 (N_6815,N_5682,N_5815);
and U6816 (N_6816,N_5067,N_5044);
nor U6817 (N_6817,N_5827,N_5759);
xor U6818 (N_6818,N_5846,N_5914);
nand U6819 (N_6819,N_5110,N_5675);
and U6820 (N_6820,N_5691,N_5575);
nor U6821 (N_6821,N_5881,N_5343);
or U6822 (N_6822,N_5298,N_5815);
or U6823 (N_6823,N_5875,N_5725);
or U6824 (N_6824,N_5927,N_5840);
or U6825 (N_6825,N_5670,N_5956);
nand U6826 (N_6826,N_5411,N_5758);
and U6827 (N_6827,N_5629,N_5516);
and U6828 (N_6828,N_5300,N_5536);
or U6829 (N_6829,N_5165,N_5701);
nor U6830 (N_6830,N_5721,N_5035);
or U6831 (N_6831,N_5690,N_5419);
nor U6832 (N_6832,N_5454,N_5356);
or U6833 (N_6833,N_5542,N_5380);
or U6834 (N_6834,N_5663,N_5544);
nor U6835 (N_6835,N_5720,N_5591);
nand U6836 (N_6836,N_5876,N_5991);
nand U6837 (N_6837,N_5652,N_5365);
nand U6838 (N_6838,N_5749,N_5485);
and U6839 (N_6839,N_5424,N_5792);
nor U6840 (N_6840,N_5626,N_5643);
and U6841 (N_6841,N_5560,N_5178);
nor U6842 (N_6842,N_5430,N_5006);
and U6843 (N_6843,N_5323,N_5846);
nor U6844 (N_6844,N_5807,N_5304);
nand U6845 (N_6845,N_5123,N_5224);
or U6846 (N_6846,N_5392,N_5775);
or U6847 (N_6847,N_5658,N_5309);
or U6848 (N_6848,N_5820,N_5953);
nor U6849 (N_6849,N_5184,N_5446);
nand U6850 (N_6850,N_5019,N_5581);
nand U6851 (N_6851,N_5996,N_5790);
nor U6852 (N_6852,N_5722,N_5336);
or U6853 (N_6853,N_5387,N_5786);
nand U6854 (N_6854,N_5454,N_5754);
nor U6855 (N_6855,N_5984,N_5906);
nor U6856 (N_6856,N_5666,N_5829);
nand U6857 (N_6857,N_5329,N_5520);
and U6858 (N_6858,N_5116,N_5938);
or U6859 (N_6859,N_5359,N_5453);
nor U6860 (N_6860,N_5209,N_5804);
nand U6861 (N_6861,N_5846,N_5105);
and U6862 (N_6862,N_5327,N_5844);
nand U6863 (N_6863,N_5151,N_5677);
or U6864 (N_6864,N_5088,N_5819);
nand U6865 (N_6865,N_5182,N_5820);
nand U6866 (N_6866,N_5255,N_5447);
nor U6867 (N_6867,N_5505,N_5581);
or U6868 (N_6868,N_5009,N_5327);
and U6869 (N_6869,N_5459,N_5837);
and U6870 (N_6870,N_5587,N_5980);
nand U6871 (N_6871,N_5381,N_5794);
and U6872 (N_6872,N_5088,N_5191);
nand U6873 (N_6873,N_5431,N_5677);
nand U6874 (N_6874,N_5581,N_5168);
nand U6875 (N_6875,N_5475,N_5654);
nand U6876 (N_6876,N_5098,N_5477);
nand U6877 (N_6877,N_5741,N_5500);
nor U6878 (N_6878,N_5676,N_5811);
and U6879 (N_6879,N_5031,N_5686);
and U6880 (N_6880,N_5309,N_5290);
and U6881 (N_6881,N_5963,N_5734);
nand U6882 (N_6882,N_5500,N_5874);
nand U6883 (N_6883,N_5656,N_5032);
nor U6884 (N_6884,N_5929,N_5355);
nand U6885 (N_6885,N_5155,N_5367);
and U6886 (N_6886,N_5421,N_5182);
and U6887 (N_6887,N_5963,N_5500);
xnor U6888 (N_6888,N_5479,N_5584);
or U6889 (N_6889,N_5821,N_5752);
nor U6890 (N_6890,N_5166,N_5105);
nor U6891 (N_6891,N_5774,N_5037);
nor U6892 (N_6892,N_5863,N_5758);
nand U6893 (N_6893,N_5462,N_5764);
nor U6894 (N_6894,N_5314,N_5774);
nor U6895 (N_6895,N_5830,N_5326);
nor U6896 (N_6896,N_5780,N_5120);
or U6897 (N_6897,N_5864,N_5992);
and U6898 (N_6898,N_5909,N_5808);
or U6899 (N_6899,N_5817,N_5555);
nand U6900 (N_6900,N_5662,N_5663);
or U6901 (N_6901,N_5227,N_5163);
or U6902 (N_6902,N_5541,N_5268);
nor U6903 (N_6903,N_5757,N_5360);
nor U6904 (N_6904,N_5975,N_5045);
nand U6905 (N_6905,N_5652,N_5382);
nor U6906 (N_6906,N_5876,N_5699);
nor U6907 (N_6907,N_5589,N_5798);
or U6908 (N_6908,N_5227,N_5521);
or U6909 (N_6909,N_5137,N_5428);
nand U6910 (N_6910,N_5310,N_5368);
nand U6911 (N_6911,N_5683,N_5092);
and U6912 (N_6912,N_5423,N_5436);
nor U6913 (N_6913,N_5676,N_5066);
and U6914 (N_6914,N_5397,N_5584);
nand U6915 (N_6915,N_5617,N_5893);
nor U6916 (N_6916,N_5528,N_5263);
nor U6917 (N_6917,N_5302,N_5034);
or U6918 (N_6918,N_5444,N_5932);
and U6919 (N_6919,N_5243,N_5268);
and U6920 (N_6920,N_5348,N_5416);
nor U6921 (N_6921,N_5322,N_5452);
and U6922 (N_6922,N_5963,N_5354);
and U6923 (N_6923,N_5795,N_5296);
or U6924 (N_6924,N_5526,N_5996);
or U6925 (N_6925,N_5509,N_5521);
nor U6926 (N_6926,N_5797,N_5200);
or U6927 (N_6927,N_5051,N_5409);
nand U6928 (N_6928,N_5645,N_5212);
nand U6929 (N_6929,N_5516,N_5355);
or U6930 (N_6930,N_5913,N_5106);
or U6931 (N_6931,N_5602,N_5728);
or U6932 (N_6932,N_5606,N_5850);
and U6933 (N_6933,N_5495,N_5064);
or U6934 (N_6934,N_5423,N_5766);
nand U6935 (N_6935,N_5128,N_5106);
and U6936 (N_6936,N_5836,N_5588);
or U6937 (N_6937,N_5404,N_5801);
and U6938 (N_6938,N_5354,N_5685);
and U6939 (N_6939,N_5873,N_5449);
or U6940 (N_6940,N_5988,N_5000);
and U6941 (N_6941,N_5315,N_5408);
and U6942 (N_6942,N_5403,N_5220);
nand U6943 (N_6943,N_5517,N_5171);
and U6944 (N_6944,N_5167,N_5178);
nand U6945 (N_6945,N_5209,N_5807);
nand U6946 (N_6946,N_5763,N_5658);
and U6947 (N_6947,N_5702,N_5412);
or U6948 (N_6948,N_5320,N_5328);
nor U6949 (N_6949,N_5045,N_5318);
and U6950 (N_6950,N_5502,N_5331);
nor U6951 (N_6951,N_5341,N_5871);
nor U6952 (N_6952,N_5962,N_5797);
nand U6953 (N_6953,N_5773,N_5298);
and U6954 (N_6954,N_5906,N_5095);
and U6955 (N_6955,N_5842,N_5080);
nand U6956 (N_6956,N_5735,N_5065);
and U6957 (N_6957,N_5901,N_5198);
or U6958 (N_6958,N_5353,N_5323);
and U6959 (N_6959,N_5785,N_5355);
or U6960 (N_6960,N_5887,N_5851);
nand U6961 (N_6961,N_5050,N_5044);
and U6962 (N_6962,N_5036,N_5923);
and U6963 (N_6963,N_5217,N_5179);
nand U6964 (N_6964,N_5368,N_5470);
and U6965 (N_6965,N_5834,N_5986);
and U6966 (N_6966,N_5236,N_5710);
nand U6967 (N_6967,N_5433,N_5222);
nand U6968 (N_6968,N_5533,N_5936);
nand U6969 (N_6969,N_5661,N_5268);
nor U6970 (N_6970,N_5585,N_5221);
nor U6971 (N_6971,N_5133,N_5002);
nand U6972 (N_6972,N_5625,N_5759);
or U6973 (N_6973,N_5737,N_5040);
nand U6974 (N_6974,N_5823,N_5925);
nor U6975 (N_6975,N_5419,N_5782);
and U6976 (N_6976,N_5442,N_5378);
nor U6977 (N_6977,N_5718,N_5215);
nand U6978 (N_6978,N_5825,N_5155);
and U6979 (N_6979,N_5736,N_5990);
or U6980 (N_6980,N_5123,N_5310);
and U6981 (N_6981,N_5333,N_5564);
nand U6982 (N_6982,N_5049,N_5443);
and U6983 (N_6983,N_5321,N_5258);
and U6984 (N_6984,N_5259,N_5866);
and U6985 (N_6985,N_5261,N_5331);
and U6986 (N_6986,N_5622,N_5650);
or U6987 (N_6987,N_5330,N_5731);
nor U6988 (N_6988,N_5502,N_5225);
or U6989 (N_6989,N_5469,N_5997);
nor U6990 (N_6990,N_5487,N_5416);
or U6991 (N_6991,N_5227,N_5748);
nor U6992 (N_6992,N_5241,N_5906);
and U6993 (N_6993,N_5457,N_5578);
nor U6994 (N_6994,N_5444,N_5987);
nor U6995 (N_6995,N_5381,N_5999);
and U6996 (N_6996,N_5293,N_5462);
and U6997 (N_6997,N_5542,N_5850);
nor U6998 (N_6998,N_5499,N_5246);
nor U6999 (N_6999,N_5542,N_5986);
nor U7000 (N_7000,N_6691,N_6049);
and U7001 (N_7001,N_6760,N_6060);
nand U7002 (N_7002,N_6004,N_6882);
and U7003 (N_7003,N_6427,N_6542);
nor U7004 (N_7004,N_6536,N_6237);
and U7005 (N_7005,N_6675,N_6300);
or U7006 (N_7006,N_6965,N_6162);
or U7007 (N_7007,N_6916,N_6180);
or U7008 (N_7008,N_6490,N_6591);
nor U7009 (N_7009,N_6243,N_6870);
nand U7010 (N_7010,N_6374,N_6354);
or U7011 (N_7011,N_6346,N_6469);
nand U7012 (N_7012,N_6589,N_6830);
and U7013 (N_7013,N_6301,N_6550);
or U7014 (N_7014,N_6266,N_6358);
or U7015 (N_7015,N_6417,N_6385);
nor U7016 (N_7016,N_6624,N_6126);
nor U7017 (N_7017,N_6295,N_6885);
and U7018 (N_7018,N_6154,N_6523);
or U7019 (N_7019,N_6808,N_6616);
nand U7020 (N_7020,N_6373,N_6191);
and U7021 (N_7021,N_6176,N_6547);
nand U7022 (N_7022,N_6930,N_6002);
and U7023 (N_7023,N_6102,N_6441);
nand U7024 (N_7024,N_6360,N_6630);
and U7025 (N_7025,N_6357,N_6424);
nor U7026 (N_7026,N_6751,N_6397);
nand U7027 (N_7027,N_6474,N_6680);
nand U7028 (N_7028,N_6316,N_6085);
nor U7029 (N_7029,N_6826,N_6746);
xor U7030 (N_7030,N_6075,N_6911);
nor U7031 (N_7031,N_6655,N_6140);
nand U7032 (N_7032,N_6784,N_6718);
or U7033 (N_7033,N_6155,N_6650);
nand U7034 (N_7034,N_6643,N_6872);
nor U7035 (N_7035,N_6725,N_6976);
or U7036 (N_7036,N_6802,N_6782);
nand U7037 (N_7037,N_6289,N_6907);
or U7038 (N_7038,N_6721,N_6320);
nand U7039 (N_7039,N_6804,N_6009);
or U7040 (N_7040,N_6475,N_6188);
or U7041 (N_7041,N_6132,N_6539);
nand U7042 (N_7042,N_6489,N_6257);
nand U7043 (N_7043,N_6325,N_6311);
nand U7044 (N_7044,N_6747,N_6897);
nand U7045 (N_7045,N_6118,N_6278);
nor U7046 (N_7046,N_6090,N_6665);
and U7047 (N_7047,N_6919,N_6207);
and U7048 (N_7048,N_6444,N_6792);
xnor U7049 (N_7049,N_6184,N_6866);
and U7050 (N_7050,N_6371,N_6971);
and U7051 (N_7051,N_6669,N_6906);
or U7052 (N_7052,N_6969,N_6127);
and U7053 (N_7053,N_6964,N_6342);
and U7054 (N_7054,N_6011,N_6671);
xnor U7055 (N_7055,N_6921,N_6698);
nand U7056 (N_7056,N_6059,N_6776);
or U7057 (N_7057,N_6929,N_6046);
or U7058 (N_7058,N_6568,N_6533);
or U7059 (N_7059,N_6379,N_6816);
nor U7060 (N_7060,N_6734,N_6933);
nor U7061 (N_7061,N_6493,N_6708);
nand U7062 (N_7062,N_6491,N_6611);
nor U7063 (N_7063,N_6564,N_6666);
and U7064 (N_7064,N_6774,N_6309);
nor U7065 (N_7065,N_6876,N_6974);
or U7066 (N_7066,N_6306,N_6412);
and U7067 (N_7067,N_6731,N_6948);
nor U7068 (N_7068,N_6196,N_6399);
or U7069 (N_7069,N_6436,N_6101);
and U7070 (N_7070,N_6054,N_6363);
or U7071 (N_7071,N_6558,N_6231);
nor U7072 (N_7072,N_6451,N_6038);
or U7073 (N_7073,N_6852,N_6248);
and U7074 (N_7074,N_6323,N_6141);
and U7075 (N_7075,N_6472,N_6365);
and U7076 (N_7076,N_6604,N_6805);
nand U7077 (N_7077,N_6878,N_6771);
and U7078 (N_7078,N_6061,N_6211);
and U7079 (N_7079,N_6166,N_6429);
and U7080 (N_7080,N_6297,N_6647);
nor U7081 (N_7081,N_6256,N_6007);
or U7082 (N_7082,N_6736,N_6482);
or U7083 (N_7083,N_6039,N_6845);
or U7084 (N_7084,N_6202,N_6450);
nor U7085 (N_7085,N_6409,N_6770);
or U7086 (N_7086,N_6863,N_6064);
nor U7087 (N_7087,N_6631,N_6754);
and U7088 (N_7088,N_6087,N_6957);
and U7089 (N_7089,N_6821,N_6364);
and U7090 (N_7090,N_6795,N_6268);
and U7091 (N_7091,N_6983,N_6728);
or U7092 (N_7092,N_6672,N_6682);
nand U7093 (N_7093,N_6827,N_6464);
and U7094 (N_7094,N_6463,N_6065);
or U7095 (N_7095,N_6388,N_6701);
nor U7096 (N_7096,N_6926,N_6757);
and U7097 (N_7097,N_6572,N_6435);
or U7098 (N_7098,N_6766,N_6074);
or U7099 (N_7099,N_6567,N_6538);
nor U7100 (N_7100,N_6036,N_6692);
and U7101 (N_7101,N_6438,N_6648);
and U7102 (N_7102,N_6884,N_6186);
or U7103 (N_7103,N_6270,N_6258);
nor U7104 (N_7104,N_6273,N_6642);
and U7105 (N_7105,N_6952,N_6333);
and U7106 (N_7106,N_6857,N_6232);
nor U7107 (N_7107,N_6607,N_6503);
or U7108 (N_7108,N_6769,N_6540);
or U7109 (N_7109,N_6419,N_6145);
xor U7110 (N_7110,N_6891,N_6511);
nand U7111 (N_7111,N_6587,N_6578);
nor U7112 (N_7112,N_6645,N_6044);
or U7113 (N_7113,N_6218,N_6873);
and U7114 (N_7114,N_6430,N_6632);
and U7115 (N_7115,N_6886,N_6149);
nor U7116 (N_7116,N_6050,N_6513);
or U7117 (N_7117,N_6302,N_6308);
nor U7118 (N_7118,N_6019,N_6707);
nand U7119 (N_7119,N_6812,N_6209);
nor U7120 (N_7120,N_6849,N_6889);
and U7121 (N_7121,N_6673,N_6913);
and U7122 (N_7122,N_6329,N_6042);
nor U7123 (N_7123,N_6080,N_6192);
and U7124 (N_7124,N_6678,N_6481);
or U7125 (N_7125,N_6091,N_6428);
nor U7126 (N_7126,N_6875,N_6247);
xor U7127 (N_7127,N_6659,N_6510);
nand U7128 (N_7128,N_6381,N_6227);
and U7129 (N_7129,N_6025,N_6506);
and U7130 (N_7130,N_6996,N_6670);
and U7131 (N_7131,N_6076,N_6834);
nor U7132 (N_7132,N_6944,N_6173);
and U7133 (N_7133,N_6953,N_6923);
nor U7134 (N_7134,N_6825,N_6726);
nor U7135 (N_7135,N_6703,N_6443);
nor U7136 (N_7136,N_6226,N_6560);
nor U7137 (N_7137,N_6158,N_6146);
nor U7138 (N_7138,N_6597,N_6620);
or U7139 (N_7139,N_6844,N_6762);
or U7140 (N_7140,N_6487,N_6779);
nor U7141 (N_7141,N_6377,N_6148);
nand U7142 (N_7142,N_6265,N_6394);
or U7143 (N_7143,N_6240,N_6741);
or U7144 (N_7144,N_6445,N_6261);
or U7145 (N_7145,N_6110,N_6018);
and U7146 (N_7146,N_6874,N_6233);
or U7147 (N_7147,N_6125,N_6674);
and U7148 (N_7148,N_6775,N_6915);
nand U7149 (N_7149,N_6705,N_6330);
or U7150 (N_7150,N_6313,N_6225);
and U7151 (N_7151,N_6783,N_6425);
or U7152 (N_7152,N_6868,N_6937);
nand U7153 (N_7153,N_6350,N_6212);
nor U7154 (N_7154,N_6024,N_6794);
nor U7155 (N_7155,N_6910,N_6129);
nand U7156 (N_7156,N_6548,N_6835);
and U7157 (N_7157,N_6823,N_6153);
nand U7158 (N_7158,N_6294,N_6927);
nor U7159 (N_7159,N_6378,N_6277);
nand U7160 (N_7160,N_6848,N_6667);
and U7161 (N_7161,N_6987,N_6663);
and U7162 (N_7162,N_6175,N_6133);
and U7163 (N_7163,N_6956,N_6562);
or U7164 (N_7164,N_6405,N_6104);
and U7165 (N_7165,N_6094,N_6473);
nor U7166 (N_7166,N_6052,N_6841);
or U7167 (N_7167,N_6573,N_6727);
and U7168 (N_7168,N_6190,N_6807);
nand U7169 (N_7169,N_6738,N_6255);
nor U7170 (N_7170,N_6679,N_6084);
nand U7171 (N_7171,N_6189,N_6326);
or U7172 (N_7172,N_6390,N_6344);
and U7173 (N_7173,N_6434,N_6622);
nor U7174 (N_7174,N_6668,N_6809);
and U7175 (N_7175,N_6235,N_6498);
and U7176 (N_7176,N_6789,N_6496);
or U7177 (N_7177,N_6454,N_6341);
and U7178 (N_7178,N_6855,N_6459);
and U7179 (N_7179,N_6950,N_6415);
or U7180 (N_7180,N_6860,N_6994);
or U7181 (N_7181,N_6034,N_6281);
and U7182 (N_7182,N_6216,N_6082);
nor U7183 (N_7183,N_6628,N_6989);
nor U7184 (N_7184,N_6467,N_6858);
and U7185 (N_7185,N_6375,N_6296);
nor U7186 (N_7186,N_6546,N_6468);
and U7187 (N_7187,N_6995,N_6108);
and U7188 (N_7188,N_6970,N_6939);
nor U7189 (N_7189,N_6031,N_6136);
nor U7190 (N_7190,N_6793,N_6515);
nand U7191 (N_7191,N_6600,N_6709);
nor U7192 (N_7192,N_6520,N_6317);
nor U7193 (N_7193,N_6924,N_6095);
nand U7194 (N_7194,N_6383,N_6862);
nand U7195 (N_7195,N_6576,N_6071);
xnor U7196 (N_7196,N_6197,N_6951);
and U7197 (N_7197,N_6098,N_6206);
and U7198 (N_7198,N_6321,N_6656);
nand U7199 (N_7199,N_6012,N_6109);
and U7200 (N_7200,N_6492,N_6979);
or U7201 (N_7201,N_6410,N_6403);
or U7202 (N_7202,N_6456,N_6603);
or U7203 (N_7203,N_6017,N_6903);
nor U7204 (N_7204,N_6033,N_6078);
or U7205 (N_7205,N_6112,N_6635);
nor U7206 (N_7206,N_6246,N_6179);
or U7207 (N_7207,N_6391,N_6015);
nor U7208 (N_7208,N_6723,N_6219);
and U7209 (N_7209,N_6800,N_6097);
or U7210 (N_7210,N_6070,N_6422);
nand U7211 (N_7211,N_6137,N_6942);
nand U7212 (N_7212,N_6864,N_6174);
or U7213 (N_7213,N_6617,N_6646);
nor U7214 (N_7214,N_6879,N_6695);
or U7215 (N_7215,N_6462,N_6592);
and U7216 (N_7216,N_6595,N_6704);
nor U7217 (N_7217,N_6194,N_6157);
or U7218 (N_7218,N_6504,N_6765);
and U7219 (N_7219,N_6773,N_6267);
or U7220 (N_7220,N_6909,N_6096);
nand U7221 (N_7221,N_6437,N_6213);
and U7222 (N_7222,N_6735,N_6535);
and U7223 (N_7223,N_6022,N_6159);
nor U7224 (N_7224,N_6187,N_6615);
nor U7225 (N_7225,N_6103,N_6986);
nor U7226 (N_7226,N_6938,N_6528);
and U7227 (N_7227,N_6978,N_6601);
nand U7228 (N_7228,N_6421,N_6029);
nand U7229 (N_7229,N_6480,N_6495);
nand U7230 (N_7230,N_6963,N_6193);
nand U7231 (N_7231,N_6623,N_6918);
or U7232 (N_7232,N_6432,N_6846);
or U7233 (N_7233,N_6057,N_6003);
nand U7234 (N_7234,N_6423,N_6006);
or U7235 (N_7235,N_6961,N_6814);
or U7236 (N_7236,N_6890,N_6477);
nand U7237 (N_7237,N_6171,N_6355);
and U7238 (N_7238,N_6688,N_6224);
nor U7239 (N_7239,N_6988,N_6549);
nor U7240 (N_7240,N_6447,N_6730);
nor U7241 (N_7241,N_6899,N_6169);
or U7242 (N_7242,N_6962,N_6831);
nor U7243 (N_7243,N_6780,N_6120);
and U7244 (N_7244,N_6522,N_6276);
nor U7245 (N_7245,N_6954,N_6856);
nand U7246 (N_7246,N_6543,N_6099);
nand U7247 (N_7247,N_6113,N_6259);
and U7248 (N_7248,N_6370,N_6693);
xnor U7249 (N_7249,N_6063,N_6135);
or U7250 (N_7250,N_6991,N_6943);
and U7251 (N_7251,N_6998,N_6458);
nand U7252 (N_7252,N_6048,N_6588);
and U7253 (N_7253,N_6284,N_6497);
and U7254 (N_7254,N_6293,N_6230);
nand U7255 (N_7255,N_6696,N_6037);
and U7256 (N_7256,N_6122,N_6392);
and U7257 (N_7257,N_6594,N_6781);
nor U7258 (N_7258,N_6686,N_6756);
or U7259 (N_7259,N_6067,N_6446);
nand U7260 (N_7260,N_6433,N_6901);
nor U7261 (N_7261,N_6271,N_6502);
and U7262 (N_7262,N_6056,N_6404);
nand U7263 (N_7263,N_6791,N_6252);
and U7264 (N_7264,N_6465,N_6740);
nand U7265 (N_7265,N_6694,N_6920);
nor U7266 (N_7266,N_6985,N_6574);
nor U7267 (N_7267,N_6797,N_6400);
nor U7268 (N_7268,N_6984,N_6999);
nand U7269 (N_7269,N_6941,N_6384);
or U7270 (N_7270,N_6351,N_6500);
and U7271 (N_7271,N_6026,N_6199);
and U7272 (N_7272,N_6343,N_6637);
nand U7273 (N_7273,N_6229,N_6752);
nand U7274 (N_7274,N_6505,N_6517);
nor U7275 (N_7275,N_6164,N_6334);
nand U7276 (N_7276,N_6908,N_6580);
nor U7277 (N_7277,N_6319,N_6712);
nand U7278 (N_7278,N_6716,N_6072);
nand U7279 (N_7279,N_6362,N_6593);
or U7280 (N_7280,N_6205,N_6016);
nand U7281 (N_7281,N_6361,N_6501);
nand U7282 (N_7282,N_6838,N_6069);
or U7283 (N_7283,N_6488,N_6531);
nand U7284 (N_7284,N_6554,N_6530);
nor U7285 (N_7285,N_6402,N_6749);
and U7286 (N_7286,N_6453,N_6117);
or U7287 (N_7287,N_6013,N_6144);
or U7288 (N_7288,N_6743,N_6521);
nor U7289 (N_7289,N_6955,N_6982);
nor U7290 (N_7290,N_6291,N_6380);
nor U7291 (N_7291,N_6093,N_6577);
nand U7292 (N_7292,N_6238,N_6245);
nand U7293 (N_7293,N_6820,N_6610);
nor U7294 (N_7294,N_6398,N_6681);
nand U7295 (N_7295,N_6555,N_6755);
nor U7296 (N_7296,N_6829,N_6406);
and U7297 (N_7297,N_6566,N_6796);
nor U7298 (N_7298,N_6386,N_6902);
nor U7299 (N_7299,N_6925,N_6684);
and U7300 (N_7300,N_6124,N_6803);
or U7301 (N_7301,N_6336,N_6575);
or U7302 (N_7302,N_6449,N_6785);
or U7303 (N_7303,N_6839,N_6150);
or U7304 (N_7304,N_6223,N_6853);
nand U7305 (N_7305,N_6579,N_6008);
nor U7306 (N_7306,N_6967,N_6977);
or U7307 (N_7307,N_6368,N_6275);
nor U7308 (N_7308,N_6761,N_6337);
nand U7309 (N_7309,N_6625,N_6285);
or U7310 (N_7310,N_6509,N_6960);
or U7311 (N_7311,N_6215,N_6478);
or U7312 (N_7312,N_6128,N_6966);
nand U7313 (N_7313,N_6972,N_6387);
nor U7314 (N_7314,N_6633,N_6214);
nor U7315 (N_7315,N_6614,N_6111);
or U7316 (N_7316,N_6653,N_6338);
and U7317 (N_7317,N_6524,N_6051);
nand U7318 (N_7318,N_6758,N_6431);
and U7319 (N_7319,N_6819,N_6345);
and U7320 (N_7320,N_6249,N_6945);
nand U7321 (N_7321,N_6516,N_6990);
and U7322 (N_7322,N_6833,N_6356);
and U7323 (N_7323,N_6790,N_6619);
and U7324 (N_7324,N_6160,N_6685);
and U7325 (N_7325,N_6228,N_6331);
nor U7326 (N_7326,N_6298,N_6073);
xor U7327 (N_7327,N_6408,N_6420);
or U7328 (N_7328,N_6283,N_6843);
nor U7329 (N_7329,N_6676,N_6332);
or U7330 (N_7330,N_6651,N_6824);
or U7331 (N_7331,N_6720,N_6895);
nor U7332 (N_7332,N_6750,N_6556);
and U7333 (N_7333,N_6759,N_6609);
nand U7334 (N_7334,N_6706,N_6198);
nor U7335 (N_7335,N_6114,N_6687);
nor U7336 (N_7336,N_6634,N_6959);
or U7337 (N_7337,N_6151,N_6606);
nor U7338 (N_7338,N_6367,N_6045);
nand U7339 (N_7339,N_6900,N_6565);
or U7340 (N_7340,N_6658,N_6359);
and U7341 (N_7341,N_6935,N_6279);
nor U7342 (N_7342,N_6742,N_6369);
and U7343 (N_7343,N_6946,N_6305);
nand U7344 (N_7344,N_6260,N_6382);
nor U7345 (N_7345,N_6733,N_6881);
nand U7346 (N_7346,N_6264,N_6893);
nor U7347 (N_7347,N_6828,N_6263);
nor U7348 (N_7348,N_6106,N_6299);
nand U7349 (N_7349,N_6203,N_6813);
nand U7350 (N_7350,N_6585,N_6638);
nor U7351 (N_7351,N_6799,N_6777);
nor U7352 (N_7352,N_6888,N_6711);
and U7353 (N_7353,N_6088,N_6286);
nor U7354 (N_7354,N_6657,N_6272);
nor U7355 (N_7355,N_6220,N_6001);
or U7356 (N_7356,N_6241,N_6183);
nor U7357 (N_7357,N_6280,N_6934);
or U7358 (N_7358,N_6865,N_6200);
nand U7359 (N_7359,N_6786,N_6494);
or U7360 (N_7360,N_6697,N_6055);
nor U7361 (N_7361,N_6376,N_6563);
nor U7362 (N_7362,N_6307,N_6763);
nand U7363 (N_7363,N_6871,N_6806);
and U7364 (N_7364,N_6242,N_6239);
or U7365 (N_7365,N_6639,N_6119);
nand U7366 (N_7366,N_6968,N_6217);
or U7367 (N_7367,N_6958,N_6583);
nand U7368 (N_7368,N_6581,N_6683);
or U7369 (N_7369,N_6618,N_6401);
nor U7370 (N_7370,N_6652,N_6032);
and U7371 (N_7371,N_6748,N_6143);
or U7372 (N_7372,N_6470,N_6156);
nor U7373 (N_7373,N_6836,N_6527);
nor U7374 (N_7374,N_6714,N_6123);
and U7375 (N_7375,N_6715,N_6917);
nand U7376 (N_7376,N_6167,N_6928);
nand U7377 (N_7377,N_6304,N_6485);
or U7378 (N_7378,N_6641,N_6744);
nor U7379 (N_7379,N_6288,N_6629);
and U7380 (N_7380,N_6177,N_6185);
xor U7381 (N_7381,N_6798,N_6349);
nor U7382 (N_7382,N_6262,N_6810);
or U7383 (N_7383,N_6534,N_6292);
nor U7384 (N_7384,N_6713,N_6598);
nor U7385 (N_7385,N_6318,N_6605);
nor U7386 (N_7386,N_6168,N_6590);
nand U7387 (N_7387,N_6654,N_6532);
and U7388 (N_7388,N_6040,N_6274);
nor U7389 (N_7389,N_6980,N_6702);
or U7390 (N_7390,N_6584,N_6621);
nand U7391 (N_7391,N_6700,N_6973);
and U7392 (N_7392,N_6788,N_6608);
or U7393 (N_7393,N_6322,N_6570);
or U7394 (N_7394,N_6596,N_6195);
nor U7395 (N_7395,N_6352,N_6269);
nor U7396 (N_7396,N_6208,N_6418);
nor U7397 (N_7397,N_6887,N_6324);
or U7398 (N_7398,N_6058,N_6340);
or U7399 (N_7399,N_6142,N_6466);
nor U7400 (N_7400,N_6479,N_6507);
and U7401 (N_7401,N_6559,N_6483);
nand U7402 (N_7402,N_6471,N_6077);
xor U7403 (N_7403,N_6250,N_6722);
nor U7404 (N_7404,N_6021,N_6499);
or U7405 (N_7405,N_6877,N_6204);
nor U7406 (N_7406,N_6627,N_6163);
nand U7407 (N_7407,N_6883,N_6290);
nand U7408 (N_7408,N_6636,N_6936);
xor U7409 (N_7409,N_6710,N_6541);
nor U7410 (N_7410,N_6832,N_6030);
nor U7411 (N_7411,N_6170,N_6005);
and U7412 (N_7412,N_6644,N_6089);
and U7413 (N_7413,N_6537,N_6287);
or U7414 (N_7414,N_6582,N_6457);
and U7415 (N_7415,N_6842,N_6442);
or U7416 (N_7416,N_6339,N_6586);
or U7417 (N_7417,N_6066,N_6426);
nand U7418 (N_7418,N_6455,N_6366);
and U7419 (N_7419,N_6914,N_6772);
xnor U7420 (N_7420,N_6314,N_6222);
nand U7421 (N_7421,N_6152,N_6869);
or U7422 (N_7422,N_6664,N_6850);
and U7423 (N_7423,N_6414,N_6745);
or U7424 (N_7424,N_6854,N_6732);
or U7425 (N_7425,N_6801,N_6130);
and U7426 (N_7426,N_6518,N_6898);
or U7427 (N_7427,N_6372,N_6023);
nor U7428 (N_7428,N_6100,N_6310);
and U7429 (N_7429,N_6121,N_6859);
nand U7430 (N_7430,N_6131,N_6689);
or U7431 (N_7431,N_6181,N_6000);
or U7432 (N_7432,N_6416,N_6880);
and U7433 (N_7433,N_6905,N_6787);
nor U7434 (N_7434,N_6811,N_6043);
or U7435 (N_7435,N_6079,N_6851);
nand U7436 (N_7436,N_6303,N_6353);
nor U7437 (N_7437,N_6545,N_6161);
or U7438 (N_7438,N_6460,N_6396);
nand U7439 (N_7439,N_6699,N_6514);
nand U7440 (N_7440,N_6753,N_6327);
or U7441 (N_7441,N_6690,N_6931);
nand U7442 (N_7442,N_6551,N_6837);
nand U7443 (N_7443,N_6020,N_6138);
nor U7444 (N_7444,N_6440,N_6894);
nor U7445 (N_7445,N_6461,N_6395);
and U7446 (N_7446,N_6993,N_6640);
or U7447 (N_7447,N_6840,N_6661);
nand U7448 (N_7448,N_6107,N_6519);
nand U7449 (N_7449,N_6892,N_6407);
and U7450 (N_7450,N_6997,N_6847);
nand U7451 (N_7451,N_6254,N_6393);
and U7452 (N_7452,N_6053,N_6347);
or U7453 (N_7453,N_6922,N_6602);
and U7454 (N_7454,N_6717,N_6508);
and U7455 (N_7455,N_6348,N_6613);
and U7456 (N_7456,N_6086,N_6569);
or U7457 (N_7457,N_6571,N_6981);
and U7458 (N_7458,N_6912,N_6815);
and U7459 (N_7459,N_6027,N_6083);
nand U7460 (N_7460,N_6737,N_6940);
and U7461 (N_7461,N_6210,N_6768);
and U7462 (N_7462,N_6861,N_6244);
nor U7463 (N_7463,N_6817,N_6649);
nand U7464 (N_7464,N_6764,N_6992);
nor U7465 (N_7465,N_6932,N_6662);
nand U7466 (N_7466,N_6896,N_6047);
nor U7467 (N_7467,N_6544,N_6139);
and U7468 (N_7468,N_6660,N_6014);
or U7469 (N_7469,N_6526,N_6312);
xnor U7470 (N_7470,N_6476,N_6822);
nand U7471 (N_7471,N_6201,N_6134);
or U7472 (N_7472,N_6335,N_6068);
and U7473 (N_7473,N_6178,N_6512);
nor U7474 (N_7474,N_6484,N_6729);
and U7475 (N_7475,N_6035,N_6867);
and U7476 (N_7476,N_6282,N_6081);
nand U7477 (N_7477,N_6529,N_6818);
or U7478 (N_7478,N_6739,N_6010);
nand U7479 (N_7479,N_6552,N_6328);
or U7480 (N_7480,N_6778,N_6452);
and U7481 (N_7481,N_6975,N_6525);
or U7482 (N_7482,N_6028,N_6553);
and U7483 (N_7483,N_6612,N_6561);
and U7484 (N_7484,N_6949,N_6904);
and U7485 (N_7485,N_6724,N_6947);
or U7486 (N_7486,N_6115,N_6062);
and U7487 (N_7487,N_6599,N_6234);
nor U7488 (N_7488,N_6315,N_6486);
or U7489 (N_7489,N_6092,N_6221);
nor U7490 (N_7490,N_6251,N_6116);
and U7491 (N_7491,N_6147,N_6041);
and U7492 (N_7492,N_6389,N_6626);
and U7493 (N_7493,N_6677,N_6557);
xor U7494 (N_7494,N_6448,N_6236);
nand U7495 (N_7495,N_6105,N_6182);
nor U7496 (N_7496,N_6411,N_6439);
nand U7497 (N_7497,N_6413,N_6767);
nor U7498 (N_7498,N_6172,N_6253);
nor U7499 (N_7499,N_6719,N_6165);
nor U7500 (N_7500,N_6652,N_6495);
nand U7501 (N_7501,N_6893,N_6964);
nand U7502 (N_7502,N_6164,N_6711);
nor U7503 (N_7503,N_6607,N_6414);
or U7504 (N_7504,N_6609,N_6322);
nand U7505 (N_7505,N_6319,N_6803);
nor U7506 (N_7506,N_6451,N_6534);
nand U7507 (N_7507,N_6454,N_6066);
nand U7508 (N_7508,N_6783,N_6673);
nor U7509 (N_7509,N_6673,N_6000);
nand U7510 (N_7510,N_6405,N_6152);
or U7511 (N_7511,N_6738,N_6010);
or U7512 (N_7512,N_6363,N_6200);
nand U7513 (N_7513,N_6847,N_6480);
and U7514 (N_7514,N_6383,N_6527);
nor U7515 (N_7515,N_6385,N_6493);
and U7516 (N_7516,N_6648,N_6903);
or U7517 (N_7517,N_6270,N_6149);
xnor U7518 (N_7518,N_6621,N_6060);
or U7519 (N_7519,N_6002,N_6928);
or U7520 (N_7520,N_6757,N_6454);
nor U7521 (N_7521,N_6202,N_6192);
nand U7522 (N_7522,N_6008,N_6150);
nand U7523 (N_7523,N_6264,N_6303);
or U7524 (N_7524,N_6483,N_6387);
and U7525 (N_7525,N_6128,N_6875);
or U7526 (N_7526,N_6129,N_6506);
and U7527 (N_7527,N_6655,N_6451);
xor U7528 (N_7528,N_6527,N_6676);
or U7529 (N_7529,N_6836,N_6124);
and U7530 (N_7530,N_6732,N_6723);
and U7531 (N_7531,N_6036,N_6100);
nor U7532 (N_7532,N_6449,N_6662);
nor U7533 (N_7533,N_6995,N_6880);
nor U7534 (N_7534,N_6841,N_6641);
and U7535 (N_7535,N_6484,N_6800);
and U7536 (N_7536,N_6105,N_6886);
nor U7537 (N_7537,N_6203,N_6613);
or U7538 (N_7538,N_6874,N_6321);
or U7539 (N_7539,N_6368,N_6454);
and U7540 (N_7540,N_6902,N_6375);
nand U7541 (N_7541,N_6249,N_6125);
and U7542 (N_7542,N_6291,N_6213);
and U7543 (N_7543,N_6483,N_6103);
nor U7544 (N_7544,N_6895,N_6102);
or U7545 (N_7545,N_6853,N_6876);
nand U7546 (N_7546,N_6864,N_6572);
or U7547 (N_7547,N_6165,N_6506);
nand U7548 (N_7548,N_6796,N_6073);
or U7549 (N_7549,N_6145,N_6175);
nor U7550 (N_7550,N_6899,N_6235);
or U7551 (N_7551,N_6893,N_6015);
or U7552 (N_7552,N_6977,N_6746);
nand U7553 (N_7553,N_6593,N_6099);
and U7554 (N_7554,N_6512,N_6279);
nor U7555 (N_7555,N_6483,N_6421);
nor U7556 (N_7556,N_6517,N_6748);
or U7557 (N_7557,N_6363,N_6317);
or U7558 (N_7558,N_6528,N_6590);
nand U7559 (N_7559,N_6507,N_6297);
nor U7560 (N_7560,N_6690,N_6694);
and U7561 (N_7561,N_6873,N_6390);
and U7562 (N_7562,N_6579,N_6806);
nand U7563 (N_7563,N_6120,N_6322);
nor U7564 (N_7564,N_6474,N_6687);
nand U7565 (N_7565,N_6765,N_6752);
nor U7566 (N_7566,N_6747,N_6973);
or U7567 (N_7567,N_6278,N_6133);
nor U7568 (N_7568,N_6541,N_6772);
nor U7569 (N_7569,N_6317,N_6282);
nand U7570 (N_7570,N_6428,N_6790);
nor U7571 (N_7571,N_6446,N_6370);
nor U7572 (N_7572,N_6750,N_6817);
nor U7573 (N_7573,N_6983,N_6567);
and U7574 (N_7574,N_6661,N_6094);
or U7575 (N_7575,N_6404,N_6957);
nand U7576 (N_7576,N_6731,N_6187);
and U7577 (N_7577,N_6823,N_6931);
nor U7578 (N_7578,N_6632,N_6890);
and U7579 (N_7579,N_6661,N_6734);
or U7580 (N_7580,N_6146,N_6358);
or U7581 (N_7581,N_6234,N_6009);
and U7582 (N_7582,N_6695,N_6603);
or U7583 (N_7583,N_6709,N_6715);
xor U7584 (N_7584,N_6053,N_6612);
or U7585 (N_7585,N_6134,N_6953);
and U7586 (N_7586,N_6915,N_6271);
nor U7587 (N_7587,N_6773,N_6548);
nor U7588 (N_7588,N_6552,N_6730);
or U7589 (N_7589,N_6368,N_6143);
or U7590 (N_7590,N_6418,N_6275);
nor U7591 (N_7591,N_6068,N_6109);
or U7592 (N_7592,N_6217,N_6608);
or U7593 (N_7593,N_6939,N_6380);
nand U7594 (N_7594,N_6920,N_6580);
and U7595 (N_7595,N_6120,N_6677);
nand U7596 (N_7596,N_6518,N_6503);
and U7597 (N_7597,N_6592,N_6887);
or U7598 (N_7598,N_6420,N_6349);
nand U7599 (N_7599,N_6069,N_6040);
nor U7600 (N_7600,N_6232,N_6143);
nor U7601 (N_7601,N_6424,N_6252);
nor U7602 (N_7602,N_6176,N_6376);
or U7603 (N_7603,N_6893,N_6445);
nor U7604 (N_7604,N_6647,N_6503);
nor U7605 (N_7605,N_6562,N_6732);
or U7606 (N_7606,N_6065,N_6113);
nor U7607 (N_7607,N_6379,N_6373);
nand U7608 (N_7608,N_6600,N_6636);
or U7609 (N_7609,N_6177,N_6730);
nor U7610 (N_7610,N_6204,N_6520);
nand U7611 (N_7611,N_6303,N_6739);
nand U7612 (N_7612,N_6184,N_6709);
or U7613 (N_7613,N_6302,N_6392);
and U7614 (N_7614,N_6056,N_6707);
and U7615 (N_7615,N_6040,N_6476);
or U7616 (N_7616,N_6456,N_6166);
or U7617 (N_7617,N_6547,N_6047);
nor U7618 (N_7618,N_6635,N_6288);
nor U7619 (N_7619,N_6022,N_6391);
and U7620 (N_7620,N_6223,N_6886);
nand U7621 (N_7621,N_6056,N_6158);
nand U7622 (N_7622,N_6829,N_6699);
and U7623 (N_7623,N_6427,N_6628);
or U7624 (N_7624,N_6223,N_6850);
and U7625 (N_7625,N_6673,N_6439);
nand U7626 (N_7626,N_6704,N_6788);
nand U7627 (N_7627,N_6943,N_6319);
and U7628 (N_7628,N_6892,N_6139);
nand U7629 (N_7629,N_6497,N_6718);
xnor U7630 (N_7630,N_6350,N_6635);
or U7631 (N_7631,N_6062,N_6749);
xnor U7632 (N_7632,N_6196,N_6707);
nand U7633 (N_7633,N_6278,N_6535);
or U7634 (N_7634,N_6699,N_6936);
nand U7635 (N_7635,N_6455,N_6206);
nand U7636 (N_7636,N_6918,N_6941);
nor U7637 (N_7637,N_6021,N_6404);
or U7638 (N_7638,N_6740,N_6479);
nand U7639 (N_7639,N_6703,N_6152);
nor U7640 (N_7640,N_6943,N_6439);
or U7641 (N_7641,N_6811,N_6050);
nor U7642 (N_7642,N_6177,N_6269);
nand U7643 (N_7643,N_6725,N_6555);
and U7644 (N_7644,N_6915,N_6149);
and U7645 (N_7645,N_6395,N_6700);
and U7646 (N_7646,N_6775,N_6456);
nand U7647 (N_7647,N_6780,N_6665);
nand U7648 (N_7648,N_6909,N_6715);
and U7649 (N_7649,N_6856,N_6971);
and U7650 (N_7650,N_6098,N_6423);
and U7651 (N_7651,N_6990,N_6623);
and U7652 (N_7652,N_6151,N_6627);
or U7653 (N_7653,N_6905,N_6227);
nor U7654 (N_7654,N_6546,N_6858);
or U7655 (N_7655,N_6940,N_6419);
nor U7656 (N_7656,N_6205,N_6424);
and U7657 (N_7657,N_6483,N_6948);
or U7658 (N_7658,N_6425,N_6770);
nand U7659 (N_7659,N_6861,N_6199);
nor U7660 (N_7660,N_6792,N_6491);
or U7661 (N_7661,N_6440,N_6168);
and U7662 (N_7662,N_6687,N_6700);
or U7663 (N_7663,N_6168,N_6844);
nor U7664 (N_7664,N_6955,N_6462);
nand U7665 (N_7665,N_6998,N_6726);
nor U7666 (N_7666,N_6498,N_6532);
nand U7667 (N_7667,N_6303,N_6050);
nor U7668 (N_7668,N_6084,N_6920);
or U7669 (N_7669,N_6786,N_6405);
nor U7670 (N_7670,N_6559,N_6358);
and U7671 (N_7671,N_6636,N_6998);
or U7672 (N_7672,N_6062,N_6697);
and U7673 (N_7673,N_6732,N_6669);
nor U7674 (N_7674,N_6151,N_6888);
nand U7675 (N_7675,N_6389,N_6451);
nand U7676 (N_7676,N_6337,N_6891);
nor U7677 (N_7677,N_6007,N_6569);
and U7678 (N_7678,N_6241,N_6962);
nand U7679 (N_7679,N_6220,N_6838);
and U7680 (N_7680,N_6369,N_6020);
and U7681 (N_7681,N_6015,N_6558);
nor U7682 (N_7682,N_6450,N_6632);
nand U7683 (N_7683,N_6806,N_6041);
or U7684 (N_7684,N_6118,N_6558);
or U7685 (N_7685,N_6948,N_6595);
or U7686 (N_7686,N_6835,N_6598);
nor U7687 (N_7687,N_6158,N_6623);
nor U7688 (N_7688,N_6722,N_6783);
nor U7689 (N_7689,N_6865,N_6825);
and U7690 (N_7690,N_6253,N_6426);
or U7691 (N_7691,N_6547,N_6515);
nor U7692 (N_7692,N_6799,N_6967);
and U7693 (N_7693,N_6673,N_6598);
and U7694 (N_7694,N_6992,N_6032);
or U7695 (N_7695,N_6618,N_6456);
nand U7696 (N_7696,N_6615,N_6938);
and U7697 (N_7697,N_6448,N_6429);
and U7698 (N_7698,N_6221,N_6341);
and U7699 (N_7699,N_6445,N_6405);
and U7700 (N_7700,N_6755,N_6144);
nor U7701 (N_7701,N_6918,N_6482);
xnor U7702 (N_7702,N_6538,N_6627);
or U7703 (N_7703,N_6369,N_6804);
nand U7704 (N_7704,N_6746,N_6810);
or U7705 (N_7705,N_6820,N_6927);
nand U7706 (N_7706,N_6235,N_6204);
or U7707 (N_7707,N_6027,N_6589);
and U7708 (N_7708,N_6078,N_6404);
nand U7709 (N_7709,N_6539,N_6884);
nand U7710 (N_7710,N_6940,N_6501);
nand U7711 (N_7711,N_6321,N_6172);
and U7712 (N_7712,N_6437,N_6028);
and U7713 (N_7713,N_6547,N_6509);
nand U7714 (N_7714,N_6143,N_6950);
or U7715 (N_7715,N_6235,N_6621);
and U7716 (N_7716,N_6624,N_6643);
nand U7717 (N_7717,N_6233,N_6149);
or U7718 (N_7718,N_6933,N_6525);
nor U7719 (N_7719,N_6919,N_6156);
and U7720 (N_7720,N_6498,N_6787);
nand U7721 (N_7721,N_6191,N_6157);
nand U7722 (N_7722,N_6851,N_6397);
or U7723 (N_7723,N_6753,N_6577);
or U7724 (N_7724,N_6194,N_6444);
nor U7725 (N_7725,N_6047,N_6479);
nand U7726 (N_7726,N_6255,N_6207);
nor U7727 (N_7727,N_6790,N_6543);
nand U7728 (N_7728,N_6349,N_6407);
and U7729 (N_7729,N_6560,N_6419);
and U7730 (N_7730,N_6142,N_6834);
nor U7731 (N_7731,N_6657,N_6308);
and U7732 (N_7732,N_6442,N_6563);
xnor U7733 (N_7733,N_6872,N_6919);
nor U7734 (N_7734,N_6488,N_6445);
nand U7735 (N_7735,N_6365,N_6207);
and U7736 (N_7736,N_6608,N_6514);
nand U7737 (N_7737,N_6313,N_6505);
nand U7738 (N_7738,N_6650,N_6054);
or U7739 (N_7739,N_6355,N_6287);
or U7740 (N_7740,N_6821,N_6493);
nand U7741 (N_7741,N_6579,N_6336);
nand U7742 (N_7742,N_6801,N_6085);
nand U7743 (N_7743,N_6253,N_6096);
and U7744 (N_7744,N_6428,N_6055);
nand U7745 (N_7745,N_6913,N_6923);
and U7746 (N_7746,N_6393,N_6200);
and U7747 (N_7747,N_6282,N_6973);
and U7748 (N_7748,N_6564,N_6105);
nor U7749 (N_7749,N_6279,N_6941);
nand U7750 (N_7750,N_6003,N_6680);
nor U7751 (N_7751,N_6222,N_6947);
and U7752 (N_7752,N_6081,N_6052);
and U7753 (N_7753,N_6871,N_6465);
and U7754 (N_7754,N_6664,N_6151);
nor U7755 (N_7755,N_6233,N_6660);
and U7756 (N_7756,N_6262,N_6582);
or U7757 (N_7757,N_6137,N_6441);
and U7758 (N_7758,N_6767,N_6193);
nand U7759 (N_7759,N_6824,N_6534);
or U7760 (N_7760,N_6480,N_6283);
nor U7761 (N_7761,N_6142,N_6525);
nor U7762 (N_7762,N_6265,N_6166);
nand U7763 (N_7763,N_6801,N_6087);
or U7764 (N_7764,N_6420,N_6075);
nand U7765 (N_7765,N_6368,N_6768);
and U7766 (N_7766,N_6204,N_6341);
or U7767 (N_7767,N_6493,N_6864);
nand U7768 (N_7768,N_6001,N_6616);
nor U7769 (N_7769,N_6256,N_6621);
and U7770 (N_7770,N_6011,N_6370);
and U7771 (N_7771,N_6522,N_6489);
nand U7772 (N_7772,N_6134,N_6518);
nand U7773 (N_7773,N_6865,N_6765);
and U7774 (N_7774,N_6042,N_6641);
nand U7775 (N_7775,N_6173,N_6476);
nand U7776 (N_7776,N_6534,N_6218);
and U7777 (N_7777,N_6631,N_6767);
and U7778 (N_7778,N_6595,N_6943);
or U7779 (N_7779,N_6563,N_6807);
or U7780 (N_7780,N_6372,N_6032);
nand U7781 (N_7781,N_6888,N_6624);
and U7782 (N_7782,N_6348,N_6337);
nor U7783 (N_7783,N_6779,N_6087);
nor U7784 (N_7784,N_6029,N_6146);
and U7785 (N_7785,N_6441,N_6756);
nor U7786 (N_7786,N_6034,N_6858);
and U7787 (N_7787,N_6368,N_6614);
nor U7788 (N_7788,N_6385,N_6679);
or U7789 (N_7789,N_6885,N_6488);
or U7790 (N_7790,N_6889,N_6176);
nand U7791 (N_7791,N_6978,N_6546);
nand U7792 (N_7792,N_6140,N_6925);
or U7793 (N_7793,N_6447,N_6117);
nand U7794 (N_7794,N_6938,N_6713);
nor U7795 (N_7795,N_6744,N_6177);
xnor U7796 (N_7796,N_6419,N_6475);
nor U7797 (N_7797,N_6560,N_6820);
nand U7798 (N_7798,N_6119,N_6672);
or U7799 (N_7799,N_6099,N_6957);
nor U7800 (N_7800,N_6303,N_6068);
and U7801 (N_7801,N_6526,N_6710);
nor U7802 (N_7802,N_6490,N_6693);
or U7803 (N_7803,N_6590,N_6122);
or U7804 (N_7804,N_6769,N_6081);
and U7805 (N_7805,N_6321,N_6149);
and U7806 (N_7806,N_6440,N_6386);
nand U7807 (N_7807,N_6065,N_6523);
nor U7808 (N_7808,N_6344,N_6569);
nand U7809 (N_7809,N_6059,N_6635);
nor U7810 (N_7810,N_6659,N_6614);
nand U7811 (N_7811,N_6254,N_6917);
or U7812 (N_7812,N_6195,N_6470);
and U7813 (N_7813,N_6249,N_6762);
or U7814 (N_7814,N_6980,N_6277);
and U7815 (N_7815,N_6934,N_6116);
or U7816 (N_7816,N_6995,N_6303);
nor U7817 (N_7817,N_6182,N_6312);
and U7818 (N_7818,N_6601,N_6255);
or U7819 (N_7819,N_6546,N_6539);
nand U7820 (N_7820,N_6926,N_6157);
nand U7821 (N_7821,N_6165,N_6027);
nor U7822 (N_7822,N_6909,N_6666);
nor U7823 (N_7823,N_6327,N_6914);
and U7824 (N_7824,N_6976,N_6742);
and U7825 (N_7825,N_6160,N_6279);
and U7826 (N_7826,N_6426,N_6592);
or U7827 (N_7827,N_6943,N_6733);
or U7828 (N_7828,N_6631,N_6931);
nand U7829 (N_7829,N_6840,N_6109);
or U7830 (N_7830,N_6260,N_6302);
or U7831 (N_7831,N_6805,N_6130);
nor U7832 (N_7832,N_6733,N_6919);
nor U7833 (N_7833,N_6843,N_6256);
or U7834 (N_7834,N_6588,N_6736);
nand U7835 (N_7835,N_6851,N_6461);
and U7836 (N_7836,N_6913,N_6424);
and U7837 (N_7837,N_6675,N_6607);
nand U7838 (N_7838,N_6675,N_6586);
and U7839 (N_7839,N_6133,N_6537);
nor U7840 (N_7840,N_6181,N_6603);
nand U7841 (N_7841,N_6854,N_6506);
nand U7842 (N_7842,N_6772,N_6277);
or U7843 (N_7843,N_6565,N_6886);
nor U7844 (N_7844,N_6569,N_6751);
or U7845 (N_7845,N_6759,N_6100);
nor U7846 (N_7846,N_6478,N_6398);
nor U7847 (N_7847,N_6787,N_6264);
and U7848 (N_7848,N_6178,N_6700);
or U7849 (N_7849,N_6167,N_6756);
nand U7850 (N_7850,N_6132,N_6427);
and U7851 (N_7851,N_6009,N_6166);
or U7852 (N_7852,N_6034,N_6425);
nand U7853 (N_7853,N_6039,N_6231);
or U7854 (N_7854,N_6962,N_6501);
nand U7855 (N_7855,N_6745,N_6475);
or U7856 (N_7856,N_6900,N_6211);
nand U7857 (N_7857,N_6276,N_6067);
or U7858 (N_7858,N_6999,N_6431);
nand U7859 (N_7859,N_6230,N_6950);
nor U7860 (N_7860,N_6264,N_6855);
nor U7861 (N_7861,N_6825,N_6150);
nor U7862 (N_7862,N_6912,N_6965);
nand U7863 (N_7863,N_6998,N_6461);
nor U7864 (N_7864,N_6077,N_6685);
nand U7865 (N_7865,N_6202,N_6008);
nor U7866 (N_7866,N_6810,N_6235);
and U7867 (N_7867,N_6504,N_6216);
and U7868 (N_7868,N_6945,N_6595);
nor U7869 (N_7869,N_6773,N_6714);
or U7870 (N_7870,N_6783,N_6477);
nor U7871 (N_7871,N_6282,N_6690);
xnor U7872 (N_7872,N_6581,N_6342);
or U7873 (N_7873,N_6398,N_6464);
nand U7874 (N_7874,N_6980,N_6521);
or U7875 (N_7875,N_6935,N_6074);
and U7876 (N_7876,N_6697,N_6849);
or U7877 (N_7877,N_6074,N_6955);
nor U7878 (N_7878,N_6165,N_6212);
or U7879 (N_7879,N_6730,N_6726);
or U7880 (N_7880,N_6091,N_6912);
nor U7881 (N_7881,N_6398,N_6688);
nor U7882 (N_7882,N_6061,N_6934);
and U7883 (N_7883,N_6096,N_6829);
and U7884 (N_7884,N_6244,N_6694);
or U7885 (N_7885,N_6501,N_6014);
and U7886 (N_7886,N_6427,N_6336);
nor U7887 (N_7887,N_6480,N_6448);
and U7888 (N_7888,N_6916,N_6526);
nor U7889 (N_7889,N_6641,N_6162);
nand U7890 (N_7890,N_6790,N_6942);
nor U7891 (N_7891,N_6463,N_6573);
nor U7892 (N_7892,N_6619,N_6487);
and U7893 (N_7893,N_6000,N_6193);
and U7894 (N_7894,N_6583,N_6691);
nand U7895 (N_7895,N_6034,N_6510);
nor U7896 (N_7896,N_6675,N_6037);
and U7897 (N_7897,N_6723,N_6186);
nor U7898 (N_7898,N_6569,N_6099);
nor U7899 (N_7899,N_6782,N_6546);
nor U7900 (N_7900,N_6414,N_6070);
nand U7901 (N_7901,N_6299,N_6989);
and U7902 (N_7902,N_6760,N_6113);
or U7903 (N_7903,N_6473,N_6465);
nand U7904 (N_7904,N_6399,N_6101);
nor U7905 (N_7905,N_6008,N_6688);
nand U7906 (N_7906,N_6865,N_6778);
and U7907 (N_7907,N_6956,N_6899);
or U7908 (N_7908,N_6877,N_6977);
nand U7909 (N_7909,N_6506,N_6963);
nand U7910 (N_7910,N_6260,N_6965);
nand U7911 (N_7911,N_6036,N_6149);
and U7912 (N_7912,N_6302,N_6305);
nand U7913 (N_7913,N_6759,N_6812);
nand U7914 (N_7914,N_6407,N_6724);
xor U7915 (N_7915,N_6262,N_6191);
or U7916 (N_7916,N_6760,N_6252);
and U7917 (N_7917,N_6023,N_6406);
and U7918 (N_7918,N_6143,N_6762);
or U7919 (N_7919,N_6705,N_6096);
nor U7920 (N_7920,N_6561,N_6816);
nand U7921 (N_7921,N_6469,N_6615);
nor U7922 (N_7922,N_6688,N_6517);
or U7923 (N_7923,N_6625,N_6187);
nand U7924 (N_7924,N_6481,N_6390);
and U7925 (N_7925,N_6056,N_6530);
nand U7926 (N_7926,N_6892,N_6330);
and U7927 (N_7927,N_6090,N_6368);
or U7928 (N_7928,N_6092,N_6505);
and U7929 (N_7929,N_6188,N_6394);
nor U7930 (N_7930,N_6654,N_6087);
nor U7931 (N_7931,N_6171,N_6494);
nand U7932 (N_7932,N_6560,N_6008);
and U7933 (N_7933,N_6035,N_6545);
and U7934 (N_7934,N_6409,N_6227);
nor U7935 (N_7935,N_6552,N_6424);
nor U7936 (N_7936,N_6203,N_6321);
nor U7937 (N_7937,N_6372,N_6449);
and U7938 (N_7938,N_6210,N_6469);
nand U7939 (N_7939,N_6401,N_6689);
nand U7940 (N_7940,N_6295,N_6935);
or U7941 (N_7941,N_6384,N_6303);
nand U7942 (N_7942,N_6626,N_6147);
and U7943 (N_7943,N_6263,N_6539);
and U7944 (N_7944,N_6352,N_6735);
or U7945 (N_7945,N_6351,N_6599);
and U7946 (N_7946,N_6836,N_6878);
and U7947 (N_7947,N_6808,N_6539);
and U7948 (N_7948,N_6872,N_6655);
nor U7949 (N_7949,N_6481,N_6685);
and U7950 (N_7950,N_6843,N_6076);
nor U7951 (N_7951,N_6464,N_6541);
or U7952 (N_7952,N_6945,N_6398);
and U7953 (N_7953,N_6114,N_6303);
xor U7954 (N_7954,N_6593,N_6143);
or U7955 (N_7955,N_6177,N_6845);
and U7956 (N_7956,N_6097,N_6649);
nor U7957 (N_7957,N_6620,N_6628);
nand U7958 (N_7958,N_6049,N_6179);
or U7959 (N_7959,N_6073,N_6923);
nand U7960 (N_7960,N_6389,N_6851);
or U7961 (N_7961,N_6430,N_6486);
or U7962 (N_7962,N_6036,N_6250);
or U7963 (N_7963,N_6333,N_6591);
or U7964 (N_7964,N_6532,N_6417);
and U7965 (N_7965,N_6328,N_6789);
nor U7966 (N_7966,N_6189,N_6201);
nand U7967 (N_7967,N_6694,N_6519);
or U7968 (N_7968,N_6673,N_6397);
or U7969 (N_7969,N_6378,N_6673);
or U7970 (N_7970,N_6345,N_6691);
nor U7971 (N_7971,N_6974,N_6334);
or U7972 (N_7972,N_6639,N_6792);
and U7973 (N_7973,N_6559,N_6874);
nor U7974 (N_7974,N_6181,N_6223);
or U7975 (N_7975,N_6914,N_6048);
nor U7976 (N_7976,N_6577,N_6436);
and U7977 (N_7977,N_6431,N_6516);
nor U7978 (N_7978,N_6192,N_6578);
or U7979 (N_7979,N_6867,N_6327);
nand U7980 (N_7980,N_6680,N_6416);
or U7981 (N_7981,N_6858,N_6060);
nor U7982 (N_7982,N_6060,N_6219);
nand U7983 (N_7983,N_6408,N_6557);
or U7984 (N_7984,N_6585,N_6237);
nand U7985 (N_7985,N_6558,N_6895);
nor U7986 (N_7986,N_6129,N_6932);
nor U7987 (N_7987,N_6238,N_6180);
nor U7988 (N_7988,N_6802,N_6928);
and U7989 (N_7989,N_6866,N_6917);
and U7990 (N_7990,N_6813,N_6038);
and U7991 (N_7991,N_6953,N_6703);
nand U7992 (N_7992,N_6844,N_6834);
nor U7993 (N_7993,N_6280,N_6296);
and U7994 (N_7994,N_6980,N_6426);
or U7995 (N_7995,N_6158,N_6833);
or U7996 (N_7996,N_6612,N_6493);
or U7997 (N_7997,N_6962,N_6068);
nor U7998 (N_7998,N_6346,N_6500);
and U7999 (N_7999,N_6560,N_6188);
nor U8000 (N_8000,N_7508,N_7707);
or U8001 (N_8001,N_7908,N_7644);
nor U8002 (N_8002,N_7536,N_7299);
or U8003 (N_8003,N_7065,N_7492);
or U8004 (N_8004,N_7434,N_7360);
nor U8005 (N_8005,N_7342,N_7616);
nor U8006 (N_8006,N_7645,N_7481);
nand U8007 (N_8007,N_7449,N_7829);
nor U8008 (N_8008,N_7384,N_7767);
nand U8009 (N_8009,N_7049,N_7109);
and U8010 (N_8010,N_7812,N_7361);
nand U8011 (N_8011,N_7529,N_7665);
or U8012 (N_8012,N_7824,N_7994);
nor U8013 (N_8013,N_7674,N_7501);
nor U8014 (N_8014,N_7455,N_7175);
nor U8015 (N_8015,N_7459,N_7278);
or U8016 (N_8016,N_7060,N_7474);
nand U8017 (N_8017,N_7599,N_7298);
or U8018 (N_8018,N_7652,N_7901);
or U8019 (N_8019,N_7123,N_7098);
nor U8020 (N_8020,N_7122,N_7348);
nor U8021 (N_8021,N_7408,N_7965);
and U8022 (N_8022,N_7376,N_7976);
nand U8023 (N_8023,N_7225,N_7437);
nor U8024 (N_8024,N_7654,N_7717);
nand U8025 (N_8025,N_7914,N_7280);
or U8026 (N_8026,N_7683,N_7450);
nor U8027 (N_8027,N_7176,N_7843);
nor U8028 (N_8028,N_7062,N_7261);
nor U8029 (N_8029,N_7152,N_7135);
and U8030 (N_8030,N_7833,N_7378);
nand U8031 (N_8031,N_7301,N_7485);
nand U8032 (N_8032,N_7722,N_7945);
nand U8033 (N_8033,N_7798,N_7682);
or U8034 (N_8034,N_7518,N_7887);
and U8035 (N_8035,N_7334,N_7258);
nand U8036 (N_8036,N_7647,N_7712);
or U8037 (N_8037,N_7364,N_7149);
and U8038 (N_8038,N_7007,N_7130);
and U8039 (N_8039,N_7684,N_7369);
nor U8040 (N_8040,N_7776,N_7004);
nand U8041 (N_8041,N_7181,N_7643);
and U8042 (N_8042,N_7605,N_7351);
nor U8043 (N_8043,N_7442,N_7942);
nand U8044 (N_8044,N_7509,N_7451);
or U8045 (N_8045,N_7831,N_7753);
nand U8046 (N_8046,N_7297,N_7467);
and U8047 (N_8047,N_7472,N_7483);
or U8048 (N_8048,N_7563,N_7055);
and U8049 (N_8049,N_7448,N_7465);
nor U8050 (N_8050,N_7441,N_7533);
nor U8051 (N_8051,N_7872,N_7346);
and U8052 (N_8052,N_7096,N_7950);
and U8053 (N_8053,N_7866,N_7341);
and U8054 (N_8054,N_7039,N_7074);
or U8055 (N_8055,N_7736,N_7354);
nand U8056 (N_8056,N_7457,N_7191);
nand U8057 (N_8057,N_7575,N_7745);
nor U8058 (N_8058,N_7419,N_7819);
nand U8059 (N_8059,N_7580,N_7940);
or U8060 (N_8060,N_7597,N_7446);
nor U8061 (N_8061,N_7761,N_7876);
nand U8062 (N_8062,N_7784,N_7325);
nor U8063 (N_8063,N_7841,N_7358);
nand U8064 (N_8064,N_7579,N_7964);
or U8065 (N_8065,N_7105,N_7461);
or U8066 (N_8066,N_7005,N_7430);
nor U8067 (N_8067,N_7547,N_7813);
and U8068 (N_8068,N_7852,N_7912);
nor U8069 (N_8069,N_7303,N_7290);
nand U8070 (N_8070,N_7087,N_7828);
nand U8071 (N_8071,N_7083,N_7827);
or U8072 (N_8072,N_7853,N_7101);
or U8073 (N_8073,N_7700,N_7246);
and U8074 (N_8074,N_7751,N_7935);
or U8075 (N_8075,N_7770,N_7304);
and U8076 (N_8076,N_7171,N_7830);
nand U8077 (N_8077,N_7642,N_7242);
or U8078 (N_8078,N_7691,N_7400);
nor U8079 (N_8079,N_7545,N_7047);
nor U8080 (N_8080,N_7765,N_7661);
and U8081 (N_8081,N_7424,N_7092);
nand U8082 (N_8082,N_7061,N_7207);
or U8083 (N_8083,N_7911,N_7601);
xor U8084 (N_8084,N_7374,N_7425);
nand U8085 (N_8085,N_7633,N_7045);
and U8086 (N_8086,N_7054,N_7411);
and U8087 (N_8087,N_7962,N_7118);
nor U8088 (N_8088,N_7561,N_7470);
xor U8089 (N_8089,N_7755,N_7956);
nor U8090 (N_8090,N_7287,N_7627);
nand U8091 (N_8091,N_7114,N_7532);
and U8092 (N_8092,N_7131,N_7581);
or U8093 (N_8093,N_7918,N_7163);
nand U8094 (N_8094,N_7495,N_7702);
and U8095 (N_8095,N_7133,N_7903);
nand U8096 (N_8096,N_7398,N_7650);
and U8097 (N_8097,N_7069,N_7775);
nand U8098 (N_8098,N_7452,N_7143);
or U8099 (N_8099,N_7615,N_7228);
and U8100 (N_8100,N_7933,N_7145);
and U8101 (N_8101,N_7955,N_7139);
or U8102 (N_8102,N_7531,N_7931);
nor U8103 (N_8103,N_7733,N_7677);
nor U8104 (N_8104,N_7631,N_7924);
nor U8105 (N_8105,N_7182,N_7944);
nand U8106 (N_8106,N_7111,N_7002);
or U8107 (N_8107,N_7428,N_7453);
or U8108 (N_8108,N_7013,N_7844);
nor U8109 (N_8109,N_7479,N_7790);
and U8110 (N_8110,N_7574,N_7116);
or U8111 (N_8111,N_7210,N_7797);
nor U8112 (N_8112,N_7542,N_7205);
nand U8113 (N_8113,N_7867,N_7778);
or U8114 (N_8114,N_7059,N_7134);
or U8115 (N_8115,N_7110,N_7953);
nand U8116 (N_8116,N_7715,N_7128);
xnor U8117 (N_8117,N_7774,N_7332);
and U8118 (N_8118,N_7626,N_7727);
nand U8119 (N_8119,N_7880,N_7477);
nor U8120 (N_8120,N_7008,N_7443);
or U8121 (N_8121,N_7392,N_7796);
or U8122 (N_8122,N_7347,N_7390);
and U8123 (N_8123,N_7629,N_7198);
nor U8124 (N_8124,N_7578,N_7126);
nand U8125 (N_8125,N_7664,N_7362);
and U8126 (N_8126,N_7502,N_7638);
and U8127 (N_8127,N_7077,N_7668);
or U8128 (N_8128,N_7865,N_7373);
or U8129 (N_8129,N_7789,N_7612);
nor U8130 (N_8130,N_7585,N_7241);
nor U8131 (N_8131,N_7276,N_7388);
nor U8132 (N_8132,N_7602,N_7153);
nand U8133 (N_8133,N_7413,N_7517);
nor U8134 (N_8134,N_7310,N_7167);
and U8135 (N_8135,N_7566,N_7150);
nor U8136 (N_8136,N_7040,N_7669);
nor U8137 (N_8137,N_7544,N_7913);
and U8138 (N_8138,N_7019,N_7211);
or U8139 (N_8139,N_7394,N_7187);
and U8140 (N_8140,N_7357,N_7735);
or U8141 (N_8141,N_7571,N_7878);
nor U8142 (N_8142,N_7267,N_7857);
or U8143 (N_8143,N_7487,N_7995);
or U8144 (N_8144,N_7052,N_7260);
or U8145 (N_8145,N_7811,N_7064);
or U8146 (N_8146,N_7845,N_7078);
nand U8147 (N_8147,N_7537,N_7024);
nor U8148 (N_8148,N_7314,N_7899);
nor U8149 (N_8149,N_7174,N_7368);
nand U8150 (N_8150,N_7404,N_7917);
nor U8151 (N_8151,N_7510,N_7317);
nand U8152 (N_8152,N_7838,N_7277);
nor U8153 (N_8153,N_7800,N_7099);
nand U8154 (N_8154,N_7941,N_7618);
nor U8155 (N_8155,N_7226,N_7009);
and U8156 (N_8156,N_7598,N_7649);
or U8157 (N_8157,N_7249,N_7195);
xnor U8158 (N_8158,N_7726,N_7673);
and U8159 (N_8159,N_7929,N_7016);
and U8160 (N_8160,N_7244,N_7904);
or U8161 (N_8161,N_7666,N_7340);
nor U8162 (N_8162,N_7766,N_7791);
or U8163 (N_8163,N_7081,N_7902);
nand U8164 (N_8164,N_7939,N_7273);
or U8165 (N_8165,N_7527,N_7621);
and U8166 (N_8166,N_7706,N_7910);
nor U8167 (N_8167,N_7391,N_7719);
or U8168 (N_8168,N_7926,N_7234);
or U8169 (N_8169,N_7383,N_7137);
and U8170 (N_8170,N_7604,N_7403);
and U8171 (N_8171,N_7639,N_7560);
or U8172 (N_8172,N_7456,N_7557);
nand U8173 (N_8173,N_7180,N_7498);
or U8174 (N_8174,N_7316,N_7309);
or U8175 (N_8175,N_7091,N_7406);
nand U8176 (N_8176,N_7164,N_7259);
and U8177 (N_8177,N_7822,N_7991);
or U8178 (N_8178,N_7895,N_7967);
nor U8179 (N_8179,N_7037,N_7250);
or U8180 (N_8180,N_7792,N_7603);
and U8181 (N_8181,N_7846,N_7795);
nor U8182 (N_8182,N_7363,N_7355);
or U8183 (N_8183,N_7708,N_7240);
nor U8184 (N_8184,N_7885,N_7286);
nand U8185 (N_8185,N_7562,N_7782);
or U8186 (N_8186,N_7659,N_7239);
nor U8187 (N_8187,N_7178,N_7971);
or U8188 (N_8188,N_7500,N_7594);
and U8189 (N_8189,N_7608,N_7840);
nor U8190 (N_8190,N_7539,N_7206);
nor U8191 (N_8191,N_7113,N_7970);
or U8192 (N_8192,N_7805,N_7610);
nor U8193 (N_8193,N_7697,N_7407);
and U8194 (N_8194,N_7720,N_7086);
and U8195 (N_8195,N_7530,N_7628);
or U8196 (N_8196,N_7252,N_7035);
nand U8197 (N_8197,N_7658,N_7980);
nand U8198 (N_8198,N_7826,N_7284);
nor U8199 (N_8199,N_7193,N_7236);
nor U8200 (N_8200,N_7888,N_7714);
and U8201 (N_8201,N_7809,N_7352);
and U8202 (N_8202,N_7979,N_7093);
nor U8203 (N_8203,N_7963,N_7385);
nand U8204 (N_8204,N_7146,N_7716);
and U8205 (N_8205,N_7046,N_7184);
or U8206 (N_8206,N_7972,N_7932);
nand U8207 (N_8207,N_7022,N_7353);
nor U8208 (N_8208,N_7762,N_7523);
nor U8209 (N_8209,N_7670,N_7288);
or U8210 (N_8210,N_7999,N_7414);
and U8211 (N_8211,N_7337,N_7613);
or U8212 (N_8212,N_7395,N_7693);
and U8213 (N_8213,N_7033,N_7333);
or U8214 (N_8214,N_7835,N_7094);
and U8215 (N_8215,N_7738,N_7151);
and U8216 (N_8216,N_7179,N_7213);
or U8217 (N_8217,N_7891,N_7640);
or U8218 (N_8218,N_7127,N_7998);
or U8219 (N_8219,N_7773,N_7512);
and U8220 (N_8220,N_7366,N_7922);
and U8221 (N_8221,N_7282,N_7711);
and U8222 (N_8222,N_7051,N_7102);
nor U8223 (N_8223,N_7582,N_7189);
nor U8224 (N_8224,N_7936,N_7412);
or U8225 (N_8225,N_7973,N_7896);
nor U8226 (N_8226,N_7919,N_7739);
or U8227 (N_8227,N_7982,N_7464);
nand U8228 (N_8228,N_7737,N_7272);
or U8229 (N_8229,N_7769,N_7921);
and U8230 (N_8230,N_7806,N_7641);
nand U8231 (N_8231,N_7987,N_7511);
and U8232 (N_8232,N_7196,N_7505);
or U8233 (N_8233,N_7928,N_7943);
nand U8234 (N_8234,N_7281,N_7787);
and U8235 (N_8235,N_7625,N_7496);
nand U8236 (N_8236,N_7006,N_7817);
nor U8237 (N_8237,N_7072,N_7522);
nand U8238 (N_8238,N_7981,N_7854);
nor U8239 (N_8239,N_7156,N_7012);
nor U8240 (N_8240,N_7723,N_7731);
or U8241 (N_8241,N_7148,N_7832);
and U8242 (N_8242,N_7201,N_7185);
nand U8243 (N_8243,N_7001,N_7961);
and U8244 (N_8244,N_7836,N_7025);
nand U8245 (N_8245,N_7313,N_7401);
nand U8246 (N_8246,N_7144,N_7433);
and U8247 (N_8247,N_7418,N_7721);
nor U8248 (N_8248,N_7576,N_7021);
or U8249 (N_8249,N_7785,N_7690);
or U8250 (N_8250,N_7068,N_7324);
and U8251 (N_8251,N_7820,N_7458);
or U8252 (N_8252,N_7084,N_7382);
and U8253 (N_8253,N_7513,N_7538);
or U8254 (N_8254,N_7043,N_7744);
or U8255 (N_8255,N_7592,N_7223);
or U8256 (N_8256,N_7938,N_7516);
nor U8257 (N_8257,N_7473,N_7356);
nor U8258 (N_8258,N_7154,N_7426);
nor U8259 (N_8259,N_7554,N_7906);
and U8260 (N_8260,N_7847,N_7044);
nor U8261 (N_8261,N_7937,N_7491);
nor U8262 (N_8262,N_7793,N_7480);
or U8263 (N_8263,N_7494,N_7889);
nor U8264 (N_8264,N_7851,N_7296);
nand U8265 (N_8265,N_7555,N_7230);
nor U8266 (N_8266,N_7947,N_7088);
nand U8267 (N_8267,N_7816,N_7588);
and U8268 (N_8268,N_7989,N_7689);
nand U8269 (N_8269,N_7370,N_7015);
nor U8270 (N_8270,N_7763,N_7089);
or U8271 (N_8271,N_7869,N_7166);
or U8272 (N_8272,N_7850,N_7387);
nor U8273 (N_8273,N_7359,N_7233);
nor U8274 (N_8274,N_7235,N_7256);
and U8275 (N_8275,N_7915,N_7710);
nand U8276 (N_8276,N_7680,N_7067);
or U8277 (N_8277,N_7493,N_7031);
nor U8278 (N_8278,N_7595,N_7243);
and U8279 (N_8279,N_7229,N_7524);
nand U8280 (N_8280,N_7409,N_7344);
xnor U8281 (N_8281,N_7893,N_7609);
or U8282 (N_8282,N_7186,N_7968);
nor U8283 (N_8283,N_7808,N_7294);
and U8284 (N_8284,N_7028,N_7440);
nand U8285 (N_8285,N_7142,N_7815);
nor U8286 (N_8286,N_7573,N_7882);
nand U8287 (N_8287,N_7020,N_7283);
or U8288 (N_8288,N_7900,N_7541);
or U8289 (N_8289,N_7696,N_7104);
nor U8290 (N_8290,N_7558,N_7985);
nand U8291 (N_8291,N_7534,N_7471);
and U8292 (N_8292,N_7549,N_7781);
or U8293 (N_8293,N_7097,N_7986);
or U8294 (N_8294,N_7975,N_7402);
nor U8295 (N_8295,N_7279,N_7112);
nor U8296 (N_8296,N_7803,N_7892);
nand U8297 (N_8297,N_7320,N_7870);
and U8298 (N_8298,N_7063,N_7162);
nand U8299 (N_8299,N_7553,N_7075);
nor U8300 (N_8300,N_7772,N_7307);
or U8301 (N_8301,N_7219,N_7671);
or U8302 (N_8302,N_7161,N_7934);
nor U8303 (N_8303,N_7393,N_7519);
nand U8304 (N_8304,N_7750,N_7916);
nor U8305 (N_8305,N_7397,N_7860);
nor U8306 (N_8306,N_7606,N_7909);
nor U8307 (N_8307,N_7515,N_7322);
nand U8308 (N_8308,N_7957,N_7199);
nand U8309 (N_8309,N_7336,N_7319);
and U8310 (N_8310,N_7974,N_7218);
nor U8311 (N_8311,N_7572,N_7056);
or U8312 (N_8312,N_7466,N_7890);
nor U8313 (N_8313,N_7192,N_7202);
or U8314 (N_8314,N_7687,N_7864);
nor U8315 (N_8315,N_7818,N_7447);
nand U8316 (N_8316,N_7117,N_7312);
nor U8317 (N_8317,N_7535,N_7564);
nand U8318 (N_8318,N_7997,N_7521);
or U8319 (N_8319,N_7905,N_7489);
nand U8320 (N_8320,N_7565,N_7600);
nor U8321 (N_8321,N_7326,N_7315);
nand U8322 (N_8322,N_7630,N_7377);
nand U8323 (N_8323,N_7779,N_7255);
nand U8324 (N_8324,N_7220,N_7462);
nor U8325 (N_8325,N_7331,N_7183);
nand U8326 (N_8326,N_7268,N_7788);
and U8327 (N_8327,N_7197,N_7300);
and U8328 (N_8328,N_7100,N_7129);
nand U8329 (N_8329,N_7807,N_7329);
nor U8330 (N_8330,N_7958,N_7125);
and U8331 (N_8331,N_7431,N_7308);
or U8332 (N_8332,N_7619,N_7930);
nor U8333 (N_8333,N_7405,N_7748);
or U8334 (N_8334,N_7646,N_7237);
or U8335 (N_8335,N_7698,N_7768);
nand U8336 (N_8336,N_7757,N_7038);
and U8337 (N_8337,N_7699,N_7396);
or U8338 (N_8338,N_7266,N_7732);
nand U8339 (N_8339,N_7875,N_7648);
and U8340 (N_8340,N_7634,N_7525);
nor U8341 (N_8341,N_7507,N_7747);
and U8342 (N_8342,N_7718,N_7799);
nor U8343 (N_8343,N_7275,N_7041);
nand U8344 (N_8344,N_7679,N_7678);
nand U8345 (N_8345,N_7996,N_7478);
nand U8346 (N_8346,N_7454,N_7551);
nor U8347 (N_8347,N_7389,N_7855);
and U8348 (N_8348,N_7071,N_7338);
or U8349 (N_8349,N_7381,N_7871);
nand U8350 (N_8350,N_7724,N_7756);
or U8351 (N_8351,N_7584,N_7429);
or U8352 (N_8352,N_7490,N_7586);
nor U8353 (N_8353,N_7849,N_7079);
nor U8354 (N_8354,N_7264,N_7951);
nor U8355 (N_8355,N_7777,N_7221);
or U8356 (N_8356,N_7657,N_7147);
nor U8357 (N_8357,N_7794,N_7444);
nand U8358 (N_8358,N_7879,N_7141);
or U8359 (N_8359,N_7057,N_7058);
or U8360 (N_8360,N_7222,N_7497);
and U8361 (N_8361,N_7983,N_7090);
nor U8362 (N_8362,N_7421,N_7548);
xnor U8363 (N_8363,N_7651,N_7017);
nor U8364 (N_8364,N_7704,N_7371);
nor U8365 (N_8365,N_7839,N_7617);
nor U8366 (N_8366,N_7119,N_7177);
and U8367 (N_8367,N_7969,N_7506);
and U8368 (N_8368,N_7593,N_7224);
nand U8369 (N_8369,N_7837,N_7165);
or U8370 (N_8370,N_7685,N_7254);
and U8371 (N_8371,N_7380,N_7103);
and U8372 (N_8372,N_7596,N_7232);
nor U8373 (N_8373,N_7923,N_7365);
nand U8374 (N_8374,N_7760,N_7345);
nand U8375 (N_8375,N_7881,N_7567);
nand U8376 (N_8376,N_7804,N_7475);
nor U8377 (N_8377,N_7245,N_7591);
nand U8378 (N_8378,N_7349,N_7856);
nor U8379 (N_8379,N_7293,N_7120);
nand U8380 (N_8380,N_7422,N_7759);
and U8381 (N_8381,N_7469,N_7416);
nand U8382 (N_8382,N_7692,N_7672);
or U8383 (N_8383,N_7321,N_7786);
or U8384 (N_8384,N_7468,N_7948);
nor U8385 (N_8385,N_7884,N_7350);
nor U8386 (N_8386,N_7003,N_7898);
nor U8387 (N_8387,N_7694,N_7877);
or U8388 (N_8388,N_7611,N_7705);
or U8389 (N_8389,N_7925,N_7011);
nand U8390 (N_8390,N_7514,N_7417);
nand U8391 (N_8391,N_7379,N_7569);
nor U8392 (N_8392,N_7883,N_7543);
nand U8393 (N_8393,N_7372,N_7834);
and U8394 (N_8394,N_7399,N_7614);
nand U8395 (N_8395,N_7343,N_7676);
nand U8396 (N_8396,N_7209,N_7023);
nand U8397 (N_8397,N_7066,N_7291);
nand U8398 (N_8398,N_7095,N_7034);
nor U8399 (N_8399,N_7713,N_7305);
nor U8400 (N_8400,N_7076,N_7227);
and U8401 (N_8401,N_7960,N_7862);
xor U8402 (N_8402,N_7771,N_7460);
and U8403 (N_8403,N_7620,N_7026);
or U8404 (N_8404,N_7107,N_7559);
nor U8405 (N_8405,N_7946,N_7725);
and U8406 (N_8406,N_7675,N_7863);
nand U8407 (N_8407,N_7520,N_7010);
nand U8408 (N_8408,N_7907,N_7526);
and U8409 (N_8409,N_7636,N_7635);
or U8410 (N_8410,N_7550,N_7825);
and U8411 (N_8411,N_7159,N_7036);
or U8412 (N_8412,N_7295,N_7200);
nand U8413 (N_8413,N_7590,N_7624);
nand U8414 (N_8414,N_7709,N_7386);
nor U8415 (N_8415,N_7570,N_7688);
nor U8416 (N_8416,N_7050,N_7587);
nand U8417 (N_8417,N_7173,N_7842);
or U8418 (N_8418,N_7027,N_7265);
nand U8419 (N_8419,N_7194,N_7138);
nor U8420 (N_8420,N_7000,N_7740);
nand U8421 (N_8421,N_7848,N_7990);
or U8422 (N_8422,N_7445,N_7729);
or U8423 (N_8423,N_7106,N_7623);
nand U8424 (N_8424,N_7306,N_7552);
nand U8425 (N_8425,N_7783,N_7780);
and U8426 (N_8426,N_7318,N_7742);
nor U8427 (N_8427,N_7124,N_7504);
nand U8428 (N_8428,N_7311,N_7217);
and U8429 (N_8429,N_7568,N_7858);
nor U8430 (N_8430,N_7660,N_7018);
and U8431 (N_8431,N_7410,N_7172);
nor U8432 (N_8432,N_7741,N_7438);
nor U8433 (N_8433,N_7622,N_7662);
or U8434 (N_8434,N_7208,N_7375);
nor U8435 (N_8435,N_7752,N_7262);
nor U8436 (N_8436,N_7484,N_7814);
nand U8437 (N_8437,N_7894,N_7663);
or U8438 (N_8438,N_7269,N_7121);
or U8439 (N_8439,N_7632,N_7108);
or U8440 (N_8440,N_7435,N_7873);
or U8441 (N_8441,N_7992,N_7897);
nor U8442 (N_8442,N_7810,N_7667);
nor U8443 (N_8443,N_7053,N_7528);
nand U8444 (N_8444,N_7328,N_7977);
nor U8445 (N_8445,N_7082,N_7556);
nand U8446 (N_8446,N_7966,N_7204);
and U8447 (N_8447,N_7032,N_7730);
and U8448 (N_8448,N_7285,N_7695);
nor U8449 (N_8449,N_7203,N_7248);
nor U8450 (N_8450,N_7802,N_7423);
nand U8451 (N_8451,N_7169,N_7188);
or U8452 (N_8452,N_7140,N_7030);
nor U8453 (N_8453,N_7263,N_7271);
nor U8454 (N_8454,N_7463,N_7251);
or U8455 (N_8455,N_7157,N_7978);
and U8456 (N_8456,N_7886,N_7868);
nand U8457 (N_8457,N_7214,N_7253);
nand U8458 (N_8458,N_7503,N_7216);
xnor U8459 (N_8459,N_7168,N_7546);
nand U8460 (N_8460,N_7984,N_7655);
nor U8461 (N_8461,N_7215,N_7292);
nand U8462 (N_8462,N_7540,N_7436);
nand U8463 (N_8463,N_7247,N_7577);
nor U8464 (N_8464,N_7170,N_7014);
nor U8465 (N_8465,N_7637,N_7653);
and U8466 (N_8466,N_7160,N_7073);
nand U8467 (N_8467,N_7432,N_7339);
nor U8468 (N_8468,N_7080,N_7367);
nor U8469 (N_8469,N_7607,N_7212);
nand U8470 (N_8470,N_7801,N_7959);
or U8471 (N_8471,N_7927,N_7952);
and U8472 (N_8472,N_7743,N_7029);
nand U8473 (N_8473,N_7330,N_7238);
nand U8474 (N_8474,N_7764,N_7949);
nand U8475 (N_8475,N_7746,N_7085);
nand U8476 (N_8476,N_7048,N_7420);
nor U8477 (N_8477,N_7859,N_7993);
nor U8478 (N_8478,N_7758,N_7439);
or U8479 (N_8479,N_7482,N_7499);
nand U8480 (N_8480,N_7042,N_7920);
nor U8481 (N_8481,N_7583,N_7289);
and U8482 (N_8482,N_7703,N_7681);
nand U8483 (N_8483,N_7821,N_7115);
nand U8484 (N_8484,N_7754,N_7231);
nor U8485 (N_8485,N_7988,N_7158);
or U8486 (N_8486,N_7323,N_7327);
nor U8487 (N_8487,N_7190,N_7070);
and U8488 (N_8488,N_7486,N_7136);
or U8489 (N_8489,N_7823,N_7861);
nand U8490 (N_8490,N_7954,N_7749);
nor U8491 (N_8491,N_7270,N_7701);
or U8492 (N_8492,N_7302,N_7656);
and U8493 (N_8493,N_7589,N_7874);
nor U8494 (N_8494,N_7155,N_7415);
or U8495 (N_8495,N_7427,N_7488);
and U8496 (N_8496,N_7257,N_7274);
nand U8497 (N_8497,N_7734,N_7728);
nand U8498 (N_8498,N_7686,N_7132);
nand U8499 (N_8499,N_7335,N_7476);
nand U8500 (N_8500,N_7189,N_7383);
and U8501 (N_8501,N_7213,N_7065);
and U8502 (N_8502,N_7069,N_7391);
nand U8503 (N_8503,N_7980,N_7779);
nand U8504 (N_8504,N_7735,N_7725);
nor U8505 (N_8505,N_7608,N_7454);
nor U8506 (N_8506,N_7084,N_7746);
and U8507 (N_8507,N_7784,N_7919);
or U8508 (N_8508,N_7418,N_7667);
and U8509 (N_8509,N_7269,N_7005);
or U8510 (N_8510,N_7898,N_7477);
and U8511 (N_8511,N_7735,N_7302);
nor U8512 (N_8512,N_7283,N_7796);
and U8513 (N_8513,N_7795,N_7128);
and U8514 (N_8514,N_7845,N_7668);
or U8515 (N_8515,N_7223,N_7682);
nand U8516 (N_8516,N_7203,N_7413);
or U8517 (N_8517,N_7007,N_7495);
or U8518 (N_8518,N_7046,N_7300);
or U8519 (N_8519,N_7160,N_7291);
nor U8520 (N_8520,N_7610,N_7489);
and U8521 (N_8521,N_7680,N_7521);
and U8522 (N_8522,N_7267,N_7721);
nand U8523 (N_8523,N_7912,N_7202);
or U8524 (N_8524,N_7070,N_7376);
and U8525 (N_8525,N_7761,N_7268);
or U8526 (N_8526,N_7031,N_7468);
nand U8527 (N_8527,N_7027,N_7005);
nor U8528 (N_8528,N_7910,N_7224);
nor U8529 (N_8529,N_7265,N_7256);
nor U8530 (N_8530,N_7433,N_7361);
nand U8531 (N_8531,N_7086,N_7509);
or U8532 (N_8532,N_7736,N_7855);
and U8533 (N_8533,N_7185,N_7172);
and U8534 (N_8534,N_7581,N_7127);
nor U8535 (N_8535,N_7438,N_7686);
nor U8536 (N_8536,N_7878,N_7458);
and U8537 (N_8537,N_7115,N_7783);
nand U8538 (N_8538,N_7977,N_7217);
or U8539 (N_8539,N_7134,N_7671);
or U8540 (N_8540,N_7856,N_7987);
nand U8541 (N_8541,N_7817,N_7965);
nand U8542 (N_8542,N_7491,N_7060);
or U8543 (N_8543,N_7095,N_7409);
nor U8544 (N_8544,N_7301,N_7819);
nand U8545 (N_8545,N_7977,N_7848);
nor U8546 (N_8546,N_7397,N_7264);
and U8547 (N_8547,N_7929,N_7021);
and U8548 (N_8548,N_7432,N_7713);
or U8549 (N_8549,N_7833,N_7730);
or U8550 (N_8550,N_7464,N_7506);
or U8551 (N_8551,N_7611,N_7571);
nand U8552 (N_8552,N_7917,N_7447);
and U8553 (N_8553,N_7966,N_7369);
and U8554 (N_8554,N_7251,N_7538);
and U8555 (N_8555,N_7431,N_7905);
or U8556 (N_8556,N_7200,N_7117);
nand U8557 (N_8557,N_7741,N_7181);
nand U8558 (N_8558,N_7140,N_7246);
nand U8559 (N_8559,N_7007,N_7737);
nand U8560 (N_8560,N_7159,N_7083);
or U8561 (N_8561,N_7265,N_7765);
nand U8562 (N_8562,N_7636,N_7417);
nor U8563 (N_8563,N_7048,N_7343);
nor U8564 (N_8564,N_7770,N_7607);
nand U8565 (N_8565,N_7553,N_7854);
nand U8566 (N_8566,N_7697,N_7617);
and U8567 (N_8567,N_7394,N_7097);
and U8568 (N_8568,N_7883,N_7303);
nand U8569 (N_8569,N_7356,N_7640);
and U8570 (N_8570,N_7034,N_7903);
nand U8571 (N_8571,N_7369,N_7109);
or U8572 (N_8572,N_7772,N_7896);
and U8573 (N_8573,N_7491,N_7677);
nor U8574 (N_8574,N_7160,N_7989);
and U8575 (N_8575,N_7087,N_7519);
nor U8576 (N_8576,N_7319,N_7034);
and U8577 (N_8577,N_7700,N_7363);
or U8578 (N_8578,N_7444,N_7517);
and U8579 (N_8579,N_7750,N_7207);
nor U8580 (N_8580,N_7512,N_7935);
nor U8581 (N_8581,N_7537,N_7357);
or U8582 (N_8582,N_7959,N_7330);
nor U8583 (N_8583,N_7606,N_7062);
and U8584 (N_8584,N_7619,N_7899);
nand U8585 (N_8585,N_7649,N_7572);
nor U8586 (N_8586,N_7739,N_7778);
nand U8587 (N_8587,N_7222,N_7545);
nor U8588 (N_8588,N_7668,N_7797);
and U8589 (N_8589,N_7009,N_7177);
nand U8590 (N_8590,N_7369,N_7560);
nor U8591 (N_8591,N_7021,N_7850);
nor U8592 (N_8592,N_7105,N_7929);
or U8593 (N_8593,N_7493,N_7508);
and U8594 (N_8594,N_7987,N_7483);
or U8595 (N_8595,N_7099,N_7139);
and U8596 (N_8596,N_7398,N_7123);
nand U8597 (N_8597,N_7361,N_7876);
or U8598 (N_8598,N_7779,N_7752);
and U8599 (N_8599,N_7233,N_7781);
and U8600 (N_8600,N_7505,N_7432);
or U8601 (N_8601,N_7739,N_7950);
nor U8602 (N_8602,N_7008,N_7201);
or U8603 (N_8603,N_7137,N_7284);
or U8604 (N_8604,N_7940,N_7146);
nor U8605 (N_8605,N_7285,N_7591);
nor U8606 (N_8606,N_7961,N_7295);
nand U8607 (N_8607,N_7326,N_7618);
nand U8608 (N_8608,N_7478,N_7079);
nand U8609 (N_8609,N_7316,N_7905);
nand U8610 (N_8610,N_7927,N_7538);
nand U8611 (N_8611,N_7104,N_7834);
nor U8612 (N_8612,N_7792,N_7207);
and U8613 (N_8613,N_7060,N_7410);
nand U8614 (N_8614,N_7516,N_7171);
nand U8615 (N_8615,N_7708,N_7235);
or U8616 (N_8616,N_7486,N_7996);
and U8617 (N_8617,N_7264,N_7037);
nor U8618 (N_8618,N_7750,N_7075);
or U8619 (N_8619,N_7622,N_7282);
nor U8620 (N_8620,N_7350,N_7006);
or U8621 (N_8621,N_7574,N_7367);
nand U8622 (N_8622,N_7197,N_7995);
nor U8623 (N_8623,N_7636,N_7254);
or U8624 (N_8624,N_7359,N_7530);
or U8625 (N_8625,N_7613,N_7551);
nand U8626 (N_8626,N_7569,N_7859);
nor U8627 (N_8627,N_7351,N_7610);
nor U8628 (N_8628,N_7568,N_7346);
or U8629 (N_8629,N_7322,N_7427);
or U8630 (N_8630,N_7002,N_7030);
nor U8631 (N_8631,N_7046,N_7853);
nor U8632 (N_8632,N_7290,N_7247);
nor U8633 (N_8633,N_7599,N_7034);
nor U8634 (N_8634,N_7957,N_7515);
nand U8635 (N_8635,N_7291,N_7030);
and U8636 (N_8636,N_7496,N_7240);
nand U8637 (N_8637,N_7064,N_7146);
or U8638 (N_8638,N_7715,N_7134);
nor U8639 (N_8639,N_7520,N_7640);
and U8640 (N_8640,N_7110,N_7350);
nand U8641 (N_8641,N_7436,N_7182);
or U8642 (N_8642,N_7336,N_7549);
nand U8643 (N_8643,N_7007,N_7958);
nand U8644 (N_8644,N_7117,N_7308);
and U8645 (N_8645,N_7737,N_7616);
nand U8646 (N_8646,N_7358,N_7965);
and U8647 (N_8647,N_7386,N_7001);
nor U8648 (N_8648,N_7954,N_7373);
nor U8649 (N_8649,N_7037,N_7659);
nor U8650 (N_8650,N_7913,N_7677);
nor U8651 (N_8651,N_7001,N_7194);
and U8652 (N_8652,N_7447,N_7267);
and U8653 (N_8653,N_7065,N_7814);
and U8654 (N_8654,N_7761,N_7285);
and U8655 (N_8655,N_7601,N_7530);
and U8656 (N_8656,N_7849,N_7865);
nor U8657 (N_8657,N_7624,N_7792);
and U8658 (N_8658,N_7764,N_7441);
xnor U8659 (N_8659,N_7064,N_7973);
and U8660 (N_8660,N_7115,N_7306);
nor U8661 (N_8661,N_7616,N_7231);
nor U8662 (N_8662,N_7474,N_7377);
nor U8663 (N_8663,N_7554,N_7529);
nand U8664 (N_8664,N_7172,N_7571);
or U8665 (N_8665,N_7973,N_7934);
nor U8666 (N_8666,N_7879,N_7289);
nor U8667 (N_8667,N_7140,N_7910);
nand U8668 (N_8668,N_7519,N_7624);
nor U8669 (N_8669,N_7603,N_7029);
or U8670 (N_8670,N_7032,N_7551);
or U8671 (N_8671,N_7198,N_7855);
nor U8672 (N_8672,N_7182,N_7679);
nand U8673 (N_8673,N_7436,N_7902);
nor U8674 (N_8674,N_7198,N_7066);
nor U8675 (N_8675,N_7350,N_7888);
and U8676 (N_8676,N_7109,N_7879);
and U8677 (N_8677,N_7049,N_7966);
or U8678 (N_8678,N_7913,N_7997);
or U8679 (N_8679,N_7507,N_7022);
or U8680 (N_8680,N_7545,N_7880);
and U8681 (N_8681,N_7920,N_7010);
and U8682 (N_8682,N_7321,N_7050);
or U8683 (N_8683,N_7244,N_7272);
or U8684 (N_8684,N_7521,N_7612);
or U8685 (N_8685,N_7976,N_7098);
nor U8686 (N_8686,N_7193,N_7024);
nor U8687 (N_8687,N_7661,N_7603);
nand U8688 (N_8688,N_7834,N_7207);
nor U8689 (N_8689,N_7058,N_7926);
and U8690 (N_8690,N_7058,N_7251);
and U8691 (N_8691,N_7165,N_7907);
nand U8692 (N_8692,N_7660,N_7354);
and U8693 (N_8693,N_7477,N_7436);
and U8694 (N_8694,N_7759,N_7107);
nand U8695 (N_8695,N_7495,N_7820);
or U8696 (N_8696,N_7910,N_7526);
nor U8697 (N_8697,N_7486,N_7118);
nand U8698 (N_8698,N_7150,N_7850);
nand U8699 (N_8699,N_7897,N_7671);
and U8700 (N_8700,N_7521,N_7883);
or U8701 (N_8701,N_7375,N_7471);
or U8702 (N_8702,N_7638,N_7084);
nand U8703 (N_8703,N_7335,N_7329);
or U8704 (N_8704,N_7850,N_7993);
nand U8705 (N_8705,N_7574,N_7927);
or U8706 (N_8706,N_7396,N_7312);
nor U8707 (N_8707,N_7150,N_7353);
and U8708 (N_8708,N_7487,N_7043);
or U8709 (N_8709,N_7080,N_7172);
nand U8710 (N_8710,N_7312,N_7235);
or U8711 (N_8711,N_7408,N_7615);
nor U8712 (N_8712,N_7074,N_7896);
nor U8713 (N_8713,N_7827,N_7078);
nand U8714 (N_8714,N_7725,N_7631);
nand U8715 (N_8715,N_7061,N_7669);
or U8716 (N_8716,N_7279,N_7803);
nor U8717 (N_8717,N_7249,N_7992);
nor U8718 (N_8718,N_7605,N_7556);
nor U8719 (N_8719,N_7132,N_7663);
nor U8720 (N_8720,N_7033,N_7834);
nor U8721 (N_8721,N_7973,N_7484);
xor U8722 (N_8722,N_7995,N_7793);
nand U8723 (N_8723,N_7135,N_7376);
or U8724 (N_8724,N_7483,N_7544);
or U8725 (N_8725,N_7020,N_7419);
and U8726 (N_8726,N_7299,N_7476);
nand U8727 (N_8727,N_7974,N_7020);
and U8728 (N_8728,N_7479,N_7667);
and U8729 (N_8729,N_7451,N_7556);
and U8730 (N_8730,N_7253,N_7673);
nor U8731 (N_8731,N_7443,N_7879);
or U8732 (N_8732,N_7501,N_7682);
or U8733 (N_8733,N_7067,N_7213);
and U8734 (N_8734,N_7484,N_7937);
or U8735 (N_8735,N_7140,N_7827);
nand U8736 (N_8736,N_7096,N_7274);
nor U8737 (N_8737,N_7084,N_7481);
or U8738 (N_8738,N_7661,N_7997);
nand U8739 (N_8739,N_7388,N_7498);
nand U8740 (N_8740,N_7493,N_7364);
or U8741 (N_8741,N_7810,N_7983);
nor U8742 (N_8742,N_7760,N_7099);
and U8743 (N_8743,N_7596,N_7848);
or U8744 (N_8744,N_7396,N_7921);
xnor U8745 (N_8745,N_7374,N_7028);
nor U8746 (N_8746,N_7142,N_7762);
and U8747 (N_8747,N_7425,N_7324);
nand U8748 (N_8748,N_7969,N_7523);
or U8749 (N_8749,N_7172,N_7654);
nand U8750 (N_8750,N_7336,N_7621);
nor U8751 (N_8751,N_7398,N_7221);
or U8752 (N_8752,N_7159,N_7470);
nor U8753 (N_8753,N_7715,N_7886);
nor U8754 (N_8754,N_7253,N_7007);
or U8755 (N_8755,N_7991,N_7623);
and U8756 (N_8756,N_7149,N_7667);
nor U8757 (N_8757,N_7064,N_7126);
nor U8758 (N_8758,N_7239,N_7767);
and U8759 (N_8759,N_7988,N_7756);
nand U8760 (N_8760,N_7554,N_7881);
nand U8761 (N_8761,N_7800,N_7590);
nand U8762 (N_8762,N_7556,N_7334);
or U8763 (N_8763,N_7885,N_7428);
or U8764 (N_8764,N_7263,N_7831);
or U8765 (N_8765,N_7476,N_7310);
nand U8766 (N_8766,N_7747,N_7479);
and U8767 (N_8767,N_7156,N_7612);
nor U8768 (N_8768,N_7019,N_7797);
nand U8769 (N_8769,N_7900,N_7661);
or U8770 (N_8770,N_7821,N_7728);
nand U8771 (N_8771,N_7159,N_7860);
or U8772 (N_8772,N_7440,N_7387);
or U8773 (N_8773,N_7736,N_7546);
or U8774 (N_8774,N_7139,N_7825);
nand U8775 (N_8775,N_7620,N_7224);
nor U8776 (N_8776,N_7720,N_7128);
or U8777 (N_8777,N_7797,N_7454);
and U8778 (N_8778,N_7991,N_7771);
nor U8779 (N_8779,N_7289,N_7642);
nor U8780 (N_8780,N_7409,N_7529);
nor U8781 (N_8781,N_7135,N_7474);
nand U8782 (N_8782,N_7599,N_7598);
nand U8783 (N_8783,N_7669,N_7966);
nand U8784 (N_8784,N_7040,N_7584);
nor U8785 (N_8785,N_7029,N_7755);
nor U8786 (N_8786,N_7214,N_7616);
nor U8787 (N_8787,N_7928,N_7094);
nand U8788 (N_8788,N_7873,N_7314);
or U8789 (N_8789,N_7701,N_7064);
and U8790 (N_8790,N_7873,N_7740);
or U8791 (N_8791,N_7123,N_7734);
nand U8792 (N_8792,N_7368,N_7073);
nand U8793 (N_8793,N_7320,N_7024);
nand U8794 (N_8794,N_7114,N_7368);
nor U8795 (N_8795,N_7498,N_7957);
or U8796 (N_8796,N_7128,N_7013);
nand U8797 (N_8797,N_7915,N_7401);
and U8798 (N_8798,N_7111,N_7523);
and U8799 (N_8799,N_7466,N_7900);
nor U8800 (N_8800,N_7133,N_7812);
nor U8801 (N_8801,N_7166,N_7006);
and U8802 (N_8802,N_7971,N_7111);
or U8803 (N_8803,N_7828,N_7351);
xor U8804 (N_8804,N_7853,N_7339);
and U8805 (N_8805,N_7905,N_7566);
nor U8806 (N_8806,N_7112,N_7368);
and U8807 (N_8807,N_7266,N_7275);
xor U8808 (N_8808,N_7421,N_7467);
nand U8809 (N_8809,N_7877,N_7315);
nor U8810 (N_8810,N_7740,N_7496);
nand U8811 (N_8811,N_7744,N_7038);
nand U8812 (N_8812,N_7892,N_7586);
nor U8813 (N_8813,N_7974,N_7078);
and U8814 (N_8814,N_7560,N_7113);
nor U8815 (N_8815,N_7588,N_7694);
or U8816 (N_8816,N_7781,N_7150);
nand U8817 (N_8817,N_7039,N_7596);
nor U8818 (N_8818,N_7540,N_7041);
and U8819 (N_8819,N_7564,N_7566);
and U8820 (N_8820,N_7432,N_7911);
and U8821 (N_8821,N_7101,N_7675);
xor U8822 (N_8822,N_7813,N_7783);
and U8823 (N_8823,N_7218,N_7068);
or U8824 (N_8824,N_7306,N_7546);
or U8825 (N_8825,N_7377,N_7311);
or U8826 (N_8826,N_7718,N_7360);
and U8827 (N_8827,N_7137,N_7296);
or U8828 (N_8828,N_7909,N_7723);
nor U8829 (N_8829,N_7487,N_7681);
or U8830 (N_8830,N_7759,N_7187);
nor U8831 (N_8831,N_7631,N_7715);
nor U8832 (N_8832,N_7471,N_7257);
nand U8833 (N_8833,N_7991,N_7083);
or U8834 (N_8834,N_7731,N_7769);
or U8835 (N_8835,N_7180,N_7123);
nor U8836 (N_8836,N_7446,N_7662);
or U8837 (N_8837,N_7158,N_7324);
nor U8838 (N_8838,N_7684,N_7987);
or U8839 (N_8839,N_7023,N_7989);
or U8840 (N_8840,N_7440,N_7109);
or U8841 (N_8841,N_7662,N_7046);
or U8842 (N_8842,N_7992,N_7709);
nor U8843 (N_8843,N_7444,N_7516);
and U8844 (N_8844,N_7671,N_7604);
nand U8845 (N_8845,N_7447,N_7561);
or U8846 (N_8846,N_7726,N_7036);
nand U8847 (N_8847,N_7514,N_7227);
or U8848 (N_8848,N_7343,N_7582);
and U8849 (N_8849,N_7499,N_7571);
and U8850 (N_8850,N_7092,N_7992);
or U8851 (N_8851,N_7827,N_7753);
nor U8852 (N_8852,N_7014,N_7842);
and U8853 (N_8853,N_7924,N_7364);
nand U8854 (N_8854,N_7853,N_7151);
and U8855 (N_8855,N_7197,N_7273);
or U8856 (N_8856,N_7250,N_7941);
and U8857 (N_8857,N_7827,N_7939);
nand U8858 (N_8858,N_7925,N_7647);
nand U8859 (N_8859,N_7109,N_7173);
nor U8860 (N_8860,N_7230,N_7644);
or U8861 (N_8861,N_7531,N_7309);
or U8862 (N_8862,N_7161,N_7127);
nor U8863 (N_8863,N_7659,N_7450);
and U8864 (N_8864,N_7583,N_7723);
nand U8865 (N_8865,N_7599,N_7294);
or U8866 (N_8866,N_7987,N_7164);
nand U8867 (N_8867,N_7322,N_7679);
or U8868 (N_8868,N_7279,N_7400);
nor U8869 (N_8869,N_7635,N_7303);
and U8870 (N_8870,N_7709,N_7296);
nor U8871 (N_8871,N_7921,N_7927);
nor U8872 (N_8872,N_7941,N_7985);
nor U8873 (N_8873,N_7166,N_7097);
or U8874 (N_8874,N_7975,N_7822);
nand U8875 (N_8875,N_7827,N_7648);
nor U8876 (N_8876,N_7498,N_7005);
nor U8877 (N_8877,N_7082,N_7367);
nor U8878 (N_8878,N_7579,N_7856);
or U8879 (N_8879,N_7079,N_7908);
and U8880 (N_8880,N_7478,N_7138);
or U8881 (N_8881,N_7464,N_7395);
and U8882 (N_8882,N_7406,N_7478);
nor U8883 (N_8883,N_7941,N_7305);
and U8884 (N_8884,N_7149,N_7695);
or U8885 (N_8885,N_7786,N_7463);
or U8886 (N_8886,N_7402,N_7798);
nand U8887 (N_8887,N_7731,N_7428);
or U8888 (N_8888,N_7484,N_7445);
nand U8889 (N_8889,N_7796,N_7657);
and U8890 (N_8890,N_7920,N_7304);
and U8891 (N_8891,N_7498,N_7583);
and U8892 (N_8892,N_7253,N_7504);
nand U8893 (N_8893,N_7016,N_7226);
or U8894 (N_8894,N_7687,N_7351);
and U8895 (N_8895,N_7217,N_7340);
and U8896 (N_8896,N_7399,N_7899);
nand U8897 (N_8897,N_7597,N_7897);
xor U8898 (N_8898,N_7039,N_7191);
nor U8899 (N_8899,N_7319,N_7110);
nor U8900 (N_8900,N_7406,N_7515);
and U8901 (N_8901,N_7492,N_7782);
nand U8902 (N_8902,N_7112,N_7683);
nor U8903 (N_8903,N_7750,N_7296);
or U8904 (N_8904,N_7731,N_7624);
and U8905 (N_8905,N_7863,N_7833);
and U8906 (N_8906,N_7464,N_7912);
nor U8907 (N_8907,N_7797,N_7640);
nand U8908 (N_8908,N_7291,N_7767);
nand U8909 (N_8909,N_7735,N_7856);
nand U8910 (N_8910,N_7621,N_7839);
and U8911 (N_8911,N_7914,N_7024);
nand U8912 (N_8912,N_7761,N_7916);
and U8913 (N_8913,N_7840,N_7918);
nor U8914 (N_8914,N_7839,N_7981);
or U8915 (N_8915,N_7957,N_7421);
or U8916 (N_8916,N_7306,N_7689);
nor U8917 (N_8917,N_7049,N_7121);
or U8918 (N_8918,N_7580,N_7401);
nor U8919 (N_8919,N_7129,N_7429);
or U8920 (N_8920,N_7819,N_7381);
nor U8921 (N_8921,N_7757,N_7747);
nor U8922 (N_8922,N_7033,N_7415);
and U8923 (N_8923,N_7797,N_7998);
and U8924 (N_8924,N_7308,N_7957);
nor U8925 (N_8925,N_7862,N_7968);
and U8926 (N_8926,N_7302,N_7881);
nor U8927 (N_8927,N_7318,N_7564);
nand U8928 (N_8928,N_7160,N_7377);
and U8929 (N_8929,N_7358,N_7160);
nor U8930 (N_8930,N_7933,N_7773);
nand U8931 (N_8931,N_7407,N_7316);
or U8932 (N_8932,N_7430,N_7686);
or U8933 (N_8933,N_7203,N_7772);
or U8934 (N_8934,N_7629,N_7847);
nand U8935 (N_8935,N_7542,N_7655);
nand U8936 (N_8936,N_7204,N_7802);
or U8937 (N_8937,N_7342,N_7072);
nor U8938 (N_8938,N_7665,N_7979);
and U8939 (N_8939,N_7602,N_7730);
nand U8940 (N_8940,N_7460,N_7845);
or U8941 (N_8941,N_7736,N_7808);
or U8942 (N_8942,N_7206,N_7016);
or U8943 (N_8943,N_7121,N_7161);
nand U8944 (N_8944,N_7660,N_7058);
and U8945 (N_8945,N_7739,N_7281);
or U8946 (N_8946,N_7155,N_7068);
nor U8947 (N_8947,N_7760,N_7590);
nand U8948 (N_8948,N_7793,N_7401);
nor U8949 (N_8949,N_7813,N_7317);
and U8950 (N_8950,N_7989,N_7574);
nor U8951 (N_8951,N_7399,N_7774);
and U8952 (N_8952,N_7990,N_7001);
nor U8953 (N_8953,N_7493,N_7410);
nand U8954 (N_8954,N_7171,N_7025);
or U8955 (N_8955,N_7821,N_7490);
nor U8956 (N_8956,N_7420,N_7248);
and U8957 (N_8957,N_7777,N_7602);
and U8958 (N_8958,N_7600,N_7997);
or U8959 (N_8959,N_7605,N_7625);
nor U8960 (N_8960,N_7826,N_7416);
or U8961 (N_8961,N_7129,N_7098);
nand U8962 (N_8962,N_7700,N_7900);
or U8963 (N_8963,N_7479,N_7165);
or U8964 (N_8964,N_7242,N_7574);
or U8965 (N_8965,N_7069,N_7689);
nor U8966 (N_8966,N_7166,N_7308);
or U8967 (N_8967,N_7754,N_7293);
or U8968 (N_8968,N_7034,N_7923);
nand U8969 (N_8969,N_7218,N_7989);
nor U8970 (N_8970,N_7298,N_7876);
or U8971 (N_8971,N_7226,N_7315);
nor U8972 (N_8972,N_7933,N_7931);
nor U8973 (N_8973,N_7311,N_7652);
nor U8974 (N_8974,N_7512,N_7985);
or U8975 (N_8975,N_7272,N_7805);
nand U8976 (N_8976,N_7659,N_7124);
and U8977 (N_8977,N_7651,N_7641);
or U8978 (N_8978,N_7046,N_7880);
nor U8979 (N_8979,N_7752,N_7075);
and U8980 (N_8980,N_7581,N_7871);
and U8981 (N_8981,N_7099,N_7673);
nor U8982 (N_8982,N_7671,N_7468);
nor U8983 (N_8983,N_7253,N_7938);
nor U8984 (N_8984,N_7246,N_7477);
nand U8985 (N_8985,N_7888,N_7602);
nor U8986 (N_8986,N_7132,N_7582);
nor U8987 (N_8987,N_7309,N_7405);
nand U8988 (N_8988,N_7561,N_7954);
or U8989 (N_8989,N_7141,N_7860);
nand U8990 (N_8990,N_7412,N_7935);
nor U8991 (N_8991,N_7700,N_7345);
nand U8992 (N_8992,N_7107,N_7467);
and U8993 (N_8993,N_7451,N_7656);
or U8994 (N_8994,N_7624,N_7035);
or U8995 (N_8995,N_7638,N_7786);
and U8996 (N_8996,N_7831,N_7403);
nand U8997 (N_8997,N_7144,N_7560);
or U8998 (N_8998,N_7122,N_7182);
or U8999 (N_8999,N_7457,N_7715);
xnor U9000 (N_9000,N_8605,N_8460);
nor U9001 (N_9001,N_8894,N_8471);
nand U9002 (N_9002,N_8767,N_8038);
nor U9003 (N_9003,N_8808,N_8656);
and U9004 (N_9004,N_8765,N_8698);
nand U9005 (N_9005,N_8457,N_8020);
nor U9006 (N_9006,N_8695,N_8996);
and U9007 (N_9007,N_8660,N_8077);
and U9008 (N_9008,N_8167,N_8347);
nand U9009 (N_9009,N_8396,N_8845);
and U9010 (N_9010,N_8659,N_8434);
nor U9011 (N_9011,N_8991,N_8854);
nor U9012 (N_9012,N_8777,N_8910);
nor U9013 (N_9013,N_8941,N_8979);
nor U9014 (N_9014,N_8814,N_8934);
nand U9015 (N_9015,N_8776,N_8165);
and U9016 (N_9016,N_8542,N_8795);
nor U9017 (N_9017,N_8568,N_8056);
and U9018 (N_9018,N_8464,N_8268);
or U9019 (N_9019,N_8549,N_8309);
nand U9020 (N_9020,N_8633,N_8490);
and U9021 (N_9021,N_8320,N_8972);
nand U9022 (N_9022,N_8405,N_8872);
nor U9023 (N_9023,N_8703,N_8376);
nor U9024 (N_9024,N_8031,N_8499);
nor U9025 (N_9025,N_8519,N_8939);
nand U9026 (N_9026,N_8640,N_8015);
or U9027 (N_9027,N_8737,N_8770);
nand U9028 (N_9028,N_8212,N_8055);
and U9029 (N_9029,N_8476,N_8412);
nand U9030 (N_9030,N_8775,N_8738);
and U9031 (N_9031,N_8148,N_8159);
nor U9032 (N_9032,N_8319,N_8743);
and U9033 (N_9033,N_8564,N_8867);
xor U9034 (N_9034,N_8379,N_8544);
and U9035 (N_9035,N_8646,N_8806);
nand U9036 (N_9036,N_8558,N_8086);
or U9037 (N_9037,N_8535,N_8235);
nor U9038 (N_9038,N_8006,N_8959);
nand U9039 (N_9039,N_8198,N_8132);
or U9040 (N_9040,N_8181,N_8900);
or U9041 (N_9041,N_8245,N_8270);
or U9042 (N_9042,N_8740,N_8197);
nor U9043 (N_9043,N_8053,N_8114);
nor U9044 (N_9044,N_8855,N_8919);
nor U9045 (N_9045,N_8373,N_8302);
or U9046 (N_9046,N_8019,N_8751);
and U9047 (N_9047,N_8926,N_8849);
nand U9048 (N_9048,N_8012,N_8248);
nor U9049 (N_9049,N_8966,N_8526);
and U9050 (N_9050,N_8068,N_8456);
and U9051 (N_9051,N_8290,N_8547);
nand U9052 (N_9052,N_8760,N_8316);
nand U9053 (N_9053,N_8579,N_8378);
or U9054 (N_9054,N_8258,N_8073);
or U9055 (N_9055,N_8291,N_8754);
nor U9056 (N_9056,N_8466,N_8237);
and U9057 (N_9057,N_8361,N_8022);
and U9058 (N_9058,N_8955,N_8193);
or U9059 (N_9059,N_8483,N_8602);
or U9060 (N_9060,N_8037,N_8699);
nor U9061 (N_9061,N_8064,N_8920);
or U9062 (N_9062,N_8469,N_8723);
xor U9063 (N_9063,N_8997,N_8447);
xor U9064 (N_9064,N_8732,N_8834);
nor U9065 (N_9065,N_8311,N_8087);
or U9066 (N_9066,N_8324,N_8016);
or U9067 (N_9067,N_8488,N_8416);
or U9068 (N_9068,N_8848,N_8817);
nand U9069 (N_9069,N_8911,N_8799);
or U9070 (N_9070,N_8244,N_8837);
nor U9071 (N_9071,N_8642,N_8724);
and U9072 (N_9072,N_8620,N_8190);
and U9073 (N_9073,N_8062,N_8216);
nor U9074 (N_9074,N_8601,N_8250);
nor U9075 (N_9075,N_8442,N_8709);
and U9076 (N_9076,N_8338,N_8096);
nor U9077 (N_9077,N_8074,N_8040);
nor U9078 (N_9078,N_8662,N_8501);
nor U9079 (N_9079,N_8293,N_8890);
nand U9080 (N_9080,N_8921,N_8836);
nand U9081 (N_9081,N_8851,N_8233);
and U9082 (N_9082,N_8679,N_8344);
nor U9083 (N_9083,N_8119,N_8339);
nor U9084 (N_9084,N_8079,N_8722);
or U9085 (N_9085,N_8830,N_8175);
nor U9086 (N_9086,N_8155,N_8051);
and U9087 (N_9087,N_8671,N_8002);
and U9088 (N_9088,N_8788,N_8430);
or U9089 (N_9089,N_8294,N_8478);
nand U9090 (N_9090,N_8906,N_8154);
and U9091 (N_9091,N_8680,N_8880);
nor U9092 (N_9092,N_8385,N_8368);
and U9093 (N_9093,N_8990,N_8752);
and U9094 (N_9094,N_8323,N_8701);
and U9095 (N_9095,N_8661,N_8308);
or U9096 (N_9096,N_8357,N_8214);
or U9097 (N_9097,N_8869,N_8759);
nor U9098 (N_9098,N_8611,N_8513);
or U9099 (N_9099,N_8637,N_8971);
nor U9100 (N_9100,N_8596,N_8439);
nor U9101 (N_9101,N_8774,N_8994);
and U9102 (N_9102,N_8942,N_8280);
nor U9103 (N_9103,N_8683,N_8711);
nor U9104 (N_9104,N_8871,N_8390);
nand U9105 (N_9105,N_8438,N_8185);
nand U9106 (N_9106,N_8599,N_8807);
nand U9107 (N_9107,N_8341,N_8678);
nor U9108 (N_9108,N_8206,N_8420);
and U9109 (N_9109,N_8322,N_8133);
nor U9110 (N_9110,N_8715,N_8780);
nor U9111 (N_9111,N_8809,N_8204);
nand U9112 (N_9112,N_8103,N_8383);
and U9113 (N_9113,N_8419,N_8962);
nand U9114 (N_9114,N_8164,N_8853);
xor U9115 (N_9115,N_8335,N_8034);
nor U9116 (N_9116,N_8652,N_8271);
nor U9117 (N_9117,N_8575,N_8340);
nor U9118 (N_9118,N_8741,N_8153);
nor U9119 (N_9119,N_8627,N_8350);
nand U9120 (N_9120,N_8023,N_8584);
nand U9121 (N_9121,N_8411,N_8744);
nor U9122 (N_9122,N_8102,N_8884);
and U9123 (N_9123,N_8098,N_8036);
nand U9124 (N_9124,N_8733,N_8076);
nor U9125 (N_9125,N_8054,N_8839);
nand U9126 (N_9126,N_8730,N_8172);
and U9127 (N_9127,N_8630,N_8757);
and U9128 (N_9128,N_8707,N_8009);
nand U9129 (N_9129,N_8859,N_8567);
nor U9130 (N_9130,N_8060,N_8590);
or U9131 (N_9131,N_8746,N_8232);
nand U9132 (N_9132,N_8915,N_8951);
nor U9133 (N_9133,N_8146,N_8262);
nand U9134 (N_9134,N_8509,N_8496);
and U9135 (N_9135,N_8812,N_8937);
nand U9136 (N_9136,N_8604,N_8672);
nor U9137 (N_9137,N_8913,N_8677);
nand U9138 (N_9138,N_8532,N_8755);
nor U9139 (N_9139,N_8446,N_8901);
or U9140 (N_9140,N_8981,N_8092);
nand U9141 (N_9141,N_8902,N_8935);
nor U9142 (N_9142,N_8515,N_8107);
nor U9143 (N_9143,N_8097,N_8441);
and U9144 (N_9144,N_8173,N_8522);
nand U9145 (N_9145,N_8862,N_8682);
or U9146 (N_9146,N_8521,N_8230);
and U9147 (N_9147,N_8348,N_8993);
nor U9148 (N_9148,N_8083,N_8003);
and U9149 (N_9149,N_8943,N_8893);
nor U9150 (N_9150,N_8622,N_8534);
nor U9151 (N_9151,N_8169,N_8388);
and U9152 (N_9152,N_8613,N_8988);
nand U9153 (N_9153,N_8857,N_8525);
nand U9154 (N_9154,N_8545,N_8649);
nor U9155 (N_9155,N_8641,N_8600);
nor U9156 (N_9156,N_8463,N_8465);
nand U9157 (N_9157,N_8093,N_8475);
or U9158 (N_9158,N_8426,N_8796);
nor U9159 (N_9159,N_8461,N_8885);
nand U9160 (N_9160,N_8219,N_8980);
nor U9161 (N_9161,N_8790,N_8462);
or U9162 (N_9162,N_8355,N_8178);
nand U9163 (N_9163,N_8592,N_8061);
nor U9164 (N_9164,N_8793,N_8213);
and U9165 (N_9165,N_8399,N_8126);
or U9166 (N_9166,N_8139,N_8726);
nand U9167 (N_9167,N_8041,N_8143);
nor U9168 (N_9168,N_8422,N_8868);
nand U9169 (N_9169,N_8612,N_8909);
and U9170 (N_9170,N_8514,N_8756);
and U9171 (N_9171,N_8505,N_8653);
and U9172 (N_9172,N_8846,N_8259);
nor U9173 (N_9173,N_8905,N_8066);
and U9174 (N_9174,N_8960,N_8331);
nor U9175 (N_9175,N_8318,N_8288);
nand U9176 (N_9176,N_8301,N_8931);
nand U9177 (N_9177,N_8595,N_8289);
or U9178 (N_9178,N_8574,N_8778);
or U9179 (N_9179,N_8229,N_8130);
nand U9180 (N_9180,N_8372,N_8576);
nor U9181 (N_9181,N_8184,N_8435);
or U9182 (N_9182,N_8110,N_8918);
and U9183 (N_9183,N_8543,N_8149);
and U9184 (N_9184,N_8401,N_8030);
nand U9185 (N_9185,N_8182,N_8117);
nand U9186 (N_9186,N_8263,N_8847);
nor U9187 (N_9187,N_8587,N_8384);
nor U9188 (N_9188,N_8518,N_8382);
nand U9189 (N_9189,N_8142,N_8690);
or U9190 (N_9190,N_8581,N_8560);
nand U9191 (N_9191,N_8156,N_8897);
or U9192 (N_9192,N_8976,N_8398);
nand U9193 (N_9193,N_8414,N_8606);
nand U9194 (N_9194,N_8970,N_8503);
nand U9195 (N_9195,N_8516,N_8432);
and U9196 (N_9196,N_8748,N_8450);
or U9197 (N_9197,N_8222,N_8561);
nand U9198 (N_9198,N_8000,N_8436);
nor U9199 (N_9199,N_8598,N_8639);
nor U9200 (N_9200,N_8850,N_8704);
nand U9201 (N_9201,N_8231,N_8785);
and U9202 (N_9202,N_8786,N_8789);
nand U9203 (N_9203,N_8654,N_8234);
and U9204 (N_9204,N_8424,N_8122);
and U9205 (N_9205,N_8591,N_8202);
nor U9206 (N_9206,N_8467,N_8138);
nor U9207 (N_9207,N_8710,N_8914);
nand U9208 (N_9208,N_8615,N_8895);
nand U9209 (N_9209,N_8278,N_8174);
and U9210 (N_9210,N_8004,N_8444);
nor U9211 (N_9211,N_8618,N_8391);
nor U9212 (N_9212,N_8029,N_8645);
nand U9213 (N_9213,N_8882,N_8665);
nand U9214 (N_9214,N_8792,N_8180);
or U9215 (N_9215,N_8694,N_8314);
and U9216 (N_9216,N_8084,N_8731);
nor U9217 (N_9217,N_8876,N_8326);
nand U9218 (N_9218,N_8129,N_8067);
or U9219 (N_9219,N_8527,N_8987);
or U9220 (N_9220,N_8151,N_8137);
nor U9221 (N_9221,N_8860,N_8533);
xnor U9222 (N_9222,N_8844,N_8824);
nand U9223 (N_9223,N_8228,N_8394);
or U9224 (N_9224,N_8688,N_8157);
nand U9225 (N_9225,N_8619,N_8063);
nand U9226 (N_9226,N_8801,N_8307);
or U9227 (N_9227,N_8523,N_8431);
nand U9228 (N_9228,N_8573,N_8927);
nor U9229 (N_9229,N_8256,N_8337);
or U9230 (N_9230,N_8395,N_8546);
or U9231 (N_9231,N_8091,N_8603);
nor U9232 (N_9232,N_8205,N_8236);
or U9233 (N_9233,N_8100,N_8451);
nand U9234 (N_9234,N_8626,N_8531);
nand U9235 (N_9235,N_8183,N_8470);
xor U9236 (N_9236,N_8945,N_8891);
and U9237 (N_9237,N_8624,N_8948);
or U9238 (N_9238,N_8220,N_8021);
and U9239 (N_9239,N_8866,N_8032);
and U9240 (N_9240,N_8249,N_8026);
and U9241 (N_9241,N_8362,N_8582);
nand U9242 (N_9242,N_8179,N_8402);
nor U9243 (N_9243,N_8804,N_8769);
and U9244 (N_9244,N_8717,N_8186);
nor U9245 (N_9245,N_8768,N_8306);
or U9246 (N_9246,N_8359,N_8145);
or U9247 (N_9247,N_8540,N_8089);
or U9248 (N_9248,N_8049,N_8713);
nor U9249 (N_9249,N_8681,N_8930);
or U9250 (N_9250,N_8856,N_8989);
and U9251 (N_9251,N_8152,N_8124);
or U9252 (N_9252,N_8017,N_8517);
and U9253 (N_9253,N_8504,N_8265);
or U9254 (N_9254,N_8371,N_8276);
nor U9255 (N_9255,N_8115,N_8965);
nand U9256 (N_9256,N_8865,N_8936);
and U9257 (N_9257,N_8254,N_8933);
nand U9258 (N_9258,N_8208,N_8749);
and U9259 (N_9259,N_8636,N_8668);
and U9260 (N_9260,N_8059,N_8566);
or U9261 (N_9261,N_8123,N_8223);
and U9262 (N_9262,N_8246,N_8329);
or U9263 (N_9263,N_8712,N_8508);
nor U9264 (N_9264,N_8226,N_8369);
nor U9265 (N_9265,N_8800,N_8492);
or U9266 (N_9266,N_8118,N_8045);
or U9267 (N_9267,N_8417,N_8629);
nor U9268 (N_9268,N_8367,N_8632);
nand U9269 (N_9269,N_8728,N_8039);
or U9270 (N_9270,N_8950,N_8113);
and U9271 (N_9271,N_8947,N_8954);
and U9272 (N_9272,N_8802,N_8833);
nand U9273 (N_9273,N_8095,N_8365);
nand U9274 (N_9274,N_8283,N_8445);
and U9275 (N_9275,N_8716,N_8433);
or U9276 (N_9276,N_8821,N_8116);
nor U9277 (N_9277,N_8614,N_8840);
xor U9278 (N_9278,N_8239,N_8969);
or U9279 (N_9279,N_8010,N_8718);
nand U9280 (N_9280,N_8489,N_8277);
and U9281 (N_9281,N_8071,N_8287);
nand U9282 (N_9282,N_8696,N_8764);
or U9283 (N_9283,N_8571,N_8562);
nor U9284 (N_9284,N_8984,N_8404);
and U9285 (N_9285,N_8697,N_8664);
or U9286 (N_9286,N_8192,N_8413);
or U9287 (N_9287,N_8007,N_8082);
nor U9288 (N_9288,N_8843,N_8336);
nand U9289 (N_9289,N_8274,N_8468);
nor U9290 (N_9290,N_8787,N_8537);
nor U9291 (N_9291,N_8272,N_8810);
and U9292 (N_9292,N_8131,N_8354);
nor U9293 (N_9293,N_8013,N_8472);
and U9294 (N_9294,N_8104,N_8892);
and U9295 (N_9295,N_8052,N_8766);
and U9296 (N_9296,N_8304,N_8218);
and U9297 (N_9297,N_8838,N_8588);
and U9298 (N_9298,N_8721,N_8739);
nor U9299 (N_9299,N_8403,N_8841);
nand U9300 (N_9300,N_8940,N_8473);
nand U9301 (N_9301,N_8455,N_8597);
and U9302 (N_9302,N_8529,N_8783);
or U9303 (N_9303,N_8480,N_8791);
or U9304 (N_9304,N_8929,N_8474);
nand U9305 (N_9305,N_8485,N_8794);
and U9306 (N_9306,N_8158,N_8747);
nor U9307 (N_9307,N_8200,N_8727);
or U9308 (N_9308,N_8896,N_8166);
or U9309 (N_9309,N_8745,N_8899);
nor U9310 (N_9310,N_8201,N_8638);
nand U9311 (N_9311,N_8643,N_8247);
and U9312 (N_9312,N_8211,N_8978);
and U9313 (N_9313,N_8631,N_8539);
nor U9314 (N_9314,N_8387,N_8108);
or U9315 (N_9315,N_8685,N_8608);
and U9316 (N_9316,N_8317,N_8085);
or U9317 (N_9317,N_8963,N_8903);
nand U9318 (N_9318,N_8275,N_8454);
nand U9319 (N_9319,N_8360,N_8938);
nor U9320 (N_9320,N_8874,N_8332);
nor U9321 (N_9321,N_8285,N_8177);
or U9322 (N_9322,N_8328,N_8556);
xor U9323 (N_9323,N_8070,N_8825);
nand U9324 (N_9324,N_8621,N_8415);
or U9325 (N_9325,N_8586,N_8033);
or U9326 (N_9326,N_8589,N_8363);
and U9327 (N_9327,N_8481,N_8330);
nand U9328 (N_9328,N_8418,N_8816);
nand U9329 (N_9329,N_8958,N_8452);
and U9330 (N_9330,N_8565,N_8554);
nor U9331 (N_9331,N_8553,N_8080);
nor U9332 (N_9332,N_8313,N_8267);
and U9333 (N_9333,N_8502,N_8907);
nand U9334 (N_9334,N_8956,N_8510);
or U9335 (N_9335,N_8644,N_8861);
and U9336 (N_9336,N_8163,N_8299);
nand U9337 (N_9337,N_8583,N_8224);
nor U9338 (N_9338,N_8141,N_8714);
or U9339 (N_9339,N_8106,N_8983);
and U9340 (N_9340,N_8407,N_8101);
xor U9341 (N_9341,N_8982,N_8803);
nand U9342 (N_9342,N_8282,N_8736);
and U9343 (N_9343,N_8691,N_8975);
nand U9344 (N_9344,N_8058,N_8784);
nand U9345 (N_9345,N_8829,N_8551);
nand U9346 (N_9346,N_8449,N_8011);
or U9347 (N_9347,N_8917,N_8044);
or U9348 (N_9348,N_8345,N_8273);
nand U9349 (N_9349,N_8392,N_8797);
nor U9350 (N_9350,N_8353,N_8873);
nand U9351 (N_9351,N_8078,N_8497);
and U9352 (N_9352,N_8925,N_8400);
nand U9353 (N_9353,N_8827,N_8512);
xor U9354 (N_9354,N_8842,N_8238);
and U9355 (N_9355,N_8686,N_8027);
nand U9356 (N_9356,N_8831,N_8374);
and U9357 (N_9357,N_8014,N_8187);
nand U9358 (N_9358,N_8150,N_8541);
or U9359 (N_9359,N_8781,N_8176);
nor U9360 (N_9360,N_8072,N_8203);
and U9361 (N_9361,N_8050,N_8487);
nand U9362 (N_9362,N_8875,N_8753);
nor U9363 (N_9363,N_8295,N_8952);
and U9364 (N_9364,N_8048,N_8559);
nand U9365 (N_9365,N_8887,N_8823);
and U9366 (N_9366,N_8210,N_8321);
nand U9367 (N_9367,N_8425,N_8194);
and U9368 (N_9368,N_8818,N_8820);
and U9369 (N_9369,N_8358,N_8477);
nand U9370 (N_9370,N_8973,N_8813);
nand U9371 (N_9371,N_8008,N_8486);
and U9372 (N_9372,N_8908,N_8577);
and U9373 (N_9373,N_8189,N_8269);
nor U9374 (N_9374,N_8491,N_8162);
and U9375 (N_9375,N_8042,N_8377);
nor U9376 (N_9376,N_8112,N_8782);
or U9377 (N_9377,N_8779,N_8427);
or U9378 (N_9378,N_8440,N_8932);
or U9379 (N_9379,N_8196,N_8720);
or U9380 (N_9380,N_8999,N_8437);
nand U9381 (N_9381,N_8687,N_8370);
nand U9382 (N_9382,N_8610,N_8260);
nand U9383 (N_9383,N_8957,N_8209);
nand U9384 (N_9384,N_8443,N_8284);
or U9385 (N_9385,N_8507,N_8099);
and U9386 (N_9386,N_8240,N_8028);
or U9387 (N_9387,N_8702,N_8120);
or U9388 (N_9388,N_8160,N_8352);
or U9389 (N_9389,N_8161,N_8410);
or U9390 (N_9390,N_8217,N_8429);
nand U9391 (N_9391,N_8018,N_8735);
or U9392 (N_9392,N_8327,N_8296);
and U9393 (N_9393,N_8625,N_8111);
nand U9394 (N_9394,N_8255,N_8889);
and U9395 (N_9395,N_8105,N_8992);
or U9396 (N_9396,N_8944,N_8563);
and U9397 (N_9397,N_8428,N_8761);
nand U9398 (N_9398,N_8758,N_8835);
or U9399 (N_9399,N_8995,N_8725);
and U9400 (N_9400,N_8397,N_8538);
and U9401 (N_9401,N_8572,N_8708);
nand U9402 (N_9402,N_8195,N_8593);
and U9403 (N_9403,N_8257,N_8922);
nor U9404 (N_9404,N_8852,N_8252);
nand U9405 (N_9405,N_8985,N_8520);
nor U9406 (N_9406,N_8121,N_8227);
nand U9407 (N_9407,N_8705,N_8675);
or U9408 (N_9408,N_8670,N_8706);
or U9409 (N_9409,N_8580,N_8171);
or U9410 (N_9410,N_8136,N_8953);
and U9411 (N_9411,N_8500,N_8170);
nand U9412 (N_9412,N_8719,N_8094);
nor U9413 (N_9413,N_8135,N_8334);
nand U9414 (N_9414,N_8511,N_8081);
nand U9415 (N_9415,N_8798,N_8811);
nand U9416 (N_9416,N_8570,N_8912);
nor U9417 (N_9417,N_8729,N_8090);
or U9418 (N_9418,N_8552,N_8634);
and U9419 (N_9419,N_8569,N_8967);
and U9420 (N_9420,N_8264,N_8870);
or U9421 (N_9421,N_8221,N_8968);
nor U9422 (N_9422,N_8286,N_8663);
xnor U9423 (N_9423,N_8127,N_8998);
and U9424 (N_9424,N_8692,N_8312);
or U9425 (N_9425,N_8075,N_8506);
and U9426 (N_9426,N_8303,N_8253);
xnor U9427 (N_9427,N_8858,N_8923);
nor U9428 (N_9428,N_8555,N_8878);
or U9429 (N_9429,N_8024,N_8356);
nor U9430 (N_9430,N_8964,N_8946);
and U9431 (N_9431,N_8346,N_8916);
nor U9432 (N_9432,N_8928,N_8088);
nand U9433 (N_9433,N_8207,N_8977);
nor U9434 (N_9434,N_8125,N_8279);
or U9435 (N_9435,N_8381,N_8025);
nor U9436 (N_9436,N_8199,N_8635);
nand U9437 (N_9437,N_8351,N_8828);
or U9438 (N_9438,N_8616,N_8557);
and U9439 (N_9439,N_8674,N_8188);
xor U9440 (N_9440,N_8864,N_8409);
nor U9441 (N_9441,N_8607,N_8883);
nor U9442 (N_9442,N_8243,N_8225);
xor U9443 (N_9443,N_8375,N_8667);
and U9444 (N_9444,N_8453,N_8536);
nand U9445 (N_9445,N_8310,N_8408);
or U9446 (N_9446,N_8684,N_8648);
and U9447 (N_9447,N_8421,N_8251);
or U9448 (N_9448,N_8147,N_8005);
and U9449 (N_9449,N_8924,N_8881);
or U9450 (N_9450,N_8578,N_8046);
nand U9451 (N_9451,N_8266,N_8647);
and U9452 (N_9452,N_8047,N_8380);
nand U9453 (N_9453,N_8655,N_8949);
nor U9454 (N_9454,N_8689,N_8528);
nand U9455 (N_9455,N_8657,N_8617);
or U9456 (N_9456,N_8134,N_8550);
or U9457 (N_9457,N_8734,N_8886);
and U9458 (N_9458,N_8482,N_8001);
and U9459 (N_9459,N_8065,N_8877);
nor U9460 (N_9460,N_8298,N_8548);
nor U9461 (N_9461,N_8609,N_8458);
nand U9462 (N_9462,N_8494,N_8495);
or U9463 (N_9463,N_8423,N_8666);
or U9464 (N_9464,N_8292,N_8676);
nand U9465 (N_9465,N_8585,N_8822);
nor U9466 (N_9466,N_8628,N_8524);
nor U9467 (N_9467,N_8364,N_8043);
and U9468 (N_9468,N_8389,N_8366);
or U9469 (N_9469,N_8815,N_8281);
nor U9470 (N_9470,N_8493,N_8623);
and U9471 (N_9471,N_8832,N_8888);
or U9472 (N_9472,N_8826,N_8772);
nor U9473 (N_9473,N_8315,N_8140);
and U9474 (N_9474,N_8773,N_8898);
and U9475 (N_9475,N_8771,N_8325);
and U9476 (N_9476,N_8386,N_8673);
xor U9477 (N_9477,N_8594,N_8700);
and U9478 (N_9478,N_8242,N_8762);
or U9479 (N_9479,N_8069,N_8763);
nor U9480 (N_9480,N_8658,N_8669);
or U9481 (N_9481,N_8057,N_8168);
or U9482 (N_9482,N_8448,N_8342);
nor U9483 (N_9483,N_8819,N_8459);
or U9484 (N_9484,N_8693,N_8333);
or U9485 (N_9485,N_8144,N_8128);
or U9486 (N_9486,N_8479,N_8484);
or U9487 (N_9487,N_8191,N_8863);
and U9488 (N_9488,N_8742,N_8498);
nand U9489 (N_9489,N_8530,N_8297);
and U9490 (N_9490,N_8261,N_8974);
nor U9491 (N_9491,N_8651,N_8343);
and U9492 (N_9492,N_8879,N_8035);
and U9493 (N_9493,N_8961,N_8393);
nand U9494 (N_9494,N_8750,N_8406);
or U9495 (N_9495,N_8109,N_8904);
nor U9496 (N_9496,N_8805,N_8650);
nor U9497 (N_9497,N_8215,N_8300);
and U9498 (N_9498,N_8349,N_8986);
nor U9499 (N_9499,N_8241,N_8305);
and U9500 (N_9500,N_8454,N_8918);
nor U9501 (N_9501,N_8686,N_8307);
nand U9502 (N_9502,N_8845,N_8050);
and U9503 (N_9503,N_8725,N_8488);
or U9504 (N_9504,N_8513,N_8708);
or U9505 (N_9505,N_8109,N_8985);
nor U9506 (N_9506,N_8792,N_8407);
or U9507 (N_9507,N_8508,N_8872);
or U9508 (N_9508,N_8605,N_8458);
xnor U9509 (N_9509,N_8826,N_8167);
nand U9510 (N_9510,N_8386,N_8124);
nor U9511 (N_9511,N_8689,N_8548);
nor U9512 (N_9512,N_8583,N_8853);
or U9513 (N_9513,N_8904,N_8493);
nand U9514 (N_9514,N_8202,N_8346);
and U9515 (N_9515,N_8209,N_8897);
or U9516 (N_9516,N_8603,N_8721);
and U9517 (N_9517,N_8767,N_8598);
and U9518 (N_9518,N_8490,N_8946);
and U9519 (N_9519,N_8308,N_8970);
nand U9520 (N_9520,N_8752,N_8682);
or U9521 (N_9521,N_8149,N_8380);
nand U9522 (N_9522,N_8160,N_8344);
or U9523 (N_9523,N_8037,N_8603);
or U9524 (N_9524,N_8158,N_8005);
and U9525 (N_9525,N_8585,N_8494);
nand U9526 (N_9526,N_8767,N_8757);
and U9527 (N_9527,N_8979,N_8333);
nand U9528 (N_9528,N_8604,N_8958);
and U9529 (N_9529,N_8970,N_8155);
or U9530 (N_9530,N_8729,N_8582);
nor U9531 (N_9531,N_8085,N_8525);
nand U9532 (N_9532,N_8557,N_8539);
nand U9533 (N_9533,N_8522,N_8843);
nor U9534 (N_9534,N_8999,N_8474);
nor U9535 (N_9535,N_8842,N_8756);
nand U9536 (N_9536,N_8649,N_8945);
nand U9537 (N_9537,N_8599,N_8154);
nor U9538 (N_9538,N_8507,N_8706);
and U9539 (N_9539,N_8959,N_8891);
nor U9540 (N_9540,N_8810,N_8745);
or U9541 (N_9541,N_8770,N_8174);
and U9542 (N_9542,N_8115,N_8279);
nor U9543 (N_9543,N_8477,N_8093);
nand U9544 (N_9544,N_8247,N_8561);
or U9545 (N_9545,N_8634,N_8729);
and U9546 (N_9546,N_8949,N_8271);
nand U9547 (N_9547,N_8489,N_8215);
and U9548 (N_9548,N_8427,N_8302);
and U9549 (N_9549,N_8810,N_8379);
or U9550 (N_9550,N_8785,N_8133);
nor U9551 (N_9551,N_8263,N_8186);
nor U9552 (N_9552,N_8777,N_8438);
and U9553 (N_9553,N_8229,N_8579);
nand U9554 (N_9554,N_8989,N_8060);
and U9555 (N_9555,N_8108,N_8907);
nand U9556 (N_9556,N_8608,N_8092);
or U9557 (N_9557,N_8886,N_8055);
or U9558 (N_9558,N_8742,N_8531);
or U9559 (N_9559,N_8626,N_8548);
and U9560 (N_9560,N_8922,N_8501);
and U9561 (N_9561,N_8826,N_8868);
nand U9562 (N_9562,N_8933,N_8693);
or U9563 (N_9563,N_8721,N_8966);
and U9564 (N_9564,N_8618,N_8177);
nand U9565 (N_9565,N_8483,N_8063);
nand U9566 (N_9566,N_8536,N_8114);
and U9567 (N_9567,N_8620,N_8015);
or U9568 (N_9568,N_8698,N_8509);
nor U9569 (N_9569,N_8509,N_8618);
nand U9570 (N_9570,N_8913,N_8650);
and U9571 (N_9571,N_8039,N_8315);
nor U9572 (N_9572,N_8444,N_8943);
nor U9573 (N_9573,N_8166,N_8855);
or U9574 (N_9574,N_8783,N_8137);
or U9575 (N_9575,N_8531,N_8581);
nand U9576 (N_9576,N_8823,N_8351);
nand U9577 (N_9577,N_8013,N_8314);
or U9578 (N_9578,N_8443,N_8696);
nor U9579 (N_9579,N_8569,N_8961);
and U9580 (N_9580,N_8002,N_8362);
and U9581 (N_9581,N_8841,N_8308);
nand U9582 (N_9582,N_8438,N_8839);
or U9583 (N_9583,N_8877,N_8898);
and U9584 (N_9584,N_8369,N_8419);
and U9585 (N_9585,N_8631,N_8402);
and U9586 (N_9586,N_8376,N_8199);
or U9587 (N_9587,N_8626,N_8520);
nand U9588 (N_9588,N_8685,N_8615);
nand U9589 (N_9589,N_8665,N_8473);
or U9590 (N_9590,N_8593,N_8495);
and U9591 (N_9591,N_8119,N_8962);
xnor U9592 (N_9592,N_8822,N_8692);
nand U9593 (N_9593,N_8079,N_8007);
nor U9594 (N_9594,N_8438,N_8019);
and U9595 (N_9595,N_8331,N_8667);
and U9596 (N_9596,N_8914,N_8338);
nor U9597 (N_9597,N_8431,N_8420);
nand U9598 (N_9598,N_8324,N_8864);
nand U9599 (N_9599,N_8452,N_8734);
nand U9600 (N_9600,N_8801,N_8300);
nor U9601 (N_9601,N_8415,N_8159);
nand U9602 (N_9602,N_8660,N_8192);
and U9603 (N_9603,N_8904,N_8780);
nand U9604 (N_9604,N_8959,N_8947);
or U9605 (N_9605,N_8217,N_8948);
nor U9606 (N_9606,N_8241,N_8301);
and U9607 (N_9607,N_8437,N_8733);
or U9608 (N_9608,N_8742,N_8798);
and U9609 (N_9609,N_8530,N_8750);
or U9610 (N_9610,N_8100,N_8255);
and U9611 (N_9611,N_8595,N_8484);
nor U9612 (N_9612,N_8106,N_8689);
nor U9613 (N_9613,N_8565,N_8129);
nor U9614 (N_9614,N_8052,N_8175);
nor U9615 (N_9615,N_8186,N_8052);
xor U9616 (N_9616,N_8390,N_8855);
and U9617 (N_9617,N_8073,N_8455);
nor U9618 (N_9618,N_8084,N_8275);
nand U9619 (N_9619,N_8607,N_8875);
and U9620 (N_9620,N_8065,N_8146);
and U9621 (N_9621,N_8898,N_8311);
nand U9622 (N_9622,N_8349,N_8151);
or U9623 (N_9623,N_8955,N_8628);
nand U9624 (N_9624,N_8353,N_8401);
nor U9625 (N_9625,N_8306,N_8889);
or U9626 (N_9626,N_8230,N_8545);
nand U9627 (N_9627,N_8635,N_8558);
and U9628 (N_9628,N_8526,N_8019);
nand U9629 (N_9629,N_8586,N_8453);
and U9630 (N_9630,N_8816,N_8790);
nand U9631 (N_9631,N_8224,N_8809);
and U9632 (N_9632,N_8183,N_8374);
nand U9633 (N_9633,N_8403,N_8285);
nand U9634 (N_9634,N_8775,N_8855);
or U9635 (N_9635,N_8654,N_8073);
nor U9636 (N_9636,N_8761,N_8342);
and U9637 (N_9637,N_8259,N_8385);
nand U9638 (N_9638,N_8864,N_8135);
nand U9639 (N_9639,N_8799,N_8910);
and U9640 (N_9640,N_8706,N_8258);
and U9641 (N_9641,N_8551,N_8882);
xor U9642 (N_9642,N_8974,N_8262);
or U9643 (N_9643,N_8712,N_8569);
and U9644 (N_9644,N_8298,N_8338);
nor U9645 (N_9645,N_8100,N_8165);
nand U9646 (N_9646,N_8076,N_8050);
and U9647 (N_9647,N_8374,N_8434);
or U9648 (N_9648,N_8214,N_8688);
or U9649 (N_9649,N_8663,N_8327);
and U9650 (N_9650,N_8135,N_8622);
nand U9651 (N_9651,N_8688,N_8147);
or U9652 (N_9652,N_8495,N_8638);
nand U9653 (N_9653,N_8702,N_8728);
nor U9654 (N_9654,N_8214,N_8739);
nor U9655 (N_9655,N_8299,N_8585);
or U9656 (N_9656,N_8336,N_8917);
nor U9657 (N_9657,N_8184,N_8474);
or U9658 (N_9658,N_8478,N_8731);
and U9659 (N_9659,N_8953,N_8985);
or U9660 (N_9660,N_8155,N_8863);
or U9661 (N_9661,N_8455,N_8364);
nand U9662 (N_9662,N_8154,N_8343);
and U9663 (N_9663,N_8759,N_8108);
and U9664 (N_9664,N_8829,N_8848);
or U9665 (N_9665,N_8724,N_8284);
xnor U9666 (N_9666,N_8952,N_8298);
and U9667 (N_9667,N_8800,N_8459);
and U9668 (N_9668,N_8052,N_8402);
nand U9669 (N_9669,N_8353,N_8114);
and U9670 (N_9670,N_8047,N_8111);
nor U9671 (N_9671,N_8761,N_8079);
or U9672 (N_9672,N_8619,N_8027);
nor U9673 (N_9673,N_8779,N_8662);
nand U9674 (N_9674,N_8506,N_8503);
nor U9675 (N_9675,N_8197,N_8478);
nor U9676 (N_9676,N_8252,N_8308);
or U9677 (N_9677,N_8859,N_8346);
and U9678 (N_9678,N_8241,N_8322);
and U9679 (N_9679,N_8505,N_8070);
nor U9680 (N_9680,N_8901,N_8152);
nor U9681 (N_9681,N_8983,N_8977);
or U9682 (N_9682,N_8834,N_8902);
or U9683 (N_9683,N_8958,N_8348);
or U9684 (N_9684,N_8262,N_8327);
nor U9685 (N_9685,N_8427,N_8193);
or U9686 (N_9686,N_8403,N_8169);
or U9687 (N_9687,N_8522,N_8213);
nand U9688 (N_9688,N_8321,N_8522);
or U9689 (N_9689,N_8910,N_8295);
or U9690 (N_9690,N_8017,N_8765);
or U9691 (N_9691,N_8260,N_8361);
or U9692 (N_9692,N_8168,N_8802);
nor U9693 (N_9693,N_8059,N_8357);
xor U9694 (N_9694,N_8441,N_8635);
and U9695 (N_9695,N_8109,N_8295);
nand U9696 (N_9696,N_8897,N_8216);
and U9697 (N_9697,N_8738,N_8595);
nor U9698 (N_9698,N_8328,N_8070);
and U9699 (N_9699,N_8236,N_8492);
or U9700 (N_9700,N_8574,N_8146);
nor U9701 (N_9701,N_8050,N_8538);
nand U9702 (N_9702,N_8576,N_8220);
or U9703 (N_9703,N_8056,N_8667);
and U9704 (N_9704,N_8465,N_8455);
or U9705 (N_9705,N_8236,N_8346);
and U9706 (N_9706,N_8871,N_8616);
or U9707 (N_9707,N_8175,N_8155);
or U9708 (N_9708,N_8697,N_8728);
or U9709 (N_9709,N_8534,N_8655);
or U9710 (N_9710,N_8096,N_8190);
xor U9711 (N_9711,N_8957,N_8351);
nor U9712 (N_9712,N_8867,N_8534);
or U9713 (N_9713,N_8381,N_8129);
nor U9714 (N_9714,N_8597,N_8169);
or U9715 (N_9715,N_8850,N_8686);
nor U9716 (N_9716,N_8018,N_8411);
and U9717 (N_9717,N_8038,N_8546);
and U9718 (N_9718,N_8386,N_8467);
nand U9719 (N_9719,N_8934,N_8565);
or U9720 (N_9720,N_8614,N_8338);
nand U9721 (N_9721,N_8072,N_8638);
and U9722 (N_9722,N_8368,N_8278);
or U9723 (N_9723,N_8989,N_8449);
and U9724 (N_9724,N_8122,N_8062);
nor U9725 (N_9725,N_8146,N_8095);
and U9726 (N_9726,N_8320,N_8571);
nand U9727 (N_9727,N_8752,N_8519);
nand U9728 (N_9728,N_8759,N_8727);
or U9729 (N_9729,N_8591,N_8285);
nand U9730 (N_9730,N_8227,N_8490);
nor U9731 (N_9731,N_8932,N_8580);
nor U9732 (N_9732,N_8098,N_8679);
or U9733 (N_9733,N_8671,N_8221);
or U9734 (N_9734,N_8647,N_8240);
and U9735 (N_9735,N_8525,N_8331);
and U9736 (N_9736,N_8258,N_8608);
nor U9737 (N_9737,N_8043,N_8965);
nand U9738 (N_9738,N_8673,N_8201);
or U9739 (N_9739,N_8294,N_8700);
or U9740 (N_9740,N_8556,N_8374);
and U9741 (N_9741,N_8515,N_8604);
nand U9742 (N_9742,N_8664,N_8306);
and U9743 (N_9743,N_8553,N_8092);
or U9744 (N_9744,N_8156,N_8164);
or U9745 (N_9745,N_8237,N_8208);
nor U9746 (N_9746,N_8296,N_8855);
and U9747 (N_9747,N_8554,N_8031);
or U9748 (N_9748,N_8906,N_8406);
or U9749 (N_9749,N_8996,N_8762);
nand U9750 (N_9750,N_8123,N_8676);
nor U9751 (N_9751,N_8689,N_8466);
nand U9752 (N_9752,N_8033,N_8245);
nor U9753 (N_9753,N_8427,N_8493);
nor U9754 (N_9754,N_8184,N_8171);
nor U9755 (N_9755,N_8242,N_8126);
nand U9756 (N_9756,N_8173,N_8551);
nand U9757 (N_9757,N_8528,N_8584);
nor U9758 (N_9758,N_8171,N_8207);
nand U9759 (N_9759,N_8979,N_8291);
and U9760 (N_9760,N_8503,N_8778);
nand U9761 (N_9761,N_8759,N_8008);
or U9762 (N_9762,N_8863,N_8136);
or U9763 (N_9763,N_8003,N_8111);
nand U9764 (N_9764,N_8526,N_8392);
or U9765 (N_9765,N_8995,N_8390);
nor U9766 (N_9766,N_8388,N_8088);
nand U9767 (N_9767,N_8681,N_8077);
nor U9768 (N_9768,N_8087,N_8644);
or U9769 (N_9769,N_8298,N_8721);
or U9770 (N_9770,N_8545,N_8483);
nand U9771 (N_9771,N_8780,N_8081);
nor U9772 (N_9772,N_8393,N_8104);
or U9773 (N_9773,N_8738,N_8158);
nand U9774 (N_9774,N_8870,N_8136);
nor U9775 (N_9775,N_8930,N_8421);
nor U9776 (N_9776,N_8992,N_8183);
nor U9777 (N_9777,N_8270,N_8460);
or U9778 (N_9778,N_8559,N_8444);
or U9779 (N_9779,N_8474,N_8775);
nor U9780 (N_9780,N_8083,N_8626);
nor U9781 (N_9781,N_8465,N_8467);
and U9782 (N_9782,N_8002,N_8598);
and U9783 (N_9783,N_8259,N_8188);
nand U9784 (N_9784,N_8529,N_8675);
nand U9785 (N_9785,N_8426,N_8941);
or U9786 (N_9786,N_8814,N_8923);
nand U9787 (N_9787,N_8535,N_8787);
or U9788 (N_9788,N_8256,N_8946);
and U9789 (N_9789,N_8712,N_8782);
and U9790 (N_9790,N_8256,N_8112);
nor U9791 (N_9791,N_8564,N_8107);
nor U9792 (N_9792,N_8517,N_8444);
or U9793 (N_9793,N_8182,N_8185);
and U9794 (N_9794,N_8728,N_8034);
nand U9795 (N_9795,N_8993,N_8538);
and U9796 (N_9796,N_8289,N_8829);
or U9797 (N_9797,N_8198,N_8325);
and U9798 (N_9798,N_8170,N_8365);
nand U9799 (N_9799,N_8578,N_8401);
nand U9800 (N_9800,N_8129,N_8221);
or U9801 (N_9801,N_8472,N_8505);
nor U9802 (N_9802,N_8719,N_8840);
and U9803 (N_9803,N_8594,N_8502);
and U9804 (N_9804,N_8584,N_8882);
nand U9805 (N_9805,N_8586,N_8723);
or U9806 (N_9806,N_8410,N_8454);
nand U9807 (N_9807,N_8951,N_8709);
nor U9808 (N_9808,N_8605,N_8428);
and U9809 (N_9809,N_8723,N_8961);
nand U9810 (N_9810,N_8513,N_8035);
or U9811 (N_9811,N_8237,N_8832);
and U9812 (N_9812,N_8076,N_8406);
or U9813 (N_9813,N_8191,N_8136);
or U9814 (N_9814,N_8871,N_8306);
nor U9815 (N_9815,N_8091,N_8052);
nand U9816 (N_9816,N_8294,N_8736);
nor U9817 (N_9817,N_8101,N_8460);
nand U9818 (N_9818,N_8977,N_8437);
nor U9819 (N_9819,N_8822,N_8232);
nand U9820 (N_9820,N_8415,N_8837);
nand U9821 (N_9821,N_8962,N_8505);
and U9822 (N_9822,N_8550,N_8777);
or U9823 (N_9823,N_8551,N_8760);
or U9824 (N_9824,N_8163,N_8961);
nor U9825 (N_9825,N_8271,N_8528);
or U9826 (N_9826,N_8535,N_8747);
nand U9827 (N_9827,N_8899,N_8618);
nor U9828 (N_9828,N_8847,N_8341);
or U9829 (N_9829,N_8688,N_8415);
or U9830 (N_9830,N_8836,N_8217);
and U9831 (N_9831,N_8643,N_8360);
and U9832 (N_9832,N_8141,N_8267);
nand U9833 (N_9833,N_8400,N_8569);
and U9834 (N_9834,N_8524,N_8572);
or U9835 (N_9835,N_8428,N_8366);
or U9836 (N_9836,N_8126,N_8467);
and U9837 (N_9837,N_8644,N_8664);
and U9838 (N_9838,N_8556,N_8383);
or U9839 (N_9839,N_8494,N_8132);
and U9840 (N_9840,N_8936,N_8334);
nand U9841 (N_9841,N_8887,N_8198);
nor U9842 (N_9842,N_8768,N_8565);
nand U9843 (N_9843,N_8537,N_8095);
nand U9844 (N_9844,N_8742,N_8381);
and U9845 (N_9845,N_8942,N_8329);
and U9846 (N_9846,N_8755,N_8192);
nand U9847 (N_9847,N_8266,N_8965);
nor U9848 (N_9848,N_8009,N_8731);
or U9849 (N_9849,N_8047,N_8920);
nand U9850 (N_9850,N_8373,N_8939);
and U9851 (N_9851,N_8876,N_8359);
or U9852 (N_9852,N_8212,N_8739);
or U9853 (N_9853,N_8494,N_8311);
nand U9854 (N_9854,N_8951,N_8067);
nand U9855 (N_9855,N_8825,N_8870);
nor U9856 (N_9856,N_8760,N_8166);
nand U9857 (N_9857,N_8868,N_8404);
and U9858 (N_9858,N_8437,N_8688);
and U9859 (N_9859,N_8056,N_8755);
or U9860 (N_9860,N_8804,N_8705);
and U9861 (N_9861,N_8769,N_8423);
or U9862 (N_9862,N_8141,N_8180);
and U9863 (N_9863,N_8625,N_8147);
nor U9864 (N_9864,N_8000,N_8386);
or U9865 (N_9865,N_8738,N_8774);
nand U9866 (N_9866,N_8823,N_8174);
nand U9867 (N_9867,N_8071,N_8527);
nand U9868 (N_9868,N_8578,N_8119);
nand U9869 (N_9869,N_8042,N_8433);
nor U9870 (N_9870,N_8485,N_8567);
nor U9871 (N_9871,N_8478,N_8918);
nand U9872 (N_9872,N_8662,N_8336);
or U9873 (N_9873,N_8903,N_8344);
nand U9874 (N_9874,N_8842,N_8797);
nor U9875 (N_9875,N_8721,N_8931);
or U9876 (N_9876,N_8724,N_8049);
nand U9877 (N_9877,N_8312,N_8225);
nand U9878 (N_9878,N_8181,N_8340);
nor U9879 (N_9879,N_8566,N_8569);
and U9880 (N_9880,N_8834,N_8307);
and U9881 (N_9881,N_8154,N_8317);
or U9882 (N_9882,N_8440,N_8779);
or U9883 (N_9883,N_8545,N_8728);
and U9884 (N_9884,N_8682,N_8463);
or U9885 (N_9885,N_8304,N_8107);
or U9886 (N_9886,N_8431,N_8680);
or U9887 (N_9887,N_8327,N_8824);
nor U9888 (N_9888,N_8632,N_8620);
and U9889 (N_9889,N_8554,N_8532);
or U9890 (N_9890,N_8814,N_8545);
or U9891 (N_9891,N_8048,N_8121);
or U9892 (N_9892,N_8587,N_8552);
nand U9893 (N_9893,N_8198,N_8106);
nand U9894 (N_9894,N_8421,N_8855);
or U9895 (N_9895,N_8162,N_8917);
nand U9896 (N_9896,N_8307,N_8854);
and U9897 (N_9897,N_8005,N_8576);
or U9898 (N_9898,N_8497,N_8764);
and U9899 (N_9899,N_8176,N_8997);
or U9900 (N_9900,N_8944,N_8507);
nand U9901 (N_9901,N_8146,N_8477);
nand U9902 (N_9902,N_8211,N_8589);
nor U9903 (N_9903,N_8250,N_8873);
and U9904 (N_9904,N_8718,N_8553);
nor U9905 (N_9905,N_8723,N_8962);
or U9906 (N_9906,N_8617,N_8675);
nand U9907 (N_9907,N_8927,N_8610);
and U9908 (N_9908,N_8258,N_8149);
or U9909 (N_9909,N_8535,N_8504);
and U9910 (N_9910,N_8472,N_8146);
nor U9911 (N_9911,N_8893,N_8783);
and U9912 (N_9912,N_8250,N_8364);
and U9913 (N_9913,N_8886,N_8255);
and U9914 (N_9914,N_8460,N_8352);
nor U9915 (N_9915,N_8035,N_8276);
nor U9916 (N_9916,N_8205,N_8015);
nand U9917 (N_9917,N_8717,N_8929);
nand U9918 (N_9918,N_8438,N_8814);
and U9919 (N_9919,N_8589,N_8717);
or U9920 (N_9920,N_8233,N_8185);
nor U9921 (N_9921,N_8488,N_8080);
nor U9922 (N_9922,N_8680,N_8336);
and U9923 (N_9923,N_8685,N_8987);
nor U9924 (N_9924,N_8649,N_8742);
or U9925 (N_9925,N_8895,N_8608);
or U9926 (N_9926,N_8152,N_8581);
nand U9927 (N_9927,N_8408,N_8132);
nor U9928 (N_9928,N_8810,N_8505);
or U9929 (N_9929,N_8585,N_8805);
and U9930 (N_9930,N_8469,N_8518);
nand U9931 (N_9931,N_8417,N_8634);
nand U9932 (N_9932,N_8148,N_8053);
or U9933 (N_9933,N_8680,N_8286);
nor U9934 (N_9934,N_8946,N_8348);
or U9935 (N_9935,N_8424,N_8408);
and U9936 (N_9936,N_8171,N_8645);
nor U9937 (N_9937,N_8976,N_8992);
or U9938 (N_9938,N_8264,N_8789);
or U9939 (N_9939,N_8870,N_8225);
nor U9940 (N_9940,N_8762,N_8690);
and U9941 (N_9941,N_8510,N_8590);
and U9942 (N_9942,N_8299,N_8487);
and U9943 (N_9943,N_8513,N_8074);
and U9944 (N_9944,N_8862,N_8866);
nand U9945 (N_9945,N_8904,N_8299);
nand U9946 (N_9946,N_8982,N_8053);
nand U9947 (N_9947,N_8605,N_8899);
or U9948 (N_9948,N_8293,N_8925);
or U9949 (N_9949,N_8249,N_8498);
or U9950 (N_9950,N_8666,N_8157);
and U9951 (N_9951,N_8773,N_8181);
or U9952 (N_9952,N_8230,N_8276);
and U9953 (N_9953,N_8301,N_8059);
nand U9954 (N_9954,N_8617,N_8478);
or U9955 (N_9955,N_8912,N_8137);
and U9956 (N_9956,N_8007,N_8644);
or U9957 (N_9957,N_8124,N_8110);
or U9958 (N_9958,N_8569,N_8570);
or U9959 (N_9959,N_8294,N_8854);
nand U9960 (N_9960,N_8380,N_8298);
nand U9961 (N_9961,N_8602,N_8118);
nand U9962 (N_9962,N_8942,N_8158);
or U9963 (N_9963,N_8670,N_8693);
nand U9964 (N_9964,N_8590,N_8776);
nand U9965 (N_9965,N_8024,N_8136);
nor U9966 (N_9966,N_8299,N_8501);
or U9967 (N_9967,N_8320,N_8927);
and U9968 (N_9968,N_8922,N_8437);
nor U9969 (N_9969,N_8517,N_8759);
nand U9970 (N_9970,N_8695,N_8308);
xnor U9971 (N_9971,N_8878,N_8846);
nor U9972 (N_9972,N_8308,N_8184);
and U9973 (N_9973,N_8238,N_8393);
and U9974 (N_9974,N_8458,N_8630);
nor U9975 (N_9975,N_8973,N_8598);
nor U9976 (N_9976,N_8528,N_8554);
nand U9977 (N_9977,N_8433,N_8947);
nand U9978 (N_9978,N_8932,N_8024);
nor U9979 (N_9979,N_8172,N_8358);
or U9980 (N_9980,N_8358,N_8871);
nor U9981 (N_9981,N_8152,N_8183);
nor U9982 (N_9982,N_8003,N_8807);
or U9983 (N_9983,N_8391,N_8808);
and U9984 (N_9984,N_8323,N_8516);
or U9985 (N_9985,N_8658,N_8955);
and U9986 (N_9986,N_8006,N_8121);
or U9987 (N_9987,N_8792,N_8182);
and U9988 (N_9988,N_8324,N_8922);
or U9989 (N_9989,N_8323,N_8237);
and U9990 (N_9990,N_8446,N_8742);
nand U9991 (N_9991,N_8434,N_8349);
nand U9992 (N_9992,N_8541,N_8922);
and U9993 (N_9993,N_8217,N_8889);
nand U9994 (N_9994,N_8834,N_8603);
nand U9995 (N_9995,N_8207,N_8694);
nand U9996 (N_9996,N_8632,N_8190);
or U9997 (N_9997,N_8765,N_8411);
nand U9998 (N_9998,N_8850,N_8547);
or U9999 (N_9999,N_8976,N_8664);
nor UO_0 (O_0,N_9238,N_9075);
nand UO_1 (O_1,N_9486,N_9466);
and UO_2 (O_2,N_9590,N_9972);
nor UO_3 (O_3,N_9498,N_9838);
nand UO_4 (O_4,N_9257,N_9183);
and UO_5 (O_5,N_9686,N_9336);
nand UO_6 (O_6,N_9845,N_9579);
and UO_7 (O_7,N_9279,N_9405);
xor UO_8 (O_8,N_9872,N_9292);
nand UO_9 (O_9,N_9180,N_9837);
and UO_10 (O_10,N_9153,N_9791);
nor UO_11 (O_11,N_9555,N_9148);
or UO_12 (O_12,N_9120,N_9668);
nand UO_13 (O_13,N_9309,N_9922);
nand UO_14 (O_14,N_9777,N_9174);
or UO_15 (O_15,N_9417,N_9918);
and UO_16 (O_16,N_9287,N_9199);
and UO_17 (O_17,N_9364,N_9000);
nand UO_18 (O_18,N_9423,N_9484);
nor UO_19 (O_19,N_9981,N_9418);
or UO_20 (O_20,N_9687,N_9913);
nand UO_21 (O_21,N_9820,N_9600);
or UO_22 (O_22,N_9210,N_9568);
xor UO_23 (O_23,N_9878,N_9780);
nor UO_24 (O_24,N_9882,N_9227);
or UO_25 (O_25,N_9809,N_9784);
and UO_26 (O_26,N_9944,N_9294);
nand UO_27 (O_27,N_9750,N_9827);
and UO_28 (O_28,N_9375,N_9302);
or UO_29 (O_29,N_9306,N_9860);
and UO_30 (O_30,N_9900,N_9269);
nand UO_31 (O_31,N_9663,N_9304);
and UO_32 (O_32,N_9112,N_9281);
and UO_33 (O_33,N_9818,N_9501);
nand UO_34 (O_34,N_9795,N_9111);
nor UO_35 (O_35,N_9458,N_9132);
and UO_36 (O_36,N_9718,N_9400);
or UO_37 (O_37,N_9066,N_9695);
nor UO_38 (O_38,N_9530,N_9587);
nor UO_39 (O_39,N_9315,N_9758);
and UO_40 (O_40,N_9320,N_9940);
and UO_41 (O_41,N_9689,N_9298);
or UO_42 (O_42,N_9342,N_9467);
and UO_43 (O_43,N_9850,N_9139);
nor UO_44 (O_44,N_9003,N_9631);
nand UO_45 (O_45,N_9046,N_9463);
and UO_46 (O_46,N_9394,N_9581);
and UO_47 (O_47,N_9673,N_9268);
nor UO_48 (O_48,N_9403,N_9543);
and UO_49 (O_49,N_9688,N_9738);
nor UO_50 (O_50,N_9973,N_9789);
nor UO_51 (O_51,N_9170,N_9052);
nand UO_52 (O_52,N_9121,N_9327);
nor UO_53 (O_53,N_9214,N_9636);
or UO_54 (O_54,N_9879,N_9915);
nand UO_55 (O_55,N_9176,N_9022);
and UO_56 (O_56,N_9651,N_9021);
nand UO_57 (O_57,N_9493,N_9436);
and UO_58 (O_58,N_9246,N_9189);
nand UO_59 (O_59,N_9805,N_9071);
nor UO_60 (O_60,N_9062,N_9027);
and UO_61 (O_61,N_9407,N_9144);
and UO_62 (O_62,N_9124,N_9316);
and UO_63 (O_63,N_9811,N_9782);
and UO_64 (O_64,N_9875,N_9717);
nor UO_65 (O_65,N_9070,N_9841);
and UO_66 (O_66,N_9365,N_9151);
nand UO_67 (O_67,N_9649,N_9218);
nand UO_68 (O_68,N_9094,N_9964);
or UO_69 (O_69,N_9479,N_9605);
and UO_70 (O_70,N_9938,N_9025);
nand UO_71 (O_71,N_9426,N_9353);
nor UO_72 (O_72,N_9813,N_9357);
nand UO_73 (O_73,N_9080,N_9201);
or UO_74 (O_74,N_9993,N_9444);
and UO_75 (O_75,N_9943,N_9006);
or UO_76 (O_76,N_9997,N_9868);
nand UO_77 (O_77,N_9095,N_9736);
and UO_78 (O_78,N_9776,N_9886);
nor UO_79 (O_79,N_9657,N_9010);
nor UO_80 (O_80,N_9472,N_9457);
nor UO_81 (O_81,N_9917,N_9039);
and UO_82 (O_82,N_9290,N_9044);
or UO_83 (O_83,N_9354,N_9296);
nor UO_84 (O_84,N_9241,N_9130);
nand UO_85 (O_85,N_9952,N_9164);
or UO_86 (O_86,N_9544,N_9936);
nand UO_87 (O_87,N_9710,N_9732);
or UO_88 (O_88,N_9951,N_9197);
nand UO_89 (O_89,N_9172,N_9009);
or UO_90 (O_90,N_9234,N_9090);
or UO_91 (O_91,N_9017,N_9715);
nor UO_92 (O_92,N_9550,N_9100);
xor UO_93 (O_93,N_9894,N_9666);
nand UO_94 (O_94,N_9464,N_9435);
nand UO_95 (O_95,N_9671,N_9286);
and UO_96 (O_96,N_9561,N_9096);
or UO_97 (O_97,N_9216,N_9098);
or UO_98 (O_98,N_9415,N_9935);
or UO_99 (O_99,N_9230,N_9803);
nand UO_100 (O_100,N_9051,N_9976);
or UO_101 (O_101,N_9907,N_9473);
nor UO_102 (O_102,N_9142,N_9889);
nor UO_103 (O_103,N_9157,N_9669);
and UO_104 (O_104,N_9674,N_9728);
nand UO_105 (O_105,N_9508,N_9723);
nor UO_106 (O_106,N_9001,N_9564);
nand UO_107 (O_107,N_9185,N_9541);
or UO_108 (O_108,N_9380,N_9162);
nor UO_109 (O_109,N_9761,N_9042);
nor UO_110 (O_110,N_9988,N_9680);
nor UO_111 (O_111,N_9252,N_9184);
and UO_112 (O_112,N_9746,N_9884);
and UO_113 (O_113,N_9140,N_9652);
or UO_114 (O_114,N_9529,N_9667);
or UO_115 (O_115,N_9333,N_9540);
nand UO_116 (O_116,N_9087,N_9491);
nand UO_117 (O_117,N_9076,N_9612);
nor UO_118 (O_118,N_9574,N_9043);
or UO_119 (O_119,N_9836,N_9069);
nor UO_120 (O_120,N_9725,N_9378);
nand UO_121 (O_121,N_9735,N_9707);
nor UO_122 (O_122,N_9460,N_9105);
nand UO_123 (O_123,N_9510,N_9566);
and UO_124 (O_124,N_9851,N_9248);
nand UO_125 (O_125,N_9921,N_9711);
nor UO_126 (O_126,N_9618,N_9452);
and UO_127 (O_127,N_9977,N_9928);
nand UO_128 (O_128,N_9825,N_9389);
nor UO_129 (O_129,N_9200,N_9503);
nor UO_130 (O_130,N_9855,N_9202);
nor UO_131 (O_131,N_9792,N_9549);
and UO_132 (O_132,N_9571,N_9509);
nor UO_133 (O_133,N_9276,N_9726);
and UO_134 (O_134,N_9408,N_9262);
nor UO_135 (O_135,N_9358,N_9932);
and UO_136 (O_136,N_9584,N_9527);
nor UO_137 (O_137,N_9756,N_9368);
nand UO_138 (O_138,N_9429,N_9363);
nand UO_139 (O_139,N_9237,N_9862);
or UO_140 (O_140,N_9152,N_9954);
or UO_141 (O_141,N_9606,N_9034);
nand UO_142 (O_142,N_9611,N_9459);
or UO_143 (O_143,N_9329,N_9175);
or UO_144 (O_144,N_9482,N_9854);
nor UO_145 (O_145,N_9496,N_9297);
nand UO_146 (O_146,N_9961,N_9401);
and UO_147 (O_147,N_9194,N_9817);
nand UO_148 (O_148,N_9545,N_9712);
nor UO_149 (O_149,N_9767,N_9171);
and UO_150 (O_150,N_9299,N_9620);
and UO_151 (O_151,N_9583,N_9312);
and UO_152 (O_152,N_9546,N_9195);
and UO_153 (O_153,N_9942,N_9821);
and UO_154 (O_154,N_9567,N_9513);
and UO_155 (O_155,N_9059,N_9433);
or UO_156 (O_156,N_9804,N_9522);
xor UO_157 (O_157,N_9523,N_9766);
or UO_158 (O_158,N_9923,N_9578);
and UO_159 (O_159,N_9672,N_9236);
and UO_160 (O_160,N_9274,N_9266);
and UO_161 (O_161,N_9588,N_9639);
or UO_162 (O_162,N_9582,N_9926);
xor UO_163 (O_163,N_9664,N_9058);
and UO_164 (O_164,N_9867,N_9117);
nand UO_165 (O_165,N_9849,N_9154);
or UO_166 (O_166,N_9440,N_9863);
or UO_167 (O_167,N_9119,N_9901);
nand UO_168 (O_168,N_9409,N_9012);
nand UO_169 (O_169,N_9278,N_9122);
and UO_170 (O_170,N_9370,N_9225);
and UO_171 (O_171,N_9648,N_9437);
or UO_172 (O_172,N_9771,N_9073);
or UO_173 (O_173,N_9992,N_9330);
nor UO_174 (O_174,N_9681,N_9019);
or UO_175 (O_175,N_9797,N_9514);
nor UO_176 (O_176,N_9957,N_9243);
and UO_177 (O_177,N_9719,N_9026);
or UO_178 (O_178,N_9764,N_9990);
nor UO_179 (O_179,N_9832,N_9441);
nand UO_180 (O_180,N_9413,N_9843);
xnor UO_181 (O_181,N_9307,N_9374);
or UO_182 (O_182,N_9968,N_9844);
and UO_183 (O_183,N_9824,N_9790);
nor UO_184 (O_184,N_9799,N_9233);
nor UO_185 (O_185,N_9453,N_9118);
and UO_186 (O_186,N_9348,N_9709);
nor UO_187 (O_187,N_9125,N_9888);
and UO_188 (O_188,N_9753,N_9659);
and UO_189 (O_189,N_9643,N_9676);
or UO_190 (O_190,N_9812,N_9303);
nor UO_191 (O_191,N_9684,N_9301);
and UO_192 (O_192,N_9173,N_9924);
nand UO_193 (O_193,N_9074,N_9211);
nor UO_194 (O_194,N_9984,N_9904);
and UO_195 (O_195,N_9891,N_9391);
nand UO_196 (O_196,N_9128,N_9222);
or UO_197 (O_197,N_9321,N_9018);
nor UO_198 (O_198,N_9318,N_9506);
and UO_199 (O_199,N_9332,N_9633);
nand UO_200 (O_200,N_9902,N_9032);
or UO_201 (O_201,N_9589,N_9806);
or UO_202 (O_202,N_9469,N_9536);
or UO_203 (O_203,N_9630,N_9187);
or UO_204 (O_204,N_9341,N_9533);
or UO_205 (O_205,N_9226,N_9215);
nand UO_206 (O_206,N_9406,N_9617);
nand UO_207 (O_207,N_9311,N_9896);
and UO_208 (O_208,N_9305,N_9203);
nand UO_209 (O_209,N_9192,N_9865);
nand UO_210 (O_210,N_9272,N_9691);
nand UO_211 (O_211,N_9532,N_9123);
nor UO_212 (O_212,N_9056,N_9344);
nand UO_213 (O_213,N_9335,N_9677);
and UO_214 (O_214,N_9956,N_9786);
and UO_215 (O_215,N_9049,N_9864);
nor UO_216 (O_216,N_9283,N_9787);
nand UO_217 (O_217,N_9740,N_9656);
or UO_218 (O_218,N_9774,N_9859);
and UO_219 (O_219,N_9616,N_9892);
xor UO_220 (O_220,N_9704,N_9737);
nand UO_221 (O_221,N_9511,N_9840);
and UO_222 (O_222,N_9037,N_9377);
or UO_223 (O_223,N_9393,N_9240);
nand UO_224 (O_224,N_9937,N_9228);
and UO_225 (O_225,N_9562,N_9439);
or UO_226 (O_226,N_9165,N_9250);
nand UO_227 (O_227,N_9903,N_9819);
nand UO_228 (O_228,N_9586,N_9188);
or UO_229 (O_229,N_9356,N_9492);
and UO_230 (O_230,N_9325,N_9431);
and UO_231 (O_231,N_9137,N_9271);
nand UO_232 (O_232,N_9950,N_9597);
or UO_233 (O_233,N_9455,N_9699);
nand UO_234 (O_234,N_9016,N_9592);
nand UO_235 (O_235,N_9392,N_9480);
or UO_236 (O_236,N_9534,N_9390);
and UO_237 (O_237,N_9067,N_9632);
and UO_238 (O_238,N_9885,N_9623);
nor UO_239 (O_239,N_9412,N_9594);
and UO_240 (O_240,N_9637,N_9793);
nor UO_241 (O_241,N_9270,N_9906);
nand UO_242 (O_242,N_9313,N_9823);
nor UO_243 (O_243,N_9528,N_9654);
nand UO_244 (O_244,N_9982,N_9399);
and UO_245 (O_245,N_9739,N_9499);
nand UO_246 (O_246,N_9899,N_9232);
nand UO_247 (O_247,N_9224,N_9384);
xor UO_248 (O_248,N_9385,N_9519);
and UO_249 (O_249,N_9833,N_9846);
nor UO_250 (O_250,N_9595,N_9770);
or UO_251 (O_251,N_9524,N_9502);
nor UO_252 (O_252,N_9743,N_9221);
nand UO_253 (O_253,N_9072,N_9101);
nand UO_254 (O_254,N_9983,N_9267);
or UO_255 (O_255,N_9995,N_9449);
nand UO_256 (O_256,N_9229,N_9989);
or UO_257 (O_257,N_9470,N_9602);
nor UO_258 (O_258,N_9490,N_9223);
nor UO_259 (O_259,N_9505,N_9317);
or UO_260 (O_260,N_9880,N_9871);
or UO_261 (O_261,N_9036,N_9929);
and UO_262 (O_262,N_9115,N_9217);
nor UO_263 (O_263,N_9816,N_9166);
nand UO_264 (O_264,N_9538,N_9638);
nand UO_265 (O_265,N_9382,N_9347);
or UO_266 (O_266,N_9839,N_9461);
and UO_267 (O_267,N_9714,N_9295);
or UO_268 (O_268,N_9661,N_9488);
nor UO_269 (O_269,N_9476,N_9186);
and UO_270 (O_270,N_9376,N_9077);
or UO_271 (O_271,N_9969,N_9149);
or UO_272 (O_272,N_9763,N_9518);
or UO_273 (O_273,N_9696,N_9085);
and UO_274 (O_274,N_9856,N_9554);
and UO_275 (O_275,N_9191,N_9081);
or UO_276 (O_276,N_9319,N_9834);
nand UO_277 (O_277,N_9655,N_9177);
and UO_278 (O_278,N_9068,N_9108);
and UO_279 (O_279,N_9722,N_9822);
nor UO_280 (O_280,N_9873,N_9883);
nor UO_281 (O_281,N_9783,N_9798);
nor UO_282 (O_282,N_9471,N_9702);
nor UO_283 (O_283,N_9323,N_9093);
nor UO_284 (O_284,N_9448,N_9570);
nor UO_285 (O_285,N_9553,N_9733);
nor UO_286 (O_286,N_9563,N_9011);
nand UO_287 (O_287,N_9542,N_9958);
and UO_288 (O_288,N_9345,N_9360);
nand UO_289 (O_289,N_9193,N_9745);
nor UO_290 (O_290,N_9261,N_9023);
or UO_291 (O_291,N_9099,N_9462);
and UO_292 (O_292,N_9454,N_9547);
or UO_293 (O_293,N_9031,N_9731);
and UO_294 (O_294,N_9349,N_9744);
nand UO_295 (O_295,N_9014,N_9456);
and UO_296 (O_296,N_9285,N_9451);
and UO_297 (O_297,N_9251,N_9665);
nand UO_298 (O_298,N_9640,N_9960);
nor UO_299 (O_299,N_9404,N_9551);
nand UO_300 (O_300,N_9500,N_9963);
nand UO_301 (O_301,N_9328,N_9607);
nor UO_302 (O_302,N_9662,N_9015);
nand UO_303 (O_303,N_9552,N_9483);
and UO_304 (O_304,N_9577,N_9359);
or UO_305 (O_305,N_9495,N_9697);
or UO_306 (O_306,N_9231,N_9531);
and UO_307 (O_307,N_9653,N_9701);
nor UO_308 (O_308,N_9082,N_9870);
or UO_309 (O_309,N_9916,N_9604);
or UO_310 (O_310,N_9198,N_9035);
nand UO_311 (O_311,N_9948,N_9007);
nor UO_312 (O_312,N_9213,N_9572);
nand UO_313 (O_313,N_9999,N_9078);
nor UO_314 (O_314,N_9835,N_9040);
and UO_315 (O_315,N_9994,N_9720);
or UO_316 (O_316,N_9986,N_9253);
and UO_317 (O_317,N_9422,N_9881);
nor UO_318 (O_318,N_9383,N_9730);
and UO_319 (O_319,N_9371,N_9084);
nand UO_320 (O_320,N_9537,N_9603);
and UO_321 (O_321,N_9548,N_9249);
and UO_322 (O_322,N_9160,N_9324);
or UO_323 (O_323,N_9996,N_9614);
nand UO_324 (O_324,N_9092,N_9351);
nand UO_325 (O_325,N_9178,N_9381);
nand UO_326 (O_326,N_9102,N_9933);
nor UO_327 (O_327,N_9494,N_9979);
or UO_328 (O_328,N_9497,N_9182);
and UO_329 (O_329,N_9289,N_9516);
or UO_330 (O_330,N_9398,N_9800);
and UO_331 (O_331,N_9421,N_9755);
nor UO_332 (O_332,N_9033,N_9361);
nand UO_333 (O_333,N_9340,N_9772);
and UO_334 (O_334,N_9350,N_9779);
nand UO_335 (O_335,N_9310,N_9559);
or UO_336 (O_336,N_9047,N_9974);
and UO_337 (O_337,N_9858,N_9445);
and UO_338 (O_338,N_9338,N_9450);
nand UO_339 (O_339,N_9395,N_9326);
nor UO_340 (O_340,N_9212,N_9038);
nor UO_341 (O_341,N_9914,N_9775);
or UO_342 (O_342,N_9877,N_9920);
nand UO_343 (O_343,N_9005,N_9866);
nor UO_344 (O_344,N_9028,N_9599);
or UO_345 (O_345,N_9369,N_9355);
and UO_346 (O_346,N_9131,N_9721);
nor UO_347 (O_347,N_9959,N_9438);
or UO_348 (O_348,N_9282,N_9158);
nand UO_349 (O_349,N_9129,N_9086);
nand UO_350 (O_350,N_9646,N_9520);
or UO_351 (O_351,N_9810,N_9893);
or UO_352 (O_352,N_9678,N_9754);
nor UO_353 (O_353,N_9362,N_9145);
and UO_354 (O_354,N_9205,N_9953);
or UO_355 (O_355,N_9489,N_9163);
nor UO_356 (O_356,N_9768,N_9742);
nand UO_357 (O_357,N_9991,N_9379);
and UO_358 (O_358,N_9343,N_9708);
or UO_359 (O_359,N_9558,N_9475);
and UO_360 (O_360,N_9474,N_9179);
and UO_361 (O_361,N_9402,N_9556);
and UO_362 (O_362,N_9419,N_9367);
or UO_363 (O_363,N_9919,N_9635);
xnor UO_364 (O_364,N_9209,N_9945);
and UO_365 (O_365,N_9741,N_9970);
nand UO_366 (O_366,N_9083,N_9366);
and UO_367 (O_367,N_9626,N_9314);
and UO_368 (O_368,N_9265,N_9557);
nor UO_369 (O_369,N_9966,N_9247);
and UO_370 (O_370,N_9258,N_9430);
nand UO_371 (O_371,N_9927,N_9239);
and UO_372 (O_372,N_9930,N_9055);
nand UO_373 (O_373,N_9416,N_9387);
or UO_374 (O_374,N_9946,N_9598);
nor UO_375 (O_375,N_9831,N_9693);
nor UO_376 (O_376,N_9619,N_9934);
or UO_377 (O_377,N_9156,N_9339);
nand UO_378 (O_378,N_9807,N_9065);
and UO_379 (O_379,N_9079,N_9255);
or UO_380 (O_380,N_9373,N_9887);
nand UO_381 (O_381,N_9045,N_9245);
nor UO_382 (O_382,N_9135,N_9002);
and UO_383 (O_383,N_9106,N_9104);
nor UO_384 (O_384,N_9781,N_9670);
nor UO_385 (O_385,N_9155,N_9425);
or UO_386 (O_386,N_9748,N_9751);
or UO_387 (O_387,N_9971,N_9219);
or UO_388 (O_388,N_9091,N_9912);
and UO_389 (O_389,N_9207,N_9585);
nand UO_390 (O_390,N_9909,N_9847);
nor UO_391 (O_391,N_9048,N_9987);
or UO_392 (O_392,N_9828,N_9280);
and UO_393 (O_393,N_9911,N_9698);
or UO_394 (O_394,N_9752,N_9565);
or UO_395 (O_395,N_9220,N_9388);
or UO_396 (O_396,N_9650,N_9628);
nand UO_397 (O_397,N_9609,N_9580);
and UO_398 (O_398,N_9277,N_9507);
nor UO_399 (O_399,N_9288,N_9869);
nor UO_400 (O_400,N_9446,N_9759);
nor UO_401 (O_401,N_9939,N_9254);
nand UO_402 (O_402,N_9658,N_9396);
nor UO_403 (O_403,N_9814,N_9346);
nor UO_404 (O_404,N_9263,N_9110);
nand UO_405 (O_405,N_9024,N_9168);
nor UO_406 (O_406,N_9700,N_9898);
nand UO_407 (O_407,N_9621,N_9291);
or UO_408 (O_408,N_9727,N_9244);
and UO_409 (O_409,N_9190,N_9284);
nand UO_410 (O_410,N_9608,N_9808);
and UO_411 (O_411,N_9114,N_9949);
or UO_412 (O_412,N_9647,N_9041);
and UO_413 (O_413,N_9517,N_9029);
nand UO_414 (O_414,N_9064,N_9679);
nand UO_415 (O_415,N_9300,N_9925);
nand UO_416 (O_416,N_9103,N_9716);
and UO_417 (O_417,N_9874,N_9985);
nor UO_418 (O_418,N_9420,N_9682);
and UO_419 (O_419,N_9256,N_9905);
nand UO_420 (O_420,N_9465,N_9613);
nor UO_421 (O_421,N_9829,N_9136);
and UO_422 (O_422,N_9428,N_9848);
or UO_423 (O_423,N_9908,N_9685);
nand UO_424 (O_424,N_9694,N_9645);
nand UO_425 (O_425,N_9634,N_9683);
or UO_426 (O_426,N_9260,N_9975);
and UO_427 (O_427,N_9167,N_9539);
nor UO_428 (O_428,N_9447,N_9801);
or UO_429 (O_429,N_9424,N_9629);
nand UO_430 (O_430,N_9113,N_9411);
nand UO_431 (O_431,N_9169,N_9150);
or UO_432 (O_432,N_9747,N_9206);
nor UO_433 (O_433,N_9061,N_9126);
nor UO_434 (O_434,N_9147,N_9978);
and UO_435 (O_435,N_9852,N_9627);
nand UO_436 (O_436,N_9208,N_9138);
or UO_437 (O_437,N_9515,N_9762);
nor UO_438 (O_438,N_9008,N_9641);
and UO_439 (O_439,N_9088,N_9050);
nor UO_440 (O_440,N_9760,N_9512);
nand UO_441 (O_441,N_9487,N_9706);
and UO_442 (O_442,N_9773,N_9410);
nor UO_443 (O_443,N_9235,N_9372);
nand UO_444 (O_444,N_9861,N_9259);
nor UO_445 (O_445,N_9196,N_9432);
or UO_446 (O_446,N_9794,N_9352);
or UO_447 (O_447,N_9596,N_9644);
or UO_448 (O_448,N_9876,N_9013);
or UO_449 (O_449,N_9030,N_9967);
nor UO_450 (O_450,N_9097,N_9690);
or UO_451 (O_451,N_9397,N_9442);
and UO_452 (O_452,N_9573,N_9890);
or UO_453 (O_453,N_9133,N_9109);
and UO_454 (O_454,N_9089,N_9624);
and UO_455 (O_455,N_9713,N_9116);
nand UO_456 (O_456,N_9264,N_9796);
and UO_457 (O_457,N_9560,N_9788);
nor UO_458 (O_458,N_9535,N_9308);
nor UO_459 (O_459,N_9729,N_9443);
and UO_460 (O_460,N_9143,N_9337);
and UO_461 (O_461,N_9322,N_9830);
nor UO_462 (O_462,N_9477,N_9275);
nand UO_463 (O_463,N_9063,N_9895);
nor UO_464 (O_464,N_9057,N_9159);
or UO_465 (O_465,N_9675,N_9610);
and UO_466 (O_466,N_9575,N_9427);
nand UO_467 (O_467,N_9593,N_9526);
nand UO_468 (O_468,N_9749,N_9053);
nand UO_469 (O_469,N_9910,N_9434);
nand UO_470 (O_470,N_9334,N_9802);
nand UO_471 (O_471,N_9724,N_9734);
nor UO_472 (O_472,N_9504,N_9965);
nand UO_473 (O_473,N_9204,N_9569);
or UO_474 (O_474,N_9692,N_9468);
and UO_475 (O_475,N_9757,N_9842);
nand UO_476 (O_476,N_9181,N_9955);
and UO_477 (O_477,N_9778,N_9521);
or UO_478 (O_478,N_9591,N_9857);
nand UO_479 (O_479,N_9897,N_9931);
or UO_480 (O_480,N_9941,N_9962);
nor UO_481 (O_481,N_9054,N_9947);
and UO_482 (O_482,N_9293,N_9141);
and UO_483 (O_483,N_9127,N_9622);
and UO_484 (O_484,N_9785,N_9769);
nand UO_485 (O_485,N_9004,N_9525);
and UO_486 (O_486,N_9386,N_9331);
or UO_487 (O_487,N_9107,N_9485);
xnor UO_488 (O_488,N_9601,N_9134);
or UO_489 (O_489,N_9060,N_9815);
nor UO_490 (O_490,N_9765,N_9980);
and UO_491 (O_491,N_9478,N_9660);
nor UO_492 (O_492,N_9703,N_9642);
or UO_493 (O_493,N_9826,N_9020);
and UO_494 (O_494,N_9625,N_9615);
and UO_495 (O_495,N_9481,N_9414);
or UO_496 (O_496,N_9853,N_9576);
nor UO_497 (O_497,N_9705,N_9273);
nor UO_498 (O_498,N_9242,N_9998);
and UO_499 (O_499,N_9161,N_9146);
nor UO_500 (O_500,N_9398,N_9665);
and UO_501 (O_501,N_9975,N_9086);
nor UO_502 (O_502,N_9637,N_9415);
nor UO_503 (O_503,N_9635,N_9674);
nor UO_504 (O_504,N_9235,N_9797);
nand UO_505 (O_505,N_9627,N_9848);
nor UO_506 (O_506,N_9431,N_9937);
nand UO_507 (O_507,N_9398,N_9243);
nand UO_508 (O_508,N_9621,N_9412);
nand UO_509 (O_509,N_9022,N_9469);
nand UO_510 (O_510,N_9769,N_9638);
or UO_511 (O_511,N_9099,N_9124);
nor UO_512 (O_512,N_9159,N_9629);
nand UO_513 (O_513,N_9711,N_9662);
nand UO_514 (O_514,N_9135,N_9931);
nor UO_515 (O_515,N_9514,N_9326);
nand UO_516 (O_516,N_9030,N_9212);
nand UO_517 (O_517,N_9206,N_9616);
and UO_518 (O_518,N_9367,N_9555);
and UO_519 (O_519,N_9331,N_9589);
nor UO_520 (O_520,N_9951,N_9479);
or UO_521 (O_521,N_9251,N_9531);
nor UO_522 (O_522,N_9971,N_9860);
or UO_523 (O_523,N_9461,N_9929);
nor UO_524 (O_524,N_9716,N_9551);
or UO_525 (O_525,N_9053,N_9106);
and UO_526 (O_526,N_9930,N_9148);
or UO_527 (O_527,N_9995,N_9574);
or UO_528 (O_528,N_9169,N_9221);
or UO_529 (O_529,N_9076,N_9818);
and UO_530 (O_530,N_9173,N_9639);
nor UO_531 (O_531,N_9854,N_9452);
and UO_532 (O_532,N_9187,N_9965);
nor UO_533 (O_533,N_9000,N_9049);
and UO_534 (O_534,N_9982,N_9079);
nor UO_535 (O_535,N_9462,N_9585);
nor UO_536 (O_536,N_9725,N_9107);
or UO_537 (O_537,N_9854,N_9779);
nand UO_538 (O_538,N_9877,N_9930);
nor UO_539 (O_539,N_9066,N_9359);
and UO_540 (O_540,N_9687,N_9147);
and UO_541 (O_541,N_9947,N_9062);
and UO_542 (O_542,N_9565,N_9157);
nand UO_543 (O_543,N_9386,N_9729);
nand UO_544 (O_544,N_9416,N_9449);
and UO_545 (O_545,N_9544,N_9013);
and UO_546 (O_546,N_9259,N_9318);
nor UO_547 (O_547,N_9114,N_9217);
and UO_548 (O_548,N_9021,N_9731);
nand UO_549 (O_549,N_9908,N_9710);
and UO_550 (O_550,N_9615,N_9214);
and UO_551 (O_551,N_9020,N_9754);
and UO_552 (O_552,N_9513,N_9787);
and UO_553 (O_553,N_9912,N_9437);
nor UO_554 (O_554,N_9694,N_9918);
and UO_555 (O_555,N_9503,N_9090);
nand UO_556 (O_556,N_9244,N_9071);
nor UO_557 (O_557,N_9430,N_9928);
and UO_558 (O_558,N_9871,N_9036);
and UO_559 (O_559,N_9458,N_9200);
nor UO_560 (O_560,N_9294,N_9236);
and UO_561 (O_561,N_9342,N_9022);
nand UO_562 (O_562,N_9671,N_9534);
nor UO_563 (O_563,N_9839,N_9475);
nand UO_564 (O_564,N_9845,N_9044);
and UO_565 (O_565,N_9922,N_9733);
or UO_566 (O_566,N_9168,N_9415);
nor UO_567 (O_567,N_9146,N_9118);
or UO_568 (O_568,N_9499,N_9760);
nor UO_569 (O_569,N_9134,N_9543);
nor UO_570 (O_570,N_9716,N_9307);
nand UO_571 (O_571,N_9353,N_9486);
or UO_572 (O_572,N_9723,N_9329);
or UO_573 (O_573,N_9706,N_9104);
nand UO_574 (O_574,N_9817,N_9044);
nand UO_575 (O_575,N_9734,N_9657);
or UO_576 (O_576,N_9865,N_9789);
and UO_577 (O_577,N_9728,N_9103);
nor UO_578 (O_578,N_9509,N_9418);
and UO_579 (O_579,N_9490,N_9460);
xor UO_580 (O_580,N_9134,N_9322);
nor UO_581 (O_581,N_9029,N_9440);
or UO_582 (O_582,N_9232,N_9421);
and UO_583 (O_583,N_9015,N_9480);
and UO_584 (O_584,N_9082,N_9793);
nand UO_585 (O_585,N_9785,N_9978);
nor UO_586 (O_586,N_9555,N_9870);
and UO_587 (O_587,N_9062,N_9469);
and UO_588 (O_588,N_9860,N_9479);
nor UO_589 (O_589,N_9414,N_9555);
nor UO_590 (O_590,N_9368,N_9313);
or UO_591 (O_591,N_9219,N_9510);
and UO_592 (O_592,N_9218,N_9614);
and UO_593 (O_593,N_9530,N_9111);
nand UO_594 (O_594,N_9529,N_9931);
nor UO_595 (O_595,N_9383,N_9261);
and UO_596 (O_596,N_9465,N_9061);
or UO_597 (O_597,N_9547,N_9026);
nand UO_598 (O_598,N_9483,N_9197);
nor UO_599 (O_599,N_9879,N_9566);
or UO_600 (O_600,N_9372,N_9555);
and UO_601 (O_601,N_9024,N_9416);
nand UO_602 (O_602,N_9972,N_9499);
nand UO_603 (O_603,N_9057,N_9917);
and UO_604 (O_604,N_9843,N_9486);
or UO_605 (O_605,N_9721,N_9946);
nand UO_606 (O_606,N_9354,N_9568);
or UO_607 (O_607,N_9062,N_9051);
or UO_608 (O_608,N_9140,N_9707);
nor UO_609 (O_609,N_9907,N_9377);
nand UO_610 (O_610,N_9727,N_9226);
nor UO_611 (O_611,N_9035,N_9762);
nor UO_612 (O_612,N_9273,N_9405);
and UO_613 (O_613,N_9356,N_9697);
nor UO_614 (O_614,N_9793,N_9133);
nand UO_615 (O_615,N_9488,N_9683);
or UO_616 (O_616,N_9574,N_9028);
nand UO_617 (O_617,N_9319,N_9985);
nor UO_618 (O_618,N_9539,N_9341);
and UO_619 (O_619,N_9683,N_9068);
nor UO_620 (O_620,N_9355,N_9574);
nor UO_621 (O_621,N_9131,N_9544);
and UO_622 (O_622,N_9067,N_9465);
or UO_623 (O_623,N_9063,N_9064);
and UO_624 (O_624,N_9117,N_9182);
or UO_625 (O_625,N_9142,N_9395);
nand UO_626 (O_626,N_9371,N_9486);
or UO_627 (O_627,N_9115,N_9199);
and UO_628 (O_628,N_9784,N_9603);
nand UO_629 (O_629,N_9720,N_9942);
nor UO_630 (O_630,N_9157,N_9509);
or UO_631 (O_631,N_9725,N_9018);
nand UO_632 (O_632,N_9974,N_9723);
nor UO_633 (O_633,N_9992,N_9884);
and UO_634 (O_634,N_9604,N_9114);
or UO_635 (O_635,N_9160,N_9568);
nor UO_636 (O_636,N_9767,N_9573);
nand UO_637 (O_637,N_9938,N_9714);
and UO_638 (O_638,N_9537,N_9577);
or UO_639 (O_639,N_9686,N_9323);
nor UO_640 (O_640,N_9178,N_9676);
nand UO_641 (O_641,N_9996,N_9036);
or UO_642 (O_642,N_9663,N_9017);
or UO_643 (O_643,N_9581,N_9799);
nor UO_644 (O_644,N_9118,N_9732);
and UO_645 (O_645,N_9674,N_9962);
nor UO_646 (O_646,N_9897,N_9154);
or UO_647 (O_647,N_9141,N_9876);
nor UO_648 (O_648,N_9934,N_9609);
or UO_649 (O_649,N_9422,N_9269);
nor UO_650 (O_650,N_9539,N_9853);
or UO_651 (O_651,N_9501,N_9634);
nor UO_652 (O_652,N_9410,N_9396);
and UO_653 (O_653,N_9244,N_9725);
or UO_654 (O_654,N_9797,N_9334);
and UO_655 (O_655,N_9252,N_9020);
or UO_656 (O_656,N_9091,N_9173);
or UO_657 (O_657,N_9825,N_9655);
or UO_658 (O_658,N_9327,N_9362);
or UO_659 (O_659,N_9183,N_9039);
and UO_660 (O_660,N_9070,N_9364);
or UO_661 (O_661,N_9780,N_9242);
nand UO_662 (O_662,N_9851,N_9540);
and UO_663 (O_663,N_9856,N_9139);
nor UO_664 (O_664,N_9110,N_9155);
nand UO_665 (O_665,N_9161,N_9472);
nor UO_666 (O_666,N_9783,N_9222);
and UO_667 (O_667,N_9924,N_9724);
or UO_668 (O_668,N_9112,N_9736);
nand UO_669 (O_669,N_9338,N_9540);
and UO_670 (O_670,N_9857,N_9617);
nor UO_671 (O_671,N_9614,N_9499);
or UO_672 (O_672,N_9201,N_9293);
or UO_673 (O_673,N_9220,N_9753);
nor UO_674 (O_674,N_9571,N_9401);
nand UO_675 (O_675,N_9297,N_9966);
and UO_676 (O_676,N_9956,N_9015);
and UO_677 (O_677,N_9638,N_9003);
nor UO_678 (O_678,N_9158,N_9389);
or UO_679 (O_679,N_9957,N_9083);
and UO_680 (O_680,N_9816,N_9882);
or UO_681 (O_681,N_9001,N_9781);
nand UO_682 (O_682,N_9157,N_9135);
nand UO_683 (O_683,N_9110,N_9389);
nand UO_684 (O_684,N_9211,N_9552);
nor UO_685 (O_685,N_9605,N_9873);
and UO_686 (O_686,N_9282,N_9850);
nand UO_687 (O_687,N_9884,N_9231);
nor UO_688 (O_688,N_9988,N_9698);
nor UO_689 (O_689,N_9410,N_9998);
xnor UO_690 (O_690,N_9657,N_9485);
nor UO_691 (O_691,N_9609,N_9268);
nand UO_692 (O_692,N_9747,N_9473);
nand UO_693 (O_693,N_9333,N_9962);
and UO_694 (O_694,N_9605,N_9080);
or UO_695 (O_695,N_9026,N_9822);
nor UO_696 (O_696,N_9751,N_9121);
or UO_697 (O_697,N_9457,N_9617);
or UO_698 (O_698,N_9256,N_9762);
and UO_699 (O_699,N_9914,N_9698);
or UO_700 (O_700,N_9422,N_9301);
or UO_701 (O_701,N_9901,N_9932);
or UO_702 (O_702,N_9759,N_9896);
and UO_703 (O_703,N_9066,N_9945);
and UO_704 (O_704,N_9809,N_9246);
nand UO_705 (O_705,N_9022,N_9238);
and UO_706 (O_706,N_9592,N_9441);
nand UO_707 (O_707,N_9276,N_9918);
or UO_708 (O_708,N_9628,N_9555);
nor UO_709 (O_709,N_9162,N_9686);
nor UO_710 (O_710,N_9465,N_9994);
nand UO_711 (O_711,N_9600,N_9485);
nand UO_712 (O_712,N_9429,N_9878);
nor UO_713 (O_713,N_9710,N_9744);
or UO_714 (O_714,N_9592,N_9867);
nor UO_715 (O_715,N_9559,N_9501);
and UO_716 (O_716,N_9965,N_9044);
or UO_717 (O_717,N_9965,N_9630);
nand UO_718 (O_718,N_9365,N_9041);
nor UO_719 (O_719,N_9004,N_9572);
or UO_720 (O_720,N_9000,N_9727);
and UO_721 (O_721,N_9141,N_9765);
or UO_722 (O_722,N_9133,N_9049);
nand UO_723 (O_723,N_9642,N_9985);
and UO_724 (O_724,N_9375,N_9785);
nand UO_725 (O_725,N_9703,N_9373);
and UO_726 (O_726,N_9753,N_9476);
nor UO_727 (O_727,N_9180,N_9327);
nand UO_728 (O_728,N_9127,N_9543);
nand UO_729 (O_729,N_9686,N_9361);
nand UO_730 (O_730,N_9050,N_9666);
and UO_731 (O_731,N_9382,N_9716);
and UO_732 (O_732,N_9466,N_9124);
and UO_733 (O_733,N_9724,N_9903);
and UO_734 (O_734,N_9483,N_9282);
and UO_735 (O_735,N_9832,N_9180);
and UO_736 (O_736,N_9399,N_9117);
or UO_737 (O_737,N_9917,N_9496);
and UO_738 (O_738,N_9707,N_9329);
nand UO_739 (O_739,N_9493,N_9045);
and UO_740 (O_740,N_9018,N_9278);
and UO_741 (O_741,N_9155,N_9703);
and UO_742 (O_742,N_9462,N_9849);
nand UO_743 (O_743,N_9869,N_9212);
nand UO_744 (O_744,N_9124,N_9251);
nand UO_745 (O_745,N_9257,N_9659);
and UO_746 (O_746,N_9192,N_9581);
and UO_747 (O_747,N_9971,N_9249);
nor UO_748 (O_748,N_9559,N_9894);
nand UO_749 (O_749,N_9798,N_9252);
nand UO_750 (O_750,N_9138,N_9074);
or UO_751 (O_751,N_9570,N_9955);
or UO_752 (O_752,N_9444,N_9675);
and UO_753 (O_753,N_9890,N_9510);
and UO_754 (O_754,N_9540,N_9943);
nor UO_755 (O_755,N_9761,N_9110);
or UO_756 (O_756,N_9458,N_9213);
or UO_757 (O_757,N_9631,N_9301);
nand UO_758 (O_758,N_9219,N_9469);
nor UO_759 (O_759,N_9005,N_9333);
and UO_760 (O_760,N_9719,N_9654);
nand UO_761 (O_761,N_9820,N_9710);
and UO_762 (O_762,N_9417,N_9944);
nor UO_763 (O_763,N_9913,N_9002);
nor UO_764 (O_764,N_9026,N_9041);
nor UO_765 (O_765,N_9064,N_9398);
and UO_766 (O_766,N_9537,N_9134);
or UO_767 (O_767,N_9118,N_9134);
and UO_768 (O_768,N_9450,N_9947);
nor UO_769 (O_769,N_9372,N_9128);
nand UO_770 (O_770,N_9727,N_9067);
nor UO_771 (O_771,N_9957,N_9107);
nand UO_772 (O_772,N_9746,N_9286);
and UO_773 (O_773,N_9246,N_9872);
and UO_774 (O_774,N_9692,N_9225);
and UO_775 (O_775,N_9261,N_9985);
or UO_776 (O_776,N_9814,N_9258);
nand UO_777 (O_777,N_9921,N_9922);
or UO_778 (O_778,N_9154,N_9026);
or UO_779 (O_779,N_9992,N_9325);
or UO_780 (O_780,N_9119,N_9766);
or UO_781 (O_781,N_9585,N_9814);
nor UO_782 (O_782,N_9445,N_9438);
nor UO_783 (O_783,N_9145,N_9115);
or UO_784 (O_784,N_9750,N_9299);
nor UO_785 (O_785,N_9109,N_9088);
and UO_786 (O_786,N_9850,N_9720);
and UO_787 (O_787,N_9350,N_9469);
and UO_788 (O_788,N_9334,N_9021);
and UO_789 (O_789,N_9383,N_9555);
and UO_790 (O_790,N_9482,N_9087);
nor UO_791 (O_791,N_9035,N_9308);
nand UO_792 (O_792,N_9566,N_9915);
nand UO_793 (O_793,N_9678,N_9688);
nor UO_794 (O_794,N_9454,N_9879);
nor UO_795 (O_795,N_9830,N_9275);
and UO_796 (O_796,N_9413,N_9400);
nand UO_797 (O_797,N_9944,N_9605);
nand UO_798 (O_798,N_9519,N_9850);
or UO_799 (O_799,N_9532,N_9731);
nor UO_800 (O_800,N_9936,N_9992);
and UO_801 (O_801,N_9720,N_9710);
nor UO_802 (O_802,N_9647,N_9908);
or UO_803 (O_803,N_9794,N_9290);
nand UO_804 (O_804,N_9262,N_9971);
nand UO_805 (O_805,N_9889,N_9640);
or UO_806 (O_806,N_9761,N_9213);
nand UO_807 (O_807,N_9945,N_9001);
nand UO_808 (O_808,N_9433,N_9309);
nand UO_809 (O_809,N_9726,N_9787);
or UO_810 (O_810,N_9706,N_9489);
nor UO_811 (O_811,N_9754,N_9018);
nor UO_812 (O_812,N_9703,N_9180);
and UO_813 (O_813,N_9951,N_9888);
and UO_814 (O_814,N_9454,N_9826);
or UO_815 (O_815,N_9997,N_9934);
and UO_816 (O_816,N_9203,N_9184);
xor UO_817 (O_817,N_9337,N_9440);
and UO_818 (O_818,N_9813,N_9624);
and UO_819 (O_819,N_9680,N_9172);
nand UO_820 (O_820,N_9802,N_9156);
and UO_821 (O_821,N_9946,N_9211);
and UO_822 (O_822,N_9045,N_9569);
or UO_823 (O_823,N_9527,N_9941);
nor UO_824 (O_824,N_9347,N_9546);
nand UO_825 (O_825,N_9432,N_9180);
or UO_826 (O_826,N_9786,N_9403);
and UO_827 (O_827,N_9489,N_9244);
nand UO_828 (O_828,N_9583,N_9614);
nand UO_829 (O_829,N_9936,N_9105);
nor UO_830 (O_830,N_9190,N_9848);
nor UO_831 (O_831,N_9324,N_9878);
and UO_832 (O_832,N_9664,N_9444);
or UO_833 (O_833,N_9589,N_9923);
nor UO_834 (O_834,N_9942,N_9658);
and UO_835 (O_835,N_9604,N_9814);
nand UO_836 (O_836,N_9418,N_9970);
and UO_837 (O_837,N_9529,N_9564);
or UO_838 (O_838,N_9563,N_9786);
nand UO_839 (O_839,N_9810,N_9282);
and UO_840 (O_840,N_9810,N_9539);
or UO_841 (O_841,N_9529,N_9286);
nor UO_842 (O_842,N_9302,N_9934);
nand UO_843 (O_843,N_9804,N_9853);
nand UO_844 (O_844,N_9688,N_9079);
nor UO_845 (O_845,N_9336,N_9473);
and UO_846 (O_846,N_9535,N_9056);
or UO_847 (O_847,N_9901,N_9029);
nand UO_848 (O_848,N_9837,N_9210);
nor UO_849 (O_849,N_9640,N_9451);
or UO_850 (O_850,N_9436,N_9947);
nand UO_851 (O_851,N_9492,N_9640);
and UO_852 (O_852,N_9460,N_9048);
and UO_853 (O_853,N_9576,N_9328);
nor UO_854 (O_854,N_9235,N_9587);
or UO_855 (O_855,N_9183,N_9237);
and UO_856 (O_856,N_9901,N_9299);
nand UO_857 (O_857,N_9154,N_9051);
xor UO_858 (O_858,N_9552,N_9093);
nor UO_859 (O_859,N_9856,N_9897);
nor UO_860 (O_860,N_9166,N_9654);
and UO_861 (O_861,N_9471,N_9783);
and UO_862 (O_862,N_9878,N_9203);
nor UO_863 (O_863,N_9177,N_9136);
nor UO_864 (O_864,N_9602,N_9050);
nor UO_865 (O_865,N_9535,N_9334);
nand UO_866 (O_866,N_9346,N_9067);
nor UO_867 (O_867,N_9234,N_9700);
or UO_868 (O_868,N_9718,N_9599);
nor UO_869 (O_869,N_9398,N_9469);
or UO_870 (O_870,N_9796,N_9341);
xor UO_871 (O_871,N_9271,N_9141);
nand UO_872 (O_872,N_9559,N_9592);
nor UO_873 (O_873,N_9860,N_9521);
or UO_874 (O_874,N_9348,N_9350);
nand UO_875 (O_875,N_9418,N_9346);
nand UO_876 (O_876,N_9899,N_9864);
and UO_877 (O_877,N_9728,N_9415);
or UO_878 (O_878,N_9037,N_9967);
nor UO_879 (O_879,N_9494,N_9388);
and UO_880 (O_880,N_9460,N_9895);
nor UO_881 (O_881,N_9015,N_9239);
nor UO_882 (O_882,N_9819,N_9506);
nor UO_883 (O_883,N_9876,N_9507);
nor UO_884 (O_884,N_9183,N_9016);
nor UO_885 (O_885,N_9886,N_9088);
nor UO_886 (O_886,N_9934,N_9961);
nor UO_887 (O_887,N_9886,N_9488);
and UO_888 (O_888,N_9002,N_9146);
and UO_889 (O_889,N_9925,N_9030);
nor UO_890 (O_890,N_9776,N_9477);
and UO_891 (O_891,N_9134,N_9226);
nor UO_892 (O_892,N_9715,N_9990);
or UO_893 (O_893,N_9684,N_9037);
nand UO_894 (O_894,N_9151,N_9208);
or UO_895 (O_895,N_9744,N_9048);
or UO_896 (O_896,N_9627,N_9244);
and UO_897 (O_897,N_9586,N_9215);
nor UO_898 (O_898,N_9008,N_9355);
or UO_899 (O_899,N_9164,N_9682);
or UO_900 (O_900,N_9699,N_9599);
and UO_901 (O_901,N_9292,N_9631);
nand UO_902 (O_902,N_9292,N_9217);
and UO_903 (O_903,N_9877,N_9770);
nand UO_904 (O_904,N_9158,N_9064);
and UO_905 (O_905,N_9192,N_9800);
nand UO_906 (O_906,N_9742,N_9716);
or UO_907 (O_907,N_9537,N_9755);
and UO_908 (O_908,N_9790,N_9725);
and UO_909 (O_909,N_9806,N_9820);
nand UO_910 (O_910,N_9895,N_9767);
nand UO_911 (O_911,N_9615,N_9822);
or UO_912 (O_912,N_9400,N_9785);
nor UO_913 (O_913,N_9076,N_9382);
or UO_914 (O_914,N_9178,N_9119);
or UO_915 (O_915,N_9626,N_9129);
nor UO_916 (O_916,N_9891,N_9733);
or UO_917 (O_917,N_9738,N_9986);
nor UO_918 (O_918,N_9408,N_9384);
nand UO_919 (O_919,N_9344,N_9608);
nor UO_920 (O_920,N_9817,N_9833);
and UO_921 (O_921,N_9047,N_9257);
and UO_922 (O_922,N_9959,N_9395);
nand UO_923 (O_923,N_9919,N_9545);
nor UO_924 (O_924,N_9832,N_9288);
nand UO_925 (O_925,N_9953,N_9115);
nor UO_926 (O_926,N_9596,N_9337);
nor UO_927 (O_927,N_9584,N_9224);
and UO_928 (O_928,N_9421,N_9143);
nand UO_929 (O_929,N_9042,N_9362);
nor UO_930 (O_930,N_9397,N_9355);
nor UO_931 (O_931,N_9802,N_9928);
nor UO_932 (O_932,N_9914,N_9272);
and UO_933 (O_933,N_9412,N_9365);
nand UO_934 (O_934,N_9463,N_9833);
nand UO_935 (O_935,N_9983,N_9701);
or UO_936 (O_936,N_9566,N_9217);
nand UO_937 (O_937,N_9340,N_9149);
and UO_938 (O_938,N_9359,N_9607);
and UO_939 (O_939,N_9069,N_9434);
nand UO_940 (O_940,N_9470,N_9564);
nand UO_941 (O_941,N_9707,N_9625);
nor UO_942 (O_942,N_9932,N_9191);
and UO_943 (O_943,N_9574,N_9222);
or UO_944 (O_944,N_9143,N_9445);
nor UO_945 (O_945,N_9402,N_9467);
and UO_946 (O_946,N_9584,N_9578);
nand UO_947 (O_947,N_9581,N_9514);
nand UO_948 (O_948,N_9536,N_9366);
nand UO_949 (O_949,N_9933,N_9067);
and UO_950 (O_950,N_9386,N_9097);
and UO_951 (O_951,N_9914,N_9986);
and UO_952 (O_952,N_9170,N_9341);
or UO_953 (O_953,N_9131,N_9527);
or UO_954 (O_954,N_9589,N_9470);
nor UO_955 (O_955,N_9797,N_9698);
nand UO_956 (O_956,N_9358,N_9053);
nor UO_957 (O_957,N_9037,N_9695);
nand UO_958 (O_958,N_9347,N_9363);
and UO_959 (O_959,N_9351,N_9560);
and UO_960 (O_960,N_9872,N_9172);
or UO_961 (O_961,N_9954,N_9297);
or UO_962 (O_962,N_9088,N_9611);
nand UO_963 (O_963,N_9163,N_9562);
or UO_964 (O_964,N_9323,N_9755);
nor UO_965 (O_965,N_9595,N_9926);
or UO_966 (O_966,N_9889,N_9877);
and UO_967 (O_967,N_9142,N_9234);
nor UO_968 (O_968,N_9856,N_9586);
nand UO_969 (O_969,N_9535,N_9512);
nor UO_970 (O_970,N_9729,N_9422);
nand UO_971 (O_971,N_9278,N_9787);
nor UO_972 (O_972,N_9842,N_9369);
or UO_973 (O_973,N_9345,N_9150);
or UO_974 (O_974,N_9223,N_9088);
or UO_975 (O_975,N_9281,N_9295);
or UO_976 (O_976,N_9495,N_9442);
nand UO_977 (O_977,N_9628,N_9925);
nand UO_978 (O_978,N_9314,N_9278);
nand UO_979 (O_979,N_9971,N_9412);
xor UO_980 (O_980,N_9821,N_9502);
or UO_981 (O_981,N_9118,N_9573);
or UO_982 (O_982,N_9723,N_9864);
nand UO_983 (O_983,N_9580,N_9806);
nor UO_984 (O_984,N_9979,N_9351);
nand UO_985 (O_985,N_9819,N_9525);
nor UO_986 (O_986,N_9648,N_9236);
or UO_987 (O_987,N_9145,N_9060);
nand UO_988 (O_988,N_9587,N_9082);
or UO_989 (O_989,N_9097,N_9392);
and UO_990 (O_990,N_9735,N_9447);
nor UO_991 (O_991,N_9235,N_9278);
and UO_992 (O_992,N_9317,N_9712);
nand UO_993 (O_993,N_9458,N_9025);
nand UO_994 (O_994,N_9655,N_9802);
nand UO_995 (O_995,N_9636,N_9988);
nand UO_996 (O_996,N_9828,N_9181);
and UO_997 (O_997,N_9493,N_9352);
or UO_998 (O_998,N_9204,N_9257);
xnor UO_999 (O_999,N_9792,N_9910);
nand UO_1000 (O_1000,N_9906,N_9386);
and UO_1001 (O_1001,N_9624,N_9777);
nor UO_1002 (O_1002,N_9329,N_9062);
nand UO_1003 (O_1003,N_9565,N_9524);
nand UO_1004 (O_1004,N_9026,N_9759);
nor UO_1005 (O_1005,N_9806,N_9267);
nand UO_1006 (O_1006,N_9613,N_9569);
nor UO_1007 (O_1007,N_9443,N_9597);
or UO_1008 (O_1008,N_9365,N_9880);
nand UO_1009 (O_1009,N_9157,N_9909);
or UO_1010 (O_1010,N_9594,N_9992);
and UO_1011 (O_1011,N_9666,N_9342);
and UO_1012 (O_1012,N_9564,N_9694);
or UO_1013 (O_1013,N_9262,N_9310);
xor UO_1014 (O_1014,N_9037,N_9060);
nor UO_1015 (O_1015,N_9165,N_9163);
and UO_1016 (O_1016,N_9915,N_9251);
and UO_1017 (O_1017,N_9275,N_9638);
or UO_1018 (O_1018,N_9173,N_9703);
nor UO_1019 (O_1019,N_9688,N_9990);
nor UO_1020 (O_1020,N_9540,N_9111);
and UO_1021 (O_1021,N_9708,N_9396);
nand UO_1022 (O_1022,N_9664,N_9202);
nand UO_1023 (O_1023,N_9183,N_9262);
and UO_1024 (O_1024,N_9645,N_9728);
nand UO_1025 (O_1025,N_9624,N_9797);
nor UO_1026 (O_1026,N_9497,N_9690);
or UO_1027 (O_1027,N_9260,N_9403);
nor UO_1028 (O_1028,N_9342,N_9477);
nor UO_1029 (O_1029,N_9098,N_9491);
and UO_1030 (O_1030,N_9841,N_9479);
nor UO_1031 (O_1031,N_9748,N_9432);
and UO_1032 (O_1032,N_9973,N_9518);
nand UO_1033 (O_1033,N_9962,N_9057);
or UO_1034 (O_1034,N_9513,N_9798);
nand UO_1035 (O_1035,N_9500,N_9909);
nor UO_1036 (O_1036,N_9638,N_9049);
xor UO_1037 (O_1037,N_9194,N_9064);
nor UO_1038 (O_1038,N_9617,N_9932);
nand UO_1039 (O_1039,N_9579,N_9555);
nor UO_1040 (O_1040,N_9862,N_9430);
nand UO_1041 (O_1041,N_9725,N_9268);
and UO_1042 (O_1042,N_9600,N_9769);
nor UO_1043 (O_1043,N_9204,N_9463);
or UO_1044 (O_1044,N_9022,N_9145);
or UO_1045 (O_1045,N_9763,N_9197);
or UO_1046 (O_1046,N_9816,N_9654);
and UO_1047 (O_1047,N_9499,N_9096);
nand UO_1048 (O_1048,N_9426,N_9217);
nor UO_1049 (O_1049,N_9715,N_9493);
nand UO_1050 (O_1050,N_9218,N_9123);
nand UO_1051 (O_1051,N_9456,N_9797);
and UO_1052 (O_1052,N_9926,N_9359);
nor UO_1053 (O_1053,N_9994,N_9008);
or UO_1054 (O_1054,N_9729,N_9718);
or UO_1055 (O_1055,N_9514,N_9609);
or UO_1056 (O_1056,N_9448,N_9379);
and UO_1057 (O_1057,N_9459,N_9861);
or UO_1058 (O_1058,N_9647,N_9058);
and UO_1059 (O_1059,N_9363,N_9501);
nand UO_1060 (O_1060,N_9087,N_9092);
and UO_1061 (O_1061,N_9175,N_9511);
or UO_1062 (O_1062,N_9837,N_9963);
nor UO_1063 (O_1063,N_9296,N_9583);
nor UO_1064 (O_1064,N_9576,N_9375);
and UO_1065 (O_1065,N_9372,N_9422);
nand UO_1066 (O_1066,N_9782,N_9780);
nand UO_1067 (O_1067,N_9558,N_9208);
nand UO_1068 (O_1068,N_9333,N_9446);
nor UO_1069 (O_1069,N_9522,N_9498);
nor UO_1070 (O_1070,N_9668,N_9025);
or UO_1071 (O_1071,N_9633,N_9140);
or UO_1072 (O_1072,N_9225,N_9822);
and UO_1073 (O_1073,N_9676,N_9920);
nand UO_1074 (O_1074,N_9066,N_9473);
or UO_1075 (O_1075,N_9355,N_9671);
or UO_1076 (O_1076,N_9279,N_9526);
or UO_1077 (O_1077,N_9567,N_9261);
or UO_1078 (O_1078,N_9996,N_9883);
nand UO_1079 (O_1079,N_9899,N_9314);
and UO_1080 (O_1080,N_9042,N_9753);
or UO_1081 (O_1081,N_9651,N_9915);
nand UO_1082 (O_1082,N_9519,N_9548);
nand UO_1083 (O_1083,N_9521,N_9732);
and UO_1084 (O_1084,N_9057,N_9406);
nor UO_1085 (O_1085,N_9481,N_9747);
or UO_1086 (O_1086,N_9343,N_9989);
nand UO_1087 (O_1087,N_9148,N_9360);
nor UO_1088 (O_1088,N_9406,N_9630);
or UO_1089 (O_1089,N_9113,N_9597);
or UO_1090 (O_1090,N_9620,N_9176);
or UO_1091 (O_1091,N_9600,N_9890);
nand UO_1092 (O_1092,N_9018,N_9374);
and UO_1093 (O_1093,N_9464,N_9968);
or UO_1094 (O_1094,N_9736,N_9244);
nand UO_1095 (O_1095,N_9245,N_9667);
or UO_1096 (O_1096,N_9290,N_9180);
or UO_1097 (O_1097,N_9065,N_9343);
or UO_1098 (O_1098,N_9873,N_9122);
and UO_1099 (O_1099,N_9191,N_9904);
or UO_1100 (O_1100,N_9669,N_9580);
and UO_1101 (O_1101,N_9702,N_9541);
and UO_1102 (O_1102,N_9422,N_9621);
nand UO_1103 (O_1103,N_9630,N_9016);
or UO_1104 (O_1104,N_9274,N_9364);
nor UO_1105 (O_1105,N_9392,N_9349);
or UO_1106 (O_1106,N_9009,N_9991);
or UO_1107 (O_1107,N_9403,N_9869);
nand UO_1108 (O_1108,N_9106,N_9702);
nor UO_1109 (O_1109,N_9870,N_9007);
and UO_1110 (O_1110,N_9089,N_9939);
nor UO_1111 (O_1111,N_9226,N_9123);
nand UO_1112 (O_1112,N_9894,N_9032);
or UO_1113 (O_1113,N_9572,N_9664);
nand UO_1114 (O_1114,N_9043,N_9544);
nor UO_1115 (O_1115,N_9808,N_9451);
nor UO_1116 (O_1116,N_9998,N_9337);
nand UO_1117 (O_1117,N_9081,N_9729);
and UO_1118 (O_1118,N_9243,N_9771);
and UO_1119 (O_1119,N_9836,N_9192);
nand UO_1120 (O_1120,N_9464,N_9513);
nor UO_1121 (O_1121,N_9484,N_9850);
or UO_1122 (O_1122,N_9887,N_9643);
and UO_1123 (O_1123,N_9256,N_9122);
or UO_1124 (O_1124,N_9001,N_9247);
and UO_1125 (O_1125,N_9009,N_9136);
nor UO_1126 (O_1126,N_9966,N_9221);
nand UO_1127 (O_1127,N_9626,N_9034);
or UO_1128 (O_1128,N_9919,N_9474);
nand UO_1129 (O_1129,N_9616,N_9984);
or UO_1130 (O_1130,N_9064,N_9866);
or UO_1131 (O_1131,N_9892,N_9360);
nand UO_1132 (O_1132,N_9627,N_9319);
or UO_1133 (O_1133,N_9733,N_9630);
nand UO_1134 (O_1134,N_9940,N_9361);
nor UO_1135 (O_1135,N_9992,N_9663);
or UO_1136 (O_1136,N_9831,N_9860);
and UO_1137 (O_1137,N_9051,N_9001);
nand UO_1138 (O_1138,N_9715,N_9251);
nor UO_1139 (O_1139,N_9453,N_9633);
nor UO_1140 (O_1140,N_9153,N_9846);
nor UO_1141 (O_1141,N_9801,N_9516);
or UO_1142 (O_1142,N_9324,N_9801);
nand UO_1143 (O_1143,N_9428,N_9811);
nor UO_1144 (O_1144,N_9856,N_9216);
nand UO_1145 (O_1145,N_9916,N_9215);
nor UO_1146 (O_1146,N_9061,N_9797);
nor UO_1147 (O_1147,N_9374,N_9781);
nor UO_1148 (O_1148,N_9903,N_9747);
and UO_1149 (O_1149,N_9573,N_9804);
nand UO_1150 (O_1150,N_9959,N_9549);
nand UO_1151 (O_1151,N_9423,N_9253);
nand UO_1152 (O_1152,N_9204,N_9472);
nand UO_1153 (O_1153,N_9862,N_9616);
nor UO_1154 (O_1154,N_9185,N_9371);
and UO_1155 (O_1155,N_9954,N_9331);
and UO_1156 (O_1156,N_9317,N_9073);
nand UO_1157 (O_1157,N_9890,N_9130);
and UO_1158 (O_1158,N_9159,N_9851);
nand UO_1159 (O_1159,N_9351,N_9840);
xnor UO_1160 (O_1160,N_9347,N_9857);
nor UO_1161 (O_1161,N_9030,N_9815);
nor UO_1162 (O_1162,N_9928,N_9036);
or UO_1163 (O_1163,N_9996,N_9756);
nor UO_1164 (O_1164,N_9965,N_9257);
nor UO_1165 (O_1165,N_9472,N_9934);
and UO_1166 (O_1166,N_9537,N_9258);
and UO_1167 (O_1167,N_9946,N_9428);
and UO_1168 (O_1168,N_9951,N_9583);
and UO_1169 (O_1169,N_9897,N_9691);
and UO_1170 (O_1170,N_9261,N_9725);
and UO_1171 (O_1171,N_9107,N_9520);
nand UO_1172 (O_1172,N_9690,N_9855);
or UO_1173 (O_1173,N_9738,N_9507);
or UO_1174 (O_1174,N_9781,N_9630);
and UO_1175 (O_1175,N_9994,N_9746);
or UO_1176 (O_1176,N_9139,N_9601);
nor UO_1177 (O_1177,N_9895,N_9755);
nor UO_1178 (O_1178,N_9289,N_9438);
nor UO_1179 (O_1179,N_9085,N_9043);
and UO_1180 (O_1180,N_9695,N_9608);
and UO_1181 (O_1181,N_9250,N_9011);
nand UO_1182 (O_1182,N_9488,N_9769);
nor UO_1183 (O_1183,N_9830,N_9187);
nor UO_1184 (O_1184,N_9187,N_9881);
and UO_1185 (O_1185,N_9611,N_9899);
nand UO_1186 (O_1186,N_9130,N_9083);
and UO_1187 (O_1187,N_9455,N_9443);
nor UO_1188 (O_1188,N_9666,N_9091);
or UO_1189 (O_1189,N_9657,N_9001);
nor UO_1190 (O_1190,N_9874,N_9243);
and UO_1191 (O_1191,N_9663,N_9551);
or UO_1192 (O_1192,N_9888,N_9454);
and UO_1193 (O_1193,N_9932,N_9335);
or UO_1194 (O_1194,N_9412,N_9189);
nor UO_1195 (O_1195,N_9711,N_9089);
nand UO_1196 (O_1196,N_9564,N_9020);
nand UO_1197 (O_1197,N_9725,N_9559);
and UO_1198 (O_1198,N_9197,N_9745);
and UO_1199 (O_1199,N_9575,N_9012);
or UO_1200 (O_1200,N_9409,N_9865);
and UO_1201 (O_1201,N_9198,N_9348);
nor UO_1202 (O_1202,N_9372,N_9468);
nand UO_1203 (O_1203,N_9075,N_9590);
nand UO_1204 (O_1204,N_9241,N_9524);
nand UO_1205 (O_1205,N_9810,N_9252);
nand UO_1206 (O_1206,N_9506,N_9584);
nand UO_1207 (O_1207,N_9500,N_9511);
nor UO_1208 (O_1208,N_9242,N_9900);
or UO_1209 (O_1209,N_9109,N_9257);
nor UO_1210 (O_1210,N_9881,N_9821);
nor UO_1211 (O_1211,N_9529,N_9853);
or UO_1212 (O_1212,N_9238,N_9442);
nor UO_1213 (O_1213,N_9107,N_9622);
nor UO_1214 (O_1214,N_9854,N_9267);
and UO_1215 (O_1215,N_9957,N_9016);
or UO_1216 (O_1216,N_9719,N_9847);
or UO_1217 (O_1217,N_9524,N_9080);
and UO_1218 (O_1218,N_9950,N_9429);
and UO_1219 (O_1219,N_9705,N_9361);
and UO_1220 (O_1220,N_9829,N_9406);
nand UO_1221 (O_1221,N_9420,N_9324);
nand UO_1222 (O_1222,N_9471,N_9001);
and UO_1223 (O_1223,N_9492,N_9324);
and UO_1224 (O_1224,N_9056,N_9420);
nand UO_1225 (O_1225,N_9080,N_9958);
nor UO_1226 (O_1226,N_9107,N_9800);
nand UO_1227 (O_1227,N_9027,N_9544);
nand UO_1228 (O_1228,N_9976,N_9605);
or UO_1229 (O_1229,N_9263,N_9690);
nand UO_1230 (O_1230,N_9224,N_9624);
and UO_1231 (O_1231,N_9553,N_9929);
or UO_1232 (O_1232,N_9361,N_9202);
or UO_1233 (O_1233,N_9861,N_9270);
or UO_1234 (O_1234,N_9670,N_9188);
nor UO_1235 (O_1235,N_9836,N_9601);
nand UO_1236 (O_1236,N_9841,N_9787);
nor UO_1237 (O_1237,N_9494,N_9427);
nand UO_1238 (O_1238,N_9076,N_9868);
or UO_1239 (O_1239,N_9904,N_9995);
nand UO_1240 (O_1240,N_9309,N_9313);
or UO_1241 (O_1241,N_9434,N_9990);
xor UO_1242 (O_1242,N_9101,N_9012);
nand UO_1243 (O_1243,N_9476,N_9369);
nor UO_1244 (O_1244,N_9355,N_9704);
nand UO_1245 (O_1245,N_9369,N_9855);
and UO_1246 (O_1246,N_9045,N_9281);
or UO_1247 (O_1247,N_9916,N_9485);
and UO_1248 (O_1248,N_9392,N_9129);
nand UO_1249 (O_1249,N_9312,N_9294);
and UO_1250 (O_1250,N_9735,N_9047);
nor UO_1251 (O_1251,N_9978,N_9620);
xnor UO_1252 (O_1252,N_9922,N_9257);
nor UO_1253 (O_1253,N_9072,N_9777);
and UO_1254 (O_1254,N_9771,N_9097);
or UO_1255 (O_1255,N_9162,N_9726);
nand UO_1256 (O_1256,N_9879,N_9481);
nand UO_1257 (O_1257,N_9720,N_9798);
nor UO_1258 (O_1258,N_9044,N_9313);
nand UO_1259 (O_1259,N_9111,N_9719);
nor UO_1260 (O_1260,N_9097,N_9354);
or UO_1261 (O_1261,N_9334,N_9937);
or UO_1262 (O_1262,N_9545,N_9032);
and UO_1263 (O_1263,N_9567,N_9791);
and UO_1264 (O_1264,N_9453,N_9833);
or UO_1265 (O_1265,N_9997,N_9687);
or UO_1266 (O_1266,N_9047,N_9435);
and UO_1267 (O_1267,N_9214,N_9200);
nor UO_1268 (O_1268,N_9022,N_9283);
and UO_1269 (O_1269,N_9769,N_9971);
and UO_1270 (O_1270,N_9085,N_9432);
nand UO_1271 (O_1271,N_9580,N_9720);
nor UO_1272 (O_1272,N_9932,N_9759);
nor UO_1273 (O_1273,N_9360,N_9103);
and UO_1274 (O_1274,N_9654,N_9030);
nand UO_1275 (O_1275,N_9655,N_9320);
nand UO_1276 (O_1276,N_9242,N_9508);
nand UO_1277 (O_1277,N_9372,N_9548);
and UO_1278 (O_1278,N_9877,N_9984);
or UO_1279 (O_1279,N_9201,N_9409);
nor UO_1280 (O_1280,N_9349,N_9157);
and UO_1281 (O_1281,N_9719,N_9987);
or UO_1282 (O_1282,N_9253,N_9586);
or UO_1283 (O_1283,N_9946,N_9517);
or UO_1284 (O_1284,N_9382,N_9264);
and UO_1285 (O_1285,N_9406,N_9665);
nor UO_1286 (O_1286,N_9012,N_9877);
nor UO_1287 (O_1287,N_9168,N_9544);
nor UO_1288 (O_1288,N_9597,N_9173);
nor UO_1289 (O_1289,N_9415,N_9393);
nor UO_1290 (O_1290,N_9094,N_9992);
nor UO_1291 (O_1291,N_9102,N_9521);
and UO_1292 (O_1292,N_9711,N_9258);
nand UO_1293 (O_1293,N_9179,N_9816);
and UO_1294 (O_1294,N_9394,N_9810);
or UO_1295 (O_1295,N_9682,N_9568);
or UO_1296 (O_1296,N_9997,N_9972);
or UO_1297 (O_1297,N_9251,N_9798);
and UO_1298 (O_1298,N_9846,N_9346);
and UO_1299 (O_1299,N_9566,N_9206);
nand UO_1300 (O_1300,N_9971,N_9414);
or UO_1301 (O_1301,N_9460,N_9927);
and UO_1302 (O_1302,N_9763,N_9442);
nor UO_1303 (O_1303,N_9566,N_9603);
and UO_1304 (O_1304,N_9015,N_9816);
nor UO_1305 (O_1305,N_9726,N_9799);
and UO_1306 (O_1306,N_9045,N_9822);
nor UO_1307 (O_1307,N_9049,N_9027);
or UO_1308 (O_1308,N_9505,N_9973);
or UO_1309 (O_1309,N_9738,N_9319);
and UO_1310 (O_1310,N_9130,N_9385);
or UO_1311 (O_1311,N_9412,N_9613);
and UO_1312 (O_1312,N_9226,N_9794);
nor UO_1313 (O_1313,N_9955,N_9023);
nor UO_1314 (O_1314,N_9897,N_9281);
nor UO_1315 (O_1315,N_9366,N_9856);
nand UO_1316 (O_1316,N_9234,N_9139);
and UO_1317 (O_1317,N_9260,N_9409);
and UO_1318 (O_1318,N_9038,N_9307);
or UO_1319 (O_1319,N_9390,N_9461);
nand UO_1320 (O_1320,N_9047,N_9138);
or UO_1321 (O_1321,N_9279,N_9681);
and UO_1322 (O_1322,N_9023,N_9466);
or UO_1323 (O_1323,N_9965,N_9447);
nand UO_1324 (O_1324,N_9560,N_9203);
nor UO_1325 (O_1325,N_9933,N_9985);
xnor UO_1326 (O_1326,N_9804,N_9756);
nor UO_1327 (O_1327,N_9074,N_9294);
nor UO_1328 (O_1328,N_9970,N_9389);
nand UO_1329 (O_1329,N_9616,N_9376);
and UO_1330 (O_1330,N_9879,N_9615);
nor UO_1331 (O_1331,N_9196,N_9632);
and UO_1332 (O_1332,N_9175,N_9243);
nand UO_1333 (O_1333,N_9996,N_9021);
nor UO_1334 (O_1334,N_9294,N_9980);
or UO_1335 (O_1335,N_9793,N_9313);
nor UO_1336 (O_1336,N_9578,N_9028);
nor UO_1337 (O_1337,N_9192,N_9425);
and UO_1338 (O_1338,N_9508,N_9782);
or UO_1339 (O_1339,N_9795,N_9783);
and UO_1340 (O_1340,N_9042,N_9311);
or UO_1341 (O_1341,N_9869,N_9371);
and UO_1342 (O_1342,N_9998,N_9477);
nand UO_1343 (O_1343,N_9458,N_9800);
nor UO_1344 (O_1344,N_9816,N_9848);
nor UO_1345 (O_1345,N_9293,N_9340);
nand UO_1346 (O_1346,N_9487,N_9992);
nand UO_1347 (O_1347,N_9581,N_9540);
and UO_1348 (O_1348,N_9733,N_9126);
nor UO_1349 (O_1349,N_9055,N_9258);
or UO_1350 (O_1350,N_9879,N_9463);
or UO_1351 (O_1351,N_9563,N_9308);
and UO_1352 (O_1352,N_9914,N_9816);
nor UO_1353 (O_1353,N_9249,N_9307);
nand UO_1354 (O_1354,N_9056,N_9982);
and UO_1355 (O_1355,N_9178,N_9846);
nor UO_1356 (O_1356,N_9704,N_9353);
or UO_1357 (O_1357,N_9270,N_9433);
nand UO_1358 (O_1358,N_9265,N_9758);
or UO_1359 (O_1359,N_9832,N_9736);
and UO_1360 (O_1360,N_9983,N_9662);
and UO_1361 (O_1361,N_9882,N_9225);
nor UO_1362 (O_1362,N_9879,N_9128);
nor UO_1363 (O_1363,N_9404,N_9035);
nand UO_1364 (O_1364,N_9539,N_9014);
nor UO_1365 (O_1365,N_9110,N_9946);
nor UO_1366 (O_1366,N_9945,N_9297);
and UO_1367 (O_1367,N_9886,N_9244);
nor UO_1368 (O_1368,N_9506,N_9721);
or UO_1369 (O_1369,N_9671,N_9493);
and UO_1370 (O_1370,N_9548,N_9974);
nor UO_1371 (O_1371,N_9835,N_9288);
and UO_1372 (O_1372,N_9635,N_9350);
or UO_1373 (O_1373,N_9473,N_9407);
and UO_1374 (O_1374,N_9660,N_9698);
nor UO_1375 (O_1375,N_9086,N_9464);
nor UO_1376 (O_1376,N_9999,N_9351);
nand UO_1377 (O_1377,N_9713,N_9171);
nand UO_1378 (O_1378,N_9529,N_9490);
or UO_1379 (O_1379,N_9432,N_9214);
nand UO_1380 (O_1380,N_9295,N_9638);
nor UO_1381 (O_1381,N_9066,N_9745);
and UO_1382 (O_1382,N_9360,N_9093);
nor UO_1383 (O_1383,N_9789,N_9939);
and UO_1384 (O_1384,N_9155,N_9118);
nor UO_1385 (O_1385,N_9675,N_9229);
and UO_1386 (O_1386,N_9782,N_9838);
nand UO_1387 (O_1387,N_9292,N_9668);
or UO_1388 (O_1388,N_9102,N_9803);
or UO_1389 (O_1389,N_9984,N_9673);
nor UO_1390 (O_1390,N_9599,N_9908);
nand UO_1391 (O_1391,N_9425,N_9825);
nand UO_1392 (O_1392,N_9085,N_9684);
and UO_1393 (O_1393,N_9005,N_9027);
and UO_1394 (O_1394,N_9355,N_9550);
nand UO_1395 (O_1395,N_9049,N_9458);
nand UO_1396 (O_1396,N_9137,N_9992);
nor UO_1397 (O_1397,N_9151,N_9446);
nand UO_1398 (O_1398,N_9829,N_9317);
nor UO_1399 (O_1399,N_9929,N_9257);
or UO_1400 (O_1400,N_9150,N_9413);
and UO_1401 (O_1401,N_9697,N_9436);
nand UO_1402 (O_1402,N_9765,N_9245);
nor UO_1403 (O_1403,N_9229,N_9159);
nand UO_1404 (O_1404,N_9093,N_9428);
and UO_1405 (O_1405,N_9587,N_9346);
or UO_1406 (O_1406,N_9036,N_9706);
nand UO_1407 (O_1407,N_9826,N_9172);
and UO_1408 (O_1408,N_9970,N_9342);
or UO_1409 (O_1409,N_9656,N_9411);
and UO_1410 (O_1410,N_9562,N_9991);
nand UO_1411 (O_1411,N_9386,N_9484);
nand UO_1412 (O_1412,N_9365,N_9978);
nand UO_1413 (O_1413,N_9080,N_9269);
nand UO_1414 (O_1414,N_9800,N_9146);
nor UO_1415 (O_1415,N_9492,N_9853);
or UO_1416 (O_1416,N_9650,N_9593);
or UO_1417 (O_1417,N_9400,N_9182);
and UO_1418 (O_1418,N_9659,N_9809);
nor UO_1419 (O_1419,N_9451,N_9434);
or UO_1420 (O_1420,N_9346,N_9248);
xnor UO_1421 (O_1421,N_9256,N_9678);
and UO_1422 (O_1422,N_9502,N_9212);
and UO_1423 (O_1423,N_9103,N_9132);
or UO_1424 (O_1424,N_9057,N_9804);
nand UO_1425 (O_1425,N_9998,N_9937);
nor UO_1426 (O_1426,N_9625,N_9830);
nand UO_1427 (O_1427,N_9388,N_9058);
nor UO_1428 (O_1428,N_9336,N_9584);
and UO_1429 (O_1429,N_9864,N_9821);
nand UO_1430 (O_1430,N_9531,N_9893);
nand UO_1431 (O_1431,N_9735,N_9325);
nand UO_1432 (O_1432,N_9879,N_9813);
nand UO_1433 (O_1433,N_9773,N_9464);
nor UO_1434 (O_1434,N_9120,N_9596);
or UO_1435 (O_1435,N_9748,N_9659);
or UO_1436 (O_1436,N_9217,N_9381);
nand UO_1437 (O_1437,N_9720,N_9977);
nand UO_1438 (O_1438,N_9227,N_9055);
or UO_1439 (O_1439,N_9403,N_9325);
or UO_1440 (O_1440,N_9876,N_9928);
or UO_1441 (O_1441,N_9017,N_9877);
and UO_1442 (O_1442,N_9417,N_9044);
and UO_1443 (O_1443,N_9179,N_9945);
and UO_1444 (O_1444,N_9790,N_9037);
nor UO_1445 (O_1445,N_9851,N_9486);
and UO_1446 (O_1446,N_9594,N_9966);
nor UO_1447 (O_1447,N_9851,N_9599);
and UO_1448 (O_1448,N_9628,N_9050);
or UO_1449 (O_1449,N_9223,N_9981);
or UO_1450 (O_1450,N_9006,N_9146);
or UO_1451 (O_1451,N_9582,N_9830);
or UO_1452 (O_1452,N_9216,N_9658);
nand UO_1453 (O_1453,N_9856,N_9222);
nor UO_1454 (O_1454,N_9387,N_9758);
nor UO_1455 (O_1455,N_9361,N_9897);
nand UO_1456 (O_1456,N_9469,N_9035);
nand UO_1457 (O_1457,N_9583,N_9358);
and UO_1458 (O_1458,N_9335,N_9439);
nand UO_1459 (O_1459,N_9659,N_9270);
or UO_1460 (O_1460,N_9175,N_9534);
nand UO_1461 (O_1461,N_9363,N_9971);
or UO_1462 (O_1462,N_9641,N_9069);
or UO_1463 (O_1463,N_9276,N_9986);
nand UO_1464 (O_1464,N_9452,N_9844);
nor UO_1465 (O_1465,N_9055,N_9578);
nor UO_1466 (O_1466,N_9944,N_9709);
nand UO_1467 (O_1467,N_9115,N_9356);
nand UO_1468 (O_1468,N_9562,N_9789);
nand UO_1469 (O_1469,N_9451,N_9045);
nor UO_1470 (O_1470,N_9381,N_9284);
or UO_1471 (O_1471,N_9036,N_9419);
xnor UO_1472 (O_1472,N_9365,N_9062);
nand UO_1473 (O_1473,N_9213,N_9094);
nand UO_1474 (O_1474,N_9700,N_9333);
and UO_1475 (O_1475,N_9639,N_9413);
nor UO_1476 (O_1476,N_9172,N_9635);
nand UO_1477 (O_1477,N_9010,N_9134);
or UO_1478 (O_1478,N_9134,N_9394);
nand UO_1479 (O_1479,N_9965,N_9515);
nand UO_1480 (O_1480,N_9000,N_9588);
nor UO_1481 (O_1481,N_9156,N_9402);
or UO_1482 (O_1482,N_9659,N_9360);
or UO_1483 (O_1483,N_9728,N_9953);
nor UO_1484 (O_1484,N_9350,N_9096);
nor UO_1485 (O_1485,N_9204,N_9287);
and UO_1486 (O_1486,N_9381,N_9275);
or UO_1487 (O_1487,N_9225,N_9011);
and UO_1488 (O_1488,N_9490,N_9842);
or UO_1489 (O_1489,N_9582,N_9129);
and UO_1490 (O_1490,N_9764,N_9745);
nand UO_1491 (O_1491,N_9518,N_9540);
nor UO_1492 (O_1492,N_9511,N_9033);
nand UO_1493 (O_1493,N_9170,N_9630);
and UO_1494 (O_1494,N_9931,N_9002);
and UO_1495 (O_1495,N_9089,N_9464);
nor UO_1496 (O_1496,N_9914,N_9137);
and UO_1497 (O_1497,N_9084,N_9721);
nor UO_1498 (O_1498,N_9905,N_9265);
nor UO_1499 (O_1499,N_9091,N_9266);
endmodule