module basic_500_3000_500_30_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_484,In_249);
nand U1 (N_1,In_310,In_261);
nand U2 (N_2,In_430,In_102);
or U3 (N_3,In_356,In_133);
and U4 (N_4,In_23,In_213);
xnor U5 (N_5,In_383,In_331);
xor U6 (N_6,In_347,In_245);
nor U7 (N_7,In_62,In_175);
or U8 (N_8,In_312,In_16);
and U9 (N_9,In_176,In_151);
and U10 (N_10,In_147,In_264);
nor U11 (N_11,In_355,In_468);
or U12 (N_12,In_266,In_348);
nor U13 (N_13,In_464,In_224);
xnor U14 (N_14,In_72,In_30);
and U15 (N_15,In_271,In_453);
or U16 (N_16,In_214,In_193);
nand U17 (N_17,In_218,In_126);
and U18 (N_18,In_398,In_64);
xnor U19 (N_19,In_56,In_119);
or U20 (N_20,In_40,In_365);
or U21 (N_21,In_286,In_387);
nand U22 (N_22,In_444,In_194);
or U23 (N_23,In_199,In_483);
nand U24 (N_24,In_88,In_159);
or U25 (N_25,In_423,In_259);
or U26 (N_26,In_183,In_225);
and U27 (N_27,In_234,In_118);
nor U28 (N_28,In_201,In_309);
and U29 (N_29,In_390,In_306);
nor U30 (N_30,In_180,In_343);
nor U31 (N_31,In_366,In_247);
nor U32 (N_32,In_212,In_408);
nor U33 (N_33,In_168,In_152);
nand U34 (N_34,In_163,In_221);
and U35 (N_35,In_396,In_144);
or U36 (N_36,In_295,In_113);
nand U37 (N_37,In_27,In_217);
and U38 (N_38,In_307,In_139);
or U39 (N_39,In_31,In_303);
nor U40 (N_40,In_291,In_110);
nor U41 (N_41,In_389,In_246);
nand U42 (N_42,In_50,In_316);
and U43 (N_43,In_281,In_216);
nand U44 (N_44,In_162,In_374);
or U45 (N_45,In_317,In_82);
nor U46 (N_46,In_459,In_388);
nor U47 (N_47,In_172,In_420);
xor U48 (N_48,In_380,In_449);
and U49 (N_49,In_495,In_385);
nor U50 (N_50,In_4,In_368);
and U51 (N_51,In_418,In_447);
nor U52 (N_52,In_196,In_65);
nand U53 (N_53,In_9,In_74);
or U54 (N_54,In_223,In_392);
xor U55 (N_55,In_142,In_498);
or U56 (N_56,In_215,In_43);
and U57 (N_57,In_230,In_240);
xnor U58 (N_58,In_367,In_149);
nor U59 (N_59,In_269,In_238);
nor U60 (N_60,In_260,In_128);
nor U61 (N_61,In_273,In_283);
and U62 (N_62,In_340,In_421);
nor U63 (N_63,In_78,In_476);
nand U64 (N_64,In_403,In_422);
and U65 (N_65,In_58,In_85);
nand U66 (N_66,In_485,In_177);
or U67 (N_67,In_333,In_148);
nor U68 (N_68,In_101,In_410);
xor U69 (N_69,In_41,In_222);
nor U70 (N_70,In_233,In_258);
or U71 (N_71,In_252,In_256);
or U72 (N_72,In_489,In_397);
nand U73 (N_73,In_37,In_141);
nand U74 (N_74,In_15,In_318);
nand U75 (N_75,In_63,In_446);
or U76 (N_76,In_254,In_10);
and U77 (N_77,In_253,In_198);
and U78 (N_78,In_154,In_315);
or U79 (N_79,In_123,In_12);
or U80 (N_80,In_106,In_320);
nand U81 (N_81,In_170,In_61);
and U82 (N_82,In_125,In_300);
or U83 (N_83,In_376,In_470);
or U84 (N_84,In_436,In_441);
nand U85 (N_85,In_293,In_25);
or U86 (N_86,In_130,In_332);
nand U87 (N_87,In_54,In_33);
and U88 (N_88,In_44,In_276);
and U89 (N_89,In_415,In_275);
nor U90 (N_90,In_490,In_330);
and U91 (N_91,In_465,In_399);
or U92 (N_92,In_463,In_229);
and U93 (N_93,In_478,In_429);
or U94 (N_94,In_475,In_250);
nor U95 (N_95,In_143,In_450);
xnor U96 (N_96,In_69,In_140);
and U97 (N_97,In_358,In_416);
xor U98 (N_98,In_265,In_278);
nor U99 (N_99,In_158,In_34);
nand U100 (N_100,In_442,In_192);
or U101 (N_101,In_112,N_84);
nand U102 (N_102,In_386,N_69);
nand U103 (N_103,N_86,In_499);
nand U104 (N_104,In_481,In_434);
nor U105 (N_105,In_104,In_406);
or U106 (N_106,In_182,In_328);
and U107 (N_107,N_90,N_99);
or U108 (N_108,In_482,In_301);
and U109 (N_109,In_381,N_18);
nand U110 (N_110,In_155,In_277);
or U111 (N_111,In_362,In_363);
and U112 (N_112,In_53,N_43);
and U113 (N_113,In_164,In_136);
or U114 (N_114,In_279,In_288);
nand U115 (N_115,In_89,In_471);
nand U116 (N_116,In_129,In_409);
or U117 (N_117,N_32,N_98);
or U118 (N_118,In_68,In_13);
or U119 (N_119,In_174,In_60);
nand U120 (N_120,N_93,In_157);
nor U121 (N_121,In_431,N_73);
nor U122 (N_122,In_357,In_339);
nor U123 (N_123,In_379,N_56);
and U124 (N_124,In_86,N_16);
nor U125 (N_125,In_166,N_10);
or U126 (N_126,In_137,In_179);
nand U127 (N_127,In_91,In_97);
or U128 (N_128,In_92,In_469);
and U129 (N_129,In_462,In_372);
nand U130 (N_130,In_395,In_351);
nor U131 (N_131,In_268,N_29);
or U132 (N_132,In_321,In_493);
xnor U133 (N_133,In_116,In_94);
nand U134 (N_134,In_435,In_2);
nand U135 (N_135,In_319,In_121);
and U136 (N_136,In_427,In_346);
xor U137 (N_137,In_134,In_364);
and U138 (N_138,In_373,In_243);
or U139 (N_139,In_454,N_92);
or U140 (N_140,In_1,In_477);
nor U141 (N_141,In_443,In_298);
or U142 (N_142,In_71,In_494);
or U143 (N_143,In_207,N_2);
nor U144 (N_144,In_313,In_325);
xnor U145 (N_145,In_404,N_85);
or U146 (N_146,In_305,In_83);
or U147 (N_147,In_57,In_46);
and U148 (N_148,In_248,N_44);
and U149 (N_149,In_341,N_26);
nor U150 (N_150,In_433,N_70);
or U151 (N_151,In_208,In_28);
nand U152 (N_152,N_39,In_487);
nor U153 (N_153,N_4,N_95);
and U154 (N_154,N_5,In_20);
nor U155 (N_155,N_80,In_178);
nand U156 (N_156,In_210,N_20);
and U157 (N_157,In_496,In_282);
xor U158 (N_158,In_29,In_336);
nor U159 (N_159,N_82,N_81);
xor U160 (N_160,In_255,In_107);
or U161 (N_161,In_439,In_456);
nor U162 (N_162,N_61,In_426);
nand U163 (N_163,In_437,In_287);
or U164 (N_164,In_231,In_272);
nor U165 (N_165,In_417,In_105);
or U166 (N_166,In_262,In_70);
nor U167 (N_167,N_36,In_93);
nand U168 (N_168,In_311,In_251);
and U169 (N_169,In_467,In_304);
nand U170 (N_170,In_413,In_81);
nor U171 (N_171,In_244,In_349);
and U172 (N_172,In_146,In_440);
nand U173 (N_173,N_3,In_38);
nand U174 (N_174,In_18,In_200);
or U175 (N_175,In_377,N_96);
and U176 (N_176,In_438,N_79);
nand U177 (N_177,In_480,In_322);
nand U178 (N_178,N_47,In_411);
or U179 (N_179,N_64,N_67);
nor U180 (N_180,In_263,In_184);
or U181 (N_181,N_30,In_384);
and U182 (N_182,N_57,In_202);
xor U183 (N_183,In_36,In_419);
nor U184 (N_184,In_460,In_370);
nand U185 (N_185,In_100,In_32);
nor U186 (N_186,In_451,N_34);
and U187 (N_187,N_31,In_90);
nor U188 (N_188,N_9,In_189);
nand U189 (N_189,In_219,In_492);
nor U190 (N_190,In_242,In_472);
or U191 (N_191,In_48,In_227);
xnor U192 (N_192,In_375,In_280);
nand U193 (N_193,In_235,In_402);
and U194 (N_194,N_8,N_51);
nand U195 (N_195,In_17,In_424);
and U196 (N_196,In_455,N_83);
or U197 (N_197,In_486,In_80);
and U198 (N_198,In_488,In_160);
nor U199 (N_199,In_205,In_432);
nand U200 (N_200,In_120,In_117);
and U201 (N_201,N_193,In_84);
and U202 (N_202,N_40,N_144);
nand U203 (N_203,In_302,In_173);
nand U204 (N_204,In_3,N_161);
or U205 (N_205,In_87,N_19);
and U206 (N_206,N_177,In_285);
and U207 (N_207,In_382,In_352);
nand U208 (N_208,In_24,In_479);
nand U209 (N_209,In_314,N_75);
nand U210 (N_210,N_163,In_145);
and U211 (N_211,N_198,In_354);
and U212 (N_212,In_337,In_115);
nor U213 (N_213,N_120,In_491);
nand U214 (N_214,N_171,N_111);
nand U215 (N_215,N_78,In_39);
nor U216 (N_216,N_185,In_239);
nor U217 (N_217,In_21,N_188);
and U218 (N_218,In_49,In_26);
and U219 (N_219,N_141,In_414);
nor U220 (N_220,N_88,In_114);
or U221 (N_221,N_89,N_172);
nand U222 (N_222,N_13,N_128);
and U223 (N_223,N_117,N_129);
and U224 (N_224,N_174,N_194);
nor U225 (N_225,N_71,In_323);
nor U226 (N_226,N_11,In_237);
nor U227 (N_227,N_156,N_136);
nor U228 (N_228,In_11,In_324);
and U229 (N_229,In_42,N_33);
or U230 (N_230,In_452,In_35);
xor U231 (N_231,N_189,N_178);
and U232 (N_232,N_27,N_76);
nor U233 (N_233,N_22,N_41);
xor U234 (N_234,In_47,In_197);
nor U235 (N_235,In_77,In_400);
nor U236 (N_236,In_156,N_175);
or U237 (N_237,In_445,In_191);
and U238 (N_238,N_133,N_25);
xor U239 (N_239,N_182,N_153);
or U240 (N_240,N_199,N_157);
nor U241 (N_241,N_52,In_6);
nor U242 (N_242,In_359,In_0);
nand U243 (N_243,In_206,N_151);
nand U244 (N_244,In_329,In_232);
or U245 (N_245,N_147,In_211);
xnor U246 (N_246,N_110,N_107);
nand U247 (N_247,In_59,In_96);
nor U248 (N_248,N_169,N_58);
nor U249 (N_249,In_103,In_108);
and U250 (N_250,N_100,In_76);
nor U251 (N_251,In_360,In_122);
and U252 (N_252,In_52,N_145);
nor U253 (N_253,In_45,N_130);
nand U254 (N_254,In_161,In_135);
nor U255 (N_255,N_134,In_289);
and U256 (N_256,N_118,N_104);
nand U257 (N_257,N_24,In_371);
nor U258 (N_258,N_17,N_127);
xnor U259 (N_259,In_66,N_168);
nor U260 (N_260,N_46,N_102);
nand U261 (N_261,In_308,N_101);
and U262 (N_262,N_28,N_195);
xor U263 (N_263,In_497,In_267);
or U264 (N_264,In_342,In_401);
nor U265 (N_265,N_126,N_38);
or U266 (N_266,In_187,In_131);
nor U267 (N_267,N_77,In_220);
nor U268 (N_268,N_137,N_119);
nand U269 (N_269,In_353,In_473);
nand U270 (N_270,N_91,In_284);
nor U271 (N_271,N_87,In_350);
nor U272 (N_272,In_296,N_63);
xor U273 (N_273,In_7,In_378);
and U274 (N_274,N_105,N_186);
nor U275 (N_275,N_113,In_407);
nand U276 (N_276,N_184,In_190);
nor U277 (N_277,N_150,N_165);
or U278 (N_278,N_109,N_158);
nand U279 (N_279,In_369,In_270);
nor U280 (N_280,N_135,N_162);
or U281 (N_281,In_458,In_292);
or U282 (N_282,N_42,N_121);
or U283 (N_283,In_405,N_74);
xnor U284 (N_284,In_150,N_176);
nor U285 (N_285,In_299,N_191);
nand U286 (N_286,N_143,In_75);
nor U287 (N_287,In_412,In_297);
and U288 (N_288,In_393,In_165);
nor U289 (N_289,N_116,In_361);
and U290 (N_290,N_54,In_290);
or U291 (N_291,In_274,N_125);
and U292 (N_292,In_195,N_12);
nor U293 (N_293,In_391,In_394);
and U294 (N_294,N_45,N_66);
xnor U295 (N_295,N_123,N_72);
or U296 (N_296,N_149,N_68);
nor U297 (N_297,In_55,N_140);
and U298 (N_298,In_19,In_204);
or U299 (N_299,In_127,N_164);
or U300 (N_300,In_109,In_448);
nand U301 (N_301,N_231,N_299);
nor U302 (N_302,N_192,N_211);
and U303 (N_303,N_112,In_5);
nand U304 (N_304,N_228,N_205);
xnor U305 (N_305,In_334,In_132);
nor U306 (N_306,N_196,N_94);
xnor U307 (N_307,N_97,N_212);
and U308 (N_308,N_114,N_279);
or U309 (N_309,In_338,In_186);
and U310 (N_310,In_203,N_260);
nand U311 (N_311,N_284,N_255);
xor U312 (N_312,In_188,N_122);
nor U313 (N_313,N_293,In_185);
nand U314 (N_314,N_197,N_257);
nor U315 (N_315,In_327,N_282);
nand U316 (N_316,In_95,N_225);
or U317 (N_317,N_187,N_274);
nor U318 (N_318,N_222,N_138);
nand U319 (N_319,N_55,In_51);
or U320 (N_320,N_287,N_170);
nand U321 (N_321,N_270,N_243);
nor U322 (N_322,N_209,N_294);
nand U323 (N_323,In_344,N_227);
nand U324 (N_324,N_290,In_171);
and U325 (N_325,N_297,In_79);
nand U326 (N_326,N_234,In_457);
or U327 (N_327,N_263,N_60);
and U328 (N_328,N_232,N_264);
nand U329 (N_329,In_345,N_259);
or U330 (N_330,N_167,N_59);
nand U331 (N_331,N_217,N_155);
or U332 (N_332,N_131,N_224);
nand U333 (N_333,N_160,N_292);
nor U334 (N_334,N_179,N_190);
or U335 (N_335,In_67,N_166);
nor U336 (N_336,In_474,N_249);
or U337 (N_337,N_220,N_244);
nand U338 (N_338,N_237,N_236);
and U339 (N_339,In_8,In_241);
or U340 (N_340,N_298,N_6);
or U341 (N_341,N_267,In_138);
nand U342 (N_342,N_247,N_254);
and U343 (N_343,In_73,N_251);
nand U344 (N_344,N_124,N_278);
and U345 (N_345,N_230,In_167);
or U346 (N_346,In_22,N_139);
and U347 (N_347,N_245,N_277);
nand U348 (N_348,N_65,N_281);
nor U349 (N_349,In_257,N_203);
nor U350 (N_350,N_200,N_288);
or U351 (N_351,N_248,N_62);
and U352 (N_352,In_228,N_233);
and U353 (N_353,N_48,In_466);
nor U354 (N_354,N_23,N_202);
nand U355 (N_355,N_108,N_272);
nand U356 (N_356,N_214,N_173);
nor U357 (N_357,N_271,N_280);
nand U358 (N_358,In_428,N_0);
or U359 (N_359,N_265,In_335);
and U360 (N_360,N_37,N_268);
nand U361 (N_361,N_159,N_49);
nor U362 (N_362,N_204,N_14);
or U363 (N_363,In_14,N_180);
xnor U364 (N_364,N_296,In_111);
nor U365 (N_365,N_242,N_266);
and U366 (N_366,N_286,N_148);
or U367 (N_367,N_7,N_223);
or U368 (N_368,N_207,N_276);
and U369 (N_369,In_294,In_98);
nor U370 (N_370,N_35,N_183);
or U371 (N_371,In_169,N_262);
xnor U372 (N_372,In_226,In_461);
and U373 (N_373,N_239,N_50);
nor U374 (N_374,N_246,N_154);
or U375 (N_375,N_215,N_221);
nand U376 (N_376,N_226,N_285);
nor U377 (N_377,In_236,N_210);
nor U378 (N_378,N_146,N_240);
nor U379 (N_379,N_213,N_208);
and U380 (N_380,N_289,N_229);
or U381 (N_381,In_326,In_153);
nor U382 (N_382,N_142,N_261);
xnor U383 (N_383,In_181,N_269);
nor U384 (N_384,N_201,N_106);
and U385 (N_385,In_209,N_275);
and U386 (N_386,N_218,N_252);
nand U387 (N_387,In_99,N_235);
nor U388 (N_388,N_253,N_295);
nor U389 (N_389,N_219,N_241);
nor U390 (N_390,N_258,N_291);
or U391 (N_391,N_15,N_21);
xnor U392 (N_392,N_206,N_53);
nand U393 (N_393,N_256,N_181);
nor U394 (N_394,N_1,In_425);
nor U395 (N_395,In_124,N_152);
or U396 (N_396,N_103,N_115);
or U397 (N_397,N_238,N_216);
xnor U398 (N_398,N_283,N_273);
and U399 (N_399,N_250,N_132);
nand U400 (N_400,N_367,N_358);
nor U401 (N_401,N_334,N_308);
and U402 (N_402,N_369,N_366);
or U403 (N_403,N_365,N_363);
or U404 (N_404,N_332,N_321);
and U405 (N_405,N_330,N_300);
nor U406 (N_406,N_372,N_325);
nor U407 (N_407,N_318,N_379);
xnor U408 (N_408,N_315,N_364);
and U409 (N_409,N_314,N_347);
xnor U410 (N_410,N_370,N_380);
or U411 (N_411,N_335,N_377);
and U412 (N_412,N_337,N_399);
and U413 (N_413,N_305,N_336);
nor U414 (N_414,N_385,N_386);
nor U415 (N_415,N_313,N_339);
or U416 (N_416,N_357,N_304);
or U417 (N_417,N_307,N_371);
nor U418 (N_418,N_397,N_303);
xor U419 (N_419,N_394,N_343);
or U420 (N_420,N_338,N_348);
xor U421 (N_421,N_353,N_333);
or U422 (N_422,N_355,N_317);
and U423 (N_423,N_387,N_324);
and U424 (N_424,N_352,N_354);
nand U425 (N_425,N_316,N_345);
nor U426 (N_426,N_320,N_349);
and U427 (N_427,N_329,N_327);
nand U428 (N_428,N_309,N_374);
or U429 (N_429,N_312,N_395);
or U430 (N_430,N_375,N_392);
nand U431 (N_431,N_361,N_378);
nand U432 (N_432,N_342,N_368);
nand U433 (N_433,N_328,N_359);
nand U434 (N_434,N_362,N_350);
and U435 (N_435,N_391,N_346);
or U436 (N_436,N_310,N_381);
and U437 (N_437,N_383,N_306);
nand U438 (N_438,N_398,N_389);
nor U439 (N_439,N_311,N_356);
and U440 (N_440,N_384,N_376);
nor U441 (N_441,N_322,N_331);
and U442 (N_442,N_396,N_360);
nand U443 (N_443,N_373,N_390);
xnor U444 (N_444,N_344,N_319);
xor U445 (N_445,N_302,N_341);
or U446 (N_446,N_340,N_388);
nand U447 (N_447,N_323,N_326);
or U448 (N_448,N_351,N_301);
and U449 (N_449,N_393,N_382);
or U450 (N_450,N_326,N_363);
nor U451 (N_451,N_379,N_349);
or U452 (N_452,N_394,N_325);
nor U453 (N_453,N_360,N_355);
xor U454 (N_454,N_346,N_357);
or U455 (N_455,N_310,N_347);
xnor U456 (N_456,N_399,N_315);
xnor U457 (N_457,N_324,N_326);
or U458 (N_458,N_395,N_376);
and U459 (N_459,N_340,N_352);
or U460 (N_460,N_346,N_318);
or U461 (N_461,N_393,N_384);
and U462 (N_462,N_375,N_341);
or U463 (N_463,N_303,N_335);
or U464 (N_464,N_311,N_375);
nor U465 (N_465,N_365,N_376);
and U466 (N_466,N_370,N_304);
or U467 (N_467,N_306,N_398);
nand U468 (N_468,N_344,N_399);
or U469 (N_469,N_334,N_384);
or U470 (N_470,N_394,N_384);
nand U471 (N_471,N_307,N_385);
nand U472 (N_472,N_332,N_353);
nor U473 (N_473,N_366,N_328);
xor U474 (N_474,N_309,N_398);
or U475 (N_475,N_322,N_315);
or U476 (N_476,N_379,N_344);
nand U477 (N_477,N_387,N_334);
or U478 (N_478,N_367,N_305);
nor U479 (N_479,N_356,N_380);
xnor U480 (N_480,N_320,N_352);
and U481 (N_481,N_376,N_361);
or U482 (N_482,N_323,N_351);
or U483 (N_483,N_360,N_308);
nor U484 (N_484,N_381,N_385);
or U485 (N_485,N_395,N_310);
xnor U486 (N_486,N_384,N_357);
or U487 (N_487,N_385,N_371);
and U488 (N_488,N_384,N_324);
nor U489 (N_489,N_332,N_362);
xor U490 (N_490,N_341,N_381);
and U491 (N_491,N_347,N_320);
and U492 (N_492,N_373,N_364);
or U493 (N_493,N_394,N_323);
and U494 (N_494,N_352,N_338);
and U495 (N_495,N_374,N_315);
nor U496 (N_496,N_313,N_377);
nor U497 (N_497,N_350,N_308);
nand U498 (N_498,N_336,N_318);
nor U499 (N_499,N_379,N_350);
nand U500 (N_500,N_489,N_495);
and U501 (N_501,N_464,N_437);
nor U502 (N_502,N_413,N_456);
nand U503 (N_503,N_491,N_414);
or U504 (N_504,N_453,N_482);
nor U505 (N_505,N_472,N_462);
and U506 (N_506,N_496,N_481);
nand U507 (N_507,N_442,N_412);
and U508 (N_508,N_410,N_436);
and U509 (N_509,N_475,N_465);
xor U510 (N_510,N_468,N_490);
or U511 (N_511,N_433,N_457);
nand U512 (N_512,N_455,N_476);
and U513 (N_513,N_429,N_497);
and U514 (N_514,N_424,N_486);
and U515 (N_515,N_469,N_423);
and U516 (N_516,N_441,N_443);
nand U517 (N_517,N_480,N_417);
or U518 (N_518,N_485,N_473);
xnor U519 (N_519,N_404,N_467);
nor U520 (N_520,N_411,N_419);
nor U521 (N_521,N_409,N_438);
xnor U522 (N_522,N_493,N_406);
nor U523 (N_523,N_405,N_488);
and U524 (N_524,N_458,N_479);
nor U525 (N_525,N_432,N_449);
nor U526 (N_526,N_445,N_471);
nor U527 (N_527,N_439,N_401);
xnor U528 (N_528,N_454,N_416);
nand U529 (N_529,N_427,N_498);
nor U530 (N_530,N_444,N_492);
nand U531 (N_531,N_403,N_460);
or U532 (N_532,N_422,N_466);
nand U533 (N_533,N_415,N_448);
and U534 (N_534,N_430,N_440);
nor U535 (N_535,N_447,N_450);
nand U536 (N_536,N_434,N_420);
or U537 (N_537,N_499,N_484);
and U538 (N_538,N_494,N_461);
nor U539 (N_539,N_487,N_459);
nand U540 (N_540,N_478,N_435);
or U541 (N_541,N_418,N_463);
nand U542 (N_542,N_452,N_425);
or U543 (N_543,N_402,N_428);
and U544 (N_544,N_431,N_421);
nand U545 (N_545,N_426,N_407);
and U546 (N_546,N_477,N_400);
or U547 (N_547,N_451,N_474);
and U548 (N_548,N_446,N_483);
or U549 (N_549,N_408,N_470);
or U550 (N_550,N_406,N_490);
nor U551 (N_551,N_461,N_467);
xor U552 (N_552,N_405,N_413);
or U553 (N_553,N_441,N_417);
xor U554 (N_554,N_448,N_460);
nor U555 (N_555,N_422,N_463);
and U556 (N_556,N_442,N_408);
xor U557 (N_557,N_492,N_441);
nand U558 (N_558,N_457,N_486);
nand U559 (N_559,N_489,N_404);
nand U560 (N_560,N_477,N_413);
and U561 (N_561,N_462,N_488);
and U562 (N_562,N_412,N_471);
nand U563 (N_563,N_417,N_432);
xor U564 (N_564,N_471,N_464);
nor U565 (N_565,N_465,N_482);
or U566 (N_566,N_434,N_489);
nand U567 (N_567,N_466,N_429);
nand U568 (N_568,N_496,N_411);
and U569 (N_569,N_494,N_432);
nand U570 (N_570,N_415,N_499);
and U571 (N_571,N_433,N_489);
nor U572 (N_572,N_498,N_484);
or U573 (N_573,N_465,N_471);
nand U574 (N_574,N_423,N_436);
xor U575 (N_575,N_448,N_406);
or U576 (N_576,N_467,N_471);
or U577 (N_577,N_413,N_417);
nor U578 (N_578,N_450,N_458);
nor U579 (N_579,N_443,N_424);
nand U580 (N_580,N_411,N_470);
nand U581 (N_581,N_428,N_430);
nand U582 (N_582,N_465,N_416);
and U583 (N_583,N_469,N_461);
nor U584 (N_584,N_405,N_465);
nor U585 (N_585,N_473,N_451);
and U586 (N_586,N_418,N_446);
nor U587 (N_587,N_483,N_494);
nand U588 (N_588,N_467,N_435);
and U589 (N_589,N_498,N_471);
nor U590 (N_590,N_448,N_400);
or U591 (N_591,N_403,N_402);
nor U592 (N_592,N_491,N_465);
nor U593 (N_593,N_465,N_443);
xor U594 (N_594,N_499,N_471);
or U595 (N_595,N_478,N_433);
and U596 (N_596,N_400,N_494);
nand U597 (N_597,N_478,N_492);
or U598 (N_598,N_415,N_436);
or U599 (N_599,N_416,N_414);
nand U600 (N_600,N_516,N_536);
or U601 (N_601,N_566,N_511);
or U602 (N_602,N_553,N_584);
xnor U603 (N_603,N_545,N_573);
or U604 (N_604,N_509,N_592);
and U605 (N_605,N_580,N_519);
nor U606 (N_606,N_530,N_586);
nand U607 (N_607,N_598,N_503);
nand U608 (N_608,N_578,N_507);
nor U609 (N_609,N_548,N_587);
or U610 (N_610,N_557,N_554);
or U611 (N_611,N_569,N_577);
nor U612 (N_612,N_506,N_588);
or U613 (N_613,N_561,N_502);
xnor U614 (N_614,N_527,N_581);
nor U615 (N_615,N_513,N_547);
nand U616 (N_616,N_543,N_518);
and U617 (N_617,N_528,N_575);
or U618 (N_618,N_538,N_514);
xnor U619 (N_619,N_582,N_560);
nor U620 (N_620,N_500,N_552);
nand U621 (N_621,N_549,N_534);
nand U622 (N_622,N_526,N_537);
nor U623 (N_623,N_517,N_550);
nor U624 (N_624,N_521,N_558);
xnor U625 (N_625,N_594,N_576);
nand U626 (N_626,N_564,N_535);
nor U627 (N_627,N_520,N_541);
or U628 (N_628,N_510,N_504);
xor U629 (N_629,N_529,N_544);
nor U630 (N_630,N_546,N_501);
or U631 (N_631,N_539,N_571);
nand U632 (N_632,N_597,N_591);
nor U633 (N_633,N_556,N_567);
and U634 (N_634,N_562,N_515);
or U635 (N_635,N_533,N_579);
and U636 (N_636,N_522,N_525);
and U637 (N_637,N_551,N_523);
nor U638 (N_638,N_531,N_524);
or U639 (N_639,N_565,N_508);
or U640 (N_640,N_583,N_542);
nor U641 (N_641,N_532,N_505);
xnor U642 (N_642,N_593,N_563);
xor U643 (N_643,N_574,N_596);
or U644 (N_644,N_599,N_559);
nand U645 (N_645,N_589,N_512);
xnor U646 (N_646,N_585,N_590);
or U647 (N_647,N_572,N_570);
and U648 (N_648,N_555,N_568);
and U649 (N_649,N_595,N_540);
xor U650 (N_650,N_526,N_587);
nand U651 (N_651,N_557,N_573);
nor U652 (N_652,N_559,N_540);
or U653 (N_653,N_596,N_587);
and U654 (N_654,N_571,N_583);
and U655 (N_655,N_590,N_544);
nor U656 (N_656,N_501,N_516);
or U657 (N_657,N_530,N_562);
or U658 (N_658,N_551,N_584);
or U659 (N_659,N_538,N_596);
and U660 (N_660,N_595,N_531);
and U661 (N_661,N_509,N_593);
nand U662 (N_662,N_548,N_529);
and U663 (N_663,N_533,N_512);
nand U664 (N_664,N_583,N_521);
xor U665 (N_665,N_577,N_560);
and U666 (N_666,N_560,N_595);
nor U667 (N_667,N_532,N_559);
or U668 (N_668,N_525,N_509);
and U669 (N_669,N_587,N_543);
nor U670 (N_670,N_572,N_591);
nand U671 (N_671,N_576,N_539);
xnor U672 (N_672,N_537,N_595);
and U673 (N_673,N_560,N_551);
and U674 (N_674,N_565,N_520);
and U675 (N_675,N_525,N_577);
xor U676 (N_676,N_595,N_553);
nor U677 (N_677,N_588,N_565);
nand U678 (N_678,N_510,N_591);
and U679 (N_679,N_535,N_509);
and U680 (N_680,N_547,N_599);
nor U681 (N_681,N_586,N_591);
nor U682 (N_682,N_504,N_596);
xnor U683 (N_683,N_568,N_559);
nand U684 (N_684,N_523,N_550);
nor U685 (N_685,N_538,N_560);
nor U686 (N_686,N_519,N_510);
xor U687 (N_687,N_506,N_551);
or U688 (N_688,N_557,N_576);
and U689 (N_689,N_519,N_578);
xnor U690 (N_690,N_592,N_585);
or U691 (N_691,N_551,N_510);
nand U692 (N_692,N_504,N_554);
nand U693 (N_693,N_527,N_585);
nand U694 (N_694,N_511,N_500);
xnor U695 (N_695,N_546,N_553);
nor U696 (N_696,N_513,N_577);
xor U697 (N_697,N_563,N_599);
nor U698 (N_698,N_563,N_535);
and U699 (N_699,N_571,N_547);
and U700 (N_700,N_619,N_610);
nand U701 (N_701,N_602,N_672);
nand U702 (N_702,N_674,N_627);
or U703 (N_703,N_655,N_690);
or U704 (N_704,N_696,N_661);
and U705 (N_705,N_676,N_623);
nor U706 (N_706,N_626,N_648);
nor U707 (N_707,N_614,N_645);
and U708 (N_708,N_673,N_637);
or U709 (N_709,N_621,N_657);
nor U710 (N_710,N_603,N_612);
or U711 (N_711,N_699,N_600);
or U712 (N_712,N_670,N_669);
nand U713 (N_713,N_606,N_671);
nand U714 (N_714,N_682,N_639);
nor U715 (N_715,N_692,N_636);
or U716 (N_716,N_634,N_675);
nand U717 (N_717,N_664,N_654);
nor U718 (N_718,N_601,N_697);
and U719 (N_719,N_644,N_658);
and U720 (N_720,N_668,N_622);
nor U721 (N_721,N_611,N_686);
nand U722 (N_722,N_698,N_632);
and U723 (N_723,N_631,N_618);
nand U724 (N_724,N_646,N_643);
and U725 (N_725,N_684,N_604);
or U726 (N_726,N_656,N_679);
nor U727 (N_727,N_681,N_624);
nor U728 (N_728,N_638,N_653);
or U729 (N_729,N_641,N_680);
xor U730 (N_730,N_683,N_642);
nor U731 (N_731,N_620,N_666);
nor U732 (N_732,N_613,N_647);
nand U733 (N_733,N_607,N_652);
nor U734 (N_734,N_695,N_689);
or U735 (N_735,N_650,N_693);
and U736 (N_736,N_629,N_628);
or U737 (N_737,N_677,N_615);
xor U738 (N_738,N_625,N_605);
and U739 (N_739,N_688,N_691);
and U740 (N_740,N_665,N_609);
nor U741 (N_741,N_667,N_617);
nand U742 (N_742,N_663,N_635);
nand U743 (N_743,N_633,N_685);
and U744 (N_744,N_640,N_662);
or U745 (N_745,N_616,N_651);
nand U746 (N_746,N_608,N_630);
nand U747 (N_747,N_649,N_687);
nor U748 (N_748,N_659,N_678);
and U749 (N_749,N_660,N_694);
or U750 (N_750,N_659,N_627);
nor U751 (N_751,N_614,N_689);
or U752 (N_752,N_695,N_628);
nand U753 (N_753,N_637,N_687);
or U754 (N_754,N_673,N_655);
nor U755 (N_755,N_698,N_669);
xor U756 (N_756,N_643,N_622);
and U757 (N_757,N_657,N_637);
and U758 (N_758,N_610,N_624);
nand U759 (N_759,N_684,N_616);
or U760 (N_760,N_667,N_611);
and U761 (N_761,N_625,N_611);
nand U762 (N_762,N_686,N_677);
and U763 (N_763,N_640,N_607);
nand U764 (N_764,N_621,N_666);
and U765 (N_765,N_681,N_623);
xor U766 (N_766,N_690,N_627);
and U767 (N_767,N_694,N_600);
nand U768 (N_768,N_686,N_610);
nand U769 (N_769,N_655,N_643);
xnor U770 (N_770,N_642,N_673);
nor U771 (N_771,N_601,N_634);
or U772 (N_772,N_658,N_667);
or U773 (N_773,N_639,N_691);
nand U774 (N_774,N_628,N_634);
or U775 (N_775,N_646,N_679);
xnor U776 (N_776,N_635,N_652);
or U777 (N_777,N_683,N_664);
nand U778 (N_778,N_609,N_681);
nand U779 (N_779,N_675,N_688);
nor U780 (N_780,N_699,N_648);
nand U781 (N_781,N_642,N_653);
and U782 (N_782,N_602,N_698);
nor U783 (N_783,N_678,N_665);
or U784 (N_784,N_616,N_673);
nand U785 (N_785,N_644,N_682);
nand U786 (N_786,N_619,N_641);
and U787 (N_787,N_625,N_614);
nor U788 (N_788,N_652,N_699);
and U789 (N_789,N_676,N_656);
nor U790 (N_790,N_656,N_638);
and U791 (N_791,N_674,N_678);
nor U792 (N_792,N_627,N_676);
or U793 (N_793,N_680,N_618);
and U794 (N_794,N_679,N_677);
and U795 (N_795,N_645,N_600);
nor U796 (N_796,N_661,N_604);
nor U797 (N_797,N_612,N_618);
nand U798 (N_798,N_678,N_676);
xnor U799 (N_799,N_660,N_621);
nand U800 (N_800,N_720,N_778);
nand U801 (N_801,N_709,N_767);
nor U802 (N_802,N_701,N_797);
or U803 (N_803,N_707,N_781);
xor U804 (N_804,N_703,N_744);
and U805 (N_805,N_754,N_761);
and U806 (N_806,N_723,N_788);
nand U807 (N_807,N_741,N_757);
and U808 (N_808,N_798,N_724);
nor U809 (N_809,N_708,N_752);
xnor U810 (N_810,N_766,N_704);
or U811 (N_811,N_710,N_783);
and U812 (N_812,N_748,N_729);
nand U813 (N_813,N_700,N_779);
nor U814 (N_814,N_759,N_776);
nand U815 (N_815,N_790,N_719);
and U816 (N_816,N_751,N_718);
and U817 (N_817,N_702,N_732);
and U818 (N_818,N_736,N_784);
or U819 (N_819,N_743,N_764);
nand U820 (N_820,N_711,N_731);
nand U821 (N_821,N_737,N_787);
nand U822 (N_822,N_742,N_745);
nor U823 (N_823,N_717,N_728);
and U824 (N_824,N_771,N_772);
or U825 (N_825,N_756,N_760);
or U826 (N_826,N_730,N_777);
xor U827 (N_827,N_739,N_746);
nand U828 (N_828,N_722,N_735);
nand U829 (N_829,N_795,N_716);
nand U830 (N_830,N_738,N_727);
and U831 (N_831,N_714,N_793);
nor U832 (N_832,N_749,N_715);
and U833 (N_833,N_782,N_786);
and U834 (N_834,N_791,N_789);
nand U835 (N_835,N_750,N_796);
and U836 (N_836,N_765,N_706);
xnor U837 (N_837,N_799,N_725);
or U838 (N_838,N_763,N_755);
xor U839 (N_839,N_758,N_773);
and U840 (N_840,N_768,N_792);
nand U841 (N_841,N_780,N_712);
nor U842 (N_842,N_753,N_785);
xnor U843 (N_843,N_794,N_774);
nand U844 (N_844,N_740,N_747);
and U845 (N_845,N_769,N_733);
and U846 (N_846,N_705,N_721);
or U847 (N_847,N_770,N_734);
nor U848 (N_848,N_775,N_713);
nand U849 (N_849,N_726,N_762);
nor U850 (N_850,N_719,N_724);
nor U851 (N_851,N_747,N_704);
and U852 (N_852,N_717,N_766);
xor U853 (N_853,N_787,N_727);
or U854 (N_854,N_736,N_743);
or U855 (N_855,N_712,N_735);
or U856 (N_856,N_777,N_720);
nand U857 (N_857,N_736,N_767);
or U858 (N_858,N_725,N_724);
or U859 (N_859,N_712,N_764);
and U860 (N_860,N_745,N_789);
xnor U861 (N_861,N_773,N_766);
and U862 (N_862,N_722,N_760);
nor U863 (N_863,N_791,N_783);
nand U864 (N_864,N_785,N_704);
nor U865 (N_865,N_724,N_764);
nor U866 (N_866,N_785,N_766);
xor U867 (N_867,N_765,N_708);
nand U868 (N_868,N_737,N_750);
nor U869 (N_869,N_708,N_748);
nor U870 (N_870,N_738,N_767);
and U871 (N_871,N_707,N_744);
nand U872 (N_872,N_787,N_776);
and U873 (N_873,N_763,N_754);
nor U874 (N_874,N_760,N_700);
and U875 (N_875,N_703,N_793);
and U876 (N_876,N_731,N_720);
xnor U877 (N_877,N_731,N_776);
xor U878 (N_878,N_718,N_739);
or U879 (N_879,N_789,N_792);
or U880 (N_880,N_795,N_751);
nand U881 (N_881,N_788,N_780);
nand U882 (N_882,N_707,N_735);
xor U883 (N_883,N_716,N_729);
and U884 (N_884,N_750,N_742);
and U885 (N_885,N_778,N_779);
nand U886 (N_886,N_749,N_779);
xor U887 (N_887,N_713,N_752);
nor U888 (N_888,N_778,N_734);
nor U889 (N_889,N_795,N_771);
and U890 (N_890,N_790,N_707);
and U891 (N_891,N_796,N_774);
or U892 (N_892,N_752,N_741);
or U893 (N_893,N_769,N_711);
nor U894 (N_894,N_753,N_732);
nand U895 (N_895,N_744,N_799);
nor U896 (N_896,N_764,N_731);
nor U897 (N_897,N_790,N_740);
or U898 (N_898,N_779,N_759);
and U899 (N_899,N_718,N_728);
nor U900 (N_900,N_887,N_810);
and U901 (N_901,N_860,N_893);
nor U902 (N_902,N_827,N_894);
nand U903 (N_903,N_825,N_823);
or U904 (N_904,N_806,N_870);
nor U905 (N_905,N_867,N_804);
and U906 (N_906,N_817,N_820);
or U907 (N_907,N_815,N_895);
and U908 (N_908,N_819,N_828);
nor U909 (N_909,N_868,N_813);
and U910 (N_910,N_837,N_843);
or U911 (N_911,N_809,N_863);
nor U912 (N_912,N_832,N_845);
and U913 (N_913,N_852,N_853);
and U914 (N_914,N_841,N_814);
nand U915 (N_915,N_802,N_826);
nand U916 (N_916,N_833,N_822);
or U917 (N_917,N_875,N_899);
nor U918 (N_918,N_842,N_877);
or U919 (N_919,N_840,N_850);
xnor U920 (N_920,N_897,N_882);
xnor U921 (N_921,N_800,N_896);
and U922 (N_922,N_859,N_866);
nand U923 (N_923,N_891,N_857);
or U924 (N_924,N_846,N_862);
and U925 (N_925,N_872,N_869);
or U926 (N_926,N_879,N_865);
nor U927 (N_927,N_885,N_886);
nor U928 (N_928,N_871,N_881);
nor U929 (N_929,N_874,N_824);
or U930 (N_930,N_856,N_829);
nor U931 (N_931,N_873,N_851);
nand U932 (N_932,N_888,N_880);
or U933 (N_933,N_858,N_812);
or U934 (N_934,N_830,N_834);
nand U935 (N_935,N_889,N_801);
nand U936 (N_936,N_861,N_876);
xnor U937 (N_937,N_898,N_849);
nand U938 (N_938,N_847,N_892);
or U939 (N_939,N_884,N_805);
nand U940 (N_940,N_848,N_818);
or U941 (N_941,N_835,N_803);
nor U942 (N_942,N_839,N_838);
nor U943 (N_943,N_844,N_807);
and U944 (N_944,N_855,N_811);
or U945 (N_945,N_878,N_821);
xnor U946 (N_946,N_836,N_816);
nand U947 (N_947,N_864,N_808);
and U948 (N_948,N_890,N_854);
nand U949 (N_949,N_883,N_831);
xor U950 (N_950,N_847,N_857);
nor U951 (N_951,N_824,N_858);
nor U952 (N_952,N_881,N_822);
or U953 (N_953,N_818,N_804);
nor U954 (N_954,N_848,N_817);
or U955 (N_955,N_860,N_878);
nand U956 (N_956,N_807,N_821);
or U957 (N_957,N_894,N_830);
xor U958 (N_958,N_826,N_881);
or U959 (N_959,N_896,N_849);
nand U960 (N_960,N_881,N_873);
xnor U961 (N_961,N_863,N_895);
or U962 (N_962,N_840,N_883);
nor U963 (N_963,N_810,N_873);
and U964 (N_964,N_810,N_888);
and U965 (N_965,N_807,N_845);
nor U966 (N_966,N_860,N_827);
or U967 (N_967,N_848,N_804);
nor U968 (N_968,N_823,N_829);
nand U969 (N_969,N_865,N_854);
and U970 (N_970,N_813,N_865);
or U971 (N_971,N_833,N_826);
or U972 (N_972,N_802,N_860);
nand U973 (N_973,N_829,N_847);
or U974 (N_974,N_854,N_812);
nand U975 (N_975,N_827,N_838);
nand U976 (N_976,N_881,N_866);
nand U977 (N_977,N_868,N_818);
and U978 (N_978,N_844,N_847);
nor U979 (N_979,N_863,N_836);
and U980 (N_980,N_819,N_867);
and U981 (N_981,N_851,N_867);
and U982 (N_982,N_892,N_823);
nand U983 (N_983,N_873,N_839);
or U984 (N_984,N_887,N_859);
nand U985 (N_985,N_893,N_896);
and U986 (N_986,N_813,N_850);
and U987 (N_987,N_876,N_872);
nor U988 (N_988,N_872,N_837);
nand U989 (N_989,N_878,N_805);
and U990 (N_990,N_870,N_875);
or U991 (N_991,N_807,N_852);
or U992 (N_992,N_830,N_861);
or U993 (N_993,N_823,N_864);
and U994 (N_994,N_890,N_844);
nand U995 (N_995,N_860,N_828);
nor U996 (N_996,N_849,N_893);
and U997 (N_997,N_829,N_800);
and U998 (N_998,N_897,N_848);
xnor U999 (N_999,N_894,N_831);
nor U1000 (N_1000,N_991,N_913);
or U1001 (N_1001,N_953,N_940);
and U1002 (N_1002,N_978,N_944);
nand U1003 (N_1003,N_968,N_922);
and U1004 (N_1004,N_904,N_936);
nor U1005 (N_1005,N_998,N_945);
nor U1006 (N_1006,N_965,N_906);
or U1007 (N_1007,N_973,N_972);
or U1008 (N_1008,N_933,N_901);
nand U1009 (N_1009,N_900,N_975);
nand U1010 (N_1010,N_961,N_930);
nand U1011 (N_1011,N_988,N_918);
or U1012 (N_1012,N_917,N_957);
or U1013 (N_1013,N_948,N_929);
xnor U1014 (N_1014,N_974,N_934);
or U1015 (N_1015,N_966,N_999);
xnor U1016 (N_1016,N_912,N_971);
and U1017 (N_1017,N_985,N_914);
and U1018 (N_1018,N_947,N_946);
or U1019 (N_1019,N_942,N_928);
or U1020 (N_1020,N_954,N_952);
or U1021 (N_1021,N_915,N_916);
and U1022 (N_1022,N_949,N_939);
or U1023 (N_1023,N_935,N_970);
nand U1024 (N_1024,N_969,N_996);
nor U1025 (N_1025,N_994,N_993);
xnor U1026 (N_1026,N_921,N_977);
and U1027 (N_1027,N_938,N_963);
nand U1028 (N_1028,N_937,N_995);
nand U1029 (N_1029,N_926,N_909);
xnor U1030 (N_1030,N_984,N_924);
xnor U1031 (N_1031,N_958,N_927);
nor U1032 (N_1032,N_951,N_907);
and U1033 (N_1033,N_964,N_983);
nor U1034 (N_1034,N_982,N_941);
or U1035 (N_1035,N_981,N_920);
nand U1036 (N_1036,N_910,N_919);
nor U1037 (N_1037,N_902,N_923);
nor U1038 (N_1038,N_962,N_960);
or U1039 (N_1039,N_959,N_950);
nor U1040 (N_1040,N_931,N_956);
nand U1041 (N_1041,N_987,N_989);
nand U1042 (N_1042,N_925,N_976);
and U1043 (N_1043,N_911,N_979);
nor U1044 (N_1044,N_955,N_997);
xnor U1045 (N_1045,N_908,N_903);
nand U1046 (N_1046,N_943,N_967);
xnor U1047 (N_1047,N_992,N_905);
xnor U1048 (N_1048,N_932,N_990);
or U1049 (N_1049,N_986,N_980);
nor U1050 (N_1050,N_919,N_914);
or U1051 (N_1051,N_989,N_984);
nand U1052 (N_1052,N_933,N_938);
nor U1053 (N_1053,N_991,N_932);
or U1054 (N_1054,N_914,N_976);
and U1055 (N_1055,N_915,N_994);
or U1056 (N_1056,N_924,N_910);
nand U1057 (N_1057,N_992,N_921);
or U1058 (N_1058,N_958,N_975);
or U1059 (N_1059,N_981,N_987);
and U1060 (N_1060,N_935,N_971);
nor U1061 (N_1061,N_990,N_989);
nand U1062 (N_1062,N_956,N_915);
and U1063 (N_1063,N_928,N_960);
xnor U1064 (N_1064,N_969,N_959);
nor U1065 (N_1065,N_990,N_950);
or U1066 (N_1066,N_909,N_995);
xnor U1067 (N_1067,N_924,N_930);
nand U1068 (N_1068,N_964,N_929);
or U1069 (N_1069,N_911,N_976);
xor U1070 (N_1070,N_918,N_958);
and U1071 (N_1071,N_916,N_987);
nor U1072 (N_1072,N_989,N_993);
nor U1073 (N_1073,N_993,N_947);
and U1074 (N_1074,N_916,N_939);
or U1075 (N_1075,N_962,N_919);
nand U1076 (N_1076,N_906,N_917);
or U1077 (N_1077,N_908,N_944);
nand U1078 (N_1078,N_947,N_963);
nand U1079 (N_1079,N_945,N_981);
nor U1080 (N_1080,N_920,N_940);
and U1081 (N_1081,N_999,N_926);
nand U1082 (N_1082,N_929,N_933);
or U1083 (N_1083,N_904,N_907);
nor U1084 (N_1084,N_929,N_983);
nand U1085 (N_1085,N_916,N_919);
and U1086 (N_1086,N_909,N_983);
nand U1087 (N_1087,N_994,N_972);
nor U1088 (N_1088,N_974,N_990);
or U1089 (N_1089,N_994,N_914);
xnor U1090 (N_1090,N_938,N_954);
nand U1091 (N_1091,N_991,N_955);
nor U1092 (N_1092,N_985,N_915);
and U1093 (N_1093,N_921,N_969);
nor U1094 (N_1094,N_963,N_953);
or U1095 (N_1095,N_954,N_981);
xor U1096 (N_1096,N_911,N_909);
nand U1097 (N_1097,N_951,N_967);
nor U1098 (N_1098,N_990,N_942);
nand U1099 (N_1099,N_963,N_955);
nor U1100 (N_1100,N_1085,N_1013);
xnor U1101 (N_1101,N_1011,N_1004);
xor U1102 (N_1102,N_1033,N_1063);
nor U1103 (N_1103,N_1005,N_1024);
or U1104 (N_1104,N_1023,N_1083);
or U1105 (N_1105,N_1040,N_1064);
xor U1106 (N_1106,N_1018,N_1047);
nand U1107 (N_1107,N_1087,N_1015);
or U1108 (N_1108,N_1007,N_1074);
or U1109 (N_1109,N_1052,N_1091);
and U1110 (N_1110,N_1030,N_1067);
or U1111 (N_1111,N_1060,N_1003);
xnor U1112 (N_1112,N_1088,N_1062);
nor U1113 (N_1113,N_1036,N_1043);
nor U1114 (N_1114,N_1080,N_1079);
or U1115 (N_1115,N_1069,N_1057);
nor U1116 (N_1116,N_1045,N_1029);
nor U1117 (N_1117,N_1010,N_1000);
or U1118 (N_1118,N_1026,N_1009);
and U1119 (N_1119,N_1096,N_1055);
nand U1120 (N_1120,N_1049,N_1006);
and U1121 (N_1121,N_1031,N_1099);
and U1122 (N_1122,N_1044,N_1072);
nor U1123 (N_1123,N_1092,N_1051);
nand U1124 (N_1124,N_1027,N_1037);
nor U1125 (N_1125,N_1019,N_1098);
nand U1126 (N_1126,N_1066,N_1056);
nor U1127 (N_1127,N_1077,N_1054);
nor U1128 (N_1128,N_1078,N_1002);
and U1129 (N_1129,N_1035,N_1028);
xnor U1130 (N_1130,N_1082,N_1008);
and U1131 (N_1131,N_1073,N_1071);
or U1132 (N_1132,N_1012,N_1053);
nand U1133 (N_1133,N_1059,N_1068);
and U1134 (N_1134,N_1081,N_1070);
xnor U1135 (N_1135,N_1034,N_1050);
or U1136 (N_1136,N_1089,N_1076);
and U1137 (N_1137,N_1014,N_1093);
or U1138 (N_1138,N_1095,N_1075);
nand U1139 (N_1139,N_1039,N_1042);
and U1140 (N_1140,N_1046,N_1001);
and U1141 (N_1141,N_1025,N_1097);
xor U1142 (N_1142,N_1086,N_1032);
xnor U1143 (N_1143,N_1094,N_1017);
nor U1144 (N_1144,N_1065,N_1016);
and U1145 (N_1145,N_1058,N_1022);
nand U1146 (N_1146,N_1041,N_1084);
nor U1147 (N_1147,N_1038,N_1061);
xor U1148 (N_1148,N_1090,N_1020);
or U1149 (N_1149,N_1021,N_1048);
nand U1150 (N_1150,N_1025,N_1038);
or U1151 (N_1151,N_1002,N_1083);
nand U1152 (N_1152,N_1094,N_1037);
or U1153 (N_1153,N_1001,N_1031);
nand U1154 (N_1154,N_1065,N_1028);
or U1155 (N_1155,N_1029,N_1083);
or U1156 (N_1156,N_1091,N_1002);
nor U1157 (N_1157,N_1050,N_1020);
or U1158 (N_1158,N_1096,N_1095);
and U1159 (N_1159,N_1007,N_1086);
nand U1160 (N_1160,N_1092,N_1046);
nand U1161 (N_1161,N_1098,N_1086);
and U1162 (N_1162,N_1019,N_1083);
nor U1163 (N_1163,N_1069,N_1065);
nor U1164 (N_1164,N_1000,N_1007);
or U1165 (N_1165,N_1054,N_1088);
nor U1166 (N_1166,N_1038,N_1028);
or U1167 (N_1167,N_1001,N_1061);
nand U1168 (N_1168,N_1093,N_1034);
nand U1169 (N_1169,N_1090,N_1055);
nor U1170 (N_1170,N_1089,N_1022);
nand U1171 (N_1171,N_1046,N_1004);
or U1172 (N_1172,N_1006,N_1036);
nand U1173 (N_1173,N_1098,N_1036);
nand U1174 (N_1174,N_1021,N_1046);
or U1175 (N_1175,N_1027,N_1019);
and U1176 (N_1176,N_1007,N_1005);
nand U1177 (N_1177,N_1086,N_1042);
nand U1178 (N_1178,N_1053,N_1033);
and U1179 (N_1179,N_1015,N_1070);
or U1180 (N_1180,N_1063,N_1051);
nor U1181 (N_1181,N_1049,N_1092);
or U1182 (N_1182,N_1065,N_1038);
and U1183 (N_1183,N_1018,N_1078);
and U1184 (N_1184,N_1084,N_1040);
and U1185 (N_1185,N_1083,N_1040);
nor U1186 (N_1186,N_1009,N_1099);
or U1187 (N_1187,N_1062,N_1054);
and U1188 (N_1188,N_1083,N_1077);
or U1189 (N_1189,N_1062,N_1024);
nor U1190 (N_1190,N_1018,N_1040);
or U1191 (N_1191,N_1071,N_1024);
nor U1192 (N_1192,N_1093,N_1096);
xor U1193 (N_1193,N_1073,N_1080);
nor U1194 (N_1194,N_1079,N_1062);
nor U1195 (N_1195,N_1002,N_1055);
nor U1196 (N_1196,N_1048,N_1006);
or U1197 (N_1197,N_1013,N_1098);
nor U1198 (N_1198,N_1034,N_1051);
nor U1199 (N_1199,N_1045,N_1091);
or U1200 (N_1200,N_1149,N_1107);
nand U1201 (N_1201,N_1161,N_1121);
nor U1202 (N_1202,N_1164,N_1180);
nand U1203 (N_1203,N_1110,N_1165);
and U1204 (N_1204,N_1198,N_1181);
nor U1205 (N_1205,N_1144,N_1178);
or U1206 (N_1206,N_1142,N_1191);
xnor U1207 (N_1207,N_1113,N_1132);
xnor U1208 (N_1208,N_1128,N_1133);
xor U1209 (N_1209,N_1129,N_1103);
xnor U1210 (N_1210,N_1158,N_1123);
xnor U1211 (N_1211,N_1101,N_1171);
and U1212 (N_1212,N_1193,N_1188);
nor U1213 (N_1213,N_1184,N_1156);
nor U1214 (N_1214,N_1100,N_1186);
and U1215 (N_1215,N_1197,N_1130);
nand U1216 (N_1216,N_1166,N_1176);
or U1217 (N_1217,N_1170,N_1177);
nor U1218 (N_1218,N_1192,N_1114);
or U1219 (N_1219,N_1131,N_1106);
nand U1220 (N_1220,N_1104,N_1190);
nor U1221 (N_1221,N_1147,N_1117);
nand U1222 (N_1222,N_1134,N_1120);
nor U1223 (N_1223,N_1127,N_1138);
and U1224 (N_1224,N_1141,N_1153);
nand U1225 (N_1225,N_1116,N_1145);
and U1226 (N_1226,N_1111,N_1163);
and U1227 (N_1227,N_1136,N_1183);
nand U1228 (N_1228,N_1119,N_1102);
xnor U1229 (N_1229,N_1135,N_1162);
nor U1230 (N_1230,N_1152,N_1169);
nand U1231 (N_1231,N_1194,N_1125);
and U1232 (N_1232,N_1168,N_1146);
or U1233 (N_1233,N_1148,N_1124);
nand U1234 (N_1234,N_1143,N_1196);
xnor U1235 (N_1235,N_1172,N_1122);
nand U1236 (N_1236,N_1167,N_1189);
and U1237 (N_1237,N_1155,N_1199);
nor U1238 (N_1238,N_1173,N_1108);
nor U1239 (N_1239,N_1105,N_1157);
or U1240 (N_1240,N_1187,N_1179);
or U1241 (N_1241,N_1174,N_1151);
or U1242 (N_1242,N_1154,N_1112);
or U1243 (N_1243,N_1126,N_1175);
or U1244 (N_1244,N_1182,N_1137);
and U1245 (N_1245,N_1185,N_1159);
nand U1246 (N_1246,N_1109,N_1150);
and U1247 (N_1247,N_1140,N_1160);
and U1248 (N_1248,N_1115,N_1139);
and U1249 (N_1249,N_1195,N_1118);
and U1250 (N_1250,N_1194,N_1178);
nand U1251 (N_1251,N_1162,N_1163);
and U1252 (N_1252,N_1177,N_1187);
or U1253 (N_1253,N_1189,N_1177);
nor U1254 (N_1254,N_1165,N_1188);
or U1255 (N_1255,N_1118,N_1170);
xnor U1256 (N_1256,N_1113,N_1160);
and U1257 (N_1257,N_1195,N_1119);
nand U1258 (N_1258,N_1161,N_1118);
and U1259 (N_1259,N_1107,N_1128);
and U1260 (N_1260,N_1153,N_1196);
and U1261 (N_1261,N_1120,N_1194);
nor U1262 (N_1262,N_1119,N_1127);
nor U1263 (N_1263,N_1155,N_1107);
nand U1264 (N_1264,N_1102,N_1135);
or U1265 (N_1265,N_1187,N_1102);
or U1266 (N_1266,N_1144,N_1188);
nor U1267 (N_1267,N_1198,N_1168);
nand U1268 (N_1268,N_1122,N_1146);
or U1269 (N_1269,N_1121,N_1114);
xor U1270 (N_1270,N_1146,N_1140);
nor U1271 (N_1271,N_1140,N_1122);
xnor U1272 (N_1272,N_1163,N_1183);
or U1273 (N_1273,N_1181,N_1115);
or U1274 (N_1274,N_1109,N_1152);
nor U1275 (N_1275,N_1183,N_1101);
or U1276 (N_1276,N_1186,N_1141);
or U1277 (N_1277,N_1130,N_1157);
nand U1278 (N_1278,N_1186,N_1102);
nor U1279 (N_1279,N_1107,N_1166);
xor U1280 (N_1280,N_1138,N_1144);
nor U1281 (N_1281,N_1114,N_1171);
and U1282 (N_1282,N_1178,N_1154);
and U1283 (N_1283,N_1107,N_1179);
and U1284 (N_1284,N_1155,N_1167);
or U1285 (N_1285,N_1184,N_1188);
nand U1286 (N_1286,N_1157,N_1177);
nor U1287 (N_1287,N_1147,N_1185);
xnor U1288 (N_1288,N_1173,N_1117);
nor U1289 (N_1289,N_1104,N_1154);
and U1290 (N_1290,N_1160,N_1162);
and U1291 (N_1291,N_1114,N_1154);
nand U1292 (N_1292,N_1140,N_1186);
nand U1293 (N_1293,N_1123,N_1130);
or U1294 (N_1294,N_1192,N_1138);
or U1295 (N_1295,N_1174,N_1102);
nor U1296 (N_1296,N_1171,N_1118);
and U1297 (N_1297,N_1114,N_1106);
nand U1298 (N_1298,N_1174,N_1149);
nand U1299 (N_1299,N_1111,N_1148);
nor U1300 (N_1300,N_1292,N_1212);
nand U1301 (N_1301,N_1265,N_1299);
xnor U1302 (N_1302,N_1235,N_1229);
nand U1303 (N_1303,N_1250,N_1200);
or U1304 (N_1304,N_1240,N_1243);
xor U1305 (N_1305,N_1272,N_1204);
or U1306 (N_1306,N_1263,N_1251);
nand U1307 (N_1307,N_1257,N_1201);
xnor U1308 (N_1308,N_1232,N_1217);
or U1309 (N_1309,N_1287,N_1258);
or U1310 (N_1310,N_1249,N_1225);
xor U1311 (N_1311,N_1289,N_1276);
and U1312 (N_1312,N_1260,N_1226);
nor U1313 (N_1313,N_1291,N_1262);
or U1314 (N_1314,N_1254,N_1237);
and U1315 (N_1315,N_1239,N_1206);
nand U1316 (N_1316,N_1278,N_1293);
nand U1317 (N_1317,N_1261,N_1284);
xor U1318 (N_1318,N_1238,N_1283);
and U1319 (N_1319,N_1253,N_1202);
xor U1320 (N_1320,N_1203,N_1208);
nand U1321 (N_1321,N_1288,N_1221);
or U1322 (N_1322,N_1266,N_1285);
nor U1323 (N_1323,N_1282,N_1209);
and U1324 (N_1324,N_1270,N_1223);
or U1325 (N_1325,N_1268,N_1271);
xnor U1326 (N_1326,N_1246,N_1205);
nand U1327 (N_1327,N_1286,N_1236);
nand U1328 (N_1328,N_1218,N_1222);
or U1329 (N_1329,N_1273,N_1279);
xnor U1330 (N_1330,N_1255,N_1298);
xor U1331 (N_1331,N_1297,N_1277);
or U1332 (N_1332,N_1220,N_1233);
nor U1333 (N_1333,N_1215,N_1296);
nor U1334 (N_1334,N_1227,N_1247);
and U1335 (N_1335,N_1252,N_1230);
nand U1336 (N_1336,N_1211,N_1234);
nor U1337 (N_1337,N_1245,N_1295);
xnor U1338 (N_1338,N_1294,N_1274);
nor U1339 (N_1339,N_1214,N_1248);
and U1340 (N_1340,N_1244,N_1241);
nor U1341 (N_1341,N_1213,N_1269);
nand U1342 (N_1342,N_1207,N_1264);
and U1343 (N_1343,N_1259,N_1275);
nor U1344 (N_1344,N_1280,N_1281);
or U1345 (N_1345,N_1216,N_1290);
and U1346 (N_1346,N_1231,N_1256);
and U1347 (N_1347,N_1219,N_1224);
nand U1348 (N_1348,N_1242,N_1228);
or U1349 (N_1349,N_1267,N_1210);
nor U1350 (N_1350,N_1207,N_1258);
nor U1351 (N_1351,N_1257,N_1267);
or U1352 (N_1352,N_1221,N_1234);
nand U1353 (N_1353,N_1278,N_1204);
nand U1354 (N_1354,N_1204,N_1228);
nand U1355 (N_1355,N_1222,N_1215);
and U1356 (N_1356,N_1204,N_1236);
or U1357 (N_1357,N_1225,N_1201);
nand U1358 (N_1358,N_1249,N_1251);
nand U1359 (N_1359,N_1281,N_1250);
nand U1360 (N_1360,N_1263,N_1239);
nor U1361 (N_1361,N_1279,N_1200);
and U1362 (N_1362,N_1281,N_1203);
or U1363 (N_1363,N_1292,N_1281);
nor U1364 (N_1364,N_1275,N_1283);
or U1365 (N_1365,N_1291,N_1298);
xor U1366 (N_1366,N_1271,N_1298);
and U1367 (N_1367,N_1202,N_1257);
xor U1368 (N_1368,N_1259,N_1250);
or U1369 (N_1369,N_1297,N_1282);
and U1370 (N_1370,N_1264,N_1203);
nor U1371 (N_1371,N_1204,N_1218);
and U1372 (N_1372,N_1236,N_1255);
and U1373 (N_1373,N_1293,N_1256);
or U1374 (N_1374,N_1297,N_1292);
nor U1375 (N_1375,N_1297,N_1220);
or U1376 (N_1376,N_1256,N_1243);
and U1377 (N_1377,N_1215,N_1292);
or U1378 (N_1378,N_1265,N_1287);
nor U1379 (N_1379,N_1251,N_1228);
nor U1380 (N_1380,N_1281,N_1231);
and U1381 (N_1381,N_1299,N_1232);
nand U1382 (N_1382,N_1216,N_1217);
nand U1383 (N_1383,N_1232,N_1243);
nor U1384 (N_1384,N_1202,N_1247);
nand U1385 (N_1385,N_1221,N_1248);
xnor U1386 (N_1386,N_1233,N_1296);
nand U1387 (N_1387,N_1221,N_1283);
or U1388 (N_1388,N_1219,N_1254);
nand U1389 (N_1389,N_1238,N_1268);
nand U1390 (N_1390,N_1241,N_1287);
nor U1391 (N_1391,N_1205,N_1241);
nand U1392 (N_1392,N_1239,N_1277);
nand U1393 (N_1393,N_1200,N_1238);
and U1394 (N_1394,N_1226,N_1232);
or U1395 (N_1395,N_1266,N_1210);
or U1396 (N_1396,N_1273,N_1268);
and U1397 (N_1397,N_1272,N_1248);
nand U1398 (N_1398,N_1274,N_1291);
xnor U1399 (N_1399,N_1258,N_1255);
nor U1400 (N_1400,N_1303,N_1321);
nor U1401 (N_1401,N_1351,N_1319);
nor U1402 (N_1402,N_1368,N_1334);
xnor U1403 (N_1403,N_1385,N_1313);
and U1404 (N_1404,N_1307,N_1373);
and U1405 (N_1405,N_1300,N_1360);
nor U1406 (N_1406,N_1324,N_1359);
xnor U1407 (N_1407,N_1371,N_1386);
or U1408 (N_1408,N_1357,N_1315);
nor U1409 (N_1409,N_1397,N_1390);
or U1410 (N_1410,N_1328,N_1394);
nand U1411 (N_1411,N_1344,N_1356);
nor U1412 (N_1412,N_1389,N_1388);
nand U1413 (N_1413,N_1302,N_1339);
or U1414 (N_1414,N_1345,N_1354);
or U1415 (N_1415,N_1304,N_1367);
and U1416 (N_1416,N_1301,N_1379);
nand U1417 (N_1417,N_1375,N_1322);
or U1418 (N_1418,N_1378,N_1333);
nor U1419 (N_1419,N_1347,N_1399);
nor U1420 (N_1420,N_1325,N_1336);
xor U1421 (N_1421,N_1393,N_1374);
xor U1422 (N_1422,N_1392,N_1384);
and U1423 (N_1423,N_1330,N_1363);
or U1424 (N_1424,N_1350,N_1342);
nand U1425 (N_1425,N_1355,N_1396);
or U1426 (N_1426,N_1376,N_1377);
nand U1427 (N_1427,N_1369,N_1306);
nor U1428 (N_1428,N_1318,N_1381);
and U1429 (N_1429,N_1364,N_1372);
nor U1430 (N_1430,N_1395,N_1348);
or U1431 (N_1431,N_1343,N_1308);
nand U1432 (N_1432,N_1305,N_1332);
nand U1433 (N_1433,N_1335,N_1331);
nor U1434 (N_1434,N_1387,N_1340);
and U1435 (N_1435,N_1362,N_1311);
nor U1436 (N_1436,N_1380,N_1310);
and U1437 (N_1437,N_1391,N_1365);
or U1438 (N_1438,N_1320,N_1341);
and U1439 (N_1439,N_1327,N_1317);
or U1440 (N_1440,N_1312,N_1382);
xor U1441 (N_1441,N_1316,N_1398);
xor U1442 (N_1442,N_1358,N_1326);
and U1443 (N_1443,N_1370,N_1338);
xnor U1444 (N_1444,N_1366,N_1329);
nand U1445 (N_1445,N_1361,N_1309);
nand U1446 (N_1446,N_1349,N_1314);
or U1447 (N_1447,N_1353,N_1352);
and U1448 (N_1448,N_1346,N_1323);
nor U1449 (N_1449,N_1337,N_1383);
nand U1450 (N_1450,N_1353,N_1348);
nor U1451 (N_1451,N_1355,N_1382);
or U1452 (N_1452,N_1373,N_1382);
and U1453 (N_1453,N_1348,N_1386);
xnor U1454 (N_1454,N_1356,N_1382);
nand U1455 (N_1455,N_1389,N_1332);
or U1456 (N_1456,N_1327,N_1356);
nand U1457 (N_1457,N_1327,N_1322);
nor U1458 (N_1458,N_1399,N_1316);
nor U1459 (N_1459,N_1319,N_1359);
nand U1460 (N_1460,N_1362,N_1327);
nor U1461 (N_1461,N_1376,N_1301);
nor U1462 (N_1462,N_1383,N_1339);
and U1463 (N_1463,N_1356,N_1391);
or U1464 (N_1464,N_1309,N_1335);
or U1465 (N_1465,N_1337,N_1338);
xor U1466 (N_1466,N_1311,N_1319);
xor U1467 (N_1467,N_1316,N_1310);
nand U1468 (N_1468,N_1321,N_1328);
and U1469 (N_1469,N_1323,N_1325);
and U1470 (N_1470,N_1384,N_1342);
nor U1471 (N_1471,N_1317,N_1378);
nand U1472 (N_1472,N_1312,N_1363);
and U1473 (N_1473,N_1307,N_1394);
nand U1474 (N_1474,N_1343,N_1388);
nor U1475 (N_1475,N_1359,N_1303);
xnor U1476 (N_1476,N_1367,N_1311);
or U1477 (N_1477,N_1383,N_1326);
and U1478 (N_1478,N_1362,N_1368);
or U1479 (N_1479,N_1329,N_1365);
nor U1480 (N_1480,N_1311,N_1344);
and U1481 (N_1481,N_1306,N_1376);
and U1482 (N_1482,N_1337,N_1392);
or U1483 (N_1483,N_1319,N_1364);
and U1484 (N_1484,N_1355,N_1343);
or U1485 (N_1485,N_1330,N_1313);
and U1486 (N_1486,N_1345,N_1389);
nand U1487 (N_1487,N_1304,N_1332);
and U1488 (N_1488,N_1330,N_1336);
or U1489 (N_1489,N_1342,N_1397);
or U1490 (N_1490,N_1337,N_1302);
or U1491 (N_1491,N_1321,N_1326);
and U1492 (N_1492,N_1330,N_1351);
or U1493 (N_1493,N_1305,N_1307);
nand U1494 (N_1494,N_1352,N_1315);
nor U1495 (N_1495,N_1336,N_1333);
or U1496 (N_1496,N_1367,N_1322);
nor U1497 (N_1497,N_1371,N_1345);
and U1498 (N_1498,N_1358,N_1307);
xor U1499 (N_1499,N_1351,N_1341);
and U1500 (N_1500,N_1435,N_1444);
and U1501 (N_1501,N_1472,N_1461);
or U1502 (N_1502,N_1438,N_1430);
nand U1503 (N_1503,N_1403,N_1490);
xnor U1504 (N_1504,N_1478,N_1485);
nand U1505 (N_1505,N_1451,N_1458);
xnor U1506 (N_1506,N_1417,N_1426);
or U1507 (N_1507,N_1415,N_1421);
nand U1508 (N_1508,N_1464,N_1475);
nand U1509 (N_1509,N_1480,N_1491);
and U1510 (N_1510,N_1476,N_1405);
nand U1511 (N_1511,N_1410,N_1404);
and U1512 (N_1512,N_1470,N_1446);
xor U1513 (N_1513,N_1413,N_1482);
nor U1514 (N_1514,N_1440,N_1442);
nor U1515 (N_1515,N_1459,N_1473);
nand U1516 (N_1516,N_1474,N_1487);
nor U1517 (N_1517,N_1496,N_1489);
and U1518 (N_1518,N_1419,N_1429);
nand U1519 (N_1519,N_1424,N_1411);
xnor U1520 (N_1520,N_1462,N_1420);
nand U1521 (N_1521,N_1432,N_1467);
and U1522 (N_1522,N_1441,N_1439);
nor U1523 (N_1523,N_1437,N_1416);
and U1524 (N_1524,N_1401,N_1402);
or U1525 (N_1525,N_1428,N_1466);
nor U1526 (N_1526,N_1455,N_1448);
and U1527 (N_1527,N_1425,N_1409);
or U1528 (N_1528,N_1449,N_1406);
and U1529 (N_1529,N_1468,N_1443);
and U1530 (N_1530,N_1463,N_1422);
nand U1531 (N_1531,N_1447,N_1427);
and U1532 (N_1532,N_1434,N_1469);
nor U1533 (N_1533,N_1493,N_1481);
and U1534 (N_1534,N_1423,N_1484);
nor U1535 (N_1535,N_1498,N_1452);
nor U1536 (N_1536,N_1477,N_1407);
or U1537 (N_1537,N_1433,N_1471);
or U1538 (N_1538,N_1488,N_1456);
nand U1539 (N_1539,N_1431,N_1453);
xnor U1540 (N_1540,N_1499,N_1418);
or U1541 (N_1541,N_1483,N_1492);
nand U1542 (N_1542,N_1479,N_1497);
or U1543 (N_1543,N_1400,N_1457);
nand U1544 (N_1544,N_1436,N_1460);
nand U1545 (N_1545,N_1465,N_1486);
and U1546 (N_1546,N_1450,N_1494);
and U1547 (N_1547,N_1408,N_1412);
and U1548 (N_1548,N_1495,N_1454);
and U1549 (N_1549,N_1445,N_1414);
or U1550 (N_1550,N_1413,N_1472);
or U1551 (N_1551,N_1438,N_1476);
and U1552 (N_1552,N_1448,N_1469);
or U1553 (N_1553,N_1446,N_1452);
or U1554 (N_1554,N_1486,N_1488);
and U1555 (N_1555,N_1454,N_1437);
xor U1556 (N_1556,N_1451,N_1450);
or U1557 (N_1557,N_1447,N_1490);
nand U1558 (N_1558,N_1412,N_1495);
nor U1559 (N_1559,N_1412,N_1419);
nor U1560 (N_1560,N_1447,N_1457);
and U1561 (N_1561,N_1494,N_1411);
xor U1562 (N_1562,N_1402,N_1448);
nor U1563 (N_1563,N_1468,N_1492);
or U1564 (N_1564,N_1407,N_1456);
xnor U1565 (N_1565,N_1445,N_1403);
nand U1566 (N_1566,N_1468,N_1421);
nor U1567 (N_1567,N_1454,N_1409);
and U1568 (N_1568,N_1449,N_1473);
nor U1569 (N_1569,N_1417,N_1420);
nor U1570 (N_1570,N_1499,N_1426);
nor U1571 (N_1571,N_1466,N_1498);
nand U1572 (N_1572,N_1429,N_1473);
nand U1573 (N_1573,N_1486,N_1431);
nand U1574 (N_1574,N_1458,N_1417);
and U1575 (N_1575,N_1418,N_1411);
and U1576 (N_1576,N_1410,N_1471);
nand U1577 (N_1577,N_1473,N_1487);
nor U1578 (N_1578,N_1457,N_1409);
xor U1579 (N_1579,N_1445,N_1489);
nand U1580 (N_1580,N_1463,N_1421);
and U1581 (N_1581,N_1447,N_1464);
and U1582 (N_1582,N_1406,N_1485);
nor U1583 (N_1583,N_1463,N_1439);
and U1584 (N_1584,N_1416,N_1418);
nand U1585 (N_1585,N_1423,N_1425);
or U1586 (N_1586,N_1402,N_1435);
and U1587 (N_1587,N_1425,N_1478);
nand U1588 (N_1588,N_1448,N_1420);
nor U1589 (N_1589,N_1408,N_1435);
nor U1590 (N_1590,N_1442,N_1498);
or U1591 (N_1591,N_1409,N_1476);
nand U1592 (N_1592,N_1449,N_1447);
nand U1593 (N_1593,N_1422,N_1484);
and U1594 (N_1594,N_1402,N_1447);
and U1595 (N_1595,N_1473,N_1485);
and U1596 (N_1596,N_1422,N_1460);
or U1597 (N_1597,N_1447,N_1426);
and U1598 (N_1598,N_1447,N_1463);
xnor U1599 (N_1599,N_1458,N_1431);
and U1600 (N_1600,N_1593,N_1525);
xnor U1601 (N_1601,N_1500,N_1552);
or U1602 (N_1602,N_1522,N_1506);
xnor U1603 (N_1603,N_1585,N_1504);
nor U1604 (N_1604,N_1573,N_1536);
nand U1605 (N_1605,N_1578,N_1590);
or U1606 (N_1606,N_1532,N_1543);
and U1607 (N_1607,N_1598,N_1541);
or U1608 (N_1608,N_1571,N_1545);
or U1609 (N_1609,N_1512,N_1526);
nor U1610 (N_1610,N_1565,N_1519);
and U1611 (N_1611,N_1547,N_1594);
nand U1612 (N_1612,N_1549,N_1535);
and U1613 (N_1613,N_1508,N_1516);
or U1614 (N_1614,N_1507,N_1537);
or U1615 (N_1615,N_1557,N_1534);
nor U1616 (N_1616,N_1515,N_1599);
nand U1617 (N_1617,N_1540,N_1538);
nor U1618 (N_1618,N_1559,N_1591);
nor U1619 (N_1619,N_1530,N_1580);
nor U1620 (N_1620,N_1584,N_1509);
or U1621 (N_1621,N_1527,N_1503);
nand U1622 (N_1622,N_1539,N_1572);
nor U1623 (N_1623,N_1555,N_1595);
nor U1624 (N_1624,N_1510,N_1511);
xnor U1625 (N_1625,N_1514,N_1553);
and U1626 (N_1626,N_1579,N_1529);
nor U1627 (N_1627,N_1558,N_1533);
and U1628 (N_1628,N_1554,N_1562);
and U1629 (N_1629,N_1556,N_1505);
nor U1630 (N_1630,N_1560,N_1521);
nor U1631 (N_1631,N_1520,N_1577);
nor U1632 (N_1632,N_1586,N_1546);
nand U1633 (N_1633,N_1528,N_1596);
nand U1634 (N_1634,N_1551,N_1574);
nand U1635 (N_1635,N_1588,N_1570);
and U1636 (N_1636,N_1518,N_1575);
or U1637 (N_1637,N_1548,N_1502);
nor U1638 (N_1638,N_1513,N_1542);
nor U1639 (N_1639,N_1531,N_1524);
xor U1640 (N_1640,N_1544,N_1581);
nand U1641 (N_1641,N_1550,N_1561);
nand U1642 (N_1642,N_1564,N_1517);
nand U1643 (N_1643,N_1583,N_1566);
nand U1644 (N_1644,N_1567,N_1569);
and U1645 (N_1645,N_1501,N_1589);
and U1646 (N_1646,N_1597,N_1563);
or U1647 (N_1647,N_1568,N_1587);
or U1648 (N_1648,N_1592,N_1582);
nand U1649 (N_1649,N_1523,N_1576);
nor U1650 (N_1650,N_1522,N_1524);
nand U1651 (N_1651,N_1554,N_1552);
nor U1652 (N_1652,N_1564,N_1562);
nor U1653 (N_1653,N_1522,N_1542);
nand U1654 (N_1654,N_1521,N_1522);
nor U1655 (N_1655,N_1507,N_1525);
or U1656 (N_1656,N_1572,N_1509);
xnor U1657 (N_1657,N_1554,N_1599);
nand U1658 (N_1658,N_1593,N_1598);
and U1659 (N_1659,N_1503,N_1572);
and U1660 (N_1660,N_1572,N_1587);
nand U1661 (N_1661,N_1561,N_1569);
nor U1662 (N_1662,N_1511,N_1585);
or U1663 (N_1663,N_1540,N_1576);
nand U1664 (N_1664,N_1502,N_1518);
nand U1665 (N_1665,N_1522,N_1541);
and U1666 (N_1666,N_1537,N_1531);
nand U1667 (N_1667,N_1516,N_1555);
nand U1668 (N_1668,N_1578,N_1510);
and U1669 (N_1669,N_1580,N_1587);
and U1670 (N_1670,N_1525,N_1536);
and U1671 (N_1671,N_1580,N_1591);
and U1672 (N_1672,N_1593,N_1542);
nor U1673 (N_1673,N_1596,N_1512);
or U1674 (N_1674,N_1554,N_1568);
and U1675 (N_1675,N_1569,N_1514);
or U1676 (N_1676,N_1501,N_1518);
nor U1677 (N_1677,N_1512,N_1583);
nor U1678 (N_1678,N_1549,N_1567);
nand U1679 (N_1679,N_1565,N_1516);
nor U1680 (N_1680,N_1548,N_1572);
and U1681 (N_1681,N_1502,N_1553);
or U1682 (N_1682,N_1595,N_1550);
nand U1683 (N_1683,N_1569,N_1588);
or U1684 (N_1684,N_1514,N_1521);
nand U1685 (N_1685,N_1559,N_1505);
xnor U1686 (N_1686,N_1530,N_1548);
or U1687 (N_1687,N_1554,N_1521);
nor U1688 (N_1688,N_1552,N_1568);
nor U1689 (N_1689,N_1566,N_1528);
xnor U1690 (N_1690,N_1599,N_1503);
nand U1691 (N_1691,N_1542,N_1567);
nor U1692 (N_1692,N_1521,N_1523);
nor U1693 (N_1693,N_1542,N_1538);
nor U1694 (N_1694,N_1526,N_1541);
and U1695 (N_1695,N_1553,N_1549);
or U1696 (N_1696,N_1554,N_1567);
nor U1697 (N_1697,N_1538,N_1558);
and U1698 (N_1698,N_1596,N_1527);
or U1699 (N_1699,N_1571,N_1532);
and U1700 (N_1700,N_1655,N_1631);
or U1701 (N_1701,N_1606,N_1692);
and U1702 (N_1702,N_1687,N_1649);
or U1703 (N_1703,N_1634,N_1638);
nor U1704 (N_1704,N_1664,N_1617);
nand U1705 (N_1705,N_1632,N_1676);
or U1706 (N_1706,N_1680,N_1627);
xnor U1707 (N_1707,N_1679,N_1630);
nor U1708 (N_1708,N_1677,N_1619);
nand U1709 (N_1709,N_1645,N_1697);
or U1710 (N_1710,N_1635,N_1612);
and U1711 (N_1711,N_1628,N_1625);
and U1712 (N_1712,N_1626,N_1681);
or U1713 (N_1713,N_1646,N_1663);
xor U1714 (N_1714,N_1682,N_1667);
and U1715 (N_1715,N_1699,N_1672);
nand U1716 (N_1716,N_1661,N_1674);
or U1717 (N_1717,N_1642,N_1670);
xnor U1718 (N_1718,N_1648,N_1605);
nand U1719 (N_1719,N_1691,N_1618);
nand U1720 (N_1720,N_1621,N_1693);
or U1721 (N_1721,N_1600,N_1657);
nand U1722 (N_1722,N_1636,N_1611);
or U1723 (N_1723,N_1601,N_1666);
nor U1724 (N_1724,N_1629,N_1613);
and U1725 (N_1725,N_1668,N_1689);
or U1726 (N_1726,N_1637,N_1608);
nand U1727 (N_1727,N_1683,N_1633);
or U1728 (N_1728,N_1665,N_1622);
or U1729 (N_1729,N_1644,N_1616);
or U1730 (N_1730,N_1656,N_1671);
or U1731 (N_1731,N_1651,N_1659);
and U1732 (N_1732,N_1678,N_1669);
and U1733 (N_1733,N_1652,N_1607);
nand U1734 (N_1734,N_1641,N_1658);
nor U1735 (N_1735,N_1650,N_1686);
nor U1736 (N_1736,N_1654,N_1609);
nand U1737 (N_1737,N_1615,N_1640);
and U1738 (N_1738,N_1647,N_1675);
nor U1739 (N_1739,N_1603,N_1604);
nand U1740 (N_1740,N_1660,N_1610);
nor U1741 (N_1741,N_1639,N_1695);
nand U1742 (N_1742,N_1694,N_1684);
and U1743 (N_1743,N_1643,N_1673);
or U1744 (N_1744,N_1620,N_1624);
or U1745 (N_1745,N_1690,N_1698);
nand U1746 (N_1746,N_1602,N_1685);
xnor U1747 (N_1747,N_1653,N_1688);
nor U1748 (N_1748,N_1696,N_1623);
nor U1749 (N_1749,N_1614,N_1662);
and U1750 (N_1750,N_1621,N_1687);
nor U1751 (N_1751,N_1622,N_1626);
nor U1752 (N_1752,N_1618,N_1633);
nand U1753 (N_1753,N_1634,N_1667);
and U1754 (N_1754,N_1678,N_1625);
xor U1755 (N_1755,N_1681,N_1622);
nand U1756 (N_1756,N_1629,N_1658);
or U1757 (N_1757,N_1640,N_1628);
nor U1758 (N_1758,N_1644,N_1662);
nor U1759 (N_1759,N_1613,N_1611);
nor U1760 (N_1760,N_1664,N_1652);
nand U1761 (N_1761,N_1691,N_1670);
nand U1762 (N_1762,N_1652,N_1651);
or U1763 (N_1763,N_1641,N_1642);
and U1764 (N_1764,N_1687,N_1651);
xor U1765 (N_1765,N_1613,N_1601);
or U1766 (N_1766,N_1681,N_1664);
xnor U1767 (N_1767,N_1697,N_1648);
nand U1768 (N_1768,N_1660,N_1618);
and U1769 (N_1769,N_1648,N_1638);
xnor U1770 (N_1770,N_1694,N_1628);
and U1771 (N_1771,N_1657,N_1682);
or U1772 (N_1772,N_1609,N_1642);
nand U1773 (N_1773,N_1635,N_1610);
and U1774 (N_1774,N_1682,N_1651);
xor U1775 (N_1775,N_1622,N_1605);
nand U1776 (N_1776,N_1641,N_1601);
nand U1777 (N_1777,N_1616,N_1639);
nor U1778 (N_1778,N_1634,N_1689);
or U1779 (N_1779,N_1611,N_1642);
nand U1780 (N_1780,N_1660,N_1602);
nor U1781 (N_1781,N_1674,N_1656);
or U1782 (N_1782,N_1626,N_1683);
nand U1783 (N_1783,N_1678,N_1630);
nand U1784 (N_1784,N_1667,N_1685);
or U1785 (N_1785,N_1694,N_1662);
or U1786 (N_1786,N_1649,N_1663);
xnor U1787 (N_1787,N_1656,N_1669);
and U1788 (N_1788,N_1635,N_1625);
xnor U1789 (N_1789,N_1639,N_1663);
nor U1790 (N_1790,N_1676,N_1604);
or U1791 (N_1791,N_1613,N_1618);
or U1792 (N_1792,N_1635,N_1634);
nand U1793 (N_1793,N_1642,N_1674);
or U1794 (N_1794,N_1610,N_1665);
nor U1795 (N_1795,N_1668,N_1662);
and U1796 (N_1796,N_1642,N_1634);
nor U1797 (N_1797,N_1629,N_1677);
nand U1798 (N_1798,N_1645,N_1600);
nor U1799 (N_1799,N_1637,N_1694);
xor U1800 (N_1800,N_1754,N_1799);
nand U1801 (N_1801,N_1740,N_1772);
nor U1802 (N_1802,N_1704,N_1738);
nand U1803 (N_1803,N_1712,N_1723);
nand U1804 (N_1804,N_1785,N_1730);
nand U1805 (N_1805,N_1790,N_1789);
nor U1806 (N_1806,N_1721,N_1744);
and U1807 (N_1807,N_1747,N_1726);
nand U1808 (N_1808,N_1759,N_1749);
and U1809 (N_1809,N_1719,N_1776);
nand U1810 (N_1810,N_1797,N_1716);
nor U1811 (N_1811,N_1717,N_1718);
and U1812 (N_1812,N_1722,N_1782);
and U1813 (N_1813,N_1798,N_1771);
nand U1814 (N_1814,N_1724,N_1769);
nor U1815 (N_1815,N_1703,N_1714);
or U1816 (N_1816,N_1702,N_1786);
and U1817 (N_1817,N_1710,N_1791);
xnor U1818 (N_1818,N_1732,N_1755);
xnor U1819 (N_1819,N_1793,N_1745);
or U1820 (N_1820,N_1767,N_1757);
nor U1821 (N_1821,N_1752,N_1788);
nor U1822 (N_1822,N_1762,N_1725);
nor U1823 (N_1823,N_1779,N_1763);
nand U1824 (N_1824,N_1746,N_1795);
and U1825 (N_1825,N_1792,N_1758);
or U1826 (N_1826,N_1766,N_1743);
nor U1827 (N_1827,N_1741,N_1713);
or U1828 (N_1828,N_1708,N_1709);
nand U1829 (N_1829,N_1742,N_1735);
nor U1830 (N_1830,N_1715,N_1728);
nand U1831 (N_1831,N_1729,N_1773);
and U1832 (N_1832,N_1796,N_1707);
and U1833 (N_1833,N_1783,N_1761);
and U1834 (N_1834,N_1737,N_1727);
nand U1835 (N_1835,N_1768,N_1784);
and U1836 (N_1836,N_1739,N_1700);
or U1837 (N_1837,N_1781,N_1774);
nor U1838 (N_1838,N_1753,N_1778);
nand U1839 (N_1839,N_1765,N_1760);
nor U1840 (N_1840,N_1780,N_1756);
nor U1841 (N_1841,N_1701,N_1736);
and U1842 (N_1842,N_1734,N_1750);
nor U1843 (N_1843,N_1777,N_1711);
nor U1844 (N_1844,N_1748,N_1705);
nor U1845 (N_1845,N_1787,N_1706);
and U1846 (N_1846,N_1794,N_1764);
nand U1847 (N_1847,N_1770,N_1751);
xnor U1848 (N_1848,N_1733,N_1720);
nand U1849 (N_1849,N_1775,N_1731);
and U1850 (N_1850,N_1759,N_1710);
nand U1851 (N_1851,N_1749,N_1788);
xnor U1852 (N_1852,N_1706,N_1782);
and U1853 (N_1853,N_1796,N_1776);
and U1854 (N_1854,N_1729,N_1750);
nor U1855 (N_1855,N_1719,N_1795);
xor U1856 (N_1856,N_1793,N_1711);
xnor U1857 (N_1857,N_1719,N_1752);
nand U1858 (N_1858,N_1739,N_1732);
or U1859 (N_1859,N_1761,N_1784);
nor U1860 (N_1860,N_1705,N_1704);
nand U1861 (N_1861,N_1711,N_1773);
nor U1862 (N_1862,N_1717,N_1745);
nand U1863 (N_1863,N_1727,N_1763);
nor U1864 (N_1864,N_1710,N_1726);
nand U1865 (N_1865,N_1749,N_1762);
and U1866 (N_1866,N_1754,N_1793);
or U1867 (N_1867,N_1771,N_1708);
nand U1868 (N_1868,N_1756,N_1760);
nor U1869 (N_1869,N_1780,N_1707);
or U1870 (N_1870,N_1733,N_1751);
nand U1871 (N_1871,N_1796,N_1751);
nor U1872 (N_1872,N_1731,N_1750);
nor U1873 (N_1873,N_1782,N_1756);
nor U1874 (N_1874,N_1782,N_1783);
nor U1875 (N_1875,N_1752,N_1750);
or U1876 (N_1876,N_1705,N_1796);
or U1877 (N_1877,N_1792,N_1784);
and U1878 (N_1878,N_1723,N_1769);
nor U1879 (N_1879,N_1709,N_1763);
xnor U1880 (N_1880,N_1791,N_1777);
nor U1881 (N_1881,N_1711,N_1768);
or U1882 (N_1882,N_1725,N_1738);
or U1883 (N_1883,N_1704,N_1730);
or U1884 (N_1884,N_1701,N_1747);
nand U1885 (N_1885,N_1770,N_1742);
or U1886 (N_1886,N_1709,N_1793);
nand U1887 (N_1887,N_1749,N_1764);
nor U1888 (N_1888,N_1764,N_1755);
and U1889 (N_1889,N_1710,N_1717);
nor U1890 (N_1890,N_1704,N_1747);
and U1891 (N_1891,N_1704,N_1792);
or U1892 (N_1892,N_1727,N_1760);
nand U1893 (N_1893,N_1770,N_1716);
nand U1894 (N_1894,N_1765,N_1725);
nand U1895 (N_1895,N_1701,N_1733);
xnor U1896 (N_1896,N_1780,N_1732);
and U1897 (N_1897,N_1731,N_1776);
nor U1898 (N_1898,N_1715,N_1795);
nor U1899 (N_1899,N_1771,N_1791);
xnor U1900 (N_1900,N_1844,N_1866);
and U1901 (N_1901,N_1896,N_1857);
and U1902 (N_1902,N_1819,N_1875);
nand U1903 (N_1903,N_1852,N_1889);
nor U1904 (N_1904,N_1862,N_1861);
or U1905 (N_1905,N_1895,N_1810);
nand U1906 (N_1906,N_1884,N_1848);
nor U1907 (N_1907,N_1877,N_1878);
and U1908 (N_1908,N_1841,N_1855);
and U1909 (N_1909,N_1820,N_1859);
nor U1910 (N_1910,N_1879,N_1829);
xnor U1911 (N_1911,N_1802,N_1803);
nor U1912 (N_1912,N_1850,N_1863);
nor U1913 (N_1913,N_1860,N_1835);
nor U1914 (N_1914,N_1864,N_1887);
xor U1915 (N_1915,N_1833,N_1826);
nand U1916 (N_1916,N_1899,N_1886);
and U1917 (N_1917,N_1842,N_1806);
nor U1918 (N_1918,N_1873,N_1897);
nor U1919 (N_1919,N_1871,N_1815);
nor U1920 (N_1920,N_1839,N_1830);
or U1921 (N_1921,N_1812,N_1832);
or U1922 (N_1922,N_1880,N_1813);
nand U1923 (N_1923,N_1872,N_1885);
nor U1924 (N_1924,N_1828,N_1838);
xor U1925 (N_1925,N_1808,N_1814);
or U1926 (N_1926,N_1869,N_1854);
nand U1927 (N_1927,N_1865,N_1804);
nor U1928 (N_1928,N_1823,N_1892);
and U1929 (N_1929,N_1822,N_1811);
xor U1930 (N_1930,N_1818,N_1868);
nor U1931 (N_1931,N_1893,N_1816);
or U1932 (N_1932,N_1824,N_1853);
nand U1933 (N_1933,N_1840,N_1870);
nor U1934 (N_1934,N_1874,N_1834);
nand U1935 (N_1935,N_1894,N_1836);
and U1936 (N_1936,N_1817,N_1881);
or U1937 (N_1937,N_1867,N_1856);
nand U1938 (N_1938,N_1849,N_1845);
nor U1939 (N_1939,N_1888,N_1851);
nor U1940 (N_1940,N_1898,N_1846);
nor U1941 (N_1941,N_1825,N_1843);
or U1942 (N_1942,N_1809,N_1831);
nor U1943 (N_1943,N_1805,N_1827);
nand U1944 (N_1944,N_1800,N_1847);
nand U1945 (N_1945,N_1890,N_1876);
or U1946 (N_1946,N_1891,N_1821);
nor U1947 (N_1947,N_1807,N_1801);
nor U1948 (N_1948,N_1837,N_1883);
xnor U1949 (N_1949,N_1882,N_1858);
nand U1950 (N_1950,N_1840,N_1830);
or U1951 (N_1951,N_1874,N_1899);
nand U1952 (N_1952,N_1849,N_1808);
xor U1953 (N_1953,N_1894,N_1877);
nand U1954 (N_1954,N_1898,N_1815);
xnor U1955 (N_1955,N_1859,N_1845);
nand U1956 (N_1956,N_1821,N_1887);
or U1957 (N_1957,N_1822,N_1858);
nor U1958 (N_1958,N_1891,N_1823);
nor U1959 (N_1959,N_1844,N_1890);
or U1960 (N_1960,N_1885,N_1887);
xor U1961 (N_1961,N_1869,N_1882);
nand U1962 (N_1962,N_1867,N_1894);
nand U1963 (N_1963,N_1845,N_1897);
or U1964 (N_1964,N_1841,N_1833);
or U1965 (N_1965,N_1835,N_1808);
or U1966 (N_1966,N_1873,N_1887);
or U1967 (N_1967,N_1890,N_1858);
or U1968 (N_1968,N_1891,N_1839);
and U1969 (N_1969,N_1816,N_1857);
xnor U1970 (N_1970,N_1805,N_1863);
and U1971 (N_1971,N_1891,N_1842);
nand U1972 (N_1972,N_1874,N_1804);
and U1973 (N_1973,N_1877,N_1830);
or U1974 (N_1974,N_1831,N_1824);
xnor U1975 (N_1975,N_1812,N_1852);
nand U1976 (N_1976,N_1847,N_1868);
or U1977 (N_1977,N_1828,N_1850);
nand U1978 (N_1978,N_1885,N_1836);
nor U1979 (N_1979,N_1828,N_1821);
nand U1980 (N_1980,N_1894,N_1860);
nand U1981 (N_1981,N_1858,N_1877);
xor U1982 (N_1982,N_1891,N_1831);
or U1983 (N_1983,N_1851,N_1871);
and U1984 (N_1984,N_1849,N_1841);
or U1985 (N_1985,N_1855,N_1890);
nand U1986 (N_1986,N_1802,N_1816);
nand U1987 (N_1987,N_1893,N_1852);
nor U1988 (N_1988,N_1801,N_1852);
nor U1989 (N_1989,N_1827,N_1849);
nand U1990 (N_1990,N_1883,N_1862);
nor U1991 (N_1991,N_1873,N_1884);
or U1992 (N_1992,N_1865,N_1817);
and U1993 (N_1993,N_1843,N_1806);
or U1994 (N_1994,N_1818,N_1852);
nor U1995 (N_1995,N_1885,N_1846);
and U1996 (N_1996,N_1869,N_1867);
nor U1997 (N_1997,N_1844,N_1808);
and U1998 (N_1998,N_1830,N_1873);
nor U1999 (N_1999,N_1898,N_1849);
and U2000 (N_2000,N_1951,N_1908);
nand U2001 (N_2001,N_1924,N_1937);
and U2002 (N_2002,N_1910,N_1950);
and U2003 (N_2003,N_1994,N_1912);
nand U2004 (N_2004,N_1992,N_1962);
nor U2005 (N_2005,N_1943,N_1961);
or U2006 (N_2006,N_1972,N_1927);
nor U2007 (N_2007,N_1959,N_1925);
xnor U2008 (N_2008,N_1918,N_1963);
or U2009 (N_2009,N_1979,N_1958);
nand U2010 (N_2010,N_1967,N_1960);
nor U2011 (N_2011,N_1901,N_1933);
xnor U2012 (N_2012,N_1942,N_1936);
and U2013 (N_2013,N_1983,N_1929);
nand U2014 (N_2014,N_1965,N_1909);
xnor U2015 (N_2015,N_1903,N_1939);
and U2016 (N_2016,N_1984,N_1982);
or U2017 (N_2017,N_1921,N_1911);
and U2018 (N_2018,N_1949,N_1906);
xor U2019 (N_2019,N_1941,N_1934);
or U2020 (N_2020,N_1986,N_1914);
or U2021 (N_2021,N_1902,N_1953);
nor U2022 (N_2022,N_1900,N_1969);
nor U2023 (N_2023,N_1976,N_1947);
nand U2024 (N_2024,N_1916,N_1997);
nand U2025 (N_2025,N_1985,N_1931);
nand U2026 (N_2026,N_1930,N_1991);
nor U2027 (N_2027,N_1964,N_1940);
nand U2028 (N_2028,N_1957,N_1974);
and U2029 (N_2029,N_1996,N_1988);
or U2030 (N_2030,N_1920,N_1932);
nand U2031 (N_2031,N_1975,N_1995);
and U2032 (N_2032,N_1999,N_1990);
and U2033 (N_2033,N_1955,N_1954);
and U2034 (N_2034,N_1907,N_1993);
and U2035 (N_2035,N_1980,N_1948);
nor U2036 (N_2036,N_1989,N_1915);
and U2037 (N_2037,N_1923,N_1904);
xnor U2038 (N_2038,N_1926,N_1977);
nand U2039 (N_2039,N_1919,N_1956);
nor U2040 (N_2040,N_1968,N_1913);
nor U2041 (N_2041,N_1973,N_1987);
or U2042 (N_2042,N_1917,N_1970);
nor U2043 (N_2043,N_1922,N_1998);
or U2044 (N_2044,N_1945,N_1952);
or U2045 (N_2045,N_1966,N_1944);
and U2046 (N_2046,N_1981,N_1928);
nand U2047 (N_2047,N_1946,N_1971);
nor U2048 (N_2048,N_1905,N_1938);
or U2049 (N_2049,N_1935,N_1978);
or U2050 (N_2050,N_1971,N_1922);
nand U2051 (N_2051,N_1949,N_1994);
nor U2052 (N_2052,N_1959,N_1932);
xor U2053 (N_2053,N_1988,N_1926);
nand U2054 (N_2054,N_1958,N_1905);
nand U2055 (N_2055,N_1924,N_1923);
and U2056 (N_2056,N_1991,N_1978);
nand U2057 (N_2057,N_1970,N_1903);
or U2058 (N_2058,N_1968,N_1966);
nor U2059 (N_2059,N_1990,N_1970);
xnor U2060 (N_2060,N_1902,N_1926);
nand U2061 (N_2061,N_1999,N_1945);
nand U2062 (N_2062,N_1938,N_1915);
xnor U2063 (N_2063,N_1965,N_1935);
or U2064 (N_2064,N_1932,N_1964);
nand U2065 (N_2065,N_1968,N_1975);
and U2066 (N_2066,N_1930,N_1927);
and U2067 (N_2067,N_1908,N_1922);
or U2068 (N_2068,N_1988,N_1937);
nand U2069 (N_2069,N_1949,N_1917);
nor U2070 (N_2070,N_1974,N_1904);
and U2071 (N_2071,N_1988,N_1920);
or U2072 (N_2072,N_1988,N_1989);
nand U2073 (N_2073,N_1922,N_1952);
nand U2074 (N_2074,N_1984,N_1901);
nor U2075 (N_2075,N_1964,N_1970);
nor U2076 (N_2076,N_1912,N_1902);
or U2077 (N_2077,N_1933,N_1979);
nor U2078 (N_2078,N_1904,N_1985);
and U2079 (N_2079,N_1968,N_1992);
and U2080 (N_2080,N_1924,N_1933);
nor U2081 (N_2081,N_1967,N_1934);
nand U2082 (N_2082,N_1966,N_1916);
nor U2083 (N_2083,N_1906,N_1987);
or U2084 (N_2084,N_1963,N_1911);
nor U2085 (N_2085,N_1937,N_1932);
nor U2086 (N_2086,N_1913,N_1991);
xor U2087 (N_2087,N_1971,N_1992);
nand U2088 (N_2088,N_1910,N_1921);
nor U2089 (N_2089,N_1916,N_1961);
nand U2090 (N_2090,N_1970,N_1934);
nor U2091 (N_2091,N_1970,N_1908);
or U2092 (N_2092,N_1968,N_1945);
nor U2093 (N_2093,N_1930,N_1905);
or U2094 (N_2094,N_1957,N_1938);
nand U2095 (N_2095,N_1980,N_1934);
nor U2096 (N_2096,N_1902,N_1919);
nand U2097 (N_2097,N_1943,N_1909);
xor U2098 (N_2098,N_1946,N_1930);
nand U2099 (N_2099,N_1935,N_1971);
and U2100 (N_2100,N_2050,N_2083);
or U2101 (N_2101,N_2017,N_2013);
nor U2102 (N_2102,N_2021,N_2028);
or U2103 (N_2103,N_2027,N_2046);
or U2104 (N_2104,N_2029,N_2000);
or U2105 (N_2105,N_2052,N_2063);
nand U2106 (N_2106,N_2019,N_2067);
nor U2107 (N_2107,N_2047,N_2071);
and U2108 (N_2108,N_2082,N_2089);
xor U2109 (N_2109,N_2056,N_2051);
and U2110 (N_2110,N_2045,N_2044);
and U2111 (N_2111,N_2031,N_2015);
nor U2112 (N_2112,N_2001,N_2042);
or U2113 (N_2113,N_2005,N_2043);
nand U2114 (N_2114,N_2049,N_2020);
nor U2115 (N_2115,N_2087,N_2084);
and U2116 (N_2116,N_2034,N_2072);
and U2117 (N_2117,N_2026,N_2039);
nand U2118 (N_2118,N_2095,N_2010);
nor U2119 (N_2119,N_2097,N_2036);
or U2120 (N_2120,N_2090,N_2003);
xnor U2121 (N_2121,N_2041,N_2030);
nor U2122 (N_2122,N_2055,N_2061);
nand U2123 (N_2123,N_2091,N_2088);
nor U2124 (N_2124,N_2085,N_2033);
or U2125 (N_2125,N_2011,N_2023);
or U2126 (N_2126,N_2040,N_2057);
nand U2127 (N_2127,N_2062,N_2032);
and U2128 (N_2128,N_2025,N_2096);
and U2129 (N_2129,N_2009,N_2073);
xor U2130 (N_2130,N_2099,N_2075);
xor U2131 (N_2131,N_2064,N_2092);
nand U2132 (N_2132,N_2094,N_2074);
or U2133 (N_2133,N_2086,N_2078);
nor U2134 (N_2134,N_2007,N_2002);
and U2135 (N_2135,N_2016,N_2014);
or U2136 (N_2136,N_2022,N_2024);
or U2137 (N_2137,N_2069,N_2066);
nand U2138 (N_2138,N_2076,N_2018);
and U2139 (N_2139,N_2012,N_2068);
or U2140 (N_2140,N_2070,N_2077);
and U2141 (N_2141,N_2008,N_2004);
nand U2142 (N_2142,N_2037,N_2038);
nor U2143 (N_2143,N_2035,N_2058);
nor U2144 (N_2144,N_2053,N_2079);
xor U2145 (N_2145,N_2065,N_2054);
or U2146 (N_2146,N_2048,N_2081);
xor U2147 (N_2147,N_2080,N_2093);
nor U2148 (N_2148,N_2098,N_2060);
nand U2149 (N_2149,N_2059,N_2006);
nand U2150 (N_2150,N_2072,N_2049);
nand U2151 (N_2151,N_2019,N_2080);
and U2152 (N_2152,N_2054,N_2074);
nand U2153 (N_2153,N_2094,N_2082);
nand U2154 (N_2154,N_2056,N_2044);
or U2155 (N_2155,N_2046,N_2031);
nor U2156 (N_2156,N_2082,N_2036);
and U2157 (N_2157,N_2095,N_2045);
and U2158 (N_2158,N_2052,N_2021);
or U2159 (N_2159,N_2043,N_2056);
or U2160 (N_2160,N_2022,N_2001);
or U2161 (N_2161,N_2048,N_2067);
nand U2162 (N_2162,N_2041,N_2052);
nand U2163 (N_2163,N_2076,N_2014);
and U2164 (N_2164,N_2067,N_2097);
nand U2165 (N_2165,N_2060,N_2062);
or U2166 (N_2166,N_2004,N_2050);
nand U2167 (N_2167,N_2001,N_2068);
nor U2168 (N_2168,N_2088,N_2045);
nor U2169 (N_2169,N_2048,N_2035);
nand U2170 (N_2170,N_2049,N_2058);
or U2171 (N_2171,N_2076,N_2049);
or U2172 (N_2172,N_2019,N_2085);
nor U2173 (N_2173,N_2039,N_2087);
or U2174 (N_2174,N_2031,N_2065);
nor U2175 (N_2175,N_2043,N_2037);
nand U2176 (N_2176,N_2030,N_2058);
xnor U2177 (N_2177,N_2097,N_2077);
nor U2178 (N_2178,N_2054,N_2008);
nor U2179 (N_2179,N_2035,N_2055);
or U2180 (N_2180,N_2035,N_2057);
or U2181 (N_2181,N_2006,N_2073);
nor U2182 (N_2182,N_2013,N_2060);
nor U2183 (N_2183,N_2068,N_2000);
or U2184 (N_2184,N_2045,N_2009);
and U2185 (N_2185,N_2042,N_2068);
nor U2186 (N_2186,N_2034,N_2080);
and U2187 (N_2187,N_2071,N_2059);
xor U2188 (N_2188,N_2014,N_2054);
and U2189 (N_2189,N_2038,N_2000);
nand U2190 (N_2190,N_2004,N_2096);
nand U2191 (N_2191,N_2056,N_2099);
nand U2192 (N_2192,N_2026,N_2088);
nand U2193 (N_2193,N_2017,N_2067);
or U2194 (N_2194,N_2039,N_2088);
or U2195 (N_2195,N_2021,N_2054);
nor U2196 (N_2196,N_2089,N_2069);
nor U2197 (N_2197,N_2009,N_2060);
nand U2198 (N_2198,N_2044,N_2003);
or U2199 (N_2199,N_2096,N_2012);
nand U2200 (N_2200,N_2156,N_2112);
nand U2201 (N_2201,N_2100,N_2150);
xnor U2202 (N_2202,N_2120,N_2108);
nor U2203 (N_2203,N_2144,N_2193);
or U2204 (N_2204,N_2178,N_2118);
nand U2205 (N_2205,N_2151,N_2181);
nand U2206 (N_2206,N_2106,N_2113);
and U2207 (N_2207,N_2117,N_2190);
nand U2208 (N_2208,N_2132,N_2173);
and U2209 (N_2209,N_2195,N_2154);
nand U2210 (N_2210,N_2184,N_2111);
and U2211 (N_2211,N_2128,N_2105);
nand U2212 (N_2212,N_2170,N_2115);
nand U2213 (N_2213,N_2186,N_2142);
nand U2214 (N_2214,N_2175,N_2185);
nand U2215 (N_2215,N_2152,N_2189);
and U2216 (N_2216,N_2194,N_2109);
or U2217 (N_2217,N_2139,N_2119);
or U2218 (N_2218,N_2183,N_2161);
nor U2219 (N_2219,N_2179,N_2135);
nand U2220 (N_2220,N_2133,N_2131);
or U2221 (N_2221,N_2104,N_2188);
and U2222 (N_2222,N_2162,N_2155);
and U2223 (N_2223,N_2147,N_2101);
nor U2224 (N_2224,N_2199,N_2180);
nor U2225 (N_2225,N_2143,N_2127);
nand U2226 (N_2226,N_2102,N_2168);
and U2227 (N_2227,N_2149,N_2174);
or U2228 (N_2228,N_2167,N_2157);
xnor U2229 (N_2229,N_2197,N_2125);
nor U2230 (N_2230,N_2176,N_2148);
or U2231 (N_2231,N_2134,N_2166);
and U2232 (N_2232,N_2163,N_2196);
nor U2233 (N_2233,N_2141,N_2191);
nand U2234 (N_2234,N_2130,N_2164);
nand U2235 (N_2235,N_2182,N_2171);
nor U2236 (N_2236,N_2138,N_2169);
and U2237 (N_2237,N_2158,N_2126);
nor U2238 (N_2238,N_2124,N_2198);
and U2239 (N_2239,N_2122,N_2107);
nor U2240 (N_2240,N_2123,N_2145);
nand U2241 (N_2241,N_2140,N_2129);
nor U2242 (N_2242,N_2165,N_2137);
nand U2243 (N_2243,N_2172,N_2116);
or U2244 (N_2244,N_2159,N_2187);
and U2245 (N_2245,N_2160,N_2146);
or U2246 (N_2246,N_2103,N_2110);
and U2247 (N_2247,N_2136,N_2121);
and U2248 (N_2248,N_2114,N_2192);
nand U2249 (N_2249,N_2153,N_2177);
nand U2250 (N_2250,N_2194,N_2127);
nor U2251 (N_2251,N_2126,N_2169);
or U2252 (N_2252,N_2158,N_2187);
and U2253 (N_2253,N_2188,N_2184);
nor U2254 (N_2254,N_2178,N_2176);
or U2255 (N_2255,N_2103,N_2171);
and U2256 (N_2256,N_2183,N_2149);
or U2257 (N_2257,N_2172,N_2178);
nor U2258 (N_2258,N_2198,N_2145);
nor U2259 (N_2259,N_2122,N_2154);
xnor U2260 (N_2260,N_2169,N_2192);
nand U2261 (N_2261,N_2124,N_2157);
xor U2262 (N_2262,N_2103,N_2101);
nor U2263 (N_2263,N_2170,N_2100);
and U2264 (N_2264,N_2147,N_2179);
or U2265 (N_2265,N_2199,N_2171);
or U2266 (N_2266,N_2160,N_2152);
and U2267 (N_2267,N_2110,N_2188);
and U2268 (N_2268,N_2184,N_2161);
or U2269 (N_2269,N_2190,N_2151);
nor U2270 (N_2270,N_2109,N_2139);
nor U2271 (N_2271,N_2118,N_2167);
and U2272 (N_2272,N_2148,N_2154);
or U2273 (N_2273,N_2145,N_2146);
nor U2274 (N_2274,N_2115,N_2149);
xnor U2275 (N_2275,N_2170,N_2166);
and U2276 (N_2276,N_2150,N_2141);
or U2277 (N_2277,N_2179,N_2146);
and U2278 (N_2278,N_2104,N_2127);
and U2279 (N_2279,N_2140,N_2152);
nand U2280 (N_2280,N_2175,N_2152);
nand U2281 (N_2281,N_2106,N_2140);
or U2282 (N_2282,N_2171,N_2120);
nand U2283 (N_2283,N_2183,N_2103);
and U2284 (N_2284,N_2130,N_2179);
and U2285 (N_2285,N_2172,N_2142);
or U2286 (N_2286,N_2105,N_2103);
nor U2287 (N_2287,N_2138,N_2125);
or U2288 (N_2288,N_2188,N_2114);
nor U2289 (N_2289,N_2114,N_2191);
and U2290 (N_2290,N_2155,N_2159);
and U2291 (N_2291,N_2135,N_2185);
nor U2292 (N_2292,N_2150,N_2169);
or U2293 (N_2293,N_2191,N_2157);
and U2294 (N_2294,N_2152,N_2124);
and U2295 (N_2295,N_2178,N_2123);
and U2296 (N_2296,N_2105,N_2113);
and U2297 (N_2297,N_2183,N_2187);
nand U2298 (N_2298,N_2148,N_2193);
and U2299 (N_2299,N_2194,N_2178);
or U2300 (N_2300,N_2216,N_2201);
nor U2301 (N_2301,N_2236,N_2280);
nor U2302 (N_2302,N_2239,N_2262);
nor U2303 (N_2303,N_2267,N_2257);
nor U2304 (N_2304,N_2221,N_2291);
or U2305 (N_2305,N_2242,N_2223);
and U2306 (N_2306,N_2283,N_2226);
and U2307 (N_2307,N_2234,N_2218);
nand U2308 (N_2308,N_2214,N_2251);
nor U2309 (N_2309,N_2230,N_2274);
xnor U2310 (N_2310,N_2287,N_2224);
and U2311 (N_2311,N_2246,N_2206);
nor U2312 (N_2312,N_2219,N_2277);
xor U2313 (N_2313,N_2215,N_2241);
or U2314 (N_2314,N_2293,N_2253);
nor U2315 (N_2315,N_2205,N_2232);
or U2316 (N_2316,N_2258,N_2254);
or U2317 (N_2317,N_2247,N_2259);
and U2318 (N_2318,N_2252,N_2288);
nand U2319 (N_2319,N_2229,N_2281);
nor U2320 (N_2320,N_2243,N_2260);
nand U2321 (N_2321,N_2240,N_2231);
xor U2322 (N_2322,N_2228,N_2220);
and U2323 (N_2323,N_2269,N_2217);
or U2324 (N_2324,N_2296,N_2208);
nor U2325 (N_2325,N_2282,N_2211);
and U2326 (N_2326,N_2285,N_2248);
nor U2327 (N_2327,N_2298,N_2290);
and U2328 (N_2328,N_2202,N_2286);
nand U2329 (N_2329,N_2266,N_2271);
nand U2330 (N_2330,N_2244,N_2204);
or U2331 (N_2331,N_2272,N_2225);
and U2332 (N_2332,N_2263,N_2207);
nand U2333 (N_2333,N_2273,N_2203);
or U2334 (N_2334,N_2297,N_2245);
nand U2335 (N_2335,N_2255,N_2249);
and U2336 (N_2336,N_2222,N_2250);
or U2337 (N_2337,N_2276,N_2299);
or U2338 (N_2338,N_2237,N_2233);
xor U2339 (N_2339,N_2289,N_2209);
nand U2340 (N_2340,N_2210,N_2227);
nor U2341 (N_2341,N_2279,N_2295);
nand U2342 (N_2342,N_2294,N_2235);
or U2343 (N_2343,N_2261,N_2275);
and U2344 (N_2344,N_2284,N_2256);
nor U2345 (N_2345,N_2278,N_2292);
nor U2346 (N_2346,N_2270,N_2200);
nand U2347 (N_2347,N_2268,N_2238);
and U2348 (N_2348,N_2213,N_2264);
nor U2349 (N_2349,N_2265,N_2212);
nor U2350 (N_2350,N_2298,N_2297);
nor U2351 (N_2351,N_2280,N_2241);
and U2352 (N_2352,N_2217,N_2219);
nand U2353 (N_2353,N_2259,N_2294);
xor U2354 (N_2354,N_2229,N_2268);
and U2355 (N_2355,N_2247,N_2272);
or U2356 (N_2356,N_2203,N_2244);
or U2357 (N_2357,N_2231,N_2224);
nor U2358 (N_2358,N_2223,N_2227);
or U2359 (N_2359,N_2200,N_2232);
and U2360 (N_2360,N_2299,N_2255);
nand U2361 (N_2361,N_2202,N_2297);
nand U2362 (N_2362,N_2252,N_2267);
or U2363 (N_2363,N_2219,N_2261);
nand U2364 (N_2364,N_2264,N_2224);
nand U2365 (N_2365,N_2282,N_2288);
or U2366 (N_2366,N_2238,N_2269);
and U2367 (N_2367,N_2258,N_2218);
nor U2368 (N_2368,N_2231,N_2203);
nand U2369 (N_2369,N_2206,N_2253);
nor U2370 (N_2370,N_2230,N_2251);
xnor U2371 (N_2371,N_2242,N_2237);
nor U2372 (N_2372,N_2295,N_2232);
and U2373 (N_2373,N_2292,N_2227);
nor U2374 (N_2374,N_2215,N_2226);
and U2375 (N_2375,N_2245,N_2244);
or U2376 (N_2376,N_2236,N_2271);
nor U2377 (N_2377,N_2236,N_2275);
nor U2378 (N_2378,N_2213,N_2237);
or U2379 (N_2379,N_2260,N_2297);
nor U2380 (N_2380,N_2219,N_2253);
xor U2381 (N_2381,N_2243,N_2240);
nor U2382 (N_2382,N_2297,N_2209);
nor U2383 (N_2383,N_2204,N_2207);
and U2384 (N_2384,N_2281,N_2219);
and U2385 (N_2385,N_2279,N_2215);
and U2386 (N_2386,N_2277,N_2209);
and U2387 (N_2387,N_2260,N_2284);
nor U2388 (N_2388,N_2273,N_2216);
nand U2389 (N_2389,N_2229,N_2299);
or U2390 (N_2390,N_2261,N_2218);
and U2391 (N_2391,N_2222,N_2288);
and U2392 (N_2392,N_2208,N_2217);
nor U2393 (N_2393,N_2234,N_2224);
nor U2394 (N_2394,N_2282,N_2273);
xnor U2395 (N_2395,N_2269,N_2235);
and U2396 (N_2396,N_2223,N_2245);
nor U2397 (N_2397,N_2223,N_2257);
xnor U2398 (N_2398,N_2272,N_2245);
nor U2399 (N_2399,N_2209,N_2284);
nor U2400 (N_2400,N_2309,N_2357);
nor U2401 (N_2401,N_2358,N_2303);
and U2402 (N_2402,N_2305,N_2343);
nand U2403 (N_2403,N_2362,N_2327);
nor U2404 (N_2404,N_2321,N_2314);
and U2405 (N_2405,N_2366,N_2352);
or U2406 (N_2406,N_2351,N_2398);
xor U2407 (N_2407,N_2323,N_2374);
and U2408 (N_2408,N_2349,N_2350);
or U2409 (N_2409,N_2337,N_2342);
xnor U2410 (N_2410,N_2382,N_2375);
nand U2411 (N_2411,N_2384,N_2301);
nor U2412 (N_2412,N_2359,N_2322);
and U2413 (N_2413,N_2361,N_2364);
or U2414 (N_2414,N_2387,N_2373);
nand U2415 (N_2415,N_2397,N_2346);
and U2416 (N_2416,N_2334,N_2307);
or U2417 (N_2417,N_2336,N_2365);
nand U2418 (N_2418,N_2344,N_2345);
nand U2419 (N_2419,N_2329,N_2339);
and U2420 (N_2420,N_2385,N_2390);
xnor U2421 (N_2421,N_2325,N_2311);
or U2422 (N_2422,N_2308,N_2340);
and U2423 (N_2423,N_2396,N_2391);
xnor U2424 (N_2424,N_2381,N_2395);
nor U2425 (N_2425,N_2317,N_2312);
and U2426 (N_2426,N_2328,N_2367);
and U2427 (N_2427,N_2306,N_2335);
xnor U2428 (N_2428,N_2333,N_2371);
nand U2429 (N_2429,N_2353,N_2310);
and U2430 (N_2430,N_2326,N_2360);
nor U2431 (N_2431,N_2348,N_2369);
nand U2432 (N_2432,N_2399,N_2332);
and U2433 (N_2433,N_2363,N_2372);
nand U2434 (N_2434,N_2378,N_2315);
xor U2435 (N_2435,N_2379,N_2354);
nor U2436 (N_2436,N_2355,N_2313);
and U2437 (N_2437,N_2304,N_2300);
nand U2438 (N_2438,N_2383,N_2388);
nor U2439 (N_2439,N_2392,N_2347);
and U2440 (N_2440,N_2389,N_2376);
or U2441 (N_2441,N_2302,N_2386);
nand U2442 (N_2442,N_2393,N_2331);
nor U2443 (N_2443,N_2380,N_2341);
nor U2444 (N_2444,N_2324,N_2377);
or U2445 (N_2445,N_2330,N_2318);
nand U2446 (N_2446,N_2338,N_2370);
xor U2447 (N_2447,N_2394,N_2319);
xor U2448 (N_2448,N_2368,N_2320);
nor U2449 (N_2449,N_2356,N_2316);
nor U2450 (N_2450,N_2309,N_2317);
nor U2451 (N_2451,N_2382,N_2327);
nand U2452 (N_2452,N_2353,N_2397);
or U2453 (N_2453,N_2320,N_2399);
nor U2454 (N_2454,N_2397,N_2340);
nand U2455 (N_2455,N_2349,N_2322);
xor U2456 (N_2456,N_2389,N_2345);
nand U2457 (N_2457,N_2304,N_2315);
and U2458 (N_2458,N_2309,N_2324);
or U2459 (N_2459,N_2354,N_2341);
nand U2460 (N_2460,N_2388,N_2333);
or U2461 (N_2461,N_2397,N_2375);
nor U2462 (N_2462,N_2301,N_2389);
and U2463 (N_2463,N_2300,N_2342);
nor U2464 (N_2464,N_2386,N_2306);
or U2465 (N_2465,N_2349,N_2315);
and U2466 (N_2466,N_2376,N_2398);
or U2467 (N_2467,N_2361,N_2399);
or U2468 (N_2468,N_2398,N_2378);
nand U2469 (N_2469,N_2376,N_2367);
and U2470 (N_2470,N_2321,N_2385);
and U2471 (N_2471,N_2315,N_2323);
nand U2472 (N_2472,N_2369,N_2330);
nor U2473 (N_2473,N_2381,N_2343);
nor U2474 (N_2474,N_2352,N_2314);
nand U2475 (N_2475,N_2322,N_2328);
and U2476 (N_2476,N_2307,N_2364);
or U2477 (N_2477,N_2300,N_2318);
or U2478 (N_2478,N_2382,N_2321);
or U2479 (N_2479,N_2329,N_2340);
nor U2480 (N_2480,N_2322,N_2324);
nand U2481 (N_2481,N_2351,N_2308);
or U2482 (N_2482,N_2338,N_2302);
and U2483 (N_2483,N_2399,N_2366);
nor U2484 (N_2484,N_2397,N_2380);
nor U2485 (N_2485,N_2391,N_2382);
nand U2486 (N_2486,N_2362,N_2300);
nor U2487 (N_2487,N_2323,N_2301);
xnor U2488 (N_2488,N_2340,N_2374);
nand U2489 (N_2489,N_2381,N_2321);
nor U2490 (N_2490,N_2345,N_2387);
nand U2491 (N_2491,N_2346,N_2304);
nand U2492 (N_2492,N_2327,N_2328);
nand U2493 (N_2493,N_2330,N_2364);
or U2494 (N_2494,N_2311,N_2361);
and U2495 (N_2495,N_2321,N_2308);
or U2496 (N_2496,N_2333,N_2350);
and U2497 (N_2497,N_2381,N_2306);
xnor U2498 (N_2498,N_2333,N_2356);
or U2499 (N_2499,N_2380,N_2332);
or U2500 (N_2500,N_2452,N_2483);
and U2501 (N_2501,N_2437,N_2499);
xor U2502 (N_2502,N_2433,N_2418);
nor U2503 (N_2503,N_2479,N_2486);
xnor U2504 (N_2504,N_2490,N_2495);
nor U2505 (N_2505,N_2407,N_2492);
nor U2506 (N_2506,N_2435,N_2493);
or U2507 (N_2507,N_2417,N_2482);
nor U2508 (N_2508,N_2453,N_2462);
nand U2509 (N_2509,N_2405,N_2401);
nor U2510 (N_2510,N_2467,N_2432);
nor U2511 (N_2511,N_2446,N_2455);
nand U2512 (N_2512,N_2445,N_2429);
or U2513 (N_2513,N_2458,N_2466);
or U2514 (N_2514,N_2424,N_2464);
and U2515 (N_2515,N_2443,N_2472);
or U2516 (N_2516,N_2402,N_2470);
and U2517 (N_2517,N_2409,N_2403);
nor U2518 (N_2518,N_2463,N_2439);
nor U2519 (N_2519,N_2461,N_2496);
nand U2520 (N_2520,N_2469,N_2430);
or U2521 (N_2521,N_2428,N_2431);
or U2522 (N_2522,N_2487,N_2471);
or U2523 (N_2523,N_2425,N_2412);
xnor U2524 (N_2524,N_2416,N_2475);
nor U2525 (N_2525,N_2449,N_2448);
nand U2526 (N_2526,N_2426,N_2415);
or U2527 (N_2527,N_2423,N_2460);
and U2528 (N_2528,N_2481,N_2498);
and U2529 (N_2529,N_2422,N_2421);
and U2530 (N_2530,N_2465,N_2456);
or U2531 (N_2531,N_2414,N_2436);
or U2532 (N_2532,N_2488,N_2438);
nand U2533 (N_2533,N_2410,N_2473);
nand U2534 (N_2534,N_2450,N_2447);
and U2535 (N_2535,N_2484,N_2444);
xnor U2536 (N_2536,N_2406,N_2413);
nor U2537 (N_2537,N_2411,N_2480);
or U2538 (N_2538,N_2468,N_2400);
and U2539 (N_2539,N_2478,N_2459);
or U2540 (N_2540,N_2420,N_2476);
nor U2541 (N_2541,N_2408,N_2442);
nand U2542 (N_2542,N_2427,N_2419);
nand U2543 (N_2543,N_2434,N_2404);
nand U2544 (N_2544,N_2491,N_2451);
or U2545 (N_2545,N_2474,N_2454);
nand U2546 (N_2546,N_2440,N_2477);
or U2547 (N_2547,N_2441,N_2494);
nand U2548 (N_2548,N_2485,N_2489);
and U2549 (N_2549,N_2497,N_2457);
nand U2550 (N_2550,N_2430,N_2468);
nor U2551 (N_2551,N_2462,N_2400);
nand U2552 (N_2552,N_2499,N_2401);
or U2553 (N_2553,N_2474,N_2462);
nand U2554 (N_2554,N_2438,N_2453);
xnor U2555 (N_2555,N_2416,N_2410);
nor U2556 (N_2556,N_2423,N_2436);
or U2557 (N_2557,N_2477,N_2452);
xor U2558 (N_2558,N_2411,N_2452);
nor U2559 (N_2559,N_2499,N_2463);
and U2560 (N_2560,N_2413,N_2431);
nand U2561 (N_2561,N_2441,N_2445);
and U2562 (N_2562,N_2401,N_2487);
nor U2563 (N_2563,N_2470,N_2406);
or U2564 (N_2564,N_2422,N_2404);
or U2565 (N_2565,N_2420,N_2441);
xor U2566 (N_2566,N_2445,N_2480);
or U2567 (N_2567,N_2441,N_2448);
xnor U2568 (N_2568,N_2455,N_2420);
nor U2569 (N_2569,N_2463,N_2402);
nand U2570 (N_2570,N_2423,N_2439);
nand U2571 (N_2571,N_2495,N_2404);
nand U2572 (N_2572,N_2439,N_2434);
nor U2573 (N_2573,N_2428,N_2488);
nand U2574 (N_2574,N_2405,N_2445);
nor U2575 (N_2575,N_2447,N_2417);
and U2576 (N_2576,N_2411,N_2406);
nand U2577 (N_2577,N_2441,N_2470);
or U2578 (N_2578,N_2422,N_2456);
or U2579 (N_2579,N_2494,N_2475);
xor U2580 (N_2580,N_2480,N_2469);
and U2581 (N_2581,N_2415,N_2473);
and U2582 (N_2582,N_2492,N_2443);
or U2583 (N_2583,N_2451,N_2408);
nor U2584 (N_2584,N_2485,N_2404);
nor U2585 (N_2585,N_2467,N_2415);
xor U2586 (N_2586,N_2451,N_2429);
xnor U2587 (N_2587,N_2443,N_2420);
nand U2588 (N_2588,N_2448,N_2434);
and U2589 (N_2589,N_2498,N_2430);
nor U2590 (N_2590,N_2460,N_2456);
or U2591 (N_2591,N_2445,N_2472);
xor U2592 (N_2592,N_2488,N_2477);
nand U2593 (N_2593,N_2450,N_2430);
nor U2594 (N_2594,N_2459,N_2403);
nand U2595 (N_2595,N_2499,N_2488);
nand U2596 (N_2596,N_2455,N_2431);
nor U2597 (N_2597,N_2430,N_2496);
or U2598 (N_2598,N_2449,N_2405);
nand U2599 (N_2599,N_2461,N_2472);
xor U2600 (N_2600,N_2560,N_2576);
or U2601 (N_2601,N_2524,N_2516);
and U2602 (N_2602,N_2587,N_2597);
xnor U2603 (N_2603,N_2579,N_2543);
nand U2604 (N_2604,N_2520,N_2574);
and U2605 (N_2605,N_2562,N_2592);
or U2606 (N_2606,N_2536,N_2572);
nor U2607 (N_2607,N_2507,N_2512);
or U2608 (N_2608,N_2521,N_2561);
and U2609 (N_2609,N_2591,N_2586);
nand U2610 (N_2610,N_2533,N_2510);
or U2611 (N_2611,N_2511,N_2509);
and U2612 (N_2612,N_2565,N_2567);
xor U2613 (N_2613,N_2588,N_2550);
nor U2614 (N_2614,N_2580,N_2559);
nand U2615 (N_2615,N_2593,N_2599);
nor U2616 (N_2616,N_2563,N_2535);
and U2617 (N_2617,N_2568,N_2502);
nor U2618 (N_2618,N_2542,N_2553);
and U2619 (N_2619,N_2551,N_2529);
nand U2620 (N_2620,N_2545,N_2538);
nor U2621 (N_2621,N_2589,N_2577);
and U2622 (N_2622,N_2517,N_2596);
nor U2623 (N_2623,N_2526,N_2528);
and U2624 (N_2624,N_2501,N_2573);
and U2625 (N_2625,N_2531,N_2530);
nor U2626 (N_2626,N_2558,N_2544);
nor U2627 (N_2627,N_2590,N_2504);
nor U2628 (N_2628,N_2569,N_2583);
or U2629 (N_2629,N_2505,N_2578);
xor U2630 (N_2630,N_2513,N_2566);
or U2631 (N_2631,N_2582,N_2503);
nand U2632 (N_2632,N_2519,N_2554);
or U2633 (N_2633,N_2525,N_2541);
nor U2634 (N_2634,N_2546,N_2584);
nor U2635 (N_2635,N_2532,N_2556);
nand U2636 (N_2636,N_2581,N_2594);
or U2637 (N_2637,N_2515,N_2518);
nand U2638 (N_2638,N_2575,N_2598);
nand U2639 (N_2639,N_2500,N_2570);
or U2640 (N_2640,N_2555,N_2540);
nor U2641 (N_2641,N_2514,N_2523);
nor U2642 (N_2642,N_2547,N_2537);
or U2643 (N_2643,N_2571,N_2534);
xnor U2644 (N_2644,N_2508,N_2522);
nor U2645 (N_2645,N_2506,N_2527);
xor U2646 (N_2646,N_2552,N_2595);
and U2647 (N_2647,N_2557,N_2539);
or U2648 (N_2648,N_2548,N_2549);
and U2649 (N_2649,N_2585,N_2564);
or U2650 (N_2650,N_2505,N_2551);
or U2651 (N_2651,N_2549,N_2539);
xor U2652 (N_2652,N_2560,N_2596);
and U2653 (N_2653,N_2570,N_2505);
nand U2654 (N_2654,N_2509,N_2546);
nand U2655 (N_2655,N_2594,N_2567);
or U2656 (N_2656,N_2523,N_2520);
nand U2657 (N_2657,N_2523,N_2560);
nor U2658 (N_2658,N_2501,N_2542);
nand U2659 (N_2659,N_2571,N_2566);
and U2660 (N_2660,N_2548,N_2592);
nor U2661 (N_2661,N_2525,N_2521);
xnor U2662 (N_2662,N_2595,N_2599);
and U2663 (N_2663,N_2515,N_2559);
and U2664 (N_2664,N_2506,N_2585);
nand U2665 (N_2665,N_2548,N_2582);
and U2666 (N_2666,N_2569,N_2519);
nand U2667 (N_2667,N_2585,N_2532);
xor U2668 (N_2668,N_2559,N_2585);
and U2669 (N_2669,N_2501,N_2534);
xnor U2670 (N_2670,N_2555,N_2560);
and U2671 (N_2671,N_2593,N_2533);
xnor U2672 (N_2672,N_2594,N_2588);
nor U2673 (N_2673,N_2590,N_2560);
xnor U2674 (N_2674,N_2570,N_2567);
or U2675 (N_2675,N_2531,N_2504);
nand U2676 (N_2676,N_2512,N_2559);
and U2677 (N_2677,N_2583,N_2500);
and U2678 (N_2678,N_2572,N_2562);
or U2679 (N_2679,N_2569,N_2575);
or U2680 (N_2680,N_2580,N_2579);
nand U2681 (N_2681,N_2547,N_2583);
nor U2682 (N_2682,N_2594,N_2527);
or U2683 (N_2683,N_2536,N_2528);
or U2684 (N_2684,N_2596,N_2553);
xor U2685 (N_2685,N_2513,N_2531);
xor U2686 (N_2686,N_2518,N_2555);
or U2687 (N_2687,N_2585,N_2533);
nand U2688 (N_2688,N_2566,N_2538);
nand U2689 (N_2689,N_2586,N_2553);
nand U2690 (N_2690,N_2522,N_2515);
xor U2691 (N_2691,N_2524,N_2545);
nand U2692 (N_2692,N_2526,N_2511);
xor U2693 (N_2693,N_2580,N_2513);
and U2694 (N_2694,N_2577,N_2518);
or U2695 (N_2695,N_2586,N_2572);
or U2696 (N_2696,N_2558,N_2565);
nand U2697 (N_2697,N_2594,N_2531);
nor U2698 (N_2698,N_2590,N_2506);
or U2699 (N_2699,N_2578,N_2525);
and U2700 (N_2700,N_2655,N_2693);
nor U2701 (N_2701,N_2664,N_2661);
nand U2702 (N_2702,N_2616,N_2682);
and U2703 (N_2703,N_2650,N_2642);
nor U2704 (N_2704,N_2606,N_2681);
and U2705 (N_2705,N_2654,N_2626);
nor U2706 (N_2706,N_2687,N_2696);
or U2707 (N_2707,N_2645,N_2691);
nor U2708 (N_2708,N_2651,N_2614);
nand U2709 (N_2709,N_2656,N_2692);
and U2710 (N_2710,N_2644,N_2653);
or U2711 (N_2711,N_2637,N_2622);
and U2712 (N_2712,N_2631,N_2649);
and U2713 (N_2713,N_2613,N_2697);
nor U2714 (N_2714,N_2625,N_2686);
or U2715 (N_2715,N_2663,N_2677);
nand U2716 (N_2716,N_2623,N_2675);
or U2717 (N_2717,N_2646,N_2619);
nor U2718 (N_2718,N_2684,N_2640);
xor U2719 (N_2719,N_2669,N_2609);
and U2720 (N_2720,N_2610,N_2647);
or U2721 (N_2721,N_2601,N_2673);
nand U2722 (N_2722,N_2603,N_2615);
nand U2723 (N_2723,N_2662,N_2628);
or U2724 (N_2724,N_2658,N_2634);
or U2725 (N_2725,N_2688,N_2629);
and U2726 (N_2726,N_2676,N_2689);
or U2727 (N_2727,N_2690,N_2698);
nor U2728 (N_2728,N_2665,N_2608);
nand U2729 (N_2729,N_2672,N_2671);
nand U2730 (N_2730,N_2604,N_2611);
or U2731 (N_2731,N_2600,N_2659);
nand U2732 (N_2732,N_2630,N_2617);
and U2733 (N_2733,N_2683,N_2605);
and U2734 (N_2734,N_2643,N_2620);
or U2735 (N_2735,N_2667,N_2618);
nor U2736 (N_2736,N_2632,N_2602);
and U2737 (N_2737,N_2670,N_2621);
nor U2738 (N_2738,N_2657,N_2624);
nand U2739 (N_2739,N_2678,N_2639);
or U2740 (N_2740,N_2627,N_2652);
nand U2741 (N_2741,N_2685,N_2636);
nor U2742 (N_2742,N_2666,N_2679);
and U2743 (N_2743,N_2694,N_2638);
nor U2744 (N_2744,N_2695,N_2680);
nor U2745 (N_2745,N_2674,N_2635);
xor U2746 (N_2746,N_2668,N_2607);
and U2747 (N_2747,N_2660,N_2612);
and U2748 (N_2748,N_2633,N_2699);
and U2749 (N_2749,N_2641,N_2648);
nand U2750 (N_2750,N_2603,N_2626);
nand U2751 (N_2751,N_2694,N_2628);
nor U2752 (N_2752,N_2673,N_2675);
or U2753 (N_2753,N_2670,N_2669);
nor U2754 (N_2754,N_2636,N_2698);
nand U2755 (N_2755,N_2613,N_2698);
and U2756 (N_2756,N_2662,N_2604);
nand U2757 (N_2757,N_2619,N_2611);
nor U2758 (N_2758,N_2640,N_2607);
nor U2759 (N_2759,N_2601,N_2649);
nand U2760 (N_2760,N_2612,N_2669);
nand U2761 (N_2761,N_2691,N_2697);
and U2762 (N_2762,N_2601,N_2658);
and U2763 (N_2763,N_2618,N_2646);
or U2764 (N_2764,N_2670,N_2620);
nand U2765 (N_2765,N_2692,N_2674);
nor U2766 (N_2766,N_2639,N_2646);
xor U2767 (N_2767,N_2685,N_2695);
nor U2768 (N_2768,N_2673,N_2646);
or U2769 (N_2769,N_2602,N_2680);
xor U2770 (N_2770,N_2627,N_2646);
nand U2771 (N_2771,N_2647,N_2668);
and U2772 (N_2772,N_2614,N_2673);
nand U2773 (N_2773,N_2694,N_2673);
and U2774 (N_2774,N_2641,N_2678);
nand U2775 (N_2775,N_2692,N_2614);
nor U2776 (N_2776,N_2651,N_2644);
xor U2777 (N_2777,N_2669,N_2695);
nand U2778 (N_2778,N_2609,N_2665);
or U2779 (N_2779,N_2624,N_2610);
nor U2780 (N_2780,N_2638,N_2615);
or U2781 (N_2781,N_2633,N_2697);
xnor U2782 (N_2782,N_2621,N_2624);
and U2783 (N_2783,N_2682,N_2629);
or U2784 (N_2784,N_2680,N_2614);
nor U2785 (N_2785,N_2622,N_2681);
and U2786 (N_2786,N_2679,N_2610);
nand U2787 (N_2787,N_2652,N_2615);
or U2788 (N_2788,N_2612,N_2640);
or U2789 (N_2789,N_2613,N_2658);
and U2790 (N_2790,N_2668,N_2688);
nor U2791 (N_2791,N_2694,N_2639);
nor U2792 (N_2792,N_2610,N_2620);
or U2793 (N_2793,N_2616,N_2650);
or U2794 (N_2794,N_2688,N_2627);
nand U2795 (N_2795,N_2648,N_2683);
and U2796 (N_2796,N_2684,N_2606);
xor U2797 (N_2797,N_2664,N_2659);
or U2798 (N_2798,N_2691,N_2641);
nor U2799 (N_2799,N_2624,N_2623);
and U2800 (N_2800,N_2773,N_2748);
nor U2801 (N_2801,N_2745,N_2718);
nand U2802 (N_2802,N_2738,N_2705);
or U2803 (N_2803,N_2727,N_2782);
nand U2804 (N_2804,N_2704,N_2708);
or U2805 (N_2805,N_2795,N_2766);
or U2806 (N_2806,N_2728,N_2781);
nor U2807 (N_2807,N_2752,N_2702);
and U2808 (N_2808,N_2751,N_2730);
or U2809 (N_2809,N_2713,N_2799);
nor U2810 (N_2810,N_2753,N_2707);
nor U2811 (N_2811,N_2716,N_2714);
and U2812 (N_2812,N_2749,N_2767);
nor U2813 (N_2813,N_2709,N_2755);
or U2814 (N_2814,N_2736,N_2763);
nand U2815 (N_2815,N_2740,N_2757);
xor U2816 (N_2816,N_2787,N_2743);
nand U2817 (N_2817,N_2756,N_2733);
nor U2818 (N_2818,N_2762,N_2722);
nor U2819 (N_2819,N_2790,N_2779);
nand U2820 (N_2820,N_2765,N_2764);
and U2821 (N_2821,N_2724,N_2711);
or U2822 (N_2822,N_2793,N_2706);
xnor U2823 (N_2823,N_2785,N_2796);
nor U2824 (N_2824,N_2798,N_2791);
nor U2825 (N_2825,N_2780,N_2777);
or U2826 (N_2826,N_2701,N_2744);
nor U2827 (N_2827,N_2784,N_2770);
nand U2828 (N_2828,N_2720,N_2786);
nand U2829 (N_2829,N_2768,N_2797);
or U2830 (N_2830,N_2760,N_2771);
nor U2831 (N_2831,N_2778,N_2739);
and U2832 (N_2832,N_2726,N_2735);
nand U2833 (N_2833,N_2732,N_2742);
or U2834 (N_2834,N_2712,N_2725);
and U2835 (N_2835,N_2717,N_2723);
and U2836 (N_2836,N_2700,N_2772);
and U2837 (N_2837,N_2729,N_2759);
nor U2838 (N_2838,N_2758,N_2703);
or U2839 (N_2839,N_2754,N_2774);
and U2840 (N_2840,N_2788,N_2783);
nor U2841 (N_2841,N_2721,N_2737);
or U2842 (N_2842,N_2747,N_2731);
nor U2843 (N_2843,N_2761,N_2776);
or U2844 (N_2844,N_2769,N_2789);
nor U2845 (N_2845,N_2792,N_2750);
and U2846 (N_2846,N_2775,N_2719);
nand U2847 (N_2847,N_2710,N_2715);
and U2848 (N_2848,N_2794,N_2746);
nor U2849 (N_2849,N_2741,N_2734);
or U2850 (N_2850,N_2759,N_2739);
and U2851 (N_2851,N_2740,N_2766);
and U2852 (N_2852,N_2794,N_2756);
or U2853 (N_2853,N_2741,N_2709);
xor U2854 (N_2854,N_2731,N_2772);
xnor U2855 (N_2855,N_2797,N_2739);
and U2856 (N_2856,N_2738,N_2724);
xor U2857 (N_2857,N_2739,N_2766);
nor U2858 (N_2858,N_2715,N_2745);
or U2859 (N_2859,N_2742,N_2799);
or U2860 (N_2860,N_2745,N_2779);
or U2861 (N_2861,N_2730,N_2725);
nand U2862 (N_2862,N_2774,N_2701);
and U2863 (N_2863,N_2744,N_2752);
or U2864 (N_2864,N_2752,N_2757);
and U2865 (N_2865,N_2731,N_2794);
and U2866 (N_2866,N_2794,N_2787);
nor U2867 (N_2867,N_2799,N_2722);
nor U2868 (N_2868,N_2782,N_2742);
or U2869 (N_2869,N_2727,N_2772);
or U2870 (N_2870,N_2712,N_2776);
and U2871 (N_2871,N_2757,N_2723);
and U2872 (N_2872,N_2745,N_2777);
and U2873 (N_2873,N_2788,N_2748);
and U2874 (N_2874,N_2772,N_2732);
xor U2875 (N_2875,N_2723,N_2752);
nor U2876 (N_2876,N_2754,N_2745);
or U2877 (N_2877,N_2707,N_2743);
nor U2878 (N_2878,N_2770,N_2728);
nand U2879 (N_2879,N_2724,N_2740);
xor U2880 (N_2880,N_2723,N_2724);
nor U2881 (N_2881,N_2719,N_2791);
nand U2882 (N_2882,N_2791,N_2705);
and U2883 (N_2883,N_2789,N_2799);
nand U2884 (N_2884,N_2767,N_2733);
and U2885 (N_2885,N_2755,N_2736);
nand U2886 (N_2886,N_2748,N_2732);
nor U2887 (N_2887,N_2757,N_2704);
xor U2888 (N_2888,N_2767,N_2781);
nor U2889 (N_2889,N_2747,N_2759);
and U2890 (N_2890,N_2793,N_2774);
and U2891 (N_2891,N_2745,N_2785);
and U2892 (N_2892,N_2744,N_2747);
and U2893 (N_2893,N_2718,N_2771);
nor U2894 (N_2894,N_2779,N_2726);
nand U2895 (N_2895,N_2775,N_2707);
and U2896 (N_2896,N_2750,N_2709);
or U2897 (N_2897,N_2742,N_2709);
nor U2898 (N_2898,N_2795,N_2736);
xnor U2899 (N_2899,N_2780,N_2745);
or U2900 (N_2900,N_2861,N_2892);
nor U2901 (N_2901,N_2893,N_2825);
xnor U2902 (N_2902,N_2820,N_2835);
xor U2903 (N_2903,N_2823,N_2867);
nor U2904 (N_2904,N_2811,N_2887);
nor U2905 (N_2905,N_2853,N_2809);
nand U2906 (N_2906,N_2882,N_2877);
xor U2907 (N_2907,N_2874,N_2840);
and U2908 (N_2908,N_2841,N_2851);
or U2909 (N_2909,N_2888,N_2824);
nor U2910 (N_2910,N_2846,N_2829);
nand U2911 (N_2911,N_2873,N_2897);
xor U2912 (N_2912,N_2859,N_2808);
or U2913 (N_2913,N_2881,N_2828);
and U2914 (N_2914,N_2844,N_2850);
nand U2915 (N_2915,N_2863,N_2884);
xor U2916 (N_2916,N_2890,N_2896);
and U2917 (N_2917,N_2845,N_2800);
nor U2918 (N_2918,N_2802,N_2880);
nor U2919 (N_2919,N_2810,N_2836);
and U2920 (N_2920,N_2813,N_2869);
nor U2921 (N_2921,N_2868,N_2807);
nor U2922 (N_2922,N_2806,N_2830);
nand U2923 (N_2923,N_2826,N_2838);
nor U2924 (N_2924,N_2821,N_2866);
or U2925 (N_2925,N_2878,N_2883);
xor U2926 (N_2926,N_2865,N_2849);
xnor U2927 (N_2927,N_2886,N_2801);
nor U2928 (N_2928,N_2832,N_2879);
xnor U2929 (N_2929,N_2889,N_2875);
and U2930 (N_2930,N_2857,N_2831);
nor U2931 (N_2931,N_2822,N_2833);
nor U2932 (N_2932,N_2812,N_2864);
and U2933 (N_2933,N_2871,N_2827);
or U2934 (N_2934,N_2894,N_2848);
nor U2935 (N_2935,N_2862,N_2842);
nand U2936 (N_2936,N_2895,N_2815);
or U2937 (N_2937,N_2803,N_2816);
nand U2938 (N_2938,N_2854,N_2805);
and U2939 (N_2939,N_2852,N_2804);
xor U2940 (N_2940,N_2843,N_2858);
and U2941 (N_2941,N_2839,N_2870);
nand U2942 (N_2942,N_2819,N_2899);
xnor U2943 (N_2943,N_2898,N_2818);
nand U2944 (N_2944,N_2837,N_2847);
nor U2945 (N_2945,N_2876,N_2885);
nand U2946 (N_2946,N_2872,N_2856);
xor U2947 (N_2947,N_2855,N_2860);
nor U2948 (N_2948,N_2891,N_2814);
and U2949 (N_2949,N_2834,N_2817);
nand U2950 (N_2950,N_2889,N_2841);
or U2951 (N_2951,N_2801,N_2832);
nand U2952 (N_2952,N_2836,N_2819);
nand U2953 (N_2953,N_2804,N_2821);
and U2954 (N_2954,N_2830,N_2839);
nand U2955 (N_2955,N_2814,N_2835);
nor U2956 (N_2956,N_2853,N_2897);
or U2957 (N_2957,N_2877,N_2821);
or U2958 (N_2958,N_2803,N_2820);
or U2959 (N_2959,N_2853,N_2839);
nor U2960 (N_2960,N_2871,N_2815);
nor U2961 (N_2961,N_2869,N_2876);
and U2962 (N_2962,N_2852,N_2898);
and U2963 (N_2963,N_2847,N_2890);
nand U2964 (N_2964,N_2807,N_2838);
nor U2965 (N_2965,N_2802,N_2889);
and U2966 (N_2966,N_2834,N_2804);
xnor U2967 (N_2967,N_2804,N_2859);
xnor U2968 (N_2968,N_2807,N_2837);
or U2969 (N_2969,N_2823,N_2857);
nand U2970 (N_2970,N_2880,N_2854);
nand U2971 (N_2971,N_2856,N_2832);
or U2972 (N_2972,N_2816,N_2828);
and U2973 (N_2973,N_2862,N_2877);
xor U2974 (N_2974,N_2873,N_2863);
and U2975 (N_2975,N_2890,N_2844);
or U2976 (N_2976,N_2887,N_2861);
or U2977 (N_2977,N_2813,N_2830);
and U2978 (N_2978,N_2832,N_2874);
or U2979 (N_2979,N_2850,N_2881);
nor U2980 (N_2980,N_2885,N_2841);
nand U2981 (N_2981,N_2819,N_2803);
and U2982 (N_2982,N_2803,N_2851);
nor U2983 (N_2983,N_2867,N_2851);
and U2984 (N_2984,N_2855,N_2882);
nand U2985 (N_2985,N_2888,N_2842);
xnor U2986 (N_2986,N_2855,N_2848);
or U2987 (N_2987,N_2832,N_2866);
or U2988 (N_2988,N_2841,N_2829);
and U2989 (N_2989,N_2863,N_2894);
and U2990 (N_2990,N_2856,N_2869);
nand U2991 (N_2991,N_2871,N_2898);
nor U2992 (N_2992,N_2831,N_2813);
nand U2993 (N_2993,N_2862,N_2882);
nor U2994 (N_2994,N_2863,N_2866);
and U2995 (N_2995,N_2895,N_2887);
nor U2996 (N_2996,N_2801,N_2835);
nor U2997 (N_2997,N_2836,N_2803);
or U2998 (N_2998,N_2878,N_2894);
or U2999 (N_2999,N_2856,N_2881);
nand UO_0 (O_0,N_2927,N_2912);
and UO_1 (O_1,N_2910,N_2983);
nor UO_2 (O_2,N_2956,N_2941);
nand UO_3 (O_3,N_2967,N_2951);
xnor UO_4 (O_4,N_2945,N_2992);
or UO_5 (O_5,N_2999,N_2977);
nor UO_6 (O_6,N_2918,N_2919);
or UO_7 (O_7,N_2990,N_2985);
or UO_8 (O_8,N_2902,N_2900);
and UO_9 (O_9,N_2955,N_2933);
or UO_10 (O_10,N_2929,N_2973);
or UO_11 (O_11,N_2980,N_2989);
nand UO_12 (O_12,N_2972,N_2964);
nand UO_13 (O_13,N_2991,N_2965);
nand UO_14 (O_14,N_2966,N_2969);
nand UO_15 (O_15,N_2911,N_2914);
nor UO_16 (O_16,N_2931,N_2930);
nor UO_17 (O_17,N_2906,N_2960);
and UO_18 (O_18,N_2908,N_2921);
nand UO_19 (O_19,N_2981,N_2909);
or UO_20 (O_20,N_2978,N_2994);
nand UO_21 (O_21,N_2950,N_2949);
or UO_22 (O_22,N_2905,N_2947);
nand UO_23 (O_23,N_2901,N_2935);
xor UO_24 (O_24,N_2971,N_2915);
nor UO_25 (O_25,N_2904,N_2913);
nor UO_26 (O_26,N_2907,N_2962);
or UO_27 (O_27,N_2963,N_2976);
nand UO_28 (O_28,N_2952,N_2953);
nor UO_29 (O_29,N_2938,N_2957);
nand UO_30 (O_30,N_2984,N_2958);
nand UO_31 (O_31,N_2988,N_2934);
and UO_32 (O_32,N_2997,N_2944);
or UO_33 (O_33,N_2995,N_2925);
nand UO_34 (O_34,N_2946,N_2942);
or UO_35 (O_35,N_2924,N_2926);
xnor UO_36 (O_36,N_2974,N_2959);
and UO_37 (O_37,N_2943,N_2916);
nor UO_38 (O_38,N_2937,N_2939);
nand UO_39 (O_39,N_2970,N_2993);
nor UO_40 (O_40,N_2968,N_2954);
nor UO_41 (O_41,N_2903,N_2940);
nor UO_42 (O_42,N_2996,N_2979);
nor UO_43 (O_43,N_2975,N_2961);
nand UO_44 (O_44,N_2920,N_2917);
and UO_45 (O_45,N_2987,N_2923);
nor UO_46 (O_46,N_2922,N_2998);
and UO_47 (O_47,N_2936,N_2986);
nor UO_48 (O_48,N_2932,N_2948);
nand UO_49 (O_49,N_2928,N_2982);
xor UO_50 (O_50,N_2910,N_2966);
or UO_51 (O_51,N_2908,N_2996);
or UO_52 (O_52,N_2985,N_2910);
nand UO_53 (O_53,N_2972,N_2906);
nor UO_54 (O_54,N_2940,N_2993);
or UO_55 (O_55,N_2932,N_2988);
nand UO_56 (O_56,N_2980,N_2927);
nor UO_57 (O_57,N_2929,N_2940);
nand UO_58 (O_58,N_2941,N_2957);
nand UO_59 (O_59,N_2996,N_2907);
xor UO_60 (O_60,N_2949,N_2966);
nand UO_61 (O_61,N_2995,N_2933);
nor UO_62 (O_62,N_2969,N_2965);
xnor UO_63 (O_63,N_2936,N_2977);
nor UO_64 (O_64,N_2994,N_2991);
nor UO_65 (O_65,N_2942,N_2965);
nor UO_66 (O_66,N_2904,N_2974);
xnor UO_67 (O_67,N_2913,N_2910);
and UO_68 (O_68,N_2988,N_2912);
nor UO_69 (O_69,N_2954,N_2985);
nor UO_70 (O_70,N_2993,N_2951);
and UO_71 (O_71,N_2909,N_2941);
nor UO_72 (O_72,N_2930,N_2912);
nor UO_73 (O_73,N_2987,N_2949);
or UO_74 (O_74,N_2913,N_2969);
nor UO_75 (O_75,N_2914,N_2916);
and UO_76 (O_76,N_2923,N_2998);
and UO_77 (O_77,N_2963,N_2937);
nand UO_78 (O_78,N_2914,N_2906);
or UO_79 (O_79,N_2934,N_2962);
and UO_80 (O_80,N_2920,N_2961);
and UO_81 (O_81,N_2914,N_2987);
or UO_82 (O_82,N_2927,N_2951);
nand UO_83 (O_83,N_2975,N_2915);
nand UO_84 (O_84,N_2981,N_2945);
nand UO_85 (O_85,N_2936,N_2901);
xnor UO_86 (O_86,N_2930,N_2913);
or UO_87 (O_87,N_2960,N_2912);
nand UO_88 (O_88,N_2986,N_2947);
nor UO_89 (O_89,N_2921,N_2920);
nor UO_90 (O_90,N_2970,N_2946);
nand UO_91 (O_91,N_2947,N_2957);
or UO_92 (O_92,N_2967,N_2955);
and UO_93 (O_93,N_2961,N_2950);
nor UO_94 (O_94,N_2931,N_2947);
or UO_95 (O_95,N_2905,N_2985);
nand UO_96 (O_96,N_2941,N_2925);
nand UO_97 (O_97,N_2913,N_2949);
nor UO_98 (O_98,N_2968,N_2900);
nor UO_99 (O_99,N_2938,N_2908);
and UO_100 (O_100,N_2912,N_2969);
nor UO_101 (O_101,N_2941,N_2966);
or UO_102 (O_102,N_2977,N_2983);
xor UO_103 (O_103,N_2954,N_2900);
xnor UO_104 (O_104,N_2981,N_2954);
nor UO_105 (O_105,N_2929,N_2979);
or UO_106 (O_106,N_2996,N_2969);
or UO_107 (O_107,N_2930,N_2940);
nand UO_108 (O_108,N_2990,N_2949);
nand UO_109 (O_109,N_2930,N_2933);
or UO_110 (O_110,N_2996,N_2992);
and UO_111 (O_111,N_2903,N_2927);
nor UO_112 (O_112,N_2985,N_2958);
nand UO_113 (O_113,N_2923,N_2928);
or UO_114 (O_114,N_2922,N_2984);
and UO_115 (O_115,N_2941,N_2921);
nand UO_116 (O_116,N_2960,N_2910);
and UO_117 (O_117,N_2967,N_2952);
or UO_118 (O_118,N_2912,N_2944);
or UO_119 (O_119,N_2923,N_2950);
nor UO_120 (O_120,N_2925,N_2932);
or UO_121 (O_121,N_2990,N_2989);
and UO_122 (O_122,N_2979,N_2992);
and UO_123 (O_123,N_2945,N_2936);
and UO_124 (O_124,N_2956,N_2967);
or UO_125 (O_125,N_2955,N_2972);
xnor UO_126 (O_126,N_2962,N_2999);
xnor UO_127 (O_127,N_2965,N_2960);
xor UO_128 (O_128,N_2927,N_2950);
or UO_129 (O_129,N_2973,N_2972);
nor UO_130 (O_130,N_2949,N_2997);
or UO_131 (O_131,N_2920,N_2996);
nand UO_132 (O_132,N_2930,N_2996);
and UO_133 (O_133,N_2940,N_2939);
or UO_134 (O_134,N_2936,N_2944);
or UO_135 (O_135,N_2920,N_2977);
or UO_136 (O_136,N_2996,N_2991);
nand UO_137 (O_137,N_2983,N_2961);
nand UO_138 (O_138,N_2966,N_2964);
and UO_139 (O_139,N_2954,N_2913);
and UO_140 (O_140,N_2985,N_2945);
or UO_141 (O_141,N_2953,N_2954);
or UO_142 (O_142,N_2999,N_2937);
nand UO_143 (O_143,N_2908,N_2919);
nand UO_144 (O_144,N_2967,N_2939);
or UO_145 (O_145,N_2955,N_2984);
and UO_146 (O_146,N_2951,N_2940);
nand UO_147 (O_147,N_2946,N_2917);
and UO_148 (O_148,N_2990,N_2991);
nor UO_149 (O_149,N_2957,N_2908);
and UO_150 (O_150,N_2936,N_2995);
and UO_151 (O_151,N_2938,N_2923);
and UO_152 (O_152,N_2950,N_2969);
and UO_153 (O_153,N_2968,N_2925);
or UO_154 (O_154,N_2954,N_2922);
nor UO_155 (O_155,N_2949,N_2958);
or UO_156 (O_156,N_2901,N_2937);
nand UO_157 (O_157,N_2998,N_2958);
nand UO_158 (O_158,N_2907,N_2944);
or UO_159 (O_159,N_2910,N_2984);
nor UO_160 (O_160,N_2989,N_2942);
nand UO_161 (O_161,N_2977,N_2941);
and UO_162 (O_162,N_2977,N_2940);
and UO_163 (O_163,N_2961,N_2971);
nor UO_164 (O_164,N_2994,N_2902);
nand UO_165 (O_165,N_2908,N_2912);
xnor UO_166 (O_166,N_2939,N_2985);
and UO_167 (O_167,N_2938,N_2998);
and UO_168 (O_168,N_2926,N_2955);
and UO_169 (O_169,N_2912,N_2998);
or UO_170 (O_170,N_2980,N_2986);
nand UO_171 (O_171,N_2979,N_2988);
or UO_172 (O_172,N_2917,N_2968);
nand UO_173 (O_173,N_2927,N_2920);
nand UO_174 (O_174,N_2954,N_2915);
and UO_175 (O_175,N_2932,N_2902);
and UO_176 (O_176,N_2934,N_2977);
or UO_177 (O_177,N_2977,N_2923);
and UO_178 (O_178,N_2919,N_2975);
or UO_179 (O_179,N_2913,N_2967);
nor UO_180 (O_180,N_2901,N_2908);
nor UO_181 (O_181,N_2944,N_2996);
and UO_182 (O_182,N_2983,N_2979);
or UO_183 (O_183,N_2948,N_2964);
nor UO_184 (O_184,N_2953,N_2995);
nor UO_185 (O_185,N_2954,N_2926);
xor UO_186 (O_186,N_2924,N_2972);
and UO_187 (O_187,N_2941,N_2927);
nor UO_188 (O_188,N_2982,N_2990);
or UO_189 (O_189,N_2943,N_2982);
and UO_190 (O_190,N_2999,N_2974);
nor UO_191 (O_191,N_2963,N_2968);
or UO_192 (O_192,N_2951,N_2904);
nand UO_193 (O_193,N_2963,N_2913);
xor UO_194 (O_194,N_2968,N_2941);
nor UO_195 (O_195,N_2966,N_2921);
and UO_196 (O_196,N_2932,N_2901);
or UO_197 (O_197,N_2976,N_2916);
nand UO_198 (O_198,N_2917,N_2928);
and UO_199 (O_199,N_2990,N_2962);
or UO_200 (O_200,N_2962,N_2944);
and UO_201 (O_201,N_2934,N_2954);
xnor UO_202 (O_202,N_2994,N_2981);
nand UO_203 (O_203,N_2955,N_2974);
nand UO_204 (O_204,N_2984,N_2912);
and UO_205 (O_205,N_2901,N_2950);
nor UO_206 (O_206,N_2994,N_2949);
xor UO_207 (O_207,N_2970,N_2913);
xor UO_208 (O_208,N_2983,N_2947);
nor UO_209 (O_209,N_2955,N_2966);
or UO_210 (O_210,N_2920,N_2900);
or UO_211 (O_211,N_2985,N_2992);
or UO_212 (O_212,N_2916,N_2959);
nor UO_213 (O_213,N_2980,N_2992);
nor UO_214 (O_214,N_2964,N_2951);
nand UO_215 (O_215,N_2993,N_2968);
nand UO_216 (O_216,N_2914,N_2986);
nor UO_217 (O_217,N_2926,N_2908);
nand UO_218 (O_218,N_2967,N_2923);
nor UO_219 (O_219,N_2971,N_2940);
or UO_220 (O_220,N_2940,N_2952);
or UO_221 (O_221,N_2974,N_2994);
nand UO_222 (O_222,N_2956,N_2929);
nor UO_223 (O_223,N_2933,N_2925);
xnor UO_224 (O_224,N_2935,N_2982);
nand UO_225 (O_225,N_2972,N_2963);
nor UO_226 (O_226,N_2956,N_2992);
or UO_227 (O_227,N_2920,N_2936);
xnor UO_228 (O_228,N_2909,N_2977);
or UO_229 (O_229,N_2958,N_2938);
nand UO_230 (O_230,N_2937,N_2933);
or UO_231 (O_231,N_2973,N_2906);
nor UO_232 (O_232,N_2970,N_2966);
and UO_233 (O_233,N_2953,N_2966);
nor UO_234 (O_234,N_2971,N_2958);
or UO_235 (O_235,N_2957,N_2914);
nand UO_236 (O_236,N_2909,N_2960);
or UO_237 (O_237,N_2992,N_2931);
and UO_238 (O_238,N_2963,N_2932);
nand UO_239 (O_239,N_2987,N_2977);
nand UO_240 (O_240,N_2972,N_2958);
xnor UO_241 (O_241,N_2916,N_2922);
nand UO_242 (O_242,N_2940,N_2972);
and UO_243 (O_243,N_2904,N_2973);
or UO_244 (O_244,N_2926,N_2962);
or UO_245 (O_245,N_2976,N_2953);
nand UO_246 (O_246,N_2977,N_2904);
nor UO_247 (O_247,N_2999,N_2924);
nor UO_248 (O_248,N_2949,N_2972);
and UO_249 (O_249,N_2945,N_2973);
nor UO_250 (O_250,N_2981,N_2998);
nand UO_251 (O_251,N_2943,N_2949);
and UO_252 (O_252,N_2966,N_2972);
and UO_253 (O_253,N_2942,N_2978);
and UO_254 (O_254,N_2915,N_2992);
nand UO_255 (O_255,N_2901,N_2921);
or UO_256 (O_256,N_2974,N_2968);
and UO_257 (O_257,N_2924,N_2990);
or UO_258 (O_258,N_2910,N_2991);
and UO_259 (O_259,N_2911,N_2934);
nand UO_260 (O_260,N_2943,N_2990);
nand UO_261 (O_261,N_2910,N_2947);
nor UO_262 (O_262,N_2992,N_2904);
and UO_263 (O_263,N_2971,N_2966);
or UO_264 (O_264,N_2917,N_2994);
or UO_265 (O_265,N_2943,N_2950);
nor UO_266 (O_266,N_2956,N_2959);
nand UO_267 (O_267,N_2993,N_2987);
nand UO_268 (O_268,N_2923,N_2956);
nand UO_269 (O_269,N_2948,N_2977);
and UO_270 (O_270,N_2921,N_2980);
nand UO_271 (O_271,N_2940,N_2908);
and UO_272 (O_272,N_2976,N_2926);
and UO_273 (O_273,N_2925,N_2904);
nor UO_274 (O_274,N_2977,N_2955);
nand UO_275 (O_275,N_2961,N_2958);
and UO_276 (O_276,N_2919,N_2956);
xor UO_277 (O_277,N_2951,N_2916);
nand UO_278 (O_278,N_2957,N_2959);
and UO_279 (O_279,N_2999,N_2932);
nand UO_280 (O_280,N_2991,N_2987);
xor UO_281 (O_281,N_2942,N_2991);
and UO_282 (O_282,N_2905,N_2902);
nand UO_283 (O_283,N_2904,N_2937);
and UO_284 (O_284,N_2908,N_2968);
nand UO_285 (O_285,N_2956,N_2930);
nand UO_286 (O_286,N_2906,N_2902);
nor UO_287 (O_287,N_2956,N_2914);
or UO_288 (O_288,N_2925,N_2916);
and UO_289 (O_289,N_2958,N_2995);
nand UO_290 (O_290,N_2974,N_2967);
nor UO_291 (O_291,N_2919,N_2930);
or UO_292 (O_292,N_2919,N_2993);
or UO_293 (O_293,N_2958,N_2956);
nand UO_294 (O_294,N_2941,N_2964);
or UO_295 (O_295,N_2916,N_2972);
nand UO_296 (O_296,N_2969,N_2947);
nand UO_297 (O_297,N_2924,N_2905);
and UO_298 (O_298,N_2998,N_2962);
or UO_299 (O_299,N_2977,N_2981);
or UO_300 (O_300,N_2971,N_2987);
nand UO_301 (O_301,N_2928,N_2904);
nand UO_302 (O_302,N_2943,N_2978);
nor UO_303 (O_303,N_2980,N_2956);
and UO_304 (O_304,N_2942,N_2971);
or UO_305 (O_305,N_2963,N_2925);
xnor UO_306 (O_306,N_2994,N_2967);
and UO_307 (O_307,N_2997,N_2907);
and UO_308 (O_308,N_2910,N_2982);
nand UO_309 (O_309,N_2974,N_2972);
nor UO_310 (O_310,N_2917,N_2955);
xor UO_311 (O_311,N_2936,N_2924);
or UO_312 (O_312,N_2996,N_2988);
nand UO_313 (O_313,N_2913,N_2991);
nand UO_314 (O_314,N_2989,N_2913);
nor UO_315 (O_315,N_2981,N_2937);
nand UO_316 (O_316,N_2981,N_2962);
or UO_317 (O_317,N_2945,N_2998);
and UO_318 (O_318,N_2957,N_2997);
or UO_319 (O_319,N_2947,N_2948);
nand UO_320 (O_320,N_2907,N_2969);
or UO_321 (O_321,N_2947,N_2977);
and UO_322 (O_322,N_2941,N_2973);
or UO_323 (O_323,N_2909,N_2963);
or UO_324 (O_324,N_2989,N_2904);
nor UO_325 (O_325,N_2986,N_2944);
and UO_326 (O_326,N_2924,N_2983);
xor UO_327 (O_327,N_2958,N_2911);
xor UO_328 (O_328,N_2936,N_2982);
and UO_329 (O_329,N_2903,N_2941);
nand UO_330 (O_330,N_2938,N_2915);
or UO_331 (O_331,N_2997,N_2999);
nand UO_332 (O_332,N_2970,N_2947);
and UO_333 (O_333,N_2919,N_2945);
and UO_334 (O_334,N_2991,N_2958);
or UO_335 (O_335,N_2917,N_2971);
or UO_336 (O_336,N_2957,N_2912);
nor UO_337 (O_337,N_2928,N_2967);
nand UO_338 (O_338,N_2989,N_2995);
nand UO_339 (O_339,N_2951,N_2996);
nand UO_340 (O_340,N_2950,N_2953);
nor UO_341 (O_341,N_2990,N_2905);
nand UO_342 (O_342,N_2925,N_2926);
nor UO_343 (O_343,N_2981,N_2956);
and UO_344 (O_344,N_2976,N_2962);
and UO_345 (O_345,N_2945,N_2976);
nor UO_346 (O_346,N_2972,N_2921);
nand UO_347 (O_347,N_2913,N_2956);
nand UO_348 (O_348,N_2935,N_2910);
and UO_349 (O_349,N_2957,N_2901);
and UO_350 (O_350,N_2925,N_2910);
nand UO_351 (O_351,N_2952,N_2970);
or UO_352 (O_352,N_2915,N_2940);
nor UO_353 (O_353,N_2928,N_2995);
nor UO_354 (O_354,N_2919,N_2907);
or UO_355 (O_355,N_2932,N_2996);
nor UO_356 (O_356,N_2967,N_2910);
nor UO_357 (O_357,N_2983,N_2999);
nand UO_358 (O_358,N_2995,N_2954);
and UO_359 (O_359,N_2937,N_2915);
or UO_360 (O_360,N_2914,N_2912);
or UO_361 (O_361,N_2907,N_2965);
xor UO_362 (O_362,N_2934,N_2994);
or UO_363 (O_363,N_2953,N_2967);
nand UO_364 (O_364,N_2959,N_2996);
nor UO_365 (O_365,N_2948,N_2910);
or UO_366 (O_366,N_2926,N_2978);
nand UO_367 (O_367,N_2948,N_2960);
and UO_368 (O_368,N_2990,N_2994);
nand UO_369 (O_369,N_2943,N_2904);
nand UO_370 (O_370,N_2937,N_2977);
nor UO_371 (O_371,N_2971,N_2908);
nor UO_372 (O_372,N_2931,N_2989);
nand UO_373 (O_373,N_2925,N_2930);
nor UO_374 (O_374,N_2974,N_2954);
and UO_375 (O_375,N_2978,N_2992);
xnor UO_376 (O_376,N_2942,N_2967);
nor UO_377 (O_377,N_2975,N_2973);
and UO_378 (O_378,N_2962,N_2904);
and UO_379 (O_379,N_2913,N_2906);
and UO_380 (O_380,N_2913,N_2957);
and UO_381 (O_381,N_2944,N_2903);
nand UO_382 (O_382,N_2961,N_2910);
nand UO_383 (O_383,N_2905,N_2987);
nand UO_384 (O_384,N_2922,N_2945);
nor UO_385 (O_385,N_2945,N_2931);
nand UO_386 (O_386,N_2966,N_2975);
nand UO_387 (O_387,N_2928,N_2965);
or UO_388 (O_388,N_2968,N_2939);
or UO_389 (O_389,N_2985,N_2947);
nand UO_390 (O_390,N_2903,N_2916);
nand UO_391 (O_391,N_2985,N_2983);
nor UO_392 (O_392,N_2934,N_2906);
nor UO_393 (O_393,N_2978,N_2920);
nor UO_394 (O_394,N_2963,N_2918);
nand UO_395 (O_395,N_2992,N_2965);
and UO_396 (O_396,N_2963,N_2982);
nand UO_397 (O_397,N_2957,N_2902);
and UO_398 (O_398,N_2911,N_2951);
nand UO_399 (O_399,N_2939,N_2966);
nand UO_400 (O_400,N_2989,N_2920);
and UO_401 (O_401,N_2994,N_2936);
nor UO_402 (O_402,N_2993,N_2912);
nand UO_403 (O_403,N_2902,N_2910);
or UO_404 (O_404,N_2980,N_2900);
or UO_405 (O_405,N_2951,N_2990);
and UO_406 (O_406,N_2958,N_2947);
nand UO_407 (O_407,N_2959,N_2930);
nand UO_408 (O_408,N_2936,N_2980);
nor UO_409 (O_409,N_2996,N_2975);
and UO_410 (O_410,N_2972,N_2928);
nand UO_411 (O_411,N_2982,N_2959);
xnor UO_412 (O_412,N_2906,N_2970);
nor UO_413 (O_413,N_2917,N_2997);
or UO_414 (O_414,N_2963,N_2908);
or UO_415 (O_415,N_2972,N_2967);
and UO_416 (O_416,N_2973,N_2986);
nor UO_417 (O_417,N_2945,N_2946);
or UO_418 (O_418,N_2986,N_2940);
nand UO_419 (O_419,N_2931,N_2994);
nor UO_420 (O_420,N_2941,N_2991);
or UO_421 (O_421,N_2991,N_2973);
and UO_422 (O_422,N_2983,N_2995);
nor UO_423 (O_423,N_2934,N_2992);
nand UO_424 (O_424,N_2989,N_2971);
nor UO_425 (O_425,N_2954,N_2904);
nor UO_426 (O_426,N_2952,N_2985);
xor UO_427 (O_427,N_2912,N_2981);
nand UO_428 (O_428,N_2913,N_2982);
nand UO_429 (O_429,N_2968,N_2916);
nand UO_430 (O_430,N_2977,N_2997);
nand UO_431 (O_431,N_2999,N_2929);
nor UO_432 (O_432,N_2906,N_2987);
nand UO_433 (O_433,N_2941,N_2989);
nand UO_434 (O_434,N_2929,N_2931);
nand UO_435 (O_435,N_2903,N_2945);
and UO_436 (O_436,N_2915,N_2984);
or UO_437 (O_437,N_2921,N_2943);
or UO_438 (O_438,N_2930,N_2980);
or UO_439 (O_439,N_2981,N_2984);
nand UO_440 (O_440,N_2987,N_2979);
or UO_441 (O_441,N_2987,N_2917);
nor UO_442 (O_442,N_2944,N_2982);
nor UO_443 (O_443,N_2989,N_2936);
or UO_444 (O_444,N_2916,N_2918);
and UO_445 (O_445,N_2922,N_2937);
and UO_446 (O_446,N_2972,N_2980);
or UO_447 (O_447,N_2960,N_2976);
and UO_448 (O_448,N_2953,N_2920);
and UO_449 (O_449,N_2901,N_2960);
nor UO_450 (O_450,N_2934,N_2996);
or UO_451 (O_451,N_2908,N_2965);
nand UO_452 (O_452,N_2992,N_2923);
nand UO_453 (O_453,N_2998,N_2930);
or UO_454 (O_454,N_2932,N_2976);
xor UO_455 (O_455,N_2932,N_2984);
or UO_456 (O_456,N_2996,N_2972);
and UO_457 (O_457,N_2915,N_2990);
and UO_458 (O_458,N_2939,N_2995);
nor UO_459 (O_459,N_2993,N_2979);
nor UO_460 (O_460,N_2985,N_2991);
xor UO_461 (O_461,N_2995,N_2961);
nor UO_462 (O_462,N_2909,N_2913);
nor UO_463 (O_463,N_2938,N_2901);
nand UO_464 (O_464,N_2917,N_2907);
nand UO_465 (O_465,N_2927,N_2916);
nand UO_466 (O_466,N_2948,N_2982);
nor UO_467 (O_467,N_2943,N_2900);
nand UO_468 (O_468,N_2984,N_2974);
and UO_469 (O_469,N_2963,N_2960);
or UO_470 (O_470,N_2998,N_2983);
and UO_471 (O_471,N_2988,N_2986);
and UO_472 (O_472,N_2918,N_2954);
and UO_473 (O_473,N_2906,N_2963);
or UO_474 (O_474,N_2999,N_2971);
or UO_475 (O_475,N_2973,N_2910);
nor UO_476 (O_476,N_2937,N_2935);
and UO_477 (O_477,N_2922,N_2974);
or UO_478 (O_478,N_2954,N_2906);
nor UO_479 (O_479,N_2910,N_2934);
xor UO_480 (O_480,N_2956,N_2936);
and UO_481 (O_481,N_2954,N_2925);
nand UO_482 (O_482,N_2924,N_2948);
nand UO_483 (O_483,N_2920,N_2931);
and UO_484 (O_484,N_2964,N_2900);
nor UO_485 (O_485,N_2921,N_2939);
or UO_486 (O_486,N_2954,N_2907);
xnor UO_487 (O_487,N_2959,N_2946);
nand UO_488 (O_488,N_2992,N_2947);
or UO_489 (O_489,N_2993,N_2974);
nor UO_490 (O_490,N_2934,N_2975);
and UO_491 (O_491,N_2909,N_2998);
or UO_492 (O_492,N_2982,N_2954);
xor UO_493 (O_493,N_2901,N_2985);
xor UO_494 (O_494,N_2979,N_2918);
and UO_495 (O_495,N_2958,N_2942);
nor UO_496 (O_496,N_2989,N_2949);
or UO_497 (O_497,N_2994,N_2957);
or UO_498 (O_498,N_2902,N_2920);
and UO_499 (O_499,N_2937,N_2913);
endmodule