module basic_1000_10000_1500_20_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_388,In_942);
nand U1 (N_1,In_825,In_225);
nor U2 (N_2,In_217,In_854);
nand U3 (N_3,In_794,In_608);
nor U4 (N_4,In_538,In_317);
nor U5 (N_5,In_630,In_656);
nor U6 (N_6,In_368,In_881);
nand U7 (N_7,In_938,In_785);
nor U8 (N_8,In_935,In_45);
nor U9 (N_9,In_232,In_112);
or U10 (N_10,In_644,In_408);
nor U11 (N_11,In_990,In_870);
nor U12 (N_12,In_985,In_426);
nor U13 (N_13,In_707,In_641);
or U14 (N_14,In_658,In_718);
nand U15 (N_15,In_47,In_552);
nor U16 (N_16,In_167,In_739);
or U17 (N_17,In_646,In_154);
nor U18 (N_18,In_254,In_163);
or U19 (N_19,In_193,In_224);
nand U20 (N_20,In_276,In_42);
nand U21 (N_21,In_671,In_149);
and U22 (N_22,In_447,In_0);
nand U23 (N_23,In_353,In_420);
nand U24 (N_24,In_151,In_141);
or U25 (N_25,In_683,In_604);
and U26 (N_26,In_863,In_356);
nor U27 (N_27,In_445,In_559);
or U28 (N_28,In_750,In_557);
or U29 (N_29,In_947,In_421);
and U30 (N_30,In_912,In_266);
nand U31 (N_31,In_34,In_511);
nor U32 (N_32,In_476,In_242);
nand U33 (N_33,In_592,In_17);
or U34 (N_34,In_313,In_335);
xnor U35 (N_35,In_410,In_439);
and U36 (N_36,In_443,In_28);
and U37 (N_37,In_13,In_312);
or U38 (N_38,In_652,In_599);
or U39 (N_39,In_324,In_689);
nor U40 (N_40,In_355,In_586);
nand U41 (N_41,In_187,In_766);
nor U42 (N_42,In_980,In_724);
nor U43 (N_43,In_855,In_301);
and U44 (N_44,In_545,In_784);
nor U45 (N_45,In_299,In_489);
nor U46 (N_46,In_648,In_591);
and U47 (N_47,In_285,In_762);
nor U48 (N_48,In_115,In_418);
nand U49 (N_49,In_73,In_199);
nand U50 (N_50,In_767,In_943);
and U51 (N_51,In_543,In_322);
and U52 (N_52,In_325,In_749);
or U53 (N_53,In_960,In_140);
and U54 (N_54,In_660,In_4);
nor U55 (N_55,In_85,In_77);
xor U56 (N_56,In_606,In_19);
or U57 (N_57,In_503,In_871);
nand U58 (N_58,In_5,In_622);
nor U59 (N_59,In_346,In_694);
and U60 (N_60,In_282,In_290);
nand U61 (N_61,In_650,In_558);
nor U62 (N_62,In_502,In_901);
or U63 (N_63,In_412,In_462);
and U64 (N_64,In_771,In_597);
xor U65 (N_65,In_130,In_835);
xnor U66 (N_66,In_508,In_348);
and U67 (N_67,In_948,In_813);
nand U68 (N_68,In_659,In_744);
nand U69 (N_69,In_603,In_968);
or U70 (N_70,In_365,In_364);
nor U71 (N_71,In_817,In_203);
and U72 (N_72,In_270,In_12);
nor U73 (N_73,In_343,In_473);
nor U74 (N_74,In_993,In_568);
or U75 (N_75,In_35,In_189);
nand U76 (N_76,In_135,In_856);
nor U77 (N_77,In_287,In_306);
nand U78 (N_78,In_915,In_676);
or U79 (N_79,In_100,In_82);
nor U80 (N_80,In_381,In_962);
nor U81 (N_81,In_207,In_878);
nor U82 (N_82,In_634,In_507);
or U83 (N_83,In_59,In_946);
and U84 (N_84,In_763,In_300);
and U85 (N_85,In_495,In_635);
or U86 (N_86,In_212,In_563);
nand U87 (N_87,In_781,In_499);
nor U88 (N_88,In_344,In_539);
and U89 (N_89,In_810,In_922);
or U90 (N_90,In_341,In_107);
or U91 (N_91,In_528,In_24);
or U92 (N_92,In_730,In_256);
or U93 (N_93,In_654,In_670);
or U94 (N_94,In_610,In_31);
xor U95 (N_95,In_778,In_743);
nand U96 (N_96,In_214,In_852);
xor U97 (N_97,In_347,In_530);
and U98 (N_98,In_433,In_99);
nor U99 (N_99,In_39,In_70);
nor U100 (N_100,In_53,In_411);
nor U101 (N_101,In_768,In_828);
or U102 (N_102,In_925,In_196);
and U103 (N_103,In_996,In_826);
nor U104 (N_104,In_936,In_847);
or U105 (N_105,In_819,In_230);
or U106 (N_106,In_640,In_564);
nand U107 (N_107,In_588,In_729);
xnor U108 (N_108,In_807,In_179);
nor U109 (N_109,In_633,In_395);
nand U110 (N_110,In_822,In_9);
nand U111 (N_111,In_468,In_406);
nor U112 (N_112,In_3,In_638);
and U113 (N_113,In_998,In_519);
and U114 (N_114,In_605,In_49);
xnor U115 (N_115,In_486,In_20);
or U116 (N_116,In_239,In_387);
or U117 (N_117,In_238,In_422);
xnor U118 (N_118,In_582,In_802);
nand U119 (N_119,In_719,In_505);
nand U120 (N_120,In_128,In_329);
nand U121 (N_121,In_772,In_970);
nand U122 (N_122,In_541,In_858);
nor U123 (N_123,In_883,In_414);
and U124 (N_124,In_715,In_704);
nand U125 (N_125,In_782,In_665);
or U126 (N_126,In_522,In_520);
nand U127 (N_127,In_271,In_367);
or U128 (N_128,In_693,In_427);
nand U129 (N_129,In_178,In_757);
nor U130 (N_130,In_165,In_832);
nand U131 (N_131,In_456,In_210);
and U132 (N_132,In_197,In_669);
nand U133 (N_133,In_288,In_245);
nor U134 (N_134,In_38,In_479);
nor U135 (N_135,In_765,In_16);
and U136 (N_136,In_567,In_303);
nand U137 (N_137,In_748,In_184);
and U138 (N_138,In_65,In_930);
and U139 (N_139,In_174,In_50);
and U140 (N_140,In_298,In_401);
nor U141 (N_141,In_352,In_231);
nand U142 (N_142,In_278,In_326);
nor U143 (N_143,In_452,In_906);
and U144 (N_144,In_399,In_553);
and U145 (N_145,In_188,In_409);
nand U146 (N_146,In_701,In_733);
nand U147 (N_147,In_916,In_872);
and U148 (N_148,In_467,In_950);
nand U149 (N_149,In_21,In_974);
or U150 (N_150,In_58,In_850);
nand U151 (N_151,In_41,In_257);
nor U152 (N_152,In_880,In_240);
nor U153 (N_153,In_517,In_655);
and U154 (N_154,In_7,In_1);
nand U155 (N_155,In_904,In_44);
nand U156 (N_156,In_809,In_376);
nor U157 (N_157,In_626,In_989);
nand U158 (N_158,In_320,In_243);
and U159 (N_159,In_860,In_492);
and U160 (N_160,In_789,In_206);
nand U161 (N_161,In_84,In_262);
nand U162 (N_162,In_80,In_562);
xnor U163 (N_163,In_125,In_192);
nand U164 (N_164,In_737,In_195);
nand U165 (N_165,In_354,In_896);
or U166 (N_166,In_653,In_350);
nand U167 (N_167,In_220,In_992);
nor U168 (N_168,In_695,In_579);
or U169 (N_169,In_818,In_751);
nor U170 (N_170,In_726,In_400);
and U171 (N_171,In_629,In_64);
nor U172 (N_172,In_675,In_758);
and U173 (N_173,In_647,In_742);
or U174 (N_174,In_155,In_919);
nand U175 (N_175,In_392,In_277);
nor U176 (N_176,In_544,In_542);
or U177 (N_177,In_865,In_685);
xor U178 (N_178,In_720,In_6);
or U179 (N_179,In_234,In_111);
or U180 (N_180,In_537,In_472);
nand U181 (N_181,In_83,In_712);
or U182 (N_182,In_803,In_910);
and U183 (N_183,In_444,In_475);
or U184 (N_184,In_645,In_815);
nand U185 (N_185,In_612,In_67);
nor U186 (N_186,In_222,In_471);
xor U187 (N_187,In_487,In_867);
nor U188 (N_188,In_194,In_183);
nand U189 (N_189,In_723,In_246);
and U190 (N_190,In_595,In_798);
nor U191 (N_191,In_459,In_569);
nand U192 (N_192,In_928,In_711);
nand U193 (N_193,In_321,In_191);
nand U194 (N_194,In_119,In_146);
and U195 (N_195,In_700,In_639);
nor U196 (N_196,In_394,In_23);
nor U197 (N_197,In_159,In_688);
nand U198 (N_198,In_390,In_580);
nor U199 (N_199,In_937,In_431);
and U200 (N_200,In_114,In_116);
or U201 (N_201,In_868,In_800);
nor U202 (N_202,In_296,In_651);
xor U203 (N_203,In_637,In_281);
and U204 (N_204,In_43,In_259);
nor U205 (N_205,In_921,In_36);
nor U206 (N_206,In_185,In_795);
or U207 (N_207,In_138,In_302);
nor U208 (N_208,In_168,In_440);
or U209 (N_209,In_846,In_811);
and U210 (N_210,In_93,In_593);
xor U211 (N_211,In_101,In_774);
and U212 (N_212,In_284,In_619);
nor U213 (N_213,In_932,In_816);
nand U214 (N_214,In_176,In_251);
nor U215 (N_215,In_535,In_864);
nor U216 (N_216,In_756,In_841);
nand U217 (N_217,In_478,In_836);
nand U218 (N_218,In_755,In_738);
and U219 (N_219,In_703,In_498);
nor U220 (N_220,In_11,In_680);
or U221 (N_221,In_859,In_370);
nor U222 (N_222,In_272,In_917);
nand U223 (N_223,In_952,In_359);
or U224 (N_224,In_265,In_741);
nand U225 (N_225,In_662,In_894);
and U226 (N_226,In_308,In_787);
nor U227 (N_227,In_790,In_86);
or U228 (N_228,In_674,In_594);
or U229 (N_229,In_63,In_903);
or U230 (N_230,In_837,In_405);
xnor U231 (N_231,In_129,In_106);
and U232 (N_232,In_263,In_229);
nand U233 (N_233,In_686,In_54);
nor U234 (N_234,In_215,In_372);
nor U235 (N_235,In_525,In_494);
xnor U236 (N_236,In_690,In_702);
nor U237 (N_237,In_485,In_382);
or U238 (N_238,In_866,In_60);
and U239 (N_239,In_839,In_792);
or U240 (N_240,In_297,In_145);
nand U241 (N_241,In_705,In_223);
nor U242 (N_242,In_967,In_14);
nor U243 (N_243,In_931,In_820);
or U244 (N_244,In_423,In_252);
and U245 (N_245,In_940,In_417);
nand U246 (N_246,In_331,In_514);
or U247 (N_247,In_746,In_150);
and U248 (N_248,In_120,In_958);
and U249 (N_249,In_74,In_158);
or U250 (N_250,In_907,In_360);
nor U251 (N_251,In_37,In_233);
nand U252 (N_252,In_337,In_428);
and U253 (N_253,In_103,In_764);
or U254 (N_254,In_736,In_975);
nor U255 (N_255,In_759,In_954);
or U256 (N_256,In_78,In_887);
or U257 (N_257,In_279,In_56);
nor U258 (N_258,In_560,In_923);
nand U259 (N_259,In_182,In_824);
nand U260 (N_260,In_779,In_170);
or U261 (N_261,In_624,In_617);
nand U262 (N_262,In_323,In_280);
or U263 (N_263,In_804,In_995);
xnor U264 (N_264,In_961,In_518);
or U265 (N_265,In_889,In_121);
or U266 (N_266,In_436,In_500);
and U267 (N_267,In_673,In_122);
xor U268 (N_268,In_441,In_814);
and U269 (N_269,In_840,In_566);
nor U270 (N_270,In_775,In_432);
or U271 (N_271,In_734,In_375);
and U272 (N_272,In_944,In_583);
and U273 (N_273,In_642,In_383);
nand U274 (N_274,In_319,In_173);
xnor U275 (N_275,In_133,In_620);
nor U276 (N_276,In_273,In_959);
nand U277 (N_277,In_117,In_777);
nor U278 (N_278,In_172,In_211);
nor U279 (N_279,In_725,In_510);
and U280 (N_280,In_536,In_219);
nor U281 (N_281,In_175,In_504);
nor U282 (N_282,In_430,In_260);
nor U283 (N_283,In_424,In_92);
and U284 (N_284,In_442,In_918);
xor U285 (N_285,In_95,In_578);
nor U286 (N_286,In_87,In_490);
and U287 (N_287,In_483,In_823);
nor U288 (N_288,In_105,In_513);
nand U289 (N_289,In_62,In_769);
nor U290 (N_290,In_732,In_349);
or U291 (N_291,In_334,In_827);
nor U292 (N_292,In_435,In_72);
xnor U293 (N_293,In_161,In_808);
xnor U294 (N_294,In_497,In_661);
and U295 (N_295,In_438,In_398);
nor U296 (N_296,In_623,In_255);
nand U297 (N_297,In_955,In_572);
and U298 (N_298,In_98,In_198);
and U299 (N_299,In_877,In_458);
nor U300 (N_300,In_523,In_351);
and U301 (N_301,In_747,In_144);
nor U302 (N_302,In_493,In_997);
nand U303 (N_303,In_988,In_470);
nor U304 (N_304,In_261,In_899);
and U305 (N_305,In_934,In_126);
xor U306 (N_306,In_909,In_68);
nor U307 (N_307,In_797,In_857);
xnor U308 (N_308,In_201,In_971);
or U309 (N_309,In_902,In_124);
nor U310 (N_310,In_831,In_27);
or U311 (N_311,In_236,In_267);
nor U312 (N_312,In_491,In_888);
or U313 (N_313,In_218,In_728);
and U314 (N_314,In_963,In_166);
and U315 (N_315,In_587,In_999);
nor U316 (N_316,In_631,In_933);
xnor U317 (N_317,In_451,In_677);
or U318 (N_318,In_241,In_806);
xor U319 (N_319,In_484,In_524);
or U320 (N_320,In_152,In_32);
and U321 (N_321,In_10,In_972);
xor U322 (N_322,In_461,In_761);
or U323 (N_323,In_799,In_793);
or U324 (N_324,In_373,In_264);
and U325 (N_325,In_136,In_76);
nand U326 (N_326,In_164,In_142);
and U327 (N_327,In_969,In_897);
nand U328 (N_328,In_407,In_735);
nand U329 (N_329,In_463,In_576);
nor U330 (N_330,In_477,In_862);
nand U331 (N_331,In_987,In_601);
nand U332 (N_332,In_891,In_118);
nand U333 (N_333,In_628,In_449);
and U334 (N_334,In_258,In_554);
nand U335 (N_335,In_228,In_466);
xnor U336 (N_336,In_632,In_253);
or U337 (N_337,In_834,In_147);
nor U338 (N_338,In_453,In_692);
nor U339 (N_339,In_316,In_534);
or U340 (N_340,In_358,In_900);
xor U341 (N_341,In_691,In_672);
or U342 (N_342,In_927,In_156);
nor U343 (N_343,In_621,In_446);
or U344 (N_344,In_851,In_908);
or U345 (N_345,In_668,In_404);
xnor U346 (N_346,In_15,In_926);
or U347 (N_347,In_550,In_327);
or U348 (N_348,In_89,In_791);
or U349 (N_349,In_310,In_190);
and U350 (N_350,In_109,In_268);
nor U351 (N_351,In_131,In_66);
nor U352 (N_352,In_708,In_796);
or U353 (N_353,In_339,In_709);
xnor U354 (N_354,In_153,In_981);
nand U355 (N_355,In_22,In_812);
and U356 (N_356,In_753,In_842);
nor U357 (N_357,In_177,In_226);
or U358 (N_358,In_55,In_314);
or U359 (N_359,In_983,In_706);
nor U360 (N_360,In_895,In_208);
nand U361 (N_361,In_636,In_25);
or U362 (N_362,In_913,In_75);
xor U363 (N_363,In_590,In_506);
nand U364 (N_364,In_283,In_786);
xor U365 (N_365,In_886,In_853);
or U366 (N_366,In_512,In_874);
and U367 (N_367,In_309,In_293);
nand U368 (N_368,In_533,In_698);
nand U369 (N_369,In_377,In_788);
nor U370 (N_370,In_571,In_664);
or U371 (N_371,In_318,In_602);
xnor U372 (N_372,In_643,In_361);
or U373 (N_373,In_269,In_911);
and U374 (N_374,In_213,In_248);
nand U375 (N_375,In_97,In_216);
or U376 (N_376,In_108,In_425);
or U377 (N_377,In_460,In_332);
nand U378 (N_378,In_385,In_46);
xor U379 (N_379,In_618,In_609);
nor U380 (N_380,In_127,In_821);
xor U381 (N_381,In_110,In_292);
and U382 (N_382,In_957,In_770);
xnor U383 (N_383,In_366,In_776);
nor U384 (N_384,In_869,In_687);
nand U385 (N_385,In_205,In_469);
or U386 (N_386,In_26,In_363);
nor U387 (N_387,In_275,In_526);
and U388 (N_388,In_682,In_879);
and U389 (N_389,In_221,In_607);
nand U390 (N_390,In_573,In_905);
nor U391 (N_391,In_362,In_966);
and U392 (N_392,In_209,In_396);
xor U393 (N_393,In_48,In_684);
and U394 (N_394,In_480,In_247);
and U395 (N_395,In_965,In_235);
and U396 (N_396,In_875,In_419);
nand U397 (N_397,In_186,In_429);
and U398 (N_398,In_596,In_890);
nor U399 (N_399,In_589,In_939);
nand U400 (N_400,In_979,In_139);
and U401 (N_401,In_978,In_876);
and U402 (N_402,In_413,In_752);
and U403 (N_403,In_379,In_949);
and U404 (N_404,In_614,In_237);
or U405 (N_405,In_556,In_305);
nor U406 (N_406,In_342,In_546);
or U407 (N_407,In_657,In_882);
and U408 (N_408,In_585,In_104);
nor U409 (N_409,In_516,In_893);
nand U410 (N_410,In_90,In_555);
nor U411 (N_411,In_102,In_171);
or U412 (N_412,In_509,In_434);
nor U413 (N_413,In_924,In_547);
and U414 (N_414,In_600,In_157);
nor U415 (N_415,In_294,In_843);
or U416 (N_416,In_338,In_973);
nand U417 (N_417,In_805,In_311);
or U418 (N_418,In_202,In_667);
nor U419 (N_419,In_540,In_96);
and U420 (N_420,In_113,In_570);
and U421 (N_421,In_951,In_204);
nor U422 (N_422,In_611,In_79);
and U423 (N_423,In_873,In_838);
nor U424 (N_424,In_717,In_666);
or U425 (N_425,In_527,In_386);
and U426 (N_426,In_465,In_501);
nor U427 (N_427,In_33,In_976);
or U428 (N_428,In_977,In_898);
nand U429 (N_429,In_389,In_391);
or U430 (N_430,In_773,In_274);
and U431 (N_431,In_953,In_956);
and U432 (N_432,In_760,In_713);
and U433 (N_433,In_181,In_829);
nor U434 (N_434,In_994,In_678);
nand U435 (N_435,In_584,In_134);
nand U436 (N_436,In_581,In_51);
nand U437 (N_437,In_548,In_450);
nor U438 (N_438,In_481,In_160);
or U439 (N_439,In_515,In_52);
or U440 (N_440,In_727,In_29);
nand U441 (N_441,In_716,In_616);
nor U442 (N_442,In_885,In_780);
xor U443 (N_443,In_696,In_455);
nor U444 (N_444,In_94,In_250);
nor U445 (N_445,In_403,In_532);
nand U446 (N_446,In_397,In_615);
nor U447 (N_447,In_137,In_577);
and U448 (N_448,In_369,In_496);
xor U449 (N_449,In_328,In_731);
and U450 (N_450,In_884,In_69);
nor U451 (N_451,In_625,In_304);
nor U452 (N_452,In_941,In_448);
or U453 (N_453,In_488,In_745);
nor U454 (N_454,In_929,In_845);
nand U455 (N_455,In_378,In_984);
nor U456 (N_456,In_357,In_699);
and U457 (N_457,In_40,In_333);
nor U458 (N_458,In_740,In_132);
nor U459 (N_459,In_180,In_991);
or U460 (N_460,In_380,In_330);
or U461 (N_461,In_200,In_315);
nand U462 (N_462,In_454,In_982);
nor U463 (N_463,In_561,In_722);
or U464 (N_464,In_91,In_340);
or U465 (N_465,In_415,In_482);
or U466 (N_466,In_371,In_521);
and U467 (N_467,In_861,In_295);
nor U468 (N_468,In_848,In_710);
nor U469 (N_469,In_437,In_575);
or U470 (N_470,In_88,In_336);
and U471 (N_471,In_61,In_162);
and U472 (N_472,In_244,In_783);
or U473 (N_473,In_345,In_289);
or U474 (N_474,In_663,In_986);
xor U475 (N_475,In_71,In_833);
nor U476 (N_476,In_531,In_551);
xor U477 (N_477,In_529,In_457);
and U478 (N_478,In_286,In_81);
nand U479 (N_479,In_57,In_892);
or U480 (N_480,In_464,In_565);
nor U481 (N_481,In_627,In_598);
nand U482 (N_482,In_681,In_474);
nor U483 (N_483,In_754,In_123);
nand U484 (N_484,In_679,In_249);
nand U485 (N_485,In_8,In_30);
or U486 (N_486,In_169,In_920);
nand U487 (N_487,In_721,In_801);
nor U488 (N_488,In_914,In_945);
and U489 (N_489,In_849,In_574);
and U490 (N_490,In_384,In_844);
nor U491 (N_491,In_830,In_714);
nand U492 (N_492,In_549,In_307);
and U493 (N_493,In_964,In_374);
nand U494 (N_494,In_649,In_613);
xnor U495 (N_495,In_697,In_227);
or U496 (N_496,In_291,In_148);
or U497 (N_497,In_416,In_2);
xnor U498 (N_498,In_18,In_143);
nor U499 (N_499,In_393,In_402);
xor U500 (N_500,N_116,N_435);
nand U501 (N_501,N_374,N_307);
and U502 (N_502,N_295,N_174);
xnor U503 (N_503,N_100,N_384);
xnor U504 (N_504,N_346,N_277);
nand U505 (N_505,N_305,N_468);
xor U506 (N_506,N_272,N_281);
nand U507 (N_507,N_254,N_43);
nand U508 (N_508,N_492,N_368);
xnor U509 (N_509,N_38,N_469);
or U510 (N_510,N_178,N_162);
nor U511 (N_511,N_21,N_355);
and U512 (N_512,N_407,N_101);
and U513 (N_513,N_484,N_20);
nor U514 (N_514,N_133,N_460);
and U515 (N_515,N_62,N_17);
or U516 (N_516,N_70,N_59);
and U517 (N_517,N_488,N_392);
nor U518 (N_518,N_191,N_112);
nand U519 (N_519,N_389,N_247);
nand U520 (N_520,N_163,N_290);
nor U521 (N_521,N_436,N_126);
nor U522 (N_522,N_98,N_202);
and U523 (N_523,N_314,N_496);
and U524 (N_524,N_422,N_379);
nor U525 (N_525,N_218,N_118);
and U526 (N_526,N_83,N_84);
nand U527 (N_527,N_275,N_63);
and U528 (N_528,N_471,N_217);
and U529 (N_529,N_61,N_244);
and U530 (N_530,N_317,N_56);
nor U531 (N_531,N_69,N_320);
or U532 (N_532,N_497,N_110);
nand U533 (N_533,N_181,N_297);
xor U534 (N_534,N_366,N_204);
nor U535 (N_535,N_145,N_196);
or U536 (N_536,N_113,N_457);
or U537 (N_537,N_296,N_219);
nand U538 (N_538,N_71,N_300);
xor U539 (N_539,N_65,N_425);
nor U540 (N_540,N_159,N_37);
and U541 (N_541,N_25,N_340);
and U542 (N_542,N_10,N_333);
nor U543 (N_543,N_195,N_115);
nor U544 (N_544,N_462,N_283);
or U545 (N_545,N_7,N_380);
nor U546 (N_546,N_417,N_171);
and U547 (N_547,N_149,N_326);
and U548 (N_548,N_201,N_28);
and U549 (N_549,N_109,N_255);
nor U550 (N_550,N_136,N_2);
and U551 (N_551,N_334,N_416);
or U552 (N_552,N_243,N_73);
or U553 (N_553,N_426,N_120);
or U554 (N_554,N_117,N_401);
or U555 (N_555,N_12,N_321);
and U556 (N_556,N_257,N_421);
nor U557 (N_557,N_106,N_31);
or U558 (N_558,N_128,N_206);
or U559 (N_559,N_342,N_68);
or U560 (N_560,N_456,N_213);
nor U561 (N_561,N_499,N_242);
or U562 (N_562,N_66,N_198);
nor U563 (N_563,N_441,N_424);
or U564 (N_564,N_104,N_375);
nor U565 (N_565,N_208,N_194);
and U566 (N_566,N_23,N_48);
and U567 (N_567,N_382,N_144);
nor U568 (N_568,N_413,N_27);
nor U569 (N_569,N_14,N_315);
nor U570 (N_570,N_430,N_483);
or U571 (N_571,N_209,N_197);
and U572 (N_572,N_312,N_179);
nor U573 (N_573,N_177,N_415);
nand U574 (N_574,N_428,N_474);
nor U575 (N_575,N_13,N_353);
and U576 (N_576,N_267,N_122);
and U577 (N_577,N_214,N_388);
nor U578 (N_578,N_367,N_36);
or U579 (N_579,N_9,N_432);
or U580 (N_580,N_184,N_400);
xnor U581 (N_581,N_154,N_402);
or U582 (N_582,N_103,N_261);
or U583 (N_583,N_107,N_124);
and U584 (N_584,N_481,N_319);
nor U585 (N_585,N_292,N_18);
and U586 (N_586,N_470,N_294);
and U587 (N_587,N_211,N_180);
xor U588 (N_588,N_466,N_454);
nor U589 (N_589,N_91,N_495);
and U590 (N_590,N_373,N_155);
nand U591 (N_591,N_35,N_238);
or U592 (N_592,N_278,N_491);
and U593 (N_593,N_97,N_11);
nand U594 (N_594,N_114,N_308);
nor U595 (N_595,N_349,N_448);
or U596 (N_596,N_186,N_207);
and U597 (N_597,N_146,N_357);
nor U598 (N_598,N_166,N_395);
nand U599 (N_599,N_350,N_192);
and U600 (N_600,N_390,N_47);
xor U601 (N_601,N_233,N_472);
and U602 (N_602,N_486,N_249);
nor U603 (N_603,N_264,N_399);
nor U604 (N_604,N_111,N_173);
nor U605 (N_605,N_182,N_311);
and U606 (N_606,N_253,N_444);
nand U607 (N_607,N_289,N_442);
xor U608 (N_608,N_405,N_434);
nor U609 (N_609,N_121,N_323);
nand U610 (N_610,N_51,N_376);
nand U611 (N_611,N_99,N_33);
xor U612 (N_612,N_158,N_190);
nand U613 (N_613,N_22,N_485);
and U614 (N_614,N_493,N_306);
and U615 (N_615,N_282,N_408);
xnor U616 (N_616,N_125,N_200);
and U617 (N_617,N_414,N_352);
xor U618 (N_618,N_193,N_372);
xor U619 (N_619,N_246,N_386);
nand U620 (N_620,N_269,N_30);
xor U621 (N_621,N_445,N_139);
nand U622 (N_622,N_330,N_67);
nand U623 (N_623,N_140,N_236);
or U624 (N_624,N_227,N_147);
and U625 (N_625,N_271,N_138);
or U626 (N_626,N_237,N_221);
and U627 (N_627,N_362,N_298);
nand U628 (N_628,N_49,N_438);
nor U629 (N_629,N_170,N_64);
xor U630 (N_630,N_303,N_224);
or U631 (N_631,N_90,N_1);
and U632 (N_632,N_383,N_250);
and U633 (N_633,N_40,N_148);
nor U634 (N_634,N_239,N_279);
nor U635 (N_635,N_354,N_54);
and U636 (N_636,N_331,N_248);
and U637 (N_637,N_370,N_260);
nand U638 (N_638,N_187,N_6);
and U639 (N_639,N_364,N_322);
or U640 (N_640,N_336,N_26);
or U641 (N_641,N_398,N_8);
nor U642 (N_642,N_262,N_153);
nand U643 (N_643,N_397,N_108);
or U644 (N_644,N_284,N_387);
or U645 (N_645,N_119,N_325);
nor U646 (N_646,N_189,N_19);
nor U647 (N_647,N_345,N_175);
xor U648 (N_648,N_285,N_229);
or U649 (N_649,N_365,N_151);
or U650 (N_650,N_385,N_404);
or U651 (N_651,N_188,N_301);
nand U652 (N_652,N_487,N_406);
nor U653 (N_653,N_453,N_419);
nor U654 (N_654,N_409,N_134);
xnor U655 (N_655,N_475,N_433);
or U656 (N_656,N_479,N_164);
and U657 (N_657,N_465,N_216);
nor U658 (N_658,N_286,N_332);
nand U659 (N_659,N_280,N_215);
nor U660 (N_660,N_412,N_143);
nand U661 (N_661,N_45,N_228);
nand U662 (N_662,N_420,N_287);
or U663 (N_663,N_489,N_161);
or U664 (N_664,N_449,N_338);
or U665 (N_665,N_427,N_266);
nand U666 (N_666,N_396,N_32);
or U667 (N_667,N_473,N_498);
or U668 (N_668,N_235,N_127);
nand U669 (N_669,N_81,N_41);
nor U670 (N_670,N_24,N_172);
or U671 (N_671,N_351,N_361);
and U672 (N_672,N_268,N_480);
nand U673 (N_673,N_309,N_381);
nor U674 (N_674,N_310,N_150);
or U675 (N_675,N_410,N_288);
xor U676 (N_676,N_57,N_299);
nand U677 (N_677,N_89,N_74);
or U678 (N_678,N_39,N_34);
or U679 (N_679,N_431,N_132);
nor U680 (N_680,N_86,N_476);
or U681 (N_681,N_92,N_358);
nand U682 (N_682,N_165,N_15);
and U683 (N_683,N_58,N_42);
xor U684 (N_684,N_220,N_259);
nand U685 (N_685,N_87,N_94);
xor U686 (N_686,N_156,N_276);
xor U687 (N_687,N_418,N_141);
and U688 (N_688,N_450,N_256);
nand U689 (N_689,N_347,N_359);
nor U690 (N_690,N_339,N_348);
xnor U691 (N_691,N_318,N_77);
nand U692 (N_692,N_490,N_212);
nand U693 (N_693,N_169,N_273);
nand U694 (N_694,N_459,N_222);
and U695 (N_695,N_93,N_225);
and U696 (N_696,N_245,N_356);
nand U697 (N_697,N_393,N_304);
nand U698 (N_698,N_78,N_46);
or U699 (N_699,N_88,N_185);
and U700 (N_700,N_241,N_291);
nand U701 (N_701,N_265,N_464);
nor U702 (N_702,N_270,N_29);
and U703 (N_703,N_203,N_439);
nor U704 (N_704,N_210,N_455);
and U705 (N_705,N_461,N_95);
and U706 (N_706,N_50,N_263);
nand U707 (N_707,N_157,N_377);
and U708 (N_708,N_60,N_429);
xnor U709 (N_709,N_160,N_316);
nand U710 (N_710,N_52,N_360);
xor U711 (N_711,N_458,N_44);
and U712 (N_712,N_0,N_76);
and U713 (N_713,N_3,N_440);
or U714 (N_714,N_176,N_80);
nand U715 (N_715,N_199,N_223);
and U716 (N_716,N_478,N_343);
nor U717 (N_717,N_168,N_463);
xnor U718 (N_718,N_226,N_230);
nand U719 (N_719,N_327,N_131);
nand U720 (N_720,N_75,N_234);
and U721 (N_721,N_403,N_123);
nor U722 (N_722,N_205,N_82);
nor U723 (N_723,N_16,N_137);
nand U724 (N_724,N_344,N_258);
and U725 (N_725,N_85,N_4);
and U726 (N_726,N_313,N_105);
and U727 (N_727,N_494,N_72);
and U728 (N_728,N_129,N_240);
nand U729 (N_729,N_102,N_55);
and U730 (N_730,N_130,N_329);
nand U731 (N_731,N_371,N_274);
nand U732 (N_732,N_53,N_167);
or U733 (N_733,N_363,N_467);
nand U734 (N_734,N_337,N_394);
nand U735 (N_735,N_391,N_423);
or U736 (N_736,N_447,N_252);
nand U737 (N_737,N_446,N_378);
or U738 (N_738,N_142,N_335);
or U739 (N_739,N_302,N_451);
nor U740 (N_740,N_135,N_232);
nor U741 (N_741,N_5,N_482);
xor U742 (N_742,N_96,N_293);
nand U743 (N_743,N_341,N_369);
or U744 (N_744,N_452,N_324);
nor U745 (N_745,N_152,N_79);
or U746 (N_746,N_328,N_231);
and U747 (N_747,N_443,N_183);
or U748 (N_748,N_411,N_477);
nand U749 (N_749,N_437,N_251);
xor U750 (N_750,N_372,N_235);
or U751 (N_751,N_17,N_431);
nor U752 (N_752,N_212,N_306);
nand U753 (N_753,N_128,N_68);
or U754 (N_754,N_393,N_21);
nor U755 (N_755,N_326,N_12);
nand U756 (N_756,N_432,N_471);
and U757 (N_757,N_64,N_80);
or U758 (N_758,N_39,N_288);
xor U759 (N_759,N_20,N_272);
nand U760 (N_760,N_25,N_122);
nor U761 (N_761,N_67,N_369);
or U762 (N_762,N_63,N_137);
nand U763 (N_763,N_242,N_337);
nor U764 (N_764,N_455,N_378);
nor U765 (N_765,N_300,N_414);
nor U766 (N_766,N_149,N_192);
xnor U767 (N_767,N_114,N_96);
or U768 (N_768,N_386,N_418);
or U769 (N_769,N_272,N_443);
and U770 (N_770,N_95,N_418);
and U771 (N_771,N_411,N_414);
and U772 (N_772,N_391,N_294);
nand U773 (N_773,N_73,N_186);
or U774 (N_774,N_31,N_73);
xor U775 (N_775,N_427,N_111);
nand U776 (N_776,N_104,N_278);
nor U777 (N_777,N_208,N_15);
xnor U778 (N_778,N_134,N_298);
nor U779 (N_779,N_441,N_187);
and U780 (N_780,N_95,N_465);
nand U781 (N_781,N_268,N_192);
xnor U782 (N_782,N_257,N_197);
nor U783 (N_783,N_54,N_275);
or U784 (N_784,N_180,N_421);
nand U785 (N_785,N_91,N_218);
or U786 (N_786,N_409,N_260);
nor U787 (N_787,N_443,N_34);
and U788 (N_788,N_223,N_348);
nor U789 (N_789,N_224,N_356);
nor U790 (N_790,N_130,N_365);
and U791 (N_791,N_290,N_94);
and U792 (N_792,N_91,N_54);
or U793 (N_793,N_355,N_461);
nand U794 (N_794,N_89,N_423);
nand U795 (N_795,N_217,N_414);
nor U796 (N_796,N_34,N_483);
xnor U797 (N_797,N_449,N_308);
nand U798 (N_798,N_330,N_28);
or U799 (N_799,N_79,N_292);
nor U800 (N_800,N_94,N_313);
nand U801 (N_801,N_101,N_465);
and U802 (N_802,N_88,N_496);
nor U803 (N_803,N_385,N_40);
nor U804 (N_804,N_192,N_120);
and U805 (N_805,N_111,N_48);
and U806 (N_806,N_317,N_158);
or U807 (N_807,N_71,N_106);
or U808 (N_808,N_25,N_222);
nor U809 (N_809,N_443,N_436);
nor U810 (N_810,N_461,N_186);
nor U811 (N_811,N_493,N_55);
nand U812 (N_812,N_423,N_82);
xor U813 (N_813,N_216,N_87);
nor U814 (N_814,N_311,N_409);
nand U815 (N_815,N_81,N_367);
nor U816 (N_816,N_177,N_137);
nand U817 (N_817,N_282,N_434);
nor U818 (N_818,N_331,N_235);
and U819 (N_819,N_36,N_91);
nand U820 (N_820,N_198,N_306);
nor U821 (N_821,N_153,N_196);
or U822 (N_822,N_218,N_285);
or U823 (N_823,N_271,N_309);
xor U824 (N_824,N_414,N_83);
and U825 (N_825,N_119,N_264);
and U826 (N_826,N_168,N_39);
nor U827 (N_827,N_194,N_321);
and U828 (N_828,N_447,N_335);
xnor U829 (N_829,N_365,N_354);
nand U830 (N_830,N_384,N_354);
nand U831 (N_831,N_474,N_383);
xor U832 (N_832,N_117,N_193);
nand U833 (N_833,N_376,N_248);
or U834 (N_834,N_40,N_313);
xor U835 (N_835,N_335,N_22);
or U836 (N_836,N_482,N_132);
nand U837 (N_837,N_302,N_37);
nand U838 (N_838,N_69,N_285);
nand U839 (N_839,N_424,N_232);
nor U840 (N_840,N_406,N_158);
or U841 (N_841,N_460,N_450);
xnor U842 (N_842,N_94,N_225);
and U843 (N_843,N_493,N_301);
or U844 (N_844,N_312,N_487);
or U845 (N_845,N_109,N_218);
nor U846 (N_846,N_144,N_246);
nor U847 (N_847,N_438,N_266);
nand U848 (N_848,N_63,N_471);
and U849 (N_849,N_414,N_119);
nor U850 (N_850,N_211,N_101);
nand U851 (N_851,N_347,N_403);
or U852 (N_852,N_245,N_62);
nor U853 (N_853,N_423,N_254);
or U854 (N_854,N_110,N_9);
and U855 (N_855,N_395,N_379);
xor U856 (N_856,N_176,N_475);
nand U857 (N_857,N_30,N_448);
nand U858 (N_858,N_277,N_244);
nand U859 (N_859,N_422,N_369);
or U860 (N_860,N_154,N_136);
nor U861 (N_861,N_39,N_272);
nor U862 (N_862,N_424,N_461);
xor U863 (N_863,N_204,N_451);
nand U864 (N_864,N_33,N_158);
nand U865 (N_865,N_301,N_135);
nor U866 (N_866,N_287,N_498);
or U867 (N_867,N_171,N_467);
nor U868 (N_868,N_105,N_137);
nand U869 (N_869,N_92,N_340);
or U870 (N_870,N_361,N_242);
xnor U871 (N_871,N_209,N_429);
nor U872 (N_872,N_323,N_245);
nand U873 (N_873,N_170,N_475);
nand U874 (N_874,N_160,N_131);
or U875 (N_875,N_218,N_190);
nor U876 (N_876,N_260,N_219);
xnor U877 (N_877,N_291,N_382);
nor U878 (N_878,N_108,N_103);
nand U879 (N_879,N_85,N_431);
nand U880 (N_880,N_13,N_316);
and U881 (N_881,N_133,N_157);
xnor U882 (N_882,N_225,N_17);
nor U883 (N_883,N_186,N_201);
nand U884 (N_884,N_238,N_205);
or U885 (N_885,N_66,N_241);
xnor U886 (N_886,N_277,N_487);
nor U887 (N_887,N_239,N_162);
nor U888 (N_888,N_35,N_36);
nand U889 (N_889,N_158,N_227);
nor U890 (N_890,N_381,N_158);
nor U891 (N_891,N_233,N_239);
nand U892 (N_892,N_249,N_150);
and U893 (N_893,N_145,N_96);
or U894 (N_894,N_253,N_200);
nor U895 (N_895,N_110,N_204);
nor U896 (N_896,N_399,N_464);
nor U897 (N_897,N_64,N_77);
nor U898 (N_898,N_312,N_238);
nor U899 (N_899,N_175,N_150);
or U900 (N_900,N_52,N_329);
and U901 (N_901,N_13,N_391);
and U902 (N_902,N_111,N_8);
or U903 (N_903,N_440,N_266);
xnor U904 (N_904,N_87,N_361);
nand U905 (N_905,N_246,N_433);
xnor U906 (N_906,N_190,N_257);
and U907 (N_907,N_12,N_202);
or U908 (N_908,N_378,N_95);
and U909 (N_909,N_296,N_88);
nor U910 (N_910,N_13,N_362);
nor U911 (N_911,N_59,N_281);
nor U912 (N_912,N_215,N_462);
nand U913 (N_913,N_54,N_408);
or U914 (N_914,N_438,N_429);
nor U915 (N_915,N_308,N_103);
and U916 (N_916,N_481,N_161);
nand U917 (N_917,N_331,N_385);
nand U918 (N_918,N_258,N_32);
and U919 (N_919,N_149,N_470);
or U920 (N_920,N_90,N_439);
nor U921 (N_921,N_452,N_365);
nand U922 (N_922,N_16,N_167);
or U923 (N_923,N_292,N_154);
nand U924 (N_924,N_109,N_415);
or U925 (N_925,N_336,N_47);
or U926 (N_926,N_289,N_213);
or U927 (N_927,N_382,N_4);
or U928 (N_928,N_91,N_65);
or U929 (N_929,N_340,N_77);
nor U930 (N_930,N_175,N_201);
nor U931 (N_931,N_311,N_217);
xnor U932 (N_932,N_345,N_78);
or U933 (N_933,N_161,N_356);
nand U934 (N_934,N_317,N_241);
nor U935 (N_935,N_58,N_104);
or U936 (N_936,N_112,N_16);
nand U937 (N_937,N_436,N_243);
xor U938 (N_938,N_43,N_42);
and U939 (N_939,N_214,N_95);
and U940 (N_940,N_484,N_345);
nand U941 (N_941,N_466,N_51);
nor U942 (N_942,N_25,N_187);
and U943 (N_943,N_141,N_459);
and U944 (N_944,N_221,N_309);
nor U945 (N_945,N_10,N_338);
or U946 (N_946,N_337,N_282);
nor U947 (N_947,N_150,N_491);
nor U948 (N_948,N_130,N_192);
and U949 (N_949,N_56,N_81);
nand U950 (N_950,N_450,N_167);
xnor U951 (N_951,N_1,N_444);
nand U952 (N_952,N_163,N_335);
or U953 (N_953,N_69,N_180);
nand U954 (N_954,N_285,N_237);
and U955 (N_955,N_469,N_69);
nand U956 (N_956,N_23,N_273);
nand U957 (N_957,N_445,N_475);
and U958 (N_958,N_100,N_319);
and U959 (N_959,N_483,N_363);
nand U960 (N_960,N_343,N_216);
nor U961 (N_961,N_498,N_277);
nand U962 (N_962,N_226,N_144);
and U963 (N_963,N_286,N_451);
and U964 (N_964,N_391,N_314);
xnor U965 (N_965,N_362,N_464);
nor U966 (N_966,N_475,N_252);
nor U967 (N_967,N_337,N_135);
nor U968 (N_968,N_143,N_98);
nor U969 (N_969,N_472,N_42);
xnor U970 (N_970,N_212,N_125);
nand U971 (N_971,N_495,N_466);
or U972 (N_972,N_90,N_142);
or U973 (N_973,N_273,N_396);
nor U974 (N_974,N_137,N_266);
nand U975 (N_975,N_293,N_406);
xnor U976 (N_976,N_470,N_357);
nor U977 (N_977,N_346,N_278);
nor U978 (N_978,N_134,N_293);
xnor U979 (N_979,N_498,N_429);
or U980 (N_980,N_428,N_450);
or U981 (N_981,N_267,N_36);
nor U982 (N_982,N_374,N_335);
nand U983 (N_983,N_114,N_379);
or U984 (N_984,N_470,N_20);
nand U985 (N_985,N_329,N_398);
or U986 (N_986,N_91,N_217);
nand U987 (N_987,N_98,N_5);
nand U988 (N_988,N_39,N_258);
nor U989 (N_989,N_58,N_186);
nor U990 (N_990,N_181,N_385);
or U991 (N_991,N_302,N_147);
or U992 (N_992,N_383,N_185);
nand U993 (N_993,N_174,N_258);
nor U994 (N_994,N_106,N_185);
nand U995 (N_995,N_72,N_245);
nor U996 (N_996,N_37,N_275);
nor U997 (N_997,N_189,N_42);
nand U998 (N_998,N_359,N_207);
nor U999 (N_999,N_102,N_72);
nor U1000 (N_1000,N_622,N_795);
nand U1001 (N_1001,N_843,N_882);
nand U1002 (N_1002,N_776,N_830);
xnor U1003 (N_1003,N_608,N_835);
nand U1004 (N_1004,N_904,N_563);
and U1005 (N_1005,N_662,N_560);
nor U1006 (N_1006,N_848,N_510);
nand U1007 (N_1007,N_894,N_568);
nor U1008 (N_1008,N_587,N_586);
xnor U1009 (N_1009,N_967,N_565);
xnor U1010 (N_1010,N_825,N_867);
nand U1011 (N_1011,N_858,N_881);
or U1012 (N_1012,N_599,N_654);
nand U1013 (N_1013,N_679,N_935);
and U1014 (N_1014,N_781,N_819);
nand U1015 (N_1015,N_520,N_911);
and U1016 (N_1016,N_986,N_585);
nor U1017 (N_1017,N_692,N_580);
or U1018 (N_1018,N_548,N_899);
or U1019 (N_1019,N_746,N_878);
nor U1020 (N_1020,N_539,N_783);
and U1021 (N_1021,N_600,N_612);
nand U1022 (N_1022,N_515,N_811);
and U1023 (N_1023,N_860,N_922);
nand U1024 (N_1024,N_556,N_616);
and U1025 (N_1025,N_660,N_755);
nor U1026 (N_1026,N_834,N_710);
nand U1027 (N_1027,N_863,N_553);
or U1028 (N_1028,N_809,N_552);
nor U1029 (N_1029,N_509,N_827);
nand U1030 (N_1030,N_963,N_674);
nor U1031 (N_1031,N_775,N_978);
nor U1032 (N_1032,N_764,N_651);
nand U1033 (N_1033,N_540,N_532);
or U1034 (N_1034,N_877,N_750);
or U1035 (N_1035,N_980,N_788);
nor U1036 (N_1036,N_533,N_595);
and U1037 (N_1037,N_665,N_803);
nand U1038 (N_1038,N_886,N_939);
and U1039 (N_1039,N_626,N_772);
and U1040 (N_1040,N_852,N_559);
nand U1041 (N_1041,N_909,N_603);
and U1042 (N_1042,N_845,N_999);
nor U1043 (N_1043,N_945,N_932);
nor U1044 (N_1044,N_791,N_928);
nand U1045 (N_1045,N_885,N_957);
xnor U1046 (N_1046,N_927,N_859);
nand U1047 (N_1047,N_681,N_972);
and U1048 (N_1048,N_814,N_657);
nand U1049 (N_1049,N_544,N_584);
xnor U1050 (N_1050,N_862,N_645);
and U1051 (N_1051,N_569,N_546);
xor U1052 (N_1052,N_673,N_638);
or U1053 (N_1053,N_865,N_832);
or U1054 (N_1054,N_870,N_854);
and U1055 (N_1055,N_912,N_817);
nand U1056 (N_1056,N_683,N_954);
and U1057 (N_1057,N_601,N_677);
and U1058 (N_1058,N_916,N_505);
or U1059 (N_1059,N_784,N_947);
nand U1060 (N_1060,N_526,N_695);
nor U1061 (N_1061,N_652,N_678);
nand U1062 (N_1062,N_786,N_979);
nor U1063 (N_1063,N_659,N_970);
nor U1064 (N_1064,N_523,N_690);
nor U1065 (N_1065,N_613,N_846);
and U1066 (N_1066,N_663,N_557);
and U1067 (N_1067,N_634,N_716);
and U1068 (N_1068,N_706,N_807);
nor U1069 (N_1069,N_768,N_770);
or U1070 (N_1070,N_721,N_696);
and U1071 (N_1071,N_876,N_769);
xor U1072 (N_1072,N_524,N_842);
nor U1073 (N_1073,N_961,N_729);
and U1074 (N_1074,N_996,N_880);
nand U1075 (N_1075,N_794,N_658);
nand U1076 (N_1076,N_531,N_720);
or U1077 (N_1077,N_888,N_938);
nand U1078 (N_1078,N_680,N_512);
or U1079 (N_1079,N_550,N_572);
and U1080 (N_1080,N_530,N_968);
or U1081 (N_1081,N_748,N_596);
nand U1082 (N_1082,N_627,N_682);
xnor U1083 (N_1083,N_715,N_558);
or U1084 (N_1084,N_619,N_933);
and U1085 (N_1085,N_661,N_797);
or U1086 (N_1086,N_982,N_751);
nand U1087 (N_1087,N_773,N_883);
nand U1088 (N_1088,N_734,N_931);
nand U1089 (N_1089,N_805,N_889);
nor U1090 (N_1090,N_921,N_753);
or U1091 (N_1091,N_749,N_983);
nand U1092 (N_1092,N_702,N_636);
nand U1093 (N_1093,N_871,N_823);
nand U1094 (N_1094,N_735,N_966);
nand U1095 (N_1095,N_762,N_977);
nand U1096 (N_1096,N_920,N_676);
nand U1097 (N_1097,N_956,N_822);
and U1098 (N_1098,N_994,N_637);
or U1099 (N_1099,N_849,N_617);
nand U1100 (N_1100,N_856,N_536);
nor U1101 (N_1101,N_703,N_688);
and U1102 (N_1102,N_527,N_718);
nand U1103 (N_1103,N_732,N_610);
or U1104 (N_1104,N_714,N_522);
or U1105 (N_1105,N_529,N_625);
or U1106 (N_1106,N_779,N_988);
nor U1107 (N_1107,N_561,N_730);
and U1108 (N_1108,N_606,N_908);
and U1109 (N_1109,N_653,N_955);
nand U1110 (N_1110,N_974,N_841);
nand U1111 (N_1111,N_687,N_949);
and U1112 (N_1112,N_689,N_892);
nor U1113 (N_1113,N_694,N_618);
or U1114 (N_1114,N_723,N_629);
nor U1115 (N_1115,N_738,N_853);
nand U1116 (N_1116,N_975,N_541);
and U1117 (N_1117,N_969,N_712);
or U1118 (N_1118,N_576,N_675);
or U1119 (N_1119,N_850,N_808);
or U1120 (N_1120,N_942,N_829);
nor U1121 (N_1121,N_693,N_727);
or U1122 (N_1122,N_826,N_635);
and U1123 (N_1123,N_567,N_806);
nand U1124 (N_1124,N_836,N_833);
xor U1125 (N_1125,N_759,N_643);
nand U1126 (N_1126,N_630,N_951);
and U1127 (N_1127,N_936,N_519);
xnor U1128 (N_1128,N_989,N_571);
nor U1129 (N_1129,N_760,N_873);
or U1130 (N_1130,N_670,N_992);
or U1131 (N_1131,N_668,N_960);
and U1132 (N_1132,N_581,N_549);
and U1133 (N_1133,N_778,N_930);
or U1134 (N_1134,N_941,N_708);
and U1135 (N_1135,N_838,N_582);
nand U1136 (N_1136,N_731,N_861);
nor U1137 (N_1137,N_518,N_538);
and U1138 (N_1138,N_801,N_649);
nand U1139 (N_1139,N_684,N_840);
nor U1140 (N_1140,N_711,N_700);
and U1141 (N_1141,N_562,N_551);
nand U1142 (N_1142,N_516,N_664);
or U1143 (N_1143,N_981,N_820);
and U1144 (N_1144,N_868,N_780);
nand U1145 (N_1145,N_993,N_574);
nand U1146 (N_1146,N_644,N_914);
xnor U1147 (N_1147,N_901,N_985);
or U1148 (N_1148,N_542,N_667);
nor U1149 (N_1149,N_761,N_802);
and U1150 (N_1150,N_507,N_605);
and U1151 (N_1151,N_705,N_879);
xnor U1152 (N_1152,N_624,N_611);
and U1153 (N_1153,N_952,N_573);
or U1154 (N_1154,N_591,N_609);
xnor U1155 (N_1155,N_646,N_895);
and U1156 (N_1156,N_953,N_621);
or U1157 (N_1157,N_698,N_719);
nand U1158 (N_1158,N_948,N_525);
nor U1159 (N_1159,N_984,N_815);
and U1160 (N_1160,N_508,N_647);
nand U1161 (N_1161,N_771,N_796);
and U1162 (N_1162,N_672,N_787);
nand U1163 (N_1163,N_891,N_650);
or U1164 (N_1164,N_570,N_500);
or U1165 (N_1165,N_813,N_633);
or U1166 (N_1166,N_566,N_890);
nor U1167 (N_1167,N_866,N_839);
nor U1168 (N_1168,N_857,N_579);
nor U1169 (N_1169,N_593,N_594);
and U1170 (N_1170,N_875,N_864);
and U1171 (N_1171,N_937,N_816);
nand U1172 (N_1172,N_925,N_722);
and U1173 (N_1173,N_717,N_792);
or U1174 (N_1174,N_824,N_583);
nor U1175 (N_1175,N_513,N_614);
and U1176 (N_1176,N_940,N_905);
xor U1177 (N_1177,N_631,N_906);
or U1178 (N_1178,N_514,N_590);
nand U1179 (N_1179,N_812,N_589);
nand U1180 (N_1180,N_987,N_944);
and U1181 (N_1181,N_884,N_628);
xnor U1182 (N_1182,N_503,N_733);
nor U1183 (N_1183,N_704,N_554);
nor U1184 (N_1184,N_521,N_758);
nand U1185 (N_1185,N_902,N_555);
or U1186 (N_1186,N_893,N_724);
and U1187 (N_1187,N_785,N_897);
or U1188 (N_1188,N_766,N_763);
nand U1189 (N_1189,N_793,N_537);
and U1190 (N_1190,N_950,N_639);
nand U1191 (N_1191,N_887,N_837);
xnor U1192 (N_1192,N_697,N_995);
nand U1193 (N_1193,N_666,N_818);
xnor U1194 (N_1194,N_898,N_973);
and U1195 (N_1195,N_543,N_501);
or U1196 (N_1196,N_741,N_725);
and U1197 (N_1197,N_640,N_804);
nor U1198 (N_1198,N_745,N_799);
or U1199 (N_1199,N_965,N_913);
nor U1200 (N_1200,N_844,N_896);
nor U1201 (N_1201,N_752,N_789);
and U1202 (N_1202,N_774,N_641);
nor U1203 (N_1203,N_828,N_713);
or U1204 (N_1204,N_997,N_943);
and U1205 (N_1205,N_685,N_900);
or U1206 (N_1206,N_598,N_777);
xnor U1207 (N_1207,N_847,N_991);
or U1208 (N_1208,N_655,N_648);
nor U1209 (N_1209,N_756,N_757);
or U1210 (N_1210,N_872,N_821);
nand U1211 (N_1211,N_528,N_669);
and U1212 (N_1212,N_604,N_535);
nor U1213 (N_1213,N_737,N_918);
or U1214 (N_1214,N_767,N_709);
nor U1215 (N_1215,N_686,N_874);
or U1216 (N_1216,N_926,N_511);
nor U1217 (N_1217,N_736,N_588);
nand U1218 (N_1218,N_740,N_592);
and U1219 (N_1219,N_578,N_726);
and U1220 (N_1220,N_575,N_504);
and U1221 (N_1221,N_642,N_701);
nor U1222 (N_1222,N_998,N_597);
and U1223 (N_1223,N_934,N_547);
xnor U1224 (N_1224,N_707,N_958);
nand U1225 (N_1225,N_728,N_671);
nand U1226 (N_1226,N_747,N_923);
nand U1227 (N_1227,N_656,N_502);
and U1228 (N_1228,N_506,N_855);
or U1229 (N_1229,N_765,N_623);
nand U1230 (N_1230,N_615,N_632);
or U1231 (N_1231,N_800,N_534);
nand U1232 (N_1232,N_903,N_971);
and U1233 (N_1233,N_782,N_564);
and U1234 (N_1234,N_915,N_620);
xor U1235 (N_1235,N_754,N_976);
xor U1236 (N_1236,N_959,N_742);
nand U1237 (N_1237,N_517,N_831);
xor U1238 (N_1238,N_946,N_607);
or U1239 (N_1239,N_810,N_929);
and U1240 (N_1240,N_739,N_798);
or U1241 (N_1241,N_545,N_964);
nand U1242 (N_1242,N_577,N_691);
nor U1243 (N_1243,N_990,N_699);
nor U1244 (N_1244,N_790,N_869);
nor U1245 (N_1245,N_910,N_851);
nor U1246 (N_1246,N_744,N_924);
and U1247 (N_1247,N_917,N_907);
and U1248 (N_1248,N_602,N_962);
or U1249 (N_1249,N_919,N_743);
nor U1250 (N_1250,N_614,N_774);
or U1251 (N_1251,N_578,N_706);
nand U1252 (N_1252,N_784,N_909);
nor U1253 (N_1253,N_636,N_612);
and U1254 (N_1254,N_531,N_897);
nand U1255 (N_1255,N_558,N_889);
and U1256 (N_1256,N_580,N_659);
nand U1257 (N_1257,N_502,N_693);
and U1258 (N_1258,N_983,N_685);
or U1259 (N_1259,N_843,N_923);
nand U1260 (N_1260,N_981,N_597);
and U1261 (N_1261,N_523,N_902);
nand U1262 (N_1262,N_668,N_685);
nor U1263 (N_1263,N_915,N_695);
nor U1264 (N_1264,N_554,N_675);
nand U1265 (N_1265,N_519,N_723);
xor U1266 (N_1266,N_622,N_791);
nand U1267 (N_1267,N_780,N_698);
nand U1268 (N_1268,N_653,N_961);
nand U1269 (N_1269,N_814,N_987);
nand U1270 (N_1270,N_504,N_999);
nor U1271 (N_1271,N_823,N_676);
nand U1272 (N_1272,N_839,N_777);
or U1273 (N_1273,N_773,N_754);
nand U1274 (N_1274,N_587,N_717);
or U1275 (N_1275,N_585,N_575);
nor U1276 (N_1276,N_797,N_992);
and U1277 (N_1277,N_638,N_688);
nand U1278 (N_1278,N_798,N_916);
and U1279 (N_1279,N_604,N_864);
nor U1280 (N_1280,N_561,N_611);
nor U1281 (N_1281,N_810,N_757);
nor U1282 (N_1282,N_690,N_667);
nor U1283 (N_1283,N_741,N_819);
or U1284 (N_1284,N_916,N_709);
and U1285 (N_1285,N_796,N_629);
and U1286 (N_1286,N_502,N_757);
or U1287 (N_1287,N_519,N_904);
nand U1288 (N_1288,N_617,N_577);
and U1289 (N_1289,N_698,N_625);
or U1290 (N_1290,N_875,N_944);
and U1291 (N_1291,N_801,N_553);
nor U1292 (N_1292,N_569,N_638);
nor U1293 (N_1293,N_740,N_984);
nand U1294 (N_1294,N_940,N_966);
nor U1295 (N_1295,N_721,N_546);
nor U1296 (N_1296,N_790,N_570);
and U1297 (N_1297,N_961,N_574);
nor U1298 (N_1298,N_944,N_598);
or U1299 (N_1299,N_909,N_872);
nor U1300 (N_1300,N_907,N_966);
and U1301 (N_1301,N_612,N_690);
and U1302 (N_1302,N_578,N_559);
and U1303 (N_1303,N_712,N_709);
nor U1304 (N_1304,N_540,N_527);
or U1305 (N_1305,N_639,N_735);
nor U1306 (N_1306,N_998,N_644);
or U1307 (N_1307,N_530,N_822);
and U1308 (N_1308,N_763,N_889);
nand U1309 (N_1309,N_823,N_562);
nor U1310 (N_1310,N_868,N_747);
nand U1311 (N_1311,N_896,N_819);
and U1312 (N_1312,N_920,N_554);
and U1313 (N_1313,N_670,N_508);
and U1314 (N_1314,N_906,N_575);
and U1315 (N_1315,N_659,N_876);
and U1316 (N_1316,N_740,N_685);
or U1317 (N_1317,N_592,N_715);
nor U1318 (N_1318,N_984,N_500);
and U1319 (N_1319,N_508,N_700);
nand U1320 (N_1320,N_910,N_661);
nor U1321 (N_1321,N_578,N_871);
or U1322 (N_1322,N_515,N_925);
or U1323 (N_1323,N_604,N_853);
or U1324 (N_1324,N_539,N_808);
or U1325 (N_1325,N_658,N_585);
nor U1326 (N_1326,N_640,N_729);
nor U1327 (N_1327,N_601,N_639);
nand U1328 (N_1328,N_644,N_543);
nand U1329 (N_1329,N_661,N_857);
or U1330 (N_1330,N_517,N_808);
nor U1331 (N_1331,N_593,N_952);
nand U1332 (N_1332,N_806,N_922);
nand U1333 (N_1333,N_640,N_644);
nand U1334 (N_1334,N_997,N_823);
or U1335 (N_1335,N_543,N_726);
and U1336 (N_1336,N_696,N_731);
nand U1337 (N_1337,N_783,N_863);
nand U1338 (N_1338,N_651,N_756);
or U1339 (N_1339,N_935,N_616);
or U1340 (N_1340,N_574,N_944);
nor U1341 (N_1341,N_501,N_866);
or U1342 (N_1342,N_780,N_590);
and U1343 (N_1343,N_515,N_600);
nand U1344 (N_1344,N_872,N_753);
or U1345 (N_1345,N_591,N_544);
and U1346 (N_1346,N_661,N_985);
and U1347 (N_1347,N_701,N_991);
and U1348 (N_1348,N_815,N_747);
xnor U1349 (N_1349,N_711,N_924);
nor U1350 (N_1350,N_781,N_665);
nor U1351 (N_1351,N_754,N_608);
nor U1352 (N_1352,N_579,N_668);
and U1353 (N_1353,N_893,N_910);
and U1354 (N_1354,N_599,N_590);
and U1355 (N_1355,N_977,N_988);
and U1356 (N_1356,N_979,N_663);
and U1357 (N_1357,N_747,N_837);
or U1358 (N_1358,N_580,N_920);
nor U1359 (N_1359,N_565,N_961);
and U1360 (N_1360,N_749,N_501);
and U1361 (N_1361,N_775,N_867);
nor U1362 (N_1362,N_933,N_991);
or U1363 (N_1363,N_588,N_876);
nor U1364 (N_1364,N_663,N_579);
or U1365 (N_1365,N_845,N_834);
and U1366 (N_1366,N_701,N_973);
xnor U1367 (N_1367,N_867,N_568);
and U1368 (N_1368,N_591,N_717);
nand U1369 (N_1369,N_508,N_942);
and U1370 (N_1370,N_553,N_731);
or U1371 (N_1371,N_555,N_867);
nand U1372 (N_1372,N_901,N_540);
nand U1373 (N_1373,N_799,N_649);
nor U1374 (N_1374,N_560,N_713);
xor U1375 (N_1375,N_542,N_985);
and U1376 (N_1376,N_641,N_732);
xor U1377 (N_1377,N_762,N_560);
nand U1378 (N_1378,N_677,N_888);
xor U1379 (N_1379,N_641,N_960);
nand U1380 (N_1380,N_543,N_987);
nand U1381 (N_1381,N_538,N_710);
and U1382 (N_1382,N_905,N_968);
or U1383 (N_1383,N_560,N_702);
nor U1384 (N_1384,N_840,N_616);
nand U1385 (N_1385,N_562,N_978);
and U1386 (N_1386,N_704,N_987);
nor U1387 (N_1387,N_509,N_669);
or U1388 (N_1388,N_506,N_778);
nor U1389 (N_1389,N_777,N_905);
or U1390 (N_1390,N_837,N_774);
and U1391 (N_1391,N_804,N_797);
nand U1392 (N_1392,N_910,N_830);
and U1393 (N_1393,N_642,N_602);
xor U1394 (N_1394,N_823,N_520);
xnor U1395 (N_1395,N_571,N_927);
nand U1396 (N_1396,N_774,N_693);
and U1397 (N_1397,N_966,N_911);
nand U1398 (N_1398,N_689,N_548);
and U1399 (N_1399,N_769,N_513);
and U1400 (N_1400,N_590,N_535);
or U1401 (N_1401,N_982,N_796);
xor U1402 (N_1402,N_716,N_937);
or U1403 (N_1403,N_616,N_944);
and U1404 (N_1404,N_622,N_947);
nand U1405 (N_1405,N_804,N_535);
nor U1406 (N_1406,N_719,N_795);
nor U1407 (N_1407,N_530,N_877);
xnor U1408 (N_1408,N_801,N_703);
or U1409 (N_1409,N_515,N_756);
and U1410 (N_1410,N_575,N_842);
or U1411 (N_1411,N_559,N_771);
and U1412 (N_1412,N_785,N_696);
nor U1413 (N_1413,N_754,N_741);
and U1414 (N_1414,N_697,N_652);
nand U1415 (N_1415,N_979,N_558);
nand U1416 (N_1416,N_626,N_730);
and U1417 (N_1417,N_652,N_515);
and U1418 (N_1418,N_716,N_616);
nand U1419 (N_1419,N_992,N_710);
nor U1420 (N_1420,N_600,N_980);
and U1421 (N_1421,N_829,N_909);
xnor U1422 (N_1422,N_793,N_758);
nand U1423 (N_1423,N_715,N_839);
nor U1424 (N_1424,N_710,N_855);
or U1425 (N_1425,N_765,N_608);
or U1426 (N_1426,N_586,N_602);
and U1427 (N_1427,N_967,N_897);
nand U1428 (N_1428,N_696,N_592);
or U1429 (N_1429,N_647,N_857);
or U1430 (N_1430,N_538,N_827);
and U1431 (N_1431,N_771,N_709);
xor U1432 (N_1432,N_627,N_666);
nor U1433 (N_1433,N_676,N_821);
or U1434 (N_1434,N_797,N_860);
or U1435 (N_1435,N_711,N_768);
nand U1436 (N_1436,N_934,N_844);
nor U1437 (N_1437,N_614,N_984);
or U1438 (N_1438,N_830,N_914);
or U1439 (N_1439,N_533,N_904);
nor U1440 (N_1440,N_590,N_554);
nor U1441 (N_1441,N_928,N_862);
and U1442 (N_1442,N_627,N_619);
or U1443 (N_1443,N_592,N_875);
or U1444 (N_1444,N_667,N_665);
nand U1445 (N_1445,N_725,N_914);
or U1446 (N_1446,N_679,N_568);
or U1447 (N_1447,N_890,N_998);
or U1448 (N_1448,N_659,N_915);
or U1449 (N_1449,N_871,N_876);
nand U1450 (N_1450,N_833,N_793);
xnor U1451 (N_1451,N_608,N_874);
or U1452 (N_1452,N_822,N_839);
and U1453 (N_1453,N_829,N_581);
nand U1454 (N_1454,N_674,N_897);
or U1455 (N_1455,N_731,N_848);
nand U1456 (N_1456,N_664,N_705);
and U1457 (N_1457,N_965,N_991);
or U1458 (N_1458,N_939,N_802);
or U1459 (N_1459,N_773,N_868);
and U1460 (N_1460,N_729,N_775);
or U1461 (N_1461,N_722,N_669);
xor U1462 (N_1462,N_556,N_734);
and U1463 (N_1463,N_596,N_590);
nand U1464 (N_1464,N_666,N_751);
or U1465 (N_1465,N_762,N_985);
nor U1466 (N_1466,N_758,N_573);
or U1467 (N_1467,N_946,N_512);
xor U1468 (N_1468,N_916,N_539);
nor U1469 (N_1469,N_838,N_892);
nor U1470 (N_1470,N_575,N_734);
or U1471 (N_1471,N_707,N_594);
nand U1472 (N_1472,N_732,N_701);
nor U1473 (N_1473,N_955,N_665);
and U1474 (N_1474,N_753,N_682);
nor U1475 (N_1475,N_984,N_957);
and U1476 (N_1476,N_647,N_755);
or U1477 (N_1477,N_879,N_865);
nand U1478 (N_1478,N_867,N_855);
nand U1479 (N_1479,N_989,N_553);
nand U1480 (N_1480,N_915,N_709);
or U1481 (N_1481,N_741,N_912);
nand U1482 (N_1482,N_941,N_680);
and U1483 (N_1483,N_585,N_509);
nand U1484 (N_1484,N_921,N_648);
and U1485 (N_1485,N_769,N_780);
and U1486 (N_1486,N_538,N_949);
nand U1487 (N_1487,N_975,N_837);
nand U1488 (N_1488,N_660,N_876);
nand U1489 (N_1489,N_832,N_789);
or U1490 (N_1490,N_925,N_629);
nand U1491 (N_1491,N_530,N_935);
and U1492 (N_1492,N_924,N_791);
or U1493 (N_1493,N_502,N_575);
and U1494 (N_1494,N_770,N_773);
nand U1495 (N_1495,N_880,N_750);
nor U1496 (N_1496,N_633,N_518);
and U1497 (N_1497,N_779,N_865);
nor U1498 (N_1498,N_872,N_962);
nor U1499 (N_1499,N_823,N_675);
and U1500 (N_1500,N_1051,N_1405);
and U1501 (N_1501,N_1333,N_1287);
or U1502 (N_1502,N_1323,N_1207);
and U1503 (N_1503,N_1200,N_1156);
and U1504 (N_1504,N_1292,N_1437);
and U1505 (N_1505,N_1003,N_1093);
or U1506 (N_1506,N_1109,N_1188);
nand U1507 (N_1507,N_1225,N_1144);
nand U1508 (N_1508,N_1103,N_1083);
nand U1509 (N_1509,N_1414,N_1187);
and U1510 (N_1510,N_1384,N_1340);
or U1511 (N_1511,N_1234,N_1043);
or U1512 (N_1512,N_1171,N_1190);
xnor U1513 (N_1513,N_1382,N_1272);
and U1514 (N_1514,N_1220,N_1249);
and U1515 (N_1515,N_1029,N_1360);
xor U1516 (N_1516,N_1367,N_1129);
or U1517 (N_1517,N_1152,N_1242);
and U1518 (N_1518,N_1130,N_1185);
and U1519 (N_1519,N_1448,N_1320);
and U1520 (N_1520,N_1010,N_1373);
nand U1521 (N_1521,N_1175,N_1270);
nand U1522 (N_1522,N_1022,N_1316);
nand U1523 (N_1523,N_1324,N_1229);
or U1524 (N_1524,N_1160,N_1069);
nand U1525 (N_1525,N_1217,N_1192);
and U1526 (N_1526,N_1304,N_1247);
nor U1527 (N_1527,N_1193,N_1283);
nor U1528 (N_1528,N_1426,N_1232);
nand U1529 (N_1529,N_1053,N_1334);
nor U1530 (N_1530,N_1268,N_1298);
and U1531 (N_1531,N_1063,N_1494);
nand U1532 (N_1532,N_1168,N_1045);
or U1533 (N_1533,N_1449,N_1089);
nand U1534 (N_1534,N_1203,N_1356);
or U1535 (N_1535,N_1418,N_1110);
or U1536 (N_1536,N_1409,N_1269);
nor U1537 (N_1537,N_1224,N_1216);
nor U1538 (N_1538,N_1050,N_1098);
nand U1539 (N_1539,N_1398,N_1389);
and U1540 (N_1540,N_1173,N_1201);
nand U1541 (N_1541,N_1372,N_1472);
and U1542 (N_1542,N_1136,N_1084);
or U1543 (N_1543,N_1261,N_1302);
nor U1544 (N_1544,N_1181,N_1231);
xnor U1545 (N_1545,N_1042,N_1403);
nor U1546 (N_1546,N_1289,N_1064);
nand U1547 (N_1547,N_1466,N_1362);
nor U1548 (N_1548,N_1195,N_1191);
nand U1549 (N_1549,N_1295,N_1417);
nor U1550 (N_1550,N_1422,N_1401);
and U1551 (N_1551,N_1392,N_1067);
nand U1552 (N_1552,N_1251,N_1213);
and U1553 (N_1553,N_1391,N_1014);
nor U1554 (N_1554,N_1206,N_1421);
nand U1555 (N_1555,N_1151,N_1178);
or U1556 (N_1556,N_1236,N_1434);
nand U1557 (N_1557,N_1126,N_1480);
or U1558 (N_1558,N_1039,N_1090);
or U1559 (N_1559,N_1326,N_1467);
xor U1560 (N_1560,N_1143,N_1263);
and U1561 (N_1561,N_1104,N_1423);
and U1562 (N_1562,N_1149,N_1106);
nor U1563 (N_1563,N_1363,N_1278);
nor U1564 (N_1564,N_1141,N_1256);
nand U1565 (N_1565,N_1390,N_1112);
nor U1566 (N_1566,N_1393,N_1325);
nand U1567 (N_1567,N_1101,N_1313);
or U1568 (N_1568,N_1006,N_1118);
nand U1569 (N_1569,N_1315,N_1442);
nor U1570 (N_1570,N_1239,N_1273);
nand U1571 (N_1571,N_1179,N_1164);
nor U1572 (N_1572,N_1317,N_1469);
nand U1573 (N_1573,N_1489,N_1461);
nor U1574 (N_1574,N_1365,N_1154);
nand U1575 (N_1575,N_1343,N_1400);
and U1576 (N_1576,N_1476,N_1092);
xnor U1577 (N_1577,N_1018,N_1412);
xnor U1578 (N_1578,N_1411,N_1265);
nor U1579 (N_1579,N_1176,N_1194);
or U1580 (N_1580,N_1385,N_1000);
and U1581 (N_1581,N_1337,N_1075);
and U1582 (N_1582,N_1493,N_1237);
nor U1583 (N_1583,N_1495,N_1311);
and U1584 (N_1584,N_1172,N_1055);
or U1585 (N_1585,N_1303,N_1379);
nand U1586 (N_1586,N_1037,N_1416);
and U1587 (N_1587,N_1452,N_1338);
xnor U1588 (N_1588,N_1142,N_1458);
or U1589 (N_1589,N_1020,N_1281);
and U1590 (N_1590,N_1297,N_1031);
nor U1591 (N_1591,N_1453,N_1262);
or U1592 (N_1592,N_1222,N_1105);
xor U1593 (N_1593,N_1062,N_1026);
nand U1594 (N_1594,N_1254,N_1087);
or U1595 (N_1595,N_1041,N_1027);
xor U1596 (N_1596,N_1072,N_1184);
xnor U1597 (N_1597,N_1139,N_1397);
and U1598 (N_1598,N_1204,N_1413);
or U1599 (N_1599,N_1260,N_1059);
and U1600 (N_1600,N_1358,N_1369);
nand U1601 (N_1601,N_1294,N_1341);
nor U1602 (N_1602,N_1219,N_1161);
nand U1603 (N_1603,N_1257,N_1076);
and U1604 (N_1604,N_1347,N_1475);
and U1605 (N_1605,N_1212,N_1486);
nand U1606 (N_1606,N_1034,N_1377);
nor U1607 (N_1607,N_1276,N_1081);
xor U1608 (N_1608,N_1399,N_1307);
xor U1609 (N_1609,N_1459,N_1226);
xnor U1610 (N_1610,N_1345,N_1396);
xnor U1611 (N_1611,N_1432,N_1335);
nand U1612 (N_1612,N_1487,N_1049);
xor U1613 (N_1613,N_1035,N_1210);
nand U1614 (N_1614,N_1128,N_1366);
nand U1615 (N_1615,N_1158,N_1196);
xnor U1616 (N_1616,N_1140,N_1074);
xor U1617 (N_1617,N_1424,N_1114);
and U1618 (N_1618,N_1174,N_1275);
nor U1619 (N_1619,N_1001,N_1197);
nand U1620 (N_1620,N_1351,N_1479);
and U1621 (N_1621,N_1013,N_1430);
or U1622 (N_1622,N_1127,N_1070);
nand U1623 (N_1623,N_1402,N_1293);
nor U1624 (N_1624,N_1056,N_1305);
nor U1625 (N_1625,N_1032,N_1123);
or U1626 (N_1626,N_1435,N_1167);
nand U1627 (N_1627,N_1025,N_1394);
nand U1628 (N_1628,N_1364,N_1387);
nand U1629 (N_1629,N_1182,N_1198);
or U1630 (N_1630,N_1329,N_1355);
nand U1631 (N_1631,N_1162,N_1497);
and U1632 (N_1632,N_1327,N_1485);
and U1633 (N_1633,N_1073,N_1071);
nand U1634 (N_1634,N_1102,N_1211);
nand U1635 (N_1635,N_1359,N_1290);
nand U1636 (N_1636,N_1177,N_1223);
xnor U1637 (N_1637,N_1410,N_1443);
xnor U1638 (N_1638,N_1146,N_1153);
or U1639 (N_1639,N_1267,N_1438);
nand U1640 (N_1640,N_1135,N_1133);
and U1641 (N_1641,N_1244,N_1166);
nand U1642 (N_1642,N_1131,N_1054);
and U1643 (N_1643,N_1012,N_1002);
and U1644 (N_1644,N_1271,N_1250);
nor U1645 (N_1645,N_1150,N_1238);
and U1646 (N_1646,N_1455,N_1404);
or U1647 (N_1647,N_1044,N_1499);
nor U1648 (N_1648,N_1374,N_1255);
nand U1649 (N_1649,N_1248,N_1202);
or U1650 (N_1650,N_1309,N_1330);
and U1651 (N_1651,N_1004,N_1339);
nand U1652 (N_1652,N_1066,N_1318);
nand U1653 (N_1653,N_1441,N_1077);
nor U1654 (N_1654,N_1286,N_1028);
nand U1655 (N_1655,N_1117,N_1348);
and U1656 (N_1656,N_1446,N_1350);
nor U1657 (N_1657,N_1147,N_1008);
or U1658 (N_1658,N_1462,N_1368);
nor U1659 (N_1659,N_1218,N_1331);
nand U1660 (N_1660,N_1189,N_1282);
nor U1661 (N_1661,N_1395,N_1259);
and U1662 (N_1662,N_1180,N_1241);
and U1663 (N_1663,N_1148,N_1230);
nor U1664 (N_1664,N_1353,N_1408);
nand U1665 (N_1665,N_1228,N_1371);
and U1666 (N_1666,N_1447,N_1381);
nor U1667 (N_1667,N_1097,N_1021);
and U1668 (N_1668,N_1484,N_1068);
nand U1669 (N_1669,N_1100,N_1376);
and U1670 (N_1670,N_1085,N_1252);
xor U1671 (N_1671,N_1346,N_1415);
nor U1672 (N_1672,N_1058,N_1349);
or U1673 (N_1673,N_1163,N_1464);
nor U1674 (N_1674,N_1233,N_1157);
or U1675 (N_1675,N_1291,N_1322);
and U1676 (N_1676,N_1496,N_1159);
xor U1677 (N_1677,N_1492,N_1111);
nor U1678 (N_1678,N_1047,N_1122);
xor U1679 (N_1679,N_1091,N_1312);
nand U1680 (N_1680,N_1407,N_1082);
or U1681 (N_1681,N_1186,N_1431);
nor U1682 (N_1682,N_1386,N_1456);
and U1683 (N_1683,N_1099,N_1245);
and U1684 (N_1684,N_1375,N_1488);
nor U1685 (N_1685,N_1080,N_1288);
nand U1686 (N_1686,N_1095,N_1454);
nor U1687 (N_1687,N_1215,N_1011);
nand U1688 (N_1688,N_1119,N_1429);
nor U1689 (N_1689,N_1296,N_1451);
nand U1690 (N_1690,N_1209,N_1457);
or U1691 (N_1691,N_1208,N_1046);
xor U1692 (N_1692,N_1113,N_1354);
nor U1693 (N_1693,N_1477,N_1380);
and U1694 (N_1694,N_1439,N_1199);
nor U1695 (N_1695,N_1036,N_1450);
and U1696 (N_1696,N_1310,N_1057);
xor U1697 (N_1697,N_1427,N_1266);
nor U1698 (N_1698,N_1246,N_1406);
and U1699 (N_1699,N_1378,N_1306);
and U1700 (N_1700,N_1352,N_1033);
and U1701 (N_1701,N_1125,N_1370);
and U1702 (N_1702,N_1332,N_1319);
nor U1703 (N_1703,N_1023,N_1498);
and U1704 (N_1704,N_1078,N_1328);
nor U1705 (N_1705,N_1468,N_1460);
nand U1706 (N_1706,N_1301,N_1165);
xor U1707 (N_1707,N_1015,N_1471);
or U1708 (N_1708,N_1463,N_1108);
or U1709 (N_1709,N_1361,N_1065);
xor U1710 (N_1710,N_1264,N_1444);
nand U1711 (N_1711,N_1470,N_1284);
nand U1712 (N_1712,N_1321,N_1240);
nand U1713 (N_1713,N_1005,N_1425);
and U1714 (N_1714,N_1478,N_1024);
or U1715 (N_1715,N_1107,N_1274);
or U1716 (N_1716,N_1383,N_1483);
or U1717 (N_1717,N_1227,N_1243);
or U1718 (N_1718,N_1019,N_1124);
or U1719 (N_1719,N_1481,N_1145);
nand U1720 (N_1720,N_1253,N_1342);
or U1721 (N_1721,N_1060,N_1205);
or U1722 (N_1722,N_1088,N_1183);
and U1723 (N_1723,N_1440,N_1115);
and U1724 (N_1724,N_1314,N_1048);
and U1725 (N_1725,N_1336,N_1096);
and U1726 (N_1726,N_1079,N_1473);
or U1727 (N_1727,N_1436,N_1445);
nand U1728 (N_1728,N_1285,N_1137);
or U1729 (N_1729,N_1121,N_1061);
nand U1730 (N_1730,N_1009,N_1017);
or U1731 (N_1731,N_1116,N_1134);
nor U1732 (N_1732,N_1214,N_1465);
and U1733 (N_1733,N_1120,N_1308);
nand U1734 (N_1734,N_1138,N_1490);
nand U1735 (N_1735,N_1491,N_1279);
and U1736 (N_1736,N_1277,N_1007);
and U1737 (N_1737,N_1170,N_1235);
and U1738 (N_1738,N_1482,N_1433);
nor U1739 (N_1739,N_1258,N_1357);
xor U1740 (N_1740,N_1094,N_1052);
nor U1741 (N_1741,N_1344,N_1419);
nor U1742 (N_1742,N_1420,N_1169);
or U1743 (N_1743,N_1040,N_1155);
or U1744 (N_1744,N_1474,N_1388);
or U1745 (N_1745,N_1016,N_1299);
nand U1746 (N_1746,N_1132,N_1300);
nand U1747 (N_1747,N_1280,N_1221);
or U1748 (N_1748,N_1086,N_1428);
nor U1749 (N_1749,N_1038,N_1030);
nor U1750 (N_1750,N_1444,N_1421);
nor U1751 (N_1751,N_1034,N_1425);
and U1752 (N_1752,N_1267,N_1154);
nor U1753 (N_1753,N_1045,N_1414);
nand U1754 (N_1754,N_1269,N_1344);
nor U1755 (N_1755,N_1150,N_1314);
nand U1756 (N_1756,N_1498,N_1062);
and U1757 (N_1757,N_1212,N_1446);
or U1758 (N_1758,N_1429,N_1329);
nand U1759 (N_1759,N_1304,N_1224);
nor U1760 (N_1760,N_1495,N_1302);
nand U1761 (N_1761,N_1296,N_1415);
or U1762 (N_1762,N_1230,N_1209);
or U1763 (N_1763,N_1472,N_1214);
nand U1764 (N_1764,N_1205,N_1351);
nand U1765 (N_1765,N_1000,N_1046);
nor U1766 (N_1766,N_1448,N_1199);
and U1767 (N_1767,N_1177,N_1228);
and U1768 (N_1768,N_1195,N_1338);
nand U1769 (N_1769,N_1221,N_1064);
xor U1770 (N_1770,N_1182,N_1332);
or U1771 (N_1771,N_1292,N_1389);
nor U1772 (N_1772,N_1417,N_1444);
nor U1773 (N_1773,N_1313,N_1355);
or U1774 (N_1774,N_1467,N_1084);
nand U1775 (N_1775,N_1344,N_1171);
and U1776 (N_1776,N_1424,N_1383);
nor U1777 (N_1777,N_1333,N_1203);
and U1778 (N_1778,N_1263,N_1165);
nand U1779 (N_1779,N_1470,N_1229);
and U1780 (N_1780,N_1250,N_1405);
nor U1781 (N_1781,N_1168,N_1016);
nand U1782 (N_1782,N_1428,N_1313);
or U1783 (N_1783,N_1368,N_1355);
or U1784 (N_1784,N_1353,N_1301);
nor U1785 (N_1785,N_1466,N_1496);
and U1786 (N_1786,N_1238,N_1396);
nor U1787 (N_1787,N_1034,N_1171);
and U1788 (N_1788,N_1233,N_1461);
nand U1789 (N_1789,N_1306,N_1179);
or U1790 (N_1790,N_1231,N_1227);
nor U1791 (N_1791,N_1283,N_1044);
and U1792 (N_1792,N_1262,N_1334);
xor U1793 (N_1793,N_1132,N_1039);
and U1794 (N_1794,N_1069,N_1120);
nor U1795 (N_1795,N_1463,N_1124);
or U1796 (N_1796,N_1119,N_1364);
or U1797 (N_1797,N_1368,N_1067);
nor U1798 (N_1798,N_1447,N_1251);
nor U1799 (N_1799,N_1218,N_1347);
nand U1800 (N_1800,N_1222,N_1417);
nand U1801 (N_1801,N_1347,N_1110);
nor U1802 (N_1802,N_1018,N_1230);
and U1803 (N_1803,N_1043,N_1056);
xor U1804 (N_1804,N_1270,N_1295);
nand U1805 (N_1805,N_1373,N_1283);
or U1806 (N_1806,N_1374,N_1059);
nand U1807 (N_1807,N_1365,N_1354);
nor U1808 (N_1808,N_1315,N_1021);
nor U1809 (N_1809,N_1181,N_1215);
and U1810 (N_1810,N_1216,N_1065);
and U1811 (N_1811,N_1178,N_1154);
and U1812 (N_1812,N_1310,N_1268);
or U1813 (N_1813,N_1161,N_1378);
nor U1814 (N_1814,N_1476,N_1083);
xor U1815 (N_1815,N_1212,N_1305);
nand U1816 (N_1816,N_1264,N_1436);
nand U1817 (N_1817,N_1220,N_1286);
nor U1818 (N_1818,N_1349,N_1422);
nand U1819 (N_1819,N_1048,N_1102);
or U1820 (N_1820,N_1351,N_1208);
nand U1821 (N_1821,N_1157,N_1402);
or U1822 (N_1822,N_1190,N_1174);
or U1823 (N_1823,N_1494,N_1440);
and U1824 (N_1824,N_1218,N_1314);
or U1825 (N_1825,N_1485,N_1075);
xor U1826 (N_1826,N_1435,N_1011);
or U1827 (N_1827,N_1172,N_1355);
or U1828 (N_1828,N_1078,N_1142);
and U1829 (N_1829,N_1161,N_1380);
and U1830 (N_1830,N_1231,N_1489);
nor U1831 (N_1831,N_1479,N_1281);
nand U1832 (N_1832,N_1149,N_1071);
or U1833 (N_1833,N_1197,N_1258);
nor U1834 (N_1834,N_1424,N_1224);
and U1835 (N_1835,N_1226,N_1372);
and U1836 (N_1836,N_1042,N_1266);
and U1837 (N_1837,N_1064,N_1150);
or U1838 (N_1838,N_1164,N_1122);
or U1839 (N_1839,N_1203,N_1384);
nand U1840 (N_1840,N_1180,N_1186);
nor U1841 (N_1841,N_1145,N_1043);
nor U1842 (N_1842,N_1446,N_1330);
nor U1843 (N_1843,N_1079,N_1378);
and U1844 (N_1844,N_1230,N_1043);
and U1845 (N_1845,N_1478,N_1073);
or U1846 (N_1846,N_1089,N_1241);
and U1847 (N_1847,N_1399,N_1326);
nand U1848 (N_1848,N_1336,N_1281);
nand U1849 (N_1849,N_1163,N_1483);
nor U1850 (N_1850,N_1132,N_1424);
xor U1851 (N_1851,N_1067,N_1037);
xnor U1852 (N_1852,N_1322,N_1249);
nor U1853 (N_1853,N_1078,N_1169);
and U1854 (N_1854,N_1326,N_1216);
or U1855 (N_1855,N_1469,N_1115);
or U1856 (N_1856,N_1250,N_1105);
or U1857 (N_1857,N_1336,N_1008);
xor U1858 (N_1858,N_1167,N_1090);
or U1859 (N_1859,N_1446,N_1217);
or U1860 (N_1860,N_1184,N_1169);
and U1861 (N_1861,N_1003,N_1312);
and U1862 (N_1862,N_1346,N_1352);
and U1863 (N_1863,N_1278,N_1396);
and U1864 (N_1864,N_1075,N_1036);
or U1865 (N_1865,N_1369,N_1495);
or U1866 (N_1866,N_1208,N_1268);
or U1867 (N_1867,N_1417,N_1475);
nor U1868 (N_1868,N_1499,N_1351);
xor U1869 (N_1869,N_1366,N_1293);
and U1870 (N_1870,N_1336,N_1261);
nor U1871 (N_1871,N_1489,N_1476);
and U1872 (N_1872,N_1041,N_1363);
nor U1873 (N_1873,N_1417,N_1259);
nor U1874 (N_1874,N_1333,N_1340);
nor U1875 (N_1875,N_1041,N_1383);
or U1876 (N_1876,N_1394,N_1303);
nand U1877 (N_1877,N_1489,N_1360);
and U1878 (N_1878,N_1076,N_1249);
nor U1879 (N_1879,N_1236,N_1362);
and U1880 (N_1880,N_1382,N_1407);
and U1881 (N_1881,N_1370,N_1026);
nor U1882 (N_1882,N_1420,N_1406);
or U1883 (N_1883,N_1028,N_1252);
nor U1884 (N_1884,N_1179,N_1131);
nand U1885 (N_1885,N_1120,N_1494);
nand U1886 (N_1886,N_1257,N_1083);
and U1887 (N_1887,N_1394,N_1495);
or U1888 (N_1888,N_1492,N_1467);
or U1889 (N_1889,N_1207,N_1401);
xor U1890 (N_1890,N_1226,N_1480);
or U1891 (N_1891,N_1204,N_1257);
nand U1892 (N_1892,N_1362,N_1205);
nand U1893 (N_1893,N_1032,N_1193);
nor U1894 (N_1894,N_1395,N_1355);
xnor U1895 (N_1895,N_1300,N_1360);
or U1896 (N_1896,N_1368,N_1326);
and U1897 (N_1897,N_1100,N_1218);
or U1898 (N_1898,N_1157,N_1381);
nand U1899 (N_1899,N_1035,N_1132);
nand U1900 (N_1900,N_1146,N_1355);
nor U1901 (N_1901,N_1465,N_1423);
nand U1902 (N_1902,N_1442,N_1140);
nor U1903 (N_1903,N_1430,N_1257);
or U1904 (N_1904,N_1153,N_1117);
or U1905 (N_1905,N_1388,N_1081);
and U1906 (N_1906,N_1323,N_1353);
nor U1907 (N_1907,N_1242,N_1376);
nand U1908 (N_1908,N_1404,N_1247);
and U1909 (N_1909,N_1102,N_1208);
and U1910 (N_1910,N_1357,N_1000);
or U1911 (N_1911,N_1414,N_1011);
or U1912 (N_1912,N_1378,N_1096);
and U1913 (N_1913,N_1254,N_1411);
xor U1914 (N_1914,N_1459,N_1452);
nor U1915 (N_1915,N_1024,N_1023);
or U1916 (N_1916,N_1040,N_1216);
nor U1917 (N_1917,N_1342,N_1118);
or U1918 (N_1918,N_1434,N_1029);
nor U1919 (N_1919,N_1456,N_1046);
nand U1920 (N_1920,N_1233,N_1154);
or U1921 (N_1921,N_1128,N_1362);
nor U1922 (N_1922,N_1491,N_1063);
and U1923 (N_1923,N_1299,N_1209);
xnor U1924 (N_1924,N_1321,N_1478);
and U1925 (N_1925,N_1012,N_1366);
or U1926 (N_1926,N_1188,N_1142);
and U1927 (N_1927,N_1074,N_1274);
xnor U1928 (N_1928,N_1422,N_1297);
nand U1929 (N_1929,N_1362,N_1417);
nor U1930 (N_1930,N_1387,N_1385);
nand U1931 (N_1931,N_1150,N_1121);
or U1932 (N_1932,N_1181,N_1108);
and U1933 (N_1933,N_1420,N_1283);
and U1934 (N_1934,N_1063,N_1184);
nor U1935 (N_1935,N_1479,N_1425);
nand U1936 (N_1936,N_1353,N_1123);
nand U1937 (N_1937,N_1237,N_1219);
nand U1938 (N_1938,N_1034,N_1167);
and U1939 (N_1939,N_1350,N_1258);
or U1940 (N_1940,N_1198,N_1158);
xnor U1941 (N_1941,N_1169,N_1323);
nand U1942 (N_1942,N_1008,N_1107);
nor U1943 (N_1943,N_1298,N_1318);
nand U1944 (N_1944,N_1219,N_1148);
or U1945 (N_1945,N_1460,N_1040);
nand U1946 (N_1946,N_1006,N_1125);
and U1947 (N_1947,N_1181,N_1450);
and U1948 (N_1948,N_1049,N_1433);
or U1949 (N_1949,N_1388,N_1273);
xor U1950 (N_1950,N_1459,N_1023);
nor U1951 (N_1951,N_1356,N_1182);
or U1952 (N_1952,N_1251,N_1422);
or U1953 (N_1953,N_1483,N_1295);
xnor U1954 (N_1954,N_1221,N_1490);
or U1955 (N_1955,N_1002,N_1470);
and U1956 (N_1956,N_1172,N_1485);
nor U1957 (N_1957,N_1323,N_1050);
and U1958 (N_1958,N_1015,N_1035);
or U1959 (N_1959,N_1442,N_1484);
nor U1960 (N_1960,N_1198,N_1420);
xor U1961 (N_1961,N_1186,N_1237);
or U1962 (N_1962,N_1142,N_1097);
and U1963 (N_1963,N_1156,N_1408);
and U1964 (N_1964,N_1023,N_1313);
or U1965 (N_1965,N_1111,N_1045);
nand U1966 (N_1966,N_1062,N_1303);
nand U1967 (N_1967,N_1107,N_1171);
or U1968 (N_1968,N_1001,N_1486);
or U1969 (N_1969,N_1281,N_1239);
or U1970 (N_1970,N_1049,N_1137);
nand U1971 (N_1971,N_1206,N_1372);
nand U1972 (N_1972,N_1368,N_1008);
and U1973 (N_1973,N_1232,N_1268);
and U1974 (N_1974,N_1011,N_1354);
nand U1975 (N_1975,N_1239,N_1012);
nor U1976 (N_1976,N_1019,N_1148);
and U1977 (N_1977,N_1167,N_1062);
nand U1978 (N_1978,N_1257,N_1173);
and U1979 (N_1979,N_1171,N_1292);
nor U1980 (N_1980,N_1488,N_1448);
nor U1981 (N_1981,N_1042,N_1069);
and U1982 (N_1982,N_1118,N_1083);
and U1983 (N_1983,N_1265,N_1063);
or U1984 (N_1984,N_1079,N_1149);
or U1985 (N_1985,N_1378,N_1190);
nand U1986 (N_1986,N_1399,N_1158);
nor U1987 (N_1987,N_1155,N_1228);
nand U1988 (N_1988,N_1001,N_1436);
and U1989 (N_1989,N_1451,N_1349);
nor U1990 (N_1990,N_1498,N_1159);
nand U1991 (N_1991,N_1272,N_1234);
nor U1992 (N_1992,N_1236,N_1020);
xnor U1993 (N_1993,N_1064,N_1330);
nand U1994 (N_1994,N_1268,N_1056);
nor U1995 (N_1995,N_1278,N_1302);
or U1996 (N_1996,N_1238,N_1326);
or U1997 (N_1997,N_1032,N_1370);
and U1998 (N_1998,N_1031,N_1242);
xnor U1999 (N_1999,N_1022,N_1157);
nand U2000 (N_2000,N_1588,N_1644);
and U2001 (N_2001,N_1628,N_1734);
or U2002 (N_2002,N_1694,N_1864);
or U2003 (N_2003,N_1551,N_1893);
or U2004 (N_2004,N_1652,N_1677);
or U2005 (N_2005,N_1689,N_1754);
nand U2006 (N_2006,N_1880,N_1662);
nor U2007 (N_2007,N_1927,N_1611);
or U2008 (N_2008,N_1943,N_1769);
xor U2009 (N_2009,N_1954,N_1862);
nor U2010 (N_2010,N_1825,N_1740);
nor U2011 (N_2011,N_1994,N_1956);
nor U2012 (N_2012,N_1868,N_1846);
or U2013 (N_2013,N_1783,N_1630);
xor U2014 (N_2014,N_1668,N_1741);
nand U2015 (N_2015,N_1791,N_1571);
or U2016 (N_2016,N_1724,N_1803);
or U2017 (N_2017,N_1530,N_1801);
nand U2018 (N_2018,N_1703,N_1505);
or U2019 (N_2019,N_1633,N_1568);
nand U2020 (N_2020,N_1701,N_1805);
or U2021 (N_2021,N_1558,N_1720);
nor U2022 (N_2022,N_1583,N_1676);
and U2023 (N_2023,N_1596,N_1716);
nand U2024 (N_2024,N_1828,N_1804);
xor U2025 (N_2025,N_1768,N_1678);
xnor U2026 (N_2026,N_1971,N_1570);
xnor U2027 (N_2027,N_1522,N_1934);
nand U2028 (N_2028,N_1939,N_1706);
nand U2029 (N_2029,N_1634,N_1746);
and U2030 (N_2030,N_1753,N_1503);
and U2031 (N_2031,N_1721,N_1714);
and U2032 (N_2032,N_1873,N_1591);
and U2033 (N_2033,N_1578,N_1580);
nor U2034 (N_2034,N_1871,N_1926);
nand U2035 (N_2035,N_1737,N_1619);
and U2036 (N_2036,N_1654,N_1625);
nor U2037 (N_2037,N_1765,N_1723);
nand U2038 (N_2038,N_1524,N_1750);
and U2039 (N_2039,N_1692,N_1974);
and U2040 (N_2040,N_1916,N_1879);
or U2041 (N_2041,N_1743,N_1539);
nand U2042 (N_2042,N_1976,N_1772);
and U2043 (N_2043,N_1798,N_1606);
nand U2044 (N_2044,N_1840,N_1730);
or U2045 (N_2045,N_1914,N_1671);
nor U2046 (N_2046,N_1639,N_1739);
nand U2047 (N_2047,N_1712,N_1529);
nor U2048 (N_2048,N_1523,N_1755);
or U2049 (N_2049,N_1520,N_1673);
nor U2050 (N_2050,N_1695,N_1502);
and U2051 (N_2051,N_1747,N_1988);
nand U2052 (N_2052,N_1777,N_1567);
or U2053 (N_2053,N_1744,N_1627);
nor U2054 (N_2054,N_1637,N_1506);
nor U2055 (N_2055,N_1655,N_1843);
nand U2056 (N_2056,N_1961,N_1715);
nor U2057 (N_2057,N_1788,N_1680);
nor U2058 (N_2058,N_1796,N_1776);
or U2059 (N_2059,N_1728,N_1733);
or U2060 (N_2060,N_1615,N_1736);
and U2061 (N_2061,N_1887,N_1582);
xnor U2062 (N_2062,N_1781,N_1667);
nor U2063 (N_2063,N_1857,N_1647);
nand U2064 (N_2064,N_1709,N_1635);
nand U2065 (N_2065,N_1561,N_1649);
xnor U2066 (N_2066,N_1885,N_1910);
or U2067 (N_2067,N_1665,N_1574);
and U2068 (N_2068,N_1812,N_1780);
nand U2069 (N_2069,N_1593,N_1684);
nor U2070 (N_2070,N_1980,N_1917);
or U2071 (N_2071,N_1653,N_1786);
nand U2072 (N_2072,N_1918,N_1831);
and U2073 (N_2073,N_1936,N_1758);
nor U2074 (N_2074,N_1845,N_1546);
nor U2075 (N_2075,N_1911,N_1981);
and U2076 (N_2076,N_1824,N_1953);
or U2077 (N_2077,N_1519,N_1802);
nand U2078 (N_2078,N_1566,N_1516);
nand U2079 (N_2079,N_1563,N_1512);
nor U2080 (N_2080,N_1973,N_1919);
nand U2081 (N_2081,N_1713,N_1995);
or U2082 (N_2082,N_1621,N_1731);
nand U2083 (N_2083,N_1617,N_1760);
and U2084 (N_2084,N_1535,N_1534);
or U2085 (N_2085,N_1807,N_1682);
or U2086 (N_2086,N_1930,N_1726);
or U2087 (N_2087,N_1874,N_1609);
or U2088 (N_2088,N_1823,N_1544);
nor U2089 (N_2089,N_1860,N_1763);
and U2090 (N_2090,N_1979,N_1827);
and U2091 (N_2091,N_1854,N_1509);
nand U2092 (N_2092,N_1842,N_1688);
nor U2093 (N_2093,N_1891,N_1945);
nor U2094 (N_2094,N_1993,N_1895);
nor U2095 (N_2095,N_1921,N_1821);
and U2096 (N_2096,N_1792,N_1810);
or U2097 (N_2097,N_1577,N_1901);
or U2098 (N_2098,N_1983,N_1996);
and U2099 (N_2099,N_1527,N_1764);
and U2100 (N_2100,N_1866,N_1686);
or U2101 (N_2101,N_1526,N_1500);
nand U2102 (N_2102,N_1614,N_1656);
or U2103 (N_2103,N_1541,N_1612);
and U2104 (N_2104,N_1896,N_1844);
nor U2105 (N_2105,N_1906,N_1705);
or U2106 (N_2106,N_1900,N_1648);
nand U2107 (N_2107,N_1597,N_1779);
nand U2108 (N_2108,N_1929,N_1587);
nor U2109 (N_2109,N_1538,N_1959);
or U2110 (N_2110,N_1757,N_1951);
and U2111 (N_2111,N_1833,N_1933);
xor U2112 (N_2112,N_1847,N_1550);
nand U2113 (N_2113,N_1972,N_1555);
nor U2114 (N_2114,N_1790,N_1602);
nor U2115 (N_2115,N_1560,N_1931);
or U2116 (N_2116,N_1987,N_1819);
nand U2117 (N_2117,N_1977,N_1870);
nor U2118 (N_2118,N_1839,N_1970);
nor U2119 (N_2119,N_1809,N_1732);
or U2120 (N_2120,N_1685,N_1638);
and U2121 (N_2121,N_1661,N_1968);
and U2122 (N_2122,N_1664,N_1909);
and U2123 (N_2123,N_1964,N_1669);
and U2124 (N_2124,N_1872,N_1863);
nor U2125 (N_2125,N_1585,N_1888);
nor U2126 (N_2126,N_1774,N_1882);
and U2127 (N_2127,N_1745,N_1898);
nand U2128 (N_2128,N_1965,N_1690);
xnor U2129 (N_2129,N_1575,N_1679);
nor U2130 (N_2130,N_1818,N_1889);
xnor U2131 (N_2131,N_1899,N_1794);
and U2132 (N_2132,N_1725,N_1511);
and U2133 (N_2133,N_1814,N_1675);
xnor U2134 (N_2134,N_1850,N_1579);
or U2135 (N_2135,N_1651,N_1576);
nand U2136 (N_2136,N_1643,N_1504);
nand U2137 (N_2137,N_1629,N_1600);
and U2138 (N_2138,N_1928,N_1806);
nand U2139 (N_2139,N_1982,N_1528);
xnor U2140 (N_2140,N_1967,N_1749);
and U2141 (N_2141,N_1663,N_1631);
and U2142 (N_2142,N_1830,N_1960);
and U2143 (N_2143,N_1607,N_1515);
nand U2144 (N_2144,N_1697,N_1729);
and U2145 (N_2145,N_1822,N_1962);
nand U2146 (N_2146,N_1955,N_1997);
and U2147 (N_2147,N_1573,N_1562);
and U2148 (N_2148,N_1838,N_1565);
or U2149 (N_2149,N_1944,N_1815);
nand U2150 (N_2150,N_1553,N_1952);
and U2151 (N_2151,N_1829,N_1589);
and U2152 (N_2152,N_1853,N_1817);
and U2153 (N_2153,N_1532,N_1811);
nor U2154 (N_2154,N_1517,N_1691);
or U2155 (N_2155,N_1892,N_1610);
and U2156 (N_2156,N_1975,N_1543);
and U2157 (N_2157,N_1640,N_1548);
xnor U2158 (N_2158,N_1702,N_1800);
nand U2159 (N_2159,N_1894,N_1700);
nor U2160 (N_2160,N_1905,N_1518);
or U2161 (N_2161,N_1549,N_1525);
or U2162 (N_2162,N_1545,N_1711);
xor U2163 (N_2163,N_1787,N_1658);
nor U2164 (N_2164,N_1698,N_1937);
nand U2165 (N_2165,N_1799,N_1957);
xor U2166 (N_2166,N_1849,N_1547);
and U2167 (N_2167,N_1837,N_1922);
and U2168 (N_2168,N_1969,N_1510);
nand U2169 (N_2169,N_1966,N_1590);
nor U2170 (N_2170,N_1521,N_1938);
or U2171 (N_2171,N_1820,N_1935);
or U2172 (N_2172,N_1657,N_1594);
nor U2173 (N_2173,N_1708,N_1950);
and U2174 (N_2174,N_1795,N_1537);
or U2175 (N_2175,N_1797,N_1855);
xor U2176 (N_2176,N_1650,N_1572);
and U2177 (N_2177,N_1598,N_1998);
or U2178 (N_2178,N_1907,N_1727);
and U2179 (N_2179,N_1766,N_1858);
nor U2180 (N_2180,N_1687,N_1989);
nor U2181 (N_2181,N_1599,N_1645);
or U2182 (N_2182,N_1681,N_1861);
and U2183 (N_2183,N_1865,N_1875);
and U2184 (N_2184,N_1641,N_1856);
and U2185 (N_2185,N_1592,N_1770);
nand U2186 (N_2186,N_1834,N_1704);
or U2187 (N_2187,N_1642,N_1913);
nor U2188 (N_2188,N_1782,N_1569);
or U2189 (N_2189,N_1948,N_1912);
nor U2190 (N_2190,N_1767,N_1603);
xnor U2191 (N_2191,N_1742,N_1696);
and U2192 (N_2192,N_1683,N_1886);
and U2193 (N_2193,N_1738,N_1883);
or U2194 (N_2194,N_1848,N_1622);
or U2195 (N_2195,N_1990,N_1958);
or U2196 (N_2196,N_1670,N_1632);
nor U2197 (N_2197,N_1775,N_1841);
and U2198 (N_2198,N_1748,N_1785);
nand U2199 (N_2199,N_1514,N_1908);
or U2200 (N_2200,N_1717,N_1897);
or U2201 (N_2201,N_1789,N_1604);
or U2202 (N_2202,N_1808,N_1608);
nor U2203 (N_2203,N_1623,N_1719);
or U2204 (N_2204,N_1867,N_1508);
nor U2205 (N_2205,N_1876,N_1626);
and U2206 (N_2206,N_1942,N_1531);
nor U2207 (N_2207,N_1816,N_1773);
nand U2208 (N_2208,N_1540,N_1923);
nand U2209 (N_2209,N_1978,N_1659);
nor U2210 (N_2210,N_1784,N_1536);
nand U2211 (N_2211,N_1693,N_1557);
nand U2212 (N_2212,N_1752,N_1559);
and U2213 (N_2213,N_1832,N_1771);
or U2214 (N_2214,N_1710,N_1722);
nor U2215 (N_2215,N_1616,N_1920);
nor U2216 (N_2216,N_1507,N_1826);
nor U2217 (N_2217,N_1904,N_1707);
nand U2218 (N_2218,N_1778,N_1533);
or U2219 (N_2219,N_1963,N_1991);
xor U2220 (N_2220,N_1984,N_1718);
nor U2221 (N_2221,N_1660,N_1890);
and U2222 (N_2222,N_1946,N_1618);
or U2223 (N_2223,N_1947,N_1554);
and U2224 (N_2224,N_1999,N_1513);
nand U2225 (N_2225,N_1556,N_1552);
nor U2226 (N_2226,N_1564,N_1601);
xor U2227 (N_2227,N_1859,N_1877);
xnor U2228 (N_2228,N_1986,N_1735);
and U2229 (N_2229,N_1620,N_1699);
nand U2230 (N_2230,N_1836,N_1636);
xnor U2231 (N_2231,N_1932,N_1613);
xor U2232 (N_2232,N_1925,N_1878);
nor U2233 (N_2233,N_1756,N_1924);
nor U2234 (N_2234,N_1852,N_1869);
nor U2235 (N_2235,N_1884,N_1605);
and U2236 (N_2236,N_1949,N_1761);
nor U2237 (N_2237,N_1666,N_1595);
nand U2238 (N_2238,N_1881,N_1586);
or U2239 (N_2239,N_1902,N_1674);
nor U2240 (N_2240,N_1646,N_1584);
xnor U2241 (N_2241,N_1851,N_1501);
and U2242 (N_2242,N_1759,N_1793);
nor U2243 (N_2243,N_1542,N_1940);
and U2244 (N_2244,N_1581,N_1915);
nand U2245 (N_2245,N_1835,N_1992);
nand U2246 (N_2246,N_1813,N_1751);
xor U2247 (N_2247,N_1941,N_1762);
nor U2248 (N_2248,N_1672,N_1985);
nand U2249 (N_2249,N_1624,N_1903);
nand U2250 (N_2250,N_1613,N_1914);
or U2251 (N_2251,N_1780,N_1916);
and U2252 (N_2252,N_1853,N_1567);
nor U2253 (N_2253,N_1628,N_1538);
nor U2254 (N_2254,N_1566,N_1563);
or U2255 (N_2255,N_1903,N_1765);
nand U2256 (N_2256,N_1578,N_1523);
and U2257 (N_2257,N_1504,N_1812);
and U2258 (N_2258,N_1590,N_1713);
nor U2259 (N_2259,N_1506,N_1814);
and U2260 (N_2260,N_1883,N_1679);
nand U2261 (N_2261,N_1834,N_1988);
nand U2262 (N_2262,N_1870,N_1678);
or U2263 (N_2263,N_1586,N_1713);
xnor U2264 (N_2264,N_1601,N_1835);
nor U2265 (N_2265,N_1685,N_1731);
and U2266 (N_2266,N_1557,N_1928);
and U2267 (N_2267,N_1574,N_1707);
xor U2268 (N_2268,N_1515,N_1981);
or U2269 (N_2269,N_1892,N_1559);
nand U2270 (N_2270,N_1621,N_1892);
and U2271 (N_2271,N_1656,N_1632);
or U2272 (N_2272,N_1902,N_1739);
nor U2273 (N_2273,N_1955,N_1986);
nand U2274 (N_2274,N_1727,N_1541);
nor U2275 (N_2275,N_1607,N_1699);
nor U2276 (N_2276,N_1832,N_1782);
or U2277 (N_2277,N_1642,N_1819);
or U2278 (N_2278,N_1714,N_1937);
and U2279 (N_2279,N_1734,N_1526);
nor U2280 (N_2280,N_1515,N_1585);
or U2281 (N_2281,N_1592,N_1522);
and U2282 (N_2282,N_1906,N_1992);
and U2283 (N_2283,N_1858,N_1853);
nand U2284 (N_2284,N_1621,N_1938);
nor U2285 (N_2285,N_1793,N_1935);
nor U2286 (N_2286,N_1868,N_1860);
nor U2287 (N_2287,N_1693,N_1622);
or U2288 (N_2288,N_1705,N_1900);
nand U2289 (N_2289,N_1684,N_1827);
or U2290 (N_2290,N_1705,N_1775);
nor U2291 (N_2291,N_1829,N_1644);
or U2292 (N_2292,N_1524,N_1755);
and U2293 (N_2293,N_1894,N_1810);
and U2294 (N_2294,N_1990,N_1987);
xor U2295 (N_2295,N_1975,N_1978);
and U2296 (N_2296,N_1797,N_1540);
nand U2297 (N_2297,N_1848,N_1738);
or U2298 (N_2298,N_1955,N_1573);
nand U2299 (N_2299,N_1937,N_1966);
or U2300 (N_2300,N_1554,N_1899);
or U2301 (N_2301,N_1990,N_1819);
or U2302 (N_2302,N_1835,N_1872);
nand U2303 (N_2303,N_1583,N_1974);
and U2304 (N_2304,N_1716,N_1675);
nand U2305 (N_2305,N_1982,N_1717);
and U2306 (N_2306,N_1537,N_1903);
xor U2307 (N_2307,N_1803,N_1507);
nand U2308 (N_2308,N_1636,N_1691);
or U2309 (N_2309,N_1873,N_1866);
or U2310 (N_2310,N_1659,N_1924);
and U2311 (N_2311,N_1608,N_1582);
and U2312 (N_2312,N_1864,N_1552);
or U2313 (N_2313,N_1560,N_1891);
nand U2314 (N_2314,N_1650,N_1622);
xor U2315 (N_2315,N_1963,N_1700);
nor U2316 (N_2316,N_1648,N_1608);
or U2317 (N_2317,N_1791,N_1614);
nor U2318 (N_2318,N_1546,N_1830);
xnor U2319 (N_2319,N_1887,N_1957);
or U2320 (N_2320,N_1637,N_1677);
and U2321 (N_2321,N_1882,N_1829);
nand U2322 (N_2322,N_1570,N_1863);
xnor U2323 (N_2323,N_1710,N_1625);
nand U2324 (N_2324,N_1811,N_1987);
or U2325 (N_2325,N_1581,N_1872);
and U2326 (N_2326,N_1908,N_1975);
nor U2327 (N_2327,N_1874,N_1580);
nor U2328 (N_2328,N_1604,N_1600);
nand U2329 (N_2329,N_1800,N_1749);
xnor U2330 (N_2330,N_1782,N_1680);
nand U2331 (N_2331,N_1917,N_1715);
xor U2332 (N_2332,N_1908,N_1703);
and U2333 (N_2333,N_1580,N_1598);
nor U2334 (N_2334,N_1794,N_1606);
or U2335 (N_2335,N_1638,N_1859);
and U2336 (N_2336,N_1823,N_1954);
and U2337 (N_2337,N_1599,N_1727);
xnor U2338 (N_2338,N_1804,N_1888);
nor U2339 (N_2339,N_1696,N_1655);
nand U2340 (N_2340,N_1935,N_1503);
nor U2341 (N_2341,N_1888,N_1799);
nor U2342 (N_2342,N_1739,N_1520);
or U2343 (N_2343,N_1986,N_1764);
nand U2344 (N_2344,N_1884,N_1549);
nand U2345 (N_2345,N_1935,N_1934);
and U2346 (N_2346,N_1562,N_1700);
or U2347 (N_2347,N_1707,N_1562);
nand U2348 (N_2348,N_1937,N_1744);
xor U2349 (N_2349,N_1783,N_1745);
and U2350 (N_2350,N_1592,N_1729);
nand U2351 (N_2351,N_1823,N_1834);
nand U2352 (N_2352,N_1698,N_1563);
nand U2353 (N_2353,N_1741,N_1765);
and U2354 (N_2354,N_1901,N_1853);
and U2355 (N_2355,N_1865,N_1910);
nand U2356 (N_2356,N_1832,N_1587);
and U2357 (N_2357,N_1676,N_1628);
and U2358 (N_2358,N_1804,N_1671);
or U2359 (N_2359,N_1828,N_1700);
and U2360 (N_2360,N_1719,N_1892);
and U2361 (N_2361,N_1942,N_1594);
nand U2362 (N_2362,N_1752,N_1994);
nor U2363 (N_2363,N_1799,N_1731);
or U2364 (N_2364,N_1987,N_1837);
and U2365 (N_2365,N_1639,N_1886);
and U2366 (N_2366,N_1850,N_1843);
nor U2367 (N_2367,N_1663,N_1940);
nor U2368 (N_2368,N_1784,N_1971);
and U2369 (N_2369,N_1628,N_1700);
nand U2370 (N_2370,N_1793,N_1916);
nor U2371 (N_2371,N_1586,N_1631);
and U2372 (N_2372,N_1768,N_1988);
xor U2373 (N_2373,N_1948,N_1985);
nor U2374 (N_2374,N_1588,N_1541);
or U2375 (N_2375,N_1646,N_1689);
and U2376 (N_2376,N_1764,N_1687);
nand U2377 (N_2377,N_1642,N_1888);
nor U2378 (N_2378,N_1699,N_1741);
nand U2379 (N_2379,N_1867,N_1852);
and U2380 (N_2380,N_1784,N_1515);
or U2381 (N_2381,N_1699,N_1772);
and U2382 (N_2382,N_1525,N_1700);
and U2383 (N_2383,N_1794,N_1932);
and U2384 (N_2384,N_1725,N_1666);
or U2385 (N_2385,N_1736,N_1707);
or U2386 (N_2386,N_1777,N_1811);
or U2387 (N_2387,N_1617,N_1766);
nand U2388 (N_2388,N_1979,N_1882);
and U2389 (N_2389,N_1943,N_1640);
nor U2390 (N_2390,N_1999,N_1595);
and U2391 (N_2391,N_1767,N_1860);
nor U2392 (N_2392,N_1852,N_1953);
nor U2393 (N_2393,N_1769,N_1633);
and U2394 (N_2394,N_1504,N_1843);
nand U2395 (N_2395,N_1917,N_1505);
nor U2396 (N_2396,N_1805,N_1668);
or U2397 (N_2397,N_1875,N_1656);
and U2398 (N_2398,N_1797,N_1760);
and U2399 (N_2399,N_1630,N_1997);
or U2400 (N_2400,N_1625,N_1634);
xor U2401 (N_2401,N_1886,N_1753);
and U2402 (N_2402,N_1864,N_1673);
nand U2403 (N_2403,N_1973,N_1528);
nand U2404 (N_2404,N_1520,N_1745);
xor U2405 (N_2405,N_1512,N_1886);
nor U2406 (N_2406,N_1958,N_1655);
nand U2407 (N_2407,N_1713,N_1598);
or U2408 (N_2408,N_1603,N_1597);
nor U2409 (N_2409,N_1885,N_1729);
nand U2410 (N_2410,N_1883,N_1529);
nand U2411 (N_2411,N_1975,N_1502);
xor U2412 (N_2412,N_1509,N_1560);
nand U2413 (N_2413,N_1597,N_1627);
or U2414 (N_2414,N_1501,N_1912);
nand U2415 (N_2415,N_1823,N_1675);
and U2416 (N_2416,N_1738,N_1922);
nor U2417 (N_2417,N_1772,N_1863);
or U2418 (N_2418,N_1789,N_1570);
nand U2419 (N_2419,N_1808,N_1806);
nor U2420 (N_2420,N_1872,N_1972);
and U2421 (N_2421,N_1684,N_1979);
xnor U2422 (N_2422,N_1913,N_1767);
and U2423 (N_2423,N_1865,N_1982);
xor U2424 (N_2424,N_1758,N_1931);
and U2425 (N_2425,N_1548,N_1930);
or U2426 (N_2426,N_1912,N_1775);
nand U2427 (N_2427,N_1867,N_1929);
or U2428 (N_2428,N_1544,N_1637);
nand U2429 (N_2429,N_1868,N_1908);
nand U2430 (N_2430,N_1915,N_1508);
or U2431 (N_2431,N_1800,N_1843);
nand U2432 (N_2432,N_1572,N_1881);
and U2433 (N_2433,N_1677,N_1859);
nand U2434 (N_2434,N_1546,N_1770);
nor U2435 (N_2435,N_1868,N_1524);
and U2436 (N_2436,N_1614,N_1521);
nor U2437 (N_2437,N_1861,N_1702);
and U2438 (N_2438,N_1955,N_1937);
nor U2439 (N_2439,N_1850,N_1518);
and U2440 (N_2440,N_1724,N_1877);
and U2441 (N_2441,N_1874,N_1925);
or U2442 (N_2442,N_1771,N_1515);
nand U2443 (N_2443,N_1866,N_1683);
nor U2444 (N_2444,N_1840,N_1876);
nor U2445 (N_2445,N_1907,N_1570);
or U2446 (N_2446,N_1534,N_1891);
and U2447 (N_2447,N_1741,N_1602);
or U2448 (N_2448,N_1896,N_1715);
xor U2449 (N_2449,N_1641,N_1973);
nand U2450 (N_2450,N_1762,N_1578);
xor U2451 (N_2451,N_1773,N_1899);
xor U2452 (N_2452,N_1706,N_1925);
or U2453 (N_2453,N_1537,N_1512);
and U2454 (N_2454,N_1685,N_1960);
and U2455 (N_2455,N_1810,N_1784);
nor U2456 (N_2456,N_1685,N_1815);
or U2457 (N_2457,N_1784,N_1808);
and U2458 (N_2458,N_1656,N_1951);
nand U2459 (N_2459,N_1994,N_1515);
xnor U2460 (N_2460,N_1717,N_1987);
and U2461 (N_2461,N_1903,N_1875);
nor U2462 (N_2462,N_1524,N_1757);
or U2463 (N_2463,N_1567,N_1997);
or U2464 (N_2464,N_1884,N_1979);
nand U2465 (N_2465,N_1924,N_1909);
or U2466 (N_2466,N_1646,N_1966);
and U2467 (N_2467,N_1574,N_1673);
nand U2468 (N_2468,N_1660,N_1520);
or U2469 (N_2469,N_1868,N_1681);
xor U2470 (N_2470,N_1560,N_1708);
nand U2471 (N_2471,N_1506,N_1685);
nand U2472 (N_2472,N_1945,N_1983);
or U2473 (N_2473,N_1948,N_1663);
nand U2474 (N_2474,N_1518,N_1595);
xor U2475 (N_2475,N_1795,N_1751);
nand U2476 (N_2476,N_1555,N_1997);
nand U2477 (N_2477,N_1760,N_1694);
nand U2478 (N_2478,N_1936,N_1547);
nand U2479 (N_2479,N_1759,N_1536);
or U2480 (N_2480,N_1783,N_1887);
nand U2481 (N_2481,N_1844,N_1996);
nand U2482 (N_2482,N_1508,N_1926);
or U2483 (N_2483,N_1975,N_1549);
nand U2484 (N_2484,N_1992,N_1859);
and U2485 (N_2485,N_1552,N_1592);
and U2486 (N_2486,N_1613,N_1706);
nand U2487 (N_2487,N_1849,N_1635);
or U2488 (N_2488,N_1834,N_1799);
and U2489 (N_2489,N_1943,N_1780);
or U2490 (N_2490,N_1718,N_1596);
nand U2491 (N_2491,N_1581,N_1628);
nand U2492 (N_2492,N_1666,N_1611);
nand U2493 (N_2493,N_1719,N_1994);
nor U2494 (N_2494,N_1964,N_1748);
or U2495 (N_2495,N_1695,N_1786);
nor U2496 (N_2496,N_1716,N_1893);
nor U2497 (N_2497,N_1919,N_1514);
nor U2498 (N_2498,N_1589,N_1552);
nor U2499 (N_2499,N_1934,N_1961);
nand U2500 (N_2500,N_2309,N_2271);
or U2501 (N_2501,N_2369,N_2331);
or U2502 (N_2502,N_2325,N_2244);
nor U2503 (N_2503,N_2249,N_2378);
xor U2504 (N_2504,N_2477,N_2110);
and U2505 (N_2505,N_2456,N_2209);
xnor U2506 (N_2506,N_2113,N_2047);
or U2507 (N_2507,N_2138,N_2350);
nand U2508 (N_2508,N_2391,N_2037);
nand U2509 (N_2509,N_2355,N_2485);
nand U2510 (N_2510,N_2275,N_2360);
and U2511 (N_2511,N_2186,N_2264);
xor U2512 (N_2512,N_2351,N_2393);
or U2513 (N_2513,N_2039,N_2321);
xor U2514 (N_2514,N_2376,N_2070);
nor U2515 (N_2515,N_2294,N_2297);
nand U2516 (N_2516,N_2493,N_2109);
and U2517 (N_2517,N_2478,N_2265);
nand U2518 (N_2518,N_2229,N_2289);
nor U2519 (N_2519,N_2329,N_2248);
xor U2520 (N_2520,N_2434,N_2164);
or U2521 (N_2521,N_2496,N_2084);
nor U2522 (N_2522,N_2214,N_2380);
and U2523 (N_2523,N_2292,N_2274);
xnor U2524 (N_2524,N_2111,N_2449);
xnor U2525 (N_2525,N_2421,N_2095);
and U2526 (N_2526,N_2147,N_2238);
xnor U2527 (N_2527,N_2291,N_2306);
and U2528 (N_2528,N_2464,N_2128);
or U2529 (N_2529,N_2323,N_2069);
xnor U2530 (N_2530,N_2447,N_2403);
and U2531 (N_2531,N_2259,N_2319);
nor U2532 (N_2532,N_2405,N_2361);
nor U2533 (N_2533,N_2232,N_2141);
and U2534 (N_2534,N_2282,N_2389);
and U2535 (N_2535,N_2311,N_2367);
nand U2536 (N_2536,N_2190,N_2416);
and U2537 (N_2537,N_2102,N_2395);
or U2538 (N_2538,N_2176,N_2153);
nor U2539 (N_2539,N_2210,N_2430);
or U2540 (N_2540,N_2051,N_2221);
or U2541 (N_2541,N_2452,N_2031);
nand U2542 (N_2542,N_2359,N_2060);
nor U2543 (N_2543,N_2363,N_2061);
nand U2544 (N_2544,N_2009,N_2412);
nor U2545 (N_2545,N_2087,N_2358);
nand U2546 (N_2546,N_2152,N_2489);
nand U2547 (N_2547,N_2383,N_2114);
nand U2548 (N_2548,N_2154,N_2415);
nor U2549 (N_2549,N_2440,N_2370);
nor U2550 (N_2550,N_2173,N_2174);
nand U2551 (N_2551,N_2242,N_2427);
and U2552 (N_2552,N_2287,N_2071);
and U2553 (N_2553,N_2143,N_2123);
nand U2554 (N_2554,N_2025,N_2027);
or U2555 (N_2555,N_2055,N_2046);
nor U2556 (N_2556,N_2068,N_2347);
nor U2557 (N_2557,N_2165,N_2345);
nor U2558 (N_2558,N_2388,N_2101);
and U2559 (N_2559,N_2012,N_2273);
nand U2560 (N_2560,N_2450,N_2014);
nand U2561 (N_2561,N_2056,N_2356);
nor U2562 (N_2562,N_2285,N_2301);
or U2563 (N_2563,N_2300,N_2092);
or U2564 (N_2564,N_2234,N_2466);
nor U2565 (N_2565,N_2467,N_2136);
nand U2566 (N_2566,N_2052,N_2451);
and U2567 (N_2567,N_2220,N_2097);
and U2568 (N_2568,N_2317,N_2327);
nor U2569 (N_2569,N_2365,N_2333);
nand U2570 (N_2570,N_2015,N_2318);
nor U2571 (N_2571,N_2353,N_2048);
and U2572 (N_2572,N_2105,N_2179);
and U2573 (N_2573,N_2150,N_2194);
or U2574 (N_2574,N_2100,N_2066);
or U2575 (N_2575,N_2419,N_2126);
and U2576 (N_2576,N_2324,N_2151);
and U2577 (N_2577,N_2235,N_2156);
and U2578 (N_2578,N_2334,N_2437);
and U2579 (N_2579,N_2423,N_2483);
or U2580 (N_2580,N_2366,N_2339);
or U2581 (N_2581,N_2187,N_2083);
nor U2582 (N_2582,N_2255,N_2304);
nor U2583 (N_2583,N_2195,N_2175);
or U2584 (N_2584,N_2094,N_2316);
nand U2585 (N_2585,N_2418,N_2044);
nor U2586 (N_2586,N_2207,N_2473);
or U2587 (N_2587,N_2426,N_2211);
nand U2588 (N_2588,N_2007,N_2305);
or U2589 (N_2589,N_2375,N_2033);
and U2590 (N_2590,N_2379,N_2402);
and U2591 (N_2591,N_2161,N_2253);
or U2592 (N_2592,N_2247,N_2251);
or U2593 (N_2593,N_2073,N_2178);
xnor U2594 (N_2594,N_2453,N_2326);
nand U2595 (N_2595,N_2429,N_2017);
and U2596 (N_2596,N_2462,N_2081);
nand U2597 (N_2597,N_2104,N_2299);
and U2598 (N_2598,N_2280,N_2112);
xnor U2599 (N_2599,N_2086,N_2307);
nand U2600 (N_2600,N_2283,N_2371);
nor U2601 (N_2601,N_2159,N_2279);
nand U2602 (N_2602,N_2240,N_2492);
nor U2603 (N_2603,N_2058,N_2257);
or U2604 (N_2604,N_2335,N_2461);
nand U2605 (N_2605,N_2116,N_2239);
xor U2606 (N_2606,N_2142,N_2144);
nand U2607 (N_2607,N_2448,N_2343);
xnor U2608 (N_2608,N_2054,N_2458);
nand U2609 (N_2609,N_2352,N_2053);
nand U2610 (N_2610,N_2133,N_2085);
nand U2611 (N_2611,N_2029,N_2124);
or U2612 (N_2612,N_2200,N_2362);
nand U2613 (N_2613,N_2459,N_2454);
nand U2614 (N_2614,N_2278,N_2432);
and U2615 (N_2615,N_2422,N_2020);
and U2616 (N_2616,N_2204,N_2106);
nand U2617 (N_2617,N_2243,N_2442);
nand U2618 (N_2618,N_2043,N_2225);
xnor U2619 (N_2619,N_2457,N_2443);
nand U2620 (N_2620,N_2246,N_2197);
nand U2621 (N_2621,N_2107,N_2099);
xnor U2622 (N_2622,N_2487,N_2199);
and U2623 (N_2623,N_2076,N_2198);
xnor U2624 (N_2624,N_2139,N_2494);
and U2625 (N_2625,N_2062,N_2320);
nor U2626 (N_2626,N_2192,N_2268);
nand U2627 (N_2627,N_2080,N_2149);
and U2628 (N_2628,N_2258,N_2172);
nor U2629 (N_2629,N_2293,N_2019);
or U2630 (N_2630,N_2188,N_2476);
nand U2631 (N_2631,N_2074,N_2120);
nor U2632 (N_2632,N_2148,N_2010);
or U2633 (N_2633,N_2469,N_2050);
and U2634 (N_2634,N_2460,N_2032);
nand U2635 (N_2635,N_2267,N_2011);
and U2636 (N_2636,N_2428,N_2330);
nor U2637 (N_2637,N_2277,N_2261);
nor U2638 (N_2638,N_2166,N_2286);
or U2639 (N_2639,N_2158,N_2129);
nor U2640 (N_2640,N_2308,N_2414);
nand U2641 (N_2641,N_2254,N_2222);
or U2642 (N_2642,N_2433,N_2404);
or U2643 (N_2643,N_2344,N_2013);
and U2644 (N_2644,N_2381,N_2018);
nand U2645 (N_2645,N_2337,N_2205);
or U2646 (N_2646,N_2130,N_2411);
or U2647 (N_2647,N_2262,N_2065);
nand U2648 (N_2648,N_2063,N_2470);
nor U2649 (N_2649,N_2218,N_2270);
nor U2650 (N_2650,N_2132,N_2193);
or U2651 (N_2651,N_2424,N_2227);
xnor U2652 (N_2652,N_2256,N_2290);
xnor U2653 (N_2653,N_2417,N_2398);
or U2654 (N_2654,N_2022,N_2226);
and U2655 (N_2655,N_2021,N_2281);
or U2656 (N_2656,N_2230,N_2185);
nor U2657 (N_2657,N_2410,N_2040);
xor U2658 (N_2658,N_2005,N_2059);
or U2659 (N_2659,N_2364,N_2328);
nand U2660 (N_2660,N_2206,N_2382);
and U2661 (N_2661,N_2446,N_2490);
or U2662 (N_2662,N_2284,N_2023);
and U2663 (N_2663,N_2409,N_2115);
xor U2664 (N_2664,N_2303,N_2224);
nor U2665 (N_2665,N_2008,N_2322);
xor U2666 (N_2666,N_2203,N_2397);
or U2667 (N_2667,N_2348,N_2310);
and U2668 (N_2668,N_2480,N_2387);
or U2669 (N_2669,N_2146,N_2042);
xor U2670 (N_2670,N_2215,N_2241);
nor U2671 (N_2671,N_2103,N_2171);
nor U2672 (N_2672,N_2245,N_2006);
xor U2673 (N_2673,N_2078,N_2368);
nor U2674 (N_2674,N_2216,N_2145);
and U2675 (N_2675,N_2400,N_2035);
nand U2676 (N_2676,N_2028,N_2436);
and U2677 (N_2677,N_2168,N_2341);
or U2678 (N_2678,N_2122,N_2385);
nor U2679 (N_2679,N_2024,N_2276);
nand U2680 (N_2680,N_2425,N_2336);
nand U2681 (N_2681,N_2497,N_2036);
or U2682 (N_2682,N_2406,N_2444);
nand U2683 (N_2683,N_2463,N_2096);
xor U2684 (N_2684,N_2498,N_2233);
nor U2685 (N_2685,N_2445,N_2413);
nand U2686 (N_2686,N_2137,N_2155);
nand U2687 (N_2687,N_2163,N_2135);
or U2688 (N_2688,N_2034,N_2202);
nand U2689 (N_2689,N_2119,N_2088);
nand U2690 (N_2690,N_2016,N_2077);
nand U2691 (N_2691,N_2495,N_2167);
xnor U2692 (N_2692,N_2396,N_2072);
and U2693 (N_2693,N_2407,N_2219);
nand U2694 (N_2694,N_2392,N_2089);
or U2695 (N_2695,N_2169,N_2184);
or U2696 (N_2696,N_2196,N_2313);
nand U2697 (N_2697,N_2468,N_2213);
or U2698 (N_2698,N_2302,N_2160);
or U2699 (N_2699,N_2482,N_2390);
nor U2700 (N_2700,N_2170,N_2486);
nor U2701 (N_2701,N_2475,N_2002);
nor U2702 (N_2702,N_2189,N_2180);
or U2703 (N_2703,N_2372,N_2228);
nor U2704 (N_2704,N_2401,N_2191);
nand U2705 (N_2705,N_2474,N_2314);
or U2706 (N_2706,N_2041,N_2374);
nand U2707 (N_2707,N_2064,N_2266);
nor U2708 (N_2708,N_2340,N_2030);
and U2709 (N_2709,N_2484,N_2026);
nand U2710 (N_2710,N_2098,N_2298);
nor U2711 (N_2711,N_2431,N_2217);
or U2712 (N_2712,N_2250,N_2231);
nand U2713 (N_2713,N_2472,N_2394);
nand U2714 (N_2714,N_2408,N_2332);
or U2715 (N_2715,N_2420,N_2399);
or U2716 (N_2716,N_2315,N_2471);
nand U2717 (N_2717,N_2288,N_2177);
nor U2718 (N_2718,N_2134,N_2342);
nand U2719 (N_2719,N_2441,N_2295);
or U2720 (N_2720,N_2237,N_2455);
nor U2721 (N_2721,N_2346,N_2201);
xnor U2722 (N_2722,N_2338,N_2272);
and U2723 (N_2723,N_2481,N_2140);
and U2724 (N_2724,N_2373,N_2349);
nand U2725 (N_2725,N_2079,N_2004);
nand U2726 (N_2726,N_2162,N_2001);
nor U2727 (N_2727,N_2183,N_2057);
nand U2728 (N_2728,N_2075,N_2263);
xor U2729 (N_2729,N_2067,N_2127);
or U2730 (N_2730,N_2049,N_2121);
or U2731 (N_2731,N_2479,N_2093);
and U2732 (N_2732,N_2045,N_2384);
xor U2733 (N_2733,N_2491,N_2090);
or U2734 (N_2734,N_2386,N_2465);
nand U2735 (N_2735,N_2223,N_2181);
nor U2736 (N_2736,N_2236,N_2312);
xor U2737 (N_2737,N_2435,N_2118);
nor U2738 (N_2738,N_2125,N_2091);
and U2739 (N_2739,N_2357,N_2000);
or U2740 (N_2740,N_2296,N_2354);
and U2741 (N_2741,N_2260,N_2182);
or U2742 (N_2742,N_2131,N_2082);
and U2743 (N_2743,N_2252,N_2269);
xor U2744 (N_2744,N_2038,N_2117);
and U2745 (N_2745,N_2003,N_2488);
or U2746 (N_2746,N_2108,N_2377);
xor U2747 (N_2747,N_2499,N_2212);
nand U2748 (N_2748,N_2439,N_2438);
nand U2749 (N_2749,N_2157,N_2208);
nand U2750 (N_2750,N_2165,N_2303);
nand U2751 (N_2751,N_2182,N_2001);
and U2752 (N_2752,N_2231,N_2385);
and U2753 (N_2753,N_2018,N_2260);
nand U2754 (N_2754,N_2438,N_2472);
nand U2755 (N_2755,N_2281,N_2232);
nand U2756 (N_2756,N_2027,N_2195);
nand U2757 (N_2757,N_2078,N_2319);
or U2758 (N_2758,N_2164,N_2430);
or U2759 (N_2759,N_2468,N_2472);
xnor U2760 (N_2760,N_2072,N_2205);
and U2761 (N_2761,N_2486,N_2151);
xor U2762 (N_2762,N_2039,N_2088);
or U2763 (N_2763,N_2096,N_2162);
nor U2764 (N_2764,N_2141,N_2112);
nor U2765 (N_2765,N_2144,N_2444);
nor U2766 (N_2766,N_2018,N_2487);
nor U2767 (N_2767,N_2434,N_2393);
and U2768 (N_2768,N_2389,N_2319);
nand U2769 (N_2769,N_2296,N_2015);
nand U2770 (N_2770,N_2258,N_2016);
and U2771 (N_2771,N_2426,N_2323);
nand U2772 (N_2772,N_2389,N_2100);
nor U2773 (N_2773,N_2173,N_2145);
xor U2774 (N_2774,N_2401,N_2358);
or U2775 (N_2775,N_2162,N_2429);
and U2776 (N_2776,N_2089,N_2214);
and U2777 (N_2777,N_2269,N_2024);
or U2778 (N_2778,N_2486,N_2439);
or U2779 (N_2779,N_2049,N_2267);
nand U2780 (N_2780,N_2399,N_2351);
or U2781 (N_2781,N_2146,N_2303);
nor U2782 (N_2782,N_2159,N_2260);
xor U2783 (N_2783,N_2283,N_2377);
and U2784 (N_2784,N_2400,N_2160);
nor U2785 (N_2785,N_2319,N_2085);
nand U2786 (N_2786,N_2065,N_2202);
xnor U2787 (N_2787,N_2359,N_2482);
and U2788 (N_2788,N_2443,N_2316);
or U2789 (N_2789,N_2453,N_2193);
nand U2790 (N_2790,N_2138,N_2447);
nor U2791 (N_2791,N_2330,N_2467);
nand U2792 (N_2792,N_2105,N_2468);
or U2793 (N_2793,N_2454,N_2298);
xnor U2794 (N_2794,N_2265,N_2243);
or U2795 (N_2795,N_2442,N_2367);
nand U2796 (N_2796,N_2114,N_2122);
xnor U2797 (N_2797,N_2284,N_2085);
nand U2798 (N_2798,N_2353,N_2294);
nor U2799 (N_2799,N_2363,N_2246);
nor U2800 (N_2800,N_2347,N_2357);
nand U2801 (N_2801,N_2495,N_2186);
and U2802 (N_2802,N_2398,N_2070);
nand U2803 (N_2803,N_2031,N_2117);
nor U2804 (N_2804,N_2205,N_2448);
xor U2805 (N_2805,N_2075,N_2375);
or U2806 (N_2806,N_2015,N_2087);
or U2807 (N_2807,N_2275,N_2180);
nand U2808 (N_2808,N_2436,N_2262);
nor U2809 (N_2809,N_2464,N_2461);
xnor U2810 (N_2810,N_2083,N_2270);
nor U2811 (N_2811,N_2308,N_2353);
or U2812 (N_2812,N_2200,N_2281);
nand U2813 (N_2813,N_2039,N_2366);
nand U2814 (N_2814,N_2286,N_2083);
or U2815 (N_2815,N_2430,N_2275);
nor U2816 (N_2816,N_2118,N_2292);
and U2817 (N_2817,N_2430,N_2241);
nor U2818 (N_2818,N_2327,N_2160);
or U2819 (N_2819,N_2443,N_2175);
or U2820 (N_2820,N_2166,N_2321);
nor U2821 (N_2821,N_2166,N_2082);
and U2822 (N_2822,N_2414,N_2415);
nor U2823 (N_2823,N_2221,N_2248);
nor U2824 (N_2824,N_2319,N_2401);
xnor U2825 (N_2825,N_2499,N_2114);
and U2826 (N_2826,N_2026,N_2311);
nor U2827 (N_2827,N_2084,N_2069);
and U2828 (N_2828,N_2166,N_2462);
nand U2829 (N_2829,N_2158,N_2330);
nand U2830 (N_2830,N_2245,N_2369);
and U2831 (N_2831,N_2153,N_2465);
nor U2832 (N_2832,N_2349,N_2438);
xnor U2833 (N_2833,N_2373,N_2362);
nor U2834 (N_2834,N_2237,N_2473);
nand U2835 (N_2835,N_2081,N_2379);
xor U2836 (N_2836,N_2286,N_2447);
nor U2837 (N_2837,N_2101,N_2014);
or U2838 (N_2838,N_2083,N_2040);
nand U2839 (N_2839,N_2463,N_2371);
nand U2840 (N_2840,N_2379,N_2279);
and U2841 (N_2841,N_2279,N_2425);
nor U2842 (N_2842,N_2030,N_2373);
and U2843 (N_2843,N_2325,N_2090);
and U2844 (N_2844,N_2034,N_2280);
and U2845 (N_2845,N_2018,N_2410);
and U2846 (N_2846,N_2483,N_2168);
or U2847 (N_2847,N_2267,N_2127);
and U2848 (N_2848,N_2020,N_2094);
nand U2849 (N_2849,N_2214,N_2258);
or U2850 (N_2850,N_2349,N_2150);
xnor U2851 (N_2851,N_2471,N_2252);
nor U2852 (N_2852,N_2341,N_2399);
nor U2853 (N_2853,N_2195,N_2021);
nand U2854 (N_2854,N_2328,N_2189);
and U2855 (N_2855,N_2140,N_2284);
nand U2856 (N_2856,N_2417,N_2081);
xnor U2857 (N_2857,N_2101,N_2349);
and U2858 (N_2858,N_2201,N_2036);
and U2859 (N_2859,N_2485,N_2411);
nand U2860 (N_2860,N_2309,N_2360);
and U2861 (N_2861,N_2325,N_2094);
xnor U2862 (N_2862,N_2253,N_2325);
nor U2863 (N_2863,N_2122,N_2079);
and U2864 (N_2864,N_2054,N_2052);
nor U2865 (N_2865,N_2458,N_2179);
xor U2866 (N_2866,N_2130,N_2391);
xor U2867 (N_2867,N_2390,N_2150);
or U2868 (N_2868,N_2231,N_2167);
nor U2869 (N_2869,N_2101,N_2294);
or U2870 (N_2870,N_2370,N_2272);
and U2871 (N_2871,N_2436,N_2037);
and U2872 (N_2872,N_2122,N_2194);
and U2873 (N_2873,N_2428,N_2315);
xnor U2874 (N_2874,N_2300,N_2323);
or U2875 (N_2875,N_2386,N_2468);
nand U2876 (N_2876,N_2076,N_2094);
nor U2877 (N_2877,N_2027,N_2061);
nor U2878 (N_2878,N_2204,N_2428);
nor U2879 (N_2879,N_2162,N_2170);
and U2880 (N_2880,N_2408,N_2234);
and U2881 (N_2881,N_2245,N_2492);
and U2882 (N_2882,N_2359,N_2129);
or U2883 (N_2883,N_2420,N_2220);
and U2884 (N_2884,N_2204,N_2025);
or U2885 (N_2885,N_2357,N_2439);
and U2886 (N_2886,N_2037,N_2204);
nor U2887 (N_2887,N_2286,N_2367);
and U2888 (N_2888,N_2094,N_2466);
and U2889 (N_2889,N_2131,N_2130);
nor U2890 (N_2890,N_2221,N_2179);
nor U2891 (N_2891,N_2325,N_2268);
nand U2892 (N_2892,N_2297,N_2269);
or U2893 (N_2893,N_2074,N_2364);
or U2894 (N_2894,N_2124,N_2175);
nor U2895 (N_2895,N_2120,N_2192);
and U2896 (N_2896,N_2056,N_2103);
or U2897 (N_2897,N_2199,N_2260);
nand U2898 (N_2898,N_2312,N_2113);
nand U2899 (N_2899,N_2353,N_2367);
nor U2900 (N_2900,N_2430,N_2168);
nor U2901 (N_2901,N_2225,N_2273);
and U2902 (N_2902,N_2037,N_2183);
xor U2903 (N_2903,N_2151,N_2086);
nor U2904 (N_2904,N_2383,N_2316);
or U2905 (N_2905,N_2292,N_2378);
nor U2906 (N_2906,N_2406,N_2370);
or U2907 (N_2907,N_2403,N_2488);
nor U2908 (N_2908,N_2335,N_2124);
nor U2909 (N_2909,N_2400,N_2334);
and U2910 (N_2910,N_2086,N_2211);
nand U2911 (N_2911,N_2124,N_2348);
nand U2912 (N_2912,N_2151,N_2262);
or U2913 (N_2913,N_2059,N_2489);
xor U2914 (N_2914,N_2445,N_2394);
nor U2915 (N_2915,N_2309,N_2273);
nor U2916 (N_2916,N_2389,N_2403);
nand U2917 (N_2917,N_2325,N_2403);
and U2918 (N_2918,N_2110,N_2444);
nor U2919 (N_2919,N_2010,N_2456);
nor U2920 (N_2920,N_2289,N_2305);
xnor U2921 (N_2921,N_2168,N_2396);
nor U2922 (N_2922,N_2323,N_2486);
and U2923 (N_2923,N_2393,N_2191);
nor U2924 (N_2924,N_2268,N_2022);
nand U2925 (N_2925,N_2461,N_2382);
nor U2926 (N_2926,N_2366,N_2262);
nand U2927 (N_2927,N_2370,N_2451);
and U2928 (N_2928,N_2307,N_2048);
nor U2929 (N_2929,N_2027,N_2235);
and U2930 (N_2930,N_2347,N_2203);
or U2931 (N_2931,N_2415,N_2326);
nand U2932 (N_2932,N_2283,N_2246);
nand U2933 (N_2933,N_2300,N_2193);
nand U2934 (N_2934,N_2303,N_2417);
and U2935 (N_2935,N_2225,N_2399);
and U2936 (N_2936,N_2117,N_2128);
nand U2937 (N_2937,N_2297,N_2328);
nor U2938 (N_2938,N_2477,N_2078);
nor U2939 (N_2939,N_2262,N_2169);
or U2940 (N_2940,N_2239,N_2418);
and U2941 (N_2941,N_2333,N_2158);
nand U2942 (N_2942,N_2033,N_2102);
nor U2943 (N_2943,N_2168,N_2164);
nor U2944 (N_2944,N_2005,N_2375);
nor U2945 (N_2945,N_2312,N_2223);
xor U2946 (N_2946,N_2439,N_2412);
or U2947 (N_2947,N_2493,N_2364);
and U2948 (N_2948,N_2156,N_2427);
nand U2949 (N_2949,N_2173,N_2441);
or U2950 (N_2950,N_2082,N_2245);
or U2951 (N_2951,N_2051,N_2444);
or U2952 (N_2952,N_2492,N_2011);
or U2953 (N_2953,N_2025,N_2166);
nand U2954 (N_2954,N_2061,N_2277);
and U2955 (N_2955,N_2493,N_2297);
nor U2956 (N_2956,N_2020,N_2031);
and U2957 (N_2957,N_2031,N_2475);
and U2958 (N_2958,N_2265,N_2301);
xnor U2959 (N_2959,N_2336,N_2080);
or U2960 (N_2960,N_2179,N_2367);
nand U2961 (N_2961,N_2473,N_2228);
xnor U2962 (N_2962,N_2259,N_2151);
and U2963 (N_2963,N_2452,N_2010);
xor U2964 (N_2964,N_2103,N_2018);
nor U2965 (N_2965,N_2174,N_2162);
nand U2966 (N_2966,N_2193,N_2195);
nor U2967 (N_2967,N_2309,N_2353);
or U2968 (N_2968,N_2366,N_2351);
nand U2969 (N_2969,N_2142,N_2070);
or U2970 (N_2970,N_2482,N_2344);
nor U2971 (N_2971,N_2257,N_2315);
nand U2972 (N_2972,N_2423,N_2196);
nand U2973 (N_2973,N_2020,N_2388);
and U2974 (N_2974,N_2430,N_2426);
or U2975 (N_2975,N_2195,N_2168);
nand U2976 (N_2976,N_2449,N_2321);
and U2977 (N_2977,N_2375,N_2245);
nand U2978 (N_2978,N_2037,N_2363);
nor U2979 (N_2979,N_2448,N_2080);
and U2980 (N_2980,N_2341,N_2088);
and U2981 (N_2981,N_2067,N_2433);
nor U2982 (N_2982,N_2004,N_2142);
nor U2983 (N_2983,N_2213,N_2479);
nand U2984 (N_2984,N_2368,N_2330);
xor U2985 (N_2985,N_2271,N_2208);
nand U2986 (N_2986,N_2015,N_2064);
nand U2987 (N_2987,N_2385,N_2073);
and U2988 (N_2988,N_2373,N_2378);
or U2989 (N_2989,N_2488,N_2373);
nor U2990 (N_2990,N_2042,N_2118);
and U2991 (N_2991,N_2028,N_2078);
or U2992 (N_2992,N_2009,N_2491);
or U2993 (N_2993,N_2360,N_2396);
or U2994 (N_2994,N_2287,N_2261);
or U2995 (N_2995,N_2485,N_2279);
and U2996 (N_2996,N_2225,N_2119);
or U2997 (N_2997,N_2079,N_2290);
nor U2998 (N_2998,N_2436,N_2265);
or U2999 (N_2999,N_2034,N_2447);
nor U3000 (N_3000,N_2524,N_2899);
nor U3001 (N_3001,N_2856,N_2979);
nand U3002 (N_3002,N_2887,N_2951);
nand U3003 (N_3003,N_2853,N_2693);
and U3004 (N_3004,N_2774,N_2850);
and U3005 (N_3005,N_2686,N_2586);
nand U3006 (N_3006,N_2698,N_2817);
nand U3007 (N_3007,N_2878,N_2789);
nand U3008 (N_3008,N_2656,N_2582);
nand U3009 (N_3009,N_2723,N_2990);
and U3010 (N_3010,N_2959,N_2761);
or U3011 (N_3011,N_2812,N_2671);
nor U3012 (N_3012,N_2712,N_2643);
and U3013 (N_3013,N_2766,N_2960);
or U3014 (N_3014,N_2517,N_2785);
nor U3015 (N_3015,N_2673,N_2934);
nor U3016 (N_3016,N_2889,N_2535);
nand U3017 (N_3017,N_2540,N_2772);
nor U3018 (N_3018,N_2971,N_2816);
nand U3019 (N_3019,N_2998,N_2962);
nor U3020 (N_3020,N_2578,N_2746);
nand U3021 (N_3021,N_2957,N_2580);
nor U3022 (N_3022,N_2811,N_2854);
or U3023 (N_3023,N_2777,N_2964);
nand U3024 (N_3024,N_2793,N_2612);
and U3025 (N_3025,N_2776,N_2759);
nor U3026 (N_3026,N_2552,N_2705);
and U3027 (N_3027,N_2700,N_2568);
nand U3028 (N_3028,N_2911,N_2558);
or U3029 (N_3029,N_2943,N_2588);
or U3030 (N_3030,N_2961,N_2839);
nor U3031 (N_3031,N_2630,N_2708);
nor U3032 (N_3032,N_2956,N_2931);
or U3033 (N_3033,N_2841,N_2559);
and U3034 (N_3034,N_2940,N_2923);
or U3035 (N_3035,N_2716,N_2946);
nor U3036 (N_3036,N_2783,N_2954);
or U3037 (N_3037,N_2676,N_2952);
or U3038 (N_3038,N_2840,N_2605);
nor U3039 (N_3039,N_2523,N_2829);
or U3040 (N_3040,N_2626,N_2884);
nor U3041 (N_3041,N_2718,N_2502);
nor U3042 (N_3042,N_2533,N_2832);
nand U3043 (N_3043,N_2751,N_2950);
nor U3044 (N_3044,N_2787,N_2925);
and U3045 (N_3045,N_2664,N_2937);
nor U3046 (N_3046,N_2989,N_2546);
or U3047 (N_3047,N_2598,N_2648);
and U3048 (N_3048,N_2596,N_2587);
or U3049 (N_3049,N_2821,N_2666);
and U3050 (N_3050,N_2973,N_2912);
and U3051 (N_3051,N_2548,N_2702);
and U3052 (N_3052,N_2567,N_2501);
or U3053 (N_3053,N_2909,N_2775);
nand U3054 (N_3054,N_2714,N_2944);
nand U3055 (N_3055,N_2541,N_2755);
or U3056 (N_3056,N_2525,N_2756);
or U3057 (N_3057,N_2624,N_2677);
nor U3058 (N_3058,N_2881,N_2851);
nor U3059 (N_3059,N_2947,N_2688);
and U3060 (N_3060,N_2830,N_2976);
nand U3061 (N_3061,N_2768,N_2527);
or U3062 (N_3062,N_2738,N_2597);
and U3063 (N_3063,N_2948,N_2575);
nand U3064 (N_3064,N_2683,N_2724);
xnor U3065 (N_3065,N_2675,N_2507);
or U3066 (N_3066,N_2823,N_2642);
nor U3067 (N_3067,N_2640,N_2604);
nand U3068 (N_3068,N_2510,N_2995);
nand U3069 (N_3069,N_2985,N_2696);
and U3070 (N_3070,N_2868,N_2584);
or U3071 (N_3071,N_2667,N_2992);
and U3072 (N_3072,N_2606,N_2543);
nand U3073 (N_3073,N_2572,N_2986);
nor U3074 (N_3074,N_2529,N_2621);
nor U3075 (N_3075,N_2844,N_2906);
and U3076 (N_3076,N_2554,N_2945);
or U3077 (N_3077,N_2625,N_2691);
nor U3078 (N_3078,N_2663,N_2734);
and U3079 (N_3079,N_2904,N_2860);
nor U3080 (N_3080,N_2503,N_2883);
nand U3081 (N_3081,N_2634,N_2874);
nand U3082 (N_3082,N_2993,N_2719);
nor U3083 (N_3083,N_2968,N_2910);
nand U3084 (N_3084,N_2707,N_2660);
and U3085 (N_3085,N_2566,N_2848);
xnor U3086 (N_3086,N_2922,N_2736);
or U3087 (N_3087,N_2530,N_2647);
xor U3088 (N_3088,N_2828,N_2873);
xor U3089 (N_3089,N_2935,N_2891);
nor U3090 (N_3090,N_2933,N_2875);
xor U3091 (N_3091,N_2689,N_2824);
or U3092 (N_3092,N_2609,N_2877);
nand U3093 (N_3093,N_2845,N_2652);
xor U3094 (N_3094,N_2542,N_2728);
or U3095 (N_3095,N_2921,N_2886);
nand U3096 (N_3096,N_2905,N_2740);
nand U3097 (N_3097,N_2651,N_2915);
xnor U3098 (N_3098,N_2966,N_2805);
and U3099 (N_3099,N_2928,N_2784);
xnor U3100 (N_3100,N_2769,N_2791);
xor U3101 (N_3101,N_2802,N_2919);
nand U3102 (N_3102,N_2749,N_2767);
nor U3103 (N_3103,N_2778,N_2722);
nand U3104 (N_3104,N_2629,N_2916);
and U3105 (N_3105,N_2846,N_2773);
xnor U3106 (N_3106,N_2720,N_2872);
or U3107 (N_3107,N_2650,N_2508);
or U3108 (N_3108,N_2879,N_2589);
or U3109 (N_3109,N_2594,N_2645);
and U3110 (N_3110,N_2654,N_2792);
nor U3111 (N_3111,N_2764,N_2936);
and U3112 (N_3112,N_2638,N_2996);
nand U3113 (N_3113,N_2975,N_2795);
xor U3114 (N_3114,N_2744,N_2796);
and U3115 (N_3115,N_2619,N_2701);
or U3116 (N_3116,N_2512,N_2521);
nor U3117 (N_3117,N_2892,N_2509);
and U3118 (N_3118,N_2893,N_2842);
and U3119 (N_3119,N_2713,N_2780);
nand U3120 (N_3120,N_2799,N_2516);
or U3121 (N_3121,N_2852,N_2843);
and U3122 (N_3122,N_2685,N_2704);
nand U3123 (N_3123,N_2513,N_2963);
and U3124 (N_3124,N_2741,N_2818);
nand U3125 (N_3125,N_2978,N_2635);
or U3126 (N_3126,N_2551,N_2731);
nor U3127 (N_3127,N_2585,N_2896);
nor U3128 (N_3128,N_2833,N_2890);
nand U3129 (N_3129,N_2574,N_2555);
nand U3130 (N_3130,N_2536,N_2939);
nor U3131 (N_3131,N_2977,N_2514);
or U3132 (N_3132,N_2620,N_2593);
nand U3133 (N_3133,N_2581,N_2646);
nor U3134 (N_3134,N_2888,N_2825);
nor U3135 (N_3135,N_2725,N_2902);
nand U3136 (N_3136,N_2537,N_2601);
or U3137 (N_3137,N_2680,N_2608);
nor U3138 (N_3138,N_2699,N_2927);
nand U3139 (N_3139,N_2562,N_2864);
or U3140 (N_3140,N_2733,N_2924);
or U3141 (N_3141,N_2897,N_2991);
nand U3142 (N_3142,N_2855,N_2579);
or U3143 (N_3143,N_2970,N_2622);
nand U3144 (N_3144,N_2511,N_2721);
or U3145 (N_3145,N_2831,N_2982);
xnor U3146 (N_3146,N_2687,N_2758);
nand U3147 (N_3147,N_2763,N_2617);
xnor U3148 (N_3148,N_2703,N_2836);
nor U3149 (N_3149,N_2506,N_2932);
or U3150 (N_3150,N_2739,N_2797);
nor U3151 (N_3151,N_2747,N_2870);
nand U3152 (N_3152,N_2637,N_2727);
and U3153 (N_3153,N_2706,N_2735);
nor U3154 (N_3154,N_2732,N_2591);
or U3155 (N_3155,N_2742,N_2900);
and U3156 (N_3156,N_2590,N_2658);
or U3157 (N_3157,N_2849,N_2710);
and U3158 (N_3158,N_2903,N_2611);
nor U3159 (N_3159,N_2561,N_2790);
nand U3160 (N_3160,N_2520,N_2965);
nand U3161 (N_3161,N_2807,N_2865);
nand U3162 (N_3162,N_2942,N_2941);
nand U3163 (N_3163,N_2798,N_2618);
or U3164 (N_3164,N_2684,N_2955);
and U3165 (N_3165,N_2500,N_2754);
xnor U3166 (N_3166,N_2743,N_2560);
nor U3167 (N_3167,N_2639,N_2837);
and U3168 (N_3168,N_2610,N_2682);
and U3169 (N_3169,N_2988,N_2665);
or U3170 (N_3170,N_2760,N_2657);
nor U3171 (N_3171,N_2649,N_2592);
nand U3172 (N_3172,N_2984,N_2859);
or U3173 (N_3173,N_2800,N_2871);
or U3174 (N_3174,N_2709,N_2869);
nor U3175 (N_3175,N_2974,N_2858);
nor U3176 (N_3176,N_2599,N_2518);
xor U3177 (N_3177,N_2697,N_2644);
nand U3178 (N_3178,N_2505,N_2679);
nand U3179 (N_3179,N_2810,N_2894);
nand U3180 (N_3180,N_2577,N_2534);
or U3181 (N_3181,N_2715,N_2573);
nor U3182 (N_3182,N_2804,N_2981);
and U3183 (N_3183,N_2822,N_2814);
xor U3184 (N_3184,N_2504,N_2930);
nor U3185 (N_3185,N_2929,N_2678);
xor U3186 (N_3186,N_2867,N_2600);
and U3187 (N_3187,N_2895,N_2813);
nand U3188 (N_3188,N_2882,N_2913);
or U3189 (N_3189,N_2987,N_2757);
nand U3190 (N_3190,N_2519,N_2616);
or U3191 (N_3191,N_2958,N_2781);
or U3192 (N_3192,N_2834,N_2603);
nand U3193 (N_3193,N_2917,N_2539);
nand U3194 (N_3194,N_2794,N_2806);
nand U3195 (N_3195,N_2627,N_2730);
nor U3196 (N_3196,N_2690,N_2711);
nor U3197 (N_3197,N_2633,N_2557);
nor U3198 (N_3198,N_2569,N_2564);
nand U3199 (N_3199,N_2655,N_2827);
and U3200 (N_3200,N_2885,N_2576);
nor U3201 (N_3201,N_2613,N_2623);
and U3202 (N_3202,N_2692,N_2726);
nor U3203 (N_3203,N_2750,N_2994);
nand U3204 (N_3204,N_2583,N_2819);
or U3205 (N_3205,N_2628,N_2661);
nand U3206 (N_3206,N_2636,N_2920);
and U3207 (N_3207,N_2570,N_2602);
nor U3208 (N_3208,N_2969,N_2967);
xor U3209 (N_3209,N_2765,N_2926);
nor U3210 (N_3210,N_2762,N_2876);
or U3211 (N_3211,N_2908,N_2820);
nand U3212 (N_3212,N_2531,N_2545);
nand U3213 (N_3213,N_2809,N_2528);
or U3214 (N_3214,N_2786,N_2808);
and U3215 (N_3215,N_2681,N_2826);
nand U3216 (N_3216,N_2753,N_2737);
nand U3217 (N_3217,N_2779,N_2641);
nand U3218 (N_3218,N_2631,N_2550);
nand U3219 (N_3219,N_2972,N_2771);
and U3220 (N_3220,N_2847,N_2953);
and U3221 (N_3221,N_2803,N_2669);
xor U3222 (N_3222,N_2632,N_2980);
nor U3223 (N_3223,N_2668,N_2788);
nor U3224 (N_3224,N_2938,N_2614);
xor U3225 (N_3225,N_2556,N_2862);
nand U3226 (N_3226,N_2752,N_2532);
nand U3227 (N_3227,N_2918,N_2695);
and U3228 (N_3228,N_2553,N_2674);
nand U3229 (N_3229,N_2729,N_2694);
nor U3230 (N_3230,N_2672,N_2983);
and U3231 (N_3231,N_2782,N_2857);
xnor U3232 (N_3232,N_2653,N_2880);
and U3233 (N_3233,N_2949,N_2999);
nand U3234 (N_3234,N_2717,N_2748);
nor U3235 (N_3235,N_2770,N_2549);
xor U3236 (N_3236,N_2866,N_2861);
or U3237 (N_3237,N_2538,N_2914);
nor U3238 (N_3238,N_2571,N_2670);
or U3239 (N_3239,N_2515,N_2526);
nand U3240 (N_3240,N_2898,N_2522);
nand U3241 (N_3241,N_2907,N_2863);
or U3242 (N_3242,N_2997,N_2835);
xor U3243 (N_3243,N_2801,N_2607);
and U3244 (N_3244,N_2565,N_2544);
nand U3245 (N_3245,N_2838,N_2662);
nand U3246 (N_3246,N_2745,N_2615);
nor U3247 (N_3247,N_2595,N_2563);
or U3248 (N_3248,N_2901,N_2815);
nand U3249 (N_3249,N_2659,N_2547);
or U3250 (N_3250,N_2993,N_2533);
nor U3251 (N_3251,N_2817,N_2694);
and U3252 (N_3252,N_2979,N_2959);
nand U3253 (N_3253,N_2586,N_2811);
nand U3254 (N_3254,N_2732,N_2716);
and U3255 (N_3255,N_2884,N_2920);
and U3256 (N_3256,N_2813,N_2569);
nor U3257 (N_3257,N_2787,N_2518);
and U3258 (N_3258,N_2838,N_2642);
nand U3259 (N_3259,N_2637,N_2677);
and U3260 (N_3260,N_2791,N_2508);
nand U3261 (N_3261,N_2748,N_2810);
and U3262 (N_3262,N_2731,N_2845);
nand U3263 (N_3263,N_2686,N_2875);
and U3264 (N_3264,N_2817,N_2897);
or U3265 (N_3265,N_2833,N_2693);
nor U3266 (N_3266,N_2679,N_2741);
and U3267 (N_3267,N_2652,N_2585);
and U3268 (N_3268,N_2703,N_2957);
or U3269 (N_3269,N_2703,N_2719);
nor U3270 (N_3270,N_2539,N_2808);
nor U3271 (N_3271,N_2985,N_2594);
xor U3272 (N_3272,N_2558,N_2854);
or U3273 (N_3273,N_2974,N_2967);
and U3274 (N_3274,N_2637,N_2661);
and U3275 (N_3275,N_2669,N_2588);
and U3276 (N_3276,N_2589,N_2631);
or U3277 (N_3277,N_2564,N_2515);
nor U3278 (N_3278,N_2540,N_2637);
nor U3279 (N_3279,N_2603,N_2946);
or U3280 (N_3280,N_2655,N_2805);
nor U3281 (N_3281,N_2593,N_2585);
nor U3282 (N_3282,N_2999,N_2501);
nand U3283 (N_3283,N_2627,N_2719);
nor U3284 (N_3284,N_2558,N_2660);
or U3285 (N_3285,N_2793,N_2535);
nor U3286 (N_3286,N_2789,N_2647);
or U3287 (N_3287,N_2936,N_2872);
and U3288 (N_3288,N_2904,N_2954);
nor U3289 (N_3289,N_2537,N_2894);
nor U3290 (N_3290,N_2803,N_2798);
nand U3291 (N_3291,N_2926,N_2712);
and U3292 (N_3292,N_2899,N_2968);
nor U3293 (N_3293,N_2975,N_2770);
or U3294 (N_3294,N_2992,N_2637);
nor U3295 (N_3295,N_2551,N_2936);
nor U3296 (N_3296,N_2924,N_2804);
and U3297 (N_3297,N_2545,N_2956);
and U3298 (N_3298,N_2585,N_2578);
nand U3299 (N_3299,N_2601,N_2783);
xor U3300 (N_3300,N_2551,N_2595);
and U3301 (N_3301,N_2534,N_2678);
nand U3302 (N_3302,N_2868,N_2514);
nand U3303 (N_3303,N_2841,N_2959);
nand U3304 (N_3304,N_2525,N_2611);
nor U3305 (N_3305,N_2901,N_2705);
nand U3306 (N_3306,N_2789,N_2521);
or U3307 (N_3307,N_2626,N_2945);
and U3308 (N_3308,N_2981,N_2978);
xor U3309 (N_3309,N_2937,N_2767);
and U3310 (N_3310,N_2749,N_2722);
and U3311 (N_3311,N_2701,N_2922);
and U3312 (N_3312,N_2663,N_2755);
nor U3313 (N_3313,N_2931,N_2656);
nor U3314 (N_3314,N_2778,N_2608);
and U3315 (N_3315,N_2999,N_2940);
xnor U3316 (N_3316,N_2645,N_2551);
nand U3317 (N_3317,N_2524,N_2816);
nand U3318 (N_3318,N_2884,N_2612);
nand U3319 (N_3319,N_2796,N_2536);
or U3320 (N_3320,N_2994,N_2797);
and U3321 (N_3321,N_2691,N_2610);
or U3322 (N_3322,N_2647,N_2600);
nor U3323 (N_3323,N_2949,N_2570);
or U3324 (N_3324,N_2706,N_2704);
or U3325 (N_3325,N_2925,N_2951);
nor U3326 (N_3326,N_2844,N_2891);
xor U3327 (N_3327,N_2768,N_2841);
nand U3328 (N_3328,N_2819,N_2827);
or U3329 (N_3329,N_2568,N_2740);
nand U3330 (N_3330,N_2751,N_2982);
nor U3331 (N_3331,N_2654,N_2517);
nand U3332 (N_3332,N_2840,N_2563);
and U3333 (N_3333,N_2634,N_2901);
nor U3334 (N_3334,N_2942,N_2972);
xnor U3335 (N_3335,N_2798,N_2511);
or U3336 (N_3336,N_2959,N_2937);
or U3337 (N_3337,N_2596,N_2757);
nor U3338 (N_3338,N_2936,N_2813);
and U3339 (N_3339,N_2769,N_2821);
nand U3340 (N_3340,N_2538,N_2539);
and U3341 (N_3341,N_2638,N_2551);
and U3342 (N_3342,N_2776,N_2620);
nor U3343 (N_3343,N_2604,N_2556);
and U3344 (N_3344,N_2783,N_2709);
and U3345 (N_3345,N_2509,N_2839);
or U3346 (N_3346,N_2744,N_2745);
nor U3347 (N_3347,N_2714,N_2642);
nand U3348 (N_3348,N_2974,N_2776);
or U3349 (N_3349,N_2524,N_2780);
and U3350 (N_3350,N_2996,N_2878);
or U3351 (N_3351,N_2865,N_2848);
or U3352 (N_3352,N_2864,N_2792);
and U3353 (N_3353,N_2519,N_2792);
and U3354 (N_3354,N_2790,N_2969);
and U3355 (N_3355,N_2879,N_2586);
or U3356 (N_3356,N_2560,N_2571);
or U3357 (N_3357,N_2943,N_2748);
and U3358 (N_3358,N_2564,N_2630);
and U3359 (N_3359,N_2790,N_2973);
and U3360 (N_3360,N_2908,N_2846);
and U3361 (N_3361,N_2778,N_2733);
and U3362 (N_3362,N_2821,N_2819);
nand U3363 (N_3363,N_2995,N_2839);
or U3364 (N_3364,N_2996,N_2907);
nand U3365 (N_3365,N_2539,N_2936);
or U3366 (N_3366,N_2577,N_2679);
xor U3367 (N_3367,N_2973,N_2621);
and U3368 (N_3368,N_2819,N_2806);
and U3369 (N_3369,N_2638,N_2833);
or U3370 (N_3370,N_2779,N_2660);
xor U3371 (N_3371,N_2771,N_2955);
nand U3372 (N_3372,N_2894,N_2987);
nor U3373 (N_3373,N_2625,N_2717);
nor U3374 (N_3374,N_2770,N_2589);
nor U3375 (N_3375,N_2652,N_2973);
and U3376 (N_3376,N_2892,N_2772);
or U3377 (N_3377,N_2642,N_2658);
and U3378 (N_3378,N_2722,N_2783);
xnor U3379 (N_3379,N_2845,N_2997);
or U3380 (N_3380,N_2595,N_2580);
nand U3381 (N_3381,N_2925,N_2893);
nor U3382 (N_3382,N_2779,N_2958);
and U3383 (N_3383,N_2900,N_2721);
or U3384 (N_3384,N_2774,N_2524);
or U3385 (N_3385,N_2715,N_2774);
nand U3386 (N_3386,N_2808,N_2834);
and U3387 (N_3387,N_2724,N_2535);
or U3388 (N_3388,N_2818,N_2680);
nor U3389 (N_3389,N_2640,N_2688);
nor U3390 (N_3390,N_2682,N_2505);
or U3391 (N_3391,N_2845,N_2512);
nor U3392 (N_3392,N_2573,N_2598);
nor U3393 (N_3393,N_2765,N_2619);
and U3394 (N_3394,N_2993,N_2858);
nor U3395 (N_3395,N_2663,N_2558);
and U3396 (N_3396,N_2654,N_2769);
nor U3397 (N_3397,N_2801,N_2940);
nand U3398 (N_3398,N_2919,N_2616);
nor U3399 (N_3399,N_2802,N_2697);
and U3400 (N_3400,N_2711,N_2573);
nor U3401 (N_3401,N_2932,N_2703);
and U3402 (N_3402,N_2542,N_2683);
nor U3403 (N_3403,N_2653,N_2681);
nor U3404 (N_3404,N_2809,N_2643);
nor U3405 (N_3405,N_2719,N_2725);
nand U3406 (N_3406,N_2675,N_2830);
nor U3407 (N_3407,N_2695,N_2791);
and U3408 (N_3408,N_2771,N_2927);
nor U3409 (N_3409,N_2560,N_2877);
nand U3410 (N_3410,N_2503,N_2512);
or U3411 (N_3411,N_2891,N_2858);
nand U3412 (N_3412,N_2924,N_2994);
nor U3413 (N_3413,N_2612,N_2636);
and U3414 (N_3414,N_2642,N_2908);
or U3415 (N_3415,N_2549,N_2531);
nand U3416 (N_3416,N_2906,N_2536);
xnor U3417 (N_3417,N_2633,N_2661);
and U3418 (N_3418,N_2803,N_2838);
nor U3419 (N_3419,N_2613,N_2544);
nor U3420 (N_3420,N_2582,N_2750);
or U3421 (N_3421,N_2649,N_2623);
and U3422 (N_3422,N_2689,N_2776);
nand U3423 (N_3423,N_2605,N_2686);
and U3424 (N_3424,N_2725,N_2588);
or U3425 (N_3425,N_2766,N_2949);
nand U3426 (N_3426,N_2601,N_2849);
nand U3427 (N_3427,N_2818,N_2728);
or U3428 (N_3428,N_2666,N_2720);
nand U3429 (N_3429,N_2783,N_2698);
nor U3430 (N_3430,N_2854,N_2848);
nand U3431 (N_3431,N_2755,N_2638);
and U3432 (N_3432,N_2752,N_2518);
and U3433 (N_3433,N_2889,N_2802);
nor U3434 (N_3434,N_2723,N_2840);
or U3435 (N_3435,N_2919,N_2801);
nor U3436 (N_3436,N_2645,N_2539);
nor U3437 (N_3437,N_2581,N_2687);
or U3438 (N_3438,N_2792,N_2934);
and U3439 (N_3439,N_2590,N_2829);
xor U3440 (N_3440,N_2654,N_2922);
and U3441 (N_3441,N_2728,N_2517);
nor U3442 (N_3442,N_2946,N_2973);
nor U3443 (N_3443,N_2613,N_2925);
nor U3444 (N_3444,N_2717,N_2937);
or U3445 (N_3445,N_2840,N_2629);
or U3446 (N_3446,N_2987,N_2996);
or U3447 (N_3447,N_2516,N_2995);
nand U3448 (N_3448,N_2832,N_2731);
or U3449 (N_3449,N_2916,N_2830);
or U3450 (N_3450,N_2862,N_2632);
nor U3451 (N_3451,N_2690,N_2516);
nand U3452 (N_3452,N_2911,N_2852);
or U3453 (N_3453,N_2579,N_2701);
nor U3454 (N_3454,N_2875,N_2527);
nand U3455 (N_3455,N_2893,N_2942);
nand U3456 (N_3456,N_2512,N_2864);
and U3457 (N_3457,N_2556,N_2528);
nand U3458 (N_3458,N_2929,N_2669);
and U3459 (N_3459,N_2980,N_2737);
xnor U3460 (N_3460,N_2631,N_2551);
nor U3461 (N_3461,N_2571,N_2887);
or U3462 (N_3462,N_2649,N_2721);
or U3463 (N_3463,N_2596,N_2841);
nand U3464 (N_3464,N_2890,N_2791);
and U3465 (N_3465,N_2957,N_2919);
nor U3466 (N_3466,N_2653,N_2826);
and U3467 (N_3467,N_2642,N_2939);
and U3468 (N_3468,N_2972,N_2867);
and U3469 (N_3469,N_2974,N_2659);
xnor U3470 (N_3470,N_2923,N_2711);
nand U3471 (N_3471,N_2796,N_2933);
or U3472 (N_3472,N_2682,N_2931);
nand U3473 (N_3473,N_2595,N_2518);
nor U3474 (N_3474,N_2983,N_2994);
nand U3475 (N_3475,N_2602,N_2731);
nor U3476 (N_3476,N_2659,N_2836);
nor U3477 (N_3477,N_2553,N_2551);
and U3478 (N_3478,N_2813,N_2829);
xor U3479 (N_3479,N_2865,N_2557);
or U3480 (N_3480,N_2851,N_2580);
or U3481 (N_3481,N_2899,N_2962);
and U3482 (N_3482,N_2554,N_2865);
or U3483 (N_3483,N_2976,N_2822);
and U3484 (N_3484,N_2565,N_2909);
or U3485 (N_3485,N_2544,N_2744);
nand U3486 (N_3486,N_2609,N_2565);
or U3487 (N_3487,N_2536,N_2698);
nand U3488 (N_3488,N_2784,N_2591);
nand U3489 (N_3489,N_2634,N_2833);
and U3490 (N_3490,N_2639,N_2919);
and U3491 (N_3491,N_2904,N_2997);
or U3492 (N_3492,N_2749,N_2744);
nor U3493 (N_3493,N_2771,N_2977);
xor U3494 (N_3494,N_2820,N_2771);
or U3495 (N_3495,N_2563,N_2907);
nand U3496 (N_3496,N_2892,N_2938);
nor U3497 (N_3497,N_2752,N_2581);
nor U3498 (N_3498,N_2965,N_2761);
nor U3499 (N_3499,N_2873,N_2911);
and U3500 (N_3500,N_3260,N_3040);
nand U3501 (N_3501,N_3097,N_3294);
or U3502 (N_3502,N_3397,N_3210);
nor U3503 (N_3503,N_3201,N_3332);
nor U3504 (N_3504,N_3217,N_3281);
or U3505 (N_3505,N_3062,N_3231);
nor U3506 (N_3506,N_3354,N_3013);
or U3507 (N_3507,N_3186,N_3096);
and U3508 (N_3508,N_3079,N_3483);
nor U3509 (N_3509,N_3041,N_3431);
and U3510 (N_3510,N_3365,N_3447);
or U3511 (N_3511,N_3232,N_3136);
and U3512 (N_3512,N_3064,N_3081);
or U3513 (N_3513,N_3463,N_3128);
and U3514 (N_3514,N_3443,N_3479);
or U3515 (N_3515,N_3492,N_3026);
and U3516 (N_3516,N_3140,N_3270);
or U3517 (N_3517,N_3047,N_3314);
or U3518 (N_3518,N_3056,N_3187);
nor U3519 (N_3519,N_3240,N_3373);
nor U3520 (N_3520,N_3082,N_3024);
nand U3521 (N_3521,N_3057,N_3122);
and U3522 (N_3522,N_3341,N_3449);
nor U3523 (N_3523,N_3366,N_3299);
and U3524 (N_3524,N_3486,N_3415);
nand U3525 (N_3525,N_3351,N_3403);
or U3526 (N_3526,N_3093,N_3285);
nand U3527 (N_3527,N_3413,N_3138);
or U3528 (N_3528,N_3021,N_3275);
nand U3529 (N_3529,N_3301,N_3368);
nor U3530 (N_3530,N_3491,N_3359);
or U3531 (N_3531,N_3429,N_3146);
nor U3532 (N_3532,N_3052,N_3267);
and U3533 (N_3533,N_3315,N_3465);
or U3534 (N_3534,N_3350,N_3302);
and U3535 (N_3535,N_3099,N_3205);
nor U3536 (N_3536,N_3139,N_3177);
and U3537 (N_3537,N_3494,N_3174);
and U3538 (N_3538,N_3110,N_3434);
nor U3539 (N_3539,N_3360,N_3002);
and U3540 (N_3540,N_3418,N_3025);
nand U3541 (N_3541,N_3220,N_3208);
nor U3542 (N_3542,N_3063,N_3305);
nor U3543 (N_3543,N_3230,N_3171);
nand U3544 (N_3544,N_3181,N_3043);
and U3545 (N_3545,N_3312,N_3286);
or U3546 (N_3546,N_3141,N_3192);
nor U3547 (N_3547,N_3420,N_3225);
or U3548 (N_3548,N_3298,N_3241);
and U3549 (N_3549,N_3103,N_3007);
nand U3550 (N_3550,N_3251,N_3334);
or U3551 (N_3551,N_3392,N_3437);
nor U3552 (N_3552,N_3129,N_3321);
and U3553 (N_3553,N_3133,N_3006);
and U3554 (N_3554,N_3318,N_3436);
xor U3555 (N_3555,N_3349,N_3358);
nor U3556 (N_3556,N_3460,N_3451);
nor U3557 (N_3557,N_3071,N_3410);
nor U3558 (N_3558,N_3094,N_3084);
and U3559 (N_3559,N_3475,N_3377);
or U3560 (N_3560,N_3073,N_3066);
nor U3561 (N_3561,N_3107,N_3467);
nand U3562 (N_3562,N_3183,N_3018);
nand U3563 (N_3563,N_3149,N_3037);
or U3564 (N_3564,N_3167,N_3031);
nor U3565 (N_3565,N_3404,N_3078);
nand U3566 (N_3566,N_3269,N_3060);
nand U3567 (N_3567,N_3009,N_3042);
nand U3568 (N_3568,N_3045,N_3379);
nand U3569 (N_3569,N_3249,N_3488);
nand U3570 (N_3570,N_3331,N_3454);
nand U3571 (N_3571,N_3384,N_3333);
and U3572 (N_3572,N_3307,N_3200);
nor U3573 (N_3573,N_3310,N_3381);
and U3574 (N_3574,N_3126,N_3123);
and U3575 (N_3575,N_3356,N_3424);
nand U3576 (N_3576,N_3320,N_3058);
or U3577 (N_3577,N_3419,N_3295);
or U3578 (N_3578,N_3154,N_3046);
xnor U3579 (N_3579,N_3471,N_3190);
or U3580 (N_3580,N_3343,N_3124);
or U3581 (N_3581,N_3109,N_3196);
nand U3582 (N_3582,N_3422,N_3452);
or U3583 (N_3583,N_3189,N_3003);
nor U3584 (N_3584,N_3014,N_3290);
or U3585 (N_3585,N_3322,N_3206);
or U3586 (N_3586,N_3474,N_3478);
nand U3587 (N_3587,N_3236,N_3409);
or U3588 (N_3588,N_3158,N_3257);
nand U3589 (N_3589,N_3383,N_3182);
and U3590 (N_3590,N_3219,N_3423);
nor U3591 (N_3591,N_3179,N_3070);
and U3592 (N_3592,N_3276,N_3498);
or U3593 (N_3593,N_3484,N_3345);
nor U3594 (N_3594,N_3222,N_3265);
xnor U3595 (N_3595,N_3145,N_3442);
and U3596 (N_3596,N_3405,N_3044);
and U3597 (N_3597,N_3076,N_3304);
nor U3598 (N_3598,N_3153,N_3135);
nor U3599 (N_3599,N_3371,N_3185);
and U3600 (N_3600,N_3395,N_3490);
nor U3601 (N_3601,N_3370,N_3472);
nand U3602 (N_3602,N_3367,N_3155);
nor U3603 (N_3603,N_3407,N_3168);
nor U3604 (N_3604,N_3184,N_3016);
nor U3605 (N_3605,N_3375,N_3316);
xor U3606 (N_3606,N_3291,N_3357);
and U3607 (N_3607,N_3271,N_3401);
xnor U3608 (N_3608,N_3117,N_3380);
or U3609 (N_3609,N_3067,N_3180);
or U3610 (N_3610,N_3289,N_3309);
and U3611 (N_3611,N_3188,N_3280);
nand U3612 (N_3612,N_3198,N_3215);
nand U3613 (N_3613,N_3085,N_3459);
or U3614 (N_3614,N_3416,N_3191);
xor U3615 (N_3615,N_3017,N_3391);
nand U3616 (N_3616,N_3378,N_3212);
and U3617 (N_3617,N_3163,N_3273);
xor U3618 (N_3618,N_3106,N_3160);
nand U3619 (N_3619,N_3150,N_3104);
nand U3620 (N_3620,N_3036,N_3015);
nand U3621 (N_3621,N_3033,N_3010);
and U3622 (N_3622,N_3469,N_3313);
and U3623 (N_3623,N_3004,N_3340);
nand U3624 (N_3624,N_3376,N_3054);
nor U3625 (N_3625,N_3468,N_3161);
or U3626 (N_3626,N_3347,N_3226);
nand U3627 (N_3627,N_3243,N_3261);
nand U3628 (N_3628,N_3132,N_3121);
nor U3629 (N_3629,N_3242,N_3252);
and U3630 (N_3630,N_3446,N_3069);
and U3631 (N_3631,N_3089,N_3458);
nor U3632 (N_3632,N_3466,N_3116);
or U3633 (N_3633,N_3450,N_3115);
nand U3634 (N_3634,N_3428,N_3142);
nor U3635 (N_3635,N_3344,N_3259);
nor U3636 (N_3636,N_3156,N_3455);
or U3637 (N_3637,N_3427,N_3120);
and U3638 (N_3638,N_3254,N_3338);
xor U3639 (N_3639,N_3329,N_3032);
or U3640 (N_3640,N_3143,N_3008);
nand U3641 (N_3641,N_3218,N_3030);
xnor U3642 (N_3642,N_3342,N_3296);
or U3643 (N_3643,N_3051,N_3087);
or U3644 (N_3644,N_3091,N_3489);
nor U3645 (N_3645,N_3176,N_3199);
xnor U3646 (N_3646,N_3300,N_3382);
nor U3647 (N_3647,N_3250,N_3207);
or U3648 (N_3648,N_3336,N_3476);
and U3649 (N_3649,N_3086,N_3435);
nor U3650 (N_3650,N_3430,N_3448);
nand U3651 (N_3651,N_3131,N_3499);
nand U3652 (N_3652,N_3134,N_3393);
nor U3653 (N_3653,N_3352,N_3480);
nand U3654 (N_3654,N_3414,N_3202);
or U3655 (N_3655,N_3213,N_3027);
and U3656 (N_3656,N_3053,N_3247);
and U3657 (N_3657,N_3330,N_3092);
xnor U3658 (N_3658,N_3111,N_3193);
xnor U3659 (N_3659,N_3119,N_3496);
nor U3660 (N_3660,N_3353,N_3012);
and U3661 (N_3661,N_3061,N_3147);
nand U3662 (N_3662,N_3152,N_3229);
nor U3663 (N_3663,N_3049,N_3438);
or U3664 (N_3664,N_3137,N_3234);
nand U3665 (N_3665,N_3464,N_3398);
or U3666 (N_3666,N_3239,N_3317);
nand U3667 (N_3667,N_3461,N_3402);
nor U3668 (N_3668,N_3172,N_3157);
nor U3669 (N_3669,N_3346,N_3385);
nor U3670 (N_3670,N_3194,N_3493);
and U3671 (N_3671,N_3195,N_3074);
and U3672 (N_3672,N_3263,N_3369);
nand U3673 (N_3673,N_3283,N_3297);
nand U3674 (N_3674,N_3266,N_3005);
nor U3675 (N_3675,N_3090,N_3439);
nor U3676 (N_3676,N_3209,N_3457);
nor U3677 (N_3677,N_3151,N_3228);
nand U3678 (N_3678,N_3374,N_3456);
nand U3679 (N_3679,N_3324,N_3125);
nand U3680 (N_3680,N_3170,N_3077);
and U3681 (N_3681,N_3068,N_3244);
or U3682 (N_3682,N_3287,N_3308);
nand U3683 (N_3683,N_3325,N_3328);
or U3684 (N_3684,N_3274,N_3178);
xnor U3685 (N_3685,N_3306,N_3337);
nor U3686 (N_3686,N_3433,N_3165);
nand U3687 (N_3687,N_3127,N_3001);
xnor U3688 (N_3688,N_3175,N_3130);
or U3689 (N_3689,N_3453,N_3164);
xnor U3690 (N_3690,N_3237,N_3028);
nor U3691 (N_3691,N_3432,N_3390);
and U3692 (N_3692,N_3264,N_3169);
xnor U3693 (N_3693,N_3497,N_3262);
nor U3694 (N_3694,N_3386,N_3412);
nor U3695 (N_3695,N_3495,N_3477);
xor U3696 (N_3696,N_3440,N_3470);
and U3697 (N_3697,N_3361,N_3098);
nor U3698 (N_3698,N_3268,N_3323);
nor U3699 (N_3699,N_3444,N_3293);
or U3700 (N_3700,N_3059,N_3114);
nor U3701 (N_3701,N_3339,N_3039);
nand U3702 (N_3702,N_3399,N_3364);
nor U3703 (N_3703,N_3288,N_3029);
nor U3704 (N_3704,N_3034,N_3481);
or U3705 (N_3705,N_3072,N_3303);
nor U3706 (N_3706,N_3023,N_3000);
or U3707 (N_3707,N_3389,N_3417);
nor U3708 (N_3708,N_3400,N_3487);
nand U3709 (N_3709,N_3105,N_3223);
or U3710 (N_3710,N_3372,N_3144);
nor U3711 (N_3711,N_3075,N_3335);
xnor U3712 (N_3712,N_3095,N_3482);
xnor U3713 (N_3713,N_3203,N_3355);
nand U3714 (N_3714,N_3396,N_3445);
and U3715 (N_3715,N_3113,N_3020);
or U3716 (N_3716,N_3035,N_3284);
or U3717 (N_3717,N_3227,N_3282);
xor U3718 (N_3718,N_3235,N_3327);
and U3719 (N_3719,N_3233,N_3473);
nor U3720 (N_3720,N_3248,N_3204);
xor U3721 (N_3721,N_3425,N_3162);
and U3722 (N_3722,N_3394,N_3362);
or U3723 (N_3723,N_3311,N_3173);
or U3724 (N_3724,N_3388,N_3148);
nand U3725 (N_3725,N_3238,N_3019);
nor U3726 (N_3726,N_3485,N_3245);
and U3727 (N_3727,N_3100,N_3216);
nand U3728 (N_3728,N_3348,N_3065);
nor U3729 (N_3729,N_3277,N_3255);
or U3730 (N_3730,N_3406,N_3278);
and U3731 (N_3731,N_3272,N_3011);
and U3732 (N_3732,N_3462,N_3197);
and U3733 (N_3733,N_3083,N_3080);
and U3734 (N_3734,N_3038,N_3022);
nor U3735 (N_3735,N_3166,N_3319);
or U3736 (N_3736,N_3214,N_3050);
or U3737 (N_3737,N_3279,N_3221);
or U3738 (N_3738,N_3112,N_3411);
or U3739 (N_3739,N_3253,N_3118);
nand U3740 (N_3740,N_3292,N_3108);
nand U3741 (N_3741,N_3102,N_3441);
or U3742 (N_3742,N_3408,N_3246);
nand U3743 (N_3743,N_3101,N_3387);
xor U3744 (N_3744,N_3055,N_3256);
or U3745 (N_3745,N_3363,N_3224);
or U3746 (N_3746,N_3088,N_3421);
and U3747 (N_3747,N_3048,N_3326);
nand U3748 (N_3748,N_3426,N_3159);
xor U3749 (N_3749,N_3258,N_3211);
and U3750 (N_3750,N_3442,N_3191);
nand U3751 (N_3751,N_3384,N_3209);
and U3752 (N_3752,N_3385,N_3384);
nor U3753 (N_3753,N_3459,N_3486);
and U3754 (N_3754,N_3498,N_3497);
nor U3755 (N_3755,N_3128,N_3364);
and U3756 (N_3756,N_3279,N_3312);
and U3757 (N_3757,N_3289,N_3304);
or U3758 (N_3758,N_3004,N_3365);
or U3759 (N_3759,N_3204,N_3190);
or U3760 (N_3760,N_3089,N_3277);
or U3761 (N_3761,N_3094,N_3225);
and U3762 (N_3762,N_3178,N_3044);
nor U3763 (N_3763,N_3355,N_3484);
or U3764 (N_3764,N_3301,N_3441);
and U3765 (N_3765,N_3155,N_3446);
xnor U3766 (N_3766,N_3203,N_3161);
or U3767 (N_3767,N_3301,N_3016);
and U3768 (N_3768,N_3311,N_3046);
or U3769 (N_3769,N_3220,N_3366);
or U3770 (N_3770,N_3223,N_3458);
nand U3771 (N_3771,N_3341,N_3377);
nand U3772 (N_3772,N_3131,N_3479);
nand U3773 (N_3773,N_3024,N_3080);
nor U3774 (N_3774,N_3219,N_3424);
nor U3775 (N_3775,N_3333,N_3072);
and U3776 (N_3776,N_3286,N_3351);
nor U3777 (N_3777,N_3225,N_3053);
nor U3778 (N_3778,N_3117,N_3418);
and U3779 (N_3779,N_3285,N_3056);
and U3780 (N_3780,N_3222,N_3133);
nand U3781 (N_3781,N_3191,N_3159);
nand U3782 (N_3782,N_3188,N_3247);
nand U3783 (N_3783,N_3336,N_3200);
nand U3784 (N_3784,N_3422,N_3405);
or U3785 (N_3785,N_3278,N_3148);
nand U3786 (N_3786,N_3289,N_3421);
nand U3787 (N_3787,N_3407,N_3239);
nand U3788 (N_3788,N_3167,N_3035);
nand U3789 (N_3789,N_3461,N_3310);
nor U3790 (N_3790,N_3144,N_3343);
and U3791 (N_3791,N_3031,N_3353);
or U3792 (N_3792,N_3220,N_3001);
or U3793 (N_3793,N_3162,N_3046);
xnor U3794 (N_3794,N_3277,N_3280);
or U3795 (N_3795,N_3154,N_3234);
or U3796 (N_3796,N_3274,N_3298);
or U3797 (N_3797,N_3438,N_3404);
or U3798 (N_3798,N_3366,N_3212);
xor U3799 (N_3799,N_3130,N_3145);
nand U3800 (N_3800,N_3355,N_3442);
nand U3801 (N_3801,N_3219,N_3233);
or U3802 (N_3802,N_3384,N_3085);
nor U3803 (N_3803,N_3146,N_3014);
nor U3804 (N_3804,N_3147,N_3412);
nor U3805 (N_3805,N_3429,N_3308);
and U3806 (N_3806,N_3065,N_3422);
and U3807 (N_3807,N_3321,N_3394);
nand U3808 (N_3808,N_3097,N_3016);
nor U3809 (N_3809,N_3360,N_3413);
and U3810 (N_3810,N_3350,N_3157);
nand U3811 (N_3811,N_3497,N_3231);
nand U3812 (N_3812,N_3250,N_3085);
or U3813 (N_3813,N_3307,N_3038);
nor U3814 (N_3814,N_3414,N_3187);
and U3815 (N_3815,N_3073,N_3206);
xnor U3816 (N_3816,N_3290,N_3162);
and U3817 (N_3817,N_3422,N_3135);
xor U3818 (N_3818,N_3388,N_3167);
xor U3819 (N_3819,N_3424,N_3047);
or U3820 (N_3820,N_3074,N_3372);
nand U3821 (N_3821,N_3036,N_3133);
or U3822 (N_3822,N_3469,N_3221);
or U3823 (N_3823,N_3174,N_3134);
nor U3824 (N_3824,N_3167,N_3257);
nor U3825 (N_3825,N_3214,N_3377);
nand U3826 (N_3826,N_3154,N_3243);
and U3827 (N_3827,N_3246,N_3256);
nand U3828 (N_3828,N_3077,N_3068);
nor U3829 (N_3829,N_3438,N_3071);
and U3830 (N_3830,N_3196,N_3209);
nand U3831 (N_3831,N_3099,N_3245);
nand U3832 (N_3832,N_3463,N_3036);
nand U3833 (N_3833,N_3165,N_3166);
nand U3834 (N_3834,N_3237,N_3425);
and U3835 (N_3835,N_3303,N_3060);
nand U3836 (N_3836,N_3373,N_3333);
nand U3837 (N_3837,N_3136,N_3414);
and U3838 (N_3838,N_3336,N_3050);
nand U3839 (N_3839,N_3231,N_3002);
nand U3840 (N_3840,N_3440,N_3389);
nand U3841 (N_3841,N_3443,N_3308);
or U3842 (N_3842,N_3236,N_3387);
nand U3843 (N_3843,N_3300,N_3090);
nand U3844 (N_3844,N_3095,N_3325);
and U3845 (N_3845,N_3200,N_3155);
or U3846 (N_3846,N_3331,N_3132);
xor U3847 (N_3847,N_3244,N_3265);
and U3848 (N_3848,N_3449,N_3096);
nor U3849 (N_3849,N_3297,N_3446);
xnor U3850 (N_3850,N_3457,N_3142);
or U3851 (N_3851,N_3300,N_3091);
nor U3852 (N_3852,N_3114,N_3433);
nand U3853 (N_3853,N_3301,N_3300);
nor U3854 (N_3854,N_3202,N_3497);
nand U3855 (N_3855,N_3243,N_3198);
or U3856 (N_3856,N_3467,N_3209);
or U3857 (N_3857,N_3401,N_3037);
or U3858 (N_3858,N_3190,N_3324);
and U3859 (N_3859,N_3104,N_3475);
and U3860 (N_3860,N_3451,N_3267);
and U3861 (N_3861,N_3001,N_3247);
xnor U3862 (N_3862,N_3233,N_3099);
nor U3863 (N_3863,N_3118,N_3172);
nand U3864 (N_3864,N_3219,N_3378);
nand U3865 (N_3865,N_3171,N_3384);
nand U3866 (N_3866,N_3330,N_3363);
nor U3867 (N_3867,N_3284,N_3073);
nand U3868 (N_3868,N_3460,N_3216);
and U3869 (N_3869,N_3261,N_3297);
and U3870 (N_3870,N_3327,N_3363);
nor U3871 (N_3871,N_3056,N_3297);
or U3872 (N_3872,N_3454,N_3355);
and U3873 (N_3873,N_3147,N_3249);
or U3874 (N_3874,N_3408,N_3248);
or U3875 (N_3875,N_3290,N_3377);
nand U3876 (N_3876,N_3345,N_3438);
and U3877 (N_3877,N_3249,N_3421);
nand U3878 (N_3878,N_3476,N_3102);
nand U3879 (N_3879,N_3315,N_3433);
nand U3880 (N_3880,N_3176,N_3150);
or U3881 (N_3881,N_3480,N_3116);
or U3882 (N_3882,N_3145,N_3267);
and U3883 (N_3883,N_3101,N_3036);
nand U3884 (N_3884,N_3068,N_3102);
nor U3885 (N_3885,N_3453,N_3060);
and U3886 (N_3886,N_3062,N_3379);
and U3887 (N_3887,N_3107,N_3138);
or U3888 (N_3888,N_3066,N_3398);
xnor U3889 (N_3889,N_3107,N_3361);
nor U3890 (N_3890,N_3424,N_3289);
and U3891 (N_3891,N_3048,N_3246);
or U3892 (N_3892,N_3059,N_3072);
and U3893 (N_3893,N_3089,N_3218);
nand U3894 (N_3894,N_3374,N_3330);
nor U3895 (N_3895,N_3036,N_3002);
nor U3896 (N_3896,N_3185,N_3397);
or U3897 (N_3897,N_3456,N_3158);
xnor U3898 (N_3898,N_3005,N_3298);
nor U3899 (N_3899,N_3464,N_3102);
nand U3900 (N_3900,N_3355,N_3381);
nand U3901 (N_3901,N_3053,N_3327);
or U3902 (N_3902,N_3034,N_3172);
and U3903 (N_3903,N_3163,N_3346);
nor U3904 (N_3904,N_3077,N_3309);
or U3905 (N_3905,N_3047,N_3456);
nand U3906 (N_3906,N_3429,N_3464);
or U3907 (N_3907,N_3140,N_3115);
nor U3908 (N_3908,N_3091,N_3299);
nand U3909 (N_3909,N_3055,N_3461);
and U3910 (N_3910,N_3156,N_3265);
nand U3911 (N_3911,N_3426,N_3409);
or U3912 (N_3912,N_3477,N_3347);
nand U3913 (N_3913,N_3240,N_3327);
or U3914 (N_3914,N_3492,N_3447);
or U3915 (N_3915,N_3441,N_3406);
or U3916 (N_3916,N_3214,N_3313);
and U3917 (N_3917,N_3113,N_3280);
and U3918 (N_3918,N_3338,N_3296);
nand U3919 (N_3919,N_3059,N_3210);
and U3920 (N_3920,N_3084,N_3060);
or U3921 (N_3921,N_3160,N_3104);
nand U3922 (N_3922,N_3175,N_3004);
and U3923 (N_3923,N_3266,N_3451);
nor U3924 (N_3924,N_3490,N_3193);
or U3925 (N_3925,N_3332,N_3471);
nor U3926 (N_3926,N_3104,N_3476);
nor U3927 (N_3927,N_3438,N_3414);
or U3928 (N_3928,N_3091,N_3376);
xnor U3929 (N_3929,N_3451,N_3177);
nor U3930 (N_3930,N_3017,N_3466);
or U3931 (N_3931,N_3156,N_3433);
nand U3932 (N_3932,N_3078,N_3396);
or U3933 (N_3933,N_3499,N_3347);
and U3934 (N_3934,N_3361,N_3362);
nand U3935 (N_3935,N_3311,N_3225);
and U3936 (N_3936,N_3081,N_3252);
and U3937 (N_3937,N_3008,N_3339);
nor U3938 (N_3938,N_3154,N_3366);
or U3939 (N_3939,N_3087,N_3323);
nand U3940 (N_3940,N_3305,N_3199);
nand U3941 (N_3941,N_3437,N_3064);
nand U3942 (N_3942,N_3114,N_3412);
nor U3943 (N_3943,N_3115,N_3408);
nand U3944 (N_3944,N_3437,N_3177);
or U3945 (N_3945,N_3186,N_3284);
and U3946 (N_3946,N_3302,N_3274);
and U3947 (N_3947,N_3444,N_3332);
or U3948 (N_3948,N_3428,N_3053);
and U3949 (N_3949,N_3488,N_3447);
nand U3950 (N_3950,N_3065,N_3354);
nor U3951 (N_3951,N_3044,N_3154);
xnor U3952 (N_3952,N_3230,N_3127);
nor U3953 (N_3953,N_3308,N_3034);
nand U3954 (N_3954,N_3073,N_3021);
and U3955 (N_3955,N_3110,N_3164);
or U3956 (N_3956,N_3133,N_3196);
and U3957 (N_3957,N_3049,N_3246);
and U3958 (N_3958,N_3261,N_3247);
nand U3959 (N_3959,N_3289,N_3122);
nor U3960 (N_3960,N_3112,N_3351);
nor U3961 (N_3961,N_3206,N_3422);
or U3962 (N_3962,N_3428,N_3476);
nor U3963 (N_3963,N_3365,N_3146);
or U3964 (N_3964,N_3221,N_3040);
and U3965 (N_3965,N_3262,N_3484);
and U3966 (N_3966,N_3318,N_3099);
or U3967 (N_3967,N_3439,N_3462);
nor U3968 (N_3968,N_3033,N_3438);
nand U3969 (N_3969,N_3396,N_3226);
xnor U3970 (N_3970,N_3012,N_3448);
xnor U3971 (N_3971,N_3409,N_3301);
nor U3972 (N_3972,N_3119,N_3205);
nand U3973 (N_3973,N_3158,N_3203);
or U3974 (N_3974,N_3263,N_3307);
nor U3975 (N_3975,N_3207,N_3276);
or U3976 (N_3976,N_3300,N_3203);
nand U3977 (N_3977,N_3248,N_3031);
nand U3978 (N_3978,N_3051,N_3193);
or U3979 (N_3979,N_3399,N_3063);
and U3980 (N_3980,N_3045,N_3370);
or U3981 (N_3981,N_3366,N_3493);
and U3982 (N_3982,N_3211,N_3012);
and U3983 (N_3983,N_3327,N_3347);
nor U3984 (N_3984,N_3329,N_3146);
and U3985 (N_3985,N_3308,N_3255);
nand U3986 (N_3986,N_3008,N_3161);
or U3987 (N_3987,N_3402,N_3354);
nand U3988 (N_3988,N_3105,N_3238);
or U3989 (N_3989,N_3039,N_3384);
nand U3990 (N_3990,N_3105,N_3227);
nor U3991 (N_3991,N_3415,N_3394);
and U3992 (N_3992,N_3372,N_3301);
nand U3993 (N_3993,N_3035,N_3231);
xor U3994 (N_3994,N_3385,N_3391);
nand U3995 (N_3995,N_3258,N_3194);
and U3996 (N_3996,N_3379,N_3432);
and U3997 (N_3997,N_3492,N_3029);
nor U3998 (N_3998,N_3038,N_3409);
nor U3999 (N_3999,N_3314,N_3260);
xor U4000 (N_4000,N_3563,N_3514);
and U4001 (N_4001,N_3924,N_3680);
nand U4002 (N_4002,N_3763,N_3685);
or U4003 (N_4003,N_3715,N_3671);
or U4004 (N_4004,N_3885,N_3678);
nand U4005 (N_4005,N_3717,N_3899);
or U4006 (N_4006,N_3747,N_3825);
or U4007 (N_4007,N_3775,N_3777);
nand U4008 (N_4008,N_3767,N_3960);
xnor U4009 (N_4009,N_3890,N_3756);
and U4010 (N_4010,N_3925,N_3605);
xor U4011 (N_4011,N_3785,N_3849);
nand U4012 (N_4012,N_3795,N_3809);
nor U4013 (N_4013,N_3604,N_3638);
or U4014 (N_4014,N_3762,N_3842);
or U4015 (N_4015,N_3700,N_3574);
nand U4016 (N_4016,N_3559,N_3919);
nor U4017 (N_4017,N_3728,N_3512);
nor U4018 (N_4018,N_3992,N_3718);
or U4019 (N_4019,N_3807,N_3534);
nand U4020 (N_4020,N_3936,N_3820);
nor U4021 (N_4021,N_3852,N_3853);
nor U4022 (N_4022,N_3546,N_3702);
xor U4023 (N_4023,N_3502,N_3964);
or U4024 (N_4024,N_3692,N_3623);
nand U4025 (N_4025,N_3694,N_3547);
and U4026 (N_4026,N_3591,N_3965);
xnor U4027 (N_4027,N_3505,N_3761);
or U4028 (N_4028,N_3799,N_3889);
xor U4029 (N_4029,N_3632,N_3804);
nor U4030 (N_4030,N_3812,N_3773);
nand U4031 (N_4031,N_3877,N_3548);
and U4032 (N_4032,N_3658,N_3770);
nand U4033 (N_4033,N_3985,N_3878);
xnor U4034 (N_4034,N_3577,N_3752);
nand U4035 (N_4035,N_3682,N_3601);
or U4036 (N_4036,N_3729,N_3945);
nand U4037 (N_4037,N_3616,N_3518);
and U4038 (N_4038,N_3581,N_3724);
or U4039 (N_4039,N_3740,N_3647);
nand U4040 (N_4040,N_3793,N_3954);
and U4041 (N_4041,N_3712,N_3674);
and U4042 (N_4042,N_3713,N_3948);
and U4043 (N_4043,N_3920,N_3608);
xor U4044 (N_4044,N_3926,N_3526);
nor U4045 (N_4045,N_3957,N_3677);
or U4046 (N_4046,N_3845,N_3725);
and U4047 (N_4047,N_3843,N_3710);
nor U4048 (N_4048,N_3558,N_3633);
nor U4049 (N_4049,N_3681,N_3754);
and U4050 (N_4050,N_3759,N_3753);
and U4051 (N_4051,N_3722,N_3566);
and U4052 (N_4052,N_3634,N_3881);
nand U4053 (N_4053,N_3982,N_3832);
and U4054 (N_4054,N_3603,N_3611);
xor U4055 (N_4055,N_3579,N_3980);
nand U4056 (N_4056,N_3739,N_3606);
nand U4057 (N_4057,N_3507,N_3934);
nand U4058 (N_4058,N_3977,N_3552);
and U4059 (N_4059,N_3983,N_3774);
or U4060 (N_4060,N_3944,N_3930);
nand U4061 (N_4061,N_3991,N_3911);
nor U4062 (N_4062,N_3769,N_3586);
or U4063 (N_4063,N_3629,N_3743);
nor U4064 (N_4064,N_3979,N_3808);
nor U4065 (N_4065,N_3646,N_3539);
nor U4066 (N_4066,N_3643,N_3856);
xor U4067 (N_4067,N_3598,N_3939);
and U4068 (N_4068,N_3587,N_3828);
nand U4069 (N_4069,N_3789,N_3571);
and U4070 (N_4070,N_3510,N_3532);
and U4071 (N_4071,N_3779,N_3971);
and U4072 (N_4072,N_3588,N_3984);
or U4073 (N_4073,N_3529,N_3708);
and U4074 (N_4074,N_3848,N_3719);
nor U4075 (N_4075,N_3766,N_3609);
nor U4076 (N_4076,N_3704,N_3916);
nand U4077 (N_4077,N_3988,N_3522);
nand U4078 (N_4078,N_3689,N_3501);
or U4079 (N_4079,N_3962,N_3963);
and U4080 (N_4080,N_3855,N_3593);
nand U4081 (N_4081,N_3627,N_3676);
nor U4082 (N_4082,N_3750,N_3691);
or U4083 (N_4083,N_3995,N_3701);
nor U4084 (N_4084,N_3851,N_3662);
and U4085 (N_4085,N_3876,N_3741);
nor U4086 (N_4086,N_3821,N_3661);
and U4087 (N_4087,N_3537,N_3891);
and U4088 (N_4088,N_3838,N_3663);
and U4089 (N_4089,N_3705,N_3645);
xnor U4090 (N_4090,N_3764,N_3961);
and U4091 (N_4091,N_3847,N_3573);
and U4092 (N_4092,N_3626,N_3567);
and U4093 (N_4093,N_3986,N_3687);
or U4094 (N_4094,N_3817,N_3822);
or U4095 (N_4095,N_3542,N_3723);
and U4096 (N_4096,N_3721,N_3543);
nand U4097 (N_4097,N_3953,N_3690);
xor U4098 (N_4098,N_3837,N_3525);
nand U4099 (N_4099,N_3778,N_3896);
xor U4100 (N_4100,N_3797,N_3655);
nand U4101 (N_4101,N_3600,N_3931);
nand U4102 (N_4102,N_3918,N_3839);
and U4103 (N_4103,N_3892,N_3744);
or U4104 (N_4104,N_3557,N_3993);
nor U4105 (N_4105,N_3783,N_3511);
nand U4106 (N_4106,N_3928,N_3862);
or U4107 (N_4107,N_3956,N_3697);
or U4108 (N_4108,N_3967,N_3905);
and U4109 (N_4109,N_3875,N_3897);
nor U4110 (N_4110,N_3914,N_3709);
nand U4111 (N_4111,N_3612,N_3902);
xnor U4112 (N_4112,N_3660,N_3698);
nand U4113 (N_4113,N_3699,N_3947);
xor U4114 (N_4114,N_3519,N_3751);
or U4115 (N_4115,N_3528,N_3866);
nor U4116 (N_4116,N_3688,N_3933);
nor U4117 (N_4117,N_3520,N_3664);
nand U4118 (N_4118,N_3870,N_3578);
or U4119 (N_4119,N_3997,N_3978);
nor U4120 (N_4120,N_3815,N_3857);
and U4121 (N_4121,N_3669,N_3927);
or U4122 (N_4122,N_3871,N_3811);
or U4123 (N_4123,N_3639,N_3860);
nand U4124 (N_4124,N_3665,N_3824);
and U4125 (N_4125,N_3565,N_3900);
and U4126 (N_4126,N_3550,N_3635);
nor U4127 (N_4127,N_3707,N_3553);
nand U4128 (N_4128,N_3938,N_3906);
and U4129 (N_4129,N_3720,N_3736);
or U4130 (N_4130,N_3966,N_3716);
nand U4131 (N_4131,N_3907,N_3904);
or U4132 (N_4132,N_3508,N_3735);
nor U4133 (N_4133,N_3940,N_3792);
nor U4134 (N_4134,N_3749,N_3950);
or U4135 (N_4135,N_3631,N_3536);
nor U4136 (N_4136,N_3901,N_3730);
and U4137 (N_4137,N_3524,N_3912);
nor U4138 (N_4138,N_3556,N_3610);
and U4139 (N_4139,N_3874,N_3863);
nand U4140 (N_4140,N_3684,N_3737);
nand U4141 (N_4141,N_3540,N_3806);
and U4142 (N_4142,N_3583,N_3672);
or U4143 (N_4143,N_3607,N_3513);
nand U4144 (N_4144,N_3597,N_3921);
and U4145 (N_4145,N_3580,N_3541);
and U4146 (N_4146,N_3654,N_3826);
or U4147 (N_4147,N_3903,N_3562);
or U4148 (N_4148,N_3516,N_3859);
nor U4149 (N_4149,N_3544,N_3584);
or U4150 (N_4150,N_3673,N_3883);
xnor U4151 (N_4151,N_3554,N_3816);
nand U4152 (N_4152,N_3706,N_3831);
or U4153 (N_4153,N_3958,N_3595);
nand U4154 (N_4154,N_3670,N_3503);
nor U4155 (N_4155,N_3652,N_3895);
or U4156 (N_4156,N_3570,N_3500);
and U4157 (N_4157,N_3854,N_3893);
and U4158 (N_4158,N_3757,N_3840);
or U4159 (N_4159,N_3803,N_3738);
nand U4160 (N_4160,N_3576,N_3810);
nor U4161 (N_4161,N_3768,N_3675);
nor U4162 (N_4162,N_3693,N_3802);
xnor U4163 (N_4163,N_3861,N_3630);
nand U4164 (N_4164,N_3935,N_3733);
and U4165 (N_4165,N_3833,N_3836);
and U4166 (N_4166,N_3758,N_3805);
xnor U4167 (N_4167,N_3644,N_3794);
xnor U4168 (N_4168,N_3755,N_3873);
and U4169 (N_4169,N_3641,N_3521);
nor U4170 (N_4170,N_3745,N_3780);
nor U4171 (N_4171,N_3594,N_3614);
and U4172 (N_4172,N_3527,N_3765);
or U4173 (N_4173,N_3642,N_3679);
nor U4174 (N_4174,N_3879,N_3929);
or U4175 (N_4175,N_3998,N_3615);
xor U4176 (N_4176,N_3656,N_3585);
nand U4177 (N_4177,N_3987,N_3649);
nor U4178 (N_4178,N_3898,N_3549);
or U4179 (N_4179,N_3731,N_3561);
nand U4180 (N_4180,N_3636,N_3533);
nor U4181 (N_4181,N_3772,N_3592);
and U4182 (N_4182,N_3886,N_3640);
nand U4183 (N_4183,N_3932,N_3538);
nand U4184 (N_4184,N_3796,N_3726);
nand U4185 (N_4185,N_3732,N_3653);
nor U4186 (N_4186,N_3894,N_3968);
and U4187 (N_4187,N_3887,N_3504);
or U4188 (N_4188,N_3959,N_3545);
or U4189 (N_4189,N_3798,N_3990);
or U4190 (N_4190,N_3996,N_3790);
and U4191 (N_4191,N_3989,N_3711);
and U4192 (N_4192,N_3823,N_3517);
and U4193 (N_4193,N_3589,N_3923);
or U4194 (N_4194,N_3868,N_3830);
or U4195 (N_4195,N_3858,N_3835);
or U4196 (N_4196,N_3872,N_3869);
and U4197 (N_4197,N_3949,N_3791);
nor U4198 (N_4198,N_3976,N_3974);
or U4199 (N_4199,N_3523,N_3551);
nor U4200 (N_4200,N_3703,N_3575);
nor U4201 (N_4201,N_3952,N_3613);
and U4202 (N_4202,N_3695,N_3867);
and U4203 (N_4203,N_3813,N_3908);
xor U4204 (N_4204,N_3746,N_3865);
or U4205 (N_4205,N_3624,N_3909);
nor U4206 (N_4206,N_3955,N_3776);
or U4207 (N_4207,N_3727,N_3827);
nand U4208 (N_4208,N_3617,N_3981);
or U4209 (N_4209,N_3683,N_3941);
nor U4210 (N_4210,N_3942,N_3973);
nand U4211 (N_4211,N_3560,N_3910);
and U4212 (N_4212,N_3782,N_3922);
and U4213 (N_4213,N_3625,N_3696);
or U4214 (N_4214,N_3844,N_3734);
nand U4215 (N_4215,N_3506,N_3651);
or U4216 (N_4216,N_3568,N_3535);
nor U4217 (N_4217,N_3572,N_3596);
or U4218 (N_4218,N_3637,N_3619);
nand U4219 (N_4219,N_3888,N_3994);
or U4220 (N_4220,N_3951,N_3800);
nand U4221 (N_4221,N_3969,N_3667);
nor U4222 (N_4222,N_3801,N_3784);
nor U4223 (N_4223,N_3846,N_3882);
or U4224 (N_4224,N_3668,N_3850);
and U4225 (N_4225,N_3564,N_3618);
xor U4226 (N_4226,N_3781,N_3582);
nand U4227 (N_4227,N_3714,N_3531);
nor U4228 (N_4228,N_3913,N_3818);
and U4229 (N_4229,N_3917,N_3760);
nor U4230 (N_4230,N_3569,N_3834);
nand U4231 (N_4231,N_3841,N_3972);
and U4232 (N_4232,N_3999,N_3686);
or U4233 (N_4233,N_3659,N_3590);
nand U4234 (N_4234,N_3943,N_3829);
and U4235 (N_4235,N_3628,N_3884);
nand U4236 (N_4236,N_3814,N_3648);
nor U4237 (N_4237,N_3937,N_3975);
or U4238 (N_4238,N_3748,N_3788);
nor U4239 (N_4239,N_3946,N_3666);
nor U4240 (N_4240,N_3970,N_3622);
or U4241 (N_4241,N_3819,N_3742);
and U4242 (N_4242,N_3771,N_3530);
nand U4243 (N_4243,N_3509,N_3787);
or U4244 (N_4244,N_3620,N_3621);
nor U4245 (N_4245,N_3657,N_3786);
xor U4246 (N_4246,N_3864,N_3515);
nand U4247 (N_4247,N_3915,N_3599);
or U4248 (N_4248,N_3602,N_3880);
nor U4249 (N_4249,N_3555,N_3650);
and U4250 (N_4250,N_3767,N_3805);
or U4251 (N_4251,N_3880,N_3879);
nor U4252 (N_4252,N_3650,N_3538);
and U4253 (N_4253,N_3901,N_3804);
nor U4254 (N_4254,N_3911,N_3539);
nor U4255 (N_4255,N_3586,N_3980);
and U4256 (N_4256,N_3864,N_3519);
nor U4257 (N_4257,N_3849,N_3740);
and U4258 (N_4258,N_3887,N_3920);
or U4259 (N_4259,N_3688,N_3655);
nand U4260 (N_4260,N_3771,N_3850);
or U4261 (N_4261,N_3827,N_3622);
and U4262 (N_4262,N_3770,N_3943);
or U4263 (N_4263,N_3580,N_3866);
and U4264 (N_4264,N_3746,N_3806);
nor U4265 (N_4265,N_3885,N_3522);
and U4266 (N_4266,N_3956,N_3983);
nand U4267 (N_4267,N_3706,N_3878);
or U4268 (N_4268,N_3530,N_3916);
nand U4269 (N_4269,N_3823,N_3952);
nor U4270 (N_4270,N_3841,N_3686);
nand U4271 (N_4271,N_3519,N_3599);
nor U4272 (N_4272,N_3786,N_3779);
and U4273 (N_4273,N_3571,N_3527);
nor U4274 (N_4274,N_3631,N_3525);
xnor U4275 (N_4275,N_3741,N_3845);
or U4276 (N_4276,N_3619,N_3635);
nor U4277 (N_4277,N_3690,N_3774);
and U4278 (N_4278,N_3824,N_3992);
and U4279 (N_4279,N_3840,N_3692);
nor U4280 (N_4280,N_3760,N_3939);
nand U4281 (N_4281,N_3516,N_3741);
nor U4282 (N_4282,N_3806,N_3838);
nand U4283 (N_4283,N_3862,N_3916);
and U4284 (N_4284,N_3755,N_3914);
or U4285 (N_4285,N_3982,N_3753);
and U4286 (N_4286,N_3863,N_3521);
and U4287 (N_4287,N_3725,N_3928);
or U4288 (N_4288,N_3712,N_3904);
nand U4289 (N_4289,N_3725,N_3590);
xor U4290 (N_4290,N_3742,N_3932);
nand U4291 (N_4291,N_3633,N_3635);
nor U4292 (N_4292,N_3697,N_3993);
and U4293 (N_4293,N_3926,N_3596);
nand U4294 (N_4294,N_3891,N_3880);
and U4295 (N_4295,N_3976,N_3623);
or U4296 (N_4296,N_3902,N_3503);
or U4297 (N_4297,N_3604,N_3520);
nor U4298 (N_4298,N_3609,N_3778);
and U4299 (N_4299,N_3647,N_3910);
xor U4300 (N_4300,N_3715,N_3965);
xor U4301 (N_4301,N_3666,N_3739);
and U4302 (N_4302,N_3812,N_3948);
or U4303 (N_4303,N_3832,N_3754);
nor U4304 (N_4304,N_3866,N_3925);
and U4305 (N_4305,N_3764,N_3980);
nand U4306 (N_4306,N_3527,N_3749);
nand U4307 (N_4307,N_3730,N_3591);
nor U4308 (N_4308,N_3978,N_3775);
or U4309 (N_4309,N_3598,N_3549);
or U4310 (N_4310,N_3998,N_3879);
or U4311 (N_4311,N_3506,N_3737);
and U4312 (N_4312,N_3950,N_3918);
nor U4313 (N_4313,N_3838,N_3724);
and U4314 (N_4314,N_3510,N_3639);
nor U4315 (N_4315,N_3970,N_3703);
and U4316 (N_4316,N_3560,N_3770);
or U4317 (N_4317,N_3878,N_3828);
or U4318 (N_4318,N_3580,N_3783);
nor U4319 (N_4319,N_3963,N_3650);
nand U4320 (N_4320,N_3539,N_3552);
nand U4321 (N_4321,N_3535,N_3810);
and U4322 (N_4322,N_3676,N_3842);
or U4323 (N_4323,N_3976,N_3579);
or U4324 (N_4324,N_3864,N_3606);
or U4325 (N_4325,N_3555,N_3599);
and U4326 (N_4326,N_3569,N_3884);
or U4327 (N_4327,N_3970,N_3840);
nand U4328 (N_4328,N_3984,N_3791);
or U4329 (N_4329,N_3831,N_3804);
and U4330 (N_4330,N_3990,N_3855);
and U4331 (N_4331,N_3828,N_3803);
nand U4332 (N_4332,N_3936,N_3878);
nor U4333 (N_4333,N_3933,N_3986);
or U4334 (N_4334,N_3870,N_3666);
xor U4335 (N_4335,N_3500,N_3956);
nand U4336 (N_4336,N_3764,N_3602);
nand U4337 (N_4337,N_3519,N_3945);
or U4338 (N_4338,N_3938,N_3915);
nand U4339 (N_4339,N_3921,N_3839);
nand U4340 (N_4340,N_3878,N_3669);
nor U4341 (N_4341,N_3739,N_3825);
or U4342 (N_4342,N_3554,N_3613);
and U4343 (N_4343,N_3793,N_3914);
and U4344 (N_4344,N_3503,N_3993);
nor U4345 (N_4345,N_3555,N_3568);
nand U4346 (N_4346,N_3627,N_3747);
and U4347 (N_4347,N_3530,N_3703);
nor U4348 (N_4348,N_3511,N_3651);
and U4349 (N_4349,N_3991,N_3790);
nor U4350 (N_4350,N_3978,N_3711);
and U4351 (N_4351,N_3921,N_3739);
xnor U4352 (N_4352,N_3797,N_3815);
nor U4353 (N_4353,N_3794,N_3609);
xor U4354 (N_4354,N_3517,N_3636);
and U4355 (N_4355,N_3865,N_3778);
or U4356 (N_4356,N_3727,N_3771);
nand U4357 (N_4357,N_3789,N_3733);
nand U4358 (N_4358,N_3924,N_3774);
and U4359 (N_4359,N_3630,N_3930);
and U4360 (N_4360,N_3786,N_3809);
nand U4361 (N_4361,N_3730,N_3767);
xor U4362 (N_4362,N_3538,N_3919);
and U4363 (N_4363,N_3658,N_3640);
and U4364 (N_4364,N_3597,N_3905);
or U4365 (N_4365,N_3867,N_3580);
and U4366 (N_4366,N_3803,N_3629);
or U4367 (N_4367,N_3827,N_3581);
nor U4368 (N_4368,N_3573,N_3882);
nand U4369 (N_4369,N_3710,N_3606);
nand U4370 (N_4370,N_3587,N_3885);
nand U4371 (N_4371,N_3910,N_3887);
or U4372 (N_4372,N_3689,N_3734);
nor U4373 (N_4373,N_3673,N_3745);
xor U4374 (N_4374,N_3863,N_3570);
nand U4375 (N_4375,N_3798,N_3677);
nand U4376 (N_4376,N_3560,N_3956);
and U4377 (N_4377,N_3999,N_3766);
nor U4378 (N_4378,N_3568,N_3706);
nand U4379 (N_4379,N_3917,N_3685);
nand U4380 (N_4380,N_3979,N_3586);
nor U4381 (N_4381,N_3933,N_3784);
nand U4382 (N_4382,N_3578,N_3826);
and U4383 (N_4383,N_3878,N_3680);
or U4384 (N_4384,N_3714,N_3762);
nand U4385 (N_4385,N_3598,N_3596);
or U4386 (N_4386,N_3686,N_3970);
nand U4387 (N_4387,N_3524,N_3726);
nor U4388 (N_4388,N_3881,N_3536);
and U4389 (N_4389,N_3500,N_3778);
and U4390 (N_4390,N_3902,N_3896);
or U4391 (N_4391,N_3873,N_3716);
and U4392 (N_4392,N_3707,N_3585);
and U4393 (N_4393,N_3636,N_3757);
nor U4394 (N_4394,N_3607,N_3661);
or U4395 (N_4395,N_3873,N_3546);
xor U4396 (N_4396,N_3875,N_3886);
or U4397 (N_4397,N_3562,N_3663);
and U4398 (N_4398,N_3875,N_3672);
nor U4399 (N_4399,N_3903,N_3515);
or U4400 (N_4400,N_3926,N_3834);
nand U4401 (N_4401,N_3786,N_3511);
nand U4402 (N_4402,N_3658,N_3627);
nand U4403 (N_4403,N_3714,N_3627);
nor U4404 (N_4404,N_3994,N_3739);
nand U4405 (N_4405,N_3772,N_3658);
nor U4406 (N_4406,N_3556,N_3810);
and U4407 (N_4407,N_3850,N_3955);
xnor U4408 (N_4408,N_3520,N_3878);
xnor U4409 (N_4409,N_3825,N_3674);
nand U4410 (N_4410,N_3640,N_3615);
nor U4411 (N_4411,N_3508,N_3651);
nor U4412 (N_4412,N_3636,N_3993);
xnor U4413 (N_4413,N_3824,N_3853);
and U4414 (N_4414,N_3539,N_3864);
nor U4415 (N_4415,N_3908,N_3530);
and U4416 (N_4416,N_3717,N_3790);
nor U4417 (N_4417,N_3707,N_3895);
or U4418 (N_4418,N_3814,N_3913);
nor U4419 (N_4419,N_3550,N_3627);
or U4420 (N_4420,N_3620,N_3897);
nor U4421 (N_4421,N_3644,N_3867);
nor U4422 (N_4422,N_3512,N_3649);
or U4423 (N_4423,N_3893,N_3523);
or U4424 (N_4424,N_3836,N_3766);
nor U4425 (N_4425,N_3662,N_3519);
and U4426 (N_4426,N_3688,N_3710);
nand U4427 (N_4427,N_3576,N_3964);
xor U4428 (N_4428,N_3501,N_3515);
nor U4429 (N_4429,N_3851,N_3519);
and U4430 (N_4430,N_3741,N_3622);
nand U4431 (N_4431,N_3944,N_3551);
nor U4432 (N_4432,N_3981,N_3836);
xnor U4433 (N_4433,N_3961,N_3874);
xnor U4434 (N_4434,N_3868,N_3846);
nor U4435 (N_4435,N_3841,N_3931);
nand U4436 (N_4436,N_3508,N_3967);
nand U4437 (N_4437,N_3788,N_3571);
nor U4438 (N_4438,N_3918,N_3929);
nor U4439 (N_4439,N_3982,N_3510);
nand U4440 (N_4440,N_3668,N_3892);
and U4441 (N_4441,N_3608,N_3988);
and U4442 (N_4442,N_3952,N_3921);
or U4443 (N_4443,N_3918,N_3697);
and U4444 (N_4444,N_3914,N_3839);
and U4445 (N_4445,N_3507,N_3514);
nand U4446 (N_4446,N_3564,N_3902);
or U4447 (N_4447,N_3770,N_3510);
nand U4448 (N_4448,N_3846,N_3709);
nand U4449 (N_4449,N_3844,N_3789);
or U4450 (N_4450,N_3907,N_3845);
nor U4451 (N_4451,N_3549,N_3968);
or U4452 (N_4452,N_3903,N_3723);
nor U4453 (N_4453,N_3501,N_3574);
and U4454 (N_4454,N_3570,N_3854);
nor U4455 (N_4455,N_3667,N_3975);
nand U4456 (N_4456,N_3757,N_3910);
nor U4457 (N_4457,N_3607,N_3861);
or U4458 (N_4458,N_3579,N_3869);
nand U4459 (N_4459,N_3900,N_3861);
nor U4460 (N_4460,N_3762,N_3961);
and U4461 (N_4461,N_3894,N_3519);
nor U4462 (N_4462,N_3935,N_3538);
nor U4463 (N_4463,N_3533,N_3821);
nand U4464 (N_4464,N_3786,N_3971);
and U4465 (N_4465,N_3985,N_3716);
or U4466 (N_4466,N_3652,N_3616);
or U4467 (N_4467,N_3586,N_3660);
nor U4468 (N_4468,N_3741,N_3695);
nand U4469 (N_4469,N_3713,N_3823);
and U4470 (N_4470,N_3669,N_3505);
nand U4471 (N_4471,N_3643,N_3935);
and U4472 (N_4472,N_3660,N_3780);
nand U4473 (N_4473,N_3964,N_3520);
nand U4474 (N_4474,N_3778,N_3855);
or U4475 (N_4475,N_3736,N_3975);
xnor U4476 (N_4476,N_3711,N_3811);
or U4477 (N_4477,N_3660,N_3817);
nor U4478 (N_4478,N_3697,N_3611);
nand U4479 (N_4479,N_3665,N_3887);
and U4480 (N_4480,N_3831,N_3705);
and U4481 (N_4481,N_3515,N_3589);
and U4482 (N_4482,N_3750,N_3792);
and U4483 (N_4483,N_3799,N_3894);
or U4484 (N_4484,N_3983,N_3787);
nand U4485 (N_4485,N_3673,N_3570);
or U4486 (N_4486,N_3500,N_3616);
nor U4487 (N_4487,N_3589,N_3982);
and U4488 (N_4488,N_3592,N_3853);
or U4489 (N_4489,N_3811,N_3889);
and U4490 (N_4490,N_3773,N_3680);
and U4491 (N_4491,N_3676,N_3788);
or U4492 (N_4492,N_3755,N_3758);
nand U4493 (N_4493,N_3992,N_3810);
xor U4494 (N_4494,N_3919,N_3673);
and U4495 (N_4495,N_3877,N_3857);
xor U4496 (N_4496,N_3943,N_3962);
or U4497 (N_4497,N_3693,N_3644);
nor U4498 (N_4498,N_3579,N_3792);
nor U4499 (N_4499,N_3819,N_3820);
nand U4500 (N_4500,N_4044,N_4251);
nor U4501 (N_4501,N_4213,N_4479);
nand U4502 (N_4502,N_4421,N_4088);
and U4503 (N_4503,N_4344,N_4194);
nor U4504 (N_4504,N_4151,N_4257);
nor U4505 (N_4505,N_4392,N_4411);
nor U4506 (N_4506,N_4167,N_4428);
nand U4507 (N_4507,N_4143,N_4082);
and U4508 (N_4508,N_4066,N_4242);
and U4509 (N_4509,N_4214,N_4229);
nor U4510 (N_4510,N_4102,N_4371);
nor U4511 (N_4511,N_4061,N_4309);
nor U4512 (N_4512,N_4494,N_4005);
nor U4513 (N_4513,N_4131,N_4000);
nor U4514 (N_4514,N_4169,N_4389);
xor U4515 (N_4515,N_4203,N_4150);
xor U4516 (N_4516,N_4087,N_4207);
and U4517 (N_4517,N_4328,N_4261);
nor U4518 (N_4518,N_4413,N_4313);
or U4519 (N_4519,N_4170,N_4033);
nand U4520 (N_4520,N_4191,N_4105);
nand U4521 (N_4521,N_4282,N_4224);
nor U4522 (N_4522,N_4304,N_4056);
nand U4523 (N_4523,N_4443,N_4117);
xor U4524 (N_4524,N_4473,N_4090);
or U4525 (N_4525,N_4454,N_4084);
and U4526 (N_4526,N_4283,N_4023);
or U4527 (N_4527,N_4260,N_4077);
and U4528 (N_4528,N_4373,N_4230);
and U4529 (N_4529,N_4244,N_4085);
or U4530 (N_4530,N_4036,N_4069);
or U4531 (N_4531,N_4152,N_4431);
or U4532 (N_4532,N_4012,N_4320);
nor U4533 (N_4533,N_4490,N_4447);
nor U4534 (N_4534,N_4441,N_4157);
nor U4535 (N_4535,N_4175,N_4202);
and U4536 (N_4536,N_4333,N_4146);
and U4537 (N_4537,N_4404,N_4334);
or U4538 (N_4538,N_4367,N_4019);
nor U4539 (N_4539,N_4226,N_4124);
and U4540 (N_4540,N_4034,N_4198);
nor U4541 (N_4541,N_4126,N_4350);
nor U4542 (N_4542,N_4075,N_4480);
nor U4543 (N_4543,N_4292,N_4439);
and U4544 (N_4544,N_4254,N_4264);
nand U4545 (N_4545,N_4402,N_4250);
nor U4546 (N_4546,N_4427,N_4255);
and U4547 (N_4547,N_4380,N_4384);
and U4548 (N_4548,N_4408,N_4100);
nand U4549 (N_4549,N_4498,N_4217);
nand U4550 (N_4550,N_4448,N_4122);
nand U4551 (N_4551,N_4187,N_4184);
or U4552 (N_4552,N_4183,N_4489);
and U4553 (N_4553,N_4359,N_4234);
nor U4554 (N_4554,N_4495,N_4430);
nand U4555 (N_4555,N_4185,N_4091);
nand U4556 (N_4556,N_4163,N_4368);
nor U4557 (N_4557,N_4468,N_4327);
and U4558 (N_4558,N_4189,N_4071);
and U4559 (N_4559,N_4115,N_4286);
nand U4560 (N_4560,N_4054,N_4032);
nand U4561 (N_4561,N_4065,N_4285);
nand U4562 (N_4562,N_4485,N_4280);
nand U4563 (N_4563,N_4021,N_4345);
and U4564 (N_4564,N_4058,N_4356);
nand U4565 (N_4565,N_4478,N_4422);
and U4566 (N_4566,N_4195,N_4365);
nor U4567 (N_4567,N_4295,N_4111);
nor U4568 (N_4568,N_4471,N_4357);
or U4569 (N_4569,N_4456,N_4381);
xor U4570 (N_4570,N_4237,N_4376);
and U4571 (N_4571,N_4140,N_4205);
xor U4572 (N_4572,N_4458,N_4319);
xnor U4573 (N_4573,N_4051,N_4089);
nor U4574 (N_4574,N_4247,N_4128);
nor U4575 (N_4575,N_4211,N_4160);
or U4576 (N_4576,N_4096,N_4063);
nor U4577 (N_4577,N_4385,N_4343);
nand U4578 (N_4578,N_4403,N_4026);
nand U4579 (N_4579,N_4446,N_4050);
nor U4580 (N_4580,N_4390,N_4437);
nor U4581 (N_4581,N_4174,N_4486);
xnor U4582 (N_4582,N_4400,N_4452);
or U4583 (N_4583,N_4149,N_4388);
and U4584 (N_4584,N_4168,N_4340);
and U4585 (N_4585,N_4308,N_4068);
nor U4586 (N_4586,N_4018,N_4451);
nor U4587 (N_4587,N_4287,N_4147);
or U4588 (N_4588,N_4316,N_4406);
or U4589 (N_4589,N_4414,N_4161);
nand U4590 (N_4590,N_4272,N_4003);
nand U4591 (N_4591,N_4281,N_4290);
nor U4592 (N_4592,N_4249,N_4154);
or U4593 (N_4593,N_4335,N_4104);
xnor U4594 (N_4594,N_4293,N_4132);
and U4595 (N_4595,N_4225,N_4097);
nor U4596 (N_4596,N_4006,N_4259);
xor U4597 (N_4597,N_4302,N_4366);
nor U4598 (N_4598,N_4346,N_4410);
or U4599 (N_4599,N_4420,N_4166);
xnor U4600 (N_4600,N_4190,N_4135);
or U4601 (N_4601,N_4138,N_4412);
nand U4602 (N_4602,N_4031,N_4011);
and U4603 (N_4603,N_4049,N_4072);
nor U4604 (N_4604,N_4052,N_4156);
nor U4605 (N_4605,N_4432,N_4141);
nor U4606 (N_4606,N_4222,N_4435);
or U4607 (N_4607,N_4337,N_4236);
or U4608 (N_4608,N_4442,N_4294);
nand U4609 (N_4609,N_4227,N_4445);
nor U4610 (N_4610,N_4277,N_4349);
nor U4611 (N_4611,N_4246,N_4475);
nor U4612 (N_4612,N_4112,N_4415);
nand U4613 (N_4613,N_4288,N_4312);
and U4614 (N_4614,N_4323,N_4332);
and U4615 (N_4615,N_4114,N_4383);
nor U4616 (N_4616,N_4035,N_4098);
nor U4617 (N_4617,N_4109,N_4177);
and U4618 (N_4618,N_4076,N_4080);
nand U4619 (N_4619,N_4296,N_4326);
or U4620 (N_4620,N_4101,N_4047);
or U4621 (N_4621,N_4284,N_4476);
or U4622 (N_4622,N_4401,N_4238);
nor U4623 (N_4623,N_4208,N_4059);
or U4624 (N_4624,N_4039,N_4375);
nor U4625 (N_4625,N_4306,N_4178);
or U4626 (N_4626,N_4221,N_4144);
or U4627 (N_4627,N_4358,N_4165);
nor U4628 (N_4628,N_4014,N_4378);
or U4629 (N_4629,N_4298,N_4215);
xor U4630 (N_4630,N_4074,N_4391);
nand U4631 (N_4631,N_4318,N_4179);
xor U4632 (N_4632,N_4274,N_4017);
or U4633 (N_4633,N_4418,N_4387);
nand U4634 (N_4634,N_4395,N_4266);
xor U4635 (N_4635,N_4271,N_4482);
nor U4636 (N_4636,N_4464,N_4315);
nand U4637 (N_4637,N_4118,N_4002);
nand U4638 (N_4638,N_4010,N_4279);
nand U4639 (N_4639,N_4305,N_4363);
and U4640 (N_4640,N_4062,N_4046);
and U4641 (N_4641,N_4436,N_4453);
and U4642 (N_4642,N_4278,N_4275);
xor U4643 (N_4643,N_4331,N_4407);
nor U4644 (N_4644,N_4450,N_4182);
or U4645 (N_4645,N_4459,N_4022);
or U4646 (N_4646,N_4488,N_4201);
nand U4647 (N_4647,N_4057,N_4270);
and U4648 (N_4648,N_4369,N_4186);
xor U4649 (N_4649,N_4125,N_4139);
nor U4650 (N_4650,N_4491,N_4078);
xnor U4651 (N_4651,N_4417,N_4322);
nor U4652 (N_4652,N_4461,N_4496);
nor U4653 (N_4653,N_4291,N_4336);
nor U4654 (N_4654,N_4253,N_4273);
or U4655 (N_4655,N_4197,N_4110);
nand U4656 (N_4656,N_4301,N_4093);
or U4657 (N_4657,N_4241,N_4045);
nor U4658 (N_4658,N_4130,N_4119);
xnor U4659 (N_4659,N_4300,N_4196);
nor U4660 (N_4660,N_4398,N_4347);
and U4661 (N_4661,N_4396,N_4268);
or U4662 (N_4662,N_4425,N_4438);
xor U4663 (N_4663,N_4397,N_4027);
or U4664 (N_4664,N_4338,N_4219);
nor U4665 (N_4665,N_4386,N_4463);
or U4666 (N_4666,N_4469,N_4209);
or U4667 (N_4667,N_4181,N_4370);
or U4668 (N_4668,N_4434,N_4307);
and U4669 (N_4669,N_4024,N_4136);
xor U4670 (N_4670,N_4393,N_4107);
and U4671 (N_4671,N_4472,N_4269);
nor U4672 (N_4672,N_4258,N_4419);
nand U4673 (N_4673,N_4341,N_4121);
nand U4674 (N_4674,N_4297,N_4113);
or U4675 (N_4675,N_4133,N_4030);
and U4676 (N_4676,N_4095,N_4233);
or U4677 (N_4677,N_4487,N_4013);
nor U4678 (N_4678,N_4499,N_4362);
or U4679 (N_4679,N_4015,N_4199);
xnor U4680 (N_4680,N_4232,N_4262);
and U4681 (N_4681,N_4204,N_4467);
nor U4682 (N_4682,N_4008,N_4321);
or U4683 (N_4683,N_4172,N_4210);
nand U4684 (N_4684,N_4470,N_4155);
nor U4685 (N_4685,N_4108,N_4355);
nor U4686 (N_4686,N_4220,N_4239);
and U4687 (N_4687,N_4218,N_4330);
nor U4688 (N_4688,N_4252,N_4192);
nand U4689 (N_4689,N_4342,N_4460);
and U4690 (N_4690,N_4497,N_4153);
xor U4691 (N_4691,N_4164,N_4399);
and U4692 (N_4692,N_4481,N_4354);
nand U4693 (N_4693,N_4042,N_4007);
nand U4694 (N_4694,N_4416,N_4099);
or U4695 (N_4695,N_4311,N_4142);
nor U4696 (N_4696,N_4041,N_4405);
or U4697 (N_4697,N_4120,N_4372);
and U4698 (N_4698,N_4070,N_4200);
or U4699 (N_4699,N_4248,N_4484);
xor U4700 (N_4700,N_4364,N_4351);
nor U4701 (N_4701,N_4081,N_4038);
nor U4702 (N_4702,N_4424,N_4231);
nand U4703 (N_4703,N_4440,N_4043);
and U4704 (N_4704,N_4073,N_4483);
xor U4705 (N_4705,N_4106,N_4352);
nand U4706 (N_4706,N_4103,N_4206);
or U4707 (N_4707,N_4116,N_4009);
or U4708 (N_4708,N_4243,N_4016);
and U4709 (N_4709,N_4159,N_4462);
and U4710 (N_4710,N_4409,N_4423);
nor U4711 (N_4711,N_4092,N_4276);
xor U4712 (N_4712,N_4158,N_4265);
nand U4713 (N_4713,N_4004,N_4348);
or U4714 (N_4714,N_4444,N_4145);
or U4715 (N_4715,N_4317,N_4429);
nand U4716 (N_4716,N_4067,N_4374);
or U4717 (N_4717,N_4377,N_4457);
nor U4718 (N_4718,N_4245,N_4493);
nor U4719 (N_4719,N_4465,N_4064);
xnor U4720 (N_4720,N_4382,N_4129);
or U4721 (N_4721,N_4361,N_4324);
and U4722 (N_4722,N_4123,N_4001);
nand U4723 (N_4723,N_4433,N_4171);
nor U4724 (N_4724,N_4310,N_4134);
nand U4725 (N_4725,N_4455,N_4256);
nor U4726 (N_4726,N_4477,N_4360);
nor U4727 (N_4727,N_4314,N_4162);
xnor U4728 (N_4728,N_4148,N_4267);
xnor U4729 (N_4729,N_4223,N_4060);
nand U4730 (N_4730,N_4492,N_4176);
nor U4731 (N_4731,N_4028,N_4094);
xnor U4732 (N_4732,N_4289,N_4086);
or U4733 (N_4733,N_4083,N_4137);
nor U4734 (N_4734,N_4353,N_4193);
xnor U4735 (N_4735,N_4474,N_4426);
nor U4736 (N_4736,N_4029,N_4299);
nand U4737 (N_4737,N_4037,N_4263);
or U4738 (N_4738,N_4180,N_4020);
and U4739 (N_4739,N_4325,N_4339);
nand U4740 (N_4740,N_4055,N_4212);
and U4741 (N_4741,N_4329,N_4449);
and U4742 (N_4742,N_4040,N_4228);
nand U4743 (N_4743,N_4079,N_4235);
nor U4744 (N_4744,N_4025,N_4303);
or U4745 (N_4745,N_4053,N_4394);
or U4746 (N_4746,N_4188,N_4466);
nor U4747 (N_4747,N_4127,N_4173);
or U4748 (N_4748,N_4216,N_4379);
nand U4749 (N_4749,N_4240,N_4048);
nor U4750 (N_4750,N_4232,N_4464);
nand U4751 (N_4751,N_4166,N_4025);
and U4752 (N_4752,N_4109,N_4046);
xnor U4753 (N_4753,N_4053,N_4184);
and U4754 (N_4754,N_4163,N_4006);
xnor U4755 (N_4755,N_4101,N_4286);
nor U4756 (N_4756,N_4286,N_4090);
and U4757 (N_4757,N_4207,N_4447);
xnor U4758 (N_4758,N_4431,N_4273);
xnor U4759 (N_4759,N_4006,N_4076);
or U4760 (N_4760,N_4270,N_4373);
nor U4761 (N_4761,N_4372,N_4337);
xor U4762 (N_4762,N_4250,N_4210);
xnor U4763 (N_4763,N_4381,N_4101);
nor U4764 (N_4764,N_4095,N_4353);
and U4765 (N_4765,N_4315,N_4124);
and U4766 (N_4766,N_4298,N_4404);
nand U4767 (N_4767,N_4069,N_4492);
nand U4768 (N_4768,N_4363,N_4055);
and U4769 (N_4769,N_4252,N_4214);
nor U4770 (N_4770,N_4328,N_4159);
nand U4771 (N_4771,N_4420,N_4036);
or U4772 (N_4772,N_4208,N_4147);
nor U4773 (N_4773,N_4068,N_4184);
nand U4774 (N_4774,N_4106,N_4475);
nor U4775 (N_4775,N_4427,N_4404);
or U4776 (N_4776,N_4144,N_4228);
nor U4777 (N_4777,N_4276,N_4061);
nor U4778 (N_4778,N_4332,N_4334);
and U4779 (N_4779,N_4368,N_4421);
and U4780 (N_4780,N_4047,N_4133);
and U4781 (N_4781,N_4049,N_4260);
or U4782 (N_4782,N_4308,N_4219);
and U4783 (N_4783,N_4159,N_4489);
xnor U4784 (N_4784,N_4037,N_4098);
nor U4785 (N_4785,N_4036,N_4243);
or U4786 (N_4786,N_4356,N_4495);
nand U4787 (N_4787,N_4018,N_4363);
nor U4788 (N_4788,N_4337,N_4106);
and U4789 (N_4789,N_4213,N_4255);
or U4790 (N_4790,N_4006,N_4269);
or U4791 (N_4791,N_4035,N_4202);
or U4792 (N_4792,N_4173,N_4063);
nand U4793 (N_4793,N_4323,N_4384);
or U4794 (N_4794,N_4015,N_4428);
nand U4795 (N_4795,N_4118,N_4163);
or U4796 (N_4796,N_4215,N_4314);
xor U4797 (N_4797,N_4158,N_4063);
or U4798 (N_4798,N_4143,N_4019);
xnor U4799 (N_4799,N_4315,N_4042);
or U4800 (N_4800,N_4039,N_4386);
or U4801 (N_4801,N_4413,N_4433);
and U4802 (N_4802,N_4489,N_4418);
nor U4803 (N_4803,N_4127,N_4070);
or U4804 (N_4804,N_4476,N_4187);
or U4805 (N_4805,N_4051,N_4024);
xor U4806 (N_4806,N_4439,N_4483);
nor U4807 (N_4807,N_4180,N_4417);
nor U4808 (N_4808,N_4181,N_4188);
and U4809 (N_4809,N_4058,N_4103);
and U4810 (N_4810,N_4061,N_4443);
nand U4811 (N_4811,N_4403,N_4475);
or U4812 (N_4812,N_4219,N_4103);
and U4813 (N_4813,N_4177,N_4358);
or U4814 (N_4814,N_4274,N_4128);
nor U4815 (N_4815,N_4256,N_4100);
and U4816 (N_4816,N_4182,N_4178);
nor U4817 (N_4817,N_4467,N_4141);
xnor U4818 (N_4818,N_4243,N_4488);
and U4819 (N_4819,N_4007,N_4420);
and U4820 (N_4820,N_4470,N_4365);
nor U4821 (N_4821,N_4219,N_4463);
nor U4822 (N_4822,N_4110,N_4303);
nand U4823 (N_4823,N_4447,N_4046);
xnor U4824 (N_4824,N_4253,N_4320);
nand U4825 (N_4825,N_4300,N_4310);
nand U4826 (N_4826,N_4165,N_4026);
nor U4827 (N_4827,N_4332,N_4301);
and U4828 (N_4828,N_4345,N_4221);
nand U4829 (N_4829,N_4246,N_4339);
xor U4830 (N_4830,N_4337,N_4047);
nand U4831 (N_4831,N_4165,N_4196);
or U4832 (N_4832,N_4448,N_4135);
and U4833 (N_4833,N_4452,N_4182);
nand U4834 (N_4834,N_4231,N_4372);
nand U4835 (N_4835,N_4022,N_4144);
nand U4836 (N_4836,N_4127,N_4454);
nor U4837 (N_4837,N_4037,N_4017);
nand U4838 (N_4838,N_4080,N_4465);
nand U4839 (N_4839,N_4205,N_4141);
nand U4840 (N_4840,N_4247,N_4359);
or U4841 (N_4841,N_4204,N_4075);
xnor U4842 (N_4842,N_4324,N_4489);
or U4843 (N_4843,N_4154,N_4356);
nor U4844 (N_4844,N_4144,N_4130);
nand U4845 (N_4845,N_4126,N_4304);
and U4846 (N_4846,N_4227,N_4393);
and U4847 (N_4847,N_4261,N_4281);
nand U4848 (N_4848,N_4220,N_4106);
nor U4849 (N_4849,N_4408,N_4136);
and U4850 (N_4850,N_4427,N_4274);
or U4851 (N_4851,N_4108,N_4228);
or U4852 (N_4852,N_4387,N_4360);
or U4853 (N_4853,N_4457,N_4126);
or U4854 (N_4854,N_4287,N_4316);
or U4855 (N_4855,N_4143,N_4123);
or U4856 (N_4856,N_4284,N_4358);
xnor U4857 (N_4857,N_4166,N_4335);
nand U4858 (N_4858,N_4077,N_4469);
and U4859 (N_4859,N_4193,N_4268);
nand U4860 (N_4860,N_4334,N_4257);
nor U4861 (N_4861,N_4131,N_4005);
nor U4862 (N_4862,N_4366,N_4498);
nor U4863 (N_4863,N_4470,N_4120);
nor U4864 (N_4864,N_4212,N_4173);
nand U4865 (N_4865,N_4334,N_4316);
and U4866 (N_4866,N_4193,N_4279);
nor U4867 (N_4867,N_4073,N_4315);
and U4868 (N_4868,N_4173,N_4076);
xnor U4869 (N_4869,N_4261,N_4235);
xnor U4870 (N_4870,N_4072,N_4336);
nand U4871 (N_4871,N_4371,N_4463);
nor U4872 (N_4872,N_4392,N_4170);
nor U4873 (N_4873,N_4278,N_4417);
nand U4874 (N_4874,N_4289,N_4297);
and U4875 (N_4875,N_4302,N_4089);
nor U4876 (N_4876,N_4003,N_4456);
or U4877 (N_4877,N_4411,N_4235);
or U4878 (N_4878,N_4144,N_4124);
nor U4879 (N_4879,N_4138,N_4233);
nor U4880 (N_4880,N_4104,N_4353);
or U4881 (N_4881,N_4065,N_4284);
and U4882 (N_4882,N_4284,N_4016);
xnor U4883 (N_4883,N_4493,N_4058);
and U4884 (N_4884,N_4338,N_4122);
nor U4885 (N_4885,N_4010,N_4225);
nand U4886 (N_4886,N_4041,N_4196);
and U4887 (N_4887,N_4150,N_4089);
and U4888 (N_4888,N_4257,N_4290);
xnor U4889 (N_4889,N_4050,N_4402);
and U4890 (N_4890,N_4177,N_4168);
and U4891 (N_4891,N_4243,N_4026);
nor U4892 (N_4892,N_4491,N_4320);
and U4893 (N_4893,N_4431,N_4101);
nand U4894 (N_4894,N_4431,N_4095);
or U4895 (N_4895,N_4339,N_4322);
or U4896 (N_4896,N_4236,N_4005);
and U4897 (N_4897,N_4266,N_4131);
nand U4898 (N_4898,N_4169,N_4049);
nand U4899 (N_4899,N_4269,N_4023);
nand U4900 (N_4900,N_4056,N_4177);
nand U4901 (N_4901,N_4283,N_4453);
nand U4902 (N_4902,N_4354,N_4447);
and U4903 (N_4903,N_4361,N_4074);
xor U4904 (N_4904,N_4261,N_4238);
or U4905 (N_4905,N_4279,N_4482);
nor U4906 (N_4906,N_4185,N_4410);
or U4907 (N_4907,N_4409,N_4252);
and U4908 (N_4908,N_4479,N_4103);
and U4909 (N_4909,N_4159,N_4318);
nor U4910 (N_4910,N_4426,N_4065);
and U4911 (N_4911,N_4332,N_4119);
or U4912 (N_4912,N_4118,N_4154);
or U4913 (N_4913,N_4419,N_4330);
nand U4914 (N_4914,N_4137,N_4134);
or U4915 (N_4915,N_4041,N_4085);
xnor U4916 (N_4916,N_4325,N_4332);
nand U4917 (N_4917,N_4351,N_4097);
nand U4918 (N_4918,N_4339,N_4259);
and U4919 (N_4919,N_4406,N_4483);
nor U4920 (N_4920,N_4322,N_4418);
and U4921 (N_4921,N_4170,N_4215);
and U4922 (N_4922,N_4365,N_4332);
and U4923 (N_4923,N_4245,N_4239);
nand U4924 (N_4924,N_4380,N_4226);
nand U4925 (N_4925,N_4173,N_4100);
nor U4926 (N_4926,N_4445,N_4039);
nor U4927 (N_4927,N_4079,N_4092);
or U4928 (N_4928,N_4091,N_4381);
xnor U4929 (N_4929,N_4442,N_4026);
and U4930 (N_4930,N_4072,N_4230);
xor U4931 (N_4931,N_4225,N_4440);
nand U4932 (N_4932,N_4025,N_4111);
or U4933 (N_4933,N_4455,N_4233);
nor U4934 (N_4934,N_4167,N_4300);
nor U4935 (N_4935,N_4056,N_4320);
nand U4936 (N_4936,N_4082,N_4256);
and U4937 (N_4937,N_4483,N_4222);
or U4938 (N_4938,N_4197,N_4215);
nand U4939 (N_4939,N_4004,N_4118);
or U4940 (N_4940,N_4336,N_4487);
nand U4941 (N_4941,N_4238,N_4045);
and U4942 (N_4942,N_4093,N_4044);
nand U4943 (N_4943,N_4237,N_4294);
or U4944 (N_4944,N_4287,N_4193);
or U4945 (N_4945,N_4372,N_4433);
xor U4946 (N_4946,N_4449,N_4321);
nor U4947 (N_4947,N_4381,N_4494);
or U4948 (N_4948,N_4215,N_4030);
nand U4949 (N_4949,N_4234,N_4278);
xnor U4950 (N_4950,N_4489,N_4042);
or U4951 (N_4951,N_4454,N_4074);
nor U4952 (N_4952,N_4053,N_4420);
nor U4953 (N_4953,N_4150,N_4016);
and U4954 (N_4954,N_4284,N_4139);
nand U4955 (N_4955,N_4023,N_4429);
xnor U4956 (N_4956,N_4132,N_4235);
and U4957 (N_4957,N_4459,N_4410);
or U4958 (N_4958,N_4268,N_4252);
xor U4959 (N_4959,N_4426,N_4107);
nand U4960 (N_4960,N_4188,N_4320);
or U4961 (N_4961,N_4332,N_4007);
nand U4962 (N_4962,N_4029,N_4119);
and U4963 (N_4963,N_4145,N_4188);
nand U4964 (N_4964,N_4393,N_4334);
and U4965 (N_4965,N_4066,N_4096);
nor U4966 (N_4966,N_4165,N_4258);
and U4967 (N_4967,N_4419,N_4479);
and U4968 (N_4968,N_4016,N_4050);
and U4969 (N_4969,N_4049,N_4251);
or U4970 (N_4970,N_4203,N_4456);
nor U4971 (N_4971,N_4166,N_4478);
nand U4972 (N_4972,N_4055,N_4204);
or U4973 (N_4973,N_4404,N_4403);
nand U4974 (N_4974,N_4405,N_4020);
and U4975 (N_4975,N_4222,N_4430);
nor U4976 (N_4976,N_4227,N_4264);
nor U4977 (N_4977,N_4238,N_4481);
nor U4978 (N_4978,N_4119,N_4112);
nand U4979 (N_4979,N_4431,N_4170);
nor U4980 (N_4980,N_4486,N_4482);
nand U4981 (N_4981,N_4133,N_4098);
and U4982 (N_4982,N_4073,N_4130);
or U4983 (N_4983,N_4499,N_4085);
and U4984 (N_4984,N_4047,N_4258);
and U4985 (N_4985,N_4046,N_4213);
and U4986 (N_4986,N_4457,N_4244);
and U4987 (N_4987,N_4051,N_4455);
and U4988 (N_4988,N_4090,N_4298);
nand U4989 (N_4989,N_4063,N_4455);
xnor U4990 (N_4990,N_4110,N_4247);
nor U4991 (N_4991,N_4163,N_4224);
nand U4992 (N_4992,N_4218,N_4353);
nand U4993 (N_4993,N_4492,N_4146);
and U4994 (N_4994,N_4347,N_4251);
nand U4995 (N_4995,N_4447,N_4229);
or U4996 (N_4996,N_4431,N_4357);
nor U4997 (N_4997,N_4201,N_4417);
nor U4998 (N_4998,N_4442,N_4049);
or U4999 (N_4999,N_4226,N_4197);
and U5000 (N_5000,N_4726,N_4903);
or U5001 (N_5001,N_4699,N_4925);
xor U5002 (N_5002,N_4666,N_4999);
and U5003 (N_5003,N_4577,N_4952);
xor U5004 (N_5004,N_4688,N_4943);
and U5005 (N_5005,N_4752,N_4632);
and U5006 (N_5006,N_4692,N_4774);
and U5007 (N_5007,N_4982,N_4503);
and U5008 (N_5008,N_4888,N_4549);
and U5009 (N_5009,N_4911,N_4875);
nor U5010 (N_5010,N_4877,N_4797);
and U5011 (N_5011,N_4651,N_4816);
nand U5012 (N_5012,N_4654,N_4957);
and U5013 (N_5013,N_4758,N_4893);
nor U5014 (N_5014,N_4514,N_4822);
nor U5015 (N_5015,N_4723,N_4621);
or U5016 (N_5016,N_4779,N_4522);
nand U5017 (N_5017,N_4773,N_4769);
and U5018 (N_5018,N_4656,N_4808);
xor U5019 (N_5019,N_4901,N_4806);
nor U5020 (N_5020,N_4883,N_4551);
nor U5021 (N_5021,N_4868,N_4947);
or U5022 (N_5022,N_4720,N_4960);
xnor U5023 (N_5023,N_4658,N_4622);
or U5024 (N_5024,N_4838,N_4961);
nor U5025 (N_5025,N_4655,N_4834);
nand U5026 (N_5026,N_4873,N_4556);
nor U5027 (N_5027,N_4983,N_4645);
nor U5028 (N_5028,N_4524,N_4867);
and U5029 (N_5029,N_4639,N_4755);
nand U5030 (N_5030,N_4970,N_4855);
and U5031 (N_5031,N_4602,N_4581);
and U5032 (N_5032,N_4563,N_4809);
or U5033 (N_5033,N_4765,N_4798);
or U5034 (N_5034,N_4704,N_4660);
and U5035 (N_5035,N_4818,N_4972);
nor U5036 (N_5036,N_4749,N_4861);
nor U5037 (N_5037,N_4730,N_4531);
and U5038 (N_5038,N_4793,N_4969);
or U5039 (N_5039,N_4968,N_4512);
or U5040 (N_5040,N_4625,N_4821);
or U5041 (N_5041,N_4711,N_4828);
nor U5042 (N_5042,N_4706,N_4600);
nor U5043 (N_5043,N_4853,N_4684);
xor U5044 (N_5044,N_4908,N_4876);
nor U5045 (N_5045,N_4772,N_4523);
or U5046 (N_5046,N_4535,N_4530);
xnor U5047 (N_5047,N_4582,N_4592);
nor U5048 (N_5048,N_4913,N_4744);
xor U5049 (N_5049,N_4653,N_4646);
or U5050 (N_5050,N_4605,N_4724);
and U5051 (N_5051,N_4912,N_4844);
nor U5052 (N_5052,N_4784,N_4538);
nand U5053 (N_5053,N_4945,N_4790);
nand U5054 (N_5054,N_4880,N_4845);
nand U5055 (N_5055,N_4751,N_4517);
nand U5056 (N_5056,N_4548,N_4515);
nor U5057 (N_5057,N_4626,N_4896);
xor U5058 (N_5058,N_4899,N_4792);
or U5059 (N_5059,N_4678,N_4995);
nand U5060 (N_5060,N_4843,N_4799);
and U5061 (N_5061,N_4963,N_4664);
nand U5062 (N_5062,N_4553,N_4987);
or U5063 (N_5063,N_4629,N_4951);
nor U5064 (N_5064,N_4782,N_4606);
and U5065 (N_5065,N_4544,N_4839);
and U5066 (N_5066,N_4895,N_4785);
nor U5067 (N_5067,N_4764,N_4540);
and U5068 (N_5068,N_4985,N_4910);
and U5069 (N_5069,N_4944,N_4650);
nand U5070 (N_5070,N_4736,N_4932);
or U5071 (N_5071,N_4815,N_4928);
xnor U5072 (N_5072,N_4949,N_4946);
or U5073 (N_5073,N_4796,N_4775);
and U5074 (N_5074,N_4921,N_4783);
xnor U5075 (N_5075,N_4975,N_4683);
and U5076 (N_5076,N_4713,N_4611);
nand U5077 (N_5077,N_4886,N_4804);
or U5078 (N_5078,N_4670,N_4830);
nor U5079 (N_5079,N_4864,N_4667);
nand U5080 (N_5080,N_4718,N_4641);
and U5081 (N_5081,N_4558,N_4703);
nor U5082 (N_5082,N_4506,N_4746);
nor U5083 (N_5083,N_4638,N_4948);
nor U5084 (N_5084,N_4608,N_4962);
nand U5085 (N_5085,N_4511,N_4978);
nand U5086 (N_5086,N_4636,N_4616);
nor U5087 (N_5087,N_4572,N_4679);
nor U5088 (N_5088,N_4567,N_4827);
nand U5089 (N_5089,N_4587,N_4627);
nand U5090 (N_5090,N_4504,N_4731);
and U5091 (N_5091,N_4974,N_4643);
nand U5092 (N_5092,N_4560,N_4574);
and U5093 (N_5093,N_4984,N_4719);
nor U5094 (N_5094,N_4689,N_4942);
and U5095 (N_5095,N_4545,N_4835);
nor U5096 (N_5096,N_4994,N_4846);
or U5097 (N_5097,N_4937,N_4938);
nand U5098 (N_5098,N_4905,N_4698);
or U5099 (N_5099,N_4585,N_4732);
xor U5100 (N_5100,N_4833,N_4979);
nor U5101 (N_5101,N_4635,N_4857);
xor U5102 (N_5102,N_4906,N_4525);
nand U5103 (N_5103,N_4794,N_4955);
nor U5104 (N_5104,N_4940,N_4771);
and U5105 (N_5105,N_4580,N_4509);
or U5106 (N_5106,N_4820,N_4856);
or U5107 (N_5107,N_4966,N_4568);
nand U5108 (N_5108,N_4673,N_4885);
nand U5109 (N_5109,N_4738,N_4848);
nor U5110 (N_5110,N_4777,N_4686);
or U5111 (N_5111,N_4756,N_4507);
nor U5112 (N_5112,N_4647,N_4702);
xor U5113 (N_5113,N_4971,N_4836);
and U5114 (N_5114,N_4935,N_4807);
nand U5115 (N_5115,N_4789,N_4863);
or U5116 (N_5116,N_4989,N_4941);
and U5117 (N_5117,N_4882,N_4677);
and U5118 (N_5118,N_4735,N_4694);
or U5119 (N_5119,N_4527,N_4902);
nand U5120 (N_5120,N_4763,N_4924);
nand U5121 (N_5121,N_4598,N_4926);
nor U5122 (N_5122,N_4976,N_4562);
nor U5123 (N_5123,N_4541,N_4813);
nor U5124 (N_5124,N_4508,N_4700);
nand U5125 (N_5125,N_4564,N_4865);
nor U5126 (N_5126,N_4591,N_4780);
xor U5127 (N_5127,N_4762,N_4781);
nand U5128 (N_5128,N_4958,N_4993);
or U5129 (N_5129,N_4546,N_4858);
or U5130 (N_5130,N_4543,N_4739);
or U5131 (N_5131,N_4554,N_4701);
nand U5132 (N_5132,N_4922,N_4840);
nor U5133 (N_5133,N_4559,N_4871);
and U5134 (N_5134,N_4892,N_4528);
nor U5135 (N_5135,N_4570,N_4753);
or U5136 (N_5136,N_4741,N_4576);
and U5137 (N_5137,N_4613,N_4642);
nand U5138 (N_5138,N_4802,N_4934);
xnor U5139 (N_5139,N_4860,N_4954);
xor U5140 (N_5140,N_4917,N_4998);
or U5141 (N_5141,N_4967,N_4536);
nor U5142 (N_5142,N_4542,N_4696);
nor U5143 (N_5143,N_4770,N_4661);
and U5144 (N_5144,N_4620,N_4884);
nor U5145 (N_5145,N_4814,N_4918);
xnor U5146 (N_5146,N_4693,N_4850);
nor U5147 (N_5147,N_4748,N_4933);
nand U5148 (N_5148,N_4537,N_4500);
nand U5149 (N_5149,N_4676,N_4672);
nand U5150 (N_5150,N_4931,N_4936);
or U5151 (N_5151,N_4852,N_4788);
xor U5152 (N_5152,N_4566,N_4854);
and U5153 (N_5153,N_4817,N_4533);
nor U5154 (N_5154,N_4829,N_4659);
and U5155 (N_5155,N_4603,N_4668);
nand U5156 (N_5156,N_4502,N_4599);
and U5157 (N_5157,N_4849,N_4589);
or U5158 (N_5158,N_4891,N_4520);
nor U5159 (N_5159,N_4878,N_4980);
nor U5160 (N_5160,N_4619,N_4550);
xnor U5161 (N_5161,N_4609,N_4604);
and U5162 (N_5162,N_4707,N_4716);
nor U5163 (N_5163,N_4964,N_4521);
and U5164 (N_5164,N_4601,N_4709);
nand U5165 (N_5165,N_4721,N_4595);
and U5166 (N_5166,N_4526,N_4519);
nand U5167 (N_5167,N_4881,N_4761);
or U5168 (N_5168,N_4991,N_4607);
or U5169 (N_5169,N_4889,N_4759);
or U5170 (N_5170,N_4740,N_4927);
nand U5171 (N_5171,N_4869,N_4823);
or U5172 (N_5172,N_4743,N_4615);
nor U5173 (N_5173,N_4826,N_4505);
or U5174 (N_5174,N_4648,N_4710);
and U5175 (N_5175,N_4939,N_4593);
or U5176 (N_5176,N_4669,N_4675);
or U5177 (N_5177,N_4539,N_4652);
nand U5178 (N_5178,N_4733,N_4717);
or U5179 (N_5179,N_4695,N_4555);
and U5180 (N_5180,N_4786,N_4907);
nor U5181 (N_5181,N_4557,N_4584);
xor U5182 (N_5182,N_4930,N_4630);
or U5183 (N_5183,N_4801,N_4811);
nand U5184 (N_5184,N_4965,N_4841);
or U5185 (N_5185,N_4640,N_4671);
and U5186 (N_5186,N_4663,N_4859);
nand U5187 (N_5187,N_4518,N_4547);
and U5188 (N_5188,N_4617,N_4819);
nor U5189 (N_5189,N_4897,N_4708);
nor U5190 (N_5190,N_4631,N_4649);
nand U5191 (N_5191,N_4812,N_4697);
nor U5192 (N_5192,N_4552,N_4579);
and U5193 (N_5193,N_4915,N_4767);
nand U5194 (N_5194,N_4997,N_4776);
nor U5195 (N_5195,N_4990,N_4824);
nand U5196 (N_5196,N_4565,N_4742);
nand U5197 (N_5197,N_4729,N_4529);
or U5198 (N_5198,N_4728,N_4900);
nor U5199 (N_5199,N_4866,N_4919);
xor U5200 (N_5200,N_4727,N_4904);
xnor U5201 (N_5201,N_4862,N_4956);
xor U5202 (N_5202,N_4778,N_4583);
or U5203 (N_5203,N_4624,N_4768);
nand U5204 (N_5204,N_4610,N_4959);
xnor U5205 (N_5205,N_4837,N_4916);
and U5206 (N_5206,N_4725,N_4687);
or U5207 (N_5207,N_4832,N_4920);
nand U5208 (N_5208,N_4665,N_4992);
or U5209 (N_5209,N_4691,N_4872);
nor U5210 (N_5210,N_4623,N_4923);
nor U5211 (N_5211,N_4810,N_4996);
xnor U5212 (N_5212,N_4745,N_4657);
xnor U5213 (N_5213,N_4532,N_4825);
nand U5214 (N_5214,N_4685,N_4805);
nand U5215 (N_5215,N_4516,N_4569);
and U5216 (N_5216,N_4662,N_4597);
nand U5217 (N_5217,N_4561,N_4594);
or U5218 (N_5218,N_4890,N_4633);
or U5219 (N_5219,N_4747,N_4575);
nand U5220 (N_5220,N_4847,N_4754);
or U5221 (N_5221,N_4628,N_4682);
xor U5222 (N_5222,N_4977,N_4909);
nor U5223 (N_5223,N_4510,N_4705);
and U5224 (N_5224,N_4795,N_4898);
nand U5225 (N_5225,N_4590,N_4874);
xor U5226 (N_5226,N_4986,N_4870);
and U5227 (N_5227,N_4894,N_4787);
and U5228 (N_5228,N_4644,N_4586);
nor U5229 (N_5229,N_4588,N_4534);
or U5230 (N_5230,N_4737,N_4722);
nand U5231 (N_5231,N_4715,N_4750);
nand U5232 (N_5232,N_4851,N_4879);
nand U5233 (N_5233,N_4766,N_4634);
nor U5234 (N_5234,N_4573,N_4803);
nor U5235 (N_5235,N_4714,N_4578);
and U5236 (N_5236,N_4680,N_4571);
xor U5237 (N_5237,N_4760,N_4501);
nor U5238 (N_5238,N_4734,N_4988);
or U5239 (N_5239,N_4757,N_4618);
xnor U5240 (N_5240,N_4614,N_4831);
nor U5241 (N_5241,N_4791,N_4973);
or U5242 (N_5242,N_4596,N_4513);
nor U5243 (N_5243,N_4929,N_4681);
and U5244 (N_5244,N_4674,N_4981);
nor U5245 (N_5245,N_4637,N_4914);
nor U5246 (N_5246,N_4950,N_4712);
nand U5247 (N_5247,N_4612,N_4800);
nor U5248 (N_5248,N_4690,N_4842);
or U5249 (N_5249,N_4887,N_4953);
xnor U5250 (N_5250,N_4989,N_4713);
nor U5251 (N_5251,N_4771,N_4704);
xor U5252 (N_5252,N_4544,N_4677);
and U5253 (N_5253,N_4647,N_4664);
xor U5254 (N_5254,N_4654,N_4736);
and U5255 (N_5255,N_4574,N_4845);
or U5256 (N_5256,N_4996,N_4597);
nand U5257 (N_5257,N_4749,N_4881);
nor U5258 (N_5258,N_4623,N_4539);
or U5259 (N_5259,N_4547,N_4667);
and U5260 (N_5260,N_4831,N_4968);
or U5261 (N_5261,N_4798,N_4746);
or U5262 (N_5262,N_4941,N_4853);
nand U5263 (N_5263,N_4685,N_4950);
and U5264 (N_5264,N_4710,N_4785);
or U5265 (N_5265,N_4521,N_4523);
nand U5266 (N_5266,N_4989,N_4601);
nand U5267 (N_5267,N_4555,N_4921);
and U5268 (N_5268,N_4669,N_4802);
or U5269 (N_5269,N_4879,N_4955);
nand U5270 (N_5270,N_4935,N_4655);
or U5271 (N_5271,N_4694,N_4955);
nor U5272 (N_5272,N_4597,N_4651);
and U5273 (N_5273,N_4959,N_4858);
nand U5274 (N_5274,N_4900,N_4837);
nand U5275 (N_5275,N_4789,N_4966);
or U5276 (N_5276,N_4595,N_4901);
xnor U5277 (N_5277,N_4917,N_4827);
and U5278 (N_5278,N_4603,N_4747);
and U5279 (N_5279,N_4710,N_4864);
or U5280 (N_5280,N_4615,N_4696);
nand U5281 (N_5281,N_4627,N_4598);
nor U5282 (N_5282,N_4607,N_4737);
and U5283 (N_5283,N_4573,N_4745);
nor U5284 (N_5284,N_4942,N_4946);
or U5285 (N_5285,N_4798,N_4573);
and U5286 (N_5286,N_4581,N_4752);
and U5287 (N_5287,N_4691,N_4656);
or U5288 (N_5288,N_4932,N_4854);
nor U5289 (N_5289,N_4711,N_4736);
or U5290 (N_5290,N_4778,N_4946);
and U5291 (N_5291,N_4813,N_4956);
nand U5292 (N_5292,N_4837,N_4593);
nand U5293 (N_5293,N_4881,N_4637);
nand U5294 (N_5294,N_4858,N_4510);
and U5295 (N_5295,N_4656,N_4799);
nand U5296 (N_5296,N_4995,N_4691);
nor U5297 (N_5297,N_4722,N_4538);
or U5298 (N_5298,N_4570,N_4878);
nand U5299 (N_5299,N_4720,N_4850);
nand U5300 (N_5300,N_4645,N_4998);
nand U5301 (N_5301,N_4930,N_4780);
nand U5302 (N_5302,N_4776,N_4981);
xor U5303 (N_5303,N_4808,N_4648);
and U5304 (N_5304,N_4508,N_4552);
or U5305 (N_5305,N_4653,N_4691);
and U5306 (N_5306,N_4650,N_4657);
nor U5307 (N_5307,N_4861,N_4667);
nand U5308 (N_5308,N_4506,N_4963);
xor U5309 (N_5309,N_4949,N_4868);
nor U5310 (N_5310,N_4680,N_4754);
and U5311 (N_5311,N_4724,N_4994);
xor U5312 (N_5312,N_4683,N_4846);
nand U5313 (N_5313,N_4951,N_4630);
nor U5314 (N_5314,N_4835,N_4616);
nor U5315 (N_5315,N_4780,N_4794);
xnor U5316 (N_5316,N_4980,N_4675);
and U5317 (N_5317,N_4993,N_4729);
nand U5318 (N_5318,N_4922,N_4754);
nand U5319 (N_5319,N_4546,N_4662);
nor U5320 (N_5320,N_4731,N_4821);
xor U5321 (N_5321,N_4815,N_4779);
and U5322 (N_5322,N_4888,N_4930);
nor U5323 (N_5323,N_4855,N_4775);
and U5324 (N_5324,N_4793,N_4638);
nand U5325 (N_5325,N_4601,N_4930);
nand U5326 (N_5326,N_4953,N_4804);
nand U5327 (N_5327,N_4911,N_4789);
and U5328 (N_5328,N_4780,N_4605);
xnor U5329 (N_5329,N_4924,N_4516);
nand U5330 (N_5330,N_4936,N_4648);
or U5331 (N_5331,N_4745,N_4760);
or U5332 (N_5332,N_4664,N_4909);
nand U5333 (N_5333,N_4650,N_4790);
xnor U5334 (N_5334,N_4640,N_4963);
and U5335 (N_5335,N_4692,N_4569);
and U5336 (N_5336,N_4704,N_4663);
nand U5337 (N_5337,N_4585,N_4986);
nand U5338 (N_5338,N_4887,N_4610);
nand U5339 (N_5339,N_4828,N_4926);
and U5340 (N_5340,N_4670,N_4615);
nor U5341 (N_5341,N_4844,N_4895);
nor U5342 (N_5342,N_4812,N_4721);
and U5343 (N_5343,N_4668,N_4583);
or U5344 (N_5344,N_4760,N_4647);
and U5345 (N_5345,N_4675,N_4939);
nor U5346 (N_5346,N_4874,N_4610);
xnor U5347 (N_5347,N_4831,N_4965);
nand U5348 (N_5348,N_4883,N_4780);
nor U5349 (N_5349,N_4883,N_4722);
and U5350 (N_5350,N_4788,N_4552);
or U5351 (N_5351,N_4993,N_4734);
and U5352 (N_5352,N_4545,N_4518);
nand U5353 (N_5353,N_4796,N_4693);
or U5354 (N_5354,N_4953,N_4505);
and U5355 (N_5355,N_4837,N_4565);
and U5356 (N_5356,N_4637,N_4991);
and U5357 (N_5357,N_4784,N_4995);
and U5358 (N_5358,N_4813,N_4683);
and U5359 (N_5359,N_4721,N_4917);
xor U5360 (N_5360,N_4543,N_4632);
nor U5361 (N_5361,N_4550,N_4781);
and U5362 (N_5362,N_4914,N_4618);
nor U5363 (N_5363,N_4583,N_4596);
and U5364 (N_5364,N_4901,N_4929);
and U5365 (N_5365,N_4516,N_4819);
xnor U5366 (N_5366,N_4653,N_4575);
nand U5367 (N_5367,N_4709,N_4507);
nor U5368 (N_5368,N_4769,N_4989);
xor U5369 (N_5369,N_4590,N_4985);
nor U5370 (N_5370,N_4976,N_4927);
nand U5371 (N_5371,N_4593,N_4860);
or U5372 (N_5372,N_4612,N_4918);
and U5373 (N_5373,N_4978,N_4615);
nor U5374 (N_5374,N_4943,N_4628);
nand U5375 (N_5375,N_4871,N_4930);
nor U5376 (N_5376,N_4950,N_4540);
nand U5377 (N_5377,N_4547,N_4648);
nor U5378 (N_5378,N_4896,N_4904);
nand U5379 (N_5379,N_4654,N_4645);
nand U5380 (N_5380,N_4536,N_4504);
and U5381 (N_5381,N_4765,N_4912);
nand U5382 (N_5382,N_4985,N_4505);
nor U5383 (N_5383,N_4702,N_4833);
and U5384 (N_5384,N_4597,N_4796);
or U5385 (N_5385,N_4827,N_4763);
nand U5386 (N_5386,N_4959,N_4987);
nor U5387 (N_5387,N_4930,N_4838);
and U5388 (N_5388,N_4930,N_4575);
nor U5389 (N_5389,N_4665,N_4638);
or U5390 (N_5390,N_4985,N_4604);
nor U5391 (N_5391,N_4908,N_4925);
xnor U5392 (N_5392,N_4550,N_4855);
xnor U5393 (N_5393,N_4787,N_4622);
xnor U5394 (N_5394,N_4504,N_4795);
and U5395 (N_5395,N_4675,N_4836);
xnor U5396 (N_5396,N_4532,N_4587);
nand U5397 (N_5397,N_4929,N_4649);
or U5398 (N_5398,N_4582,N_4926);
nand U5399 (N_5399,N_4770,N_4916);
and U5400 (N_5400,N_4693,N_4551);
xor U5401 (N_5401,N_4625,N_4911);
and U5402 (N_5402,N_4549,N_4997);
xor U5403 (N_5403,N_4574,N_4681);
nand U5404 (N_5404,N_4986,N_4698);
nor U5405 (N_5405,N_4809,N_4533);
nor U5406 (N_5406,N_4890,N_4907);
nand U5407 (N_5407,N_4544,N_4783);
or U5408 (N_5408,N_4923,N_4583);
or U5409 (N_5409,N_4789,N_4608);
and U5410 (N_5410,N_4893,N_4558);
nand U5411 (N_5411,N_4649,N_4981);
and U5412 (N_5412,N_4913,N_4565);
xor U5413 (N_5413,N_4579,N_4805);
nor U5414 (N_5414,N_4633,N_4786);
or U5415 (N_5415,N_4991,N_4685);
or U5416 (N_5416,N_4712,N_4655);
or U5417 (N_5417,N_4732,N_4721);
or U5418 (N_5418,N_4504,N_4940);
nor U5419 (N_5419,N_4961,N_4539);
and U5420 (N_5420,N_4962,N_4911);
and U5421 (N_5421,N_4624,N_4668);
and U5422 (N_5422,N_4926,N_4537);
and U5423 (N_5423,N_4727,N_4996);
or U5424 (N_5424,N_4923,N_4641);
xnor U5425 (N_5425,N_4660,N_4651);
xnor U5426 (N_5426,N_4714,N_4927);
and U5427 (N_5427,N_4964,N_4612);
nand U5428 (N_5428,N_4806,N_4977);
and U5429 (N_5429,N_4861,N_4803);
or U5430 (N_5430,N_4700,N_4973);
and U5431 (N_5431,N_4881,N_4960);
xor U5432 (N_5432,N_4779,N_4931);
and U5433 (N_5433,N_4739,N_4566);
and U5434 (N_5434,N_4910,N_4542);
nor U5435 (N_5435,N_4835,N_4533);
nor U5436 (N_5436,N_4691,N_4667);
nor U5437 (N_5437,N_4982,N_4905);
and U5438 (N_5438,N_4720,N_4980);
or U5439 (N_5439,N_4863,N_4703);
or U5440 (N_5440,N_4860,N_4976);
or U5441 (N_5441,N_4891,N_4600);
nand U5442 (N_5442,N_4658,N_4718);
or U5443 (N_5443,N_4563,N_4786);
or U5444 (N_5444,N_4805,N_4882);
nor U5445 (N_5445,N_4738,N_4934);
and U5446 (N_5446,N_4671,N_4886);
xor U5447 (N_5447,N_4583,N_4798);
and U5448 (N_5448,N_4680,N_4998);
or U5449 (N_5449,N_4782,N_4911);
and U5450 (N_5450,N_4647,N_4583);
nor U5451 (N_5451,N_4898,N_4932);
nand U5452 (N_5452,N_4664,N_4747);
nand U5453 (N_5453,N_4513,N_4948);
or U5454 (N_5454,N_4549,N_4980);
xor U5455 (N_5455,N_4787,N_4775);
and U5456 (N_5456,N_4986,N_4823);
and U5457 (N_5457,N_4903,N_4660);
nor U5458 (N_5458,N_4789,N_4987);
nand U5459 (N_5459,N_4502,N_4941);
nand U5460 (N_5460,N_4709,N_4837);
and U5461 (N_5461,N_4908,N_4649);
nor U5462 (N_5462,N_4826,N_4513);
nand U5463 (N_5463,N_4974,N_4929);
nand U5464 (N_5464,N_4880,N_4969);
nor U5465 (N_5465,N_4919,N_4847);
nor U5466 (N_5466,N_4630,N_4536);
and U5467 (N_5467,N_4956,N_4955);
nand U5468 (N_5468,N_4869,N_4646);
and U5469 (N_5469,N_4977,N_4584);
nor U5470 (N_5470,N_4670,N_4535);
xnor U5471 (N_5471,N_4730,N_4621);
xnor U5472 (N_5472,N_4870,N_4517);
or U5473 (N_5473,N_4935,N_4778);
or U5474 (N_5474,N_4841,N_4579);
nand U5475 (N_5475,N_4575,N_4669);
and U5476 (N_5476,N_4840,N_4559);
xor U5477 (N_5477,N_4662,N_4776);
and U5478 (N_5478,N_4504,N_4614);
nor U5479 (N_5479,N_4679,N_4598);
nand U5480 (N_5480,N_4960,N_4807);
nor U5481 (N_5481,N_4877,N_4623);
nand U5482 (N_5482,N_4508,N_4798);
or U5483 (N_5483,N_4851,N_4639);
nor U5484 (N_5484,N_4863,N_4748);
nor U5485 (N_5485,N_4777,N_4757);
nor U5486 (N_5486,N_4725,N_4891);
and U5487 (N_5487,N_4623,N_4882);
or U5488 (N_5488,N_4542,N_4764);
and U5489 (N_5489,N_4813,N_4573);
nor U5490 (N_5490,N_4622,N_4590);
xnor U5491 (N_5491,N_4533,N_4700);
nand U5492 (N_5492,N_4625,N_4660);
nor U5493 (N_5493,N_4988,N_4573);
and U5494 (N_5494,N_4900,N_4616);
and U5495 (N_5495,N_4903,N_4576);
nor U5496 (N_5496,N_4676,N_4802);
and U5497 (N_5497,N_4543,N_4647);
nand U5498 (N_5498,N_4777,N_4580);
and U5499 (N_5499,N_4948,N_4900);
and U5500 (N_5500,N_5166,N_5111);
nand U5501 (N_5501,N_5381,N_5206);
nor U5502 (N_5502,N_5077,N_5289);
or U5503 (N_5503,N_5321,N_5019);
nor U5504 (N_5504,N_5026,N_5461);
nor U5505 (N_5505,N_5426,N_5382);
nor U5506 (N_5506,N_5316,N_5408);
nor U5507 (N_5507,N_5148,N_5233);
nand U5508 (N_5508,N_5096,N_5116);
or U5509 (N_5509,N_5303,N_5464);
nor U5510 (N_5510,N_5147,N_5194);
nor U5511 (N_5511,N_5310,N_5252);
nand U5512 (N_5512,N_5475,N_5041);
and U5513 (N_5513,N_5199,N_5442);
nand U5514 (N_5514,N_5372,N_5169);
nand U5515 (N_5515,N_5071,N_5431);
nor U5516 (N_5516,N_5459,N_5055);
nand U5517 (N_5517,N_5030,N_5465);
and U5518 (N_5518,N_5018,N_5181);
and U5519 (N_5519,N_5208,N_5152);
or U5520 (N_5520,N_5110,N_5184);
or U5521 (N_5521,N_5005,N_5339);
nand U5522 (N_5522,N_5423,N_5183);
or U5523 (N_5523,N_5195,N_5102);
xor U5524 (N_5524,N_5226,N_5209);
nor U5525 (N_5525,N_5211,N_5378);
nor U5526 (N_5526,N_5334,N_5035);
nand U5527 (N_5527,N_5419,N_5109);
nor U5528 (N_5528,N_5292,N_5276);
nand U5529 (N_5529,N_5156,N_5369);
nor U5530 (N_5530,N_5498,N_5347);
nor U5531 (N_5531,N_5173,N_5472);
xnor U5532 (N_5532,N_5362,N_5328);
or U5533 (N_5533,N_5477,N_5298);
nand U5534 (N_5534,N_5344,N_5006);
and U5535 (N_5535,N_5064,N_5182);
or U5536 (N_5536,N_5331,N_5001);
or U5537 (N_5537,N_5097,N_5315);
nand U5538 (N_5538,N_5401,N_5313);
nand U5539 (N_5539,N_5371,N_5042);
and U5540 (N_5540,N_5420,N_5330);
or U5541 (N_5541,N_5488,N_5029);
nor U5542 (N_5542,N_5494,N_5449);
and U5543 (N_5543,N_5384,N_5463);
nor U5544 (N_5544,N_5046,N_5403);
and U5545 (N_5545,N_5450,N_5163);
xnor U5546 (N_5546,N_5044,N_5063);
or U5547 (N_5547,N_5370,N_5225);
and U5548 (N_5548,N_5312,N_5364);
nand U5549 (N_5549,N_5227,N_5022);
and U5550 (N_5550,N_5360,N_5485);
nor U5551 (N_5551,N_5231,N_5049);
nand U5552 (N_5552,N_5299,N_5455);
or U5553 (N_5553,N_5380,N_5153);
or U5554 (N_5554,N_5415,N_5348);
nor U5555 (N_5555,N_5297,N_5275);
nor U5556 (N_5556,N_5444,N_5368);
or U5557 (N_5557,N_5132,N_5058);
nor U5558 (N_5558,N_5452,N_5101);
xnor U5559 (N_5559,N_5091,N_5341);
nor U5560 (N_5560,N_5232,N_5155);
nand U5561 (N_5561,N_5363,N_5031);
xor U5562 (N_5562,N_5080,N_5090);
and U5563 (N_5563,N_5069,N_5356);
nor U5564 (N_5564,N_5220,N_5159);
xor U5565 (N_5565,N_5040,N_5456);
and U5566 (N_5566,N_5053,N_5305);
nand U5567 (N_5567,N_5346,N_5004);
or U5568 (N_5568,N_5437,N_5428);
xnor U5569 (N_5569,N_5479,N_5142);
and U5570 (N_5570,N_5061,N_5084);
or U5571 (N_5571,N_5238,N_5411);
nand U5572 (N_5572,N_5272,N_5135);
or U5573 (N_5573,N_5085,N_5447);
nor U5574 (N_5574,N_5083,N_5119);
or U5575 (N_5575,N_5260,N_5066);
or U5576 (N_5576,N_5106,N_5309);
and U5577 (N_5577,N_5244,N_5146);
or U5578 (N_5578,N_5300,N_5373);
nand U5579 (N_5579,N_5425,N_5037);
nand U5580 (N_5580,N_5377,N_5038);
or U5581 (N_5581,N_5074,N_5482);
or U5582 (N_5582,N_5210,N_5120);
nand U5583 (N_5583,N_5468,N_5311);
nand U5584 (N_5584,N_5306,N_5458);
xnor U5585 (N_5585,N_5353,N_5481);
or U5586 (N_5586,N_5251,N_5440);
or U5587 (N_5587,N_5269,N_5336);
nand U5588 (N_5588,N_5392,N_5405);
nor U5589 (N_5589,N_5361,N_5160);
nand U5590 (N_5590,N_5413,N_5154);
and U5591 (N_5591,N_5100,N_5033);
nand U5592 (N_5592,N_5376,N_5054);
and U5593 (N_5593,N_5103,N_5192);
nor U5594 (N_5594,N_5340,N_5067);
and U5595 (N_5595,N_5217,N_5158);
and U5596 (N_5596,N_5245,N_5359);
and U5597 (N_5597,N_5214,N_5234);
nand U5598 (N_5598,N_5414,N_5057);
or U5599 (N_5599,N_5247,N_5060);
and U5600 (N_5600,N_5048,N_5358);
nand U5601 (N_5601,N_5399,N_5435);
and U5602 (N_5602,N_5266,N_5200);
and U5603 (N_5603,N_5324,N_5418);
nor U5604 (N_5604,N_5150,N_5224);
nor U5605 (N_5605,N_5317,N_5137);
nor U5606 (N_5606,N_5172,N_5280);
nor U5607 (N_5607,N_5283,N_5170);
nor U5608 (N_5608,N_5355,N_5186);
nor U5609 (N_5609,N_5439,N_5205);
nand U5610 (N_5610,N_5121,N_5332);
or U5611 (N_5611,N_5079,N_5032);
and U5612 (N_5612,N_5448,N_5478);
and U5613 (N_5613,N_5221,N_5314);
nand U5614 (N_5614,N_5254,N_5015);
or U5615 (N_5615,N_5395,N_5094);
xnor U5616 (N_5616,N_5398,N_5043);
nand U5617 (N_5617,N_5168,N_5118);
or U5618 (N_5618,N_5189,N_5278);
or U5619 (N_5619,N_5213,N_5338);
xnor U5620 (N_5620,N_5255,N_5281);
and U5621 (N_5621,N_5416,N_5129);
or U5622 (N_5622,N_5286,N_5383);
or U5623 (N_5623,N_5375,N_5218);
or U5624 (N_5624,N_5075,N_5107);
nand U5625 (N_5625,N_5284,N_5351);
nor U5626 (N_5626,N_5059,N_5357);
nand U5627 (N_5627,N_5215,N_5157);
nor U5628 (N_5628,N_5323,N_5349);
xor U5629 (N_5629,N_5007,N_5127);
nor U5630 (N_5630,N_5385,N_5124);
and U5631 (N_5631,N_5335,N_5161);
or U5632 (N_5632,N_5396,N_5243);
or U5633 (N_5633,N_5402,N_5222);
xnor U5634 (N_5634,N_5446,N_5089);
nand U5635 (N_5635,N_5434,N_5151);
or U5636 (N_5636,N_5261,N_5443);
nor U5637 (N_5637,N_5268,N_5039);
and U5638 (N_5638,N_5098,N_5009);
nand U5639 (N_5639,N_5149,N_5114);
or U5640 (N_5640,N_5190,N_5493);
and U5641 (N_5641,N_5417,N_5460);
and U5642 (N_5642,N_5092,N_5010);
nor U5643 (N_5643,N_5241,N_5264);
nand U5644 (N_5644,N_5265,N_5457);
nor U5645 (N_5645,N_5027,N_5325);
nand U5646 (N_5646,N_5164,N_5393);
xnor U5647 (N_5647,N_5196,N_5282);
and U5648 (N_5648,N_5424,N_5256);
nand U5649 (N_5649,N_5487,N_5327);
nor U5650 (N_5650,N_5099,N_5014);
or U5651 (N_5651,N_5491,N_5140);
and U5652 (N_5652,N_5117,N_5469);
nand U5653 (N_5653,N_5301,N_5204);
or U5654 (N_5654,N_5145,N_5008);
and U5655 (N_5655,N_5302,N_5259);
nand U5656 (N_5656,N_5441,N_5291);
nand U5657 (N_5657,N_5198,N_5343);
and U5658 (N_5658,N_5175,N_5253);
and U5659 (N_5659,N_5193,N_5484);
nand U5660 (N_5660,N_5236,N_5492);
xnor U5661 (N_5661,N_5342,N_5451);
nand U5662 (N_5662,N_5178,N_5407);
nand U5663 (N_5663,N_5240,N_5133);
nand U5664 (N_5664,N_5017,N_5065);
nand U5665 (N_5665,N_5422,N_5379);
nand U5666 (N_5666,N_5490,N_5144);
or U5667 (N_5667,N_5087,N_5366);
nand U5668 (N_5668,N_5433,N_5390);
nand U5669 (N_5669,N_5165,N_5389);
or U5670 (N_5670,N_5050,N_5445);
or U5671 (N_5671,N_5318,N_5345);
or U5672 (N_5672,N_5427,N_5002);
nor U5673 (N_5673,N_5337,N_5480);
nor U5674 (N_5674,N_5105,N_5082);
and U5675 (N_5675,N_5277,N_5141);
and U5676 (N_5676,N_5257,N_5088);
or U5677 (N_5677,N_5023,N_5122);
or U5678 (N_5678,N_5197,N_5000);
or U5679 (N_5679,N_5179,N_5112);
and U5680 (N_5680,N_5223,N_5270);
nand U5681 (N_5681,N_5497,N_5136);
nand U5682 (N_5682,N_5134,N_5454);
or U5683 (N_5683,N_5476,N_5406);
nand U5684 (N_5684,N_5296,N_5421);
nor U5685 (N_5685,N_5410,N_5262);
nand U5686 (N_5686,N_5285,N_5081);
and U5687 (N_5687,N_5025,N_5185);
nor U5688 (N_5688,N_5430,N_5020);
or U5689 (N_5689,N_5391,N_5212);
or U5690 (N_5690,N_5139,N_5216);
and U5691 (N_5691,N_5271,N_5070);
and U5692 (N_5692,N_5201,N_5354);
and U5693 (N_5693,N_5350,N_5436);
and U5694 (N_5694,N_5219,N_5237);
or U5695 (N_5695,N_5486,N_5294);
nor U5696 (N_5696,N_5429,N_5187);
and U5697 (N_5697,N_5125,N_5052);
nor U5698 (N_5698,N_5326,N_5273);
or U5699 (N_5699,N_5320,N_5388);
and U5700 (N_5700,N_5180,N_5235);
or U5701 (N_5701,N_5086,N_5466);
and U5702 (N_5702,N_5304,N_5287);
or U5703 (N_5703,N_5267,N_5365);
xnor U5704 (N_5704,N_5467,N_5387);
nor U5705 (N_5705,N_5462,N_5228);
xnor U5706 (N_5706,N_5333,N_5489);
and U5707 (N_5707,N_5239,N_5177);
or U5708 (N_5708,N_5034,N_5138);
nand U5709 (N_5709,N_5412,N_5036);
and U5710 (N_5710,N_5246,N_5288);
nor U5711 (N_5711,N_5474,N_5352);
nor U5712 (N_5712,N_5248,N_5404);
nor U5713 (N_5713,N_5308,N_5013);
nand U5714 (N_5714,N_5113,N_5374);
and U5715 (N_5715,N_5295,N_5409);
or U5716 (N_5716,N_5095,N_5016);
nor U5717 (N_5717,N_5400,N_5191);
nor U5718 (N_5718,N_5207,N_5051);
and U5719 (N_5719,N_5068,N_5115);
xnor U5720 (N_5720,N_5062,N_5496);
nor U5721 (N_5721,N_5499,N_5078);
nand U5722 (N_5722,N_5274,N_5011);
nand U5723 (N_5723,N_5174,N_5203);
or U5724 (N_5724,N_5045,N_5230);
xnor U5725 (N_5725,N_5003,N_5495);
nand U5726 (N_5726,N_5076,N_5322);
xnor U5727 (N_5727,N_5453,N_5143);
nor U5728 (N_5728,N_5056,N_5073);
xor U5729 (N_5729,N_5471,N_5128);
nand U5730 (N_5730,N_5021,N_5394);
nor U5731 (N_5731,N_5131,N_5438);
and U5732 (N_5732,N_5483,N_5104);
and U5733 (N_5733,N_5176,N_5307);
nor U5734 (N_5734,N_5123,N_5290);
and U5735 (N_5735,N_5263,N_5047);
and U5736 (N_5736,N_5293,N_5093);
nand U5737 (N_5737,N_5386,N_5171);
nor U5738 (N_5738,N_5012,N_5329);
nand U5739 (N_5739,N_5188,N_5108);
or U5740 (N_5740,N_5072,N_5167);
or U5741 (N_5741,N_5279,N_5202);
nor U5742 (N_5742,N_5249,N_5130);
nor U5743 (N_5743,N_5028,N_5432);
or U5744 (N_5744,N_5242,N_5470);
nand U5745 (N_5745,N_5126,N_5319);
nor U5746 (N_5746,N_5258,N_5024);
xor U5747 (N_5747,N_5367,N_5397);
nand U5748 (N_5748,N_5250,N_5229);
nor U5749 (N_5749,N_5162,N_5473);
nor U5750 (N_5750,N_5143,N_5144);
and U5751 (N_5751,N_5382,N_5354);
xor U5752 (N_5752,N_5464,N_5340);
or U5753 (N_5753,N_5025,N_5445);
nor U5754 (N_5754,N_5469,N_5042);
and U5755 (N_5755,N_5443,N_5038);
or U5756 (N_5756,N_5454,N_5038);
nand U5757 (N_5757,N_5443,N_5324);
nor U5758 (N_5758,N_5483,N_5068);
and U5759 (N_5759,N_5456,N_5028);
nand U5760 (N_5760,N_5376,N_5298);
and U5761 (N_5761,N_5349,N_5338);
and U5762 (N_5762,N_5135,N_5300);
and U5763 (N_5763,N_5120,N_5452);
or U5764 (N_5764,N_5201,N_5003);
nand U5765 (N_5765,N_5298,N_5341);
nor U5766 (N_5766,N_5229,N_5002);
or U5767 (N_5767,N_5470,N_5300);
nor U5768 (N_5768,N_5074,N_5114);
or U5769 (N_5769,N_5081,N_5463);
nand U5770 (N_5770,N_5364,N_5239);
or U5771 (N_5771,N_5365,N_5021);
and U5772 (N_5772,N_5384,N_5271);
or U5773 (N_5773,N_5090,N_5159);
nor U5774 (N_5774,N_5001,N_5342);
nand U5775 (N_5775,N_5248,N_5427);
and U5776 (N_5776,N_5454,N_5239);
xor U5777 (N_5777,N_5139,N_5310);
nor U5778 (N_5778,N_5144,N_5012);
or U5779 (N_5779,N_5357,N_5015);
and U5780 (N_5780,N_5042,N_5232);
nand U5781 (N_5781,N_5308,N_5428);
nand U5782 (N_5782,N_5314,N_5449);
nor U5783 (N_5783,N_5492,N_5054);
or U5784 (N_5784,N_5070,N_5179);
nor U5785 (N_5785,N_5129,N_5017);
xnor U5786 (N_5786,N_5405,N_5112);
nor U5787 (N_5787,N_5018,N_5232);
nand U5788 (N_5788,N_5437,N_5412);
nand U5789 (N_5789,N_5306,N_5060);
and U5790 (N_5790,N_5093,N_5160);
and U5791 (N_5791,N_5380,N_5486);
nand U5792 (N_5792,N_5222,N_5036);
nand U5793 (N_5793,N_5092,N_5155);
and U5794 (N_5794,N_5461,N_5080);
and U5795 (N_5795,N_5049,N_5373);
nor U5796 (N_5796,N_5366,N_5430);
nor U5797 (N_5797,N_5080,N_5210);
nand U5798 (N_5798,N_5262,N_5118);
or U5799 (N_5799,N_5273,N_5399);
xnor U5800 (N_5800,N_5408,N_5412);
and U5801 (N_5801,N_5307,N_5361);
or U5802 (N_5802,N_5231,N_5340);
or U5803 (N_5803,N_5127,N_5175);
nor U5804 (N_5804,N_5046,N_5003);
or U5805 (N_5805,N_5119,N_5140);
nor U5806 (N_5806,N_5017,N_5009);
nor U5807 (N_5807,N_5466,N_5060);
xor U5808 (N_5808,N_5387,N_5470);
and U5809 (N_5809,N_5047,N_5382);
or U5810 (N_5810,N_5313,N_5493);
or U5811 (N_5811,N_5373,N_5219);
nand U5812 (N_5812,N_5070,N_5086);
or U5813 (N_5813,N_5283,N_5234);
and U5814 (N_5814,N_5118,N_5374);
nor U5815 (N_5815,N_5065,N_5076);
nor U5816 (N_5816,N_5370,N_5431);
nand U5817 (N_5817,N_5118,N_5460);
nand U5818 (N_5818,N_5422,N_5473);
nand U5819 (N_5819,N_5274,N_5484);
or U5820 (N_5820,N_5324,N_5257);
and U5821 (N_5821,N_5016,N_5299);
or U5822 (N_5822,N_5395,N_5211);
nand U5823 (N_5823,N_5318,N_5453);
nor U5824 (N_5824,N_5035,N_5096);
nor U5825 (N_5825,N_5175,N_5354);
and U5826 (N_5826,N_5287,N_5030);
nand U5827 (N_5827,N_5220,N_5238);
xnor U5828 (N_5828,N_5147,N_5055);
or U5829 (N_5829,N_5104,N_5184);
or U5830 (N_5830,N_5037,N_5277);
xor U5831 (N_5831,N_5192,N_5004);
or U5832 (N_5832,N_5208,N_5400);
nor U5833 (N_5833,N_5348,N_5330);
or U5834 (N_5834,N_5356,N_5498);
and U5835 (N_5835,N_5282,N_5263);
or U5836 (N_5836,N_5016,N_5307);
or U5837 (N_5837,N_5050,N_5106);
and U5838 (N_5838,N_5397,N_5231);
nor U5839 (N_5839,N_5115,N_5117);
and U5840 (N_5840,N_5120,N_5199);
nor U5841 (N_5841,N_5482,N_5327);
nand U5842 (N_5842,N_5130,N_5037);
or U5843 (N_5843,N_5143,N_5019);
nor U5844 (N_5844,N_5088,N_5210);
xnor U5845 (N_5845,N_5070,N_5327);
or U5846 (N_5846,N_5064,N_5458);
nand U5847 (N_5847,N_5227,N_5099);
and U5848 (N_5848,N_5161,N_5133);
xor U5849 (N_5849,N_5320,N_5274);
and U5850 (N_5850,N_5015,N_5088);
or U5851 (N_5851,N_5276,N_5214);
xor U5852 (N_5852,N_5003,N_5160);
and U5853 (N_5853,N_5034,N_5275);
or U5854 (N_5854,N_5306,N_5030);
nand U5855 (N_5855,N_5299,N_5473);
and U5856 (N_5856,N_5416,N_5242);
or U5857 (N_5857,N_5483,N_5099);
and U5858 (N_5858,N_5152,N_5291);
nor U5859 (N_5859,N_5140,N_5130);
xnor U5860 (N_5860,N_5346,N_5131);
or U5861 (N_5861,N_5409,N_5078);
and U5862 (N_5862,N_5000,N_5176);
nand U5863 (N_5863,N_5319,N_5286);
nor U5864 (N_5864,N_5228,N_5239);
nand U5865 (N_5865,N_5250,N_5444);
xnor U5866 (N_5866,N_5307,N_5066);
nand U5867 (N_5867,N_5153,N_5056);
nand U5868 (N_5868,N_5439,N_5095);
nand U5869 (N_5869,N_5473,N_5325);
or U5870 (N_5870,N_5146,N_5493);
nor U5871 (N_5871,N_5075,N_5032);
nand U5872 (N_5872,N_5163,N_5207);
nand U5873 (N_5873,N_5267,N_5286);
nand U5874 (N_5874,N_5402,N_5456);
nor U5875 (N_5875,N_5415,N_5181);
nand U5876 (N_5876,N_5431,N_5358);
and U5877 (N_5877,N_5476,N_5393);
nor U5878 (N_5878,N_5470,N_5184);
nor U5879 (N_5879,N_5455,N_5357);
and U5880 (N_5880,N_5302,N_5425);
nand U5881 (N_5881,N_5186,N_5078);
or U5882 (N_5882,N_5124,N_5323);
or U5883 (N_5883,N_5036,N_5268);
nor U5884 (N_5884,N_5335,N_5133);
or U5885 (N_5885,N_5011,N_5168);
xnor U5886 (N_5886,N_5034,N_5215);
nor U5887 (N_5887,N_5120,N_5461);
or U5888 (N_5888,N_5455,N_5058);
nand U5889 (N_5889,N_5372,N_5054);
or U5890 (N_5890,N_5035,N_5014);
nor U5891 (N_5891,N_5208,N_5026);
or U5892 (N_5892,N_5482,N_5302);
nor U5893 (N_5893,N_5147,N_5212);
nand U5894 (N_5894,N_5004,N_5490);
nand U5895 (N_5895,N_5487,N_5186);
or U5896 (N_5896,N_5201,N_5097);
and U5897 (N_5897,N_5144,N_5129);
and U5898 (N_5898,N_5202,N_5312);
nor U5899 (N_5899,N_5408,N_5489);
xnor U5900 (N_5900,N_5353,N_5430);
nor U5901 (N_5901,N_5259,N_5491);
or U5902 (N_5902,N_5431,N_5422);
and U5903 (N_5903,N_5259,N_5020);
or U5904 (N_5904,N_5065,N_5035);
nor U5905 (N_5905,N_5200,N_5002);
and U5906 (N_5906,N_5289,N_5172);
nor U5907 (N_5907,N_5176,N_5155);
or U5908 (N_5908,N_5198,N_5414);
nor U5909 (N_5909,N_5064,N_5291);
and U5910 (N_5910,N_5117,N_5364);
and U5911 (N_5911,N_5101,N_5112);
or U5912 (N_5912,N_5423,N_5198);
nand U5913 (N_5913,N_5400,N_5204);
and U5914 (N_5914,N_5020,N_5363);
or U5915 (N_5915,N_5402,N_5261);
nand U5916 (N_5916,N_5149,N_5198);
or U5917 (N_5917,N_5365,N_5039);
nand U5918 (N_5918,N_5383,N_5338);
nor U5919 (N_5919,N_5153,N_5157);
nor U5920 (N_5920,N_5391,N_5364);
xor U5921 (N_5921,N_5358,N_5189);
nor U5922 (N_5922,N_5141,N_5413);
nor U5923 (N_5923,N_5210,N_5199);
nor U5924 (N_5924,N_5029,N_5053);
nor U5925 (N_5925,N_5046,N_5271);
or U5926 (N_5926,N_5391,N_5016);
and U5927 (N_5927,N_5116,N_5382);
xor U5928 (N_5928,N_5056,N_5000);
or U5929 (N_5929,N_5052,N_5305);
nor U5930 (N_5930,N_5425,N_5185);
nand U5931 (N_5931,N_5332,N_5160);
and U5932 (N_5932,N_5103,N_5462);
nor U5933 (N_5933,N_5341,N_5344);
or U5934 (N_5934,N_5422,N_5105);
or U5935 (N_5935,N_5165,N_5093);
or U5936 (N_5936,N_5385,N_5178);
xnor U5937 (N_5937,N_5033,N_5342);
xor U5938 (N_5938,N_5222,N_5212);
nor U5939 (N_5939,N_5110,N_5220);
nand U5940 (N_5940,N_5231,N_5112);
xor U5941 (N_5941,N_5250,N_5333);
and U5942 (N_5942,N_5048,N_5056);
nand U5943 (N_5943,N_5231,N_5278);
nand U5944 (N_5944,N_5011,N_5396);
or U5945 (N_5945,N_5470,N_5318);
nor U5946 (N_5946,N_5452,N_5003);
or U5947 (N_5947,N_5318,N_5480);
and U5948 (N_5948,N_5262,N_5451);
xor U5949 (N_5949,N_5396,N_5205);
nand U5950 (N_5950,N_5271,N_5054);
or U5951 (N_5951,N_5028,N_5189);
nor U5952 (N_5952,N_5260,N_5335);
and U5953 (N_5953,N_5071,N_5216);
or U5954 (N_5954,N_5479,N_5287);
or U5955 (N_5955,N_5177,N_5240);
nor U5956 (N_5956,N_5490,N_5426);
or U5957 (N_5957,N_5265,N_5160);
nand U5958 (N_5958,N_5209,N_5258);
or U5959 (N_5959,N_5105,N_5362);
nand U5960 (N_5960,N_5327,N_5057);
nor U5961 (N_5961,N_5263,N_5115);
nor U5962 (N_5962,N_5459,N_5384);
and U5963 (N_5963,N_5405,N_5290);
nor U5964 (N_5964,N_5420,N_5091);
or U5965 (N_5965,N_5120,N_5251);
nor U5966 (N_5966,N_5437,N_5452);
or U5967 (N_5967,N_5431,N_5230);
nor U5968 (N_5968,N_5132,N_5195);
nor U5969 (N_5969,N_5161,N_5360);
nor U5970 (N_5970,N_5160,N_5140);
or U5971 (N_5971,N_5050,N_5184);
and U5972 (N_5972,N_5339,N_5285);
or U5973 (N_5973,N_5341,N_5474);
nand U5974 (N_5974,N_5309,N_5377);
nand U5975 (N_5975,N_5105,N_5315);
nand U5976 (N_5976,N_5080,N_5347);
and U5977 (N_5977,N_5399,N_5038);
nor U5978 (N_5978,N_5182,N_5116);
or U5979 (N_5979,N_5360,N_5246);
nor U5980 (N_5980,N_5288,N_5291);
and U5981 (N_5981,N_5295,N_5461);
or U5982 (N_5982,N_5362,N_5152);
and U5983 (N_5983,N_5452,N_5331);
and U5984 (N_5984,N_5248,N_5356);
xor U5985 (N_5985,N_5244,N_5095);
and U5986 (N_5986,N_5297,N_5193);
nand U5987 (N_5987,N_5362,N_5150);
and U5988 (N_5988,N_5182,N_5265);
nand U5989 (N_5989,N_5101,N_5357);
nand U5990 (N_5990,N_5480,N_5389);
and U5991 (N_5991,N_5150,N_5023);
or U5992 (N_5992,N_5114,N_5207);
and U5993 (N_5993,N_5058,N_5130);
xnor U5994 (N_5994,N_5337,N_5238);
nor U5995 (N_5995,N_5422,N_5080);
and U5996 (N_5996,N_5439,N_5292);
nand U5997 (N_5997,N_5385,N_5448);
and U5998 (N_5998,N_5336,N_5474);
or U5999 (N_5999,N_5279,N_5311);
nor U6000 (N_6000,N_5720,N_5916);
or U6001 (N_6001,N_5782,N_5640);
nor U6002 (N_6002,N_5899,N_5703);
or U6003 (N_6003,N_5647,N_5966);
or U6004 (N_6004,N_5862,N_5864);
and U6005 (N_6005,N_5616,N_5939);
xnor U6006 (N_6006,N_5543,N_5604);
xnor U6007 (N_6007,N_5929,N_5896);
nand U6008 (N_6008,N_5974,N_5832);
and U6009 (N_6009,N_5749,N_5557);
or U6010 (N_6010,N_5605,N_5767);
nand U6011 (N_6011,N_5865,N_5910);
nand U6012 (N_6012,N_5944,N_5622);
xor U6013 (N_6013,N_5907,N_5756);
nor U6014 (N_6014,N_5694,N_5739);
and U6015 (N_6015,N_5788,N_5702);
or U6016 (N_6016,N_5536,N_5957);
nor U6017 (N_6017,N_5844,N_5838);
nand U6018 (N_6018,N_5985,N_5823);
or U6019 (N_6019,N_5883,N_5728);
nor U6020 (N_6020,N_5869,N_5866);
or U6021 (N_6021,N_5878,N_5982);
nand U6022 (N_6022,N_5665,N_5735);
nor U6023 (N_6023,N_5804,N_5898);
and U6024 (N_6024,N_5583,N_5690);
nand U6025 (N_6025,N_5680,N_5989);
nor U6026 (N_6026,N_5537,N_5600);
or U6027 (N_6027,N_5654,N_5761);
or U6028 (N_6028,N_5691,N_5805);
nand U6029 (N_6029,N_5718,N_5556);
and U6030 (N_6030,N_5533,N_5529);
nand U6031 (N_6031,N_5777,N_5684);
and U6032 (N_6032,N_5711,N_5615);
nand U6033 (N_6033,N_5636,N_5607);
or U6034 (N_6034,N_5752,N_5858);
nor U6035 (N_6035,N_5750,N_5997);
xor U6036 (N_6036,N_5918,N_5980);
nor U6037 (N_6037,N_5975,N_5889);
nand U6038 (N_6038,N_5538,N_5669);
nor U6039 (N_6039,N_5990,N_5521);
and U6040 (N_6040,N_5826,N_5574);
nor U6041 (N_6041,N_5563,N_5504);
or U6042 (N_6042,N_5760,N_5774);
and U6043 (N_6043,N_5695,N_5955);
nand U6044 (N_6044,N_5708,N_5649);
or U6045 (N_6045,N_5935,N_5765);
and U6046 (N_6046,N_5584,N_5599);
and U6047 (N_6047,N_5792,N_5784);
nand U6048 (N_6048,N_5578,N_5836);
and U6049 (N_6049,N_5828,N_5958);
nor U6050 (N_6050,N_5778,N_5868);
nor U6051 (N_6051,N_5902,N_5780);
nor U6052 (N_6052,N_5508,N_5800);
and U6053 (N_6053,N_5895,N_5847);
or U6054 (N_6054,N_5724,N_5968);
nand U6055 (N_6055,N_5517,N_5608);
and U6056 (N_6056,N_5639,N_5839);
or U6057 (N_6057,N_5841,N_5783);
or U6058 (N_6058,N_5790,N_5603);
nand U6059 (N_6059,N_5672,N_5730);
and U6060 (N_6060,N_5950,N_5994);
nand U6061 (N_6061,N_5825,N_5822);
nor U6062 (N_6062,N_5951,N_5808);
nor U6063 (N_6063,N_5632,N_5658);
or U6064 (N_6064,N_5970,N_5803);
or U6065 (N_6065,N_5519,N_5593);
or U6066 (N_6066,N_5725,N_5996);
nand U6067 (N_6067,N_5531,N_5736);
nand U6068 (N_6068,N_5566,N_5676);
and U6069 (N_6069,N_5637,N_5641);
or U6070 (N_6070,N_5675,N_5689);
nor U6071 (N_6071,N_5701,N_5611);
or U6072 (N_6072,N_5511,N_5848);
nand U6073 (N_6073,N_5554,N_5814);
nor U6074 (N_6074,N_5683,N_5635);
and U6075 (N_6075,N_5897,N_5816);
or U6076 (N_6076,N_5522,N_5530);
nand U6077 (N_6077,N_5592,N_5705);
nand U6078 (N_6078,N_5580,N_5706);
xor U6079 (N_6079,N_5967,N_5852);
nand U6080 (N_6080,N_5983,N_5840);
or U6081 (N_6081,N_5875,N_5551);
or U6082 (N_6082,N_5633,N_5853);
nand U6083 (N_6083,N_5885,N_5945);
xor U6084 (N_6084,N_5964,N_5510);
xor U6085 (N_6085,N_5960,N_5936);
and U6086 (N_6086,N_5938,N_5567);
nor U6087 (N_6087,N_5655,N_5573);
xor U6088 (N_6088,N_5717,N_5651);
nor U6089 (N_6089,N_5810,N_5710);
and U6090 (N_6090,N_5714,N_5986);
or U6091 (N_6091,N_5671,N_5661);
or U6092 (N_6092,N_5666,N_5663);
and U6093 (N_6093,N_5667,N_5963);
or U6094 (N_6094,N_5500,N_5913);
nand U6095 (N_6095,N_5995,N_5594);
or U6096 (N_6096,N_5821,N_5894);
nand U6097 (N_6097,N_5953,N_5976);
nand U6098 (N_6098,N_5606,N_5911);
and U6099 (N_6099,N_5870,N_5993);
xnor U6100 (N_6100,N_5506,N_5670);
nand U6101 (N_6101,N_5773,N_5723);
or U6102 (N_6102,N_5771,N_5999);
xnor U6103 (N_6103,N_5571,N_5570);
and U6104 (N_6104,N_5577,N_5696);
and U6105 (N_6105,N_5659,N_5879);
nand U6106 (N_6106,N_5962,N_5729);
xnor U6107 (N_6107,N_5502,N_5795);
nand U6108 (N_6108,N_5948,N_5540);
or U6109 (N_6109,N_5835,N_5732);
nand U6110 (N_6110,N_5751,N_5909);
and U6111 (N_6111,N_5959,N_5877);
and U6112 (N_6112,N_5920,N_5552);
nor U6113 (N_6113,N_5686,N_5564);
nor U6114 (N_6114,N_5743,N_5861);
or U6115 (N_6115,N_5988,N_5890);
nor U6116 (N_6116,N_5619,N_5681);
nand U6117 (N_6117,N_5768,N_5638);
xnor U6118 (N_6118,N_5591,N_5892);
and U6119 (N_6119,N_5643,N_5534);
xor U6120 (N_6120,N_5807,N_5523);
and U6121 (N_6121,N_5933,N_5733);
and U6122 (N_6122,N_5634,N_5516);
or U6123 (N_6123,N_5561,N_5715);
nor U6124 (N_6124,N_5772,N_5785);
nor U6125 (N_6125,N_5978,N_5559);
nand U6126 (N_6126,N_5770,N_5548);
nor U6127 (N_6127,N_5520,N_5811);
and U6128 (N_6128,N_5871,N_5819);
nand U6129 (N_6129,N_5679,N_5704);
nand U6130 (N_6130,N_5941,N_5503);
and U6131 (N_6131,N_5824,N_5699);
or U6132 (N_6132,N_5830,N_5569);
and U6133 (N_6133,N_5558,N_5856);
or U6134 (N_6134,N_5582,N_5553);
nor U6135 (N_6135,N_5642,N_5940);
nor U6136 (N_6136,N_5542,N_5881);
and U6137 (N_6137,N_5812,N_5602);
nand U6138 (N_6138,N_5737,N_5906);
xnor U6139 (N_6139,N_5587,N_5646);
and U6140 (N_6140,N_5834,N_5682);
or U6141 (N_6141,N_5693,N_5707);
nand U6142 (N_6142,N_5741,N_5586);
nor U6143 (N_6143,N_5555,N_5798);
nor U6144 (N_6144,N_5727,N_5601);
and U6145 (N_6145,N_5507,N_5860);
nor U6146 (N_6146,N_5793,N_5598);
and U6147 (N_6147,N_5901,N_5747);
nor U6148 (N_6148,N_5719,N_5886);
and U6149 (N_6149,N_5796,N_5512);
or U6150 (N_6150,N_5677,N_5917);
or U6151 (N_6151,N_5734,N_5954);
and U6152 (N_6152,N_5923,N_5546);
or U6153 (N_6153,N_5596,N_5597);
and U6154 (N_6154,N_5656,N_5757);
or U6155 (N_6155,N_5755,N_5541);
and U6156 (N_6156,N_5514,N_5509);
nand U6157 (N_6157,N_5664,N_5738);
xnor U6158 (N_6158,N_5524,N_5874);
or U6159 (N_6159,N_5932,N_5905);
and U6160 (N_6160,N_5998,N_5742);
or U6161 (N_6161,N_5882,N_5891);
nor U6162 (N_6162,N_5872,N_5662);
or U6163 (N_6163,N_5972,N_5873);
and U6164 (N_6164,N_5786,N_5539);
and U6165 (N_6165,N_5965,N_5513);
nor U6166 (N_6166,N_5947,N_5745);
nand U6167 (N_6167,N_5588,N_5575);
nor U6168 (N_6168,N_5748,N_5697);
nand U6169 (N_6169,N_5722,N_5802);
or U6170 (N_6170,N_5806,N_5726);
and U6171 (N_6171,N_5781,N_5937);
nor U6172 (N_6172,N_5562,N_5903);
nor U6173 (N_6173,N_5581,N_5627);
nand U6174 (N_6174,N_5549,N_5921);
nor U6175 (N_6175,N_5831,N_5766);
nor U6176 (N_6176,N_5893,N_5992);
nor U6177 (N_6177,N_5623,N_5956);
and U6178 (N_6178,N_5618,N_5753);
nand U6179 (N_6179,N_5845,N_5759);
nand U6180 (N_6180,N_5712,N_5888);
nand U6181 (N_6181,N_5934,N_5946);
or U6182 (N_6182,N_5673,N_5762);
and U6183 (N_6183,N_5949,N_5977);
or U6184 (N_6184,N_5721,N_5652);
nand U6185 (N_6185,N_5709,N_5535);
or U6186 (N_6186,N_5688,N_5746);
or U6187 (N_6187,N_5629,N_5981);
nand U6188 (N_6188,N_5579,N_5791);
nand U6189 (N_6189,N_5769,N_5685);
and U6190 (N_6190,N_5797,N_5621);
and U6191 (N_6191,N_5501,N_5775);
xnor U6192 (N_6192,N_5943,N_5789);
or U6193 (N_6193,N_5987,N_5952);
nand U6194 (N_6194,N_5973,N_5863);
xnor U6195 (N_6195,N_5532,N_5855);
nand U6196 (N_6196,N_5813,N_5763);
and U6197 (N_6197,N_5908,N_5630);
nor U6198 (N_6198,N_5799,N_5776);
or U6199 (N_6199,N_5827,N_5713);
nand U6200 (N_6200,N_5505,N_5758);
and U6201 (N_6201,N_5809,N_5614);
xnor U6202 (N_6202,N_5849,N_5912);
xor U6203 (N_6203,N_5609,N_5590);
and U6204 (N_6204,N_5820,N_5927);
nor U6205 (N_6205,N_5731,N_5984);
or U6206 (N_6206,N_5700,N_5518);
nor U6207 (N_6207,N_5924,N_5887);
xnor U6208 (N_6208,N_5687,N_5678);
nand U6209 (N_6209,N_5931,N_5589);
nor U6210 (N_6210,N_5880,N_5926);
nand U6211 (N_6211,N_5833,N_5595);
and U6212 (N_6212,N_5648,N_5801);
nor U6213 (N_6213,N_5779,N_5744);
nor U6214 (N_6214,N_5547,N_5650);
nand U6215 (N_6215,N_5837,N_5843);
nor U6216 (N_6216,N_5613,N_5829);
nor U6217 (N_6217,N_5928,N_5617);
nand U6218 (N_6218,N_5930,N_5979);
and U6219 (N_6219,N_5526,N_5674);
and U6220 (N_6220,N_5740,N_5854);
or U6221 (N_6221,N_5969,N_5900);
nor U6222 (N_6222,N_5550,N_5585);
and U6223 (N_6223,N_5612,N_5645);
nand U6224 (N_6224,N_5942,N_5818);
and U6225 (N_6225,N_5817,N_5624);
nor U6226 (N_6226,N_5925,N_5857);
nor U6227 (N_6227,N_5787,N_5922);
nor U6228 (N_6228,N_5545,N_5884);
or U6229 (N_6229,N_5653,N_5867);
nand U6230 (N_6230,N_5568,N_5851);
nor U6231 (N_6231,N_5644,N_5914);
nand U6232 (N_6232,N_5842,N_5631);
nand U6233 (N_6233,N_5576,N_5657);
xor U6234 (N_6234,N_5692,N_5620);
and U6235 (N_6235,N_5859,N_5716);
nor U6236 (N_6236,N_5626,N_5560);
nor U6237 (N_6237,N_5991,N_5846);
nor U6238 (N_6238,N_5698,N_5660);
nand U6239 (N_6239,N_5961,N_5610);
and U6240 (N_6240,N_5544,N_5628);
or U6241 (N_6241,N_5764,N_5565);
nand U6242 (N_6242,N_5794,N_5876);
nand U6243 (N_6243,N_5625,N_5971);
nand U6244 (N_6244,N_5919,N_5915);
or U6245 (N_6245,N_5572,N_5815);
or U6246 (N_6246,N_5515,N_5850);
nor U6247 (N_6247,N_5754,N_5904);
or U6248 (N_6248,N_5528,N_5668);
nor U6249 (N_6249,N_5527,N_5525);
nand U6250 (N_6250,N_5747,N_5634);
or U6251 (N_6251,N_5761,N_5525);
nor U6252 (N_6252,N_5821,N_5513);
or U6253 (N_6253,N_5965,N_5842);
or U6254 (N_6254,N_5693,N_5639);
nand U6255 (N_6255,N_5868,N_5949);
or U6256 (N_6256,N_5577,N_5521);
and U6257 (N_6257,N_5958,N_5942);
nor U6258 (N_6258,N_5611,N_5928);
nand U6259 (N_6259,N_5988,N_5525);
and U6260 (N_6260,N_5838,N_5898);
or U6261 (N_6261,N_5695,N_5971);
nand U6262 (N_6262,N_5608,N_5682);
xor U6263 (N_6263,N_5840,N_5979);
nand U6264 (N_6264,N_5884,N_5757);
or U6265 (N_6265,N_5869,N_5782);
xor U6266 (N_6266,N_5814,N_5857);
and U6267 (N_6267,N_5662,N_5817);
and U6268 (N_6268,N_5895,N_5666);
xor U6269 (N_6269,N_5969,N_5509);
and U6270 (N_6270,N_5725,N_5559);
and U6271 (N_6271,N_5598,N_5799);
and U6272 (N_6272,N_5930,N_5677);
nand U6273 (N_6273,N_5528,N_5597);
nor U6274 (N_6274,N_5575,N_5528);
xor U6275 (N_6275,N_5914,N_5517);
xnor U6276 (N_6276,N_5973,N_5609);
and U6277 (N_6277,N_5873,N_5776);
and U6278 (N_6278,N_5759,N_5558);
nor U6279 (N_6279,N_5570,N_5697);
and U6280 (N_6280,N_5918,N_5740);
nor U6281 (N_6281,N_5606,N_5585);
nand U6282 (N_6282,N_5983,N_5804);
and U6283 (N_6283,N_5866,N_5888);
and U6284 (N_6284,N_5563,N_5942);
or U6285 (N_6285,N_5987,N_5509);
nand U6286 (N_6286,N_5672,N_5777);
xnor U6287 (N_6287,N_5578,N_5714);
nand U6288 (N_6288,N_5785,N_5748);
and U6289 (N_6289,N_5971,N_5513);
nand U6290 (N_6290,N_5649,N_5963);
or U6291 (N_6291,N_5739,N_5955);
nor U6292 (N_6292,N_5927,N_5908);
nand U6293 (N_6293,N_5596,N_5688);
xnor U6294 (N_6294,N_5814,N_5786);
or U6295 (N_6295,N_5508,N_5624);
and U6296 (N_6296,N_5811,N_5659);
nor U6297 (N_6297,N_5660,N_5999);
nand U6298 (N_6298,N_5591,N_5933);
nor U6299 (N_6299,N_5942,N_5789);
nand U6300 (N_6300,N_5939,N_5628);
nor U6301 (N_6301,N_5702,N_5676);
or U6302 (N_6302,N_5653,N_5594);
or U6303 (N_6303,N_5550,N_5972);
and U6304 (N_6304,N_5821,N_5993);
and U6305 (N_6305,N_5780,N_5626);
nor U6306 (N_6306,N_5565,N_5550);
and U6307 (N_6307,N_5873,N_5768);
nor U6308 (N_6308,N_5718,N_5982);
nor U6309 (N_6309,N_5826,N_5972);
or U6310 (N_6310,N_5736,N_5805);
or U6311 (N_6311,N_5630,N_5771);
or U6312 (N_6312,N_5645,N_5708);
nand U6313 (N_6313,N_5630,N_5653);
xnor U6314 (N_6314,N_5959,N_5626);
and U6315 (N_6315,N_5529,N_5892);
nand U6316 (N_6316,N_5767,N_5985);
and U6317 (N_6317,N_5955,N_5724);
nand U6318 (N_6318,N_5975,N_5781);
nor U6319 (N_6319,N_5609,N_5597);
and U6320 (N_6320,N_5772,N_5627);
and U6321 (N_6321,N_5758,N_5646);
nor U6322 (N_6322,N_5998,N_5932);
nor U6323 (N_6323,N_5817,N_5763);
nor U6324 (N_6324,N_5655,N_5510);
nand U6325 (N_6325,N_5794,N_5910);
nor U6326 (N_6326,N_5602,N_5965);
or U6327 (N_6327,N_5847,N_5765);
or U6328 (N_6328,N_5935,N_5949);
or U6329 (N_6329,N_5882,N_5611);
nor U6330 (N_6330,N_5941,N_5595);
and U6331 (N_6331,N_5557,N_5660);
nor U6332 (N_6332,N_5749,N_5604);
nor U6333 (N_6333,N_5897,N_5975);
xor U6334 (N_6334,N_5650,N_5973);
xor U6335 (N_6335,N_5581,N_5615);
xnor U6336 (N_6336,N_5859,N_5660);
or U6337 (N_6337,N_5683,N_5523);
and U6338 (N_6338,N_5872,N_5816);
and U6339 (N_6339,N_5640,N_5639);
nor U6340 (N_6340,N_5975,N_5627);
or U6341 (N_6341,N_5708,N_5772);
nor U6342 (N_6342,N_5816,N_5892);
and U6343 (N_6343,N_5537,N_5990);
or U6344 (N_6344,N_5513,N_5892);
nand U6345 (N_6345,N_5757,N_5736);
nand U6346 (N_6346,N_5764,N_5762);
nand U6347 (N_6347,N_5865,N_5593);
and U6348 (N_6348,N_5839,N_5860);
nor U6349 (N_6349,N_5811,N_5531);
nand U6350 (N_6350,N_5923,N_5531);
xor U6351 (N_6351,N_5741,N_5779);
nand U6352 (N_6352,N_5915,N_5631);
nor U6353 (N_6353,N_5589,N_5600);
nand U6354 (N_6354,N_5820,N_5960);
and U6355 (N_6355,N_5666,N_5599);
nor U6356 (N_6356,N_5963,N_5535);
and U6357 (N_6357,N_5952,N_5983);
xnor U6358 (N_6358,N_5609,N_5936);
nand U6359 (N_6359,N_5546,N_5975);
xor U6360 (N_6360,N_5778,N_5871);
nor U6361 (N_6361,N_5928,N_5942);
nand U6362 (N_6362,N_5932,N_5986);
nand U6363 (N_6363,N_5790,N_5550);
nand U6364 (N_6364,N_5963,N_5651);
nand U6365 (N_6365,N_5694,N_5749);
nor U6366 (N_6366,N_5938,N_5940);
nor U6367 (N_6367,N_5940,N_5932);
and U6368 (N_6368,N_5851,N_5977);
nor U6369 (N_6369,N_5858,N_5736);
nor U6370 (N_6370,N_5507,N_5744);
and U6371 (N_6371,N_5749,N_5960);
or U6372 (N_6372,N_5690,N_5542);
or U6373 (N_6373,N_5750,N_5671);
and U6374 (N_6374,N_5815,N_5984);
nand U6375 (N_6375,N_5763,N_5709);
and U6376 (N_6376,N_5845,N_5911);
nand U6377 (N_6377,N_5924,N_5566);
nor U6378 (N_6378,N_5801,N_5850);
or U6379 (N_6379,N_5714,N_5616);
or U6380 (N_6380,N_5553,N_5724);
nand U6381 (N_6381,N_5705,N_5965);
and U6382 (N_6382,N_5965,N_5680);
xor U6383 (N_6383,N_5517,N_5576);
nor U6384 (N_6384,N_5515,N_5969);
nand U6385 (N_6385,N_5851,N_5633);
xor U6386 (N_6386,N_5813,N_5575);
and U6387 (N_6387,N_5863,N_5706);
and U6388 (N_6388,N_5938,N_5805);
nand U6389 (N_6389,N_5709,N_5698);
nor U6390 (N_6390,N_5995,N_5753);
or U6391 (N_6391,N_5581,N_5728);
xnor U6392 (N_6392,N_5763,N_5659);
nor U6393 (N_6393,N_5795,N_5851);
nor U6394 (N_6394,N_5825,N_5859);
or U6395 (N_6395,N_5574,N_5985);
nand U6396 (N_6396,N_5746,N_5957);
xnor U6397 (N_6397,N_5982,N_5665);
and U6398 (N_6398,N_5826,N_5517);
nand U6399 (N_6399,N_5615,N_5765);
or U6400 (N_6400,N_5989,N_5801);
or U6401 (N_6401,N_5979,N_5914);
and U6402 (N_6402,N_5681,N_5978);
nor U6403 (N_6403,N_5553,N_5578);
nor U6404 (N_6404,N_5761,N_5698);
nand U6405 (N_6405,N_5847,N_5967);
nand U6406 (N_6406,N_5855,N_5773);
nor U6407 (N_6407,N_5726,N_5689);
or U6408 (N_6408,N_5939,N_5851);
xnor U6409 (N_6409,N_5787,N_5520);
nand U6410 (N_6410,N_5646,N_5849);
nor U6411 (N_6411,N_5763,N_5625);
or U6412 (N_6412,N_5884,N_5982);
nand U6413 (N_6413,N_5908,N_5529);
and U6414 (N_6414,N_5921,N_5784);
xnor U6415 (N_6415,N_5697,N_5523);
xnor U6416 (N_6416,N_5667,N_5641);
nor U6417 (N_6417,N_5662,N_5737);
nor U6418 (N_6418,N_5972,N_5982);
or U6419 (N_6419,N_5641,N_5557);
nand U6420 (N_6420,N_5705,N_5851);
and U6421 (N_6421,N_5687,N_5890);
nor U6422 (N_6422,N_5902,N_5512);
nor U6423 (N_6423,N_5502,N_5705);
and U6424 (N_6424,N_5662,N_5516);
or U6425 (N_6425,N_5862,N_5528);
nor U6426 (N_6426,N_5696,N_5693);
nor U6427 (N_6427,N_5932,N_5776);
or U6428 (N_6428,N_5650,N_5572);
nand U6429 (N_6429,N_5697,N_5568);
nor U6430 (N_6430,N_5604,N_5522);
and U6431 (N_6431,N_5568,N_5603);
and U6432 (N_6432,N_5813,N_5794);
nand U6433 (N_6433,N_5807,N_5524);
nand U6434 (N_6434,N_5755,N_5811);
or U6435 (N_6435,N_5584,N_5721);
nand U6436 (N_6436,N_5736,N_5893);
nor U6437 (N_6437,N_5560,N_5859);
and U6438 (N_6438,N_5724,N_5785);
nor U6439 (N_6439,N_5984,N_5587);
or U6440 (N_6440,N_5906,N_5825);
or U6441 (N_6441,N_5736,N_5987);
nor U6442 (N_6442,N_5933,N_5688);
nand U6443 (N_6443,N_5575,N_5584);
nor U6444 (N_6444,N_5513,N_5551);
and U6445 (N_6445,N_5775,N_5894);
nor U6446 (N_6446,N_5996,N_5965);
nand U6447 (N_6447,N_5500,N_5566);
nor U6448 (N_6448,N_5540,N_5722);
and U6449 (N_6449,N_5834,N_5914);
and U6450 (N_6450,N_5552,N_5714);
or U6451 (N_6451,N_5963,N_5844);
nor U6452 (N_6452,N_5976,N_5999);
nor U6453 (N_6453,N_5919,N_5837);
nor U6454 (N_6454,N_5535,N_5739);
nor U6455 (N_6455,N_5769,N_5947);
nand U6456 (N_6456,N_5730,N_5958);
or U6457 (N_6457,N_5839,N_5812);
or U6458 (N_6458,N_5568,N_5503);
or U6459 (N_6459,N_5784,N_5741);
nand U6460 (N_6460,N_5861,N_5622);
xor U6461 (N_6461,N_5873,N_5652);
and U6462 (N_6462,N_5651,N_5761);
nor U6463 (N_6463,N_5674,N_5888);
or U6464 (N_6464,N_5943,N_5831);
nand U6465 (N_6465,N_5963,N_5592);
or U6466 (N_6466,N_5763,N_5560);
nor U6467 (N_6467,N_5998,N_5570);
nand U6468 (N_6468,N_5582,N_5605);
or U6469 (N_6469,N_5614,N_5530);
nor U6470 (N_6470,N_5669,N_5867);
nor U6471 (N_6471,N_5696,N_5900);
and U6472 (N_6472,N_5912,N_5949);
xor U6473 (N_6473,N_5731,N_5676);
xnor U6474 (N_6474,N_5530,N_5544);
nor U6475 (N_6475,N_5503,N_5579);
nor U6476 (N_6476,N_5544,N_5722);
or U6477 (N_6477,N_5550,N_5599);
and U6478 (N_6478,N_5938,N_5875);
or U6479 (N_6479,N_5703,N_5865);
nor U6480 (N_6480,N_5571,N_5884);
nand U6481 (N_6481,N_5669,N_5597);
or U6482 (N_6482,N_5616,N_5575);
and U6483 (N_6483,N_5986,N_5841);
and U6484 (N_6484,N_5959,N_5923);
nor U6485 (N_6485,N_5771,N_5622);
or U6486 (N_6486,N_5821,N_5566);
xnor U6487 (N_6487,N_5636,N_5753);
and U6488 (N_6488,N_5620,N_5759);
nor U6489 (N_6489,N_5980,N_5898);
nand U6490 (N_6490,N_5785,N_5693);
or U6491 (N_6491,N_5598,N_5994);
and U6492 (N_6492,N_5563,N_5532);
nand U6493 (N_6493,N_5869,N_5725);
nor U6494 (N_6494,N_5822,N_5687);
and U6495 (N_6495,N_5980,N_5574);
nand U6496 (N_6496,N_5575,N_5782);
nor U6497 (N_6497,N_5560,N_5548);
or U6498 (N_6498,N_5748,N_5714);
and U6499 (N_6499,N_5536,N_5848);
or U6500 (N_6500,N_6454,N_6027);
or U6501 (N_6501,N_6046,N_6243);
or U6502 (N_6502,N_6094,N_6053);
and U6503 (N_6503,N_6019,N_6186);
or U6504 (N_6504,N_6484,N_6364);
nor U6505 (N_6505,N_6340,N_6300);
nor U6506 (N_6506,N_6209,N_6302);
and U6507 (N_6507,N_6346,N_6149);
nand U6508 (N_6508,N_6301,N_6341);
and U6509 (N_6509,N_6328,N_6334);
or U6510 (N_6510,N_6026,N_6411);
nand U6511 (N_6511,N_6034,N_6146);
nand U6512 (N_6512,N_6425,N_6329);
xor U6513 (N_6513,N_6137,N_6294);
nand U6514 (N_6514,N_6433,N_6219);
or U6515 (N_6515,N_6192,N_6071);
nor U6516 (N_6516,N_6499,N_6273);
or U6517 (N_6517,N_6223,N_6274);
nor U6518 (N_6518,N_6405,N_6005);
nor U6519 (N_6519,N_6410,N_6076);
or U6520 (N_6520,N_6052,N_6020);
and U6521 (N_6521,N_6197,N_6256);
or U6522 (N_6522,N_6464,N_6196);
nor U6523 (N_6523,N_6038,N_6259);
xor U6524 (N_6524,N_6080,N_6171);
or U6525 (N_6525,N_6230,N_6073);
xnor U6526 (N_6526,N_6323,N_6443);
or U6527 (N_6527,N_6482,N_6498);
nand U6528 (N_6528,N_6155,N_6078);
nand U6529 (N_6529,N_6041,N_6474);
or U6530 (N_6530,N_6444,N_6199);
and U6531 (N_6531,N_6013,N_6456);
or U6532 (N_6532,N_6287,N_6412);
and U6533 (N_6533,N_6249,N_6255);
and U6534 (N_6534,N_6140,N_6248);
and U6535 (N_6535,N_6158,N_6090);
nor U6536 (N_6536,N_6125,N_6461);
nor U6537 (N_6537,N_6115,N_6106);
nand U6538 (N_6538,N_6194,N_6429);
nand U6539 (N_6539,N_6169,N_6148);
and U6540 (N_6540,N_6067,N_6393);
nand U6541 (N_6541,N_6111,N_6063);
nor U6542 (N_6542,N_6486,N_6206);
xnor U6543 (N_6543,N_6193,N_6124);
and U6544 (N_6544,N_6264,N_6174);
or U6545 (N_6545,N_6320,N_6048);
xor U6546 (N_6546,N_6143,N_6398);
xor U6547 (N_6547,N_6138,N_6134);
nor U6548 (N_6548,N_6350,N_6437);
or U6549 (N_6549,N_6012,N_6254);
nand U6550 (N_6550,N_6397,N_6391);
and U6551 (N_6551,N_6039,N_6387);
and U6552 (N_6552,N_6162,N_6139);
and U6553 (N_6553,N_6372,N_6144);
or U6554 (N_6554,N_6338,N_6316);
nor U6555 (N_6555,N_6151,N_6369);
or U6556 (N_6556,N_6352,N_6252);
or U6557 (N_6557,N_6105,N_6092);
nand U6558 (N_6558,N_6191,N_6023);
nand U6559 (N_6559,N_6070,N_6481);
nor U6560 (N_6560,N_6436,N_6333);
or U6561 (N_6561,N_6044,N_6419);
or U6562 (N_6562,N_6470,N_6003);
and U6563 (N_6563,N_6275,N_6210);
nand U6564 (N_6564,N_6431,N_6430);
nor U6565 (N_6565,N_6141,N_6371);
and U6566 (N_6566,N_6295,N_6326);
or U6567 (N_6567,N_6221,N_6282);
nor U6568 (N_6568,N_6042,N_6361);
and U6569 (N_6569,N_6008,N_6491);
nand U6570 (N_6570,N_6277,N_6135);
xor U6571 (N_6571,N_6228,N_6427);
nor U6572 (N_6572,N_6131,N_6118);
nor U6573 (N_6573,N_6225,N_6406);
or U6574 (N_6574,N_6036,N_6299);
and U6575 (N_6575,N_6010,N_6313);
xor U6576 (N_6576,N_6353,N_6024);
nor U6577 (N_6577,N_6331,N_6347);
nand U6578 (N_6578,N_6428,N_6025);
nor U6579 (N_6579,N_6285,N_6203);
and U6580 (N_6580,N_6463,N_6289);
nand U6581 (N_6581,N_6086,N_6177);
or U6582 (N_6582,N_6385,N_6496);
and U6583 (N_6583,N_6279,N_6460);
xnor U6584 (N_6584,N_6362,N_6327);
or U6585 (N_6585,N_6359,N_6424);
nand U6586 (N_6586,N_6290,N_6104);
nor U6587 (N_6587,N_6168,N_6442);
or U6588 (N_6588,N_6272,N_6035);
and U6589 (N_6589,N_6314,N_6400);
and U6590 (N_6590,N_6207,N_6394);
xnor U6591 (N_6591,N_6417,N_6292);
nand U6592 (N_6592,N_6358,N_6163);
xor U6593 (N_6593,N_6365,N_6257);
nand U6594 (N_6594,N_6122,N_6095);
and U6595 (N_6595,N_6262,N_6332);
or U6596 (N_6596,N_6179,N_6091);
nor U6597 (N_6597,N_6242,N_6483);
or U6598 (N_6598,N_6267,N_6375);
or U6599 (N_6599,N_6176,N_6355);
or U6600 (N_6600,N_6253,N_6478);
xor U6601 (N_6601,N_6445,N_6233);
nor U6602 (N_6602,N_6471,N_6190);
nand U6603 (N_6603,N_6488,N_6297);
nand U6604 (N_6604,N_6084,N_6349);
or U6605 (N_6605,N_6200,N_6421);
nor U6606 (N_6606,N_6093,N_6281);
nor U6607 (N_6607,N_6284,N_6234);
and U6608 (N_6608,N_6455,N_6175);
nor U6609 (N_6609,N_6055,N_6101);
and U6610 (N_6610,N_6344,N_6009);
nor U6611 (N_6611,N_6251,N_6420);
and U6612 (N_6612,N_6030,N_6280);
nand U6613 (N_6613,N_6153,N_6466);
and U6614 (N_6614,N_6475,N_6473);
nor U6615 (N_6615,N_6401,N_6451);
or U6616 (N_6616,N_6107,N_6426);
nor U6617 (N_6617,N_6432,N_6108);
and U6618 (N_6618,N_6268,N_6060);
nand U6619 (N_6619,N_6037,N_6100);
nor U6620 (N_6620,N_6367,N_6172);
or U6621 (N_6621,N_6178,N_6269);
nand U6622 (N_6622,N_6096,N_6380);
and U6623 (N_6623,N_6271,N_6062);
nor U6624 (N_6624,N_6418,N_6069);
and U6625 (N_6625,N_6232,N_6479);
xnor U6626 (N_6626,N_6396,N_6321);
nand U6627 (N_6627,N_6303,N_6258);
nand U6628 (N_6628,N_6363,N_6130);
xor U6629 (N_6629,N_6343,N_6018);
and U6630 (N_6630,N_6117,N_6322);
and U6631 (N_6631,N_6276,N_6357);
nor U6632 (N_6632,N_6377,N_6061);
nand U6633 (N_6633,N_6047,N_6278);
and U6634 (N_6634,N_6469,N_6435);
and U6635 (N_6635,N_6098,N_6029);
or U6636 (N_6636,N_6116,N_6170);
nor U6637 (N_6637,N_6492,N_6182);
nand U6638 (N_6638,N_6497,N_6450);
and U6639 (N_6639,N_6157,N_6184);
and U6640 (N_6640,N_6127,N_6495);
and U6641 (N_6641,N_6214,N_6305);
and U6642 (N_6642,N_6261,N_6065);
and U6643 (N_6643,N_6395,N_6288);
nor U6644 (N_6644,N_6159,N_6336);
and U6645 (N_6645,N_6112,N_6360);
or U6646 (N_6646,N_6114,N_6083);
and U6647 (N_6647,N_6081,N_6054);
and U6648 (N_6648,N_6001,N_6057);
nor U6649 (N_6649,N_6480,N_6485);
or U6650 (N_6650,N_6213,N_6309);
or U6651 (N_6651,N_6216,N_6386);
and U6652 (N_6652,N_6319,N_6468);
and U6653 (N_6653,N_6458,N_6097);
nor U6654 (N_6654,N_6446,N_6247);
and U6655 (N_6655,N_6079,N_6150);
nor U6656 (N_6656,N_6351,N_6298);
xor U6657 (N_6657,N_6066,N_6129);
nand U6658 (N_6658,N_6204,N_6188);
nor U6659 (N_6659,N_6244,N_6161);
nor U6660 (N_6660,N_6465,N_6286);
or U6661 (N_6661,N_6154,N_6235);
nor U6662 (N_6662,N_6147,N_6068);
nor U6663 (N_6663,N_6181,N_6000);
nand U6664 (N_6664,N_6379,N_6021);
or U6665 (N_6665,N_6049,N_6402);
and U6666 (N_6666,N_6490,N_6059);
or U6667 (N_6667,N_6074,N_6165);
and U6668 (N_6668,N_6220,N_6082);
xnor U6669 (N_6669,N_6408,N_6373);
and U6670 (N_6670,N_6310,N_6390);
or U6671 (N_6671,N_6241,N_6342);
nand U6672 (N_6672,N_6102,N_6293);
nor U6673 (N_6673,N_6308,N_6007);
nor U6674 (N_6674,N_6403,N_6245);
nor U6675 (N_6675,N_6337,N_6226);
or U6676 (N_6676,N_6016,N_6173);
nor U6677 (N_6677,N_6006,N_6058);
xnor U6678 (N_6678,N_6325,N_6185);
nand U6679 (N_6679,N_6467,N_6164);
nor U6680 (N_6680,N_6413,N_6315);
or U6681 (N_6681,N_6189,N_6384);
nor U6682 (N_6682,N_6032,N_6142);
xnor U6683 (N_6683,N_6422,N_6453);
nand U6684 (N_6684,N_6033,N_6368);
and U6685 (N_6685,N_6416,N_6156);
nand U6686 (N_6686,N_6407,N_6366);
or U6687 (N_6687,N_6113,N_6075);
or U6688 (N_6688,N_6238,N_6345);
nor U6689 (N_6689,N_6014,N_6447);
or U6690 (N_6690,N_6388,N_6448);
xnor U6691 (N_6691,N_6160,N_6404);
xor U6692 (N_6692,N_6476,N_6123);
nor U6693 (N_6693,N_6459,N_6376);
or U6694 (N_6694,N_6414,N_6283);
and U6695 (N_6695,N_6152,N_6462);
nand U6696 (N_6696,N_6439,N_6103);
nor U6697 (N_6697,N_6056,N_6109);
nor U6698 (N_6698,N_6072,N_6265);
or U6699 (N_6699,N_6227,N_6217);
and U6700 (N_6700,N_6215,N_6064);
or U6701 (N_6701,N_6304,N_6415);
and U6702 (N_6702,N_6317,N_6087);
or U6703 (N_6703,N_6004,N_6354);
nor U6704 (N_6704,N_6452,N_6211);
and U6705 (N_6705,N_6051,N_6240);
nor U6706 (N_6706,N_6339,N_6423);
nand U6707 (N_6707,N_6077,N_6441);
and U6708 (N_6708,N_6399,N_6180);
or U6709 (N_6709,N_6409,N_6183);
xnor U6710 (N_6710,N_6088,N_6166);
nand U6711 (N_6711,N_6040,N_6085);
and U6712 (N_6712,N_6382,N_6002);
or U6713 (N_6713,N_6318,N_6208);
and U6714 (N_6714,N_6434,N_6028);
nand U6715 (N_6715,N_6231,N_6477);
nand U6716 (N_6716,N_6236,N_6187);
nor U6717 (N_6717,N_6222,N_6017);
nor U6718 (N_6718,N_6045,N_6311);
nor U6719 (N_6719,N_6260,N_6306);
nor U6720 (N_6720,N_6120,N_6440);
nand U6721 (N_6721,N_6218,N_6335);
and U6722 (N_6722,N_6145,N_6381);
xor U6723 (N_6723,N_6198,N_6099);
and U6724 (N_6724,N_6121,N_6312);
or U6725 (N_6725,N_6266,N_6307);
or U6726 (N_6726,N_6472,N_6128);
or U6727 (N_6727,N_6229,N_6132);
nand U6728 (N_6728,N_6224,N_6383);
nand U6729 (N_6729,N_6270,N_6202);
or U6730 (N_6730,N_6250,N_6212);
nor U6731 (N_6731,N_6374,N_6126);
or U6732 (N_6732,N_6263,N_6136);
or U6733 (N_6733,N_6296,N_6389);
or U6734 (N_6734,N_6119,N_6457);
nand U6735 (N_6735,N_6205,N_6493);
nor U6736 (N_6736,N_6089,N_6449);
or U6737 (N_6737,N_6167,N_6370);
nand U6738 (N_6738,N_6050,N_6110);
xnor U6739 (N_6739,N_6015,N_6201);
nor U6740 (N_6740,N_6237,N_6489);
nand U6741 (N_6741,N_6392,N_6487);
and U6742 (N_6742,N_6494,N_6239);
xor U6743 (N_6743,N_6246,N_6011);
or U6744 (N_6744,N_6438,N_6356);
and U6745 (N_6745,N_6378,N_6022);
xnor U6746 (N_6746,N_6291,N_6324);
and U6747 (N_6747,N_6133,N_6195);
or U6748 (N_6748,N_6330,N_6348);
nand U6749 (N_6749,N_6031,N_6043);
or U6750 (N_6750,N_6207,N_6078);
nand U6751 (N_6751,N_6081,N_6087);
nor U6752 (N_6752,N_6056,N_6315);
nor U6753 (N_6753,N_6485,N_6002);
and U6754 (N_6754,N_6390,N_6056);
nand U6755 (N_6755,N_6383,N_6122);
nand U6756 (N_6756,N_6409,N_6427);
nand U6757 (N_6757,N_6308,N_6348);
xnor U6758 (N_6758,N_6212,N_6361);
nand U6759 (N_6759,N_6387,N_6240);
or U6760 (N_6760,N_6240,N_6313);
nor U6761 (N_6761,N_6223,N_6288);
and U6762 (N_6762,N_6173,N_6166);
nand U6763 (N_6763,N_6058,N_6132);
nor U6764 (N_6764,N_6277,N_6154);
or U6765 (N_6765,N_6010,N_6378);
and U6766 (N_6766,N_6002,N_6040);
nand U6767 (N_6767,N_6476,N_6222);
or U6768 (N_6768,N_6486,N_6493);
nor U6769 (N_6769,N_6222,N_6434);
and U6770 (N_6770,N_6201,N_6318);
nor U6771 (N_6771,N_6397,N_6178);
nor U6772 (N_6772,N_6189,N_6413);
nor U6773 (N_6773,N_6108,N_6225);
and U6774 (N_6774,N_6104,N_6376);
nor U6775 (N_6775,N_6168,N_6073);
xor U6776 (N_6776,N_6081,N_6286);
nand U6777 (N_6777,N_6011,N_6192);
or U6778 (N_6778,N_6033,N_6221);
or U6779 (N_6779,N_6153,N_6369);
or U6780 (N_6780,N_6156,N_6069);
or U6781 (N_6781,N_6250,N_6156);
xnor U6782 (N_6782,N_6284,N_6486);
nor U6783 (N_6783,N_6479,N_6446);
and U6784 (N_6784,N_6114,N_6480);
nand U6785 (N_6785,N_6204,N_6200);
or U6786 (N_6786,N_6353,N_6151);
nor U6787 (N_6787,N_6305,N_6488);
nor U6788 (N_6788,N_6229,N_6336);
nor U6789 (N_6789,N_6110,N_6489);
and U6790 (N_6790,N_6426,N_6408);
nand U6791 (N_6791,N_6160,N_6440);
nand U6792 (N_6792,N_6134,N_6489);
and U6793 (N_6793,N_6056,N_6395);
nor U6794 (N_6794,N_6471,N_6034);
and U6795 (N_6795,N_6449,N_6159);
nand U6796 (N_6796,N_6311,N_6102);
nand U6797 (N_6797,N_6098,N_6355);
xor U6798 (N_6798,N_6079,N_6165);
or U6799 (N_6799,N_6375,N_6191);
and U6800 (N_6800,N_6113,N_6127);
and U6801 (N_6801,N_6156,N_6383);
nand U6802 (N_6802,N_6437,N_6071);
nand U6803 (N_6803,N_6383,N_6321);
or U6804 (N_6804,N_6118,N_6433);
xor U6805 (N_6805,N_6487,N_6094);
nor U6806 (N_6806,N_6143,N_6406);
or U6807 (N_6807,N_6292,N_6015);
and U6808 (N_6808,N_6427,N_6161);
xor U6809 (N_6809,N_6017,N_6489);
or U6810 (N_6810,N_6476,N_6149);
and U6811 (N_6811,N_6093,N_6096);
and U6812 (N_6812,N_6088,N_6023);
nor U6813 (N_6813,N_6199,N_6401);
or U6814 (N_6814,N_6147,N_6402);
nor U6815 (N_6815,N_6132,N_6481);
nor U6816 (N_6816,N_6474,N_6140);
nand U6817 (N_6817,N_6441,N_6242);
nand U6818 (N_6818,N_6450,N_6454);
nand U6819 (N_6819,N_6188,N_6101);
xor U6820 (N_6820,N_6199,N_6369);
nand U6821 (N_6821,N_6247,N_6226);
nor U6822 (N_6822,N_6010,N_6255);
or U6823 (N_6823,N_6348,N_6415);
nor U6824 (N_6824,N_6431,N_6406);
nor U6825 (N_6825,N_6282,N_6463);
and U6826 (N_6826,N_6219,N_6454);
or U6827 (N_6827,N_6202,N_6486);
and U6828 (N_6828,N_6438,N_6490);
or U6829 (N_6829,N_6411,N_6164);
xnor U6830 (N_6830,N_6452,N_6350);
or U6831 (N_6831,N_6137,N_6362);
and U6832 (N_6832,N_6154,N_6226);
nor U6833 (N_6833,N_6045,N_6088);
or U6834 (N_6834,N_6064,N_6110);
nor U6835 (N_6835,N_6493,N_6341);
or U6836 (N_6836,N_6092,N_6261);
or U6837 (N_6837,N_6260,N_6066);
nand U6838 (N_6838,N_6145,N_6131);
and U6839 (N_6839,N_6463,N_6011);
or U6840 (N_6840,N_6029,N_6441);
and U6841 (N_6841,N_6173,N_6113);
nor U6842 (N_6842,N_6434,N_6354);
nand U6843 (N_6843,N_6258,N_6409);
xnor U6844 (N_6844,N_6163,N_6237);
nor U6845 (N_6845,N_6110,N_6112);
nor U6846 (N_6846,N_6139,N_6257);
nand U6847 (N_6847,N_6288,N_6200);
xor U6848 (N_6848,N_6363,N_6384);
or U6849 (N_6849,N_6167,N_6259);
and U6850 (N_6850,N_6087,N_6305);
xor U6851 (N_6851,N_6049,N_6310);
nor U6852 (N_6852,N_6230,N_6131);
nor U6853 (N_6853,N_6475,N_6364);
nand U6854 (N_6854,N_6158,N_6203);
nor U6855 (N_6855,N_6243,N_6318);
or U6856 (N_6856,N_6117,N_6452);
nor U6857 (N_6857,N_6220,N_6371);
nand U6858 (N_6858,N_6073,N_6475);
xor U6859 (N_6859,N_6049,N_6355);
or U6860 (N_6860,N_6354,N_6351);
nand U6861 (N_6861,N_6293,N_6124);
nor U6862 (N_6862,N_6395,N_6244);
and U6863 (N_6863,N_6379,N_6358);
or U6864 (N_6864,N_6402,N_6030);
and U6865 (N_6865,N_6370,N_6274);
and U6866 (N_6866,N_6025,N_6090);
and U6867 (N_6867,N_6434,N_6006);
nand U6868 (N_6868,N_6400,N_6069);
nor U6869 (N_6869,N_6388,N_6420);
nor U6870 (N_6870,N_6354,N_6262);
nand U6871 (N_6871,N_6239,N_6341);
nor U6872 (N_6872,N_6470,N_6463);
and U6873 (N_6873,N_6073,N_6467);
or U6874 (N_6874,N_6119,N_6120);
xnor U6875 (N_6875,N_6444,N_6467);
xor U6876 (N_6876,N_6018,N_6426);
nor U6877 (N_6877,N_6009,N_6318);
or U6878 (N_6878,N_6464,N_6090);
and U6879 (N_6879,N_6451,N_6165);
nor U6880 (N_6880,N_6095,N_6156);
or U6881 (N_6881,N_6473,N_6201);
nor U6882 (N_6882,N_6079,N_6133);
and U6883 (N_6883,N_6274,N_6039);
and U6884 (N_6884,N_6347,N_6498);
or U6885 (N_6885,N_6200,N_6435);
or U6886 (N_6886,N_6101,N_6355);
and U6887 (N_6887,N_6393,N_6294);
nand U6888 (N_6888,N_6070,N_6352);
xnor U6889 (N_6889,N_6277,N_6234);
and U6890 (N_6890,N_6454,N_6134);
nand U6891 (N_6891,N_6484,N_6190);
and U6892 (N_6892,N_6364,N_6208);
nand U6893 (N_6893,N_6365,N_6070);
or U6894 (N_6894,N_6224,N_6476);
or U6895 (N_6895,N_6177,N_6339);
or U6896 (N_6896,N_6434,N_6454);
xor U6897 (N_6897,N_6224,N_6436);
or U6898 (N_6898,N_6035,N_6159);
nor U6899 (N_6899,N_6334,N_6206);
nor U6900 (N_6900,N_6457,N_6305);
xnor U6901 (N_6901,N_6404,N_6221);
nor U6902 (N_6902,N_6460,N_6105);
or U6903 (N_6903,N_6343,N_6147);
xor U6904 (N_6904,N_6149,N_6056);
nand U6905 (N_6905,N_6041,N_6097);
or U6906 (N_6906,N_6177,N_6375);
or U6907 (N_6907,N_6389,N_6195);
or U6908 (N_6908,N_6259,N_6350);
and U6909 (N_6909,N_6112,N_6077);
nand U6910 (N_6910,N_6313,N_6226);
nor U6911 (N_6911,N_6293,N_6041);
and U6912 (N_6912,N_6110,N_6097);
or U6913 (N_6913,N_6450,N_6046);
or U6914 (N_6914,N_6107,N_6343);
or U6915 (N_6915,N_6217,N_6335);
and U6916 (N_6916,N_6103,N_6486);
nand U6917 (N_6917,N_6001,N_6296);
or U6918 (N_6918,N_6253,N_6434);
and U6919 (N_6919,N_6038,N_6101);
and U6920 (N_6920,N_6399,N_6278);
and U6921 (N_6921,N_6155,N_6016);
nand U6922 (N_6922,N_6383,N_6273);
and U6923 (N_6923,N_6103,N_6219);
nand U6924 (N_6924,N_6479,N_6177);
or U6925 (N_6925,N_6411,N_6177);
or U6926 (N_6926,N_6287,N_6051);
and U6927 (N_6927,N_6454,N_6273);
nand U6928 (N_6928,N_6359,N_6296);
and U6929 (N_6929,N_6383,N_6313);
or U6930 (N_6930,N_6034,N_6311);
or U6931 (N_6931,N_6277,N_6033);
xnor U6932 (N_6932,N_6122,N_6295);
and U6933 (N_6933,N_6308,N_6227);
nand U6934 (N_6934,N_6112,N_6030);
or U6935 (N_6935,N_6432,N_6325);
and U6936 (N_6936,N_6151,N_6281);
or U6937 (N_6937,N_6317,N_6198);
nand U6938 (N_6938,N_6100,N_6380);
nor U6939 (N_6939,N_6364,N_6195);
and U6940 (N_6940,N_6067,N_6112);
nand U6941 (N_6941,N_6163,N_6274);
or U6942 (N_6942,N_6432,N_6074);
nor U6943 (N_6943,N_6187,N_6060);
nand U6944 (N_6944,N_6064,N_6311);
or U6945 (N_6945,N_6288,N_6098);
and U6946 (N_6946,N_6407,N_6063);
and U6947 (N_6947,N_6359,N_6099);
nand U6948 (N_6948,N_6012,N_6164);
or U6949 (N_6949,N_6167,N_6130);
and U6950 (N_6950,N_6119,N_6143);
nor U6951 (N_6951,N_6306,N_6240);
and U6952 (N_6952,N_6494,N_6309);
nor U6953 (N_6953,N_6407,N_6308);
or U6954 (N_6954,N_6228,N_6199);
nand U6955 (N_6955,N_6334,N_6300);
and U6956 (N_6956,N_6386,N_6203);
and U6957 (N_6957,N_6219,N_6438);
nor U6958 (N_6958,N_6496,N_6434);
nand U6959 (N_6959,N_6360,N_6333);
or U6960 (N_6960,N_6489,N_6465);
nand U6961 (N_6961,N_6320,N_6082);
or U6962 (N_6962,N_6297,N_6475);
nor U6963 (N_6963,N_6077,N_6277);
nor U6964 (N_6964,N_6142,N_6053);
or U6965 (N_6965,N_6139,N_6446);
or U6966 (N_6966,N_6069,N_6462);
nor U6967 (N_6967,N_6296,N_6031);
xor U6968 (N_6968,N_6321,N_6154);
and U6969 (N_6969,N_6150,N_6192);
and U6970 (N_6970,N_6489,N_6163);
xnor U6971 (N_6971,N_6062,N_6371);
nand U6972 (N_6972,N_6242,N_6399);
or U6973 (N_6973,N_6278,N_6033);
nand U6974 (N_6974,N_6434,N_6050);
or U6975 (N_6975,N_6156,N_6306);
nand U6976 (N_6976,N_6142,N_6019);
nor U6977 (N_6977,N_6230,N_6096);
nand U6978 (N_6978,N_6105,N_6330);
and U6979 (N_6979,N_6401,N_6470);
nand U6980 (N_6980,N_6034,N_6177);
nand U6981 (N_6981,N_6242,N_6011);
nand U6982 (N_6982,N_6390,N_6336);
nor U6983 (N_6983,N_6320,N_6425);
nand U6984 (N_6984,N_6347,N_6220);
nor U6985 (N_6985,N_6469,N_6048);
nor U6986 (N_6986,N_6328,N_6369);
nor U6987 (N_6987,N_6307,N_6296);
and U6988 (N_6988,N_6497,N_6030);
and U6989 (N_6989,N_6032,N_6209);
or U6990 (N_6990,N_6390,N_6348);
and U6991 (N_6991,N_6105,N_6229);
nor U6992 (N_6992,N_6216,N_6461);
or U6993 (N_6993,N_6071,N_6360);
and U6994 (N_6994,N_6311,N_6374);
or U6995 (N_6995,N_6499,N_6393);
and U6996 (N_6996,N_6126,N_6290);
and U6997 (N_6997,N_6474,N_6471);
nand U6998 (N_6998,N_6103,N_6475);
xor U6999 (N_6999,N_6159,N_6274);
xor U7000 (N_7000,N_6501,N_6701);
xor U7001 (N_7001,N_6585,N_6611);
xor U7002 (N_7002,N_6949,N_6562);
nor U7003 (N_7003,N_6983,N_6583);
nand U7004 (N_7004,N_6979,N_6581);
or U7005 (N_7005,N_6943,N_6755);
nor U7006 (N_7006,N_6894,N_6758);
and U7007 (N_7007,N_6822,N_6871);
nand U7008 (N_7008,N_6750,N_6884);
xor U7009 (N_7009,N_6877,N_6751);
nand U7010 (N_7010,N_6856,N_6941);
xnor U7011 (N_7011,N_6766,N_6610);
and U7012 (N_7012,N_6502,N_6759);
nor U7013 (N_7013,N_6688,N_6764);
and U7014 (N_7014,N_6656,N_6623);
or U7015 (N_7015,N_6748,N_6885);
or U7016 (N_7016,N_6593,N_6878);
and U7017 (N_7017,N_6837,N_6754);
nand U7018 (N_7018,N_6620,N_6913);
and U7019 (N_7019,N_6836,N_6829);
xnor U7020 (N_7020,N_6769,N_6544);
nand U7021 (N_7021,N_6843,N_6712);
nand U7022 (N_7022,N_6537,N_6638);
nand U7023 (N_7023,N_6900,N_6783);
nand U7024 (N_7024,N_6902,N_6917);
xnor U7025 (N_7025,N_6929,N_6503);
or U7026 (N_7026,N_6919,N_6960);
nand U7027 (N_7027,N_6824,N_6765);
nor U7028 (N_7028,N_6592,N_6794);
and U7029 (N_7029,N_6945,N_6613);
and U7030 (N_7030,N_6806,N_6669);
nor U7031 (N_7031,N_6541,N_6668);
and U7032 (N_7032,N_6576,N_6978);
nand U7033 (N_7033,N_6568,N_6863);
nand U7034 (N_7034,N_6851,N_6787);
and U7035 (N_7035,N_6803,N_6634);
and U7036 (N_7036,N_6805,N_6584);
and U7037 (N_7037,N_6704,N_6905);
nand U7038 (N_7038,N_6838,N_6504);
and U7039 (N_7039,N_6814,N_6790);
nand U7040 (N_7040,N_6834,N_6521);
xor U7041 (N_7041,N_6591,N_6912);
nand U7042 (N_7042,N_6703,N_6904);
and U7043 (N_7043,N_6664,N_6647);
and U7044 (N_7044,N_6689,N_6672);
and U7045 (N_7045,N_6670,N_6552);
or U7046 (N_7046,N_6990,N_6626);
nor U7047 (N_7047,N_6791,N_6639);
nor U7048 (N_7048,N_6967,N_6883);
and U7049 (N_7049,N_6932,N_6586);
nand U7050 (N_7050,N_6555,N_6940);
nand U7051 (N_7051,N_6823,N_6588);
xnor U7052 (N_7052,N_6707,N_6965);
nor U7053 (N_7053,N_6994,N_6854);
or U7054 (N_7054,N_6618,N_6529);
or U7055 (N_7055,N_6615,N_6686);
or U7056 (N_7056,N_6849,N_6673);
and U7057 (N_7057,N_6820,N_6525);
nand U7058 (N_7058,N_6880,N_6881);
or U7059 (N_7059,N_6736,N_6889);
nor U7060 (N_7060,N_6564,N_6784);
nand U7061 (N_7061,N_6812,N_6869);
nand U7062 (N_7062,N_6524,N_6977);
nand U7063 (N_7063,N_6918,N_6813);
and U7064 (N_7064,N_6649,N_6685);
and U7065 (N_7065,N_6518,N_6528);
xnor U7066 (N_7066,N_6998,N_6855);
nand U7067 (N_7067,N_6522,N_6780);
nor U7068 (N_7068,N_6507,N_6950);
nand U7069 (N_7069,N_6752,N_6663);
or U7070 (N_7070,N_6538,N_6989);
or U7071 (N_7071,N_6640,N_6879);
nor U7072 (N_7072,N_6840,N_6716);
and U7073 (N_7073,N_6760,N_6852);
or U7074 (N_7074,N_6903,N_6825);
nor U7075 (N_7075,N_6771,N_6891);
and U7076 (N_7076,N_6559,N_6778);
xor U7077 (N_7077,N_6906,N_6582);
nor U7078 (N_7078,N_6832,N_6675);
nand U7079 (N_7079,N_6865,N_6734);
or U7080 (N_7080,N_6898,N_6680);
and U7081 (N_7081,N_6789,N_6678);
and U7082 (N_7082,N_6691,N_6534);
nor U7083 (N_7083,N_6850,N_6733);
or U7084 (N_7084,N_6857,N_6866);
nand U7085 (N_7085,N_6557,N_6775);
nor U7086 (N_7086,N_6781,N_6969);
nand U7087 (N_7087,N_6953,N_6684);
nand U7088 (N_7088,N_6908,N_6531);
nor U7089 (N_7089,N_6819,N_6726);
nand U7090 (N_7090,N_6625,N_6692);
or U7091 (N_7091,N_6946,N_6999);
nand U7092 (N_7092,N_6715,N_6772);
and U7093 (N_7093,N_6867,N_6596);
or U7094 (N_7094,N_6930,N_6710);
or U7095 (N_7095,N_6645,N_6683);
or U7096 (N_7096,N_6594,N_6756);
nor U7097 (N_7097,N_6597,N_6539);
nand U7098 (N_7098,N_6991,N_6655);
or U7099 (N_7099,N_6551,N_6514);
or U7100 (N_7100,N_6792,N_6722);
nand U7101 (N_7101,N_6631,N_6740);
and U7102 (N_7102,N_6810,N_6955);
nand U7103 (N_7103,N_6619,N_6933);
nand U7104 (N_7104,N_6711,N_6926);
nand U7105 (N_7105,N_6637,N_6598);
and U7106 (N_7106,N_6928,N_6723);
nor U7107 (N_7107,N_6509,N_6846);
and U7108 (N_7108,N_6739,N_6616);
or U7109 (N_7109,N_6963,N_6667);
or U7110 (N_7110,N_6811,N_6700);
nand U7111 (N_7111,N_6986,N_6914);
or U7112 (N_7112,N_6817,N_6605);
nand U7113 (N_7113,N_6572,N_6858);
nor U7114 (N_7114,N_6934,N_6951);
or U7115 (N_7115,N_6561,N_6621);
or U7116 (N_7116,N_6779,N_6526);
xnor U7117 (N_7117,N_6622,N_6921);
nor U7118 (N_7118,N_6679,N_6942);
or U7119 (N_7119,N_6705,N_6608);
nor U7120 (N_7120,N_6996,N_6571);
nand U7121 (N_7121,N_6614,N_6962);
and U7122 (N_7122,N_6718,N_6890);
nor U7123 (N_7123,N_6601,N_6827);
nor U7124 (N_7124,N_6872,N_6808);
nand U7125 (N_7125,N_6976,N_6948);
xnor U7126 (N_7126,N_6579,N_6577);
and U7127 (N_7127,N_6801,N_6549);
nor U7128 (N_7128,N_6512,N_6944);
nand U7129 (N_7129,N_6937,N_6882);
and U7130 (N_7130,N_6599,N_6595);
nand U7131 (N_7131,N_6844,N_6627);
or U7132 (N_7132,N_6510,N_6886);
and U7133 (N_7133,N_6785,N_6674);
nand U7134 (N_7134,N_6743,N_6511);
nand U7135 (N_7135,N_6527,N_6578);
nor U7136 (N_7136,N_6624,N_6920);
xor U7137 (N_7137,N_6818,N_6706);
xor U7138 (N_7138,N_6617,N_6687);
and U7139 (N_7139,N_6763,N_6915);
and U7140 (N_7140,N_6826,N_6975);
and U7141 (N_7141,N_6661,N_6516);
or U7142 (N_7142,N_6749,N_6732);
nand U7143 (N_7143,N_6859,N_6606);
and U7144 (N_7144,N_6795,N_6848);
and U7145 (N_7145,N_6609,N_6633);
xnor U7146 (N_7146,N_6652,N_6542);
nor U7147 (N_7147,N_6797,N_6612);
or U7148 (N_7148,N_6788,N_6958);
nand U7149 (N_7149,N_6636,N_6982);
and U7150 (N_7150,N_6782,N_6860);
and U7151 (N_7151,N_6809,N_6676);
and U7152 (N_7152,N_6887,N_6570);
and U7153 (N_7153,N_6554,N_6833);
nand U7154 (N_7154,N_6972,N_6660);
or U7155 (N_7155,N_6657,N_6861);
xnor U7156 (N_7156,N_6658,N_6985);
and U7157 (N_7157,N_6892,N_6796);
and U7158 (N_7158,N_6721,N_6807);
xor U7159 (N_7159,N_6922,N_6973);
nand U7160 (N_7160,N_6517,N_6729);
xnor U7161 (N_7161,N_6506,N_6847);
nand U7162 (N_7162,N_6802,N_6768);
nor U7163 (N_7163,N_6540,N_6747);
nor U7164 (N_7164,N_6776,N_6745);
nor U7165 (N_7165,N_6695,N_6547);
and U7166 (N_7166,N_6635,N_6927);
nand U7167 (N_7167,N_6556,N_6589);
or U7168 (N_7168,N_6828,N_6935);
nor U7169 (N_7169,N_6773,N_6786);
nand U7170 (N_7170,N_6911,N_6862);
xor U7171 (N_7171,N_6909,N_6742);
nor U7172 (N_7172,N_6709,N_6741);
nand U7173 (N_7173,N_6924,N_6961);
nand U7174 (N_7174,N_6799,N_6735);
or U7175 (N_7175,N_6650,N_6800);
nor U7176 (N_7176,N_6708,N_6830);
or U7177 (N_7177,N_6845,N_6519);
and U7178 (N_7178,N_6993,N_6603);
or U7179 (N_7179,N_6550,N_6939);
or U7180 (N_7180,N_6630,N_6984);
nand U7181 (N_7181,N_6901,N_6730);
xnor U7182 (N_7182,N_6717,N_6520);
and U7183 (N_7183,N_6992,N_6746);
and U7184 (N_7184,N_6895,N_6575);
xor U7185 (N_7185,N_6966,N_6956);
nor U7186 (N_7186,N_6697,N_6690);
nand U7187 (N_7187,N_6870,N_6694);
nand U7188 (N_7188,N_6798,N_6565);
and U7189 (N_7189,N_6699,N_6727);
and U7190 (N_7190,N_6713,N_6607);
nand U7191 (N_7191,N_6839,N_6545);
nand U7192 (N_7192,N_6532,N_6659);
nand U7193 (N_7193,N_6767,N_6632);
or U7194 (N_7194,N_6600,N_6648);
or U7195 (N_7195,N_6831,N_6841);
nor U7196 (N_7196,N_6995,N_6896);
nor U7197 (N_7197,N_6629,N_6968);
nand U7198 (N_7198,N_6602,N_6720);
nor U7199 (N_7199,N_6970,N_6677);
and U7200 (N_7200,N_6888,N_6923);
nor U7201 (N_7201,N_6876,N_6777);
or U7202 (N_7202,N_6653,N_6696);
xnor U7203 (N_7203,N_6543,N_6774);
xnor U7204 (N_7204,N_6662,N_6604);
nand U7205 (N_7205,N_6804,N_6580);
nand U7206 (N_7206,N_6558,N_6744);
nor U7207 (N_7207,N_6714,N_6842);
nor U7208 (N_7208,N_6925,N_6573);
nand U7209 (N_7209,N_6642,N_6907);
nor U7210 (N_7210,N_6793,N_6997);
and U7211 (N_7211,N_6931,N_6864);
nor U7212 (N_7212,N_6569,N_6500);
or U7213 (N_7213,N_6553,N_6563);
nor U7214 (N_7214,N_6954,N_6567);
or U7215 (N_7215,N_6587,N_6590);
xor U7216 (N_7216,N_6505,N_6651);
nor U7217 (N_7217,N_6988,N_6835);
nor U7218 (N_7218,N_6853,N_6548);
or U7219 (N_7219,N_6693,N_6974);
or U7220 (N_7220,N_6643,N_6523);
and U7221 (N_7221,N_6654,N_6665);
nor U7222 (N_7222,N_6644,N_6628);
nor U7223 (N_7223,N_6513,N_6536);
nand U7224 (N_7224,N_6725,N_6666);
nor U7225 (N_7225,N_6728,N_6641);
or U7226 (N_7226,N_6761,N_6671);
or U7227 (N_7227,N_6936,N_6508);
or U7228 (N_7228,N_6873,N_6533);
nand U7229 (N_7229,N_6964,N_6702);
nand U7230 (N_7230,N_6762,N_6731);
xnor U7231 (N_7231,N_6770,N_6698);
nand U7232 (N_7232,N_6947,N_6971);
nand U7233 (N_7233,N_6987,N_6959);
and U7234 (N_7234,N_6952,N_6874);
or U7235 (N_7235,N_6899,N_6682);
nor U7236 (N_7236,N_6897,N_6957);
and U7237 (N_7237,N_6560,N_6821);
xor U7238 (N_7238,N_6530,N_6566);
and U7239 (N_7239,N_6681,N_6893);
nand U7240 (N_7240,N_6910,N_6535);
and U7241 (N_7241,N_6719,N_6515);
nand U7242 (N_7242,N_6916,N_6981);
nand U7243 (N_7243,N_6753,N_6646);
nand U7244 (N_7244,N_6724,N_6574);
nand U7245 (N_7245,N_6737,N_6875);
nor U7246 (N_7246,N_6738,N_6816);
or U7247 (N_7247,N_6546,N_6868);
or U7248 (N_7248,N_6938,N_6815);
nand U7249 (N_7249,N_6757,N_6980);
nor U7250 (N_7250,N_6957,N_6507);
and U7251 (N_7251,N_6937,N_6556);
nor U7252 (N_7252,N_6995,N_6808);
nor U7253 (N_7253,N_6504,N_6808);
or U7254 (N_7254,N_6945,N_6857);
nor U7255 (N_7255,N_6895,N_6979);
xnor U7256 (N_7256,N_6876,N_6712);
nor U7257 (N_7257,N_6787,N_6868);
nor U7258 (N_7258,N_6941,N_6629);
and U7259 (N_7259,N_6528,N_6929);
nand U7260 (N_7260,N_6783,N_6986);
and U7261 (N_7261,N_6906,N_6670);
or U7262 (N_7262,N_6820,N_6906);
or U7263 (N_7263,N_6886,N_6712);
or U7264 (N_7264,N_6899,N_6987);
nand U7265 (N_7265,N_6937,N_6894);
or U7266 (N_7266,N_6652,N_6870);
and U7267 (N_7267,N_6615,N_6614);
nor U7268 (N_7268,N_6836,N_6516);
nand U7269 (N_7269,N_6742,N_6548);
nand U7270 (N_7270,N_6532,N_6518);
and U7271 (N_7271,N_6818,N_6880);
or U7272 (N_7272,N_6653,N_6785);
xnor U7273 (N_7273,N_6544,N_6569);
or U7274 (N_7274,N_6721,N_6682);
or U7275 (N_7275,N_6998,N_6694);
nor U7276 (N_7276,N_6553,N_6517);
and U7277 (N_7277,N_6708,N_6759);
or U7278 (N_7278,N_6933,N_6813);
nand U7279 (N_7279,N_6892,N_6872);
nand U7280 (N_7280,N_6597,N_6538);
and U7281 (N_7281,N_6843,N_6541);
xnor U7282 (N_7282,N_6617,N_6916);
nand U7283 (N_7283,N_6934,N_6694);
nor U7284 (N_7284,N_6943,N_6661);
and U7285 (N_7285,N_6863,N_6517);
and U7286 (N_7286,N_6957,N_6509);
nor U7287 (N_7287,N_6976,N_6969);
or U7288 (N_7288,N_6918,N_6730);
nand U7289 (N_7289,N_6706,N_6663);
nor U7290 (N_7290,N_6846,N_6973);
xor U7291 (N_7291,N_6517,N_6921);
or U7292 (N_7292,N_6602,N_6721);
and U7293 (N_7293,N_6920,N_6915);
or U7294 (N_7294,N_6792,N_6754);
nand U7295 (N_7295,N_6537,N_6963);
xnor U7296 (N_7296,N_6633,N_6632);
and U7297 (N_7297,N_6958,N_6847);
xor U7298 (N_7298,N_6778,N_6787);
xnor U7299 (N_7299,N_6668,N_6764);
nand U7300 (N_7300,N_6921,N_6959);
nor U7301 (N_7301,N_6639,N_6711);
nor U7302 (N_7302,N_6621,N_6976);
or U7303 (N_7303,N_6669,N_6723);
and U7304 (N_7304,N_6711,N_6613);
and U7305 (N_7305,N_6634,N_6999);
nand U7306 (N_7306,N_6849,N_6567);
or U7307 (N_7307,N_6867,N_6506);
nor U7308 (N_7308,N_6677,N_6805);
nand U7309 (N_7309,N_6915,N_6555);
or U7310 (N_7310,N_6656,N_6937);
xor U7311 (N_7311,N_6623,N_6969);
and U7312 (N_7312,N_6658,N_6679);
xnor U7313 (N_7313,N_6611,N_6761);
nor U7314 (N_7314,N_6675,N_6831);
or U7315 (N_7315,N_6703,N_6623);
nor U7316 (N_7316,N_6796,N_6671);
or U7317 (N_7317,N_6871,N_6625);
xor U7318 (N_7318,N_6984,N_6840);
or U7319 (N_7319,N_6719,N_6976);
nand U7320 (N_7320,N_6800,N_6691);
and U7321 (N_7321,N_6866,N_6973);
nand U7322 (N_7322,N_6853,N_6925);
or U7323 (N_7323,N_6746,N_6965);
nor U7324 (N_7324,N_6810,N_6563);
and U7325 (N_7325,N_6858,N_6554);
and U7326 (N_7326,N_6507,N_6571);
nand U7327 (N_7327,N_6534,N_6501);
xor U7328 (N_7328,N_6553,N_6509);
nor U7329 (N_7329,N_6532,N_6736);
nor U7330 (N_7330,N_6902,N_6769);
nor U7331 (N_7331,N_6946,N_6826);
or U7332 (N_7332,N_6809,N_6629);
or U7333 (N_7333,N_6654,N_6917);
nand U7334 (N_7334,N_6729,N_6681);
nand U7335 (N_7335,N_6587,N_6659);
and U7336 (N_7336,N_6817,N_6715);
nand U7337 (N_7337,N_6965,N_6827);
nand U7338 (N_7338,N_6792,N_6758);
nor U7339 (N_7339,N_6965,N_6589);
and U7340 (N_7340,N_6852,N_6924);
xor U7341 (N_7341,N_6692,N_6600);
or U7342 (N_7342,N_6992,N_6574);
xor U7343 (N_7343,N_6630,N_6602);
nand U7344 (N_7344,N_6725,N_6967);
nor U7345 (N_7345,N_6961,N_6750);
nor U7346 (N_7346,N_6612,N_6515);
xor U7347 (N_7347,N_6806,N_6850);
or U7348 (N_7348,N_6811,N_6947);
nand U7349 (N_7349,N_6868,N_6792);
nand U7350 (N_7350,N_6878,N_6803);
and U7351 (N_7351,N_6637,N_6646);
or U7352 (N_7352,N_6834,N_6920);
nor U7353 (N_7353,N_6718,N_6903);
and U7354 (N_7354,N_6957,N_6662);
and U7355 (N_7355,N_6589,N_6582);
xnor U7356 (N_7356,N_6736,N_6688);
and U7357 (N_7357,N_6502,N_6728);
xor U7358 (N_7358,N_6673,N_6635);
nand U7359 (N_7359,N_6644,N_6939);
nor U7360 (N_7360,N_6537,N_6989);
or U7361 (N_7361,N_6900,N_6534);
nor U7362 (N_7362,N_6605,N_6865);
or U7363 (N_7363,N_6755,N_6890);
and U7364 (N_7364,N_6968,N_6931);
nor U7365 (N_7365,N_6622,N_6951);
nand U7366 (N_7366,N_6598,N_6883);
or U7367 (N_7367,N_6535,N_6955);
nor U7368 (N_7368,N_6666,N_6844);
nor U7369 (N_7369,N_6573,N_6585);
nand U7370 (N_7370,N_6886,N_6861);
nor U7371 (N_7371,N_6847,N_6712);
nand U7372 (N_7372,N_6569,N_6730);
nor U7373 (N_7373,N_6593,N_6846);
or U7374 (N_7374,N_6574,N_6546);
and U7375 (N_7375,N_6757,N_6700);
nand U7376 (N_7376,N_6705,N_6793);
or U7377 (N_7377,N_6846,N_6576);
or U7378 (N_7378,N_6986,N_6851);
or U7379 (N_7379,N_6620,N_6618);
nand U7380 (N_7380,N_6746,N_6721);
nor U7381 (N_7381,N_6857,N_6969);
or U7382 (N_7382,N_6582,N_6553);
nor U7383 (N_7383,N_6863,N_6687);
and U7384 (N_7384,N_6774,N_6843);
or U7385 (N_7385,N_6899,N_6546);
and U7386 (N_7386,N_6987,N_6782);
or U7387 (N_7387,N_6858,N_6822);
xor U7388 (N_7388,N_6528,N_6710);
or U7389 (N_7389,N_6737,N_6980);
and U7390 (N_7390,N_6874,N_6889);
nand U7391 (N_7391,N_6916,N_6639);
or U7392 (N_7392,N_6565,N_6989);
or U7393 (N_7393,N_6823,N_6822);
or U7394 (N_7394,N_6503,N_6962);
or U7395 (N_7395,N_6901,N_6906);
nor U7396 (N_7396,N_6849,N_6544);
nand U7397 (N_7397,N_6686,N_6563);
nand U7398 (N_7398,N_6828,N_6504);
or U7399 (N_7399,N_6557,N_6862);
or U7400 (N_7400,N_6836,N_6823);
nor U7401 (N_7401,N_6791,N_6687);
nand U7402 (N_7402,N_6812,N_6538);
nand U7403 (N_7403,N_6591,N_6903);
xnor U7404 (N_7404,N_6969,N_6814);
xor U7405 (N_7405,N_6790,N_6656);
nor U7406 (N_7406,N_6957,N_6605);
nand U7407 (N_7407,N_6691,N_6728);
and U7408 (N_7408,N_6683,N_6778);
nand U7409 (N_7409,N_6982,N_6603);
nor U7410 (N_7410,N_6749,N_6596);
or U7411 (N_7411,N_6796,N_6896);
and U7412 (N_7412,N_6612,N_6923);
or U7413 (N_7413,N_6957,N_6693);
and U7414 (N_7414,N_6880,N_6707);
xnor U7415 (N_7415,N_6580,N_6946);
and U7416 (N_7416,N_6702,N_6791);
nand U7417 (N_7417,N_6699,N_6797);
nor U7418 (N_7418,N_6900,N_6562);
xnor U7419 (N_7419,N_6986,N_6647);
xor U7420 (N_7420,N_6913,N_6706);
nand U7421 (N_7421,N_6860,N_6781);
or U7422 (N_7422,N_6877,N_6565);
nor U7423 (N_7423,N_6721,N_6914);
nand U7424 (N_7424,N_6507,N_6883);
and U7425 (N_7425,N_6708,N_6552);
and U7426 (N_7426,N_6673,N_6686);
nor U7427 (N_7427,N_6758,N_6513);
nor U7428 (N_7428,N_6711,N_6650);
or U7429 (N_7429,N_6765,N_6510);
and U7430 (N_7430,N_6671,N_6641);
and U7431 (N_7431,N_6593,N_6782);
and U7432 (N_7432,N_6875,N_6835);
or U7433 (N_7433,N_6608,N_6914);
nand U7434 (N_7434,N_6878,N_6779);
or U7435 (N_7435,N_6818,N_6984);
and U7436 (N_7436,N_6723,N_6982);
or U7437 (N_7437,N_6703,N_6728);
nor U7438 (N_7438,N_6872,N_6718);
and U7439 (N_7439,N_6724,N_6735);
nand U7440 (N_7440,N_6921,N_6544);
nand U7441 (N_7441,N_6813,N_6919);
or U7442 (N_7442,N_6677,N_6799);
nor U7443 (N_7443,N_6655,N_6807);
nand U7444 (N_7444,N_6533,N_6571);
and U7445 (N_7445,N_6633,N_6764);
nor U7446 (N_7446,N_6898,N_6820);
and U7447 (N_7447,N_6720,N_6641);
or U7448 (N_7448,N_6502,N_6738);
and U7449 (N_7449,N_6793,N_6748);
nor U7450 (N_7450,N_6858,N_6680);
or U7451 (N_7451,N_6653,N_6682);
and U7452 (N_7452,N_6974,N_6915);
or U7453 (N_7453,N_6932,N_6745);
nand U7454 (N_7454,N_6765,N_6737);
or U7455 (N_7455,N_6963,N_6916);
or U7456 (N_7456,N_6500,N_6833);
nor U7457 (N_7457,N_6595,N_6721);
nand U7458 (N_7458,N_6523,N_6838);
and U7459 (N_7459,N_6848,N_6971);
and U7460 (N_7460,N_6748,N_6690);
nor U7461 (N_7461,N_6592,N_6737);
or U7462 (N_7462,N_6919,N_6852);
nand U7463 (N_7463,N_6673,N_6696);
or U7464 (N_7464,N_6721,N_6707);
or U7465 (N_7465,N_6646,N_6853);
nor U7466 (N_7466,N_6795,N_6650);
nand U7467 (N_7467,N_6695,N_6702);
or U7468 (N_7468,N_6671,N_6941);
or U7469 (N_7469,N_6761,N_6711);
nor U7470 (N_7470,N_6657,N_6856);
and U7471 (N_7471,N_6916,N_6568);
or U7472 (N_7472,N_6835,N_6643);
nor U7473 (N_7473,N_6740,N_6577);
and U7474 (N_7474,N_6726,N_6570);
or U7475 (N_7475,N_6721,N_6936);
nor U7476 (N_7476,N_6706,N_6573);
or U7477 (N_7477,N_6512,N_6548);
and U7478 (N_7478,N_6692,N_6718);
nor U7479 (N_7479,N_6718,N_6576);
or U7480 (N_7480,N_6843,N_6933);
and U7481 (N_7481,N_6524,N_6690);
nor U7482 (N_7482,N_6786,N_6681);
nand U7483 (N_7483,N_6554,N_6875);
or U7484 (N_7484,N_6873,N_6643);
or U7485 (N_7485,N_6884,N_6629);
or U7486 (N_7486,N_6835,N_6527);
and U7487 (N_7487,N_6713,N_6753);
and U7488 (N_7488,N_6505,N_6729);
and U7489 (N_7489,N_6846,N_6770);
xor U7490 (N_7490,N_6836,N_6755);
xnor U7491 (N_7491,N_6831,N_6815);
nor U7492 (N_7492,N_6846,N_6904);
and U7493 (N_7493,N_6967,N_6690);
and U7494 (N_7494,N_6742,N_6715);
and U7495 (N_7495,N_6738,N_6721);
xor U7496 (N_7496,N_6807,N_6783);
and U7497 (N_7497,N_6988,N_6650);
and U7498 (N_7498,N_6845,N_6850);
xor U7499 (N_7499,N_6505,N_6837);
xnor U7500 (N_7500,N_7336,N_7431);
nand U7501 (N_7501,N_7258,N_7332);
nand U7502 (N_7502,N_7022,N_7048);
nand U7503 (N_7503,N_7040,N_7047);
nand U7504 (N_7504,N_7223,N_7144);
nand U7505 (N_7505,N_7326,N_7139);
nor U7506 (N_7506,N_7013,N_7145);
or U7507 (N_7507,N_7498,N_7006);
nand U7508 (N_7508,N_7333,N_7403);
and U7509 (N_7509,N_7276,N_7103);
or U7510 (N_7510,N_7073,N_7296);
nand U7511 (N_7511,N_7226,N_7133);
nor U7512 (N_7512,N_7000,N_7009);
nand U7513 (N_7513,N_7147,N_7212);
xnor U7514 (N_7514,N_7157,N_7086);
or U7515 (N_7515,N_7135,N_7181);
xor U7516 (N_7516,N_7032,N_7209);
or U7517 (N_7517,N_7076,N_7128);
nand U7518 (N_7518,N_7455,N_7119);
or U7519 (N_7519,N_7480,N_7391);
xnor U7520 (N_7520,N_7429,N_7063);
nand U7521 (N_7521,N_7183,N_7028);
xor U7522 (N_7522,N_7214,N_7065);
nor U7523 (N_7523,N_7051,N_7057);
nand U7524 (N_7524,N_7250,N_7054);
or U7525 (N_7525,N_7140,N_7002);
xor U7526 (N_7526,N_7362,N_7464);
nand U7527 (N_7527,N_7413,N_7395);
nand U7528 (N_7528,N_7421,N_7149);
xnor U7529 (N_7529,N_7487,N_7083);
and U7530 (N_7530,N_7445,N_7475);
and U7531 (N_7531,N_7004,N_7298);
and U7532 (N_7532,N_7059,N_7294);
nor U7533 (N_7533,N_7220,N_7109);
nand U7534 (N_7534,N_7188,N_7217);
and U7535 (N_7535,N_7253,N_7447);
nand U7536 (N_7536,N_7432,N_7330);
or U7537 (N_7537,N_7020,N_7417);
nand U7538 (N_7538,N_7290,N_7191);
nand U7539 (N_7539,N_7353,N_7248);
nor U7540 (N_7540,N_7015,N_7068);
nand U7541 (N_7541,N_7321,N_7152);
nor U7542 (N_7542,N_7104,N_7366);
nor U7543 (N_7543,N_7003,N_7066);
nor U7544 (N_7544,N_7118,N_7303);
nand U7545 (N_7545,N_7268,N_7305);
or U7546 (N_7546,N_7224,N_7393);
and U7547 (N_7547,N_7313,N_7309);
nand U7548 (N_7548,N_7449,N_7189);
nor U7549 (N_7549,N_7277,N_7379);
nand U7550 (N_7550,N_7058,N_7195);
and U7551 (N_7551,N_7461,N_7050);
xor U7552 (N_7552,N_7098,N_7396);
nor U7553 (N_7553,N_7182,N_7237);
or U7554 (N_7554,N_7031,N_7367);
xor U7555 (N_7555,N_7180,N_7433);
or U7556 (N_7556,N_7225,N_7374);
or U7557 (N_7557,N_7018,N_7027);
and U7558 (N_7558,N_7372,N_7173);
and U7559 (N_7559,N_7350,N_7265);
xnor U7560 (N_7560,N_7089,N_7138);
nor U7561 (N_7561,N_7325,N_7358);
nor U7562 (N_7562,N_7206,N_7357);
or U7563 (N_7563,N_7371,N_7067);
xnor U7564 (N_7564,N_7377,N_7151);
and U7565 (N_7565,N_7252,N_7163);
nand U7566 (N_7566,N_7192,N_7115);
xor U7567 (N_7567,N_7482,N_7404);
and U7568 (N_7568,N_7291,N_7084);
xor U7569 (N_7569,N_7438,N_7019);
nand U7570 (N_7570,N_7361,N_7370);
and U7571 (N_7571,N_7123,N_7166);
or U7572 (N_7572,N_7384,N_7196);
nand U7573 (N_7573,N_7499,N_7400);
and U7574 (N_7574,N_7324,N_7427);
nor U7575 (N_7575,N_7478,N_7107);
or U7576 (N_7576,N_7244,N_7348);
and U7577 (N_7577,N_7219,N_7090);
nor U7578 (N_7578,N_7315,N_7342);
xor U7579 (N_7579,N_7130,N_7261);
xnor U7580 (N_7580,N_7092,N_7495);
or U7581 (N_7581,N_7311,N_7402);
and U7582 (N_7582,N_7091,N_7339);
and U7583 (N_7583,N_7093,N_7299);
nor U7584 (N_7584,N_7469,N_7278);
or U7585 (N_7585,N_7233,N_7238);
nand U7586 (N_7586,N_7453,N_7346);
nor U7587 (N_7587,N_7490,N_7352);
nor U7588 (N_7588,N_7046,N_7132);
nor U7589 (N_7589,N_7284,N_7271);
nand U7590 (N_7590,N_7165,N_7312);
and U7591 (N_7591,N_7376,N_7155);
nor U7592 (N_7592,N_7005,N_7425);
xnor U7593 (N_7593,N_7283,N_7441);
nor U7594 (N_7594,N_7460,N_7319);
or U7595 (N_7595,N_7021,N_7443);
nor U7596 (N_7596,N_7125,N_7127);
nand U7597 (N_7597,N_7045,N_7049);
xnor U7598 (N_7598,N_7236,N_7409);
or U7599 (N_7599,N_7136,N_7327);
nand U7600 (N_7600,N_7080,N_7255);
nand U7601 (N_7601,N_7078,N_7288);
nand U7602 (N_7602,N_7269,N_7077);
and U7603 (N_7603,N_7012,N_7286);
or U7604 (N_7604,N_7345,N_7369);
and U7605 (N_7605,N_7412,N_7307);
xor U7606 (N_7606,N_7041,N_7451);
nor U7607 (N_7607,N_7450,N_7401);
or U7608 (N_7608,N_7257,N_7456);
nand U7609 (N_7609,N_7164,N_7174);
or U7610 (N_7610,N_7383,N_7126);
nor U7611 (N_7611,N_7184,N_7198);
nor U7612 (N_7612,N_7231,N_7389);
nand U7613 (N_7613,N_7150,N_7044);
and U7614 (N_7614,N_7017,N_7203);
and U7615 (N_7615,N_7249,N_7262);
nor U7616 (N_7616,N_7210,N_7341);
and U7617 (N_7617,N_7375,N_7197);
nand U7618 (N_7618,N_7070,N_7142);
nand U7619 (N_7619,N_7496,N_7360);
and U7620 (N_7620,N_7486,N_7242);
nor U7621 (N_7621,N_7227,N_7300);
nor U7622 (N_7622,N_7423,N_7484);
or U7623 (N_7623,N_7062,N_7408);
and U7624 (N_7624,N_7069,N_7170);
and U7625 (N_7625,N_7293,N_7179);
or U7626 (N_7626,N_7102,N_7388);
and U7627 (N_7627,N_7285,N_7075);
nor U7628 (N_7628,N_7359,N_7101);
and U7629 (N_7629,N_7010,N_7458);
nor U7630 (N_7630,N_7292,N_7037);
nor U7631 (N_7631,N_7351,N_7052);
nor U7632 (N_7632,N_7426,N_7060);
or U7633 (N_7633,N_7399,N_7202);
or U7634 (N_7634,N_7272,N_7008);
xor U7635 (N_7635,N_7467,N_7082);
nand U7636 (N_7636,N_7323,N_7282);
nor U7637 (N_7637,N_7095,N_7222);
nor U7638 (N_7638,N_7185,N_7161);
nor U7639 (N_7639,N_7235,N_7158);
xnor U7640 (N_7640,N_7175,N_7207);
xor U7641 (N_7641,N_7452,N_7172);
or U7642 (N_7642,N_7422,N_7308);
nor U7643 (N_7643,N_7094,N_7056);
or U7644 (N_7644,N_7039,N_7122);
xor U7645 (N_7645,N_7087,N_7344);
or U7646 (N_7646,N_7477,N_7190);
and U7647 (N_7647,N_7406,N_7025);
and U7648 (N_7648,N_7338,N_7208);
nor U7649 (N_7649,N_7105,N_7167);
xor U7650 (N_7650,N_7416,N_7186);
and U7651 (N_7651,N_7382,N_7218);
and U7652 (N_7652,N_7134,N_7131);
and U7653 (N_7653,N_7430,N_7213);
nor U7654 (N_7654,N_7100,N_7442);
and U7655 (N_7655,N_7153,N_7373);
and U7656 (N_7656,N_7485,N_7034);
and U7657 (N_7657,N_7241,N_7444);
or U7658 (N_7658,N_7042,N_7141);
xor U7659 (N_7659,N_7386,N_7492);
or U7660 (N_7660,N_7378,N_7038);
nor U7661 (N_7661,N_7240,N_7322);
or U7662 (N_7662,N_7023,N_7483);
and U7663 (N_7663,N_7279,N_7194);
and U7664 (N_7664,N_7440,N_7295);
xor U7665 (N_7665,N_7270,N_7439);
and U7666 (N_7666,N_7390,N_7316);
nor U7667 (N_7667,N_7234,N_7494);
xor U7668 (N_7668,N_7178,N_7159);
nand U7669 (N_7669,N_7215,N_7410);
xnor U7670 (N_7670,N_7071,N_7465);
and U7671 (N_7671,N_7053,N_7281);
or U7672 (N_7672,N_7334,N_7424);
nand U7673 (N_7673,N_7074,N_7110);
nor U7674 (N_7674,N_7097,N_7111);
nor U7675 (N_7675,N_7329,N_7267);
xor U7676 (N_7676,N_7437,N_7488);
or U7677 (N_7677,N_7113,N_7474);
nand U7678 (N_7678,N_7254,N_7381);
or U7679 (N_7679,N_7463,N_7304);
nand U7680 (N_7680,N_7489,N_7462);
or U7681 (N_7681,N_7302,N_7435);
or U7682 (N_7682,N_7251,N_7392);
nand U7683 (N_7683,N_7273,N_7448);
nor U7684 (N_7684,N_7216,N_7394);
and U7685 (N_7685,N_7026,N_7274);
nor U7686 (N_7686,N_7414,N_7035);
nor U7687 (N_7687,N_7001,N_7124);
xnor U7688 (N_7688,N_7356,N_7407);
nor U7689 (N_7689,N_7472,N_7201);
and U7690 (N_7690,N_7137,N_7014);
nand U7691 (N_7691,N_7471,N_7232);
nand U7692 (N_7692,N_7256,N_7297);
nand U7693 (N_7693,N_7405,N_7211);
nand U7694 (N_7694,N_7029,N_7385);
and U7695 (N_7695,N_7310,N_7364);
and U7696 (N_7696,N_7036,N_7129);
xor U7697 (N_7697,N_7205,N_7411);
nor U7698 (N_7698,N_7200,N_7317);
nor U7699 (N_7699,N_7148,N_7347);
and U7700 (N_7700,N_7112,N_7363);
nor U7701 (N_7701,N_7055,N_7280);
nor U7702 (N_7702,N_7024,N_7229);
nor U7703 (N_7703,N_7354,N_7072);
nand U7704 (N_7704,N_7420,N_7030);
nor U7705 (N_7705,N_7337,N_7007);
nand U7706 (N_7706,N_7419,N_7289);
or U7707 (N_7707,N_7146,N_7491);
nor U7708 (N_7708,N_7243,N_7368);
and U7709 (N_7709,N_7230,N_7221);
and U7710 (N_7710,N_7454,N_7415);
nand U7711 (N_7711,N_7457,N_7061);
nand U7712 (N_7712,N_7154,N_7320);
nor U7713 (N_7713,N_7318,N_7266);
or U7714 (N_7714,N_7355,N_7120);
or U7715 (N_7715,N_7428,N_7343);
nor U7716 (N_7716,N_7228,N_7088);
or U7717 (N_7717,N_7156,N_7085);
and U7718 (N_7718,N_7239,N_7446);
or U7719 (N_7719,N_7033,N_7116);
and U7720 (N_7720,N_7459,N_7340);
nand U7721 (N_7721,N_7468,N_7177);
and U7722 (N_7722,N_7176,N_7204);
nand U7723 (N_7723,N_7171,N_7143);
nand U7724 (N_7724,N_7434,N_7121);
and U7725 (N_7725,N_7397,N_7479);
nor U7726 (N_7726,N_7466,N_7335);
and U7727 (N_7727,N_7199,N_7011);
or U7728 (N_7728,N_7168,N_7481);
nand U7729 (N_7729,N_7314,N_7247);
nand U7730 (N_7730,N_7064,N_7287);
and U7731 (N_7731,N_7114,N_7260);
xor U7732 (N_7732,N_7436,N_7245);
nor U7733 (N_7733,N_7162,N_7016);
nor U7734 (N_7734,N_7246,N_7263);
nor U7735 (N_7735,N_7328,N_7380);
nor U7736 (N_7736,N_7096,N_7473);
nand U7737 (N_7737,N_7259,N_7476);
and U7738 (N_7738,N_7470,N_7264);
or U7739 (N_7739,N_7160,N_7193);
and U7740 (N_7740,N_7187,N_7306);
or U7741 (N_7741,N_7493,N_7387);
or U7742 (N_7742,N_7108,N_7331);
or U7743 (N_7743,N_7349,N_7081);
nor U7744 (N_7744,N_7497,N_7365);
or U7745 (N_7745,N_7099,N_7043);
nor U7746 (N_7746,N_7301,N_7275);
nand U7747 (N_7747,N_7106,N_7079);
and U7748 (N_7748,N_7169,N_7418);
or U7749 (N_7749,N_7117,N_7398);
and U7750 (N_7750,N_7076,N_7331);
nor U7751 (N_7751,N_7236,N_7294);
nor U7752 (N_7752,N_7139,N_7306);
and U7753 (N_7753,N_7159,N_7055);
or U7754 (N_7754,N_7114,N_7342);
or U7755 (N_7755,N_7116,N_7150);
nand U7756 (N_7756,N_7215,N_7214);
nand U7757 (N_7757,N_7342,N_7162);
or U7758 (N_7758,N_7419,N_7220);
nand U7759 (N_7759,N_7394,N_7085);
nor U7760 (N_7760,N_7451,N_7475);
nand U7761 (N_7761,N_7441,N_7384);
and U7762 (N_7762,N_7267,N_7121);
nor U7763 (N_7763,N_7400,N_7445);
nand U7764 (N_7764,N_7227,N_7242);
and U7765 (N_7765,N_7458,N_7403);
or U7766 (N_7766,N_7209,N_7027);
or U7767 (N_7767,N_7428,N_7223);
or U7768 (N_7768,N_7168,N_7204);
nor U7769 (N_7769,N_7318,N_7079);
xnor U7770 (N_7770,N_7320,N_7092);
or U7771 (N_7771,N_7293,N_7122);
and U7772 (N_7772,N_7201,N_7358);
or U7773 (N_7773,N_7335,N_7032);
or U7774 (N_7774,N_7332,N_7172);
xnor U7775 (N_7775,N_7197,N_7143);
or U7776 (N_7776,N_7397,N_7487);
nand U7777 (N_7777,N_7068,N_7118);
or U7778 (N_7778,N_7490,N_7116);
nand U7779 (N_7779,N_7018,N_7325);
nand U7780 (N_7780,N_7252,N_7414);
and U7781 (N_7781,N_7313,N_7355);
nand U7782 (N_7782,N_7237,N_7204);
nand U7783 (N_7783,N_7083,N_7188);
and U7784 (N_7784,N_7061,N_7020);
nand U7785 (N_7785,N_7429,N_7165);
and U7786 (N_7786,N_7129,N_7004);
nand U7787 (N_7787,N_7075,N_7385);
nor U7788 (N_7788,N_7074,N_7268);
nand U7789 (N_7789,N_7106,N_7363);
nor U7790 (N_7790,N_7293,N_7090);
or U7791 (N_7791,N_7270,N_7130);
or U7792 (N_7792,N_7171,N_7166);
nor U7793 (N_7793,N_7090,N_7197);
xnor U7794 (N_7794,N_7216,N_7202);
or U7795 (N_7795,N_7148,N_7193);
or U7796 (N_7796,N_7107,N_7009);
nor U7797 (N_7797,N_7350,N_7101);
and U7798 (N_7798,N_7047,N_7387);
or U7799 (N_7799,N_7147,N_7479);
or U7800 (N_7800,N_7416,N_7007);
nor U7801 (N_7801,N_7313,N_7138);
nand U7802 (N_7802,N_7335,N_7214);
nor U7803 (N_7803,N_7289,N_7175);
nor U7804 (N_7804,N_7111,N_7170);
and U7805 (N_7805,N_7046,N_7234);
and U7806 (N_7806,N_7314,N_7234);
xor U7807 (N_7807,N_7037,N_7384);
or U7808 (N_7808,N_7173,N_7085);
xor U7809 (N_7809,N_7123,N_7315);
nor U7810 (N_7810,N_7087,N_7448);
nor U7811 (N_7811,N_7129,N_7459);
and U7812 (N_7812,N_7042,N_7257);
nor U7813 (N_7813,N_7270,N_7450);
nor U7814 (N_7814,N_7122,N_7067);
nor U7815 (N_7815,N_7085,N_7269);
or U7816 (N_7816,N_7161,N_7331);
xor U7817 (N_7817,N_7379,N_7056);
nand U7818 (N_7818,N_7192,N_7450);
nor U7819 (N_7819,N_7194,N_7467);
or U7820 (N_7820,N_7222,N_7399);
and U7821 (N_7821,N_7418,N_7373);
nand U7822 (N_7822,N_7196,N_7245);
nand U7823 (N_7823,N_7274,N_7454);
and U7824 (N_7824,N_7050,N_7215);
nor U7825 (N_7825,N_7389,N_7202);
or U7826 (N_7826,N_7495,N_7288);
and U7827 (N_7827,N_7037,N_7474);
and U7828 (N_7828,N_7475,N_7174);
nand U7829 (N_7829,N_7466,N_7117);
or U7830 (N_7830,N_7485,N_7495);
nand U7831 (N_7831,N_7122,N_7040);
nand U7832 (N_7832,N_7282,N_7319);
xnor U7833 (N_7833,N_7403,N_7217);
nor U7834 (N_7834,N_7117,N_7301);
and U7835 (N_7835,N_7009,N_7044);
or U7836 (N_7836,N_7135,N_7209);
nand U7837 (N_7837,N_7496,N_7385);
xnor U7838 (N_7838,N_7187,N_7292);
nor U7839 (N_7839,N_7289,N_7132);
nor U7840 (N_7840,N_7044,N_7134);
nor U7841 (N_7841,N_7256,N_7140);
and U7842 (N_7842,N_7338,N_7440);
xor U7843 (N_7843,N_7414,N_7402);
and U7844 (N_7844,N_7203,N_7379);
nor U7845 (N_7845,N_7317,N_7160);
and U7846 (N_7846,N_7105,N_7065);
and U7847 (N_7847,N_7127,N_7188);
or U7848 (N_7848,N_7290,N_7028);
or U7849 (N_7849,N_7460,N_7055);
or U7850 (N_7850,N_7106,N_7455);
nor U7851 (N_7851,N_7193,N_7135);
nand U7852 (N_7852,N_7169,N_7186);
nand U7853 (N_7853,N_7275,N_7032);
or U7854 (N_7854,N_7393,N_7119);
or U7855 (N_7855,N_7273,N_7478);
or U7856 (N_7856,N_7445,N_7190);
nor U7857 (N_7857,N_7478,N_7117);
xor U7858 (N_7858,N_7193,N_7484);
nor U7859 (N_7859,N_7067,N_7361);
or U7860 (N_7860,N_7135,N_7044);
or U7861 (N_7861,N_7475,N_7228);
and U7862 (N_7862,N_7028,N_7079);
or U7863 (N_7863,N_7151,N_7189);
and U7864 (N_7864,N_7040,N_7471);
or U7865 (N_7865,N_7259,N_7192);
or U7866 (N_7866,N_7256,N_7023);
or U7867 (N_7867,N_7490,N_7147);
nor U7868 (N_7868,N_7488,N_7222);
and U7869 (N_7869,N_7438,N_7316);
or U7870 (N_7870,N_7490,N_7048);
or U7871 (N_7871,N_7016,N_7342);
nor U7872 (N_7872,N_7280,N_7225);
xnor U7873 (N_7873,N_7321,N_7180);
nor U7874 (N_7874,N_7013,N_7315);
or U7875 (N_7875,N_7328,N_7258);
nor U7876 (N_7876,N_7158,N_7327);
and U7877 (N_7877,N_7147,N_7313);
nor U7878 (N_7878,N_7470,N_7281);
and U7879 (N_7879,N_7276,N_7301);
xor U7880 (N_7880,N_7117,N_7330);
nand U7881 (N_7881,N_7324,N_7354);
nand U7882 (N_7882,N_7057,N_7096);
nand U7883 (N_7883,N_7058,N_7211);
and U7884 (N_7884,N_7474,N_7191);
or U7885 (N_7885,N_7169,N_7434);
or U7886 (N_7886,N_7340,N_7402);
or U7887 (N_7887,N_7284,N_7425);
nand U7888 (N_7888,N_7168,N_7438);
and U7889 (N_7889,N_7229,N_7267);
and U7890 (N_7890,N_7059,N_7217);
nor U7891 (N_7891,N_7397,N_7313);
and U7892 (N_7892,N_7273,N_7363);
nor U7893 (N_7893,N_7001,N_7193);
or U7894 (N_7894,N_7497,N_7045);
or U7895 (N_7895,N_7076,N_7045);
nand U7896 (N_7896,N_7288,N_7283);
nor U7897 (N_7897,N_7005,N_7495);
xnor U7898 (N_7898,N_7445,N_7222);
and U7899 (N_7899,N_7281,N_7051);
nor U7900 (N_7900,N_7040,N_7481);
and U7901 (N_7901,N_7499,N_7259);
and U7902 (N_7902,N_7181,N_7161);
or U7903 (N_7903,N_7043,N_7307);
nand U7904 (N_7904,N_7035,N_7209);
or U7905 (N_7905,N_7292,N_7304);
nand U7906 (N_7906,N_7457,N_7169);
and U7907 (N_7907,N_7100,N_7061);
and U7908 (N_7908,N_7144,N_7079);
or U7909 (N_7909,N_7096,N_7403);
xnor U7910 (N_7910,N_7444,N_7461);
or U7911 (N_7911,N_7461,N_7010);
or U7912 (N_7912,N_7445,N_7470);
xnor U7913 (N_7913,N_7315,N_7482);
nor U7914 (N_7914,N_7195,N_7411);
xnor U7915 (N_7915,N_7125,N_7491);
nor U7916 (N_7916,N_7084,N_7032);
and U7917 (N_7917,N_7386,N_7404);
nor U7918 (N_7918,N_7015,N_7218);
nand U7919 (N_7919,N_7209,N_7080);
nand U7920 (N_7920,N_7169,N_7454);
or U7921 (N_7921,N_7160,N_7234);
nand U7922 (N_7922,N_7251,N_7294);
nand U7923 (N_7923,N_7193,N_7036);
or U7924 (N_7924,N_7320,N_7385);
nand U7925 (N_7925,N_7205,N_7290);
xnor U7926 (N_7926,N_7283,N_7313);
nand U7927 (N_7927,N_7301,N_7088);
and U7928 (N_7928,N_7019,N_7086);
nor U7929 (N_7929,N_7401,N_7449);
nor U7930 (N_7930,N_7295,N_7107);
and U7931 (N_7931,N_7264,N_7079);
and U7932 (N_7932,N_7187,N_7048);
xnor U7933 (N_7933,N_7061,N_7488);
nor U7934 (N_7934,N_7457,N_7157);
nor U7935 (N_7935,N_7035,N_7310);
xnor U7936 (N_7936,N_7322,N_7360);
nand U7937 (N_7937,N_7083,N_7303);
and U7938 (N_7938,N_7397,N_7194);
or U7939 (N_7939,N_7005,N_7394);
nand U7940 (N_7940,N_7494,N_7072);
nor U7941 (N_7941,N_7203,N_7421);
and U7942 (N_7942,N_7240,N_7478);
nand U7943 (N_7943,N_7129,N_7381);
xor U7944 (N_7944,N_7299,N_7158);
and U7945 (N_7945,N_7204,N_7374);
nand U7946 (N_7946,N_7084,N_7126);
and U7947 (N_7947,N_7064,N_7364);
and U7948 (N_7948,N_7023,N_7169);
or U7949 (N_7949,N_7444,N_7181);
or U7950 (N_7950,N_7270,N_7109);
xor U7951 (N_7951,N_7460,N_7022);
or U7952 (N_7952,N_7364,N_7062);
nor U7953 (N_7953,N_7347,N_7201);
or U7954 (N_7954,N_7333,N_7210);
nor U7955 (N_7955,N_7148,N_7300);
nand U7956 (N_7956,N_7044,N_7322);
xor U7957 (N_7957,N_7414,N_7112);
xnor U7958 (N_7958,N_7297,N_7220);
nor U7959 (N_7959,N_7104,N_7261);
nand U7960 (N_7960,N_7445,N_7449);
nand U7961 (N_7961,N_7452,N_7318);
nor U7962 (N_7962,N_7327,N_7428);
and U7963 (N_7963,N_7156,N_7029);
nand U7964 (N_7964,N_7140,N_7417);
nand U7965 (N_7965,N_7168,N_7371);
and U7966 (N_7966,N_7474,N_7384);
or U7967 (N_7967,N_7155,N_7143);
and U7968 (N_7968,N_7015,N_7084);
and U7969 (N_7969,N_7139,N_7077);
or U7970 (N_7970,N_7462,N_7399);
and U7971 (N_7971,N_7081,N_7406);
nor U7972 (N_7972,N_7341,N_7121);
nor U7973 (N_7973,N_7435,N_7286);
and U7974 (N_7974,N_7333,N_7297);
or U7975 (N_7975,N_7003,N_7465);
and U7976 (N_7976,N_7384,N_7126);
nand U7977 (N_7977,N_7174,N_7045);
or U7978 (N_7978,N_7213,N_7272);
and U7979 (N_7979,N_7129,N_7369);
and U7980 (N_7980,N_7277,N_7421);
nor U7981 (N_7981,N_7213,N_7136);
nand U7982 (N_7982,N_7143,N_7108);
and U7983 (N_7983,N_7009,N_7013);
nor U7984 (N_7984,N_7279,N_7222);
or U7985 (N_7985,N_7297,N_7040);
or U7986 (N_7986,N_7262,N_7245);
or U7987 (N_7987,N_7164,N_7171);
and U7988 (N_7988,N_7296,N_7128);
xnor U7989 (N_7989,N_7064,N_7477);
and U7990 (N_7990,N_7263,N_7023);
nand U7991 (N_7991,N_7262,N_7391);
or U7992 (N_7992,N_7299,N_7114);
or U7993 (N_7993,N_7390,N_7231);
nor U7994 (N_7994,N_7418,N_7332);
nor U7995 (N_7995,N_7163,N_7333);
nor U7996 (N_7996,N_7108,N_7189);
nand U7997 (N_7997,N_7232,N_7127);
nor U7998 (N_7998,N_7132,N_7421);
nor U7999 (N_7999,N_7155,N_7262);
xor U8000 (N_8000,N_7818,N_7769);
nor U8001 (N_8001,N_7837,N_7752);
and U8002 (N_8002,N_7668,N_7646);
xnor U8003 (N_8003,N_7530,N_7636);
or U8004 (N_8004,N_7517,N_7859);
or U8005 (N_8005,N_7892,N_7613);
and U8006 (N_8006,N_7539,N_7969);
nor U8007 (N_8007,N_7504,N_7738);
xor U8008 (N_8008,N_7567,N_7617);
nor U8009 (N_8009,N_7707,N_7755);
and U8010 (N_8010,N_7595,N_7753);
nor U8011 (N_8011,N_7562,N_7697);
or U8012 (N_8012,N_7748,N_7661);
nor U8013 (N_8013,N_7553,N_7700);
and U8014 (N_8014,N_7672,N_7904);
or U8015 (N_8015,N_7704,N_7981);
and U8016 (N_8016,N_7608,N_7566);
or U8017 (N_8017,N_7712,N_7989);
or U8018 (N_8018,N_7946,N_7840);
nor U8019 (N_8019,N_7705,N_7898);
nor U8020 (N_8020,N_7757,N_7764);
and U8021 (N_8021,N_7938,N_7611);
nand U8022 (N_8022,N_7781,N_7895);
and U8023 (N_8023,N_7640,N_7877);
xor U8024 (N_8024,N_7863,N_7586);
or U8025 (N_8025,N_7956,N_7590);
or U8026 (N_8026,N_7835,N_7761);
and U8027 (N_8027,N_7540,N_7819);
nand U8028 (N_8028,N_7552,N_7588);
and U8029 (N_8029,N_7606,N_7524);
nor U8030 (N_8030,N_7512,N_7880);
and U8031 (N_8031,N_7943,N_7772);
xnor U8032 (N_8032,N_7777,N_7831);
nand U8033 (N_8033,N_7711,N_7920);
and U8034 (N_8034,N_7579,N_7839);
nor U8035 (N_8035,N_7805,N_7884);
nor U8036 (N_8036,N_7733,N_7622);
and U8037 (N_8037,N_7670,N_7710);
or U8038 (N_8038,N_7671,N_7536);
and U8039 (N_8039,N_7618,N_7734);
or U8040 (N_8040,N_7885,N_7692);
nor U8041 (N_8041,N_7929,N_7688);
or U8042 (N_8042,N_7997,N_7960);
nand U8043 (N_8043,N_7750,N_7693);
and U8044 (N_8044,N_7996,N_7589);
nand U8045 (N_8045,N_7675,N_7939);
xnor U8046 (N_8046,N_7809,N_7918);
nand U8047 (N_8047,N_7810,N_7975);
nand U8048 (N_8048,N_7703,N_7597);
nor U8049 (N_8049,N_7949,N_7679);
nand U8050 (N_8050,N_7947,N_7650);
nor U8051 (N_8051,N_7667,N_7745);
or U8052 (N_8052,N_7903,N_7771);
and U8053 (N_8053,N_7623,N_7846);
nor U8054 (N_8054,N_7820,N_7842);
xor U8055 (N_8055,N_7888,N_7925);
nor U8056 (N_8056,N_7766,N_7851);
and U8057 (N_8057,N_7602,N_7910);
nand U8058 (N_8058,N_7690,N_7518);
nor U8059 (N_8059,N_7736,N_7922);
or U8060 (N_8060,N_7653,N_7682);
nand U8061 (N_8061,N_7857,N_7627);
and U8062 (N_8062,N_7853,N_7545);
nand U8063 (N_8063,N_7974,N_7765);
or U8064 (N_8064,N_7987,N_7541);
nand U8065 (N_8065,N_7980,N_7911);
or U8066 (N_8066,N_7629,N_7847);
nand U8067 (N_8067,N_7855,N_7502);
nor U8068 (N_8068,N_7645,N_7664);
xnor U8069 (N_8069,N_7551,N_7506);
nand U8070 (N_8070,N_7596,N_7882);
and U8071 (N_8071,N_7767,N_7575);
nand U8072 (N_8072,N_7612,N_7585);
and U8073 (N_8073,N_7547,N_7897);
xnor U8074 (N_8074,N_7988,N_7601);
nand U8075 (N_8075,N_7937,N_7580);
and U8076 (N_8076,N_7744,N_7890);
or U8077 (N_8077,N_7919,N_7564);
nor U8078 (N_8078,N_7559,N_7715);
or U8079 (N_8079,N_7511,N_7599);
nand U8080 (N_8080,N_7637,N_7544);
nor U8081 (N_8081,N_7827,N_7543);
and U8082 (N_8082,N_7515,N_7525);
and U8083 (N_8083,N_7604,N_7776);
nor U8084 (N_8084,N_7639,N_7724);
nor U8085 (N_8085,N_7737,N_7731);
or U8086 (N_8086,N_7786,N_7647);
and U8087 (N_8087,N_7955,N_7548);
nor U8088 (N_8088,N_7915,N_7649);
xnor U8089 (N_8089,N_7965,N_7702);
and U8090 (N_8090,N_7906,N_7933);
xnor U8091 (N_8091,N_7509,N_7659);
and U8092 (N_8092,N_7522,N_7728);
nor U8093 (N_8093,N_7948,N_7773);
and U8094 (N_8094,N_7534,N_7811);
or U8095 (N_8095,N_7924,N_7665);
nand U8096 (N_8096,N_7778,N_7538);
nand U8097 (N_8097,N_7790,N_7560);
and U8098 (N_8098,N_7982,N_7964);
nor U8099 (N_8099,N_7749,N_7725);
xnor U8100 (N_8100,N_7620,N_7740);
or U8101 (N_8101,N_7927,N_7869);
and U8102 (N_8102,N_7814,N_7626);
and U8103 (N_8103,N_7901,N_7878);
nand U8104 (N_8104,N_7625,N_7848);
xor U8105 (N_8105,N_7967,N_7716);
xnor U8106 (N_8106,N_7881,N_7691);
nor U8107 (N_8107,N_7813,N_7834);
or U8108 (N_8108,N_7662,N_7935);
and U8109 (N_8109,N_7568,N_7991);
or U8110 (N_8110,N_7833,N_7746);
and U8111 (N_8111,N_7642,N_7758);
or U8112 (N_8112,N_7843,N_7526);
and U8113 (N_8113,N_7998,N_7628);
nor U8114 (N_8114,N_7598,N_7887);
and U8115 (N_8115,N_7985,N_7689);
nor U8116 (N_8116,N_7963,N_7858);
nand U8117 (N_8117,N_7576,N_7673);
nand U8118 (N_8118,N_7574,N_7635);
xor U8119 (N_8119,N_7713,N_7799);
or U8120 (N_8120,N_7591,N_7905);
nand U8121 (N_8121,N_7829,N_7708);
or U8122 (N_8122,N_7782,N_7936);
nand U8123 (N_8123,N_7893,N_7763);
and U8124 (N_8124,N_7654,N_7958);
xnor U8125 (N_8125,N_7909,N_7593);
and U8126 (N_8126,N_7605,N_7867);
and U8127 (N_8127,N_7961,N_7794);
nor U8128 (N_8128,N_7886,N_7729);
and U8129 (N_8129,N_7774,N_7584);
nand U8130 (N_8130,N_7950,N_7743);
nor U8131 (N_8131,N_7862,N_7587);
or U8132 (N_8132,N_7614,N_7816);
nor U8133 (N_8133,N_7876,N_7594);
xor U8134 (N_8134,N_7563,N_7683);
nor U8135 (N_8135,N_7657,N_7795);
nor U8136 (N_8136,N_7796,N_7986);
xnor U8137 (N_8137,N_7521,N_7788);
nor U8138 (N_8138,N_7959,N_7875);
xnor U8139 (N_8139,N_7742,N_7609);
nor U8140 (N_8140,N_7621,N_7792);
or U8141 (N_8141,N_7825,N_7994);
nor U8142 (N_8142,N_7945,N_7550);
and U8143 (N_8143,N_7694,N_7872);
nand U8144 (N_8144,N_7503,N_7808);
xnor U8145 (N_8145,N_7633,N_7505);
and U8146 (N_8146,N_7630,N_7709);
and U8147 (N_8147,N_7644,N_7856);
and U8148 (N_8148,N_7874,N_7870);
nand U8149 (N_8149,N_7804,N_7658);
and U8150 (N_8150,N_7523,N_7891);
nor U8151 (N_8151,N_7554,N_7983);
nor U8152 (N_8152,N_7914,N_7921);
nor U8153 (N_8153,N_7720,N_7836);
nor U8154 (N_8154,N_7930,N_7812);
and U8155 (N_8155,N_7569,N_7826);
and U8156 (N_8156,N_7896,N_7865);
nor U8157 (N_8157,N_7984,N_7600);
nor U8158 (N_8158,N_7655,N_7527);
and U8159 (N_8159,N_7718,N_7531);
nor U8160 (N_8160,N_7751,N_7696);
and U8161 (N_8161,N_7784,N_7864);
nand U8162 (N_8162,N_7666,N_7756);
nor U8163 (N_8163,N_7684,N_7850);
or U8164 (N_8164,N_7638,N_7535);
nor U8165 (N_8165,N_7676,N_7581);
and U8166 (N_8166,N_7508,N_7970);
and U8167 (N_8167,N_7557,N_7678);
nand U8168 (N_8168,N_7706,N_7634);
and U8169 (N_8169,N_7873,N_7866);
and U8170 (N_8170,N_7762,N_7780);
nor U8171 (N_8171,N_7723,N_7501);
and U8172 (N_8172,N_7695,N_7516);
and U8173 (N_8173,N_7942,N_7681);
and U8174 (N_8174,N_7565,N_7747);
and U8175 (N_8175,N_7871,N_7815);
nor U8176 (N_8176,N_7643,N_7912);
nand U8177 (N_8177,N_7685,N_7582);
nand U8178 (N_8178,N_7783,N_7656);
or U8179 (N_8179,N_7972,N_7714);
and U8180 (N_8180,N_7923,N_7717);
and U8181 (N_8181,N_7926,N_7798);
or U8182 (N_8182,N_7732,N_7768);
or U8183 (N_8183,N_7971,N_7507);
and U8184 (N_8184,N_7760,N_7993);
nor U8185 (N_8185,N_7698,N_7849);
nand U8186 (N_8186,N_7779,N_7883);
or U8187 (N_8187,N_7889,N_7616);
nor U8188 (N_8188,N_7828,N_7879);
nor U8189 (N_8189,N_7759,N_7868);
xor U8190 (N_8190,N_7838,N_7916);
and U8191 (N_8191,N_7932,N_7739);
nor U8192 (N_8192,N_7941,N_7861);
or U8193 (N_8193,N_7944,N_7894);
xor U8194 (N_8194,N_7513,N_7735);
nor U8195 (N_8195,N_7529,N_7677);
nand U8196 (N_8196,N_7555,N_7913);
xnor U8197 (N_8197,N_7561,N_7632);
or U8198 (N_8198,N_7854,N_7660);
or U8199 (N_8199,N_7519,N_7844);
xnor U8200 (N_8200,N_7860,N_7577);
and U8201 (N_8201,N_7823,N_7770);
and U8202 (N_8202,N_7510,N_7979);
or U8203 (N_8203,N_7954,N_7992);
nor U8204 (N_8204,N_7607,N_7680);
nand U8205 (N_8205,N_7730,N_7821);
and U8206 (N_8206,N_7801,N_7537);
nor U8207 (N_8207,N_7726,N_7940);
nor U8208 (N_8208,N_7570,N_7727);
nand U8209 (N_8209,N_7977,N_7789);
nand U8210 (N_8210,N_7631,N_7845);
nand U8211 (N_8211,N_7800,N_7663);
or U8212 (N_8212,N_7990,N_7907);
nor U8213 (N_8213,N_7719,N_7546);
or U8214 (N_8214,N_7999,N_7520);
or U8215 (N_8215,N_7651,N_7934);
or U8216 (N_8216,N_7830,N_7686);
or U8217 (N_8217,N_7533,N_7900);
xnor U8218 (N_8218,N_7841,N_7573);
xor U8219 (N_8219,N_7558,N_7592);
nand U8220 (N_8220,N_7931,N_7951);
or U8221 (N_8221,N_7791,N_7785);
nor U8222 (N_8222,N_7978,N_7803);
xor U8223 (N_8223,N_7962,N_7674);
or U8224 (N_8224,N_7775,N_7556);
nand U8225 (N_8225,N_7701,N_7583);
and U8226 (N_8226,N_7572,N_7669);
nand U8227 (N_8227,N_7817,N_7802);
nor U8228 (N_8228,N_7852,N_7754);
or U8229 (N_8229,N_7957,N_7952);
nand U8230 (N_8230,N_7549,N_7652);
nand U8231 (N_8231,N_7571,N_7741);
nand U8232 (N_8232,N_7603,N_7902);
or U8233 (N_8233,N_7953,N_7722);
or U8234 (N_8234,N_7793,N_7532);
and U8235 (N_8235,N_7615,N_7721);
xnor U8236 (N_8236,N_7807,N_7797);
and U8237 (N_8237,N_7610,N_7806);
and U8238 (N_8238,N_7624,N_7917);
nor U8239 (N_8239,N_7787,N_7968);
nand U8240 (N_8240,N_7976,N_7699);
nor U8241 (N_8241,N_7908,N_7899);
nor U8242 (N_8242,N_7648,N_7973);
or U8243 (N_8243,N_7514,N_7832);
nand U8244 (N_8244,N_7928,N_7822);
and U8245 (N_8245,N_7500,N_7578);
or U8246 (N_8246,N_7528,N_7824);
or U8247 (N_8247,N_7542,N_7619);
nor U8248 (N_8248,N_7966,N_7641);
xor U8249 (N_8249,N_7995,N_7687);
or U8250 (N_8250,N_7785,N_7824);
and U8251 (N_8251,N_7567,N_7644);
or U8252 (N_8252,N_7860,N_7576);
nand U8253 (N_8253,N_7858,N_7880);
and U8254 (N_8254,N_7648,N_7786);
xnor U8255 (N_8255,N_7723,N_7812);
nand U8256 (N_8256,N_7981,N_7653);
or U8257 (N_8257,N_7853,N_7985);
and U8258 (N_8258,N_7668,N_7876);
or U8259 (N_8259,N_7736,N_7645);
nand U8260 (N_8260,N_7577,N_7887);
nand U8261 (N_8261,N_7576,N_7827);
or U8262 (N_8262,N_7835,N_7886);
or U8263 (N_8263,N_7776,N_7778);
nor U8264 (N_8264,N_7757,N_7815);
nor U8265 (N_8265,N_7705,N_7947);
or U8266 (N_8266,N_7572,N_7882);
and U8267 (N_8267,N_7563,N_7984);
nor U8268 (N_8268,N_7528,N_7947);
and U8269 (N_8269,N_7598,N_7869);
or U8270 (N_8270,N_7948,N_7660);
nor U8271 (N_8271,N_7968,N_7821);
or U8272 (N_8272,N_7617,N_7591);
nor U8273 (N_8273,N_7619,N_7898);
and U8274 (N_8274,N_7774,N_7659);
and U8275 (N_8275,N_7716,N_7833);
nor U8276 (N_8276,N_7719,N_7834);
nand U8277 (N_8277,N_7677,N_7688);
nand U8278 (N_8278,N_7717,N_7995);
nand U8279 (N_8279,N_7511,N_7655);
nor U8280 (N_8280,N_7852,N_7648);
or U8281 (N_8281,N_7854,N_7585);
and U8282 (N_8282,N_7928,N_7598);
and U8283 (N_8283,N_7581,N_7635);
and U8284 (N_8284,N_7908,N_7795);
or U8285 (N_8285,N_7610,N_7800);
nand U8286 (N_8286,N_7900,N_7681);
nand U8287 (N_8287,N_7661,N_7699);
xor U8288 (N_8288,N_7529,N_7682);
nand U8289 (N_8289,N_7887,N_7939);
and U8290 (N_8290,N_7511,N_7906);
or U8291 (N_8291,N_7718,N_7925);
or U8292 (N_8292,N_7690,N_7576);
and U8293 (N_8293,N_7914,N_7684);
or U8294 (N_8294,N_7878,N_7829);
nand U8295 (N_8295,N_7760,N_7604);
nand U8296 (N_8296,N_7615,N_7654);
and U8297 (N_8297,N_7981,N_7707);
nand U8298 (N_8298,N_7718,N_7714);
and U8299 (N_8299,N_7744,N_7915);
nand U8300 (N_8300,N_7675,N_7839);
and U8301 (N_8301,N_7986,N_7693);
and U8302 (N_8302,N_7859,N_7588);
or U8303 (N_8303,N_7876,N_7752);
nor U8304 (N_8304,N_7879,N_7808);
nand U8305 (N_8305,N_7992,N_7819);
nand U8306 (N_8306,N_7803,N_7576);
nor U8307 (N_8307,N_7671,N_7585);
nand U8308 (N_8308,N_7554,N_7888);
nand U8309 (N_8309,N_7974,N_7799);
nor U8310 (N_8310,N_7566,N_7976);
or U8311 (N_8311,N_7590,N_7731);
xor U8312 (N_8312,N_7599,N_7527);
nand U8313 (N_8313,N_7558,N_7604);
xor U8314 (N_8314,N_7894,N_7608);
and U8315 (N_8315,N_7738,N_7861);
nand U8316 (N_8316,N_7925,N_7941);
or U8317 (N_8317,N_7793,N_7895);
and U8318 (N_8318,N_7733,N_7512);
xnor U8319 (N_8319,N_7809,N_7776);
nor U8320 (N_8320,N_7871,N_7713);
nor U8321 (N_8321,N_7643,N_7928);
or U8322 (N_8322,N_7770,N_7627);
nor U8323 (N_8323,N_7619,N_7746);
nand U8324 (N_8324,N_7743,N_7580);
or U8325 (N_8325,N_7614,N_7883);
nor U8326 (N_8326,N_7685,N_7859);
or U8327 (N_8327,N_7693,N_7926);
and U8328 (N_8328,N_7565,N_7810);
nand U8329 (N_8329,N_7722,N_7934);
nor U8330 (N_8330,N_7903,N_7557);
nand U8331 (N_8331,N_7529,N_7543);
nor U8332 (N_8332,N_7899,N_7830);
nor U8333 (N_8333,N_7612,N_7726);
and U8334 (N_8334,N_7582,N_7946);
nand U8335 (N_8335,N_7517,N_7796);
nor U8336 (N_8336,N_7823,N_7930);
and U8337 (N_8337,N_7669,N_7741);
and U8338 (N_8338,N_7765,N_7712);
nand U8339 (N_8339,N_7619,N_7710);
and U8340 (N_8340,N_7679,N_7960);
or U8341 (N_8341,N_7672,N_7759);
nand U8342 (N_8342,N_7666,N_7986);
nand U8343 (N_8343,N_7898,N_7732);
nand U8344 (N_8344,N_7625,N_7795);
nand U8345 (N_8345,N_7594,N_7854);
and U8346 (N_8346,N_7669,N_7853);
nand U8347 (N_8347,N_7789,N_7918);
nor U8348 (N_8348,N_7924,N_7786);
nand U8349 (N_8349,N_7738,N_7804);
nand U8350 (N_8350,N_7626,N_7887);
nor U8351 (N_8351,N_7677,N_7994);
and U8352 (N_8352,N_7607,N_7867);
nand U8353 (N_8353,N_7771,N_7512);
or U8354 (N_8354,N_7630,N_7696);
nor U8355 (N_8355,N_7892,N_7915);
xor U8356 (N_8356,N_7805,N_7730);
and U8357 (N_8357,N_7931,N_7884);
nand U8358 (N_8358,N_7583,N_7990);
nand U8359 (N_8359,N_7570,N_7613);
nor U8360 (N_8360,N_7661,N_7923);
or U8361 (N_8361,N_7722,N_7854);
or U8362 (N_8362,N_7693,N_7974);
nor U8363 (N_8363,N_7967,N_7650);
xnor U8364 (N_8364,N_7568,N_7736);
nand U8365 (N_8365,N_7725,N_7516);
or U8366 (N_8366,N_7510,N_7895);
or U8367 (N_8367,N_7720,N_7527);
nand U8368 (N_8368,N_7868,N_7943);
nand U8369 (N_8369,N_7946,N_7821);
and U8370 (N_8370,N_7961,N_7689);
nand U8371 (N_8371,N_7859,N_7789);
xor U8372 (N_8372,N_7895,N_7971);
xnor U8373 (N_8373,N_7826,N_7654);
nand U8374 (N_8374,N_7913,N_7568);
nand U8375 (N_8375,N_7671,N_7603);
or U8376 (N_8376,N_7516,N_7618);
nand U8377 (N_8377,N_7961,N_7869);
nor U8378 (N_8378,N_7691,N_7722);
or U8379 (N_8379,N_7687,N_7532);
and U8380 (N_8380,N_7859,N_7814);
nand U8381 (N_8381,N_7968,N_7560);
or U8382 (N_8382,N_7577,N_7726);
or U8383 (N_8383,N_7626,N_7631);
and U8384 (N_8384,N_7729,N_7980);
or U8385 (N_8385,N_7822,N_7596);
and U8386 (N_8386,N_7953,N_7968);
nor U8387 (N_8387,N_7596,N_7752);
and U8388 (N_8388,N_7993,N_7871);
and U8389 (N_8389,N_7971,N_7811);
nand U8390 (N_8390,N_7761,N_7940);
nand U8391 (N_8391,N_7830,N_7979);
and U8392 (N_8392,N_7944,N_7950);
or U8393 (N_8393,N_7528,N_7842);
or U8394 (N_8394,N_7628,N_7743);
nor U8395 (N_8395,N_7504,N_7897);
nor U8396 (N_8396,N_7725,N_7845);
nor U8397 (N_8397,N_7540,N_7984);
nor U8398 (N_8398,N_7718,N_7923);
and U8399 (N_8399,N_7995,N_7641);
or U8400 (N_8400,N_7933,N_7617);
and U8401 (N_8401,N_7575,N_7932);
and U8402 (N_8402,N_7767,N_7853);
nor U8403 (N_8403,N_7835,N_7704);
and U8404 (N_8404,N_7921,N_7845);
or U8405 (N_8405,N_7897,N_7551);
or U8406 (N_8406,N_7718,N_7813);
or U8407 (N_8407,N_7542,N_7755);
and U8408 (N_8408,N_7798,N_7773);
nand U8409 (N_8409,N_7708,N_7585);
nor U8410 (N_8410,N_7730,N_7741);
or U8411 (N_8411,N_7976,N_7597);
nor U8412 (N_8412,N_7929,N_7787);
and U8413 (N_8413,N_7542,N_7538);
and U8414 (N_8414,N_7963,N_7548);
or U8415 (N_8415,N_7842,N_7909);
xnor U8416 (N_8416,N_7673,N_7594);
or U8417 (N_8417,N_7800,N_7964);
nand U8418 (N_8418,N_7594,N_7910);
nor U8419 (N_8419,N_7767,N_7677);
xnor U8420 (N_8420,N_7953,N_7808);
or U8421 (N_8421,N_7642,N_7968);
or U8422 (N_8422,N_7788,N_7537);
nor U8423 (N_8423,N_7715,N_7518);
and U8424 (N_8424,N_7820,N_7645);
and U8425 (N_8425,N_7637,N_7990);
or U8426 (N_8426,N_7730,N_7508);
nor U8427 (N_8427,N_7908,N_7780);
nand U8428 (N_8428,N_7893,N_7582);
and U8429 (N_8429,N_7686,N_7647);
nand U8430 (N_8430,N_7625,N_7727);
nor U8431 (N_8431,N_7566,N_7573);
xnor U8432 (N_8432,N_7810,N_7660);
and U8433 (N_8433,N_7643,N_7836);
nor U8434 (N_8434,N_7898,N_7865);
nor U8435 (N_8435,N_7794,N_7806);
nor U8436 (N_8436,N_7672,N_7886);
and U8437 (N_8437,N_7867,N_7557);
nor U8438 (N_8438,N_7709,N_7702);
and U8439 (N_8439,N_7691,N_7540);
nor U8440 (N_8440,N_7849,N_7701);
nor U8441 (N_8441,N_7762,N_7991);
nand U8442 (N_8442,N_7753,N_7712);
and U8443 (N_8443,N_7819,N_7705);
and U8444 (N_8444,N_7830,N_7887);
nand U8445 (N_8445,N_7788,N_7911);
nor U8446 (N_8446,N_7909,N_7559);
or U8447 (N_8447,N_7905,N_7793);
and U8448 (N_8448,N_7630,N_7576);
or U8449 (N_8449,N_7843,N_7716);
nor U8450 (N_8450,N_7696,N_7814);
nor U8451 (N_8451,N_7952,N_7552);
and U8452 (N_8452,N_7904,N_7859);
or U8453 (N_8453,N_7630,N_7974);
or U8454 (N_8454,N_7727,N_7809);
nor U8455 (N_8455,N_7766,N_7938);
nor U8456 (N_8456,N_7690,N_7712);
and U8457 (N_8457,N_7558,N_7784);
nor U8458 (N_8458,N_7527,N_7744);
xor U8459 (N_8459,N_7511,N_7652);
and U8460 (N_8460,N_7973,N_7620);
and U8461 (N_8461,N_7541,N_7991);
xnor U8462 (N_8462,N_7997,N_7900);
nor U8463 (N_8463,N_7560,N_7835);
or U8464 (N_8464,N_7651,N_7890);
nand U8465 (N_8465,N_7790,N_7651);
nor U8466 (N_8466,N_7736,N_7702);
and U8467 (N_8467,N_7553,N_7851);
or U8468 (N_8468,N_7588,N_7918);
nor U8469 (N_8469,N_7961,N_7548);
nor U8470 (N_8470,N_7720,N_7844);
nand U8471 (N_8471,N_7974,N_7729);
nand U8472 (N_8472,N_7780,N_7735);
nor U8473 (N_8473,N_7505,N_7907);
or U8474 (N_8474,N_7916,N_7516);
nand U8475 (N_8475,N_7964,N_7892);
or U8476 (N_8476,N_7958,N_7868);
or U8477 (N_8477,N_7548,N_7641);
and U8478 (N_8478,N_7639,N_7845);
nand U8479 (N_8479,N_7696,N_7938);
nor U8480 (N_8480,N_7636,N_7761);
and U8481 (N_8481,N_7959,N_7840);
nor U8482 (N_8482,N_7585,N_7579);
or U8483 (N_8483,N_7727,N_7691);
nor U8484 (N_8484,N_7939,N_7972);
nor U8485 (N_8485,N_7997,N_7849);
nor U8486 (N_8486,N_7832,N_7987);
or U8487 (N_8487,N_7509,N_7709);
and U8488 (N_8488,N_7967,N_7808);
nor U8489 (N_8489,N_7839,N_7789);
or U8490 (N_8490,N_7873,N_7590);
or U8491 (N_8491,N_7695,N_7791);
nor U8492 (N_8492,N_7567,N_7564);
and U8493 (N_8493,N_7797,N_7554);
or U8494 (N_8494,N_7681,N_7731);
and U8495 (N_8495,N_7875,N_7544);
nand U8496 (N_8496,N_7506,N_7951);
and U8497 (N_8497,N_7766,N_7538);
nand U8498 (N_8498,N_7908,N_7562);
nor U8499 (N_8499,N_7679,N_7895);
and U8500 (N_8500,N_8359,N_8183);
nor U8501 (N_8501,N_8103,N_8019);
nand U8502 (N_8502,N_8277,N_8199);
or U8503 (N_8503,N_8222,N_8257);
and U8504 (N_8504,N_8050,N_8329);
nand U8505 (N_8505,N_8098,N_8068);
or U8506 (N_8506,N_8356,N_8353);
nand U8507 (N_8507,N_8201,N_8399);
and U8508 (N_8508,N_8345,N_8185);
nand U8509 (N_8509,N_8247,N_8173);
nor U8510 (N_8510,N_8436,N_8351);
or U8511 (N_8511,N_8018,N_8271);
nand U8512 (N_8512,N_8057,N_8147);
nand U8513 (N_8513,N_8381,N_8390);
nor U8514 (N_8514,N_8287,N_8422);
or U8515 (N_8515,N_8358,N_8062);
and U8516 (N_8516,N_8022,N_8065);
or U8517 (N_8517,N_8090,N_8442);
nor U8518 (N_8518,N_8140,N_8413);
and U8519 (N_8519,N_8301,N_8216);
or U8520 (N_8520,N_8434,N_8258);
and U8521 (N_8521,N_8094,N_8034);
or U8522 (N_8522,N_8272,N_8417);
or U8523 (N_8523,N_8451,N_8058);
nand U8524 (N_8524,N_8446,N_8273);
or U8525 (N_8525,N_8200,N_8328);
nor U8526 (N_8526,N_8129,N_8340);
or U8527 (N_8527,N_8212,N_8276);
nand U8528 (N_8528,N_8264,N_8189);
or U8529 (N_8529,N_8056,N_8380);
nor U8530 (N_8530,N_8071,N_8223);
nor U8531 (N_8531,N_8024,N_8453);
xor U8532 (N_8532,N_8484,N_8220);
and U8533 (N_8533,N_8360,N_8291);
and U8534 (N_8534,N_8467,N_8218);
nand U8535 (N_8535,N_8414,N_8032);
or U8536 (N_8536,N_8424,N_8375);
or U8537 (N_8537,N_8260,N_8089);
xnor U8538 (N_8538,N_8312,N_8289);
nand U8539 (N_8539,N_8462,N_8474);
or U8540 (N_8540,N_8343,N_8181);
or U8541 (N_8541,N_8002,N_8014);
nand U8542 (N_8542,N_8163,N_8315);
or U8543 (N_8543,N_8118,N_8154);
or U8544 (N_8544,N_8388,N_8338);
or U8545 (N_8545,N_8197,N_8466);
nor U8546 (N_8546,N_8003,N_8204);
or U8547 (N_8547,N_8254,N_8054);
xnor U8548 (N_8548,N_8464,N_8443);
xnor U8549 (N_8549,N_8231,N_8447);
and U8550 (N_8550,N_8468,N_8198);
or U8551 (N_8551,N_8108,N_8037);
and U8552 (N_8552,N_8490,N_8136);
xnor U8553 (N_8553,N_8366,N_8342);
xnor U8554 (N_8554,N_8431,N_8040);
nor U8555 (N_8555,N_8428,N_8126);
nand U8556 (N_8556,N_8396,N_8421);
nor U8557 (N_8557,N_8455,N_8176);
nand U8558 (N_8558,N_8210,N_8405);
nor U8559 (N_8559,N_8155,N_8426);
nand U8560 (N_8560,N_8076,N_8371);
nor U8561 (N_8561,N_8393,N_8263);
and U8562 (N_8562,N_8365,N_8344);
nor U8563 (N_8563,N_8109,N_8233);
nor U8564 (N_8564,N_8027,N_8498);
xor U8565 (N_8565,N_8253,N_8295);
and U8566 (N_8566,N_8265,N_8234);
and U8567 (N_8567,N_8317,N_8191);
nand U8568 (N_8568,N_8377,N_8382);
nand U8569 (N_8569,N_8493,N_8452);
and U8570 (N_8570,N_8100,N_8293);
and U8571 (N_8571,N_8217,N_8239);
or U8572 (N_8572,N_8385,N_8142);
nand U8573 (N_8573,N_8488,N_8111);
nor U8574 (N_8574,N_8232,N_8167);
nor U8575 (N_8575,N_8363,N_8458);
and U8576 (N_8576,N_8309,N_8159);
xnor U8577 (N_8577,N_8114,N_8066);
or U8578 (N_8578,N_8046,N_8006);
nor U8579 (N_8579,N_8193,N_8336);
xor U8580 (N_8580,N_8143,N_8456);
and U8581 (N_8581,N_8269,N_8406);
nand U8582 (N_8582,N_8387,N_8262);
nor U8583 (N_8583,N_8115,N_8367);
and U8584 (N_8584,N_8093,N_8207);
xnor U8585 (N_8585,N_8157,N_8499);
or U8586 (N_8586,N_8407,N_8482);
xor U8587 (N_8587,N_8383,N_8087);
nor U8588 (N_8588,N_8224,N_8012);
or U8589 (N_8589,N_8320,N_8432);
and U8590 (N_8590,N_8410,N_8379);
nand U8591 (N_8591,N_8300,N_8331);
or U8592 (N_8592,N_8042,N_8245);
or U8593 (N_8593,N_8226,N_8290);
nand U8594 (N_8594,N_8180,N_8445);
nor U8595 (N_8595,N_8106,N_8337);
and U8596 (N_8596,N_8013,N_8025);
and U8597 (N_8597,N_8319,N_8074);
nor U8598 (N_8598,N_8495,N_8011);
or U8599 (N_8599,N_8242,N_8280);
nand U8600 (N_8600,N_8316,N_8252);
nor U8601 (N_8601,N_8404,N_8435);
or U8602 (N_8602,N_8374,N_8219);
or U8603 (N_8603,N_8369,N_8270);
xor U8604 (N_8604,N_8151,N_8203);
or U8605 (N_8605,N_8261,N_8292);
or U8606 (N_8606,N_8297,N_8459);
or U8607 (N_8607,N_8333,N_8010);
and U8608 (N_8608,N_8067,N_8267);
nand U8609 (N_8609,N_8225,N_8251);
nor U8610 (N_8610,N_8036,N_8469);
and U8611 (N_8611,N_8243,N_8208);
and U8612 (N_8612,N_8250,N_8279);
nand U8613 (N_8613,N_8281,N_8070);
nor U8614 (N_8614,N_8470,N_8069);
and U8615 (N_8615,N_8408,N_8177);
and U8616 (N_8616,N_8327,N_8081);
or U8617 (N_8617,N_8454,N_8196);
or U8618 (N_8618,N_8433,N_8349);
and U8619 (N_8619,N_8427,N_8480);
and U8620 (N_8620,N_8078,N_8105);
nand U8621 (N_8621,N_8368,N_8357);
nand U8622 (N_8622,N_8248,N_8412);
nand U8623 (N_8623,N_8102,N_8423);
xnor U8624 (N_8624,N_8008,N_8373);
nor U8625 (N_8625,N_8313,N_8079);
nor U8626 (N_8626,N_8122,N_8311);
and U8627 (N_8627,N_8121,N_8481);
nor U8628 (N_8628,N_8494,N_8130);
nor U8629 (N_8629,N_8119,N_8463);
nor U8630 (N_8630,N_8080,N_8268);
nor U8631 (N_8631,N_8170,N_8370);
and U8632 (N_8632,N_8274,N_8063);
nor U8633 (N_8633,N_8348,N_8175);
nand U8634 (N_8634,N_8400,N_8401);
nor U8635 (N_8635,N_8149,N_8128);
or U8636 (N_8636,N_8487,N_8064);
nand U8637 (N_8637,N_8020,N_8088);
and U8638 (N_8638,N_8148,N_8117);
nor U8639 (N_8639,N_8449,N_8075);
and U8640 (N_8640,N_8214,N_8409);
nand U8641 (N_8641,N_8391,N_8285);
xor U8642 (N_8642,N_8097,N_8429);
nand U8643 (N_8643,N_8240,N_8361);
nand U8644 (N_8644,N_8236,N_8047);
nand U8645 (N_8645,N_8486,N_8221);
nor U8646 (N_8646,N_8384,N_8376);
xnor U8647 (N_8647,N_8060,N_8153);
xnor U8648 (N_8648,N_8237,N_8282);
xnor U8649 (N_8649,N_8448,N_8158);
or U8650 (N_8650,N_8127,N_8321);
or U8651 (N_8651,N_8015,N_8294);
or U8652 (N_8652,N_8402,N_8308);
nand U8653 (N_8653,N_8135,N_8156);
and U8654 (N_8654,N_8113,N_8160);
nand U8655 (N_8655,N_8283,N_8112);
or U8656 (N_8656,N_8033,N_8322);
nand U8657 (N_8657,N_8346,N_8187);
nor U8658 (N_8658,N_8403,N_8195);
or U8659 (N_8659,N_8278,N_8029);
xor U8660 (N_8660,N_8241,N_8205);
nor U8661 (N_8661,N_8229,N_8305);
nor U8662 (N_8662,N_8139,N_8465);
nor U8663 (N_8663,N_8473,N_8096);
xor U8664 (N_8664,N_8324,N_8497);
nor U8665 (N_8665,N_8124,N_8141);
nor U8666 (N_8666,N_8182,N_8031);
and U8667 (N_8667,N_8004,N_8364);
nand U8668 (N_8668,N_8132,N_8202);
or U8669 (N_8669,N_8303,N_8419);
nor U8670 (N_8670,N_8171,N_8168);
and U8671 (N_8671,N_8394,N_8044);
nor U8672 (N_8672,N_8386,N_8162);
nand U8673 (N_8673,N_8211,N_8150);
nor U8674 (N_8674,N_8209,N_8492);
nor U8675 (N_8675,N_8352,N_8334);
xor U8676 (N_8676,N_8039,N_8026);
and U8677 (N_8677,N_8137,N_8298);
and U8678 (N_8678,N_8179,N_8005);
or U8679 (N_8679,N_8304,N_8145);
or U8680 (N_8680,N_8471,N_8444);
nor U8681 (N_8681,N_8489,N_8347);
and U8682 (N_8682,N_8341,N_8073);
nor U8683 (N_8683,N_8415,N_8460);
nor U8684 (N_8684,N_8227,N_8169);
or U8685 (N_8685,N_8190,N_8104);
and U8686 (N_8686,N_8086,N_8284);
nand U8687 (N_8687,N_8131,N_8450);
xnor U8688 (N_8688,N_8302,N_8049);
xor U8689 (N_8689,N_8318,N_8418);
nor U8690 (N_8690,N_8330,N_8152);
nor U8691 (N_8691,N_8496,N_8244);
or U8692 (N_8692,N_8275,N_8085);
or U8693 (N_8693,N_8246,N_8256);
nor U8694 (N_8694,N_8165,N_8335);
xnor U8695 (N_8695,N_8192,N_8082);
nor U8696 (N_8696,N_8332,N_8099);
or U8697 (N_8697,N_8215,N_8372);
and U8698 (N_8698,N_8146,N_8072);
xor U8699 (N_8699,N_8043,N_8016);
nand U8700 (N_8700,N_8310,N_8084);
nor U8701 (N_8701,N_8411,N_8041);
and U8702 (N_8702,N_8007,N_8000);
and U8703 (N_8703,N_8172,N_8048);
nand U8704 (N_8704,N_8440,N_8350);
nor U8705 (N_8705,N_8472,N_8116);
and U8706 (N_8706,N_8306,N_8051);
xnor U8707 (N_8707,N_8420,N_8323);
nand U8708 (N_8708,N_8389,N_8266);
nand U8709 (N_8709,N_8476,N_8138);
nor U8710 (N_8710,N_8174,N_8475);
and U8711 (N_8711,N_8091,N_8430);
xor U8712 (N_8712,N_8101,N_8144);
or U8713 (N_8713,N_8438,N_8194);
nand U8714 (N_8714,N_8178,N_8230);
nor U8715 (N_8715,N_8299,N_8249);
nand U8716 (N_8716,N_8397,N_8314);
nand U8717 (N_8717,N_8123,N_8477);
or U8718 (N_8718,N_8030,N_8095);
nand U8719 (N_8719,N_8120,N_8255);
nor U8720 (N_8720,N_8441,N_8259);
or U8721 (N_8721,N_8296,N_8398);
nand U8722 (N_8722,N_8134,N_8061);
nor U8723 (N_8723,N_8362,N_8083);
nor U8724 (N_8724,N_8326,N_8038);
xnor U8725 (N_8725,N_8288,N_8478);
or U8726 (N_8726,N_8107,N_8001);
and U8727 (N_8727,N_8483,N_8021);
nor U8728 (N_8728,N_8009,N_8354);
and U8729 (N_8729,N_8184,N_8028);
or U8730 (N_8730,N_8166,N_8395);
and U8731 (N_8731,N_8213,N_8059);
nor U8732 (N_8732,N_8161,N_8235);
and U8733 (N_8733,N_8206,N_8017);
and U8734 (N_8734,N_8439,N_8491);
nor U8735 (N_8735,N_8055,N_8392);
or U8736 (N_8736,N_8307,N_8355);
and U8737 (N_8737,N_8485,N_8425);
and U8738 (N_8738,N_8164,N_8437);
nand U8739 (N_8739,N_8052,N_8053);
nor U8740 (N_8740,N_8457,N_8077);
or U8741 (N_8741,N_8416,N_8023);
nand U8742 (N_8742,N_8325,N_8092);
nor U8743 (N_8743,N_8045,N_8461);
nor U8744 (N_8744,N_8110,N_8133);
nor U8745 (N_8745,N_8479,N_8035);
nand U8746 (N_8746,N_8186,N_8286);
xnor U8747 (N_8747,N_8188,N_8238);
nand U8748 (N_8748,N_8339,N_8378);
nor U8749 (N_8749,N_8125,N_8228);
nand U8750 (N_8750,N_8465,N_8385);
and U8751 (N_8751,N_8351,N_8202);
or U8752 (N_8752,N_8182,N_8396);
nand U8753 (N_8753,N_8311,N_8492);
or U8754 (N_8754,N_8227,N_8251);
or U8755 (N_8755,N_8412,N_8474);
xnor U8756 (N_8756,N_8323,N_8034);
nor U8757 (N_8757,N_8116,N_8157);
nor U8758 (N_8758,N_8076,N_8177);
or U8759 (N_8759,N_8015,N_8417);
nand U8760 (N_8760,N_8034,N_8039);
nor U8761 (N_8761,N_8334,N_8001);
and U8762 (N_8762,N_8410,N_8318);
nand U8763 (N_8763,N_8468,N_8477);
nor U8764 (N_8764,N_8025,N_8362);
or U8765 (N_8765,N_8304,N_8032);
nand U8766 (N_8766,N_8184,N_8098);
or U8767 (N_8767,N_8046,N_8281);
nor U8768 (N_8768,N_8065,N_8432);
or U8769 (N_8769,N_8496,N_8376);
and U8770 (N_8770,N_8469,N_8300);
xor U8771 (N_8771,N_8450,N_8086);
or U8772 (N_8772,N_8410,N_8436);
and U8773 (N_8773,N_8082,N_8031);
or U8774 (N_8774,N_8283,N_8258);
nor U8775 (N_8775,N_8465,N_8092);
nor U8776 (N_8776,N_8400,N_8441);
and U8777 (N_8777,N_8289,N_8170);
nor U8778 (N_8778,N_8494,N_8223);
nor U8779 (N_8779,N_8155,N_8114);
and U8780 (N_8780,N_8336,N_8325);
nor U8781 (N_8781,N_8446,N_8331);
and U8782 (N_8782,N_8088,N_8335);
or U8783 (N_8783,N_8008,N_8311);
and U8784 (N_8784,N_8007,N_8135);
and U8785 (N_8785,N_8398,N_8058);
or U8786 (N_8786,N_8351,N_8302);
and U8787 (N_8787,N_8474,N_8162);
nand U8788 (N_8788,N_8418,N_8449);
nor U8789 (N_8789,N_8260,N_8066);
and U8790 (N_8790,N_8354,N_8312);
nor U8791 (N_8791,N_8174,N_8068);
nand U8792 (N_8792,N_8085,N_8013);
nor U8793 (N_8793,N_8415,N_8464);
or U8794 (N_8794,N_8394,N_8347);
or U8795 (N_8795,N_8126,N_8075);
nor U8796 (N_8796,N_8174,N_8208);
and U8797 (N_8797,N_8224,N_8286);
nor U8798 (N_8798,N_8298,N_8348);
or U8799 (N_8799,N_8293,N_8214);
and U8800 (N_8800,N_8023,N_8386);
or U8801 (N_8801,N_8126,N_8488);
and U8802 (N_8802,N_8134,N_8013);
nand U8803 (N_8803,N_8476,N_8130);
nor U8804 (N_8804,N_8042,N_8252);
and U8805 (N_8805,N_8254,N_8171);
nand U8806 (N_8806,N_8066,N_8236);
or U8807 (N_8807,N_8003,N_8108);
nand U8808 (N_8808,N_8457,N_8031);
nand U8809 (N_8809,N_8013,N_8142);
or U8810 (N_8810,N_8167,N_8182);
or U8811 (N_8811,N_8436,N_8227);
nand U8812 (N_8812,N_8264,N_8436);
nor U8813 (N_8813,N_8396,N_8471);
and U8814 (N_8814,N_8415,N_8127);
and U8815 (N_8815,N_8026,N_8401);
nor U8816 (N_8816,N_8072,N_8105);
nor U8817 (N_8817,N_8225,N_8450);
nand U8818 (N_8818,N_8195,N_8071);
or U8819 (N_8819,N_8476,N_8089);
and U8820 (N_8820,N_8142,N_8080);
xnor U8821 (N_8821,N_8462,N_8172);
nand U8822 (N_8822,N_8475,N_8381);
and U8823 (N_8823,N_8403,N_8049);
and U8824 (N_8824,N_8055,N_8301);
or U8825 (N_8825,N_8171,N_8201);
or U8826 (N_8826,N_8126,N_8358);
and U8827 (N_8827,N_8440,N_8264);
or U8828 (N_8828,N_8096,N_8489);
and U8829 (N_8829,N_8196,N_8108);
nand U8830 (N_8830,N_8412,N_8167);
nor U8831 (N_8831,N_8219,N_8265);
nor U8832 (N_8832,N_8373,N_8056);
and U8833 (N_8833,N_8315,N_8450);
nand U8834 (N_8834,N_8423,N_8399);
nand U8835 (N_8835,N_8454,N_8106);
nor U8836 (N_8836,N_8443,N_8189);
and U8837 (N_8837,N_8413,N_8205);
nand U8838 (N_8838,N_8103,N_8176);
nand U8839 (N_8839,N_8018,N_8302);
or U8840 (N_8840,N_8272,N_8286);
or U8841 (N_8841,N_8370,N_8213);
xnor U8842 (N_8842,N_8490,N_8409);
or U8843 (N_8843,N_8057,N_8447);
or U8844 (N_8844,N_8083,N_8386);
nor U8845 (N_8845,N_8162,N_8318);
nand U8846 (N_8846,N_8488,N_8000);
nor U8847 (N_8847,N_8403,N_8389);
nand U8848 (N_8848,N_8156,N_8040);
nand U8849 (N_8849,N_8096,N_8240);
nor U8850 (N_8850,N_8467,N_8035);
nand U8851 (N_8851,N_8457,N_8325);
nor U8852 (N_8852,N_8312,N_8414);
nor U8853 (N_8853,N_8217,N_8265);
nor U8854 (N_8854,N_8262,N_8153);
and U8855 (N_8855,N_8294,N_8060);
and U8856 (N_8856,N_8427,N_8047);
and U8857 (N_8857,N_8231,N_8367);
and U8858 (N_8858,N_8433,N_8315);
or U8859 (N_8859,N_8398,N_8005);
and U8860 (N_8860,N_8126,N_8331);
nand U8861 (N_8861,N_8308,N_8021);
or U8862 (N_8862,N_8259,N_8423);
or U8863 (N_8863,N_8400,N_8038);
or U8864 (N_8864,N_8094,N_8498);
and U8865 (N_8865,N_8219,N_8157);
nor U8866 (N_8866,N_8277,N_8039);
or U8867 (N_8867,N_8316,N_8260);
or U8868 (N_8868,N_8015,N_8333);
and U8869 (N_8869,N_8428,N_8225);
or U8870 (N_8870,N_8290,N_8427);
nand U8871 (N_8871,N_8252,N_8463);
nor U8872 (N_8872,N_8061,N_8248);
nor U8873 (N_8873,N_8304,N_8055);
nor U8874 (N_8874,N_8361,N_8060);
nand U8875 (N_8875,N_8430,N_8015);
nor U8876 (N_8876,N_8338,N_8039);
or U8877 (N_8877,N_8397,N_8013);
or U8878 (N_8878,N_8121,N_8104);
or U8879 (N_8879,N_8065,N_8431);
nand U8880 (N_8880,N_8237,N_8300);
or U8881 (N_8881,N_8379,N_8265);
nor U8882 (N_8882,N_8228,N_8426);
xor U8883 (N_8883,N_8372,N_8410);
and U8884 (N_8884,N_8244,N_8285);
nand U8885 (N_8885,N_8307,N_8010);
nand U8886 (N_8886,N_8060,N_8120);
nand U8887 (N_8887,N_8012,N_8000);
nand U8888 (N_8888,N_8103,N_8184);
and U8889 (N_8889,N_8020,N_8335);
and U8890 (N_8890,N_8381,N_8152);
or U8891 (N_8891,N_8430,N_8356);
and U8892 (N_8892,N_8193,N_8285);
and U8893 (N_8893,N_8035,N_8031);
xor U8894 (N_8894,N_8287,N_8482);
nand U8895 (N_8895,N_8287,N_8418);
and U8896 (N_8896,N_8095,N_8209);
or U8897 (N_8897,N_8028,N_8337);
and U8898 (N_8898,N_8351,N_8259);
and U8899 (N_8899,N_8203,N_8055);
nand U8900 (N_8900,N_8248,N_8378);
nor U8901 (N_8901,N_8427,N_8431);
nor U8902 (N_8902,N_8260,N_8088);
nand U8903 (N_8903,N_8375,N_8255);
and U8904 (N_8904,N_8022,N_8325);
and U8905 (N_8905,N_8108,N_8056);
and U8906 (N_8906,N_8481,N_8160);
and U8907 (N_8907,N_8415,N_8354);
nor U8908 (N_8908,N_8365,N_8473);
nand U8909 (N_8909,N_8166,N_8477);
nor U8910 (N_8910,N_8115,N_8126);
nor U8911 (N_8911,N_8057,N_8255);
or U8912 (N_8912,N_8091,N_8233);
nand U8913 (N_8913,N_8054,N_8420);
and U8914 (N_8914,N_8297,N_8347);
nand U8915 (N_8915,N_8230,N_8149);
nor U8916 (N_8916,N_8345,N_8204);
or U8917 (N_8917,N_8239,N_8490);
and U8918 (N_8918,N_8460,N_8281);
nand U8919 (N_8919,N_8096,N_8214);
and U8920 (N_8920,N_8039,N_8324);
or U8921 (N_8921,N_8471,N_8172);
nand U8922 (N_8922,N_8043,N_8172);
nand U8923 (N_8923,N_8102,N_8345);
nor U8924 (N_8924,N_8251,N_8256);
nand U8925 (N_8925,N_8171,N_8221);
and U8926 (N_8926,N_8445,N_8402);
nand U8927 (N_8927,N_8040,N_8061);
or U8928 (N_8928,N_8466,N_8200);
and U8929 (N_8929,N_8445,N_8387);
or U8930 (N_8930,N_8183,N_8271);
and U8931 (N_8931,N_8276,N_8449);
nor U8932 (N_8932,N_8059,N_8072);
nor U8933 (N_8933,N_8437,N_8249);
or U8934 (N_8934,N_8340,N_8348);
or U8935 (N_8935,N_8264,N_8105);
or U8936 (N_8936,N_8035,N_8176);
nand U8937 (N_8937,N_8120,N_8399);
or U8938 (N_8938,N_8011,N_8229);
nor U8939 (N_8939,N_8362,N_8171);
nand U8940 (N_8940,N_8400,N_8218);
nand U8941 (N_8941,N_8284,N_8381);
and U8942 (N_8942,N_8259,N_8218);
nor U8943 (N_8943,N_8022,N_8371);
xnor U8944 (N_8944,N_8030,N_8272);
nor U8945 (N_8945,N_8223,N_8082);
nor U8946 (N_8946,N_8421,N_8417);
or U8947 (N_8947,N_8492,N_8318);
nor U8948 (N_8948,N_8262,N_8250);
or U8949 (N_8949,N_8076,N_8316);
and U8950 (N_8950,N_8199,N_8203);
and U8951 (N_8951,N_8198,N_8130);
xor U8952 (N_8952,N_8338,N_8200);
or U8953 (N_8953,N_8370,N_8492);
nand U8954 (N_8954,N_8168,N_8405);
and U8955 (N_8955,N_8212,N_8116);
or U8956 (N_8956,N_8039,N_8398);
or U8957 (N_8957,N_8432,N_8242);
or U8958 (N_8958,N_8338,N_8293);
and U8959 (N_8959,N_8283,N_8380);
and U8960 (N_8960,N_8417,N_8340);
and U8961 (N_8961,N_8173,N_8437);
nand U8962 (N_8962,N_8145,N_8394);
nor U8963 (N_8963,N_8026,N_8492);
and U8964 (N_8964,N_8007,N_8363);
and U8965 (N_8965,N_8498,N_8109);
nand U8966 (N_8966,N_8270,N_8424);
nand U8967 (N_8967,N_8156,N_8433);
or U8968 (N_8968,N_8226,N_8137);
and U8969 (N_8969,N_8365,N_8413);
and U8970 (N_8970,N_8194,N_8445);
xor U8971 (N_8971,N_8453,N_8313);
and U8972 (N_8972,N_8153,N_8168);
nand U8973 (N_8973,N_8200,N_8027);
xnor U8974 (N_8974,N_8202,N_8344);
nor U8975 (N_8975,N_8436,N_8230);
or U8976 (N_8976,N_8035,N_8214);
xor U8977 (N_8977,N_8206,N_8385);
nand U8978 (N_8978,N_8105,N_8280);
xor U8979 (N_8979,N_8353,N_8293);
nor U8980 (N_8980,N_8296,N_8337);
nor U8981 (N_8981,N_8108,N_8177);
nor U8982 (N_8982,N_8316,N_8461);
or U8983 (N_8983,N_8327,N_8399);
or U8984 (N_8984,N_8115,N_8314);
or U8985 (N_8985,N_8415,N_8283);
nor U8986 (N_8986,N_8151,N_8115);
or U8987 (N_8987,N_8017,N_8077);
or U8988 (N_8988,N_8297,N_8259);
nor U8989 (N_8989,N_8320,N_8125);
xnor U8990 (N_8990,N_8288,N_8440);
and U8991 (N_8991,N_8314,N_8103);
and U8992 (N_8992,N_8407,N_8038);
xnor U8993 (N_8993,N_8103,N_8167);
nor U8994 (N_8994,N_8235,N_8285);
nor U8995 (N_8995,N_8161,N_8333);
xor U8996 (N_8996,N_8467,N_8190);
nand U8997 (N_8997,N_8243,N_8297);
nor U8998 (N_8998,N_8481,N_8233);
or U8999 (N_8999,N_8157,N_8200);
xnor U9000 (N_9000,N_8722,N_8563);
or U9001 (N_9001,N_8804,N_8645);
nor U9002 (N_9002,N_8782,N_8866);
nand U9003 (N_9003,N_8575,N_8966);
nor U9004 (N_9004,N_8868,N_8737);
xor U9005 (N_9005,N_8806,N_8714);
nand U9006 (N_9006,N_8935,N_8781);
and U9007 (N_9007,N_8573,N_8917);
nor U9008 (N_9008,N_8888,N_8723);
and U9009 (N_9009,N_8658,N_8594);
nor U9010 (N_9010,N_8717,N_8607);
and U9011 (N_9011,N_8548,N_8916);
nand U9012 (N_9012,N_8997,N_8725);
nand U9013 (N_9013,N_8923,N_8684);
or U9014 (N_9014,N_8647,N_8859);
or U9015 (N_9015,N_8551,N_8559);
xor U9016 (N_9016,N_8757,N_8834);
nand U9017 (N_9017,N_8593,N_8924);
nor U9018 (N_9018,N_8977,N_8794);
nor U9019 (N_9019,N_8553,N_8908);
or U9020 (N_9020,N_8805,N_8585);
or U9021 (N_9021,N_8976,N_8960);
nor U9022 (N_9022,N_8820,N_8926);
nor U9023 (N_9023,N_8583,N_8918);
and U9024 (N_9024,N_8589,N_8832);
nand U9025 (N_9025,N_8919,N_8743);
nor U9026 (N_9026,N_8546,N_8547);
nor U9027 (N_9027,N_8721,N_8760);
nand U9028 (N_9028,N_8767,N_8894);
nor U9029 (N_9029,N_8776,N_8680);
nand U9030 (N_9030,N_8599,N_8984);
or U9031 (N_9031,N_8909,N_8939);
or U9032 (N_9032,N_8772,N_8655);
nor U9033 (N_9033,N_8770,N_8630);
nor U9034 (N_9034,N_8611,N_8615);
and U9035 (N_9035,N_8867,N_8540);
or U9036 (N_9036,N_8839,N_8500);
and U9037 (N_9037,N_8792,N_8683);
nor U9038 (N_9038,N_8861,N_8938);
and U9039 (N_9039,N_8904,N_8696);
or U9040 (N_9040,N_8850,N_8844);
or U9041 (N_9041,N_8821,N_8727);
or U9042 (N_9042,N_8665,N_8603);
xor U9043 (N_9043,N_8505,N_8522);
nor U9044 (N_9044,N_8813,N_8527);
xnor U9045 (N_9045,N_8664,N_8638);
nand U9046 (N_9046,N_8783,N_8745);
and U9047 (N_9047,N_8712,N_8831);
nor U9048 (N_9048,N_8542,N_8619);
xnor U9049 (N_9049,N_8653,N_8959);
nand U9050 (N_9050,N_8928,N_8726);
and U9051 (N_9051,N_8856,N_8953);
or U9052 (N_9052,N_8591,N_8571);
nor U9053 (N_9053,N_8561,N_8577);
xnor U9054 (N_9054,N_8506,N_8766);
xor U9055 (N_9055,N_8948,N_8718);
and U9056 (N_9056,N_8748,N_8639);
nor U9057 (N_9057,N_8833,N_8707);
nand U9058 (N_9058,N_8596,N_8525);
or U9059 (N_9059,N_8545,N_8930);
nand U9060 (N_9060,N_8880,N_8803);
xnor U9061 (N_9061,N_8974,N_8900);
and U9062 (N_9062,N_8969,N_8534);
nor U9063 (N_9063,N_8708,N_8808);
or U9064 (N_9064,N_8719,N_8830);
nor U9065 (N_9065,N_8656,N_8628);
or U9066 (N_9066,N_8740,N_8915);
and U9067 (N_9067,N_8756,N_8807);
xnor U9068 (N_9068,N_8787,N_8568);
nor U9069 (N_9069,N_8857,N_8914);
xnor U9070 (N_9070,N_8980,N_8738);
nand U9071 (N_9071,N_8840,N_8588);
or U9072 (N_9072,N_8514,N_8846);
nand U9073 (N_9073,N_8691,N_8537);
or U9074 (N_9074,N_8780,N_8598);
nor U9075 (N_9075,N_8896,N_8934);
nand U9076 (N_9076,N_8648,N_8695);
xor U9077 (N_9077,N_8529,N_8992);
and U9078 (N_9078,N_8771,N_8795);
xor U9079 (N_9079,N_8566,N_8870);
nor U9080 (N_9080,N_8632,N_8810);
nor U9081 (N_9081,N_8822,N_8642);
nand U9082 (N_9082,N_8701,N_8586);
nor U9083 (N_9083,N_8706,N_8758);
and U9084 (N_9084,N_8574,N_8978);
and U9085 (N_9085,N_8799,N_8724);
and U9086 (N_9086,N_8692,N_8754);
xor U9087 (N_9087,N_8581,N_8560);
nand U9088 (N_9088,N_8646,N_8951);
or U9089 (N_9089,N_8823,N_8623);
nand U9090 (N_9090,N_8616,N_8815);
or U9091 (N_9091,N_8836,N_8635);
nand U9092 (N_9092,N_8773,N_8601);
nor U9093 (N_9093,N_8733,N_8582);
and U9094 (N_9094,N_8925,N_8778);
nand U9095 (N_9095,N_8643,N_8986);
nor U9096 (N_9096,N_8842,N_8981);
and U9097 (N_9097,N_8901,N_8517);
nor U9098 (N_9098,N_8891,N_8634);
and U9099 (N_9099,N_8536,N_8541);
or U9100 (N_9100,N_8796,N_8749);
or U9101 (N_9101,N_8988,N_8570);
and U9102 (N_9102,N_8873,N_8535);
xor U9103 (N_9103,N_8613,N_8967);
or U9104 (N_9104,N_8689,N_8676);
nand U9105 (N_9105,N_8637,N_8965);
or U9106 (N_9106,N_8673,N_8902);
or U9107 (N_9107,N_8595,N_8858);
or U9108 (N_9108,N_8998,N_8544);
nand U9109 (N_9109,N_8819,N_8962);
or U9110 (N_9110,N_8704,N_8662);
and U9111 (N_9111,N_8788,N_8605);
nor U9112 (N_9112,N_8814,N_8983);
or U9113 (N_9113,N_8576,N_8955);
nand U9114 (N_9114,N_8732,N_8668);
xor U9115 (N_9115,N_8843,N_8612);
nand U9116 (N_9116,N_8511,N_8513);
nand U9117 (N_9117,N_8759,N_8625);
or U9118 (N_9118,N_8829,N_8985);
or U9119 (N_9119,N_8627,N_8768);
nand U9120 (N_9120,N_8713,N_8789);
or U9121 (N_9121,N_8851,N_8636);
nand U9122 (N_9122,N_8940,N_8621);
nor U9123 (N_9123,N_8694,N_8504);
nor U9124 (N_9124,N_8569,N_8971);
nand U9125 (N_9125,N_8958,N_8933);
nor U9126 (N_9126,N_8674,N_8785);
xor U9127 (N_9127,N_8578,N_8552);
nand U9128 (N_9128,N_8644,N_8633);
nor U9129 (N_9129,N_8961,N_8963);
nand U9130 (N_9130,N_8679,N_8956);
nor U9131 (N_9131,N_8661,N_8557);
nand U9132 (N_9132,N_8512,N_8996);
nor U9133 (N_9133,N_8518,N_8747);
or U9134 (N_9134,N_8920,N_8697);
xnor U9135 (N_9135,N_8729,N_8797);
or U9136 (N_9136,N_8502,N_8949);
or U9137 (N_9137,N_8641,N_8600);
nor U9138 (N_9138,N_8886,N_8811);
nor U9139 (N_9139,N_8584,N_8622);
nor U9140 (N_9140,N_8685,N_8614);
or U9141 (N_9141,N_8554,N_8703);
nor U9142 (N_9142,N_8530,N_8824);
or U9143 (N_9143,N_8895,N_8786);
and U9144 (N_9144,N_8883,N_8539);
or U9145 (N_9145,N_8790,N_8519);
and U9146 (N_9146,N_8515,N_8825);
and U9147 (N_9147,N_8802,N_8910);
nor U9148 (N_9148,N_8762,N_8884);
nand U9149 (N_9149,N_8798,N_8675);
nand U9150 (N_9150,N_8835,N_8592);
and U9151 (N_9151,N_8555,N_8763);
nand U9152 (N_9152,N_8678,N_8887);
nor U9153 (N_9153,N_8827,N_8970);
nand U9154 (N_9154,N_8651,N_8610);
and U9155 (N_9155,N_8777,N_8954);
nor U9156 (N_9156,N_8816,N_8994);
xor U9157 (N_9157,N_8649,N_8828);
and U9158 (N_9158,N_8657,N_8746);
and U9159 (N_9159,N_8550,N_8979);
xor U9160 (N_9160,N_8660,N_8855);
xnor U9161 (N_9161,N_8838,N_8892);
nand U9162 (N_9162,N_8862,N_8693);
and U9163 (N_9163,N_8687,N_8877);
nor U9164 (N_9164,N_8730,N_8874);
and U9165 (N_9165,N_8556,N_8975);
nor U9166 (N_9166,N_8659,N_8765);
nor U9167 (N_9167,N_8872,N_8507);
and U9168 (N_9168,N_8990,N_8620);
nor U9169 (N_9169,N_8736,N_8800);
xnor U9170 (N_9170,N_8698,N_8524);
and U9171 (N_9171,N_8587,N_8670);
nor U9172 (N_9172,N_8852,N_8624);
and U9173 (N_9173,N_8750,N_8860);
or U9174 (N_9174,N_8911,N_8899);
nor U9175 (N_9175,N_8944,N_8982);
nor U9176 (N_9176,N_8993,N_8501);
or U9177 (N_9177,N_8510,N_8631);
nand U9178 (N_9178,N_8590,N_8849);
nor U9179 (N_9179,N_8818,N_8526);
xor U9180 (N_9180,N_8650,N_8931);
or U9181 (N_9181,N_8952,N_8558);
and U9182 (N_9182,N_8879,N_8779);
or U9183 (N_9183,N_8618,N_8672);
nand U9184 (N_9184,N_8580,N_8898);
nand U9185 (N_9185,N_8709,N_8715);
or U9186 (N_9186,N_8533,N_8508);
or U9187 (N_9187,N_8640,N_8671);
or U9188 (N_9188,N_8741,N_8562);
or U9189 (N_9189,N_8989,N_8769);
xnor U9190 (N_9190,N_8876,N_8865);
or U9191 (N_9191,N_8932,N_8869);
and U9192 (N_9192,N_8602,N_8654);
or U9193 (N_9193,N_8669,N_8735);
nand U9194 (N_9194,N_8503,N_8878);
and U9195 (N_9195,N_8964,N_8549);
nand U9196 (N_9196,N_8700,N_8626);
or U9197 (N_9197,N_8791,N_8841);
xor U9198 (N_9198,N_8973,N_8538);
nand U9199 (N_9199,N_8809,N_8881);
nand U9200 (N_9200,N_8532,N_8751);
nor U9201 (N_9201,N_8764,N_8528);
nor U9202 (N_9202,N_8991,N_8572);
xnor U9203 (N_9203,N_8907,N_8663);
nand U9204 (N_9204,N_8710,N_8567);
nand U9205 (N_9205,N_8731,N_8753);
nor U9206 (N_9206,N_8677,N_8711);
or U9207 (N_9207,N_8995,N_8817);
nand U9208 (N_9208,N_8837,N_8688);
or U9209 (N_9209,N_8531,N_8972);
or U9210 (N_9210,N_8942,N_8608);
nor U9211 (N_9211,N_8667,N_8609);
nor U9212 (N_9212,N_8728,N_8604);
nor U9213 (N_9213,N_8606,N_8734);
nor U9214 (N_9214,N_8929,N_8987);
or U9215 (N_9215,N_8864,N_8912);
nand U9216 (N_9216,N_8775,N_8853);
or U9217 (N_9217,N_8897,N_8937);
nor U9218 (N_9218,N_8666,N_8913);
or U9219 (N_9219,N_8682,N_8742);
nand U9220 (N_9220,N_8579,N_8686);
xor U9221 (N_9221,N_8516,N_8543);
and U9222 (N_9222,N_8957,N_8968);
nand U9223 (N_9223,N_8521,N_8885);
nand U9224 (N_9224,N_8761,N_8854);
nand U9225 (N_9225,N_8509,N_8871);
and U9226 (N_9226,N_8523,N_8716);
nor U9227 (N_9227,N_8690,N_8597);
and U9228 (N_9228,N_8739,N_8699);
xnor U9229 (N_9229,N_8702,N_8520);
nor U9230 (N_9230,N_8946,N_8617);
or U9231 (N_9231,N_8947,N_8950);
xor U9232 (N_9232,N_8863,N_8893);
or U9233 (N_9233,N_8793,N_8652);
nor U9234 (N_9234,N_8826,N_8999);
and U9235 (N_9235,N_8629,N_8845);
or U9236 (N_9236,N_8784,N_8720);
or U9237 (N_9237,N_8936,N_8705);
nor U9238 (N_9238,N_8755,N_8943);
or U9239 (N_9239,N_8889,N_8744);
or U9240 (N_9240,N_8752,N_8890);
nor U9241 (N_9241,N_8945,N_8903);
nand U9242 (N_9242,N_8774,N_8847);
nor U9243 (N_9243,N_8922,N_8681);
or U9244 (N_9244,N_8941,N_8906);
xor U9245 (N_9245,N_8927,N_8882);
or U9246 (N_9246,N_8565,N_8564);
and U9247 (N_9247,N_8921,N_8905);
nand U9248 (N_9248,N_8848,N_8812);
nor U9249 (N_9249,N_8801,N_8875);
or U9250 (N_9250,N_8988,N_8919);
nand U9251 (N_9251,N_8992,N_8568);
or U9252 (N_9252,N_8591,N_8812);
and U9253 (N_9253,N_8820,N_8694);
and U9254 (N_9254,N_8581,N_8835);
or U9255 (N_9255,N_8691,N_8855);
nand U9256 (N_9256,N_8922,N_8904);
and U9257 (N_9257,N_8926,N_8819);
or U9258 (N_9258,N_8976,N_8988);
xor U9259 (N_9259,N_8738,N_8518);
nand U9260 (N_9260,N_8732,N_8974);
nand U9261 (N_9261,N_8818,N_8722);
nor U9262 (N_9262,N_8717,N_8609);
and U9263 (N_9263,N_8791,N_8838);
xnor U9264 (N_9264,N_8990,N_8574);
nand U9265 (N_9265,N_8917,N_8934);
xor U9266 (N_9266,N_8598,N_8922);
xnor U9267 (N_9267,N_8620,N_8613);
nand U9268 (N_9268,N_8810,N_8768);
xnor U9269 (N_9269,N_8884,N_8635);
nand U9270 (N_9270,N_8646,N_8704);
nand U9271 (N_9271,N_8592,N_8949);
or U9272 (N_9272,N_8697,N_8591);
and U9273 (N_9273,N_8911,N_8821);
xor U9274 (N_9274,N_8644,N_8574);
nand U9275 (N_9275,N_8863,N_8713);
or U9276 (N_9276,N_8671,N_8760);
or U9277 (N_9277,N_8843,N_8796);
nand U9278 (N_9278,N_8675,N_8931);
and U9279 (N_9279,N_8648,N_8580);
and U9280 (N_9280,N_8759,N_8764);
nor U9281 (N_9281,N_8788,N_8534);
nor U9282 (N_9282,N_8916,N_8813);
xor U9283 (N_9283,N_8760,N_8680);
or U9284 (N_9284,N_8900,N_8530);
nor U9285 (N_9285,N_8718,N_8810);
nand U9286 (N_9286,N_8826,N_8556);
or U9287 (N_9287,N_8927,N_8671);
nor U9288 (N_9288,N_8647,N_8772);
and U9289 (N_9289,N_8964,N_8565);
nor U9290 (N_9290,N_8519,N_8772);
or U9291 (N_9291,N_8935,N_8893);
nand U9292 (N_9292,N_8777,N_8532);
nor U9293 (N_9293,N_8640,N_8930);
nand U9294 (N_9294,N_8685,N_8657);
nand U9295 (N_9295,N_8622,N_8546);
nor U9296 (N_9296,N_8731,N_8695);
nor U9297 (N_9297,N_8879,N_8784);
nor U9298 (N_9298,N_8935,N_8749);
nor U9299 (N_9299,N_8872,N_8639);
nor U9300 (N_9300,N_8885,N_8741);
nor U9301 (N_9301,N_8613,N_8984);
xor U9302 (N_9302,N_8866,N_8870);
or U9303 (N_9303,N_8896,N_8974);
nand U9304 (N_9304,N_8581,N_8938);
nor U9305 (N_9305,N_8879,N_8599);
or U9306 (N_9306,N_8722,N_8841);
nand U9307 (N_9307,N_8719,N_8574);
nand U9308 (N_9308,N_8590,N_8940);
or U9309 (N_9309,N_8624,N_8760);
nor U9310 (N_9310,N_8662,N_8543);
xnor U9311 (N_9311,N_8992,N_8523);
and U9312 (N_9312,N_8983,N_8932);
and U9313 (N_9313,N_8907,N_8598);
xnor U9314 (N_9314,N_8747,N_8886);
nand U9315 (N_9315,N_8753,N_8932);
nand U9316 (N_9316,N_8812,N_8724);
or U9317 (N_9317,N_8605,N_8558);
or U9318 (N_9318,N_8599,N_8682);
nor U9319 (N_9319,N_8881,N_8819);
nand U9320 (N_9320,N_8828,N_8953);
and U9321 (N_9321,N_8636,N_8541);
and U9322 (N_9322,N_8508,N_8620);
and U9323 (N_9323,N_8948,N_8579);
nand U9324 (N_9324,N_8740,N_8755);
and U9325 (N_9325,N_8532,N_8922);
xnor U9326 (N_9326,N_8836,N_8618);
or U9327 (N_9327,N_8604,N_8575);
nand U9328 (N_9328,N_8584,N_8926);
or U9329 (N_9329,N_8691,N_8882);
nor U9330 (N_9330,N_8682,N_8684);
xor U9331 (N_9331,N_8820,N_8981);
nor U9332 (N_9332,N_8730,N_8797);
xnor U9333 (N_9333,N_8655,N_8797);
nor U9334 (N_9334,N_8973,N_8836);
and U9335 (N_9335,N_8771,N_8752);
or U9336 (N_9336,N_8743,N_8852);
nor U9337 (N_9337,N_8724,N_8716);
nand U9338 (N_9338,N_8881,N_8563);
xor U9339 (N_9339,N_8838,N_8712);
and U9340 (N_9340,N_8989,N_8797);
and U9341 (N_9341,N_8798,N_8548);
nor U9342 (N_9342,N_8917,N_8710);
nor U9343 (N_9343,N_8603,N_8844);
nor U9344 (N_9344,N_8937,N_8903);
nand U9345 (N_9345,N_8810,N_8554);
nand U9346 (N_9346,N_8854,N_8765);
or U9347 (N_9347,N_8717,N_8818);
and U9348 (N_9348,N_8690,N_8787);
nor U9349 (N_9349,N_8557,N_8713);
nand U9350 (N_9350,N_8651,N_8780);
nor U9351 (N_9351,N_8638,N_8678);
nand U9352 (N_9352,N_8992,N_8737);
and U9353 (N_9353,N_8555,N_8718);
and U9354 (N_9354,N_8557,N_8799);
nor U9355 (N_9355,N_8663,N_8734);
or U9356 (N_9356,N_8935,N_8746);
and U9357 (N_9357,N_8644,N_8856);
xor U9358 (N_9358,N_8706,N_8969);
nor U9359 (N_9359,N_8964,N_8590);
nand U9360 (N_9360,N_8550,N_8731);
and U9361 (N_9361,N_8909,N_8559);
and U9362 (N_9362,N_8654,N_8936);
or U9363 (N_9363,N_8940,N_8956);
or U9364 (N_9364,N_8774,N_8651);
and U9365 (N_9365,N_8833,N_8830);
nor U9366 (N_9366,N_8720,N_8780);
nand U9367 (N_9367,N_8945,N_8555);
nand U9368 (N_9368,N_8553,N_8541);
nor U9369 (N_9369,N_8894,N_8527);
or U9370 (N_9370,N_8522,N_8677);
xor U9371 (N_9371,N_8781,N_8882);
and U9372 (N_9372,N_8961,N_8597);
or U9373 (N_9373,N_8573,N_8789);
nor U9374 (N_9374,N_8894,N_8577);
nand U9375 (N_9375,N_8914,N_8711);
nor U9376 (N_9376,N_8681,N_8807);
nand U9377 (N_9377,N_8858,N_8717);
or U9378 (N_9378,N_8569,N_8745);
nor U9379 (N_9379,N_8721,N_8680);
nand U9380 (N_9380,N_8641,N_8708);
or U9381 (N_9381,N_8804,N_8724);
nor U9382 (N_9382,N_8663,N_8840);
xnor U9383 (N_9383,N_8730,N_8568);
xnor U9384 (N_9384,N_8944,N_8549);
or U9385 (N_9385,N_8525,N_8717);
nand U9386 (N_9386,N_8559,N_8937);
nand U9387 (N_9387,N_8879,N_8712);
or U9388 (N_9388,N_8900,N_8556);
nor U9389 (N_9389,N_8765,N_8569);
nand U9390 (N_9390,N_8567,N_8827);
or U9391 (N_9391,N_8520,N_8954);
or U9392 (N_9392,N_8545,N_8864);
or U9393 (N_9393,N_8882,N_8976);
xor U9394 (N_9394,N_8808,N_8640);
and U9395 (N_9395,N_8554,N_8900);
nand U9396 (N_9396,N_8679,N_8508);
nor U9397 (N_9397,N_8975,N_8597);
xnor U9398 (N_9398,N_8819,N_8590);
nand U9399 (N_9399,N_8516,N_8643);
or U9400 (N_9400,N_8602,N_8692);
and U9401 (N_9401,N_8768,N_8759);
nand U9402 (N_9402,N_8565,N_8790);
and U9403 (N_9403,N_8846,N_8559);
nand U9404 (N_9404,N_8578,N_8792);
nand U9405 (N_9405,N_8638,N_8600);
or U9406 (N_9406,N_8939,N_8577);
or U9407 (N_9407,N_8888,N_8709);
nand U9408 (N_9408,N_8983,N_8605);
and U9409 (N_9409,N_8832,N_8561);
nor U9410 (N_9410,N_8590,N_8984);
nand U9411 (N_9411,N_8767,N_8782);
xor U9412 (N_9412,N_8618,N_8795);
and U9413 (N_9413,N_8541,N_8576);
nand U9414 (N_9414,N_8614,N_8920);
nand U9415 (N_9415,N_8885,N_8589);
or U9416 (N_9416,N_8924,N_8883);
xnor U9417 (N_9417,N_8858,N_8734);
nor U9418 (N_9418,N_8645,N_8872);
or U9419 (N_9419,N_8878,N_8693);
nor U9420 (N_9420,N_8658,N_8926);
and U9421 (N_9421,N_8782,N_8970);
nor U9422 (N_9422,N_8780,N_8991);
nand U9423 (N_9423,N_8582,N_8948);
and U9424 (N_9424,N_8967,N_8926);
nand U9425 (N_9425,N_8941,N_8690);
xnor U9426 (N_9426,N_8992,N_8973);
or U9427 (N_9427,N_8768,N_8813);
nor U9428 (N_9428,N_8817,N_8991);
xor U9429 (N_9429,N_8623,N_8562);
nand U9430 (N_9430,N_8649,N_8859);
nor U9431 (N_9431,N_8781,N_8878);
nand U9432 (N_9432,N_8520,N_8571);
and U9433 (N_9433,N_8880,N_8722);
and U9434 (N_9434,N_8751,N_8665);
or U9435 (N_9435,N_8826,N_8884);
nand U9436 (N_9436,N_8526,N_8639);
and U9437 (N_9437,N_8547,N_8576);
or U9438 (N_9438,N_8678,N_8637);
and U9439 (N_9439,N_8954,N_8731);
nand U9440 (N_9440,N_8785,N_8970);
nor U9441 (N_9441,N_8838,N_8773);
nand U9442 (N_9442,N_8820,N_8884);
nand U9443 (N_9443,N_8801,N_8931);
and U9444 (N_9444,N_8521,N_8581);
xor U9445 (N_9445,N_8624,N_8523);
nor U9446 (N_9446,N_8558,N_8764);
and U9447 (N_9447,N_8889,N_8871);
nand U9448 (N_9448,N_8544,N_8897);
xor U9449 (N_9449,N_8568,N_8500);
or U9450 (N_9450,N_8693,N_8896);
or U9451 (N_9451,N_8941,N_8762);
xnor U9452 (N_9452,N_8981,N_8533);
nor U9453 (N_9453,N_8908,N_8571);
xor U9454 (N_9454,N_8900,N_8582);
nor U9455 (N_9455,N_8976,N_8814);
or U9456 (N_9456,N_8680,N_8602);
and U9457 (N_9457,N_8830,N_8907);
and U9458 (N_9458,N_8689,N_8972);
or U9459 (N_9459,N_8742,N_8518);
and U9460 (N_9460,N_8596,N_8803);
or U9461 (N_9461,N_8717,N_8610);
nand U9462 (N_9462,N_8932,N_8695);
and U9463 (N_9463,N_8908,N_8678);
nor U9464 (N_9464,N_8984,N_8839);
nand U9465 (N_9465,N_8602,N_8979);
and U9466 (N_9466,N_8690,N_8942);
nand U9467 (N_9467,N_8894,N_8872);
nor U9468 (N_9468,N_8977,N_8502);
nor U9469 (N_9469,N_8808,N_8926);
nor U9470 (N_9470,N_8511,N_8608);
nor U9471 (N_9471,N_8684,N_8812);
or U9472 (N_9472,N_8882,N_8982);
and U9473 (N_9473,N_8648,N_8923);
xor U9474 (N_9474,N_8509,N_8727);
and U9475 (N_9475,N_8929,N_8718);
and U9476 (N_9476,N_8778,N_8678);
nor U9477 (N_9477,N_8617,N_8867);
nor U9478 (N_9478,N_8955,N_8558);
nor U9479 (N_9479,N_8796,N_8744);
nor U9480 (N_9480,N_8598,N_8716);
and U9481 (N_9481,N_8970,N_8786);
nand U9482 (N_9482,N_8648,N_8811);
nand U9483 (N_9483,N_8716,N_8852);
nand U9484 (N_9484,N_8517,N_8511);
and U9485 (N_9485,N_8964,N_8705);
nand U9486 (N_9486,N_8633,N_8579);
nor U9487 (N_9487,N_8880,N_8764);
nor U9488 (N_9488,N_8770,N_8627);
xnor U9489 (N_9489,N_8923,N_8960);
and U9490 (N_9490,N_8693,N_8941);
and U9491 (N_9491,N_8956,N_8571);
or U9492 (N_9492,N_8658,N_8861);
or U9493 (N_9493,N_8819,N_8725);
nor U9494 (N_9494,N_8737,N_8556);
nor U9495 (N_9495,N_8838,N_8537);
nor U9496 (N_9496,N_8669,N_8740);
nand U9497 (N_9497,N_8750,N_8794);
and U9498 (N_9498,N_8801,N_8516);
and U9499 (N_9499,N_8832,N_8606);
nand U9500 (N_9500,N_9015,N_9200);
and U9501 (N_9501,N_9075,N_9455);
or U9502 (N_9502,N_9360,N_9473);
nand U9503 (N_9503,N_9343,N_9396);
nand U9504 (N_9504,N_9158,N_9294);
and U9505 (N_9505,N_9063,N_9460);
nand U9506 (N_9506,N_9375,N_9160);
nand U9507 (N_9507,N_9273,N_9078);
or U9508 (N_9508,N_9023,N_9133);
nand U9509 (N_9509,N_9028,N_9229);
nand U9510 (N_9510,N_9144,N_9207);
or U9511 (N_9511,N_9269,N_9424);
and U9512 (N_9512,N_9202,N_9352);
and U9513 (N_9513,N_9062,N_9035);
xor U9514 (N_9514,N_9115,N_9064);
or U9515 (N_9515,N_9212,N_9445);
nor U9516 (N_9516,N_9059,N_9211);
and U9517 (N_9517,N_9174,N_9026);
and U9518 (N_9518,N_9266,N_9238);
and U9519 (N_9519,N_9070,N_9085);
nand U9520 (N_9520,N_9168,N_9272);
and U9521 (N_9521,N_9492,N_9378);
or U9522 (N_9522,N_9182,N_9317);
xor U9523 (N_9523,N_9013,N_9397);
and U9524 (N_9524,N_9476,N_9382);
and U9525 (N_9525,N_9339,N_9190);
nand U9526 (N_9526,N_9243,N_9261);
nor U9527 (N_9527,N_9322,N_9346);
xnor U9528 (N_9528,N_9415,N_9076);
and U9529 (N_9529,N_9044,N_9439);
xnor U9530 (N_9530,N_9156,N_9403);
nor U9531 (N_9531,N_9001,N_9019);
and U9532 (N_9532,N_9305,N_9010);
nor U9533 (N_9533,N_9050,N_9459);
and U9534 (N_9534,N_9047,N_9486);
and U9535 (N_9535,N_9328,N_9184);
nand U9536 (N_9536,N_9496,N_9049);
or U9537 (N_9537,N_9082,N_9451);
and U9538 (N_9538,N_9142,N_9185);
nand U9539 (N_9539,N_9327,N_9043);
xnor U9540 (N_9540,N_9435,N_9358);
and U9541 (N_9541,N_9220,N_9086);
or U9542 (N_9542,N_9127,N_9253);
nor U9543 (N_9543,N_9157,N_9463);
and U9544 (N_9544,N_9102,N_9493);
nor U9545 (N_9545,N_9310,N_9335);
nor U9546 (N_9546,N_9409,N_9377);
nand U9547 (N_9547,N_9180,N_9237);
nor U9548 (N_9548,N_9080,N_9318);
nor U9549 (N_9549,N_9119,N_9487);
nand U9550 (N_9550,N_9155,N_9203);
or U9551 (N_9551,N_9005,N_9234);
or U9552 (N_9552,N_9095,N_9458);
nor U9553 (N_9553,N_9226,N_9466);
and U9554 (N_9554,N_9242,N_9012);
nand U9555 (N_9555,N_9427,N_9150);
nand U9556 (N_9556,N_9152,N_9299);
nor U9557 (N_9557,N_9021,N_9483);
xor U9558 (N_9558,N_9280,N_9312);
nor U9559 (N_9559,N_9452,N_9347);
nor U9560 (N_9560,N_9351,N_9422);
and U9561 (N_9561,N_9368,N_9283);
nor U9562 (N_9562,N_9254,N_9364);
or U9563 (N_9563,N_9362,N_9471);
nand U9564 (N_9564,N_9292,N_9029);
xnor U9565 (N_9565,N_9033,N_9399);
nor U9566 (N_9566,N_9475,N_9104);
and U9567 (N_9567,N_9300,N_9222);
nor U9568 (N_9568,N_9416,N_9430);
and U9569 (N_9569,N_9369,N_9068);
nor U9570 (N_9570,N_9289,N_9225);
nor U9571 (N_9571,N_9365,N_9098);
or U9572 (N_9572,N_9125,N_9418);
xnor U9573 (N_9573,N_9126,N_9433);
xor U9574 (N_9574,N_9221,N_9441);
and U9575 (N_9575,N_9470,N_9281);
or U9576 (N_9576,N_9313,N_9159);
and U9577 (N_9577,N_9008,N_9214);
nor U9578 (N_9578,N_9199,N_9121);
nand U9579 (N_9579,N_9040,N_9349);
xor U9580 (N_9580,N_9355,N_9042);
nand U9581 (N_9581,N_9303,N_9301);
nand U9582 (N_9582,N_9107,N_9464);
nor U9583 (N_9583,N_9387,N_9039);
or U9584 (N_9584,N_9171,N_9112);
nand U9585 (N_9585,N_9004,N_9411);
nor U9586 (N_9586,N_9128,N_9162);
nand U9587 (N_9587,N_9089,N_9374);
or U9588 (N_9588,N_9109,N_9208);
or U9589 (N_9589,N_9041,N_9414);
and U9590 (N_9590,N_9359,N_9118);
and U9591 (N_9591,N_9498,N_9468);
and U9592 (N_9592,N_9361,N_9117);
or U9593 (N_9593,N_9205,N_9348);
nor U9594 (N_9594,N_9100,N_9077);
or U9595 (N_9595,N_9056,N_9209);
nor U9596 (N_9596,N_9438,N_9287);
and U9597 (N_9597,N_9179,N_9302);
nor U9598 (N_9598,N_9114,N_9477);
nand U9599 (N_9599,N_9259,N_9428);
or U9600 (N_9600,N_9389,N_9494);
and U9601 (N_9601,N_9055,N_9061);
or U9602 (N_9602,N_9137,N_9073);
nor U9603 (N_9603,N_9124,N_9081);
nor U9604 (N_9604,N_9123,N_9009);
and U9605 (N_9605,N_9099,N_9215);
or U9606 (N_9606,N_9405,N_9395);
or U9607 (N_9607,N_9198,N_9277);
nand U9608 (N_9608,N_9231,N_9178);
and U9609 (N_9609,N_9345,N_9290);
nor U9610 (N_9610,N_9083,N_9201);
or U9611 (N_9611,N_9412,N_9437);
nand U9612 (N_9612,N_9032,N_9265);
nor U9613 (N_9613,N_9279,N_9490);
nor U9614 (N_9614,N_9245,N_9380);
xor U9615 (N_9615,N_9181,N_9247);
or U9616 (N_9616,N_9331,N_9480);
or U9617 (N_9617,N_9274,N_9436);
nand U9618 (N_9618,N_9241,N_9461);
and U9619 (N_9619,N_9169,N_9210);
nor U9620 (N_9620,N_9097,N_9298);
and U9621 (N_9621,N_9235,N_9088);
nand U9622 (N_9622,N_9410,N_9334);
nor U9623 (N_9623,N_9110,N_9219);
nor U9624 (N_9624,N_9326,N_9014);
and U9625 (N_9625,N_9194,N_9392);
or U9626 (N_9626,N_9320,N_9297);
nand U9627 (N_9627,N_9094,N_9357);
or U9628 (N_9628,N_9367,N_9419);
nor U9629 (N_9629,N_9293,N_9046);
xor U9630 (N_9630,N_9031,N_9105);
or U9631 (N_9631,N_9193,N_9074);
or U9632 (N_9632,N_9204,N_9407);
nand U9633 (N_9633,N_9143,N_9398);
xnor U9634 (N_9634,N_9284,N_9340);
nor U9635 (N_9635,N_9051,N_9465);
and U9636 (N_9636,N_9216,N_9187);
and U9637 (N_9637,N_9354,N_9069);
nand U9638 (N_9638,N_9092,N_9079);
nand U9639 (N_9639,N_9325,N_9306);
nor U9640 (N_9640,N_9134,N_9307);
and U9641 (N_9641,N_9016,N_9191);
or U9642 (N_9642,N_9163,N_9282);
nand U9643 (N_9643,N_9379,N_9093);
and U9644 (N_9644,N_9066,N_9249);
and U9645 (N_9645,N_9034,N_9018);
nand U9646 (N_9646,N_9024,N_9206);
or U9647 (N_9647,N_9479,N_9048);
nand U9648 (N_9648,N_9006,N_9462);
or U9649 (N_9649,N_9038,N_9270);
or U9650 (N_9650,N_9329,N_9246);
xor U9651 (N_9651,N_9391,N_9295);
nor U9652 (N_9652,N_9236,N_9022);
nor U9653 (N_9653,N_9052,N_9469);
nor U9654 (N_9654,N_9091,N_9333);
nand U9655 (N_9655,N_9434,N_9218);
or U9656 (N_9656,N_9113,N_9054);
nor U9657 (N_9657,N_9332,N_9170);
nor U9658 (N_9658,N_9315,N_9224);
nor U9659 (N_9659,N_9271,N_9384);
nand U9660 (N_9660,N_9495,N_9278);
nand U9661 (N_9661,N_9154,N_9148);
nand U9662 (N_9662,N_9263,N_9372);
and U9663 (N_9663,N_9316,N_9065);
nand U9664 (N_9664,N_9344,N_9020);
nand U9665 (N_9665,N_9188,N_9256);
or U9666 (N_9666,N_9084,N_9484);
nor U9667 (N_9667,N_9267,N_9390);
nand U9668 (N_9668,N_9448,N_9239);
nor U9669 (N_9669,N_9167,N_9071);
or U9670 (N_9670,N_9120,N_9402);
and U9671 (N_9671,N_9045,N_9139);
nand U9672 (N_9672,N_9417,N_9145);
nor U9673 (N_9673,N_9406,N_9457);
nand U9674 (N_9674,N_9481,N_9251);
nand U9675 (N_9675,N_9002,N_9330);
nand U9676 (N_9676,N_9165,N_9227);
or U9677 (N_9677,N_9131,N_9108);
and U9678 (N_9678,N_9072,N_9176);
nor U9679 (N_9679,N_9175,N_9173);
nor U9680 (N_9680,N_9136,N_9447);
xor U9681 (N_9681,N_9404,N_9058);
or U9682 (N_9682,N_9250,N_9370);
and U9683 (N_9683,N_9000,N_9252);
nor U9684 (N_9684,N_9336,N_9443);
or U9685 (N_9685,N_9450,N_9177);
or U9686 (N_9686,N_9472,N_9067);
or U9687 (N_9687,N_9053,N_9423);
and U9688 (N_9688,N_9431,N_9376);
nor U9689 (N_9689,N_9444,N_9183);
nor U9690 (N_9690,N_9425,N_9116);
nor U9691 (N_9691,N_9296,N_9195);
nor U9692 (N_9692,N_9309,N_9025);
nand U9693 (N_9693,N_9166,N_9482);
nor U9694 (N_9694,N_9353,N_9401);
nor U9695 (N_9695,N_9146,N_9453);
and U9696 (N_9696,N_9103,N_9454);
or U9697 (N_9697,N_9314,N_9122);
or U9698 (N_9698,N_9230,N_9446);
or U9699 (N_9699,N_9456,N_9381);
nor U9700 (N_9700,N_9244,N_9217);
or U9701 (N_9701,N_9017,N_9090);
xnor U9702 (N_9702,N_9275,N_9385);
or U9703 (N_9703,N_9223,N_9011);
or U9704 (N_9704,N_9497,N_9311);
and U9705 (N_9705,N_9421,N_9106);
nand U9706 (N_9706,N_9262,N_9393);
nor U9707 (N_9707,N_9324,N_9149);
or U9708 (N_9708,N_9342,N_9388);
nand U9709 (N_9709,N_9386,N_9057);
and U9710 (N_9710,N_9356,N_9304);
nand U9711 (N_9711,N_9338,N_9260);
nand U9712 (N_9712,N_9132,N_9172);
nor U9713 (N_9713,N_9285,N_9140);
nand U9714 (N_9714,N_9420,N_9383);
or U9715 (N_9715,N_9192,N_9478);
nand U9716 (N_9716,N_9373,N_9488);
or U9717 (N_9717,N_9248,N_9240);
or U9718 (N_9718,N_9147,N_9485);
nor U9719 (N_9719,N_9129,N_9233);
or U9720 (N_9720,N_9196,N_9213);
xor U9721 (N_9721,N_9268,N_9060);
nor U9722 (N_9722,N_9153,N_9189);
nand U9723 (N_9723,N_9027,N_9255);
nand U9724 (N_9724,N_9291,N_9037);
and U9725 (N_9725,N_9426,N_9321);
or U9726 (N_9726,N_9489,N_9232);
nor U9727 (N_9727,N_9141,N_9432);
nor U9728 (N_9728,N_9161,N_9101);
or U9729 (N_9729,N_9130,N_9036);
xor U9730 (N_9730,N_9030,N_9197);
or U9731 (N_9731,N_9337,N_9400);
nand U9732 (N_9732,N_9366,N_9286);
nand U9733 (N_9733,N_9096,N_9264);
or U9734 (N_9734,N_9350,N_9499);
and U9735 (N_9735,N_9363,N_9491);
nand U9736 (N_9736,N_9467,N_9151);
and U9737 (N_9737,N_9449,N_9323);
and U9738 (N_9738,N_9111,N_9371);
or U9739 (N_9739,N_9288,N_9276);
nand U9740 (N_9740,N_9408,N_9164);
nand U9741 (N_9741,N_9258,N_9429);
xor U9742 (N_9742,N_9308,N_9440);
nand U9743 (N_9743,N_9007,N_9474);
nand U9744 (N_9744,N_9413,N_9186);
and U9745 (N_9745,N_9228,N_9341);
xnor U9746 (N_9746,N_9319,N_9138);
and U9747 (N_9747,N_9087,N_9257);
and U9748 (N_9748,N_9442,N_9394);
or U9749 (N_9749,N_9003,N_9135);
or U9750 (N_9750,N_9074,N_9055);
and U9751 (N_9751,N_9464,N_9060);
nor U9752 (N_9752,N_9364,N_9147);
xnor U9753 (N_9753,N_9296,N_9228);
and U9754 (N_9754,N_9273,N_9403);
or U9755 (N_9755,N_9072,N_9460);
nand U9756 (N_9756,N_9005,N_9489);
nor U9757 (N_9757,N_9239,N_9444);
nand U9758 (N_9758,N_9291,N_9169);
nor U9759 (N_9759,N_9491,N_9416);
and U9760 (N_9760,N_9496,N_9165);
nor U9761 (N_9761,N_9229,N_9416);
and U9762 (N_9762,N_9211,N_9481);
nor U9763 (N_9763,N_9007,N_9033);
or U9764 (N_9764,N_9414,N_9301);
and U9765 (N_9765,N_9119,N_9045);
nand U9766 (N_9766,N_9233,N_9014);
nand U9767 (N_9767,N_9332,N_9252);
nor U9768 (N_9768,N_9399,N_9279);
nor U9769 (N_9769,N_9478,N_9496);
or U9770 (N_9770,N_9064,N_9319);
nand U9771 (N_9771,N_9358,N_9008);
and U9772 (N_9772,N_9295,N_9091);
nand U9773 (N_9773,N_9315,N_9399);
nor U9774 (N_9774,N_9120,N_9325);
or U9775 (N_9775,N_9064,N_9182);
nor U9776 (N_9776,N_9341,N_9270);
or U9777 (N_9777,N_9275,N_9365);
nor U9778 (N_9778,N_9269,N_9154);
nand U9779 (N_9779,N_9216,N_9371);
nand U9780 (N_9780,N_9426,N_9069);
nand U9781 (N_9781,N_9368,N_9088);
and U9782 (N_9782,N_9171,N_9478);
nor U9783 (N_9783,N_9455,N_9381);
or U9784 (N_9784,N_9460,N_9393);
and U9785 (N_9785,N_9179,N_9356);
nor U9786 (N_9786,N_9100,N_9317);
nor U9787 (N_9787,N_9441,N_9296);
or U9788 (N_9788,N_9399,N_9496);
and U9789 (N_9789,N_9313,N_9377);
nand U9790 (N_9790,N_9249,N_9282);
and U9791 (N_9791,N_9375,N_9051);
nor U9792 (N_9792,N_9405,N_9387);
nand U9793 (N_9793,N_9465,N_9383);
xnor U9794 (N_9794,N_9308,N_9487);
nor U9795 (N_9795,N_9483,N_9312);
xor U9796 (N_9796,N_9093,N_9433);
and U9797 (N_9797,N_9101,N_9157);
xor U9798 (N_9798,N_9009,N_9331);
nor U9799 (N_9799,N_9209,N_9154);
nor U9800 (N_9800,N_9004,N_9277);
nand U9801 (N_9801,N_9190,N_9021);
and U9802 (N_9802,N_9386,N_9391);
nand U9803 (N_9803,N_9275,N_9016);
or U9804 (N_9804,N_9366,N_9303);
and U9805 (N_9805,N_9476,N_9255);
and U9806 (N_9806,N_9101,N_9198);
nand U9807 (N_9807,N_9325,N_9101);
nor U9808 (N_9808,N_9317,N_9202);
xnor U9809 (N_9809,N_9015,N_9423);
nand U9810 (N_9810,N_9303,N_9160);
nor U9811 (N_9811,N_9161,N_9020);
nor U9812 (N_9812,N_9282,N_9150);
nand U9813 (N_9813,N_9260,N_9292);
nor U9814 (N_9814,N_9081,N_9153);
or U9815 (N_9815,N_9121,N_9330);
nand U9816 (N_9816,N_9448,N_9486);
nor U9817 (N_9817,N_9108,N_9241);
nand U9818 (N_9818,N_9480,N_9243);
or U9819 (N_9819,N_9318,N_9245);
nand U9820 (N_9820,N_9325,N_9469);
nor U9821 (N_9821,N_9146,N_9080);
nand U9822 (N_9822,N_9425,N_9115);
or U9823 (N_9823,N_9074,N_9208);
or U9824 (N_9824,N_9206,N_9180);
and U9825 (N_9825,N_9387,N_9435);
or U9826 (N_9826,N_9467,N_9465);
or U9827 (N_9827,N_9245,N_9348);
or U9828 (N_9828,N_9334,N_9100);
nor U9829 (N_9829,N_9378,N_9441);
xor U9830 (N_9830,N_9458,N_9277);
or U9831 (N_9831,N_9196,N_9140);
or U9832 (N_9832,N_9107,N_9186);
or U9833 (N_9833,N_9055,N_9368);
or U9834 (N_9834,N_9145,N_9489);
xnor U9835 (N_9835,N_9185,N_9492);
nand U9836 (N_9836,N_9172,N_9323);
nand U9837 (N_9837,N_9495,N_9190);
nand U9838 (N_9838,N_9067,N_9073);
and U9839 (N_9839,N_9007,N_9435);
and U9840 (N_9840,N_9238,N_9316);
or U9841 (N_9841,N_9047,N_9467);
nand U9842 (N_9842,N_9377,N_9153);
nor U9843 (N_9843,N_9085,N_9040);
or U9844 (N_9844,N_9247,N_9413);
nand U9845 (N_9845,N_9407,N_9104);
nor U9846 (N_9846,N_9365,N_9356);
or U9847 (N_9847,N_9358,N_9016);
nand U9848 (N_9848,N_9008,N_9454);
nand U9849 (N_9849,N_9200,N_9063);
or U9850 (N_9850,N_9088,N_9108);
xnor U9851 (N_9851,N_9404,N_9464);
nor U9852 (N_9852,N_9189,N_9191);
and U9853 (N_9853,N_9334,N_9378);
or U9854 (N_9854,N_9396,N_9388);
and U9855 (N_9855,N_9193,N_9032);
nor U9856 (N_9856,N_9166,N_9132);
nor U9857 (N_9857,N_9199,N_9171);
xor U9858 (N_9858,N_9029,N_9406);
nor U9859 (N_9859,N_9326,N_9141);
and U9860 (N_9860,N_9226,N_9102);
or U9861 (N_9861,N_9086,N_9182);
and U9862 (N_9862,N_9034,N_9264);
xor U9863 (N_9863,N_9488,N_9491);
nand U9864 (N_9864,N_9148,N_9334);
nor U9865 (N_9865,N_9004,N_9299);
xor U9866 (N_9866,N_9197,N_9485);
and U9867 (N_9867,N_9054,N_9294);
or U9868 (N_9868,N_9429,N_9229);
xor U9869 (N_9869,N_9300,N_9139);
nand U9870 (N_9870,N_9021,N_9458);
nand U9871 (N_9871,N_9082,N_9297);
nor U9872 (N_9872,N_9238,N_9492);
nand U9873 (N_9873,N_9441,N_9320);
nor U9874 (N_9874,N_9253,N_9156);
xor U9875 (N_9875,N_9190,N_9092);
and U9876 (N_9876,N_9462,N_9011);
and U9877 (N_9877,N_9454,N_9265);
xor U9878 (N_9878,N_9072,N_9391);
xnor U9879 (N_9879,N_9410,N_9254);
nand U9880 (N_9880,N_9113,N_9296);
and U9881 (N_9881,N_9422,N_9039);
or U9882 (N_9882,N_9065,N_9079);
nor U9883 (N_9883,N_9309,N_9408);
or U9884 (N_9884,N_9428,N_9261);
xor U9885 (N_9885,N_9053,N_9374);
nand U9886 (N_9886,N_9071,N_9070);
nor U9887 (N_9887,N_9053,N_9117);
and U9888 (N_9888,N_9188,N_9084);
or U9889 (N_9889,N_9481,N_9314);
nand U9890 (N_9890,N_9401,N_9397);
and U9891 (N_9891,N_9152,N_9146);
nand U9892 (N_9892,N_9287,N_9383);
or U9893 (N_9893,N_9294,N_9377);
nor U9894 (N_9894,N_9093,N_9203);
nor U9895 (N_9895,N_9304,N_9012);
nor U9896 (N_9896,N_9332,N_9137);
or U9897 (N_9897,N_9330,N_9357);
and U9898 (N_9898,N_9200,N_9298);
nor U9899 (N_9899,N_9399,N_9347);
and U9900 (N_9900,N_9066,N_9425);
or U9901 (N_9901,N_9466,N_9045);
nor U9902 (N_9902,N_9169,N_9262);
nor U9903 (N_9903,N_9144,N_9232);
nor U9904 (N_9904,N_9488,N_9445);
and U9905 (N_9905,N_9050,N_9161);
or U9906 (N_9906,N_9365,N_9332);
xor U9907 (N_9907,N_9418,N_9274);
nor U9908 (N_9908,N_9447,N_9026);
and U9909 (N_9909,N_9397,N_9164);
nand U9910 (N_9910,N_9100,N_9276);
nand U9911 (N_9911,N_9106,N_9483);
xnor U9912 (N_9912,N_9440,N_9422);
xor U9913 (N_9913,N_9122,N_9072);
or U9914 (N_9914,N_9108,N_9135);
xor U9915 (N_9915,N_9170,N_9031);
nor U9916 (N_9916,N_9415,N_9085);
or U9917 (N_9917,N_9101,N_9298);
and U9918 (N_9918,N_9312,N_9055);
and U9919 (N_9919,N_9407,N_9175);
or U9920 (N_9920,N_9438,N_9384);
or U9921 (N_9921,N_9010,N_9123);
and U9922 (N_9922,N_9101,N_9117);
and U9923 (N_9923,N_9448,N_9324);
nor U9924 (N_9924,N_9489,N_9041);
nand U9925 (N_9925,N_9499,N_9159);
nand U9926 (N_9926,N_9256,N_9258);
or U9927 (N_9927,N_9064,N_9122);
and U9928 (N_9928,N_9219,N_9062);
nor U9929 (N_9929,N_9317,N_9093);
xnor U9930 (N_9930,N_9183,N_9308);
nand U9931 (N_9931,N_9064,N_9079);
and U9932 (N_9932,N_9162,N_9023);
and U9933 (N_9933,N_9411,N_9202);
xnor U9934 (N_9934,N_9498,N_9396);
or U9935 (N_9935,N_9338,N_9293);
and U9936 (N_9936,N_9011,N_9104);
nor U9937 (N_9937,N_9123,N_9020);
nand U9938 (N_9938,N_9230,N_9266);
nor U9939 (N_9939,N_9053,N_9429);
nor U9940 (N_9940,N_9413,N_9228);
or U9941 (N_9941,N_9127,N_9157);
and U9942 (N_9942,N_9035,N_9345);
xnor U9943 (N_9943,N_9310,N_9326);
nand U9944 (N_9944,N_9103,N_9386);
xnor U9945 (N_9945,N_9244,N_9020);
xnor U9946 (N_9946,N_9061,N_9129);
and U9947 (N_9947,N_9388,N_9190);
or U9948 (N_9948,N_9281,N_9214);
nor U9949 (N_9949,N_9369,N_9211);
nor U9950 (N_9950,N_9285,N_9065);
or U9951 (N_9951,N_9129,N_9063);
nand U9952 (N_9952,N_9220,N_9365);
nor U9953 (N_9953,N_9005,N_9372);
nand U9954 (N_9954,N_9213,N_9367);
or U9955 (N_9955,N_9110,N_9450);
xnor U9956 (N_9956,N_9282,N_9408);
or U9957 (N_9957,N_9273,N_9044);
and U9958 (N_9958,N_9141,N_9226);
and U9959 (N_9959,N_9404,N_9056);
or U9960 (N_9960,N_9038,N_9033);
nand U9961 (N_9961,N_9499,N_9077);
nor U9962 (N_9962,N_9325,N_9474);
xor U9963 (N_9963,N_9325,N_9086);
and U9964 (N_9964,N_9136,N_9287);
nor U9965 (N_9965,N_9314,N_9159);
xor U9966 (N_9966,N_9424,N_9250);
or U9967 (N_9967,N_9029,N_9457);
xnor U9968 (N_9968,N_9320,N_9087);
nand U9969 (N_9969,N_9240,N_9453);
nand U9970 (N_9970,N_9372,N_9356);
nor U9971 (N_9971,N_9162,N_9041);
nand U9972 (N_9972,N_9002,N_9110);
xnor U9973 (N_9973,N_9489,N_9428);
nor U9974 (N_9974,N_9490,N_9355);
nor U9975 (N_9975,N_9068,N_9344);
or U9976 (N_9976,N_9011,N_9323);
nor U9977 (N_9977,N_9147,N_9021);
and U9978 (N_9978,N_9231,N_9184);
and U9979 (N_9979,N_9112,N_9270);
nor U9980 (N_9980,N_9429,N_9084);
nand U9981 (N_9981,N_9036,N_9203);
nor U9982 (N_9982,N_9368,N_9227);
or U9983 (N_9983,N_9301,N_9023);
or U9984 (N_9984,N_9366,N_9157);
xnor U9985 (N_9985,N_9083,N_9473);
and U9986 (N_9986,N_9459,N_9033);
and U9987 (N_9987,N_9337,N_9368);
and U9988 (N_9988,N_9368,N_9327);
and U9989 (N_9989,N_9402,N_9140);
nand U9990 (N_9990,N_9140,N_9398);
nor U9991 (N_9991,N_9473,N_9081);
nor U9992 (N_9992,N_9229,N_9138);
nand U9993 (N_9993,N_9426,N_9108);
nor U9994 (N_9994,N_9496,N_9143);
and U9995 (N_9995,N_9294,N_9053);
and U9996 (N_9996,N_9333,N_9349);
nand U9997 (N_9997,N_9253,N_9037);
or U9998 (N_9998,N_9181,N_9376);
and U9999 (N_9999,N_9473,N_9430);
nor UO_0 (O_0,N_9632,N_9650);
nor UO_1 (O_1,N_9746,N_9622);
and UO_2 (O_2,N_9509,N_9556);
and UO_3 (O_3,N_9959,N_9812);
and UO_4 (O_4,N_9568,N_9845);
nand UO_5 (O_5,N_9712,N_9931);
nand UO_6 (O_6,N_9995,N_9641);
nand UO_7 (O_7,N_9524,N_9867);
or UO_8 (O_8,N_9715,N_9942);
nor UO_9 (O_9,N_9599,N_9777);
nor UO_10 (O_10,N_9864,N_9609);
nor UO_11 (O_11,N_9806,N_9674);
nor UO_12 (O_12,N_9789,N_9573);
nor UO_13 (O_13,N_9842,N_9802);
nor UO_14 (O_14,N_9516,N_9871);
nor UO_15 (O_15,N_9542,N_9693);
nor UO_16 (O_16,N_9587,N_9821);
or UO_17 (O_17,N_9608,N_9530);
or UO_18 (O_18,N_9730,N_9917);
and UO_19 (O_19,N_9903,N_9592);
nor UO_20 (O_20,N_9600,N_9776);
nor UO_21 (O_21,N_9831,N_9858);
and UO_22 (O_22,N_9896,N_9820);
or UO_23 (O_23,N_9668,N_9874);
and UO_24 (O_24,N_9703,N_9788);
and UO_25 (O_25,N_9898,N_9984);
and UO_26 (O_26,N_9624,N_9951);
or UO_27 (O_27,N_9676,N_9616);
nand UO_28 (O_28,N_9893,N_9673);
or UO_29 (O_29,N_9932,N_9745);
and UO_30 (O_30,N_9921,N_9866);
nor UO_31 (O_31,N_9571,N_9547);
and UO_32 (O_32,N_9907,N_9647);
nand UO_33 (O_33,N_9952,N_9737);
and UO_34 (O_34,N_9982,N_9838);
nand UO_35 (O_35,N_9805,N_9944);
or UO_36 (O_36,N_9511,N_9648);
nor UO_37 (O_37,N_9536,N_9618);
nand UO_38 (O_38,N_9878,N_9627);
nand UO_39 (O_39,N_9834,N_9644);
nor UO_40 (O_40,N_9904,N_9678);
nor UO_41 (O_41,N_9840,N_9671);
nand UO_42 (O_42,N_9625,N_9590);
and UO_43 (O_43,N_9976,N_9630);
nor UO_44 (O_44,N_9563,N_9827);
or UO_45 (O_45,N_9980,N_9537);
nand UO_46 (O_46,N_9615,N_9705);
or UO_47 (O_47,N_9817,N_9757);
or UO_48 (O_48,N_9844,N_9716);
nand UO_49 (O_49,N_9744,N_9654);
xor UO_50 (O_50,N_9800,N_9546);
nor UO_51 (O_51,N_9791,N_9635);
nor UO_52 (O_52,N_9836,N_9970);
or UO_53 (O_53,N_9819,N_9636);
and UO_54 (O_54,N_9642,N_9522);
and UO_55 (O_55,N_9728,N_9567);
or UO_56 (O_56,N_9652,N_9999);
nand UO_57 (O_57,N_9729,N_9538);
or UO_58 (O_58,N_9813,N_9792);
nor UO_59 (O_59,N_9640,N_9861);
nor UO_60 (O_60,N_9830,N_9850);
or UO_61 (O_61,N_9502,N_9753);
or UO_62 (O_62,N_9736,N_9988);
xor UO_63 (O_63,N_9755,N_9551);
and UO_64 (O_64,N_9779,N_9877);
nor UO_65 (O_65,N_9918,N_9666);
nor UO_66 (O_66,N_9963,N_9950);
nor UO_67 (O_67,N_9639,N_9684);
nor UO_68 (O_68,N_9928,N_9519);
xor UO_69 (O_69,N_9584,N_9939);
nor UO_70 (O_70,N_9555,N_9526);
or UO_71 (O_71,N_9869,N_9733);
xnor UO_72 (O_72,N_9667,N_9593);
and UO_73 (O_73,N_9930,N_9531);
nor UO_74 (O_74,N_9762,N_9771);
nor UO_75 (O_75,N_9694,N_9854);
and UO_76 (O_76,N_9832,N_9919);
xnor UO_77 (O_77,N_9882,N_9868);
nand UO_78 (O_78,N_9740,N_9911);
nor UO_79 (O_79,N_9621,N_9569);
and UO_80 (O_80,N_9612,N_9588);
nor UO_81 (O_81,N_9760,N_9646);
xnor UO_82 (O_82,N_9533,N_9848);
or UO_83 (O_83,N_9889,N_9763);
or UO_84 (O_84,N_9575,N_9698);
and UO_85 (O_85,N_9707,N_9933);
nand UO_86 (O_86,N_9752,N_9843);
nor UO_87 (O_87,N_9758,N_9875);
nand UO_88 (O_88,N_9727,N_9914);
xor UO_89 (O_89,N_9992,N_9947);
nor UO_90 (O_90,N_9987,N_9876);
or UO_91 (O_91,N_9965,N_9924);
nor UO_92 (O_92,N_9521,N_9807);
xnor UO_93 (O_93,N_9900,N_9796);
nor UO_94 (O_94,N_9535,N_9972);
or UO_95 (O_95,N_9529,N_9510);
nand UO_96 (O_96,N_9784,N_9564);
nand UO_97 (O_97,N_9525,N_9506);
xnor UO_98 (O_98,N_9815,N_9927);
nand UO_99 (O_99,N_9857,N_9895);
nor UO_100 (O_100,N_9662,N_9607);
xnor UO_101 (O_101,N_9527,N_9986);
nand UO_102 (O_102,N_9846,N_9709);
nor UO_103 (O_103,N_9899,N_9702);
nor UO_104 (O_104,N_9701,N_9532);
and UO_105 (O_105,N_9809,N_9721);
nand UO_106 (O_106,N_9724,N_9589);
and UO_107 (O_107,N_9717,N_9747);
xor UO_108 (O_108,N_9797,N_9759);
and UO_109 (O_109,N_9906,N_9946);
nand UO_110 (O_110,N_9623,N_9696);
or UO_111 (O_111,N_9826,N_9520);
and UO_112 (O_112,N_9565,N_9825);
xor UO_113 (O_113,N_9852,N_9704);
and UO_114 (O_114,N_9739,N_9656);
and UO_115 (O_115,N_9655,N_9783);
nor UO_116 (O_116,N_9505,N_9695);
xor UO_117 (O_117,N_9513,N_9808);
and UO_118 (O_118,N_9540,N_9816);
nor UO_119 (O_119,N_9598,N_9828);
and UO_120 (O_120,N_9929,N_9661);
or UO_121 (O_121,N_9708,N_9890);
nor UO_122 (O_122,N_9824,N_9572);
and UO_123 (O_123,N_9835,N_9998);
nor UO_124 (O_124,N_9734,N_9562);
and UO_125 (O_125,N_9945,N_9949);
nor UO_126 (O_126,N_9665,N_9981);
and UO_127 (O_127,N_9870,N_9672);
nor UO_128 (O_128,N_9793,N_9699);
xor UO_129 (O_129,N_9881,N_9604);
or UO_130 (O_130,N_9605,N_9971);
and UO_131 (O_131,N_9722,N_9775);
and UO_132 (O_132,N_9989,N_9691);
nor UO_133 (O_133,N_9620,N_9996);
nor UO_134 (O_134,N_9803,N_9905);
or UO_135 (O_135,N_9856,N_9968);
nand UO_136 (O_136,N_9862,N_9915);
and UO_137 (O_137,N_9580,N_9983);
or UO_138 (O_138,N_9786,N_9901);
nand UO_139 (O_139,N_9837,N_9985);
and UO_140 (O_140,N_9964,N_9660);
or UO_141 (O_141,N_9761,N_9884);
and UO_142 (O_142,N_9804,N_9500);
nor UO_143 (O_143,N_9833,N_9550);
or UO_144 (O_144,N_9934,N_9748);
xor UO_145 (O_145,N_9633,N_9956);
and UO_146 (O_146,N_9559,N_9926);
nand UO_147 (O_147,N_9766,N_9923);
nor UO_148 (O_148,N_9591,N_9799);
and UO_149 (O_149,N_9629,N_9638);
nor UO_150 (O_150,N_9891,N_9902);
or UO_151 (O_151,N_9725,N_9679);
nand UO_152 (O_152,N_9732,N_9860);
xor UO_153 (O_153,N_9936,N_9714);
nand UO_154 (O_154,N_9810,N_9941);
nor UO_155 (O_155,N_9549,N_9683);
and UO_156 (O_156,N_9570,N_9977);
and UO_157 (O_157,N_9626,N_9978);
or UO_158 (O_158,N_9953,N_9764);
and UO_159 (O_159,N_9872,N_9677);
and UO_160 (O_160,N_9610,N_9925);
xor UO_161 (O_161,N_9841,N_9628);
and UO_162 (O_162,N_9643,N_9781);
nand UO_163 (O_163,N_9670,N_9849);
xnor UO_164 (O_164,N_9504,N_9680);
or UO_165 (O_165,N_9772,N_9782);
nor UO_166 (O_166,N_9847,N_9710);
nand UO_167 (O_167,N_9664,N_9617);
nand UO_168 (O_168,N_9798,N_9773);
nor UO_169 (O_169,N_9553,N_9697);
or UO_170 (O_170,N_9961,N_9967);
and UO_171 (O_171,N_9780,N_9507);
or UO_172 (O_172,N_9853,N_9920);
nor UO_173 (O_173,N_9690,N_9974);
nor UO_174 (O_174,N_9686,N_9637);
nand UO_175 (O_175,N_9994,N_9910);
nand UO_176 (O_176,N_9885,N_9560);
and UO_177 (O_177,N_9576,N_9687);
nor UO_178 (O_178,N_9706,N_9993);
nor UO_179 (O_179,N_9916,N_9894);
or UO_180 (O_180,N_9548,N_9586);
or UO_181 (O_181,N_9514,N_9990);
and UO_182 (O_182,N_9790,N_9675);
and UO_183 (O_183,N_9606,N_9611);
and UO_184 (O_184,N_9688,N_9523);
nor UO_185 (O_185,N_9720,N_9501);
or UO_186 (O_186,N_9873,N_9958);
and UO_187 (O_187,N_9554,N_9940);
and UO_188 (O_188,N_9888,N_9508);
nor UO_189 (O_189,N_9711,N_9912);
and UO_190 (O_190,N_9863,N_9596);
and UO_191 (O_191,N_9651,N_9577);
or UO_192 (O_192,N_9887,N_9669);
nor UO_193 (O_193,N_9735,N_9613);
or UO_194 (O_194,N_9751,N_9619);
xor UO_195 (O_195,N_9908,N_9859);
nand UO_196 (O_196,N_9962,N_9597);
and UO_197 (O_197,N_9689,N_9973);
nor UO_198 (O_198,N_9685,N_9883);
or UO_199 (O_199,N_9658,N_9561);
nand UO_200 (O_200,N_9785,N_9544);
xor UO_201 (O_201,N_9659,N_9713);
nand UO_202 (O_202,N_9943,N_9566);
and UO_203 (O_203,N_9582,N_9767);
and UO_204 (O_204,N_9768,N_9997);
or UO_205 (O_205,N_9913,N_9743);
nor UO_206 (O_206,N_9517,N_9581);
and UO_207 (O_207,N_9991,N_9512);
nor UO_208 (O_208,N_9657,N_9583);
nor UO_209 (O_209,N_9634,N_9719);
nand UO_210 (O_210,N_9829,N_9794);
xor UO_211 (O_211,N_9855,N_9602);
and UO_212 (O_212,N_9811,N_9957);
nand UO_213 (O_213,N_9718,N_9543);
or UO_214 (O_214,N_9975,N_9528);
and UO_215 (O_215,N_9558,N_9534);
and UO_216 (O_216,N_9892,N_9574);
or UO_217 (O_217,N_9897,N_9594);
xnor UO_218 (O_218,N_9649,N_9922);
or UO_219 (O_219,N_9938,N_9937);
nand UO_220 (O_220,N_9778,N_9955);
nor UO_221 (O_221,N_9552,N_9738);
and UO_222 (O_222,N_9539,N_9754);
nand UO_223 (O_223,N_9700,N_9585);
or UO_224 (O_224,N_9822,N_9631);
nand UO_225 (O_225,N_9742,N_9979);
nor UO_226 (O_226,N_9503,N_9960);
and UO_227 (O_227,N_9769,N_9814);
and UO_228 (O_228,N_9595,N_9603);
or UO_229 (O_229,N_9909,N_9756);
xor UO_230 (O_230,N_9663,N_9741);
and UO_231 (O_231,N_9681,N_9614);
nand UO_232 (O_232,N_9749,N_9969);
or UO_233 (O_233,N_9865,N_9839);
nand UO_234 (O_234,N_9795,N_9774);
nand UO_235 (O_235,N_9801,N_9770);
nor UO_236 (O_236,N_9886,N_9851);
nor UO_237 (O_237,N_9731,N_9578);
and UO_238 (O_238,N_9823,N_9765);
or UO_239 (O_239,N_9750,N_9541);
nor UO_240 (O_240,N_9579,N_9787);
or UO_241 (O_241,N_9545,N_9954);
or UO_242 (O_242,N_9653,N_9645);
nand UO_243 (O_243,N_9948,N_9818);
nor UO_244 (O_244,N_9692,N_9557);
nand UO_245 (O_245,N_9682,N_9601);
xnor UO_246 (O_246,N_9518,N_9723);
and UO_247 (O_247,N_9880,N_9515);
and UO_248 (O_248,N_9879,N_9935);
and UO_249 (O_249,N_9726,N_9966);
nor UO_250 (O_250,N_9839,N_9654);
or UO_251 (O_251,N_9828,N_9525);
and UO_252 (O_252,N_9505,N_9599);
or UO_253 (O_253,N_9524,N_9619);
nor UO_254 (O_254,N_9899,N_9583);
or UO_255 (O_255,N_9551,N_9542);
nand UO_256 (O_256,N_9596,N_9520);
xnor UO_257 (O_257,N_9690,N_9525);
or UO_258 (O_258,N_9563,N_9678);
xor UO_259 (O_259,N_9547,N_9879);
and UO_260 (O_260,N_9989,N_9801);
nand UO_261 (O_261,N_9961,N_9970);
and UO_262 (O_262,N_9807,N_9897);
or UO_263 (O_263,N_9987,N_9642);
or UO_264 (O_264,N_9763,N_9789);
and UO_265 (O_265,N_9557,N_9634);
and UO_266 (O_266,N_9754,N_9826);
nor UO_267 (O_267,N_9888,N_9617);
and UO_268 (O_268,N_9516,N_9893);
or UO_269 (O_269,N_9711,N_9593);
and UO_270 (O_270,N_9849,N_9976);
and UO_271 (O_271,N_9873,N_9636);
or UO_272 (O_272,N_9709,N_9549);
or UO_273 (O_273,N_9534,N_9692);
nand UO_274 (O_274,N_9718,N_9871);
nor UO_275 (O_275,N_9881,N_9793);
nor UO_276 (O_276,N_9791,N_9604);
and UO_277 (O_277,N_9681,N_9848);
xnor UO_278 (O_278,N_9846,N_9716);
nor UO_279 (O_279,N_9527,N_9661);
or UO_280 (O_280,N_9793,N_9587);
nand UO_281 (O_281,N_9542,N_9893);
and UO_282 (O_282,N_9629,N_9848);
and UO_283 (O_283,N_9906,N_9579);
xor UO_284 (O_284,N_9702,N_9708);
nand UO_285 (O_285,N_9684,N_9879);
or UO_286 (O_286,N_9759,N_9818);
nor UO_287 (O_287,N_9725,N_9916);
nor UO_288 (O_288,N_9528,N_9622);
and UO_289 (O_289,N_9637,N_9696);
and UO_290 (O_290,N_9879,N_9699);
and UO_291 (O_291,N_9516,N_9769);
xnor UO_292 (O_292,N_9832,N_9874);
and UO_293 (O_293,N_9701,N_9994);
or UO_294 (O_294,N_9997,N_9734);
and UO_295 (O_295,N_9961,N_9917);
nor UO_296 (O_296,N_9577,N_9687);
or UO_297 (O_297,N_9582,N_9534);
nor UO_298 (O_298,N_9678,N_9748);
and UO_299 (O_299,N_9858,N_9562);
nor UO_300 (O_300,N_9981,N_9607);
or UO_301 (O_301,N_9589,N_9772);
nand UO_302 (O_302,N_9621,N_9649);
xnor UO_303 (O_303,N_9589,N_9814);
or UO_304 (O_304,N_9605,N_9821);
nor UO_305 (O_305,N_9854,N_9642);
and UO_306 (O_306,N_9827,N_9762);
nand UO_307 (O_307,N_9629,N_9657);
nor UO_308 (O_308,N_9632,N_9979);
nor UO_309 (O_309,N_9705,N_9728);
nor UO_310 (O_310,N_9562,N_9578);
or UO_311 (O_311,N_9664,N_9828);
or UO_312 (O_312,N_9726,N_9928);
nor UO_313 (O_313,N_9571,N_9990);
or UO_314 (O_314,N_9787,N_9993);
or UO_315 (O_315,N_9897,N_9715);
xnor UO_316 (O_316,N_9693,N_9751);
and UO_317 (O_317,N_9799,N_9571);
or UO_318 (O_318,N_9723,N_9952);
or UO_319 (O_319,N_9795,N_9875);
or UO_320 (O_320,N_9793,N_9825);
or UO_321 (O_321,N_9549,N_9874);
nand UO_322 (O_322,N_9855,N_9859);
or UO_323 (O_323,N_9724,N_9569);
and UO_324 (O_324,N_9847,N_9570);
or UO_325 (O_325,N_9918,N_9705);
nand UO_326 (O_326,N_9916,N_9601);
nor UO_327 (O_327,N_9669,N_9533);
nor UO_328 (O_328,N_9564,N_9693);
or UO_329 (O_329,N_9802,N_9871);
nor UO_330 (O_330,N_9591,N_9867);
xnor UO_331 (O_331,N_9569,N_9545);
nand UO_332 (O_332,N_9646,N_9725);
nand UO_333 (O_333,N_9811,N_9808);
or UO_334 (O_334,N_9762,N_9566);
xnor UO_335 (O_335,N_9957,N_9513);
or UO_336 (O_336,N_9657,N_9581);
xor UO_337 (O_337,N_9967,N_9627);
nor UO_338 (O_338,N_9989,N_9730);
and UO_339 (O_339,N_9935,N_9627);
nor UO_340 (O_340,N_9857,N_9636);
or UO_341 (O_341,N_9544,N_9960);
or UO_342 (O_342,N_9899,N_9907);
or UO_343 (O_343,N_9903,N_9611);
xnor UO_344 (O_344,N_9909,N_9686);
or UO_345 (O_345,N_9892,N_9732);
xor UO_346 (O_346,N_9828,N_9640);
nand UO_347 (O_347,N_9544,N_9737);
or UO_348 (O_348,N_9762,N_9876);
or UO_349 (O_349,N_9816,N_9859);
nand UO_350 (O_350,N_9902,N_9687);
nor UO_351 (O_351,N_9812,N_9659);
nand UO_352 (O_352,N_9996,N_9730);
nand UO_353 (O_353,N_9701,N_9833);
or UO_354 (O_354,N_9703,N_9689);
nor UO_355 (O_355,N_9984,N_9516);
or UO_356 (O_356,N_9692,N_9891);
or UO_357 (O_357,N_9917,N_9540);
nand UO_358 (O_358,N_9614,N_9732);
nand UO_359 (O_359,N_9934,N_9559);
and UO_360 (O_360,N_9917,N_9641);
nand UO_361 (O_361,N_9616,N_9631);
or UO_362 (O_362,N_9805,N_9708);
nand UO_363 (O_363,N_9634,N_9693);
and UO_364 (O_364,N_9806,N_9743);
nand UO_365 (O_365,N_9775,N_9719);
nand UO_366 (O_366,N_9925,N_9575);
and UO_367 (O_367,N_9526,N_9610);
nand UO_368 (O_368,N_9866,N_9610);
and UO_369 (O_369,N_9934,N_9943);
or UO_370 (O_370,N_9616,N_9975);
or UO_371 (O_371,N_9570,N_9643);
nor UO_372 (O_372,N_9854,N_9638);
and UO_373 (O_373,N_9554,N_9556);
and UO_374 (O_374,N_9846,N_9821);
nand UO_375 (O_375,N_9605,N_9997);
nand UO_376 (O_376,N_9832,N_9737);
nor UO_377 (O_377,N_9634,N_9951);
nor UO_378 (O_378,N_9948,N_9830);
nor UO_379 (O_379,N_9684,N_9726);
nand UO_380 (O_380,N_9861,N_9915);
nor UO_381 (O_381,N_9534,N_9578);
or UO_382 (O_382,N_9610,N_9661);
nor UO_383 (O_383,N_9914,N_9520);
and UO_384 (O_384,N_9560,N_9753);
and UO_385 (O_385,N_9571,N_9893);
nor UO_386 (O_386,N_9638,N_9795);
nor UO_387 (O_387,N_9966,N_9849);
nor UO_388 (O_388,N_9959,N_9677);
nand UO_389 (O_389,N_9662,N_9665);
nor UO_390 (O_390,N_9904,N_9677);
xor UO_391 (O_391,N_9627,N_9606);
nor UO_392 (O_392,N_9985,N_9769);
nand UO_393 (O_393,N_9967,N_9994);
or UO_394 (O_394,N_9781,N_9800);
nand UO_395 (O_395,N_9610,N_9708);
nand UO_396 (O_396,N_9759,N_9711);
or UO_397 (O_397,N_9997,N_9637);
xnor UO_398 (O_398,N_9693,N_9528);
xor UO_399 (O_399,N_9951,N_9617);
nand UO_400 (O_400,N_9837,N_9551);
or UO_401 (O_401,N_9790,N_9988);
and UO_402 (O_402,N_9533,N_9808);
nor UO_403 (O_403,N_9938,N_9578);
or UO_404 (O_404,N_9815,N_9847);
or UO_405 (O_405,N_9536,N_9738);
nor UO_406 (O_406,N_9962,N_9900);
nand UO_407 (O_407,N_9631,N_9856);
or UO_408 (O_408,N_9989,N_9591);
or UO_409 (O_409,N_9517,N_9567);
nand UO_410 (O_410,N_9618,N_9606);
nor UO_411 (O_411,N_9807,N_9759);
nor UO_412 (O_412,N_9507,N_9699);
xnor UO_413 (O_413,N_9944,N_9880);
nor UO_414 (O_414,N_9977,N_9577);
or UO_415 (O_415,N_9683,N_9616);
nand UO_416 (O_416,N_9802,N_9812);
and UO_417 (O_417,N_9769,N_9676);
and UO_418 (O_418,N_9571,N_9869);
and UO_419 (O_419,N_9951,N_9977);
and UO_420 (O_420,N_9869,N_9781);
or UO_421 (O_421,N_9515,N_9951);
nor UO_422 (O_422,N_9640,N_9744);
or UO_423 (O_423,N_9976,N_9869);
and UO_424 (O_424,N_9815,N_9705);
or UO_425 (O_425,N_9923,N_9756);
nand UO_426 (O_426,N_9605,N_9661);
and UO_427 (O_427,N_9637,N_9976);
and UO_428 (O_428,N_9812,N_9901);
and UO_429 (O_429,N_9916,N_9941);
nand UO_430 (O_430,N_9824,N_9719);
nand UO_431 (O_431,N_9903,N_9517);
and UO_432 (O_432,N_9755,N_9998);
nand UO_433 (O_433,N_9889,N_9633);
or UO_434 (O_434,N_9620,N_9512);
nand UO_435 (O_435,N_9694,N_9567);
nand UO_436 (O_436,N_9574,N_9866);
and UO_437 (O_437,N_9895,N_9784);
or UO_438 (O_438,N_9903,N_9938);
nor UO_439 (O_439,N_9685,N_9628);
xnor UO_440 (O_440,N_9505,N_9680);
nand UO_441 (O_441,N_9503,N_9793);
and UO_442 (O_442,N_9825,N_9945);
xor UO_443 (O_443,N_9852,N_9740);
nor UO_444 (O_444,N_9791,N_9538);
nor UO_445 (O_445,N_9778,N_9879);
nand UO_446 (O_446,N_9707,N_9709);
and UO_447 (O_447,N_9896,N_9699);
nand UO_448 (O_448,N_9717,N_9903);
xnor UO_449 (O_449,N_9507,N_9660);
nand UO_450 (O_450,N_9755,N_9903);
or UO_451 (O_451,N_9793,N_9758);
xnor UO_452 (O_452,N_9556,N_9750);
and UO_453 (O_453,N_9945,N_9639);
nor UO_454 (O_454,N_9972,N_9754);
and UO_455 (O_455,N_9835,N_9984);
or UO_456 (O_456,N_9820,N_9709);
and UO_457 (O_457,N_9672,N_9624);
or UO_458 (O_458,N_9731,N_9887);
nand UO_459 (O_459,N_9511,N_9729);
nand UO_460 (O_460,N_9531,N_9952);
or UO_461 (O_461,N_9944,N_9974);
nor UO_462 (O_462,N_9616,N_9633);
nor UO_463 (O_463,N_9564,N_9545);
xnor UO_464 (O_464,N_9909,N_9811);
xor UO_465 (O_465,N_9914,N_9781);
nor UO_466 (O_466,N_9919,N_9582);
nor UO_467 (O_467,N_9633,N_9965);
nand UO_468 (O_468,N_9878,N_9680);
nor UO_469 (O_469,N_9597,N_9711);
nor UO_470 (O_470,N_9668,N_9514);
and UO_471 (O_471,N_9847,N_9968);
or UO_472 (O_472,N_9669,N_9576);
nand UO_473 (O_473,N_9848,N_9796);
nand UO_474 (O_474,N_9968,N_9850);
nor UO_475 (O_475,N_9566,N_9865);
nand UO_476 (O_476,N_9784,N_9788);
nor UO_477 (O_477,N_9791,N_9658);
nand UO_478 (O_478,N_9651,N_9686);
nand UO_479 (O_479,N_9898,N_9838);
and UO_480 (O_480,N_9540,N_9864);
or UO_481 (O_481,N_9510,N_9803);
nand UO_482 (O_482,N_9967,N_9800);
and UO_483 (O_483,N_9669,N_9624);
xor UO_484 (O_484,N_9699,N_9776);
nand UO_485 (O_485,N_9722,N_9894);
xnor UO_486 (O_486,N_9876,N_9740);
and UO_487 (O_487,N_9857,N_9738);
nor UO_488 (O_488,N_9840,N_9575);
and UO_489 (O_489,N_9679,N_9793);
or UO_490 (O_490,N_9682,N_9569);
or UO_491 (O_491,N_9754,N_9571);
and UO_492 (O_492,N_9731,N_9868);
nand UO_493 (O_493,N_9535,N_9503);
and UO_494 (O_494,N_9625,N_9603);
nor UO_495 (O_495,N_9683,N_9702);
and UO_496 (O_496,N_9755,N_9687);
nor UO_497 (O_497,N_9566,N_9949);
nor UO_498 (O_498,N_9552,N_9874);
nand UO_499 (O_499,N_9960,N_9855);
nor UO_500 (O_500,N_9530,N_9879);
or UO_501 (O_501,N_9905,N_9658);
nor UO_502 (O_502,N_9987,N_9518);
nand UO_503 (O_503,N_9523,N_9559);
nor UO_504 (O_504,N_9838,N_9566);
nand UO_505 (O_505,N_9764,N_9679);
and UO_506 (O_506,N_9698,N_9930);
xor UO_507 (O_507,N_9691,N_9514);
and UO_508 (O_508,N_9895,N_9713);
nor UO_509 (O_509,N_9572,N_9874);
nor UO_510 (O_510,N_9886,N_9668);
and UO_511 (O_511,N_9550,N_9813);
nand UO_512 (O_512,N_9675,N_9676);
nand UO_513 (O_513,N_9503,N_9872);
nand UO_514 (O_514,N_9727,N_9681);
nor UO_515 (O_515,N_9939,N_9818);
nor UO_516 (O_516,N_9660,N_9817);
and UO_517 (O_517,N_9633,N_9572);
nor UO_518 (O_518,N_9756,N_9894);
and UO_519 (O_519,N_9856,N_9525);
nor UO_520 (O_520,N_9818,N_9605);
nor UO_521 (O_521,N_9617,N_9865);
nand UO_522 (O_522,N_9823,N_9772);
nor UO_523 (O_523,N_9880,N_9870);
nand UO_524 (O_524,N_9879,N_9554);
and UO_525 (O_525,N_9895,N_9798);
nand UO_526 (O_526,N_9822,N_9657);
or UO_527 (O_527,N_9805,N_9731);
nor UO_528 (O_528,N_9588,N_9682);
or UO_529 (O_529,N_9977,N_9559);
and UO_530 (O_530,N_9937,N_9688);
and UO_531 (O_531,N_9861,N_9877);
nor UO_532 (O_532,N_9625,N_9649);
nor UO_533 (O_533,N_9616,N_9970);
or UO_534 (O_534,N_9858,N_9502);
and UO_535 (O_535,N_9541,N_9514);
and UO_536 (O_536,N_9602,N_9951);
nand UO_537 (O_537,N_9870,N_9526);
and UO_538 (O_538,N_9620,N_9786);
and UO_539 (O_539,N_9642,N_9955);
nor UO_540 (O_540,N_9528,N_9826);
or UO_541 (O_541,N_9972,N_9662);
xor UO_542 (O_542,N_9909,N_9843);
or UO_543 (O_543,N_9693,N_9735);
nor UO_544 (O_544,N_9896,N_9621);
and UO_545 (O_545,N_9686,N_9781);
xor UO_546 (O_546,N_9621,N_9577);
nand UO_547 (O_547,N_9605,N_9694);
nor UO_548 (O_548,N_9762,N_9744);
xnor UO_549 (O_549,N_9865,N_9664);
and UO_550 (O_550,N_9977,N_9902);
or UO_551 (O_551,N_9565,N_9615);
and UO_552 (O_552,N_9750,N_9939);
and UO_553 (O_553,N_9869,N_9756);
nor UO_554 (O_554,N_9608,N_9962);
and UO_555 (O_555,N_9706,N_9680);
nor UO_556 (O_556,N_9612,N_9946);
nand UO_557 (O_557,N_9965,N_9573);
or UO_558 (O_558,N_9574,N_9632);
and UO_559 (O_559,N_9875,N_9952);
or UO_560 (O_560,N_9704,N_9996);
nor UO_561 (O_561,N_9786,N_9811);
and UO_562 (O_562,N_9874,N_9511);
and UO_563 (O_563,N_9586,N_9761);
nor UO_564 (O_564,N_9612,N_9747);
nand UO_565 (O_565,N_9877,N_9504);
nor UO_566 (O_566,N_9787,N_9937);
nand UO_567 (O_567,N_9551,N_9896);
nand UO_568 (O_568,N_9635,N_9714);
and UO_569 (O_569,N_9823,N_9669);
or UO_570 (O_570,N_9545,N_9999);
nand UO_571 (O_571,N_9695,N_9523);
or UO_572 (O_572,N_9524,N_9964);
or UO_573 (O_573,N_9665,N_9982);
nand UO_574 (O_574,N_9629,N_9926);
nand UO_575 (O_575,N_9702,N_9938);
nor UO_576 (O_576,N_9537,N_9971);
nand UO_577 (O_577,N_9900,N_9799);
nand UO_578 (O_578,N_9689,N_9853);
and UO_579 (O_579,N_9952,N_9517);
nor UO_580 (O_580,N_9881,N_9649);
or UO_581 (O_581,N_9763,N_9657);
nor UO_582 (O_582,N_9744,N_9761);
or UO_583 (O_583,N_9807,N_9654);
nor UO_584 (O_584,N_9631,N_9982);
or UO_585 (O_585,N_9846,N_9995);
or UO_586 (O_586,N_9753,N_9987);
nor UO_587 (O_587,N_9848,N_9819);
and UO_588 (O_588,N_9541,N_9573);
nand UO_589 (O_589,N_9537,N_9859);
or UO_590 (O_590,N_9676,N_9933);
or UO_591 (O_591,N_9993,N_9873);
xnor UO_592 (O_592,N_9869,N_9534);
or UO_593 (O_593,N_9743,N_9936);
nand UO_594 (O_594,N_9756,N_9598);
or UO_595 (O_595,N_9706,N_9646);
xnor UO_596 (O_596,N_9516,N_9604);
nand UO_597 (O_597,N_9560,N_9985);
xnor UO_598 (O_598,N_9867,N_9925);
xor UO_599 (O_599,N_9762,N_9720);
or UO_600 (O_600,N_9699,N_9579);
nand UO_601 (O_601,N_9563,N_9588);
or UO_602 (O_602,N_9683,N_9845);
or UO_603 (O_603,N_9867,N_9876);
nor UO_604 (O_604,N_9508,N_9615);
nor UO_605 (O_605,N_9529,N_9975);
nand UO_606 (O_606,N_9981,N_9653);
nand UO_607 (O_607,N_9705,N_9962);
xnor UO_608 (O_608,N_9755,N_9593);
nand UO_609 (O_609,N_9516,N_9646);
or UO_610 (O_610,N_9516,N_9928);
and UO_611 (O_611,N_9613,N_9954);
nor UO_612 (O_612,N_9894,N_9697);
nand UO_613 (O_613,N_9934,N_9643);
nor UO_614 (O_614,N_9618,N_9575);
and UO_615 (O_615,N_9607,N_9680);
nor UO_616 (O_616,N_9577,N_9949);
nand UO_617 (O_617,N_9911,N_9875);
nor UO_618 (O_618,N_9644,N_9803);
nand UO_619 (O_619,N_9517,N_9851);
and UO_620 (O_620,N_9892,N_9755);
and UO_621 (O_621,N_9859,N_9919);
and UO_622 (O_622,N_9970,N_9924);
or UO_623 (O_623,N_9784,N_9500);
or UO_624 (O_624,N_9993,N_9537);
nor UO_625 (O_625,N_9852,N_9943);
nor UO_626 (O_626,N_9580,N_9949);
and UO_627 (O_627,N_9812,N_9853);
or UO_628 (O_628,N_9855,N_9517);
or UO_629 (O_629,N_9580,N_9745);
nor UO_630 (O_630,N_9692,N_9660);
and UO_631 (O_631,N_9522,N_9772);
and UO_632 (O_632,N_9727,N_9631);
nand UO_633 (O_633,N_9813,N_9601);
nand UO_634 (O_634,N_9991,N_9942);
nand UO_635 (O_635,N_9661,N_9614);
nor UO_636 (O_636,N_9797,N_9545);
nor UO_637 (O_637,N_9927,N_9593);
and UO_638 (O_638,N_9507,N_9537);
and UO_639 (O_639,N_9732,N_9600);
nor UO_640 (O_640,N_9927,N_9727);
and UO_641 (O_641,N_9927,N_9752);
xor UO_642 (O_642,N_9851,N_9974);
or UO_643 (O_643,N_9725,N_9964);
nand UO_644 (O_644,N_9993,N_9669);
xor UO_645 (O_645,N_9740,N_9543);
or UO_646 (O_646,N_9664,N_9528);
nor UO_647 (O_647,N_9597,N_9644);
nand UO_648 (O_648,N_9630,N_9989);
xor UO_649 (O_649,N_9963,N_9822);
nor UO_650 (O_650,N_9880,N_9824);
and UO_651 (O_651,N_9782,N_9740);
nand UO_652 (O_652,N_9558,N_9737);
or UO_653 (O_653,N_9783,N_9596);
nor UO_654 (O_654,N_9696,N_9634);
or UO_655 (O_655,N_9686,N_9533);
nand UO_656 (O_656,N_9686,N_9735);
nor UO_657 (O_657,N_9897,N_9931);
and UO_658 (O_658,N_9959,N_9993);
nor UO_659 (O_659,N_9731,N_9626);
xnor UO_660 (O_660,N_9935,N_9647);
and UO_661 (O_661,N_9663,N_9593);
nor UO_662 (O_662,N_9902,N_9798);
or UO_663 (O_663,N_9654,N_9771);
and UO_664 (O_664,N_9545,N_9556);
and UO_665 (O_665,N_9775,N_9561);
and UO_666 (O_666,N_9504,N_9988);
nand UO_667 (O_667,N_9823,N_9759);
nor UO_668 (O_668,N_9798,N_9666);
xnor UO_669 (O_669,N_9928,N_9975);
nand UO_670 (O_670,N_9798,N_9916);
xnor UO_671 (O_671,N_9738,N_9887);
or UO_672 (O_672,N_9956,N_9743);
nor UO_673 (O_673,N_9799,N_9948);
xnor UO_674 (O_674,N_9821,N_9710);
nor UO_675 (O_675,N_9648,N_9896);
nand UO_676 (O_676,N_9948,N_9710);
nand UO_677 (O_677,N_9655,N_9546);
nor UO_678 (O_678,N_9523,N_9978);
xor UO_679 (O_679,N_9747,N_9835);
nand UO_680 (O_680,N_9533,N_9871);
nor UO_681 (O_681,N_9521,N_9776);
xor UO_682 (O_682,N_9944,N_9555);
and UO_683 (O_683,N_9820,N_9875);
xor UO_684 (O_684,N_9578,N_9921);
or UO_685 (O_685,N_9592,N_9729);
or UO_686 (O_686,N_9679,N_9504);
xor UO_687 (O_687,N_9828,N_9590);
or UO_688 (O_688,N_9508,N_9829);
or UO_689 (O_689,N_9881,N_9593);
and UO_690 (O_690,N_9900,N_9626);
xnor UO_691 (O_691,N_9746,N_9942);
nor UO_692 (O_692,N_9597,N_9515);
nand UO_693 (O_693,N_9748,N_9839);
nor UO_694 (O_694,N_9507,N_9737);
nand UO_695 (O_695,N_9702,N_9518);
nand UO_696 (O_696,N_9517,N_9854);
nand UO_697 (O_697,N_9884,N_9990);
and UO_698 (O_698,N_9856,N_9886);
nor UO_699 (O_699,N_9839,N_9598);
xor UO_700 (O_700,N_9963,N_9667);
nor UO_701 (O_701,N_9924,N_9663);
nor UO_702 (O_702,N_9558,N_9767);
nand UO_703 (O_703,N_9996,N_9644);
nor UO_704 (O_704,N_9758,N_9897);
nor UO_705 (O_705,N_9513,N_9542);
or UO_706 (O_706,N_9534,N_9955);
and UO_707 (O_707,N_9610,N_9918);
and UO_708 (O_708,N_9966,N_9702);
xor UO_709 (O_709,N_9930,N_9944);
and UO_710 (O_710,N_9742,N_9904);
and UO_711 (O_711,N_9968,N_9817);
nand UO_712 (O_712,N_9695,N_9511);
or UO_713 (O_713,N_9667,N_9549);
or UO_714 (O_714,N_9895,N_9619);
and UO_715 (O_715,N_9548,N_9516);
nor UO_716 (O_716,N_9652,N_9660);
nor UO_717 (O_717,N_9824,N_9689);
or UO_718 (O_718,N_9643,N_9524);
nor UO_719 (O_719,N_9699,N_9777);
xor UO_720 (O_720,N_9816,N_9745);
nor UO_721 (O_721,N_9580,N_9861);
nor UO_722 (O_722,N_9720,N_9886);
or UO_723 (O_723,N_9926,N_9567);
nor UO_724 (O_724,N_9857,N_9926);
and UO_725 (O_725,N_9687,N_9671);
nand UO_726 (O_726,N_9654,N_9631);
nand UO_727 (O_727,N_9890,N_9979);
xor UO_728 (O_728,N_9932,N_9601);
nor UO_729 (O_729,N_9973,N_9735);
or UO_730 (O_730,N_9881,N_9817);
nand UO_731 (O_731,N_9749,N_9868);
nand UO_732 (O_732,N_9535,N_9852);
nor UO_733 (O_733,N_9606,N_9520);
nand UO_734 (O_734,N_9778,N_9899);
or UO_735 (O_735,N_9962,N_9678);
nor UO_736 (O_736,N_9979,N_9653);
nor UO_737 (O_737,N_9854,N_9754);
nor UO_738 (O_738,N_9777,N_9803);
nand UO_739 (O_739,N_9907,N_9960);
nand UO_740 (O_740,N_9698,N_9957);
and UO_741 (O_741,N_9996,N_9580);
nand UO_742 (O_742,N_9956,N_9500);
xor UO_743 (O_743,N_9840,N_9991);
nor UO_744 (O_744,N_9703,N_9532);
nand UO_745 (O_745,N_9915,N_9939);
nand UO_746 (O_746,N_9647,N_9884);
nand UO_747 (O_747,N_9501,N_9960);
or UO_748 (O_748,N_9794,N_9660);
nand UO_749 (O_749,N_9529,N_9591);
and UO_750 (O_750,N_9665,N_9775);
nor UO_751 (O_751,N_9755,N_9776);
and UO_752 (O_752,N_9593,N_9958);
nor UO_753 (O_753,N_9546,N_9996);
nand UO_754 (O_754,N_9771,N_9557);
and UO_755 (O_755,N_9586,N_9838);
or UO_756 (O_756,N_9811,N_9722);
nand UO_757 (O_757,N_9880,N_9938);
or UO_758 (O_758,N_9782,N_9929);
nor UO_759 (O_759,N_9828,N_9652);
nand UO_760 (O_760,N_9724,N_9979);
or UO_761 (O_761,N_9584,N_9846);
or UO_762 (O_762,N_9964,N_9599);
and UO_763 (O_763,N_9569,N_9764);
nor UO_764 (O_764,N_9776,N_9807);
or UO_765 (O_765,N_9664,N_9898);
nand UO_766 (O_766,N_9548,N_9746);
and UO_767 (O_767,N_9923,N_9896);
xnor UO_768 (O_768,N_9940,N_9901);
nor UO_769 (O_769,N_9596,N_9981);
or UO_770 (O_770,N_9547,N_9625);
or UO_771 (O_771,N_9955,N_9670);
nand UO_772 (O_772,N_9652,N_9983);
or UO_773 (O_773,N_9667,N_9553);
and UO_774 (O_774,N_9798,N_9929);
and UO_775 (O_775,N_9984,N_9862);
and UO_776 (O_776,N_9925,N_9765);
nor UO_777 (O_777,N_9881,N_9629);
nand UO_778 (O_778,N_9965,N_9722);
nand UO_779 (O_779,N_9654,N_9795);
or UO_780 (O_780,N_9595,N_9979);
and UO_781 (O_781,N_9847,N_9584);
xnor UO_782 (O_782,N_9821,N_9992);
nor UO_783 (O_783,N_9933,N_9931);
nor UO_784 (O_784,N_9594,N_9899);
and UO_785 (O_785,N_9574,N_9641);
or UO_786 (O_786,N_9756,N_9835);
and UO_787 (O_787,N_9730,N_9799);
or UO_788 (O_788,N_9677,N_9698);
nor UO_789 (O_789,N_9971,N_9897);
nor UO_790 (O_790,N_9942,N_9947);
nand UO_791 (O_791,N_9749,N_9854);
nor UO_792 (O_792,N_9709,N_9564);
nand UO_793 (O_793,N_9979,N_9875);
nand UO_794 (O_794,N_9619,N_9759);
or UO_795 (O_795,N_9834,N_9853);
nor UO_796 (O_796,N_9823,N_9788);
or UO_797 (O_797,N_9612,N_9900);
xnor UO_798 (O_798,N_9981,N_9878);
nor UO_799 (O_799,N_9554,N_9973);
nand UO_800 (O_800,N_9739,N_9883);
and UO_801 (O_801,N_9720,N_9954);
or UO_802 (O_802,N_9675,N_9605);
or UO_803 (O_803,N_9675,N_9638);
or UO_804 (O_804,N_9654,N_9856);
and UO_805 (O_805,N_9704,N_9732);
and UO_806 (O_806,N_9606,N_9766);
and UO_807 (O_807,N_9779,N_9763);
or UO_808 (O_808,N_9507,N_9612);
nor UO_809 (O_809,N_9543,N_9766);
nand UO_810 (O_810,N_9812,N_9879);
nor UO_811 (O_811,N_9630,N_9770);
or UO_812 (O_812,N_9980,N_9652);
and UO_813 (O_813,N_9617,N_9797);
nand UO_814 (O_814,N_9669,N_9740);
xor UO_815 (O_815,N_9745,N_9644);
and UO_816 (O_816,N_9908,N_9507);
nand UO_817 (O_817,N_9999,N_9992);
nor UO_818 (O_818,N_9557,N_9716);
nor UO_819 (O_819,N_9721,N_9656);
and UO_820 (O_820,N_9692,N_9767);
nor UO_821 (O_821,N_9568,N_9500);
nand UO_822 (O_822,N_9989,N_9534);
xor UO_823 (O_823,N_9917,N_9749);
and UO_824 (O_824,N_9640,N_9837);
nand UO_825 (O_825,N_9568,N_9504);
or UO_826 (O_826,N_9907,N_9864);
nand UO_827 (O_827,N_9880,N_9781);
nor UO_828 (O_828,N_9583,N_9893);
and UO_829 (O_829,N_9633,N_9539);
nor UO_830 (O_830,N_9854,N_9783);
and UO_831 (O_831,N_9608,N_9735);
and UO_832 (O_832,N_9775,N_9783);
nand UO_833 (O_833,N_9562,N_9916);
nand UO_834 (O_834,N_9901,N_9647);
nor UO_835 (O_835,N_9971,N_9642);
nor UO_836 (O_836,N_9772,N_9570);
and UO_837 (O_837,N_9854,N_9803);
nand UO_838 (O_838,N_9939,N_9959);
nand UO_839 (O_839,N_9569,N_9968);
nor UO_840 (O_840,N_9576,N_9665);
and UO_841 (O_841,N_9959,N_9633);
or UO_842 (O_842,N_9544,N_9860);
and UO_843 (O_843,N_9572,N_9970);
nand UO_844 (O_844,N_9732,N_9797);
or UO_845 (O_845,N_9782,N_9921);
nor UO_846 (O_846,N_9500,N_9550);
xor UO_847 (O_847,N_9723,N_9790);
nor UO_848 (O_848,N_9879,N_9873);
and UO_849 (O_849,N_9896,N_9832);
nand UO_850 (O_850,N_9547,N_9856);
nand UO_851 (O_851,N_9945,N_9840);
nand UO_852 (O_852,N_9815,N_9995);
nand UO_853 (O_853,N_9746,N_9956);
nand UO_854 (O_854,N_9538,N_9659);
and UO_855 (O_855,N_9776,N_9680);
nor UO_856 (O_856,N_9998,N_9644);
nor UO_857 (O_857,N_9560,N_9610);
nand UO_858 (O_858,N_9668,N_9946);
nor UO_859 (O_859,N_9605,N_9907);
nand UO_860 (O_860,N_9528,N_9961);
or UO_861 (O_861,N_9862,N_9896);
nand UO_862 (O_862,N_9800,N_9817);
and UO_863 (O_863,N_9510,N_9519);
nor UO_864 (O_864,N_9945,N_9916);
xnor UO_865 (O_865,N_9993,N_9626);
nand UO_866 (O_866,N_9995,N_9578);
nand UO_867 (O_867,N_9541,N_9633);
or UO_868 (O_868,N_9641,N_9876);
or UO_869 (O_869,N_9891,N_9603);
or UO_870 (O_870,N_9871,N_9677);
nand UO_871 (O_871,N_9779,N_9986);
nor UO_872 (O_872,N_9915,N_9970);
and UO_873 (O_873,N_9987,N_9650);
xnor UO_874 (O_874,N_9968,N_9738);
nor UO_875 (O_875,N_9505,N_9526);
or UO_876 (O_876,N_9882,N_9721);
nand UO_877 (O_877,N_9767,N_9710);
nand UO_878 (O_878,N_9652,N_9702);
and UO_879 (O_879,N_9991,N_9947);
xnor UO_880 (O_880,N_9620,N_9764);
and UO_881 (O_881,N_9631,N_9936);
or UO_882 (O_882,N_9661,N_9628);
xor UO_883 (O_883,N_9652,N_9943);
and UO_884 (O_884,N_9719,N_9534);
nor UO_885 (O_885,N_9655,N_9940);
xnor UO_886 (O_886,N_9950,N_9971);
nor UO_887 (O_887,N_9976,N_9527);
nor UO_888 (O_888,N_9537,N_9560);
nand UO_889 (O_889,N_9834,N_9874);
nor UO_890 (O_890,N_9743,N_9700);
nand UO_891 (O_891,N_9621,N_9960);
or UO_892 (O_892,N_9568,N_9976);
or UO_893 (O_893,N_9713,N_9527);
and UO_894 (O_894,N_9937,N_9846);
or UO_895 (O_895,N_9600,N_9750);
or UO_896 (O_896,N_9650,N_9923);
xor UO_897 (O_897,N_9927,N_9920);
and UO_898 (O_898,N_9856,N_9565);
and UO_899 (O_899,N_9717,N_9518);
and UO_900 (O_900,N_9886,N_9810);
nand UO_901 (O_901,N_9740,N_9779);
nand UO_902 (O_902,N_9699,N_9758);
and UO_903 (O_903,N_9949,N_9512);
xnor UO_904 (O_904,N_9504,N_9944);
xnor UO_905 (O_905,N_9702,N_9755);
and UO_906 (O_906,N_9645,N_9888);
nor UO_907 (O_907,N_9995,N_9537);
nor UO_908 (O_908,N_9816,N_9920);
or UO_909 (O_909,N_9711,N_9680);
or UO_910 (O_910,N_9997,N_9668);
nand UO_911 (O_911,N_9756,N_9743);
or UO_912 (O_912,N_9526,N_9987);
or UO_913 (O_913,N_9733,N_9677);
xnor UO_914 (O_914,N_9819,N_9726);
and UO_915 (O_915,N_9807,N_9618);
nor UO_916 (O_916,N_9979,N_9567);
and UO_917 (O_917,N_9860,N_9753);
or UO_918 (O_918,N_9517,N_9819);
nand UO_919 (O_919,N_9524,N_9561);
nand UO_920 (O_920,N_9892,N_9629);
and UO_921 (O_921,N_9739,N_9619);
xnor UO_922 (O_922,N_9770,N_9985);
or UO_923 (O_923,N_9988,N_9574);
or UO_924 (O_924,N_9891,N_9691);
and UO_925 (O_925,N_9742,N_9822);
nor UO_926 (O_926,N_9631,N_9546);
or UO_927 (O_927,N_9537,N_9509);
or UO_928 (O_928,N_9796,N_9871);
nor UO_929 (O_929,N_9542,N_9637);
xnor UO_930 (O_930,N_9829,N_9972);
or UO_931 (O_931,N_9955,N_9611);
nor UO_932 (O_932,N_9740,N_9581);
and UO_933 (O_933,N_9838,N_9646);
nand UO_934 (O_934,N_9563,N_9899);
or UO_935 (O_935,N_9608,N_9851);
and UO_936 (O_936,N_9963,N_9990);
or UO_937 (O_937,N_9664,N_9810);
or UO_938 (O_938,N_9862,N_9621);
and UO_939 (O_939,N_9607,N_9506);
xnor UO_940 (O_940,N_9758,N_9967);
nand UO_941 (O_941,N_9848,N_9920);
and UO_942 (O_942,N_9904,N_9660);
and UO_943 (O_943,N_9795,N_9533);
nor UO_944 (O_944,N_9804,N_9868);
or UO_945 (O_945,N_9530,N_9979);
xnor UO_946 (O_946,N_9501,N_9601);
nor UO_947 (O_947,N_9510,N_9564);
or UO_948 (O_948,N_9888,N_9660);
nand UO_949 (O_949,N_9736,N_9786);
and UO_950 (O_950,N_9793,N_9963);
nor UO_951 (O_951,N_9718,N_9590);
nor UO_952 (O_952,N_9629,N_9751);
nor UO_953 (O_953,N_9927,N_9876);
and UO_954 (O_954,N_9605,N_9873);
nand UO_955 (O_955,N_9632,N_9611);
and UO_956 (O_956,N_9794,N_9854);
nand UO_957 (O_957,N_9554,N_9931);
nand UO_958 (O_958,N_9673,N_9534);
or UO_959 (O_959,N_9568,N_9867);
or UO_960 (O_960,N_9823,N_9998);
or UO_961 (O_961,N_9798,N_9621);
nand UO_962 (O_962,N_9768,N_9872);
nor UO_963 (O_963,N_9903,N_9645);
or UO_964 (O_964,N_9816,N_9822);
or UO_965 (O_965,N_9733,N_9859);
and UO_966 (O_966,N_9516,N_9751);
and UO_967 (O_967,N_9814,N_9986);
nand UO_968 (O_968,N_9710,N_9990);
nand UO_969 (O_969,N_9688,N_9951);
nand UO_970 (O_970,N_9893,N_9557);
and UO_971 (O_971,N_9731,N_9622);
nand UO_972 (O_972,N_9777,N_9784);
xor UO_973 (O_973,N_9804,N_9697);
nor UO_974 (O_974,N_9619,N_9983);
xor UO_975 (O_975,N_9875,N_9523);
nor UO_976 (O_976,N_9731,N_9634);
and UO_977 (O_977,N_9764,N_9663);
nand UO_978 (O_978,N_9689,N_9808);
nand UO_979 (O_979,N_9929,N_9988);
or UO_980 (O_980,N_9701,N_9723);
or UO_981 (O_981,N_9649,N_9805);
nand UO_982 (O_982,N_9986,N_9539);
xnor UO_983 (O_983,N_9985,N_9588);
xnor UO_984 (O_984,N_9930,N_9785);
and UO_985 (O_985,N_9672,N_9907);
or UO_986 (O_986,N_9705,N_9880);
and UO_987 (O_987,N_9719,N_9820);
xor UO_988 (O_988,N_9649,N_9757);
and UO_989 (O_989,N_9639,N_9624);
nand UO_990 (O_990,N_9746,N_9833);
and UO_991 (O_991,N_9823,N_9995);
or UO_992 (O_992,N_9597,N_9862);
nor UO_993 (O_993,N_9955,N_9863);
nor UO_994 (O_994,N_9948,N_9572);
or UO_995 (O_995,N_9963,N_9714);
and UO_996 (O_996,N_9946,N_9548);
and UO_997 (O_997,N_9588,N_9903);
nor UO_998 (O_998,N_9640,N_9593);
and UO_999 (O_999,N_9650,N_9747);
and UO_1000 (O_1000,N_9805,N_9809);
and UO_1001 (O_1001,N_9811,N_9970);
nand UO_1002 (O_1002,N_9917,N_9923);
xor UO_1003 (O_1003,N_9901,N_9781);
xor UO_1004 (O_1004,N_9584,N_9865);
or UO_1005 (O_1005,N_9839,N_9651);
or UO_1006 (O_1006,N_9733,N_9627);
nand UO_1007 (O_1007,N_9509,N_9630);
nand UO_1008 (O_1008,N_9904,N_9772);
nand UO_1009 (O_1009,N_9878,N_9715);
and UO_1010 (O_1010,N_9800,N_9902);
nand UO_1011 (O_1011,N_9674,N_9966);
nand UO_1012 (O_1012,N_9758,N_9751);
or UO_1013 (O_1013,N_9768,N_9998);
nor UO_1014 (O_1014,N_9555,N_9542);
nand UO_1015 (O_1015,N_9642,N_9502);
nand UO_1016 (O_1016,N_9792,N_9850);
or UO_1017 (O_1017,N_9542,N_9501);
and UO_1018 (O_1018,N_9796,N_9780);
nor UO_1019 (O_1019,N_9578,N_9787);
and UO_1020 (O_1020,N_9613,N_9826);
nor UO_1021 (O_1021,N_9665,N_9841);
nor UO_1022 (O_1022,N_9659,N_9974);
and UO_1023 (O_1023,N_9763,N_9945);
nor UO_1024 (O_1024,N_9714,N_9682);
nand UO_1025 (O_1025,N_9759,N_9915);
and UO_1026 (O_1026,N_9991,N_9765);
nand UO_1027 (O_1027,N_9896,N_9956);
and UO_1028 (O_1028,N_9670,N_9726);
nor UO_1029 (O_1029,N_9612,N_9532);
and UO_1030 (O_1030,N_9971,N_9761);
xor UO_1031 (O_1031,N_9845,N_9935);
or UO_1032 (O_1032,N_9506,N_9903);
and UO_1033 (O_1033,N_9591,N_9646);
nor UO_1034 (O_1034,N_9936,N_9890);
and UO_1035 (O_1035,N_9778,N_9932);
and UO_1036 (O_1036,N_9911,N_9997);
and UO_1037 (O_1037,N_9997,N_9590);
xnor UO_1038 (O_1038,N_9865,N_9905);
or UO_1039 (O_1039,N_9652,N_9870);
nor UO_1040 (O_1040,N_9522,N_9946);
nor UO_1041 (O_1041,N_9847,N_9620);
or UO_1042 (O_1042,N_9915,N_9545);
or UO_1043 (O_1043,N_9954,N_9710);
or UO_1044 (O_1044,N_9876,N_9787);
or UO_1045 (O_1045,N_9685,N_9956);
and UO_1046 (O_1046,N_9527,N_9842);
nand UO_1047 (O_1047,N_9790,N_9979);
or UO_1048 (O_1048,N_9565,N_9945);
and UO_1049 (O_1049,N_9667,N_9587);
and UO_1050 (O_1050,N_9978,N_9607);
and UO_1051 (O_1051,N_9701,N_9661);
nand UO_1052 (O_1052,N_9547,N_9752);
or UO_1053 (O_1053,N_9835,N_9852);
and UO_1054 (O_1054,N_9570,N_9684);
and UO_1055 (O_1055,N_9549,N_9899);
nand UO_1056 (O_1056,N_9831,N_9591);
and UO_1057 (O_1057,N_9812,N_9566);
or UO_1058 (O_1058,N_9972,N_9892);
or UO_1059 (O_1059,N_9792,N_9779);
or UO_1060 (O_1060,N_9866,N_9819);
nand UO_1061 (O_1061,N_9538,N_9683);
or UO_1062 (O_1062,N_9900,N_9659);
or UO_1063 (O_1063,N_9586,N_9779);
nor UO_1064 (O_1064,N_9597,N_9827);
nor UO_1065 (O_1065,N_9765,N_9552);
or UO_1066 (O_1066,N_9699,N_9670);
and UO_1067 (O_1067,N_9521,N_9541);
nor UO_1068 (O_1068,N_9703,N_9892);
and UO_1069 (O_1069,N_9510,N_9503);
or UO_1070 (O_1070,N_9713,N_9762);
nand UO_1071 (O_1071,N_9978,N_9671);
nand UO_1072 (O_1072,N_9514,N_9519);
nor UO_1073 (O_1073,N_9897,N_9530);
nor UO_1074 (O_1074,N_9690,N_9562);
or UO_1075 (O_1075,N_9855,N_9828);
nand UO_1076 (O_1076,N_9585,N_9560);
or UO_1077 (O_1077,N_9990,N_9730);
xnor UO_1078 (O_1078,N_9565,N_9688);
xnor UO_1079 (O_1079,N_9775,N_9593);
nand UO_1080 (O_1080,N_9724,N_9704);
or UO_1081 (O_1081,N_9644,N_9788);
and UO_1082 (O_1082,N_9673,N_9903);
and UO_1083 (O_1083,N_9795,N_9950);
nand UO_1084 (O_1084,N_9868,N_9819);
xor UO_1085 (O_1085,N_9600,N_9852);
or UO_1086 (O_1086,N_9604,N_9693);
and UO_1087 (O_1087,N_9543,N_9867);
and UO_1088 (O_1088,N_9812,N_9719);
nand UO_1089 (O_1089,N_9678,N_9850);
and UO_1090 (O_1090,N_9586,N_9759);
or UO_1091 (O_1091,N_9724,N_9679);
or UO_1092 (O_1092,N_9583,N_9821);
or UO_1093 (O_1093,N_9828,N_9734);
or UO_1094 (O_1094,N_9597,N_9682);
nand UO_1095 (O_1095,N_9960,N_9853);
nor UO_1096 (O_1096,N_9915,N_9793);
xnor UO_1097 (O_1097,N_9658,N_9594);
or UO_1098 (O_1098,N_9898,N_9710);
and UO_1099 (O_1099,N_9544,N_9984);
and UO_1100 (O_1100,N_9726,N_9696);
xor UO_1101 (O_1101,N_9843,N_9633);
nor UO_1102 (O_1102,N_9768,N_9747);
nand UO_1103 (O_1103,N_9696,N_9551);
and UO_1104 (O_1104,N_9821,N_9623);
nand UO_1105 (O_1105,N_9521,N_9692);
nor UO_1106 (O_1106,N_9522,N_9913);
and UO_1107 (O_1107,N_9715,N_9892);
and UO_1108 (O_1108,N_9840,N_9554);
nor UO_1109 (O_1109,N_9867,N_9644);
nand UO_1110 (O_1110,N_9559,N_9647);
nor UO_1111 (O_1111,N_9534,N_9526);
nand UO_1112 (O_1112,N_9690,N_9675);
nand UO_1113 (O_1113,N_9963,N_9612);
and UO_1114 (O_1114,N_9508,N_9843);
nor UO_1115 (O_1115,N_9912,N_9939);
xnor UO_1116 (O_1116,N_9811,N_9974);
and UO_1117 (O_1117,N_9712,N_9966);
and UO_1118 (O_1118,N_9526,N_9604);
or UO_1119 (O_1119,N_9787,N_9858);
xnor UO_1120 (O_1120,N_9508,N_9974);
and UO_1121 (O_1121,N_9634,N_9536);
and UO_1122 (O_1122,N_9821,N_9805);
or UO_1123 (O_1123,N_9933,N_9729);
nor UO_1124 (O_1124,N_9539,N_9936);
nand UO_1125 (O_1125,N_9610,N_9742);
nor UO_1126 (O_1126,N_9748,N_9977);
nand UO_1127 (O_1127,N_9882,N_9651);
nand UO_1128 (O_1128,N_9972,N_9556);
xor UO_1129 (O_1129,N_9576,N_9735);
nand UO_1130 (O_1130,N_9739,N_9917);
and UO_1131 (O_1131,N_9592,N_9564);
or UO_1132 (O_1132,N_9824,N_9928);
nand UO_1133 (O_1133,N_9862,N_9742);
xor UO_1134 (O_1134,N_9565,N_9644);
nor UO_1135 (O_1135,N_9919,N_9881);
or UO_1136 (O_1136,N_9957,N_9838);
nand UO_1137 (O_1137,N_9510,N_9876);
nor UO_1138 (O_1138,N_9615,N_9828);
or UO_1139 (O_1139,N_9697,N_9822);
xor UO_1140 (O_1140,N_9619,N_9506);
xnor UO_1141 (O_1141,N_9956,N_9529);
nor UO_1142 (O_1142,N_9571,N_9562);
and UO_1143 (O_1143,N_9528,N_9908);
and UO_1144 (O_1144,N_9792,N_9809);
nor UO_1145 (O_1145,N_9504,N_9914);
and UO_1146 (O_1146,N_9995,N_9825);
and UO_1147 (O_1147,N_9685,N_9809);
or UO_1148 (O_1148,N_9901,N_9540);
nand UO_1149 (O_1149,N_9793,N_9556);
and UO_1150 (O_1150,N_9749,N_9925);
and UO_1151 (O_1151,N_9886,N_9745);
nor UO_1152 (O_1152,N_9788,N_9579);
nand UO_1153 (O_1153,N_9658,N_9965);
or UO_1154 (O_1154,N_9516,N_9509);
nand UO_1155 (O_1155,N_9680,N_9986);
or UO_1156 (O_1156,N_9800,N_9736);
nor UO_1157 (O_1157,N_9725,N_9576);
nand UO_1158 (O_1158,N_9577,N_9503);
nand UO_1159 (O_1159,N_9727,N_9740);
or UO_1160 (O_1160,N_9559,N_9919);
nand UO_1161 (O_1161,N_9706,N_9662);
nor UO_1162 (O_1162,N_9748,N_9691);
nor UO_1163 (O_1163,N_9630,N_9881);
and UO_1164 (O_1164,N_9951,N_9836);
and UO_1165 (O_1165,N_9976,N_9530);
and UO_1166 (O_1166,N_9617,N_9687);
and UO_1167 (O_1167,N_9974,N_9967);
nand UO_1168 (O_1168,N_9680,N_9610);
nand UO_1169 (O_1169,N_9678,N_9790);
nor UO_1170 (O_1170,N_9514,N_9826);
nor UO_1171 (O_1171,N_9608,N_9964);
and UO_1172 (O_1172,N_9871,N_9887);
and UO_1173 (O_1173,N_9549,N_9693);
and UO_1174 (O_1174,N_9531,N_9681);
nor UO_1175 (O_1175,N_9659,N_9992);
xnor UO_1176 (O_1176,N_9841,N_9980);
or UO_1177 (O_1177,N_9575,N_9882);
or UO_1178 (O_1178,N_9991,N_9920);
and UO_1179 (O_1179,N_9988,N_9762);
xor UO_1180 (O_1180,N_9850,N_9819);
nor UO_1181 (O_1181,N_9593,N_9745);
nor UO_1182 (O_1182,N_9791,N_9621);
or UO_1183 (O_1183,N_9581,N_9914);
nor UO_1184 (O_1184,N_9888,N_9644);
or UO_1185 (O_1185,N_9792,N_9501);
xnor UO_1186 (O_1186,N_9898,N_9924);
or UO_1187 (O_1187,N_9827,N_9608);
or UO_1188 (O_1188,N_9971,N_9995);
or UO_1189 (O_1189,N_9684,N_9546);
or UO_1190 (O_1190,N_9534,N_9712);
nor UO_1191 (O_1191,N_9563,N_9674);
nor UO_1192 (O_1192,N_9524,N_9906);
or UO_1193 (O_1193,N_9814,N_9523);
nand UO_1194 (O_1194,N_9951,N_9744);
nor UO_1195 (O_1195,N_9979,N_9891);
nor UO_1196 (O_1196,N_9617,N_9596);
and UO_1197 (O_1197,N_9541,N_9727);
and UO_1198 (O_1198,N_9695,N_9701);
and UO_1199 (O_1199,N_9798,N_9910);
and UO_1200 (O_1200,N_9722,N_9723);
and UO_1201 (O_1201,N_9831,N_9978);
nand UO_1202 (O_1202,N_9999,N_9821);
nand UO_1203 (O_1203,N_9908,N_9861);
and UO_1204 (O_1204,N_9769,N_9741);
or UO_1205 (O_1205,N_9534,N_9739);
nor UO_1206 (O_1206,N_9558,N_9940);
nor UO_1207 (O_1207,N_9637,N_9500);
and UO_1208 (O_1208,N_9698,N_9519);
xor UO_1209 (O_1209,N_9583,N_9607);
nand UO_1210 (O_1210,N_9843,N_9645);
or UO_1211 (O_1211,N_9817,N_9691);
nand UO_1212 (O_1212,N_9571,N_9995);
nand UO_1213 (O_1213,N_9957,N_9645);
or UO_1214 (O_1214,N_9549,N_9701);
nand UO_1215 (O_1215,N_9507,N_9919);
nand UO_1216 (O_1216,N_9710,N_9809);
nor UO_1217 (O_1217,N_9749,N_9594);
or UO_1218 (O_1218,N_9607,N_9855);
and UO_1219 (O_1219,N_9727,N_9694);
or UO_1220 (O_1220,N_9869,N_9947);
or UO_1221 (O_1221,N_9578,N_9531);
nand UO_1222 (O_1222,N_9736,N_9966);
and UO_1223 (O_1223,N_9690,N_9522);
xor UO_1224 (O_1224,N_9817,N_9601);
or UO_1225 (O_1225,N_9633,N_9950);
nand UO_1226 (O_1226,N_9555,N_9765);
nand UO_1227 (O_1227,N_9619,N_9717);
and UO_1228 (O_1228,N_9727,N_9838);
and UO_1229 (O_1229,N_9539,N_9787);
xor UO_1230 (O_1230,N_9848,N_9592);
nand UO_1231 (O_1231,N_9995,N_9763);
nor UO_1232 (O_1232,N_9780,N_9863);
and UO_1233 (O_1233,N_9527,N_9963);
and UO_1234 (O_1234,N_9604,N_9742);
xnor UO_1235 (O_1235,N_9792,N_9972);
nand UO_1236 (O_1236,N_9514,N_9803);
xnor UO_1237 (O_1237,N_9741,N_9667);
or UO_1238 (O_1238,N_9938,N_9604);
or UO_1239 (O_1239,N_9575,N_9672);
and UO_1240 (O_1240,N_9536,N_9646);
and UO_1241 (O_1241,N_9893,N_9992);
and UO_1242 (O_1242,N_9855,N_9873);
and UO_1243 (O_1243,N_9853,N_9932);
and UO_1244 (O_1244,N_9501,N_9754);
nor UO_1245 (O_1245,N_9856,N_9605);
and UO_1246 (O_1246,N_9775,N_9956);
nor UO_1247 (O_1247,N_9514,N_9857);
nor UO_1248 (O_1248,N_9966,N_9834);
and UO_1249 (O_1249,N_9797,N_9935);
or UO_1250 (O_1250,N_9789,N_9857);
nor UO_1251 (O_1251,N_9905,N_9611);
nand UO_1252 (O_1252,N_9957,N_9963);
nand UO_1253 (O_1253,N_9872,N_9776);
nand UO_1254 (O_1254,N_9945,N_9816);
nand UO_1255 (O_1255,N_9571,N_9594);
nand UO_1256 (O_1256,N_9833,N_9953);
nor UO_1257 (O_1257,N_9843,N_9760);
nor UO_1258 (O_1258,N_9732,N_9606);
or UO_1259 (O_1259,N_9615,N_9643);
nor UO_1260 (O_1260,N_9982,N_9511);
nand UO_1261 (O_1261,N_9778,N_9521);
nand UO_1262 (O_1262,N_9737,N_9849);
nand UO_1263 (O_1263,N_9532,N_9720);
or UO_1264 (O_1264,N_9738,N_9795);
and UO_1265 (O_1265,N_9526,N_9749);
and UO_1266 (O_1266,N_9818,N_9828);
nand UO_1267 (O_1267,N_9973,N_9528);
and UO_1268 (O_1268,N_9608,N_9550);
or UO_1269 (O_1269,N_9593,N_9825);
or UO_1270 (O_1270,N_9839,N_9757);
and UO_1271 (O_1271,N_9960,N_9649);
nor UO_1272 (O_1272,N_9732,N_9575);
or UO_1273 (O_1273,N_9622,N_9655);
nand UO_1274 (O_1274,N_9807,N_9761);
and UO_1275 (O_1275,N_9596,N_9939);
and UO_1276 (O_1276,N_9685,N_9523);
and UO_1277 (O_1277,N_9822,N_9714);
or UO_1278 (O_1278,N_9843,N_9528);
and UO_1279 (O_1279,N_9791,N_9509);
nor UO_1280 (O_1280,N_9603,N_9532);
nor UO_1281 (O_1281,N_9866,N_9682);
nor UO_1282 (O_1282,N_9719,N_9912);
or UO_1283 (O_1283,N_9776,N_9653);
and UO_1284 (O_1284,N_9809,N_9715);
and UO_1285 (O_1285,N_9940,N_9935);
and UO_1286 (O_1286,N_9808,N_9636);
nor UO_1287 (O_1287,N_9774,N_9732);
nor UO_1288 (O_1288,N_9586,N_9511);
xnor UO_1289 (O_1289,N_9958,N_9913);
or UO_1290 (O_1290,N_9879,N_9939);
nor UO_1291 (O_1291,N_9536,N_9946);
and UO_1292 (O_1292,N_9652,N_9700);
and UO_1293 (O_1293,N_9882,N_9550);
or UO_1294 (O_1294,N_9903,N_9855);
nor UO_1295 (O_1295,N_9985,N_9642);
nor UO_1296 (O_1296,N_9764,N_9922);
and UO_1297 (O_1297,N_9706,N_9761);
xnor UO_1298 (O_1298,N_9910,N_9988);
nand UO_1299 (O_1299,N_9966,N_9782);
xor UO_1300 (O_1300,N_9540,N_9641);
or UO_1301 (O_1301,N_9895,N_9962);
nor UO_1302 (O_1302,N_9695,N_9678);
nand UO_1303 (O_1303,N_9735,N_9799);
xor UO_1304 (O_1304,N_9907,N_9758);
or UO_1305 (O_1305,N_9577,N_9901);
xnor UO_1306 (O_1306,N_9931,N_9599);
nand UO_1307 (O_1307,N_9638,N_9849);
nor UO_1308 (O_1308,N_9579,N_9718);
nand UO_1309 (O_1309,N_9629,N_9755);
nand UO_1310 (O_1310,N_9540,N_9963);
xnor UO_1311 (O_1311,N_9773,N_9900);
nand UO_1312 (O_1312,N_9558,N_9759);
nand UO_1313 (O_1313,N_9782,N_9602);
nor UO_1314 (O_1314,N_9832,N_9555);
nor UO_1315 (O_1315,N_9984,N_9577);
or UO_1316 (O_1316,N_9541,N_9856);
and UO_1317 (O_1317,N_9735,N_9728);
nand UO_1318 (O_1318,N_9527,N_9987);
and UO_1319 (O_1319,N_9869,N_9903);
xor UO_1320 (O_1320,N_9756,N_9645);
or UO_1321 (O_1321,N_9552,N_9585);
and UO_1322 (O_1322,N_9666,N_9520);
xor UO_1323 (O_1323,N_9854,N_9656);
nand UO_1324 (O_1324,N_9721,N_9733);
xnor UO_1325 (O_1325,N_9585,N_9603);
nand UO_1326 (O_1326,N_9654,N_9984);
nor UO_1327 (O_1327,N_9704,N_9938);
nand UO_1328 (O_1328,N_9661,N_9966);
and UO_1329 (O_1329,N_9733,N_9866);
xor UO_1330 (O_1330,N_9910,N_9990);
nand UO_1331 (O_1331,N_9969,N_9844);
nor UO_1332 (O_1332,N_9900,N_9995);
nand UO_1333 (O_1333,N_9831,N_9682);
nand UO_1334 (O_1334,N_9658,N_9558);
or UO_1335 (O_1335,N_9883,N_9655);
nand UO_1336 (O_1336,N_9813,N_9947);
nor UO_1337 (O_1337,N_9613,N_9821);
xor UO_1338 (O_1338,N_9592,N_9813);
nand UO_1339 (O_1339,N_9528,N_9505);
xor UO_1340 (O_1340,N_9524,N_9884);
and UO_1341 (O_1341,N_9872,N_9588);
nor UO_1342 (O_1342,N_9850,N_9571);
and UO_1343 (O_1343,N_9945,N_9646);
and UO_1344 (O_1344,N_9723,N_9561);
nand UO_1345 (O_1345,N_9697,N_9602);
and UO_1346 (O_1346,N_9532,N_9869);
nand UO_1347 (O_1347,N_9785,N_9582);
and UO_1348 (O_1348,N_9517,N_9958);
nand UO_1349 (O_1349,N_9585,N_9898);
nor UO_1350 (O_1350,N_9661,N_9943);
xnor UO_1351 (O_1351,N_9676,N_9573);
nand UO_1352 (O_1352,N_9502,N_9547);
nor UO_1353 (O_1353,N_9647,N_9874);
nand UO_1354 (O_1354,N_9932,N_9963);
nand UO_1355 (O_1355,N_9998,N_9852);
or UO_1356 (O_1356,N_9739,N_9752);
and UO_1357 (O_1357,N_9797,N_9517);
nand UO_1358 (O_1358,N_9545,N_9793);
or UO_1359 (O_1359,N_9768,N_9743);
nand UO_1360 (O_1360,N_9910,N_9604);
and UO_1361 (O_1361,N_9864,N_9729);
nand UO_1362 (O_1362,N_9505,N_9503);
nor UO_1363 (O_1363,N_9671,N_9912);
nand UO_1364 (O_1364,N_9697,N_9738);
nor UO_1365 (O_1365,N_9967,N_9811);
and UO_1366 (O_1366,N_9994,N_9755);
and UO_1367 (O_1367,N_9743,N_9631);
nor UO_1368 (O_1368,N_9644,N_9619);
nor UO_1369 (O_1369,N_9554,N_9709);
xnor UO_1370 (O_1370,N_9881,N_9780);
nor UO_1371 (O_1371,N_9691,N_9895);
nand UO_1372 (O_1372,N_9755,N_9874);
nor UO_1373 (O_1373,N_9841,N_9900);
nor UO_1374 (O_1374,N_9534,N_9944);
nor UO_1375 (O_1375,N_9635,N_9601);
or UO_1376 (O_1376,N_9608,N_9555);
and UO_1377 (O_1377,N_9971,N_9571);
or UO_1378 (O_1378,N_9814,N_9999);
nand UO_1379 (O_1379,N_9688,N_9615);
or UO_1380 (O_1380,N_9570,N_9830);
nand UO_1381 (O_1381,N_9773,N_9570);
or UO_1382 (O_1382,N_9707,N_9668);
nand UO_1383 (O_1383,N_9594,N_9723);
xnor UO_1384 (O_1384,N_9992,N_9870);
and UO_1385 (O_1385,N_9926,N_9940);
and UO_1386 (O_1386,N_9740,N_9529);
nor UO_1387 (O_1387,N_9869,N_9787);
and UO_1388 (O_1388,N_9632,N_9838);
nand UO_1389 (O_1389,N_9624,N_9882);
nor UO_1390 (O_1390,N_9931,N_9741);
xnor UO_1391 (O_1391,N_9865,N_9878);
xor UO_1392 (O_1392,N_9978,N_9946);
nor UO_1393 (O_1393,N_9542,N_9716);
or UO_1394 (O_1394,N_9819,N_9728);
or UO_1395 (O_1395,N_9757,N_9925);
nand UO_1396 (O_1396,N_9629,N_9656);
or UO_1397 (O_1397,N_9771,N_9609);
xor UO_1398 (O_1398,N_9927,N_9713);
nor UO_1399 (O_1399,N_9955,N_9525);
or UO_1400 (O_1400,N_9686,N_9503);
nand UO_1401 (O_1401,N_9601,N_9963);
nor UO_1402 (O_1402,N_9543,N_9800);
xnor UO_1403 (O_1403,N_9547,N_9638);
and UO_1404 (O_1404,N_9540,N_9668);
and UO_1405 (O_1405,N_9830,N_9727);
and UO_1406 (O_1406,N_9925,N_9964);
or UO_1407 (O_1407,N_9618,N_9707);
nor UO_1408 (O_1408,N_9886,N_9773);
nand UO_1409 (O_1409,N_9860,N_9644);
or UO_1410 (O_1410,N_9761,N_9994);
nor UO_1411 (O_1411,N_9686,N_9546);
nand UO_1412 (O_1412,N_9878,N_9975);
xnor UO_1413 (O_1413,N_9560,N_9840);
and UO_1414 (O_1414,N_9861,N_9578);
or UO_1415 (O_1415,N_9915,N_9717);
and UO_1416 (O_1416,N_9747,N_9935);
and UO_1417 (O_1417,N_9774,N_9996);
nor UO_1418 (O_1418,N_9806,N_9751);
xor UO_1419 (O_1419,N_9989,N_9504);
nand UO_1420 (O_1420,N_9504,N_9655);
and UO_1421 (O_1421,N_9754,N_9736);
nand UO_1422 (O_1422,N_9765,N_9898);
nor UO_1423 (O_1423,N_9654,N_9799);
nor UO_1424 (O_1424,N_9838,N_9888);
or UO_1425 (O_1425,N_9525,N_9897);
nor UO_1426 (O_1426,N_9961,N_9914);
nand UO_1427 (O_1427,N_9551,N_9883);
nand UO_1428 (O_1428,N_9752,N_9505);
nor UO_1429 (O_1429,N_9757,N_9884);
nand UO_1430 (O_1430,N_9630,N_9618);
or UO_1431 (O_1431,N_9765,N_9543);
and UO_1432 (O_1432,N_9966,N_9609);
and UO_1433 (O_1433,N_9628,N_9688);
and UO_1434 (O_1434,N_9769,N_9915);
or UO_1435 (O_1435,N_9952,N_9869);
xor UO_1436 (O_1436,N_9796,N_9514);
nand UO_1437 (O_1437,N_9637,N_9621);
nand UO_1438 (O_1438,N_9511,N_9629);
or UO_1439 (O_1439,N_9710,N_9619);
or UO_1440 (O_1440,N_9587,N_9847);
and UO_1441 (O_1441,N_9914,N_9958);
or UO_1442 (O_1442,N_9537,N_9949);
nand UO_1443 (O_1443,N_9564,N_9902);
nand UO_1444 (O_1444,N_9780,N_9989);
and UO_1445 (O_1445,N_9846,N_9522);
nand UO_1446 (O_1446,N_9690,N_9572);
xor UO_1447 (O_1447,N_9542,N_9998);
nand UO_1448 (O_1448,N_9747,N_9710);
xor UO_1449 (O_1449,N_9887,N_9742);
or UO_1450 (O_1450,N_9628,N_9506);
xnor UO_1451 (O_1451,N_9679,N_9706);
xor UO_1452 (O_1452,N_9545,N_9540);
and UO_1453 (O_1453,N_9786,N_9930);
xor UO_1454 (O_1454,N_9555,N_9627);
and UO_1455 (O_1455,N_9747,N_9741);
nand UO_1456 (O_1456,N_9870,N_9605);
or UO_1457 (O_1457,N_9577,N_9800);
nor UO_1458 (O_1458,N_9538,N_9924);
nand UO_1459 (O_1459,N_9897,N_9620);
and UO_1460 (O_1460,N_9825,N_9594);
nor UO_1461 (O_1461,N_9978,N_9794);
or UO_1462 (O_1462,N_9708,N_9653);
and UO_1463 (O_1463,N_9893,N_9675);
and UO_1464 (O_1464,N_9501,N_9510);
nor UO_1465 (O_1465,N_9984,N_9746);
xnor UO_1466 (O_1466,N_9783,N_9640);
xnor UO_1467 (O_1467,N_9671,N_9504);
or UO_1468 (O_1468,N_9954,N_9981);
and UO_1469 (O_1469,N_9794,N_9754);
nand UO_1470 (O_1470,N_9549,N_9538);
nor UO_1471 (O_1471,N_9988,N_9530);
nor UO_1472 (O_1472,N_9974,N_9554);
or UO_1473 (O_1473,N_9708,N_9582);
xnor UO_1474 (O_1474,N_9717,N_9900);
nand UO_1475 (O_1475,N_9504,N_9657);
or UO_1476 (O_1476,N_9677,N_9554);
nand UO_1477 (O_1477,N_9785,N_9745);
nand UO_1478 (O_1478,N_9855,N_9600);
and UO_1479 (O_1479,N_9927,N_9659);
nor UO_1480 (O_1480,N_9820,N_9706);
nor UO_1481 (O_1481,N_9839,N_9964);
and UO_1482 (O_1482,N_9964,N_9781);
nor UO_1483 (O_1483,N_9785,N_9915);
nand UO_1484 (O_1484,N_9922,N_9756);
nand UO_1485 (O_1485,N_9662,N_9759);
nor UO_1486 (O_1486,N_9715,N_9907);
nor UO_1487 (O_1487,N_9977,N_9795);
xor UO_1488 (O_1488,N_9950,N_9867);
and UO_1489 (O_1489,N_9695,N_9857);
nand UO_1490 (O_1490,N_9767,N_9734);
nor UO_1491 (O_1491,N_9719,N_9753);
nor UO_1492 (O_1492,N_9862,N_9948);
or UO_1493 (O_1493,N_9507,N_9710);
nand UO_1494 (O_1494,N_9668,N_9855);
nand UO_1495 (O_1495,N_9713,N_9715);
or UO_1496 (O_1496,N_9804,N_9687);
nor UO_1497 (O_1497,N_9522,N_9831);
nand UO_1498 (O_1498,N_9916,N_9504);
and UO_1499 (O_1499,N_9767,N_9600);
endmodule