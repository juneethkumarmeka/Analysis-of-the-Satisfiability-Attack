module basic_2000_20000_2500_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_569,In_1802);
nand U1 (N_1,In_993,In_788);
and U2 (N_2,In_339,In_1564);
nor U3 (N_3,In_425,In_1224);
nand U4 (N_4,In_252,In_680);
xnor U5 (N_5,In_1176,In_1416);
or U6 (N_6,In_599,In_954);
xnor U7 (N_7,In_846,In_1123);
and U8 (N_8,In_23,In_622);
or U9 (N_9,In_1293,In_1305);
nand U10 (N_10,In_1328,In_1028);
or U11 (N_11,In_1790,In_1589);
and U12 (N_12,In_523,In_144);
xor U13 (N_13,In_1247,In_810);
nand U14 (N_14,In_1725,In_1822);
and U15 (N_15,In_1040,In_129);
xor U16 (N_16,In_75,In_901);
nor U17 (N_17,In_1948,In_1343);
xnor U18 (N_18,In_1041,In_609);
nor U19 (N_19,In_1601,In_1435);
nor U20 (N_20,In_1508,In_227);
nand U21 (N_21,In_564,In_1715);
or U22 (N_22,In_790,In_1570);
xnor U23 (N_23,In_911,In_1905);
nand U24 (N_24,In_192,In_442);
or U25 (N_25,In_826,In_670);
xor U26 (N_26,In_408,In_1067);
nand U27 (N_27,In_516,In_1194);
or U28 (N_28,In_1654,In_81);
or U29 (N_29,In_514,In_1134);
xnor U30 (N_30,In_813,In_1494);
nand U31 (N_31,In_511,In_79);
nor U32 (N_32,In_1327,In_356);
nor U33 (N_33,In_197,In_279);
xnor U34 (N_34,In_821,In_369);
nand U35 (N_35,In_67,In_1989);
xnor U36 (N_36,In_1257,In_1088);
and U37 (N_37,In_1484,In_921);
nand U38 (N_38,In_1597,In_1277);
and U39 (N_39,In_1021,In_1395);
or U40 (N_40,In_215,In_1380);
nand U41 (N_41,In_1083,In_313);
and U42 (N_42,In_534,In_1441);
and U43 (N_43,In_684,In_1979);
nor U44 (N_44,In_449,In_709);
xnor U45 (N_45,In_865,In_1121);
nand U46 (N_46,In_1048,In_802);
and U47 (N_47,In_1396,In_988);
nand U48 (N_48,In_1735,In_1263);
nor U49 (N_49,In_1741,In_245);
and U50 (N_50,In_1865,In_1094);
xnor U51 (N_51,In_1424,In_879);
xnor U52 (N_52,In_1829,In_760);
nand U53 (N_53,In_693,In_384);
xor U54 (N_54,In_1667,In_655);
or U55 (N_55,In_460,In_1950);
nand U56 (N_56,In_509,In_1959);
xor U57 (N_57,In_1283,In_1353);
or U58 (N_58,In_397,In_1181);
xnor U59 (N_59,In_1931,In_1128);
nor U60 (N_60,In_930,In_413);
nand U61 (N_61,In_257,In_340);
nand U62 (N_62,In_515,In_1818);
xnor U63 (N_63,In_170,In_1086);
or U64 (N_64,In_36,In_1779);
and U65 (N_65,In_521,In_1666);
nor U66 (N_66,In_47,In_1981);
nor U67 (N_67,In_194,In_1440);
and U68 (N_68,In_737,In_1944);
nand U69 (N_69,In_959,In_951);
xnor U70 (N_70,In_1633,In_1275);
or U71 (N_71,In_1534,In_1924);
and U72 (N_72,In_1858,In_722);
xor U73 (N_73,In_1744,In_1334);
and U74 (N_74,In_230,In_344);
or U75 (N_75,In_1348,In_159);
or U76 (N_76,In_816,In_873);
xnor U77 (N_77,In_1005,In_763);
nand U78 (N_78,In_1600,In_309);
or U79 (N_79,In_156,In_1156);
nand U80 (N_80,In_1186,In_1155);
nand U81 (N_81,In_698,In_755);
nand U82 (N_82,In_68,In_1302);
xnor U83 (N_83,In_314,In_1296);
and U84 (N_84,In_100,In_1444);
or U85 (N_85,In_610,In_654);
and U86 (N_86,In_1388,In_1862);
nor U87 (N_87,In_1465,In_961);
and U88 (N_88,In_455,In_207);
or U89 (N_89,In_1996,In_316);
or U90 (N_90,In_782,In_64);
or U91 (N_91,In_945,In_537);
nand U92 (N_92,In_1197,In_643);
and U93 (N_93,In_1065,In_1970);
and U94 (N_94,In_371,In_910);
nand U95 (N_95,In_172,In_1462);
xor U96 (N_96,In_1482,In_1825);
nor U97 (N_97,In_1140,In_342);
and U98 (N_98,In_10,In_1179);
and U99 (N_99,In_1177,In_1908);
and U100 (N_100,In_273,In_1527);
xnor U101 (N_101,In_493,In_1798);
nand U102 (N_102,In_1234,In_1244);
xor U103 (N_103,In_1430,In_382);
or U104 (N_104,In_1382,In_1501);
or U105 (N_105,In_1524,In_386);
and U106 (N_106,In_780,In_1833);
or U107 (N_107,In_554,In_1493);
nor U108 (N_108,In_201,In_1469);
and U109 (N_109,In_948,In_541);
xnor U110 (N_110,In_1774,In_1376);
xor U111 (N_111,In_896,In_1621);
and U112 (N_112,In_398,In_1605);
nor U113 (N_113,In_1696,In_1112);
xor U114 (N_114,In_1405,In_1739);
and U115 (N_115,In_1457,In_204);
nand U116 (N_116,In_292,In_1125);
nand U117 (N_117,In_1685,In_1285);
or U118 (N_118,In_1515,In_823);
or U119 (N_119,In_1588,In_869);
nand U120 (N_120,In_40,In_1695);
nand U121 (N_121,In_1902,In_1985);
xnor U122 (N_122,In_805,In_1892);
xnor U123 (N_123,In_119,In_1066);
or U124 (N_124,In_984,In_1129);
nor U125 (N_125,In_1884,In_558);
and U126 (N_126,In_1315,In_387);
and U127 (N_127,In_1168,In_1879);
and U128 (N_128,In_1437,In_1332);
nor U129 (N_129,In_738,In_551);
nand U130 (N_130,In_1310,In_1982);
nor U131 (N_131,In_918,In_220);
nand U132 (N_132,In_1472,In_1544);
xor U133 (N_133,In_1414,In_19);
and U134 (N_134,In_1461,In_169);
or U135 (N_135,In_1312,In_97);
and U136 (N_136,In_280,In_1075);
nand U137 (N_137,In_1220,In_797);
xor U138 (N_138,In_839,In_1942);
nor U139 (N_139,In_756,In_745);
xor U140 (N_140,In_568,In_1215);
xnor U141 (N_141,In_1308,In_593);
nor U142 (N_142,In_1650,In_1370);
or U143 (N_143,In_117,In_716);
nand U144 (N_144,In_195,In_1887);
xnor U145 (N_145,In_664,In_13);
nand U146 (N_146,In_689,In_383);
and U147 (N_147,In_781,In_1624);
nand U148 (N_148,In_456,In_1772);
or U149 (N_149,In_65,In_545);
xnor U150 (N_150,In_1513,In_1039);
or U151 (N_151,In_591,In_1620);
or U152 (N_152,In_672,In_242);
and U153 (N_153,In_697,In_499);
nand U154 (N_154,In_0,In_1590);
or U155 (N_155,In_1191,In_1669);
nand U156 (N_156,In_1585,In_206);
and U157 (N_157,In_553,In_1612);
or U158 (N_158,In_140,In_601);
xnor U159 (N_159,In_1299,In_1204);
nand U160 (N_160,In_1093,In_1945);
and U161 (N_161,In_407,In_877);
xnor U162 (N_162,In_193,In_586);
and U163 (N_163,In_86,In_1517);
xnor U164 (N_164,In_1239,In_620);
nand U165 (N_165,In_1398,In_187);
and U166 (N_166,In_892,In_1660);
or U167 (N_167,In_1952,In_1602);
or U168 (N_168,In_1294,In_106);
nand U169 (N_169,In_787,In_611);
nor U170 (N_170,In_239,In_329);
nor U171 (N_171,In_641,In_368);
and U172 (N_172,In_1680,In_45);
xor U173 (N_173,In_246,In_476);
or U174 (N_174,In_1915,In_1937);
nand U175 (N_175,In_1341,In_1736);
or U176 (N_176,In_1815,In_1577);
and U177 (N_177,In_1977,In_1885);
and U178 (N_178,In_1167,In_175);
and U179 (N_179,In_1166,In_1111);
nor U180 (N_180,In_158,In_902);
nor U181 (N_181,In_1711,In_54);
or U182 (N_182,In_1831,In_1843);
or U183 (N_183,In_505,In_1848);
nor U184 (N_184,In_811,In_1228);
nor U185 (N_185,In_478,In_1158);
and U186 (N_186,In_1356,In_349);
xor U187 (N_187,In_647,In_288);
nand U188 (N_188,In_615,In_862);
nand U189 (N_189,In_1209,In_1360);
nand U190 (N_190,In_148,In_1781);
and U191 (N_191,In_830,In_1786);
and U192 (N_192,In_72,In_1704);
or U193 (N_193,In_269,In_1903);
xnor U194 (N_194,In_444,In_1639);
xor U195 (N_195,In_1288,In_366);
or U196 (N_196,In_575,In_1292);
and U197 (N_197,In_1886,In_583);
or U198 (N_198,In_1809,In_223);
nand U199 (N_199,In_947,In_603);
nor U200 (N_200,In_228,In_218);
and U201 (N_201,In_1897,In_1147);
or U202 (N_202,In_1502,In_640);
xnor U203 (N_203,In_1619,In_326);
xnor U204 (N_204,In_138,In_38);
and U205 (N_205,In_1301,In_1773);
or U206 (N_206,In_1983,In_1738);
or U207 (N_207,In_427,In_1384);
xnor U208 (N_208,In_364,In_893);
or U209 (N_209,In_39,In_1895);
nor U210 (N_210,In_888,In_799);
xnor U211 (N_211,In_999,In_149);
xor U212 (N_212,In_1801,In_713);
and U213 (N_213,In_1900,In_717);
and U214 (N_214,In_1904,In_1463);
or U215 (N_215,In_1592,In_467);
and U216 (N_216,In_1586,In_1323);
nor U217 (N_217,In_1306,In_1518);
nand U218 (N_218,In_1810,In_957);
xor U219 (N_219,In_435,In_1684);
or U220 (N_220,In_1928,In_663);
nor U221 (N_221,In_3,In_491);
or U222 (N_222,In_994,In_52);
nor U223 (N_223,In_981,In_768);
xor U224 (N_224,In_1916,In_1161);
nor U225 (N_225,In_1603,In_1813);
or U226 (N_226,In_949,In_1598);
and U227 (N_227,In_916,In_152);
xor U228 (N_228,In_1714,In_1662);
nand U229 (N_229,In_474,In_1421);
nand U230 (N_230,In_264,In_84);
or U231 (N_231,In_1631,In_1117);
and U232 (N_232,In_1847,In_1002);
nor U233 (N_233,In_750,In_437);
nand U234 (N_234,In_282,In_141);
and U235 (N_235,In_1805,In_844);
nor U236 (N_236,In_1836,In_154);
or U237 (N_237,In_325,In_1901);
and U238 (N_238,In_182,In_662);
nand U239 (N_239,In_803,In_1731);
nand U240 (N_240,In_391,In_847);
or U241 (N_241,In_319,In_1271);
xor U242 (N_242,In_1236,In_931);
nand U243 (N_243,In_868,In_1426);
and U244 (N_244,In_1372,In_446);
nor U245 (N_245,In_1648,In_1274);
or U246 (N_246,In_986,In_1876);
xnor U247 (N_247,In_617,In_898);
xnor U248 (N_248,In_644,In_645);
or U249 (N_249,In_673,In_1797);
and U250 (N_250,In_423,In_914);
nand U251 (N_251,In_347,In_1113);
and U252 (N_252,In_725,In_1890);
and U253 (N_253,In_606,In_1450);
xor U254 (N_254,In_142,In_770);
xor U255 (N_255,In_832,In_1460);
or U256 (N_256,In_1860,In_17);
or U257 (N_257,In_825,In_2);
nand U258 (N_258,In_607,In_1336);
xnor U259 (N_259,In_69,In_1403);
nand U260 (N_260,In_743,In_146);
and U261 (N_261,In_426,In_815);
and U262 (N_262,In_619,In_1536);
nand U263 (N_263,In_430,In_1057);
nand U264 (N_264,In_199,In_639);
nor U265 (N_265,In_585,In_135);
and U266 (N_266,In_1674,In_1304);
nand U267 (N_267,In_1286,In_623);
and U268 (N_268,In_590,In_1377);
nor U269 (N_269,In_1087,In_831);
xnor U270 (N_270,In_1587,In_1750);
or U271 (N_271,In_932,In_1175);
or U272 (N_272,In_963,In_1663);
xor U273 (N_273,In_1988,In_1214);
or U274 (N_274,In_1,In_300);
xnor U275 (N_275,In_1203,In_1682);
xnor U276 (N_276,In_1029,In_1474);
and U277 (N_277,In_1237,In_1510);
nor U278 (N_278,In_22,In_1069);
xnor U279 (N_279,In_127,In_1867);
nor U280 (N_280,In_1871,In_1807);
xnor U281 (N_281,In_454,In_1975);
and U282 (N_282,In_286,In_728);
nor U283 (N_283,In_1498,In_1742);
nand U284 (N_284,In_489,In_1845);
or U285 (N_285,In_1347,In_1999);
or U286 (N_286,In_1011,In_1497);
nand U287 (N_287,In_565,In_1153);
xor U288 (N_288,In_1165,In_73);
nand U289 (N_289,In_637,In_312);
xor U290 (N_290,In_51,In_633);
xor U291 (N_291,In_1701,In_1261);
nand U292 (N_292,In_1634,In_938);
xor U293 (N_293,In_628,In_1023);
xnor U294 (N_294,In_501,In_561);
or U295 (N_295,In_295,In_120);
or U296 (N_296,In_299,In_979);
and U297 (N_297,In_451,In_1507);
nor U298 (N_298,In_1138,In_1046);
xor U299 (N_299,In_604,In_1995);
nand U300 (N_300,In_504,In_379);
nor U301 (N_301,In_1986,In_539);
nand U302 (N_302,In_870,In_1231);
nor U303 (N_303,In_462,In_718);
and U304 (N_304,In_1967,In_483);
and U305 (N_305,In_967,In_710);
xor U306 (N_306,In_87,In_1914);
or U307 (N_307,In_1647,In_1008);
and U308 (N_308,In_362,In_46);
nor U309 (N_309,In_1616,In_166);
nand U310 (N_310,In_145,In_1530);
nand U311 (N_311,In_765,In_1757);
xnor U312 (N_312,In_231,In_878);
nor U313 (N_313,In_1572,In_212);
xor U314 (N_314,In_91,In_298);
and U315 (N_315,In_1922,In_438);
and U316 (N_316,In_857,In_1216);
nand U317 (N_317,In_440,In_1664);
nor U318 (N_318,In_1358,In_581);
xnor U319 (N_319,In_1595,In_107);
nand U320 (N_320,In_1939,In_1596);
xor U321 (N_321,In_167,In_675);
nor U322 (N_322,In_1042,In_1406);
and U323 (N_323,In_1351,In_528);
nor U324 (N_324,In_1980,In_1103);
or U325 (N_325,In_1099,In_1084);
nand U326 (N_326,In_283,In_1868);
and U327 (N_327,In_1455,In_112);
xnor U328 (N_328,In_432,In_1092);
or U329 (N_329,In_691,In_1415);
or U330 (N_330,In_1137,In_1635);
nor U331 (N_331,In_327,In_1264);
nor U332 (N_332,In_1339,In_646);
nor U333 (N_333,In_1297,In_776);
nor U334 (N_334,In_1157,In_85);
or U335 (N_335,In_479,In_1917);
nand U336 (N_336,In_758,In_1911);
or U337 (N_337,In_1340,In_572);
or U338 (N_338,In_1309,In_736);
xor U339 (N_339,In_306,In_1268);
or U340 (N_340,In_346,In_1559);
nand U341 (N_341,In_184,In_48);
and U342 (N_342,In_742,In_111);
nand U343 (N_343,In_1454,In_102);
and U344 (N_344,In_57,In_1599);
and U345 (N_345,In_304,In_354);
nand U346 (N_346,In_946,In_835);
and U347 (N_347,In_828,In_801);
nand U348 (N_348,In_1333,In_1737);
nor U349 (N_349,In_1245,In_1734);
xor U350 (N_350,In_1072,In_214);
nand U351 (N_351,In_176,In_1227);
and U352 (N_352,In_1218,In_1320);
nand U353 (N_353,In_348,In_1907);
nor U354 (N_354,In_1748,In_1196);
and U355 (N_355,In_248,In_66);
and U356 (N_356,In_1819,In_1107);
nor U357 (N_357,In_1483,In_1016);
and U358 (N_358,In_58,In_1089);
xnor U359 (N_359,In_1976,In_1840);
nand U360 (N_360,In_566,In_1608);
nand U361 (N_361,In_50,In_1091);
or U362 (N_362,In_1255,In_263);
xor U363 (N_363,In_114,In_671);
and U364 (N_364,In_864,In_1105);
and U365 (N_365,In_1477,In_793);
nor U366 (N_366,In_711,In_1037);
and U367 (N_367,In_1566,In_1992);
or U368 (N_368,In_1538,In_1373);
nor U369 (N_369,In_4,In_1529);
nand U370 (N_370,In_1971,In_137);
and U371 (N_371,In_1679,In_587);
nand U372 (N_372,In_1861,In_1452);
xnor U373 (N_373,In_472,In_1883);
and U374 (N_374,In_1064,In_1512);
nand U375 (N_375,In_1543,In_1875);
and U376 (N_376,In_1411,In_1390);
and U377 (N_377,In_470,In_1473);
xor U378 (N_378,In_1230,In_1240);
and U379 (N_379,In_1694,In_1703);
or U380 (N_380,In_1488,In_638);
nor U381 (N_381,In_1569,In_769);
nor U382 (N_382,In_1611,In_418);
nand U383 (N_383,In_412,In_1496);
nand U384 (N_384,In_1519,In_1198);
or U385 (N_385,In_1522,In_543);
xor U386 (N_386,In_332,In_1389);
nand U387 (N_387,In_929,In_1726);
or U388 (N_388,In_1906,In_1055);
nand U389 (N_389,In_351,In_953);
and U390 (N_390,In_126,In_420);
nand U391 (N_391,In_1854,In_399);
or U392 (N_392,In_1141,In_1765);
or U393 (N_393,In_56,In_496);
nand U394 (N_394,In_1525,In_773);
nor U395 (N_395,In_507,In_1957);
or U396 (N_396,In_1514,In_1202);
nand U397 (N_397,In_139,In_1638);
or U398 (N_398,In_840,In_250);
and U399 (N_399,In_563,In_1706);
nor U400 (N_400,In_1571,In_1943);
and U401 (N_401,In_1280,In_482);
nand U402 (N_402,In_1248,In_850);
nor U403 (N_403,In_365,In_1821);
nand U404 (N_404,In_1187,In_520);
xor U405 (N_405,In_1321,In_287);
or U406 (N_406,In_705,In_272);
nor U407 (N_407,In_855,In_612);
xnor U408 (N_408,In_1180,In_400);
nor U409 (N_409,In_1031,In_1689);
nand U410 (N_410,In_132,In_277);
nand U411 (N_411,In_1764,In_1082);
or U412 (N_412,In_1762,In_634);
nand U413 (N_413,In_99,In_903);
nand U414 (N_414,In_1934,In_178);
nand U415 (N_415,In_77,In_682);
nand U416 (N_416,In_436,In_853);
nand U417 (N_417,In_475,In_627);
xnor U418 (N_418,In_1794,In_1575);
or U419 (N_419,In_996,In_1563);
xor U420 (N_420,In_330,In_721);
or U421 (N_421,In_1729,In_1273);
xor U422 (N_422,In_1788,In_393);
nor U423 (N_423,In_343,In_1659);
or U424 (N_424,In_274,In_60);
and U425 (N_425,In_123,In_1787);
nor U426 (N_426,In_1832,In_307);
and U427 (N_427,In_1447,In_1713);
and U428 (N_428,In_1789,In_536);
and U429 (N_429,In_1213,In_410);
nand U430 (N_430,In_334,In_355);
xnor U431 (N_431,In_922,In_1724);
or U432 (N_432,In_1470,In_42);
and U433 (N_433,In_527,In_130);
xnor U434 (N_434,In_1552,In_151);
nand U435 (N_435,In_1010,In_876);
nand U436 (N_436,In_724,In_1556);
and U437 (N_437,In_920,In_1668);
nor U438 (N_438,In_1035,In_1051);
xnor U439 (N_439,In_179,In_122);
nor U440 (N_440,In_1325,In_836);
and U441 (N_441,In_1034,In_1708);
nor U442 (N_442,In_669,In_1265);
nor U443 (N_443,In_210,In_510);
or U444 (N_444,In_301,In_1256);
or U445 (N_445,In_764,In_1785);
and U446 (N_446,In_16,In_328);
nor U447 (N_447,In_1387,In_1352);
nand U448 (N_448,In_1258,In_222);
xor U449 (N_449,In_933,In_608);
or U450 (N_450,In_1160,In_1718);
nor U451 (N_451,In_1221,In_1758);
nor U452 (N_452,In_213,In_1752);
and U453 (N_453,In_1835,In_522);
or U454 (N_454,In_977,In_837);
and U455 (N_455,In_422,In_1200);
xnor U456 (N_456,In_1410,In_271);
xnor U457 (N_457,In_18,In_1173);
nand U458 (N_458,In_950,In_1281);
or U459 (N_459,In_927,In_784);
nor U460 (N_460,In_98,In_550);
nand U461 (N_461,In_829,In_1878);
or U462 (N_462,In_1812,In_1973);
and U463 (N_463,In_919,In_1386);
nand U464 (N_464,In_968,In_25);
nand U465 (N_465,In_1607,In_1109);
nor U466 (N_466,In_1178,In_1238);
or U467 (N_467,In_991,In_1657);
nor U468 (N_468,In_1471,In_1972);
and U469 (N_469,In_838,In_733);
or U470 (N_470,In_502,In_1467);
or U471 (N_471,In_956,In_1580);
nand U472 (N_472,In_1243,In_310);
nand U473 (N_473,In_1290,In_96);
and U474 (N_474,In_1350,In_59);
nor U475 (N_475,In_1661,In_648);
nor U476 (N_476,In_353,In_1375);
xnor U477 (N_477,In_1541,In_1849);
nand U478 (N_478,In_1012,In_409);
and U479 (N_479,In_208,In_785);
nand U480 (N_480,In_1349,In_1394);
or U481 (N_481,In_1850,In_741);
nor U482 (N_482,In_1442,In_1740);
nand U483 (N_483,In_155,In_602);
and U484 (N_484,In_798,In_1984);
nor U485 (N_485,In_1188,In_1941);
xor U486 (N_486,In_1054,In_1059);
xnor U487 (N_487,In_1015,In_27);
or U488 (N_488,In_1030,In_1964);
nor U489 (N_489,In_1688,In_1131);
xor U490 (N_490,In_338,In_1013);
nor U491 (N_491,In_1232,In_1716);
nand U492 (N_492,In_1374,In_302);
and U493 (N_493,In_266,In_93);
or U494 (N_494,In_621,In_969);
and U495 (N_495,In_487,In_1136);
nor U496 (N_496,In_1551,In_1401);
or U497 (N_497,In_492,In_1225);
nor U498 (N_498,In_1475,In_196);
nor U499 (N_499,In_1017,In_985);
nand U500 (N_500,In_392,In_1260);
xor U501 (N_501,In_820,In_719);
nand U502 (N_502,In_1485,In_78);
nand U503 (N_503,In_1182,In_1043);
or U504 (N_504,In_1272,In_906);
and U505 (N_505,In_1045,In_1342);
and U506 (N_506,In_1110,In_458);
nand U507 (N_507,In_1007,In_95);
xnor U508 (N_508,In_6,In_1079);
and U509 (N_509,In_157,In_1114);
or U510 (N_510,In_1656,In_1951);
nor U511 (N_511,In_225,In_1298);
xor U512 (N_512,In_359,In_1024);
xnor U513 (N_513,In_429,In_817);
nand U514 (N_514,In_229,In_529);
or U515 (N_515,In_656,In_1459);
xnor U516 (N_516,In_859,In_715);
xnor U517 (N_517,In_1617,In_1640);
xor U518 (N_518,In_1126,In_296);
and U519 (N_519,In_419,In_308);
nor U520 (N_520,In_305,In_1036);
xnor U521 (N_521,In_935,In_1211);
xor U522 (N_522,In_1687,In_582);
or U523 (N_523,In_477,In_1927);
nor U524 (N_524,In_244,In_727);
and U525 (N_525,In_1262,In_136);
or U526 (N_526,In_1116,In_1683);
nor U527 (N_527,In_291,In_1965);
and U528 (N_528,In_1503,In_1383);
xnor U529 (N_529,In_588,In_1677);
nor U530 (N_530,In_1670,In_162);
or U531 (N_531,In_1727,In_1404);
nor U532 (N_532,In_260,In_806);
nor U533 (N_533,In_1783,In_1270);
xnor U534 (N_534,In_254,In_540);
xor U535 (N_535,In_908,In_1555);
and U536 (N_536,In_448,In_1532);
or U537 (N_537,In_1705,In_453);
nor U538 (N_538,In_1314,In_989);
and U539 (N_539,In_345,In_1672);
and U540 (N_540,In_500,In_76);
or U541 (N_541,In_1642,In_404);
xnor U542 (N_542,In_983,In_1335);
xor U543 (N_543,In_1814,In_433);
xor U544 (N_544,In_1000,In_777);
xor U545 (N_545,In_595,In_90);
and U546 (N_546,In_598,In_1195);
nor U547 (N_547,In_490,In_1080);
nor U548 (N_548,In_1919,In_1623);
nand U549 (N_549,In_219,In_1506);
nand U550 (N_550,In_614,In_1267);
nor U551 (N_551,In_1052,In_1963);
nand U552 (N_552,In_415,In_960);
nor U553 (N_553,In_597,In_324);
nand U554 (N_554,In_224,In_134);
nor U555 (N_555,In_1629,In_1212);
xor U556 (N_556,In_1673,In_11);
and U557 (N_557,In_1795,In_1918);
xor U558 (N_558,In_1154,In_1330);
nor U559 (N_559,In_105,In_1085);
xnor U560 (N_560,In_1826,In_401);
nor U561 (N_561,In_1478,In_70);
and U562 (N_562,In_971,In_512);
nor U563 (N_563,In_778,In_1889);
xor U564 (N_564,In_1210,In_485);
nand U565 (N_565,In_913,In_1722);
and U566 (N_566,In_1163,In_1505);
xnor U567 (N_567,In_757,In_783);
and U568 (N_568,In_885,In_1949);
nand U569 (N_569,In_1542,In_941);
nor U570 (N_570,In_1144,In_600);
nand U571 (N_571,In_1593,In_1993);
and U572 (N_572,In_1645,In_924);
nand U573 (N_573,In_1003,In_538);
or U574 (N_574,In_1775,In_992);
nor U575 (N_575,In_936,In_642);
xor U576 (N_576,In_71,In_1800);
or U577 (N_577,In_1828,In_164);
nand U578 (N_578,In_1834,In_270);
nand U579 (N_579,In_1254,In_1974);
nor U580 (N_580,In_1096,In_1869);
xor U581 (N_581,In_1533,In_278);
nand U582 (N_582,In_377,In_1499);
and U583 (N_583,In_982,In_1958);
nor U584 (N_584,In_706,In_1449);
or U585 (N_585,In_1357,In_1978);
nand U586 (N_586,In_767,In_494);
or U587 (N_587,In_1468,In_1712);
nor U588 (N_588,In_1108,In_1863);
nor U589 (N_589,In_1063,In_676);
nand U590 (N_590,In_74,In_221);
or U591 (N_591,In_1521,In_526);
and U592 (N_592,In_1466,In_1489);
and U593 (N_593,In_357,In_209);
and U594 (N_594,In_1303,In_378);
nand U595 (N_595,In_584,In_411);
or U596 (N_596,In_488,In_276);
nand U597 (N_597,In_174,In_995);
xor U598 (N_598,In_557,In_1207);
or U599 (N_599,In_1956,In_375);
and U600 (N_600,In_211,In_874);
nor U601 (N_601,In_1751,In_952);
or U602 (N_602,In_1830,In_1899);
nor U603 (N_603,In_653,In_15);
nor U604 (N_604,In_1913,In_687);
nand U605 (N_605,In_1106,In_447);
and U606 (N_606,In_1183,In_605);
and U607 (N_607,In_1448,In_1893);
or U608 (N_608,In_1933,In_1720);
and U609 (N_609,In_791,In_1135);
xnor U610 (N_610,In_1700,In_1322);
and U611 (N_611,In_1691,In_942);
and U612 (N_612,In_1528,In_1282);
nor U613 (N_613,In_525,In_1289);
or U614 (N_614,In_1678,In_940);
nor U615 (N_615,In_1486,In_484);
or U616 (N_616,In_580,In_1119);
nand U617 (N_617,In_281,In_1778);
nand U618 (N_618,In_1759,In_1618);
xnor U619 (N_619,In_531,In_1614);
and U620 (N_620,In_1423,In_104);
nand U621 (N_621,In_1033,In_1431);
nor U622 (N_622,In_665,In_1846);
nor U623 (N_623,In_822,In_265);
nand U624 (N_624,In_116,In_1641);
and U625 (N_625,In_1269,In_970);
or U626 (N_626,In_1445,In_624);
nand U627 (N_627,In_1081,In_1791);
and U628 (N_628,In_1480,In_883);
nand U629 (N_629,In_237,In_1504);
xor U630 (N_630,In_1643,In_1938);
and U631 (N_631,In_1756,In_1553);
and U632 (N_632,In_559,In_1511);
or U633 (N_633,In_943,In_1500);
xor U634 (N_634,In_895,In_1784);
or U635 (N_635,In_1338,In_94);
nand U636 (N_636,In_1874,In_1095);
nand U637 (N_637,In_897,In_1337);
or U638 (N_638,In_1050,In_1076);
or U639 (N_639,In_1409,In_690);
xnor U640 (N_640,In_1573,In_1246);
xnor U641 (N_641,In_792,In_181);
nand U642 (N_642,In_915,In_1381);
or U643 (N_643,In_1581,In_761);
nand U644 (N_644,In_1561,In_53);
nor U645 (N_645,In_1433,In_1190);
nor U646 (N_646,In_1888,In_576);
nor U647 (N_647,In_632,In_318);
or U648 (N_648,In_1562,In_866);
nor U649 (N_649,In_1760,In_1418);
nand U650 (N_650,In_1331,In_421);
nor U651 (N_651,In_1222,In_373);
xnor U652 (N_652,In_498,In_1291);
xor U653 (N_653,In_35,In_1413);
nor U654 (N_654,In_1582,In_1393);
nand U655 (N_655,In_49,In_459);
xnor U656 (N_656,In_1920,In_1780);
nand U657 (N_657,In_546,In_1090);
xnor U658 (N_658,In_468,In_789);
or U659 (N_659,In_198,In_1921);
nand U660 (N_660,In_1019,In_1189);
and U661 (N_661,In_171,In_701);
xor U662 (N_662,In_683,In_1960);
and U663 (N_663,In_962,In_30);
xor U664 (N_664,In_461,In_1806);
xnor U665 (N_665,In_1329,In_1546);
nand U666 (N_666,In_863,In_1481);
or U667 (N_667,In_1652,In_434);
and U668 (N_668,In_720,In_26);
xnor U669 (N_669,In_1378,In_1692);
nand U670 (N_670,In_8,In_907);
xnor U671 (N_671,In_650,In_150);
nand U672 (N_672,In_1853,In_1702);
xnor U673 (N_673,In_293,In_367);
xor U674 (N_674,In_723,In_255);
xnor U675 (N_675,In_997,In_1150);
nand U676 (N_676,In_771,In_1811);
nor U677 (N_677,In_751,In_707);
nor U678 (N_678,In_463,In_341);
xnor U679 (N_679,In_794,In_1022);
or U680 (N_680,In_358,In_1910);
and U681 (N_681,In_14,In_851);
and U682 (N_682,In_571,In_1369);
nand U683 (N_683,In_1768,In_1206);
and U684 (N_684,In_44,In_1870);
or U685 (N_685,In_731,In_1615);
xnor U686 (N_686,In_1730,In_1632);
xnor U687 (N_687,In_1074,In_1266);
nand U688 (N_688,In_1078,In_966);
nor U689 (N_689,In_1891,In_1162);
and U690 (N_690,In_856,In_1199);
nor U691 (N_691,In_625,In_1531);
xnor U692 (N_692,In_1583,In_1955);
and U693 (N_693,In_1032,In_1935);
xor U694 (N_694,In_1749,In_795);
xnor U695 (N_695,In_389,In_1056);
nor U696 (N_696,In_1159,In_904);
or U697 (N_697,In_854,In_256);
and U698 (N_698,In_659,In_216);
xor U699 (N_699,In_1509,In_891);
nand U700 (N_700,In_1319,In_1193);
nand U701 (N_701,In_804,In_41);
xnor U702 (N_702,In_1792,In_1276);
nor U703 (N_703,In_188,In_578);
nand U704 (N_704,In_1295,In_1565);
and U705 (N_705,In_131,In_1962);
xnor U706 (N_706,In_833,In_695);
or U707 (N_707,In_1491,In_1873);
nand U708 (N_708,In_160,In_268);
and U709 (N_709,In_20,In_320);
xor U710 (N_710,In_189,In_1115);
nor U711 (N_711,In_964,In_1604);
xor U712 (N_712,In_61,In_699);
nor U713 (N_713,In_978,In_143);
nand U714 (N_714,In_1560,In_1776);
nand U715 (N_715,In_1646,In_1130);
xnor U716 (N_716,In_1422,In_1058);
xnor U717 (N_717,In_376,In_1550);
and U718 (N_718,In_944,In_1866);
nor U719 (N_719,In_331,In_1001);
nand U720 (N_720,In_360,In_1606);
xor U721 (N_721,In_657,In_200);
nor U722 (N_722,In_958,In_1576);
or U723 (N_723,In_1665,In_616);
nor U724 (N_724,In_1539,In_747);
nand U725 (N_725,In_7,In_1490);
nor U726 (N_726,In_1655,In_1930);
xnor U727 (N_727,In_147,In_1808);
or U728 (N_728,In_1676,In_635);
and U729 (N_729,In_703,In_800);
xnor U730 (N_730,In_1824,In_1747);
and U731 (N_731,In_1287,In_652);
xor U732 (N_732,In_297,In_702);
nor U733 (N_733,In_681,In_555);
or U734 (N_734,In_1020,In_1940);
xnor U735 (N_735,In_5,In_577);
xnor U736 (N_736,In_1120,In_1249);
nor U737 (N_737,In_1717,In_1070);
nand U738 (N_738,In_374,In_1049);
nor U739 (N_739,In_1362,In_1763);
xor U740 (N_740,In_1365,In_1613);
nor U741 (N_741,In_1894,In_1419);
nand U742 (N_742,In_1151,In_1841);
xnor U743 (N_743,In_235,In_1379);
or U744 (N_744,In_708,In_1233);
or U745 (N_745,In_1753,In_1436);
xor U746 (N_746,In_1487,In_92);
or U747 (N_747,In_688,In_1427);
xor U748 (N_748,In_180,In_109);
nand U749 (N_749,In_1719,In_284);
nand U750 (N_750,In_524,In_1367);
and U751 (N_751,In_101,In_814);
or U752 (N_752,In_1966,In_80);
nor U753 (N_753,In_1728,In_834);
nor U754 (N_754,In_1578,In_1279);
nand U755 (N_755,In_173,In_1361);
nand U756 (N_756,In_579,In_1761);
nand U757 (N_757,In_323,In_1241);
and U758 (N_758,In_1912,In_1251);
nand U759 (N_759,In_480,In_1516);
or U760 (N_760,In_858,In_1877);
or U761 (N_761,In_1252,In_226);
nor U762 (N_762,In_1609,In_517);
nand U763 (N_763,In_827,In_1098);
nor U764 (N_764,In_1743,In_183);
and U765 (N_765,In_253,In_1535);
and U766 (N_766,In_1969,In_118);
and U767 (N_767,In_1548,In_1408);
xor U768 (N_768,In_1707,In_618);
nor U769 (N_769,In_396,In_1185);
nand U770 (N_770,In_766,In_370);
nor U771 (N_771,In_465,In_352);
nand U772 (N_772,In_841,In_441);
xnor U773 (N_773,In_1675,In_1458);
nor U774 (N_774,In_849,In_1495);
nand U775 (N_775,In_466,In_1880);
or U776 (N_776,In_808,In_1420);
xnor U777 (N_777,In_1438,In_1060);
nor U778 (N_778,In_875,In_730);
nand U779 (N_779,In_1026,In_113);
and U780 (N_780,In_1453,In_243);
xnor U781 (N_781,In_955,In_450);
nor U782 (N_782,In_1681,In_232);
or U783 (N_783,In_735,In_1721);
xnor U784 (N_784,In_177,In_124);
or U785 (N_785,In_1397,In_1837);
nand U786 (N_786,In_335,In_1782);
nand U787 (N_787,In_1412,In_1823);
nand U788 (N_788,In_1793,In_1104);
xor U789 (N_789,In_191,In_1014);
nand U790 (N_790,In_613,In_889);
nand U791 (N_791,In_1953,In_402);
xor U792 (N_792,In_1425,In_726);
nand U793 (N_793,In_110,In_573);
nand U794 (N_794,In_734,In_1804);
nor U795 (N_795,In_928,In_519);
nor U796 (N_796,In_1961,In_1402);
nor U797 (N_797,In_350,In_417);
nor U798 (N_798,In_1434,In_1146);
and U799 (N_799,In_679,In_1803);
or U800 (N_800,In_752,In_469);
nor U801 (N_801,In_694,In_1354);
xor U802 (N_802,In_202,In_1170);
and U803 (N_803,In_1355,In_457);
nor U804 (N_804,In_414,In_431);
nand U805 (N_805,In_547,In_473);
nor U806 (N_806,In_1307,In_1947);
and U807 (N_807,In_1537,In_275);
and U808 (N_808,In_464,In_1346);
and U809 (N_809,In_636,In_1284);
or U810 (N_810,In_678,In_1205);
nor U811 (N_811,In_486,In_508);
xnor U812 (N_812,In_363,In_1318);
and U813 (N_813,In_506,In_1610);
nor U814 (N_814,In_1027,In_497);
nor U815 (N_815,In_186,In_238);
xnor U816 (N_816,In_133,In_361);
or U817 (N_817,In_1407,In_32);
nand U818 (N_818,In_882,In_1368);
or U819 (N_819,In_1259,In_809);
nand U820 (N_820,In_1923,In_934);
nand U821 (N_821,In_1217,In_1127);
xnor U822 (N_822,In_163,In_1859);
xor U823 (N_823,In_900,In_1102);
and U824 (N_824,In_1557,In_886);
nor U825 (N_825,In_746,In_1936);
or U826 (N_826,In_1998,In_333);
and U827 (N_827,In_372,In_1132);
nand U828 (N_828,In_1658,In_1626);
and U829 (N_829,In_1451,In_205);
and U830 (N_830,In_533,In_692);
and U831 (N_831,In_887,In_1898);
or U832 (N_832,In_1686,In_880);
xor U833 (N_833,In_1754,In_1429);
nor U834 (N_834,In_685,In_1443);
or U835 (N_835,In_33,In_1523);
nor U836 (N_836,In_1311,In_649);
or U837 (N_837,In_1313,In_1201);
nand U838 (N_838,In_824,In_285);
nand U839 (N_839,In_852,In_1851);
nor U840 (N_840,In_1417,In_1636);
xor U841 (N_841,In_704,In_428);
nor U842 (N_842,In_416,In_128);
or U843 (N_843,In_899,In_818);
or U844 (N_844,In_1842,In_1077);
nand U845 (N_845,In_1479,In_1926);
and U846 (N_846,In_651,In_1242);
xnor U847 (N_847,In_1520,In_1896);
nor U848 (N_848,In_939,In_503);
xnor U849 (N_849,In_1839,In_1746);
and U850 (N_850,In_262,In_1997);
xnor U851 (N_851,In_1316,In_1038);
or U852 (N_852,In_28,In_165);
or U853 (N_853,In_55,In_674);
nand U854 (N_854,In_1549,In_714);
xnor U855 (N_855,In_403,In_965);
nand U856 (N_856,In_1061,In_1857);
nor U857 (N_857,In_1637,In_1827);
xor U858 (N_858,In_975,In_592);
nor U859 (N_859,In_1097,In_1476);
and U860 (N_860,In_1852,In_740);
xnor U861 (N_861,In_82,In_89);
and U862 (N_862,In_153,In_1071);
or U863 (N_863,In_884,In_115);
xor U864 (N_864,In_251,In_1526);
and U865 (N_865,In_443,In_912);
nor U866 (N_866,In_1994,In_290);
xnor U867 (N_867,In_240,In_43);
and U868 (N_868,In_532,In_311);
xnor U869 (N_869,In_629,In_1693);
and U870 (N_870,In_1699,In_1456);
nor U871 (N_871,In_1649,In_1991);
nand U872 (N_872,In_1838,In_1732);
and U873 (N_873,In_1817,In_1579);
or U874 (N_874,In_589,In_861);
nor U875 (N_875,In_748,In_185);
nor U876 (N_876,In_381,In_1968);
or U877 (N_877,In_596,In_1192);
or U878 (N_878,In_1690,In_917);
nor U879 (N_879,In_1133,In_1733);
nor U880 (N_880,In_405,In_9);
or U881 (N_881,In_923,In_495);
and U882 (N_882,In_1492,In_1300);
nand U883 (N_883,In_1439,In_303);
nor U884 (N_884,In_987,In_241);
xor U885 (N_885,In_445,In_1363);
nor U886 (N_886,In_258,In_1229);
xor U887 (N_887,In_812,In_1855);
and U888 (N_888,In_626,In_1006);
xnor U889 (N_889,In_542,In_1143);
xor U890 (N_890,In_696,In_1932);
xnor U891 (N_891,In_88,In_739);
nor U892 (N_892,In_1767,In_1142);
or U893 (N_893,In_1345,In_860);
or U894 (N_894,In_1872,In_322);
or U895 (N_895,In_1009,In_1796);
nand U896 (N_896,In_990,In_1253);
nand U897 (N_897,In_894,In_1545);
or U898 (N_898,In_549,In_1651);
or U899 (N_899,In_37,In_1584);
xnor U900 (N_900,In_394,In_1391);
nor U901 (N_901,In_630,In_1392);
nand U902 (N_902,In_774,In_1547);
nand U903 (N_903,In_1172,In_552);
and U904 (N_904,In_1428,In_1755);
or U905 (N_905,In_1062,In_1710);
nor U906 (N_906,In_925,In_819);
nand U907 (N_907,In_1644,In_890);
nor U908 (N_908,In_1399,In_1856);
or U909 (N_909,In_1653,In_594);
xor U910 (N_910,In_980,In_1777);
xnor U911 (N_911,In_779,In_1219);
xor U912 (N_912,In_631,In_12);
or U913 (N_913,In_1709,In_1324);
nand U914 (N_914,In_289,In_1124);
and U915 (N_915,In_807,In_471);
or U916 (N_916,In_24,In_772);
xnor U917 (N_917,In_660,In_1174);
nor U918 (N_918,In_1044,In_848);
xnor U919 (N_919,In_668,In_1464);
and U920 (N_920,In_530,In_1169);
nand U921 (N_921,In_686,In_974);
nand U922 (N_922,In_1371,In_1769);
nor U923 (N_923,In_700,In_1446);
xnor U924 (N_924,In_909,In_1591);
nor U925 (N_925,In_729,In_315);
nor U926 (N_926,In_1025,In_1625);
nor U927 (N_927,In_1400,In_998);
xnor U928 (N_928,In_390,In_321);
nand U929 (N_929,In_1164,In_843);
xor U930 (N_930,In_259,In_570);
nand U931 (N_931,In_217,In_518);
and U932 (N_932,In_1844,In_1366);
nand U933 (N_933,In_973,In_190);
nor U934 (N_934,In_439,In_775);
and U935 (N_935,In_1100,In_1047);
or U936 (N_936,In_976,In_21);
nand U937 (N_937,In_1364,In_388);
nand U938 (N_938,In_548,In_574);
or U939 (N_939,In_1148,In_63);
and U940 (N_940,In_1987,In_168);
xnor U941 (N_941,In_926,In_1627);
xnor U942 (N_942,In_867,In_1630);
xor U943 (N_943,In_233,In_249);
or U944 (N_944,In_1820,In_762);
xnor U945 (N_945,In_336,In_1567);
xnor U946 (N_946,In_1594,In_1568);
nor U947 (N_947,In_544,In_871);
or U948 (N_948,In_1073,In_234);
xor U949 (N_949,In_62,In_1925);
nor U950 (N_950,In_1816,In_1101);
nand U951 (N_951,In_666,In_1909);
xnor U952 (N_952,In_905,In_567);
and U953 (N_953,In_1223,In_1004);
nand U954 (N_954,In_1278,In_1118);
nor U955 (N_955,In_661,In_1317);
or U956 (N_956,In_1799,In_1139);
and U957 (N_957,In_1946,In_1235);
nor U958 (N_958,In_712,In_1250);
or U959 (N_959,In_1864,In_1990);
nand U960 (N_960,In_1385,In_796);
xnor U961 (N_961,In_261,In_1152);
xor U962 (N_962,In_1554,In_759);
xor U963 (N_963,In_247,In_1226);
and U964 (N_964,In_1745,In_972);
nor U965 (N_965,In_385,In_103);
nor U966 (N_966,In_1540,In_1053);
xor U967 (N_967,In_267,In_1881);
xor U968 (N_968,In_29,In_845);
nor U969 (N_969,In_121,In_1622);
xor U970 (N_970,In_1208,In_1574);
or U971 (N_971,In_753,In_744);
xnor U972 (N_972,In_1018,In_203);
and U973 (N_973,In_337,In_881);
xnor U974 (N_974,In_1628,In_560);
and U975 (N_975,In_31,In_1671);
nor U976 (N_976,In_125,In_732);
and U977 (N_977,In_481,In_1171);
or U978 (N_978,In_667,In_1359);
nor U979 (N_979,In_1882,In_754);
or U980 (N_980,In_1122,In_294);
or U981 (N_981,In_562,In_1326);
or U982 (N_982,In_1145,In_424);
or U983 (N_983,In_452,In_83);
nor U984 (N_984,In_937,In_406);
nand U985 (N_985,In_1184,In_395);
nand U986 (N_986,In_1558,In_317);
nand U987 (N_987,In_236,In_161);
nand U988 (N_988,In_872,In_749);
nor U989 (N_989,In_1068,In_535);
and U990 (N_990,In_556,In_380);
or U991 (N_991,In_1771,In_1149);
or U992 (N_992,In_513,In_1929);
nand U993 (N_993,In_1344,In_1770);
or U994 (N_994,In_1697,In_1954);
nand U995 (N_995,In_1432,In_677);
nand U996 (N_996,In_842,In_786);
and U997 (N_997,In_1766,In_34);
and U998 (N_998,In_1723,In_658);
nor U999 (N_999,In_1698,In_108);
or U1000 (N_1000,In_710,In_19);
nor U1001 (N_1001,In_577,In_460);
and U1002 (N_1002,In_1704,In_1915);
nor U1003 (N_1003,In_1859,In_1616);
nor U1004 (N_1004,In_273,In_1632);
or U1005 (N_1005,In_1924,In_228);
xnor U1006 (N_1006,In_172,In_1878);
xor U1007 (N_1007,In_486,In_1182);
nand U1008 (N_1008,In_1259,In_505);
or U1009 (N_1009,In_423,In_260);
and U1010 (N_1010,In_1801,In_304);
and U1011 (N_1011,In_638,In_1536);
and U1012 (N_1012,In_1238,In_214);
and U1013 (N_1013,In_1415,In_140);
xor U1014 (N_1014,In_46,In_320);
or U1015 (N_1015,In_1940,In_1193);
nand U1016 (N_1016,In_1611,In_928);
xnor U1017 (N_1017,In_220,In_1699);
xnor U1018 (N_1018,In_1477,In_1520);
and U1019 (N_1019,In_1644,In_1187);
nor U1020 (N_1020,In_1959,In_925);
xor U1021 (N_1021,In_1248,In_1804);
nor U1022 (N_1022,In_963,In_475);
or U1023 (N_1023,In_511,In_1479);
xnor U1024 (N_1024,In_1499,In_1804);
xnor U1025 (N_1025,In_1081,In_1611);
or U1026 (N_1026,In_640,In_1030);
nor U1027 (N_1027,In_1606,In_1127);
and U1028 (N_1028,In_351,In_1977);
or U1029 (N_1029,In_57,In_1388);
nand U1030 (N_1030,In_1861,In_1918);
xor U1031 (N_1031,In_1315,In_1281);
and U1032 (N_1032,In_1530,In_199);
nand U1033 (N_1033,In_55,In_356);
xor U1034 (N_1034,In_1126,In_565);
or U1035 (N_1035,In_1444,In_1831);
or U1036 (N_1036,In_207,In_315);
nor U1037 (N_1037,In_637,In_1423);
nor U1038 (N_1038,In_1144,In_294);
xor U1039 (N_1039,In_130,In_1700);
xor U1040 (N_1040,In_950,In_1557);
nor U1041 (N_1041,In_616,In_1986);
or U1042 (N_1042,In_710,In_1146);
nor U1043 (N_1043,In_961,In_597);
or U1044 (N_1044,In_1300,In_964);
and U1045 (N_1045,In_864,In_1959);
nor U1046 (N_1046,In_1997,In_296);
nand U1047 (N_1047,In_385,In_577);
nor U1048 (N_1048,In_1193,In_1551);
and U1049 (N_1049,In_112,In_1651);
xor U1050 (N_1050,In_839,In_710);
nand U1051 (N_1051,In_1883,In_877);
nand U1052 (N_1052,In_1900,In_1211);
and U1053 (N_1053,In_891,In_7);
and U1054 (N_1054,In_1979,In_590);
or U1055 (N_1055,In_597,In_165);
xnor U1056 (N_1056,In_753,In_135);
and U1057 (N_1057,In_1723,In_760);
and U1058 (N_1058,In_1449,In_568);
nand U1059 (N_1059,In_1533,In_1479);
nor U1060 (N_1060,In_385,In_446);
and U1061 (N_1061,In_1474,In_1212);
nand U1062 (N_1062,In_1543,In_109);
nand U1063 (N_1063,In_216,In_1933);
nor U1064 (N_1064,In_138,In_229);
nor U1065 (N_1065,In_395,In_1035);
or U1066 (N_1066,In_117,In_225);
or U1067 (N_1067,In_1921,In_59);
nand U1068 (N_1068,In_1267,In_396);
or U1069 (N_1069,In_1589,In_18);
nand U1070 (N_1070,In_1378,In_289);
xnor U1071 (N_1071,In_1218,In_1437);
and U1072 (N_1072,In_933,In_1079);
nor U1073 (N_1073,In_850,In_478);
nand U1074 (N_1074,In_1048,In_1632);
and U1075 (N_1075,In_1361,In_1255);
xnor U1076 (N_1076,In_1679,In_1563);
or U1077 (N_1077,In_460,In_887);
and U1078 (N_1078,In_239,In_962);
nor U1079 (N_1079,In_1043,In_1491);
or U1080 (N_1080,In_1361,In_1295);
nand U1081 (N_1081,In_739,In_1318);
or U1082 (N_1082,In_962,In_1321);
or U1083 (N_1083,In_1216,In_662);
or U1084 (N_1084,In_193,In_1036);
nand U1085 (N_1085,In_115,In_1884);
nand U1086 (N_1086,In_1038,In_1002);
and U1087 (N_1087,In_1259,In_1098);
nand U1088 (N_1088,In_1196,In_1794);
and U1089 (N_1089,In_118,In_272);
xor U1090 (N_1090,In_1060,In_463);
or U1091 (N_1091,In_936,In_1909);
xnor U1092 (N_1092,In_379,In_216);
nor U1093 (N_1093,In_1861,In_1433);
xnor U1094 (N_1094,In_1061,In_1042);
or U1095 (N_1095,In_117,In_1041);
and U1096 (N_1096,In_1967,In_916);
or U1097 (N_1097,In_1719,In_263);
nand U1098 (N_1098,In_7,In_1950);
or U1099 (N_1099,In_1714,In_1946);
and U1100 (N_1100,In_297,In_815);
xnor U1101 (N_1101,In_604,In_1873);
xor U1102 (N_1102,In_1424,In_1450);
and U1103 (N_1103,In_1068,In_1502);
xor U1104 (N_1104,In_1254,In_1551);
nor U1105 (N_1105,In_890,In_1285);
nor U1106 (N_1106,In_587,In_329);
nand U1107 (N_1107,In_796,In_13);
nor U1108 (N_1108,In_240,In_1267);
or U1109 (N_1109,In_633,In_1027);
or U1110 (N_1110,In_124,In_1426);
nor U1111 (N_1111,In_6,In_432);
and U1112 (N_1112,In_782,In_1559);
nor U1113 (N_1113,In_191,In_1059);
and U1114 (N_1114,In_845,In_835);
xnor U1115 (N_1115,In_1010,In_533);
nand U1116 (N_1116,In_1595,In_1088);
nor U1117 (N_1117,In_597,In_1207);
nand U1118 (N_1118,In_480,In_788);
nand U1119 (N_1119,In_8,In_1910);
nand U1120 (N_1120,In_499,In_170);
nor U1121 (N_1121,In_599,In_1729);
or U1122 (N_1122,In_309,In_1968);
nor U1123 (N_1123,In_392,In_1958);
and U1124 (N_1124,In_159,In_166);
nand U1125 (N_1125,In_1740,In_758);
and U1126 (N_1126,In_296,In_38);
nand U1127 (N_1127,In_512,In_1667);
and U1128 (N_1128,In_1427,In_1769);
nor U1129 (N_1129,In_1814,In_164);
nor U1130 (N_1130,In_1772,In_363);
xor U1131 (N_1131,In_72,In_1238);
xnor U1132 (N_1132,In_1611,In_543);
and U1133 (N_1133,In_394,In_639);
and U1134 (N_1134,In_811,In_329);
and U1135 (N_1135,In_740,In_839);
xor U1136 (N_1136,In_37,In_1156);
and U1137 (N_1137,In_804,In_1679);
or U1138 (N_1138,In_1080,In_1513);
nand U1139 (N_1139,In_277,In_1071);
and U1140 (N_1140,In_377,In_173);
nor U1141 (N_1141,In_450,In_1926);
and U1142 (N_1142,In_1797,In_1899);
xor U1143 (N_1143,In_1153,In_595);
or U1144 (N_1144,In_1827,In_1434);
nor U1145 (N_1145,In_1116,In_1521);
or U1146 (N_1146,In_804,In_1168);
xor U1147 (N_1147,In_323,In_102);
and U1148 (N_1148,In_1889,In_437);
xor U1149 (N_1149,In_1067,In_1830);
nand U1150 (N_1150,In_892,In_331);
or U1151 (N_1151,In_1422,In_1549);
nand U1152 (N_1152,In_702,In_1503);
and U1153 (N_1153,In_557,In_1694);
or U1154 (N_1154,In_570,In_639);
nor U1155 (N_1155,In_1793,In_305);
and U1156 (N_1156,In_1248,In_1207);
nand U1157 (N_1157,In_1475,In_1149);
or U1158 (N_1158,In_248,In_956);
or U1159 (N_1159,In_401,In_186);
nand U1160 (N_1160,In_775,In_829);
or U1161 (N_1161,In_1162,In_19);
or U1162 (N_1162,In_1334,In_412);
nor U1163 (N_1163,In_1186,In_1509);
nor U1164 (N_1164,In_204,In_282);
or U1165 (N_1165,In_537,In_1823);
xnor U1166 (N_1166,In_1280,In_595);
xor U1167 (N_1167,In_1300,In_993);
or U1168 (N_1168,In_231,In_1454);
and U1169 (N_1169,In_333,In_1566);
and U1170 (N_1170,In_1625,In_1829);
nor U1171 (N_1171,In_182,In_1878);
or U1172 (N_1172,In_9,In_1175);
or U1173 (N_1173,In_1096,In_1998);
and U1174 (N_1174,In_1019,In_648);
nand U1175 (N_1175,In_497,In_1270);
nor U1176 (N_1176,In_812,In_154);
xor U1177 (N_1177,In_769,In_1517);
nand U1178 (N_1178,In_735,In_598);
xor U1179 (N_1179,In_1975,In_590);
xor U1180 (N_1180,In_1168,In_1194);
xnor U1181 (N_1181,In_1554,In_884);
xnor U1182 (N_1182,In_1710,In_129);
or U1183 (N_1183,In_1131,In_1612);
nor U1184 (N_1184,In_1957,In_1033);
nand U1185 (N_1185,In_968,In_1429);
and U1186 (N_1186,In_1281,In_1964);
nand U1187 (N_1187,In_1755,In_424);
nand U1188 (N_1188,In_297,In_1826);
nor U1189 (N_1189,In_1735,In_91);
nand U1190 (N_1190,In_1320,In_396);
xnor U1191 (N_1191,In_1657,In_1945);
and U1192 (N_1192,In_21,In_245);
or U1193 (N_1193,In_1345,In_770);
nor U1194 (N_1194,In_243,In_1623);
xnor U1195 (N_1195,In_703,In_1765);
nor U1196 (N_1196,In_1274,In_759);
xnor U1197 (N_1197,In_1110,In_270);
nor U1198 (N_1198,In_1393,In_745);
and U1199 (N_1199,In_10,In_1352);
nor U1200 (N_1200,In_1121,In_1620);
and U1201 (N_1201,In_1727,In_663);
nor U1202 (N_1202,In_542,In_965);
and U1203 (N_1203,In_1771,In_531);
and U1204 (N_1204,In_893,In_124);
nor U1205 (N_1205,In_902,In_1054);
nor U1206 (N_1206,In_915,In_457);
or U1207 (N_1207,In_472,In_1794);
and U1208 (N_1208,In_1126,In_1401);
or U1209 (N_1209,In_1920,In_672);
and U1210 (N_1210,In_790,In_1286);
xnor U1211 (N_1211,In_371,In_1661);
nor U1212 (N_1212,In_95,In_1357);
xor U1213 (N_1213,In_1035,In_278);
and U1214 (N_1214,In_577,In_453);
and U1215 (N_1215,In_476,In_47);
nand U1216 (N_1216,In_750,In_920);
and U1217 (N_1217,In_578,In_1850);
or U1218 (N_1218,In_1036,In_1154);
or U1219 (N_1219,In_26,In_246);
xor U1220 (N_1220,In_1707,In_1981);
or U1221 (N_1221,In_1404,In_530);
nor U1222 (N_1222,In_1754,In_396);
nand U1223 (N_1223,In_1509,In_1723);
or U1224 (N_1224,In_1900,In_262);
and U1225 (N_1225,In_296,In_863);
and U1226 (N_1226,In_892,In_146);
nand U1227 (N_1227,In_781,In_1058);
nor U1228 (N_1228,In_1558,In_668);
nor U1229 (N_1229,In_806,In_370);
xnor U1230 (N_1230,In_535,In_1761);
nand U1231 (N_1231,In_1837,In_900);
nor U1232 (N_1232,In_1219,In_1133);
nor U1233 (N_1233,In_687,In_623);
nand U1234 (N_1234,In_963,In_613);
and U1235 (N_1235,In_253,In_538);
or U1236 (N_1236,In_909,In_373);
nor U1237 (N_1237,In_1327,In_1077);
nor U1238 (N_1238,In_190,In_454);
xnor U1239 (N_1239,In_1229,In_986);
nor U1240 (N_1240,In_646,In_1685);
nand U1241 (N_1241,In_291,In_583);
and U1242 (N_1242,In_55,In_227);
and U1243 (N_1243,In_1609,In_432);
nand U1244 (N_1244,In_294,In_1054);
and U1245 (N_1245,In_173,In_47);
and U1246 (N_1246,In_510,In_106);
or U1247 (N_1247,In_498,In_1872);
nor U1248 (N_1248,In_1524,In_914);
xor U1249 (N_1249,In_1562,In_21);
xor U1250 (N_1250,In_1543,In_375);
nand U1251 (N_1251,In_403,In_372);
xor U1252 (N_1252,In_1899,In_1723);
nor U1253 (N_1253,In_20,In_162);
or U1254 (N_1254,In_226,In_1025);
nand U1255 (N_1255,In_766,In_270);
or U1256 (N_1256,In_1538,In_782);
xnor U1257 (N_1257,In_210,In_1504);
nor U1258 (N_1258,In_1679,In_1835);
nand U1259 (N_1259,In_1729,In_514);
and U1260 (N_1260,In_167,In_560);
and U1261 (N_1261,In_1412,In_1824);
xor U1262 (N_1262,In_361,In_1922);
xor U1263 (N_1263,In_1132,In_276);
and U1264 (N_1264,In_1008,In_1598);
and U1265 (N_1265,In_788,In_1823);
and U1266 (N_1266,In_112,In_966);
and U1267 (N_1267,In_249,In_641);
nand U1268 (N_1268,In_1362,In_1929);
nor U1269 (N_1269,In_1035,In_1796);
xnor U1270 (N_1270,In_855,In_1514);
and U1271 (N_1271,In_947,In_1539);
nand U1272 (N_1272,In_1945,In_1707);
nor U1273 (N_1273,In_1801,In_737);
nand U1274 (N_1274,In_1853,In_118);
xor U1275 (N_1275,In_1842,In_880);
or U1276 (N_1276,In_899,In_415);
xnor U1277 (N_1277,In_1272,In_149);
and U1278 (N_1278,In_1189,In_1414);
and U1279 (N_1279,In_798,In_997);
and U1280 (N_1280,In_1442,In_76);
and U1281 (N_1281,In_379,In_1672);
xnor U1282 (N_1282,In_360,In_1534);
nor U1283 (N_1283,In_59,In_329);
and U1284 (N_1284,In_1475,In_707);
nor U1285 (N_1285,In_387,In_1112);
and U1286 (N_1286,In_1871,In_1675);
nor U1287 (N_1287,In_1348,In_1911);
or U1288 (N_1288,In_1733,In_568);
nand U1289 (N_1289,In_1355,In_995);
nor U1290 (N_1290,In_583,In_1682);
nand U1291 (N_1291,In_764,In_692);
xnor U1292 (N_1292,In_1432,In_285);
nand U1293 (N_1293,In_1482,In_562);
or U1294 (N_1294,In_1689,In_916);
or U1295 (N_1295,In_261,In_780);
or U1296 (N_1296,In_29,In_351);
and U1297 (N_1297,In_515,In_1386);
nor U1298 (N_1298,In_1665,In_1383);
nor U1299 (N_1299,In_612,In_1406);
xnor U1300 (N_1300,In_971,In_1203);
xnor U1301 (N_1301,In_474,In_1813);
and U1302 (N_1302,In_888,In_1073);
or U1303 (N_1303,In_1214,In_530);
nand U1304 (N_1304,In_605,In_73);
and U1305 (N_1305,In_981,In_1034);
or U1306 (N_1306,In_1784,In_408);
nor U1307 (N_1307,In_551,In_1792);
and U1308 (N_1308,In_813,In_930);
nand U1309 (N_1309,In_533,In_165);
nor U1310 (N_1310,In_833,In_448);
and U1311 (N_1311,In_370,In_1243);
or U1312 (N_1312,In_1028,In_1591);
and U1313 (N_1313,In_1682,In_127);
xor U1314 (N_1314,In_1259,In_737);
xor U1315 (N_1315,In_1755,In_1386);
xnor U1316 (N_1316,In_1715,In_35);
or U1317 (N_1317,In_1594,In_791);
nand U1318 (N_1318,In_1463,In_1749);
and U1319 (N_1319,In_63,In_235);
nor U1320 (N_1320,In_1311,In_231);
nand U1321 (N_1321,In_1885,In_1194);
nor U1322 (N_1322,In_173,In_1098);
nand U1323 (N_1323,In_111,In_1362);
nor U1324 (N_1324,In_1175,In_579);
nor U1325 (N_1325,In_1125,In_232);
or U1326 (N_1326,In_1612,In_1984);
nor U1327 (N_1327,In_199,In_1716);
and U1328 (N_1328,In_1017,In_812);
or U1329 (N_1329,In_1128,In_390);
nor U1330 (N_1330,In_1550,In_860);
nor U1331 (N_1331,In_1416,In_1917);
xor U1332 (N_1332,In_1525,In_1478);
nor U1333 (N_1333,In_1288,In_1319);
nor U1334 (N_1334,In_495,In_223);
and U1335 (N_1335,In_1638,In_1575);
xnor U1336 (N_1336,In_1302,In_599);
nor U1337 (N_1337,In_832,In_752);
nor U1338 (N_1338,In_1189,In_1681);
or U1339 (N_1339,In_841,In_1341);
and U1340 (N_1340,In_1682,In_1912);
nor U1341 (N_1341,In_44,In_1792);
xor U1342 (N_1342,In_786,In_1758);
nand U1343 (N_1343,In_788,In_1841);
nor U1344 (N_1344,In_674,In_562);
or U1345 (N_1345,In_41,In_1847);
xnor U1346 (N_1346,In_1381,In_426);
nand U1347 (N_1347,In_1427,In_1794);
nor U1348 (N_1348,In_1423,In_1513);
nor U1349 (N_1349,In_1369,In_473);
nor U1350 (N_1350,In_531,In_1592);
nor U1351 (N_1351,In_1367,In_401);
or U1352 (N_1352,In_353,In_1906);
nor U1353 (N_1353,In_1032,In_1893);
nand U1354 (N_1354,In_1045,In_442);
nor U1355 (N_1355,In_83,In_153);
xor U1356 (N_1356,In_1386,In_1319);
nor U1357 (N_1357,In_1120,In_482);
nor U1358 (N_1358,In_33,In_747);
nand U1359 (N_1359,In_546,In_1258);
nor U1360 (N_1360,In_1292,In_1673);
or U1361 (N_1361,In_734,In_1118);
nor U1362 (N_1362,In_594,In_707);
nand U1363 (N_1363,In_108,In_1036);
nand U1364 (N_1364,In_819,In_1058);
nand U1365 (N_1365,In_138,In_1850);
and U1366 (N_1366,In_1819,In_208);
xor U1367 (N_1367,In_90,In_852);
or U1368 (N_1368,In_746,In_243);
or U1369 (N_1369,In_1174,In_67);
and U1370 (N_1370,In_941,In_457);
or U1371 (N_1371,In_1662,In_852);
and U1372 (N_1372,In_1540,In_817);
and U1373 (N_1373,In_561,In_754);
xor U1374 (N_1374,In_1861,In_1664);
or U1375 (N_1375,In_1114,In_221);
nand U1376 (N_1376,In_1133,In_1788);
nand U1377 (N_1377,In_433,In_1851);
nand U1378 (N_1378,In_179,In_698);
nand U1379 (N_1379,In_782,In_1352);
or U1380 (N_1380,In_473,In_1109);
and U1381 (N_1381,In_1271,In_722);
nand U1382 (N_1382,In_456,In_301);
nor U1383 (N_1383,In_1881,In_1445);
or U1384 (N_1384,In_368,In_10);
nor U1385 (N_1385,In_1598,In_1004);
or U1386 (N_1386,In_905,In_423);
or U1387 (N_1387,In_665,In_1713);
nor U1388 (N_1388,In_856,In_175);
xor U1389 (N_1389,In_1621,In_943);
xor U1390 (N_1390,In_575,In_1560);
nor U1391 (N_1391,In_1460,In_1492);
nand U1392 (N_1392,In_43,In_985);
and U1393 (N_1393,In_1012,In_1363);
nor U1394 (N_1394,In_237,In_1477);
nand U1395 (N_1395,In_416,In_1051);
nand U1396 (N_1396,In_297,In_1307);
nand U1397 (N_1397,In_1192,In_223);
xor U1398 (N_1398,In_8,In_1400);
nand U1399 (N_1399,In_591,In_623);
nor U1400 (N_1400,In_695,In_999);
or U1401 (N_1401,In_1568,In_451);
and U1402 (N_1402,In_1878,In_540);
nand U1403 (N_1403,In_1376,In_1808);
xor U1404 (N_1404,In_1906,In_1432);
nand U1405 (N_1405,In_1799,In_664);
and U1406 (N_1406,In_1436,In_1519);
nand U1407 (N_1407,In_493,In_402);
nor U1408 (N_1408,In_2,In_550);
nand U1409 (N_1409,In_1024,In_88);
and U1410 (N_1410,In_575,In_698);
xnor U1411 (N_1411,In_1743,In_1521);
or U1412 (N_1412,In_275,In_1784);
and U1413 (N_1413,In_1933,In_1632);
or U1414 (N_1414,In_219,In_491);
nand U1415 (N_1415,In_51,In_331);
or U1416 (N_1416,In_438,In_1824);
or U1417 (N_1417,In_684,In_410);
or U1418 (N_1418,In_154,In_196);
xor U1419 (N_1419,In_1364,In_1193);
nand U1420 (N_1420,In_76,In_1928);
or U1421 (N_1421,In_1319,In_1061);
or U1422 (N_1422,In_1579,In_1887);
and U1423 (N_1423,In_1520,In_138);
nor U1424 (N_1424,In_1800,In_312);
nand U1425 (N_1425,In_1320,In_60);
or U1426 (N_1426,In_1244,In_43);
and U1427 (N_1427,In_1728,In_220);
and U1428 (N_1428,In_937,In_483);
and U1429 (N_1429,In_610,In_1501);
or U1430 (N_1430,In_1439,In_1212);
and U1431 (N_1431,In_60,In_1348);
xnor U1432 (N_1432,In_1021,In_897);
nor U1433 (N_1433,In_1048,In_1169);
nand U1434 (N_1434,In_308,In_1350);
or U1435 (N_1435,In_50,In_1308);
or U1436 (N_1436,In_1668,In_551);
or U1437 (N_1437,In_383,In_8);
or U1438 (N_1438,In_1029,In_215);
and U1439 (N_1439,In_1547,In_850);
and U1440 (N_1440,In_938,In_413);
or U1441 (N_1441,In_357,In_1480);
nand U1442 (N_1442,In_1366,In_124);
or U1443 (N_1443,In_316,In_47);
xnor U1444 (N_1444,In_1357,In_986);
and U1445 (N_1445,In_942,In_1658);
nor U1446 (N_1446,In_683,In_908);
and U1447 (N_1447,In_495,In_1113);
xnor U1448 (N_1448,In_667,In_1675);
or U1449 (N_1449,In_1906,In_605);
and U1450 (N_1450,In_1283,In_1744);
xnor U1451 (N_1451,In_256,In_180);
nor U1452 (N_1452,In_1882,In_1297);
xor U1453 (N_1453,In_221,In_919);
nor U1454 (N_1454,In_1664,In_1187);
xor U1455 (N_1455,In_12,In_206);
and U1456 (N_1456,In_1108,In_103);
and U1457 (N_1457,In_1389,In_55);
xor U1458 (N_1458,In_6,In_660);
xnor U1459 (N_1459,In_1593,In_1541);
and U1460 (N_1460,In_749,In_1300);
nand U1461 (N_1461,In_1949,In_362);
nand U1462 (N_1462,In_1242,In_542);
nor U1463 (N_1463,In_104,In_68);
nand U1464 (N_1464,In_80,In_374);
or U1465 (N_1465,In_298,In_127);
xnor U1466 (N_1466,In_833,In_237);
nand U1467 (N_1467,In_1766,In_715);
xnor U1468 (N_1468,In_1011,In_1434);
nand U1469 (N_1469,In_970,In_1155);
or U1470 (N_1470,In_1084,In_1425);
xor U1471 (N_1471,In_436,In_811);
xnor U1472 (N_1472,In_665,In_1323);
nand U1473 (N_1473,In_1008,In_1217);
nand U1474 (N_1474,In_1735,In_730);
and U1475 (N_1475,In_1081,In_1958);
nor U1476 (N_1476,In_412,In_799);
nand U1477 (N_1477,In_730,In_425);
and U1478 (N_1478,In_1491,In_1442);
nand U1479 (N_1479,In_1590,In_264);
nor U1480 (N_1480,In_1619,In_1365);
nor U1481 (N_1481,In_327,In_936);
nand U1482 (N_1482,In_938,In_917);
and U1483 (N_1483,In_1230,In_1204);
xnor U1484 (N_1484,In_865,In_1244);
nand U1485 (N_1485,In_1770,In_1048);
and U1486 (N_1486,In_68,In_1855);
nor U1487 (N_1487,In_1750,In_1496);
nand U1488 (N_1488,In_651,In_1858);
or U1489 (N_1489,In_1885,In_1233);
nor U1490 (N_1490,In_923,In_1060);
xnor U1491 (N_1491,In_204,In_842);
and U1492 (N_1492,In_1243,In_1900);
and U1493 (N_1493,In_1355,In_1898);
or U1494 (N_1494,In_668,In_569);
or U1495 (N_1495,In_126,In_158);
nand U1496 (N_1496,In_3,In_1368);
and U1497 (N_1497,In_542,In_125);
or U1498 (N_1498,In_450,In_508);
or U1499 (N_1499,In_1238,In_1419);
nor U1500 (N_1500,In_591,In_868);
and U1501 (N_1501,In_751,In_676);
nand U1502 (N_1502,In_421,In_1983);
xnor U1503 (N_1503,In_954,In_1737);
nor U1504 (N_1504,In_18,In_49);
nand U1505 (N_1505,In_371,In_1266);
nand U1506 (N_1506,In_1513,In_1862);
nor U1507 (N_1507,In_536,In_976);
nor U1508 (N_1508,In_1203,In_1108);
nor U1509 (N_1509,In_1842,In_1806);
nand U1510 (N_1510,In_82,In_1763);
or U1511 (N_1511,In_832,In_261);
and U1512 (N_1512,In_1600,In_484);
or U1513 (N_1513,In_503,In_1953);
xnor U1514 (N_1514,In_987,In_112);
and U1515 (N_1515,In_829,In_770);
nor U1516 (N_1516,In_150,In_230);
nor U1517 (N_1517,In_639,In_217);
nor U1518 (N_1518,In_100,In_721);
and U1519 (N_1519,In_1205,In_1591);
nand U1520 (N_1520,In_1937,In_177);
xor U1521 (N_1521,In_682,In_1208);
or U1522 (N_1522,In_1464,In_519);
xnor U1523 (N_1523,In_1760,In_375);
xnor U1524 (N_1524,In_1670,In_1819);
and U1525 (N_1525,In_800,In_166);
xor U1526 (N_1526,In_849,In_1761);
nor U1527 (N_1527,In_68,In_1161);
nor U1528 (N_1528,In_607,In_702);
and U1529 (N_1529,In_1133,In_1976);
nor U1530 (N_1530,In_1639,In_162);
nand U1531 (N_1531,In_1993,In_496);
nor U1532 (N_1532,In_706,In_1287);
xnor U1533 (N_1533,In_1279,In_849);
or U1534 (N_1534,In_152,In_1900);
or U1535 (N_1535,In_629,In_1341);
nand U1536 (N_1536,In_1092,In_152);
nor U1537 (N_1537,In_608,In_563);
nor U1538 (N_1538,In_901,In_128);
nor U1539 (N_1539,In_401,In_1609);
nor U1540 (N_1540,In_1416,In_0);
or U1541 (N_1541,In_1757,In_255);
nor U1542 (N_1542,In_1060,In_530);
or U1543 (N_1543,In_1676,In_825);
or U1544 (N_1544,In_1665,In_1067);
nor U1545 (N_1545,In_318,In_534);
nand U1546 (N_1546,In_1641,In_168);
xnor U1547 (N_1547,In_1845,In_1897);
and U1548 (N_1548,In_1094,In_292);
nor U1549 (N_1549,In_659,In_1429);
nor U1550 (N_1550,In_611,In_999);
xnor U1551 (N_1551,In_793,In_93);
or U1552 (N_1552,In_962,In_1107);
or U1553 (N_1553,In_916,In_240);
nor U1554 (N_1554,In_1764,In_669);
and U1555 (N_1555,In_1838,In_156);
and U1556 (N_1556,In_1836,In_1469);
or U1557 (N_1557,In_1125,In_1359);
and U1558 (N_1558,In_778,In_470);
nand U1559 (N_1559,In_366,In_1670);
nor U1560 (N_1560,In_1163,In_796);
xor U1561 (N_1561,In_1021,In_8);
xnor U1562 (N_1562,In_1518,In_144);
or U1563 (N_1563,In_1360,In_11);
nor U1564 (N_1564,In_263,In_1506);
nor U1565 (N_1565,In_1372,In_1008);
nand U1566 (N_1566,In_363,In_1667);
nor U1567 (N_1567,In_1337,In_1949);
or U1568 (N_1568,In_1328,In_19);
and U1569 (N_1569,In_1793,In_1812);
xnor U1570 (N_1570,In_1703,In_1079);
and U1571 (N_1571,In_1474,In_1688);
and U1572 (N_1572,In_835,In_1684);
and U1573 (N_1573,In_221,In_652);
xnor U1574 (N_1574,In_444,In_1698);
and U1575 (N_1575,In_1817,In_40);
and U1576 (N_1576,In_743,In_317);
xor U1577 (N_1577,In_7,In_1250);
nand U1578 (N_1578,In_1228,In_1652);
nor U1579 (N_1579,In_267,In_762);
nand U1580 (N_1580,In_3,In_1124);
nand U1581 (N_1581,In_1040,In_485);
nor U1582 (N_1582,In_492,In_585);
and U1583 (N_1583,In_1572,In_403);
or U1584 (N_1584,In_1424,In_1587);
nand U1585 (N_1585,In_1350,In_427);
or U1586 (N_1586,In_77,In_685);
and U1587 (N_1587,In_1974,In_290);
xor U1588 (N_1588,In_592,In_1293);
and U1589 (N_1589,In_1367,In_1988);
and U1590 (N_1590,In_1010,In_201);
xnor U1591 (N_1591,In_257,In_1925);
xnor U1592 (N_1592,In_823,In_520);
and U1593 (N_1593,In_1508,In_832);
xor U1594 (N_1594,In_1393,In_1715);
nor U1595 (N_1595,In_368,In_639);
nor U1596 (N_1596,In_550,In_1408);
xor U1597 (N_1597,In_1263,In_497);
nor U1598 (N_1598,In_325,In_1453);
or U1599 (N_1599,In_12,In_513);
nand U1600 (N_1600,In_197,In_638);
and U1601 (N_1601,In_95,In_1901);
and U1602 (N_1602,In_157,In_1399);
or U1603 (N_1603,In_1063,In_742);
nor U1604 (N_1604,In_1116,In_300);
nor U1605 (N_1605,In_1526,In_185);
nor U1606 (N_1606,In_1296,In_1376);
xor U1607 (N_1607,In_197,In_107);
or U1608 (N_1608,In_1437,In_1161);
xor U1609 (N_1609,In_380,In_1339);
nand U1610 (N_1610,In_683,In_1655);
nor U1611 (N_1611,In_1166,In_1577);
nand U1612 (N_1612,In_1347,In_1081);
and U1613 (N_1613,In_1687,In_1053);
and U1614 (N_1614,In_1478,In_1402);
nand U1615 (N_1615,In_1109,In_583);
nand U1616 (N_1616,In_1703,In_732);
nor U1617 (N_1617,In_1090,In_1645);
or U1618 (N_1618,In_712,In_1639);
or U1619 (N_1619,In_741,In_563);
xnor U1620 (N_1620,In_648,In_1553);
xnor U1621 (N_1621,In_1855,In_1768);
xnor U1622 (N_1622,In_4,In_1287);
nand U1623 (N_1623,In_1024,In_1390);
xor U1624 (N_1624,In_677,In_1876);
nor U1625 (N_1625,In_474,In_1793);
and U1626 (N_1626,In_1176,In_832);
nor U1627 (N_1627,In_1509,In_186);
and U1628 (N_1628,In_1950,In_243);
nor U1629 (N_1629,In_586,In_1351);
and U1630 (N_1630,In_1251,In_958);
xor U1631 (N_1631,In_1456,In_1717);
nor U1632 (N_1632,In_848,In_631);
or U1633 (N_1633,In_1678,In_1197);
xor U1634 (N_1634,In_1450,In_891);
nor U1635 (N_1635,In_991,In_1937);
xor U1636 (N_1636,In_1411,In_1605);
or U1637 (N_1637,In_1204,In_107);
nor U1638 (N_1638,In_1673,In_1761);
and U1639 (N_1639,In_570,In_129);
and U1640 (N_1640,In_1517,In_1740);
or U1641 (N_1641,In_1458,In_769);
xnor U1642 (N_1642,In_461,In_901);
or U1643 (N_1643,In_1557,In_794);
and U1644 (N_1644,In_1136,In_717);
nor U1645 (N_1645,In_133,In_0);
nand U1646 (N_1646,In_1777,In_477);
or U1647 (N_1647,In_1817,In_1963);
and U1648 (N_1648,In_1088,In_1731);
and U1649 (N_1649,In_982,In_1254);
or U1650 (N_1650,In_1064,In_132);
and U1651 (N_1651,In_1137,In_1947);
and U1652 (N_1652,In_1461,In_313);
and U1653 (N_1653,In_1637,In_404);
nor U1654 (N_1654,In_1319,In_228);
or U1655 (N_1655,In_739,In_1612);
and U1656 (N_1656,In_255,In_389);
and U1657 (N_1657,In_881,In_985);
or U1658 (N_1658,In_664,In_1424);
xnor U1659 (N_1659,In_1798,In_1934);
nand U1660 (N_1660,In_941,In_1008);
nor U1661 (N_1661,In_1821,In_1339);
or U1662 (N_1662,In_1725,In_689);
xnor U1663 (N_1663,In_1289,In_149);
xor U1664 (N_1664,In_1190,In_509);
or U1665 (N_1665,In_1440,In_1830);
and U1666 (N_1666,In_462,In_1868);
nor U1667 (N_1667,In_821,In_376);
nor U1668 (N_1668,In_10,In_1558);
and U1669 (N_1669,In_251,In_856);
and U1670 (N_1670,In_1519,In_823);
nor U1671 (N_1671,In_64,In_1084);
and U1672 (N_1672,In_1240,In_689);
nand U1673 (N_1673,In_145,In_1578);
and U1674 (N_1674,In_393,In_182);
nand U1675 (N_1675,In_525,In_1905);
or U1676 (N_1676,In_1362,In_1783);
nor U1677 (N_1677,In_476,In_499);
nand U1678 (N_1678,In_710,In_1938);
xor U1679 (N_1679,In_1439,In_1197);
nand U1680 (N_1680,In_970,In_1548);
xor U1681 (N_1681,In_710,In_1278);
nand U1682 (N_1682,In_654,In_887);
xnor U1683 (N_1683,In_130,In_295);
and U1684 (N_1684,In_176,In_245);
xnor U1685 (N_1685,In_765,In_407);
nor U1686 (N_1686,In_1109,In_1082);
or U1687 (N_1687,In_1059,In_1732);
xnor U1688 (N_1688,In_1985,In_210);
or U1689 (N_1689,In_1310,In_542);
and U1690 (N_1690,In_1211,In_685);
or U1691 (N_1691,In_1732,In_708);
xnor U1692 (N_1692,In_83,In_1885);
or U1693 (N_1693,In_839,In_1888);
and U1694 (N_1694,In_1928,In_997);
and U1695 (N_1695,In_1865,In_245);
nor U1696 (N_1696,In_1956,In_403);
and U1697 (N_1697,In_1288,In_1453);
nand U1698 (N_1698,In_330,In_1373);
and U1699 (N_1699,In_1451,In_199);
or U1700 (N_1700,In_1553,In_79);
xnor U1701 (N_1701,In_706,In_908);
or U1702 (N_1702,In_1745,In_1155);
and U1703 (N_1703,In_50,In_503);
nor U1704 (N_1704,In_478,In_1727);
xnor U1705 (N_1705,In_1816,In_597);
xnor U1706 (N_1706,In_591,In_43);
and U1707 (N_1707,In_1194,In_715);
nor U1708 (N_1708,In_691,In_1852);
xnor U1709 (N_1709,In_1536,In_331);
and U1710 (N_1710,In_1797,In_1842);
nor U1711 (N_1711,In_489,In_1731);
nand U1712 (N_1712,In_783,In_910);
xor U1713 (N_1713,In_759,In_1298);
or U1714 (N_1714,In_363,In_1206);
xor U1715 (N_1715,In_276,In_939);
xor U1716 (N_1716,In_26,In_1408);
xor U1717 (N_1717,In_220,In_1211);
nor U1718 (N_1718,In_531,In_1380);
xnor U1719 (N_1719,In_1850,In_1241);
xnor U1720 (N_1720,In_1382,In_1383);
xor U1721 (N_1721,In_722,In_217);
or U1722 (N_1722,In_1184,In_1685);
nand U1723 (N_1723,In_742,In_1409);
nand U1724 (N_1724,In_1001,In_992);
nor U1725 (N_1725,In_1881,In_950);
and U1726 (N_1726,In_728,In_634);
or U1727 (N_1727,In_1120,In_1978);
nand U1728 (N_1728,In_1119,In_199);
or U1729 (N_1729,In_514,In_29);
nand U1730 (N_1730,In_863,In_336);
xor U1731 (N_1731,In_290,In_941);
xnor U1732 (N_1732,In_1015,In_1445);
and U1733 (N_1733,In_1616,In_663);
xor U1734 (N_1734,In_1568,In_1088);
nor U1735 (N_1735,In_178,In_1755);
and U1736 (N_1736,In_326,In_48);
or U1737 (N_1737,In_898,In_603);
nor U1738 (N_1738,In_1598,In_148);
nand U1739 (N_1739,In_958,In_486);
xor U1740 (N_1740,In_1465,In_600);
and U1741 (N_1741,In_1424,In_1082);
nor U1742 (N_1742,In_1299,In_970);
nor U1743 (N_1743,In_1319,In_618);
xnor U1744 (N_1744,In_240,In_1786);
xnor U1745 (N_1745,In_1167,In_1181);
nand U1746 (N_1746,In_432,In_41);
xor U1747 (N_1747,In_194,In_763);
xor U1748 (N_1748,In_1189,In_666);
and U1749 (N_1749,In_1434,In_1297);
nand U1750 (N_1750,In_312,In_1533);
nand U1751 (N_1751,In_1377,In_1140);
and U1752 (N_1752,In_1044,In_1087);
xnor U1753 (N_1753,In_318,In_1768);
nand U1754 (N_1754,In_1445,In_870);
nor U1755 (N_1755,In_1430,In_259);
nor U1756 (N_1756,In_1558,In_1588);
and U1757 (N_1757,In_1442,In_652);
nand U1758 (N_1758,In_746,In_1146);
xor U1759 (N_1759,In_713,In_799);
or U1760 (N_1760,In_1241,In_1150);
nor U1761 (N_1761,In_1534,In_1255);
xor U1762 (N_1762,In_1925,In_1076);
and U1763 (N_1763,In_538,In_912);
nor U1764 (N_1764,In_1247,In_876);
nand U1765 (N_1765,In_746,In_979);
and U1766 (N_1766,In_1958,In_729);
nand U1767 (N_1767,In_1308,In_708);
xnor U1768 (N_1768,In_905,In_138);
nand U1769 (N_1769,In_82,In_1846);
or U1770 (N_1770,In_621,In_1332);
or U1771 (N_1771,In_1254,In_566);
nor U1772 (N_1772,In_872,In_625);
and U1773 (N_1773,In_62,In_422);
nand U1774 (N_1774,In_342,In_511);
nor U1775 (N_1775,In_1630,In_806);
nor U1776 (N_1776,In_877,In_834);
or U1777 (N_1777,In_1543,In_920);
xnor U1778 (N_1778,In_1581,In_1911);
nor U1779 (N_1779,In_349,In_1118);
nor U1780 (N_1780,In_719,In_687);
nor U1781 (N_1781,In_1724,In_759);
nor U1782 (N_1782,In_846,In_249);
nor U1783 (N_1783,In_1336,In_763);
nor U1784 (N_1784,In_1626,In_652);
and U1785 (N_1785,In_1826,In_1032);
or U1786 (N_1786,In_134,In_811);
nand U1787 (N_1787,In_399,In_1578);
or U1788 (N_1788,In_244,In_1058);
nand U1789 (N_1789,In_188,In_1039);
nand U1790 (N_1790,In_1472,In_1406);
nor U1791 (N_1791,In_311,In_811);
nor U1792 (N_1792,In_1358,In_340);
or U1793 (N_1793,In_548,In_1412);
nand U1794 (N_1794,In_1839,In_1883);
or U1795 (N_1795,In_1401,In_519);
xnor U1796 (N_1796,In_1893,In_1546);
and U1797 (N_1797,In_1277,In_1939);
and U1798 (N_1798,In_1119,In_1810);
xor U1799 (N_1799,In_518,In_1569);
nor U1800 (N_1800,In_530,In_200);
nand U1801 (N_1801,In_1251,In_1897);
or U1802 (N_1802,In_1139,In_298);
or U1803 (N_1803,In_1445,In_606);
or U1804 (N_1804,In_1884,In_378);
nand U1805 (N_1805,In_1535,In_1242);
nand U1806 (N_1806,In_1573,In_252);
nand U1807 (N_1807,In_675,In_1455);
nor U1808 (N_1808,In_64,In_552);
nor U1809 (N_1809,In_1980,In_333);
nand U1810 (N_1810,In_1755,In_1934);
xor U1811 (N_1811,In_749,In_1211);
nand U1812 (N_1812,In_1626,In_1987);
and U1813 (N_1813,In_715,In_307);
nor U1814 (N_1814,In_1477,In_1957);
xor U1815 (N_1815,In_1618,In_1497);
and U1816 (N_1816,In_1181,In_1727);
nor U1817 (N_1817,In_1246,In_356);
xor U1818 (N_1818,In_1383,In_181);
or U1819 (N_1819,In_1373,In_1662);
xnor U1820 (N_1820,In_343,In_1005);
nor U1821 (N_1821,In_1219,In_868);
and U1822 (N_1822,In_244,In_1509);
or U1823 (N_1823,In_1287,In_149);
nor U1824 (N_1824,In_597,In_1440);
xnor U1825 (N_1825,In_1484,In_1038);
and U1826 (N_1826,In_556,In_837);
xor U1827 (N_1827,In_1548,In_1518);
or U1828 (N_1828,In_225,In_1010);
nand U1829 (N_1829,In_991,In_833);
nor U1830 (N_1830,In_894,In_1937);
xor U1831 (N_1831,In_972,In_1152);
nand U1832 (N_1832,In_1743,In_1208);
or U1833 (N_1833,In_1456,In_656);
and U1834 (N_1834,In_216,In_1210);
and U1835 (N_1835,In_1746,In_451);
or U1836 (N_1836,In_1890,In_20);
xor U1837 (N_1837,In_851,In_1626);
xor U1838 (N_1838,In_1533,In_291);
nand U1839 (N_1839,In_747,In_1795);
or U1840 (N_1840,In_831,In_871);
nor U1841 (N_1841,In_635,In_1648);
xor U1842 (N_1842,In_1746,In_148);
or U1843 (N_1843,In_26,In_438);
xnor U1844 (N_1844,In_1727,In_215);
or U1845 (N_1845,In_1214,In_1228);
nor U1846 (N_1846,In_601,In_762);
and U1847 (N_1847,In_1959,In_1904);
or U1848 (N_1848,In_1605,In_1744);
nand U1849 (N_1849,In_1805,In_608);
and U1850 (N_1850,In_474,In_399);
xor U1851 (N_1851,In_1124,In_157);
or U1852 (N_1852,In_1904,In_1523);
xnor U1853 (N_1853,In_1164,In_1763);
nand U1854 (N_1854,In_1736,In_383);
or U1855 (N_1855,In_1809,In_1820);
and U1856 (N_1856,In_1025,In_1823);
xor U1857 (N_1857,In_1099,In_1420);
nor U1858 (N_1858,In_160,In_1182);
xor U1859 (N_1859,In_589,In_1238);
or U1860 (N_1860,In_1883,In_1921);
nor U1861 (N_1861,In_1894,In_1186);
nor U1862 (N_1862,In_1819,In_1822);
nand U1863 (N_1863,In_517,In_467);
xnor U1864 (N_1864,In_78,In_1493);
nor U1865 (N_1865,In_743,In_590);
xnor U1866 (N_1866,In_1507,In_1264);
xor U1867 (N_1867,In_183,In_1334);
nand U1868 (N_1868,In_199,In_764);
or U1869 (N_1869,In_1342,In_1766);
nor U1870 (N_1870,In_1327,In_76);
xor U1871 (N_1871,In_388,In_416);
xnor U1872 (N_1872,In_562,In_812);
nand U1873 (N_1873,In_898,In_612);
nand U1874 (N_1874,In_975,In_1945);
nor U1875 (N_1875,In_977,In_1027);
and U1876 (N_1876,In_1553,In_1731);
nand U1877 (N_1877,In_555,In_608);
nor U1878 (N_1878,In_1225,In_397);
nor U1879 (N_1879,In_902,In_1247);
and U1880 (N_1880,In_1147,In_1875);
or U1881 (N_1881,In_1269,In_562);
or U1882 (N_1882,In_1636,In_1304);
or U1883 (N_1883,In_285,In_480);
nand U1884 (N_1884,In_958,In_393);
nor U1885 (N_1885,In_1735,In_1486);
and U1886 (N_1886,In_623,In_1295);
or U1887 (N_1887,In_618,In_1251);
nor U1888 (N_1888,In_547,In_25);
and U1889 (N_1889,In_1469,In_819);
nand U1890 (N_1890,In_804,In_419);
xnor U1891 (N_1891,In_964,In_1914);
nand U1892 (N_1892,In_251,In_1280);
and U1893 (N_1893,In_718,In_282);
nand U1894 (N_1894,In_300,In_380);
nand U1895 (N_1895,In_539,In_786);
nor U1896 (N_1896,In_877,In_237);
nor U1897 (N_1897,In_1533,In_1924);
and U1898 (N_1898,In_1027,In_480);
xnor U1899 (N_1899,In_1581,In_252);
nor U1900 (N_1900,In_147,In_1568);
and U1901 (N_1901,In_369,In_1407);
xnor U1902 (N_1902,In_830,In_686);
and U1903 (N_1903,In_744,In_302);
or U1904 (N_1904,In_256,In_1446);
or U1905 (N_1905,In_1263,In_153);
or U1906 (N_1906,In_1296,In_938);
xnor U1907 (N_1907,In_638,In_888);
or U1908 (N_1908,In_301,In_670);
or U1909 (N_1909,In_89,In_1604);
nor U1910 (N_1910,In_609,In_758);
nand U1911 (N_1911,In_1733,In_536);
and U1912 (N_1912,In_473,In_1174);
nor U1913 (N_1913,In_822,In_1559);
xnor U1914 (N_1914,In_1605,In_36);
nor U1915 (N_1915,In_368,In_1714);
or U1916 (N_1916,In_1929,In_1881);
and U1917 (N_1917,In_366,In_1745);
nand U1918 (N_1918,In_1301,In_742);
nand U1919 (N_1919,In_1788,In_241);
or U1920 (N_1920,In_1102,In_1158);
nand U1921 (N_1921,In_1927,In_1194);
or U1922 (N_1922,In_997,In_1794);
or U1923 (N_1923,In_1139,In_294);
or U1924 (N_1924,In_447,In_882);
and U1925 (N_1925,In_1792,In_244);
or U1926 (N_1926,In_505,In_1880);
nand U1927 (N_1927,In_1770,In_1169);
nand U1928 (N_1928,In_1641,In_1985);
or U1929 (N_1929,In_1030,In_411);
nor U1930 (N_1930,In_1828,In_698);
xnor U1931 (N_1931,In_1255,In_604);
nor U1932 (N_1932,In_161,In_1551);
nand U1933 (N_1933,In_1739,In_1038);
and U1934 (N_1934,In_1584,In_854);
and U1935 (N_1935,In_1843,In_408);
nor U1936 (N_1936,In_982,In_1420);
xnor U1937 (N_1937,In_242,In_1769);
or U1938 (N_1938,In_123,In_647);
nor U1939 (N_1939,In_1813,In_827);
or U1940 (N_1940,In_33,In_1017);
or U1941 (N_1941,In_1349,In_1795);
or U1942 (N_1942,In_523,In_1645);
nor U1943 (N_1943,In_928,In_1914);
nor U1944 (N_1944,In_1712,In_372);
xnor U1945 (N_1945,In_6,In_847);
xor U1946 (N_1946,In_770,In_624);
nor U1947 (N_1947,In_1876,In_1043);
nor U1948 (N_1948,In_20,In_895);
nand U1949 (N_1949,In_1262,In_1259);
nor U1950 (N_1950,In_529,In_560);
nor U1951 (N_1951,In_1488,In_1822);
or U1952 (N_1952,In_1525,In_1755);
nand U1953 (N_1953,In_727,In_1697);
xor U1954 (N_1954,In_1871,In_1039);
or U1955 (N_1955,In_942,In_221);
and U1956 (N_1956,In_594,In_174);
or U1957 (N_1957,In_409,In_1237);
or U1958 (N_1958,In_1149,In_1251);
and U1959 (N_1959,In_1068,In_1086);
xor U1960 (N_1960,In_1845,In_1115);
nand U1961 (N_1961,In_969,In_1681);
nand U1962 (N_1962,In_615,In_1428);
and U1963 (N_1963,In_357,In_735);
nand U1964 (N_1964,In_1093,In_181);
xnor U1965 (N_1965,In_1091,In_1852);
and U1966 (N_1966,In_710,In_199);
nor U1967 (N_1967,In_1009,In_1290);
or U1968 (N_1968,In_1655,In_1856);
or U1969 (N_1969,In_944,In_1910);
nand U1970 (N_1970,In_1969,In_1323);
nor U1971 (N_1971,In_1129,In_1866);
nand U1972 (N_1972,In_870,In_1625);
or U1973 (N_1973,In_1624,In_784);
xor U1974 (N_1974,In_1553,In_1230);
nand U1975 (N_1975,In_1699,In_700);
or U1976 (N_1976,In_695,In_259);
nor U1977 (N_1977,In_670,In_574);
nand U1978 (N_1978,In_1818,In_1731);
xor U1979 (N_1979,In_1832,In_1275);
xnor U1980 (N_1980,In_1758,In_1732);
or U1981 (N_1981,In_799,In_484);
or U1982 (N_1982,In_75,In_1912);
and U1983 (N_1983,In_1166,In_621);
nand U1984 (N_1984,In_1001,In_1200);
nand U1985 (N_1985,In_940,In_1166);
xor U1986 (N_1986,In_1511,In_842);
nor U1987 (N_1987,In_1995,In_446);
or U1988 (N_1988,In_1602,In_1925);
xnor U1989 (N_1989,In_1223,In_266);
nand U1990 (N_1990,In_289,In_987);
nor U1991 (N_1991,In_858,In_250);
nor U1992 (N_1992,In_263,In_1150);
and U1993 (N_1993,In_1959,In_1694);
nand U1994 (N_1994,In_488,In_1082);
nand U1995 (N_1995,In_431,In_1974);
nand U1996 (N_1996,In_799,In_321);
and U1997 (N_1997,In_1859,In_954);
nand U1998 (N_1998,In_1296,In_1467);
or U1999 (N_1999,In_907,In_1897);
nand U2000 (N_2000,In_852,In_1708);
xor U2001 (N_2001,In_1356,In_620);
and U2002 (N_2002,In_1756,In_1097);
xor U2003 (N_2003,In_777,In_1633);
xnor U2004 (N_2004,In_1962,In_385);
and U2005 (N_2005,In_1613,In_839);
nand U2006 (N_2006,In_1122,In_1290);
and U2007 (N_2007,In_0,In_123);
or U2008 (N_2008,In_283,In_1271);
or U2009 (N_2009,In_369,In_1296);
or U2010 (N_2010,In_1458,In_1971);
and U2011 (N_2011,In_216,In_1604);
or U2012 (N_2012,In_482,In_1449);
or U2013 (N_2013,In_1000,In_864);
or U2014 (N_2014,In_494,In_1099);
and U2015 (N_2015,In_1764,In_1147);
nor U2016 (N_2016,In_673,In_907);
nand U2017 (N_2017,In_1486,In_96);
xnor U2018 (N_2018,In_497,In_1837);
nand U2019 (N_2019,In_1655,In_1290);
and U2020 (N_2020,In_857,In_461);
nor U2021 (N_2021,In_1751,In_1072);
nand U2022 (N_2022,In_416,In_1506);
or U2023 (N_2023,In_1235,In_958);
nor U2024 (N_2024,In_1926,In_688);
or U2025 (N_2025,In_336,In_853);
and U2026 (N_2026,In_251,In_1951);
nand U2027 (N_2027,In_1662,In_128);
and U2028 (N_2028,In_908,In_1778);
nand U2029 (N_2029,In_1261,In_517);
nand U2030 (N_2030,In_1189,In_149);
or U2031 (N_2031,In_684,In_276);
xnor U2032 (N_2032,In_193,In_1670);
nand U2033 (N_2033,In_84,In_355);
nor U2034 (N_2034,In_1132,In_1505);
and U2035 (N_2035,In_1665,In_1398);
nand U2036 (N_2036,In_524,In_308);
nand U2037 (N_2037,In_384,In_1859);
or U2038 (N_2038,In_467,In_1963);
nand U2039 (N_2039,In_1224,In_50);
nand U2040 (N_2040,In_1723,In_1549);
nand U2041 (N_2041,In_569,In_1006);
nand U2042 (N_2042,In_1691,In_522);
and U2043 (N_2043,In_466,In_808);
xnor U2044 (N_2044,In_1785,In_1439);
or U2045 (N_2045,In_414,In_1697);
nor U2046 (N_2046,In_1306,In_310);
nand U2047 (N_2047,In_1450,In_1308);
xnor U2048 (N_2048,In_1409,In_466);
nand U2049 (N_2049,In_47,In_12);
xnor U2050 (N_2050,In_1786,In_206);
nor U2051 (N_2051,In_877,In_1852);
and U2052 (N_2052,In_1083,In_1755);
xnor U2053 (N_2053,In_1338,In_1802);
nand U2054 (N_2054,In_1730,In_967);
xor U2055 (N_2055,In_1993,In_756);
and U2056 (N_2056,In_68,In_663);
or U2057 (N_2057,In_1412,In_441);
or U2058 (N_2058,In_1163,In_993);
xor U2059 (N_2059,In_1673,In_1046);
xor U2060 (N_2060,In_1468,In_1093);
xor U2061 (N_2061,In_542,In_982);
or U2062 (N_2062,In_295,In_1324);
nor U2063 (N_2063,In_1242,In_1560);
nor U2064 (N_2064,In_515,In_1687);
nor U2065 (N_2065,In_1013,In_546);
nand U2066 (N_2066,In_520,In_1596);
nand U2067 (N_2067,In_1774,In_1088);
nand U2068 (N_2068,In_1532,In_344);
nand U2069 (N_2069,In_1603,In_1352);
nor U2070 (N_2070,In_1352,In_1145);
or U2071 (N_2071,In_363,In_22);
or U2072 (N_2072,In_205,In_1054);
nor U2073 (N_2073,In_1113,In_542);
nand U2074 (N_2074,In_320,In_765);
xnor U2075 (N_2075,In_1161,In_38);
or U2076 (N_2076,In_465,In_166);
or U2077 (N_2077,In_675,In_534);
nand U2078 (N_2078,In_1100,In_1192);
nand U2079 (N_2079,In_127,In_582);
nand U2080 (N_2080,In_345,In_174);
and U2081 (N_2081,In_487,In_1922);
nand U2082 (N_2082,In_886,In_905);
and U2083 (N_2083,In_1576,In_666);
or U2084 (N_2084,In_918,In_1722);
and U2085 (N_2085,In_1667,In_849);
xnor U2086 (N_2086,In_1864,In_1035);
or U2087 (N_2087,In_1329,In_1497);
or U2088 (N_2088,In_557,In_76);
xnor U2089 (N_2089,In_999,In_357);
and U2090 (N_2090,In_366,In_77);
nor U2091 (N_2091,In_1091,In_866);
xnor U2092 (N_2092,In_1594,In_1757);
xor U2093 (N_2093,In_1680,In_242);
or U2094 (N_2094,In_633,In_333);
or U2095 (N_2095,In_746,In_837);
nor U2096 (N_2096,In_412,In_878);
nor U2097 (N_2097,In_833,In_1499);
nor U2098 (N_2098,In_518,In_1638);
nor U2099 (N_2099,In_270,In_1);
xnor U2100 (N_2100,In_1711,In_1336);
nand U2101 (N_2101,In_1185,In_761);
and U2102 (N_2102,In_266,In_43);
xor U2103 (N_2103,In_1850,In_607);
and U2104 (N_2104,In_1059,In_475);
or U2105 (N_2105,In_38,In_302);
xnor U2106 (N_2106,In_926,In_654);
and U2107 (N_2107,In_358,In_700);
xor U2108 (N_2108,In_478,In_183);
or U2109 (N_2109,In_344,In_1937);
or U2110 (N_2110,In_1058,In_1552);
xor U2111 (N_2111,In_120,In_1934);
or U2112 (N_2112,In_851,In_348);
and U2113 (N_2113,In_1084,In_1323);
nor U2114 (N_2114,In_736,In_1839);
nor U2115 (N_2115,In_1250,In_1308);
and U2116 (N_2116,In_1287,In_1059);
or U2117 (N_2117,In_1320,In_68);
and U2118 (N_2118,In_196,In_1158);
or U2119 (N_2119,In_1962,In_1781);
or U2120 (N_2120,In_1313,In_618);
and U2121 (N_2121,In_517,In_99);
or U2122 (N_2122,In_1698,In_220);
nor U2123 (N_2123,In_411,In_399);
nor U2124 (N_2124,In_32,In_1638);
or U2125 (N_2125,In_572,In_1262);
xor U2126 (N_2126,In_366,In_1048);
nor U2127 (N_2127,In_538,In_1826);
xnor U2128 (N_2128,In_1138,In_27);
nor U2129 (N_2129,In_601,In_1542);
nor U2130 (N_2130,In_1174,In_954);
xor U2131 (N_2131,In_1666,In_1301);
or U2132 (N_2132,In_1040,In_1961);
or U2133 (N_2133,In_1234,In_1539);
xor U2134 (N_2134,In_222,In_130);
xor U2135 (N_2135,In_1186,In_349);
or U2136 (N_2136,In_981,In_282);
nor U2137 (N_2137,In_1654,In_506);
nand U2138 (N_2138,In_865,In_923);
xor U2139 (N_2139,In_1584,In_1732);
nand U2140 (N_2140,In_1684,In_437);
xor U2141 (N_2141,In_438,In_679);
or U2142 (N_2142,In_1055,In_1799);
nand U2143 (N_2143,In_429,In_284);
xnor U2144 (N_2144,In_1126,In_449);
xnor U2145 (N_2145,In_1932,In_861);
nor U2146 (N_2146,In_498,In_1310);
nand U2147 (N_2147,In_541,In_372);
or U2148 (N_2148,In_714,In_196);
and U2149 (N_2149,In_143,In_1192);
and U2150 (N_2150,In_555,In_1634);
and U2151 (N_2151,In_528,In_40);
nor U2152 (N_2152,In_1829,In_269);
nand U2153 (N_2153,In_27,In_62);
nand U2154 (N_2154,In_1548,In_596);
and U2155 (N_2155,In_506,In_431);
or U2156 (N_2156,In_1383,In_119);
nand U2157 (N_2157,In_1549,In_95);
nor U2158 (N_2158,In_1642,In_904);
xnor U2159 (N_2159,In_1035,In_238);
nor U2160 (N_2160,In_118,In_796);
and U2161 (N_2161,In_293,In_1847);
xor U2162 (N_2162,In_1221,In_1177);
nor U2163 (N_2163,In_1549,In_594);
nor U2164 (N_2164,In_1769,In_1032);
or U2165 (N_2165,In_152,In_1819);
or U2166 (N_2166,In_255,In_1581);
and U2167 (N_2167,In_676,In_1392);
nor U2168 (N_2168,In_106,In_480);
and U2169 (N_2169,In_810,In_1512);
and U2170 (N_2170,In_1934,In_1464);
xor U2171 (N_2171,In_386,In_894);
xor U2172 (N_2172,In_1583,In_778);
and U2173 (N_2173,In_782,In_1705);
and U2174 (N_2174,In_712,In_600);
nand U2175 (N_2175,In_1338,In_1712);
or U2176 (N_2176,In_465,In_149);
or U2177 (N_2177,In_840,In_1411);
or U2178 (N_2178,In_1616,In_1998);
nor U2179 (N_2179,In_1400,In_1909);
xor U2180 (N_2180,In_93,In_1792);
nor U2181 (N_2181,In_1998,In_793);
xnor U2182 (N_2182,In_1606,In_681);
nand U2183 (N_2183,In_672,In_914);
nand U2184 (N_2184,In_791,In_1500);
nand U2185 (N_2185,In_1641,In_318);
or U2186 (N_2186,In_930,In_1242);
or U2187 (N_2187,In_1832,In_1208);
nor U2188 (N_2188,In_695,In_1674);
or U2189 (N_2189,In_740,In_1768);
xor U2190 (N_2190,In_1112,In_1913);
nand U2191 (N_2191,In_1819,In_1436);
nor U2192 (N_2192,In_1413,In_1557);
nand U2193 (N_2193,In_1343,In_1983);
and U2194 (N_2194,In_319,In_1132);
and U2195 (N_2195,In_495,In_50);
or U2196 (N_2196,In_387,In_225);
and U2197 (N_2197,In_418,In_1803);
xnor U2198 (N_2198,In_853,In_503);
nand U2199 (N_2199,In_465,In_451);
nand U2200 (N_2200,In_1991,In_1845);
nor U2201 (N_2201,In_1411,In_1912);
nor U2202 (N_2202,In_1454,In_236);
xor U2203 (N_2203,In_847,In_203);
or U2204 (N_2204,In_1792,In_414);
xor U2205 (N_2205,In_1701,In_204);
or U2206 (N_2206,In_49,In_1975);
nor U2207 (N_2207,In_692,In_797);
xor U2208 (N_2208,In_859,In_152);
and U2209 (N_2209,In_490,In_1129);
xnor U2210 (N_2210,In_3,In_1600);
or U2211 (N_2211,In_58,In_561);
nor U2212 (N_2212,In_1761,In_176);
and U2213 (N_2213,In_208,In_1531);
nand U2214 (N_2214,In_302,In_1846);
and U2215 (N_2215,In_1340,In_944);
or U2216 (N_2216,In_769,In_1574);
nand U2217 (N_2217,In_107,In_510);
or U2218 (N_2218,In_1590,In_1023);
nor U2219 (N_2219,In_1505,In_1747);
nor U2220 (N_2220,In_424,In_996);
or U2221 (N_2221,In_279,In_404);
xnor U2222 (N_2222,In_316,In_1741);
and U2223 (N_2223,In_1304,In_536);
nor U2224 (N_2224,In_1459,In_1483);
or U2225 (N_2225,In_947,In_277);
xor U2226 (N_2226,In_63,In_1503);
xnor U2227 (N_2227,In_416,In_35);
xnor U2228 (N_2228,In_1731,In_112);
nand U2229 (N_2229,In_1497,In_580);
or U2230 (N_2230,In_1895,In_1667);
or U2231 (N_2231,In_1365,In_1328);
nand U2232 (N_2232,In_1485,In_808);
xnor U2233 (N_2233,In_1715,In_677);
nand U2234 (N_2234,In_1443,In_174);
xnor U2235 (N_2235,In_894,In_517);
nor U2236 (N_2236,In_1115,In_624);
and U2237 (N_2237,In_1813,In_1754);
and U2238 (N_2238,In_41,In_1884);
nand U2239 (N_2239,In_1038,In_1348);
nor U2240 (N_2240,In_930,In_892);
nor U2241 (N_2241,In_1847,In_75);
xnor U2242 (N_2242,In_306,In_69);
nor U2243 (N_2243,In_647,In_1206);
nand U2244 (N_2244,In_1958,In_1606);
xor U2245 (N_2245,In_1950,In_1139);
xor U2246 (N_2246,In_1927,In_162);
and U2247 (N_2247,In_1427,In_461);
xnor U2248 (N_2248,In_1202,In_571);
or U2249 (N_2249,In_914,In_60);
and U2250 (N_2250,In_378,In_1);
nor U2251 (N_2251,In_990,In_1748);
and U2252 (N_2252,In_1853,In_563);
xor U2253 (N_2253,In_1200,In_322);
and U2254 (N_2254,In_1122,In_723);
nor U2255 (N_2255,In_1464,In_172);
nor U2256 (N_2256,In_1620,In_1155);
and U2257 (N_2257,In_1573,In_1024);
and U2258 (N_2258,In_129,In_1186);
xor U2259 (N_2259,In_1894,In_446);
nor U2260 (N_2260,In_454,In_841);
and U2261 (N_2261,In_67,In_425);
xor U2262 (N_2262,In_1244,In_1750);
xnor U2263 (N_2263,In_756,In_349);
and U2264 (N_2264,In_220,In_1672);
and U2265 (N_2265,In_1805,In_1585);
or U2266 (N_2266,In_1319,In_804);
xnor U2267 (N_2267,In_874,In_977);
or U2268 (N_2268,In_955,In_1074);
and U2269 (N_2269,In_571,In_89);
nand U2270 (N_2270,In_448,In_1855);
and U2271 (N_2271,In_7,In_1216);
and U2272 (N_2272,In_1474,In_1354);
and U2273 (N_2273,In_1594,In_1538);
nand U2274 (N_2274,In_1268,In_1967);
nand U2275 (N_2275,In_1553,In_478);
xnor U2276 (N_2276,In_1662,In_1049);
and U2277 (N_2277,In_231,In_1788);
or U2278 (N_2278,In_1149,In_1869);
and U2279 (N_2279,In_651,In_1988);
or U2280 (N_2280,In_285,In_1161);
and U2281 (N_2281,In_687,In_402);
nor U2282 (N_2282,In_159,In_1545);
xor U2283 (N_2283,In_873,In_438);
xor U2284 (N_2284,In_623,In_16);
nand U2285 (N_2285,In_838,In_555);
or U2286 (N_2286,In_120,In_498);
and U2287 (N_2287,In_1439,In_1861);
and U2288 (N_2288,In_8,In_1022);
nor U2289 (N_2289,In_807,In_847);
and U2290 (N_2290,In_262,In_1993);
or U2291 (N_2291,In_560,In_1348);
nor U2292 (N_2292,In_1672,In_510);
nor U2293 (N_2293,In_10,In_476);
and U2294 (N_2294,In_1256,In_672);
or U2295 (N_2295,In_1092,In_271);
xnor U2296 (N_2296,In_520,In_246);
and U2297 (N_2297,In_1464,In_790);
nand U2298 (N_2298,In_1666,In_1919);
xor U2299 (N_2299,In_343,In_1946);
and U2300 (N_2300,In_547,In_98);
nand U2301 (N_2301,In_1710,In_1421);
xor U2302 (N_2302,In_1057,In_748);
nand U2303 (N_2303,In_290,In_838);
and U2304 (N_2304,In_1641,In_1424);
xnor U2305 (N_2305,In_1288,In_1572);
xnor U2306 (N_2306,In_573,In_1715);
nand U2307 (N_2307,In_1388,In_1949);
nor U2308 (N_2308,In_296,In_116);
or U2309 (N_2309,In_415,In_450);
and U2310 (N_2310,In_1004,In_785);
nor U2311 (N_2311,In_464,In_1071);
and U2312 (N_2312,In_1298,In_1901);
xnor U2313 (N_2313,In_1077,In_458);
and U2314 (N_2314,In_1893,In_233);
and U2315 (N_2315,In_1452,In_1187);
xnor U2316 (N_2316,In_1505,In_1254);
nand U2317 (N_2317,In_140,In_521);
or U2318 (N_2318,In_3,In_1692);
or U2319 (N_2319,In_113,In_1726);
nand U2320 (N_2320,In_1825,In_1566);
xnor U2321 (N_2321,In_740,In_330);
and U2322 (N_2322,In_1945,In_968);
nor U2323 (N_2323,In_665,In_229);
xor U2324 (N_2324,In_1919,In_1720);
xnor U2325 (N_2325,In_1311,In_1688);
nor U2326 (N_2326,In_1515,In_1823);
nor U2327 (N_2327,In_335,In_1649);
and U2328 (N_2328,In_865,In_1000);
nor U2329 (N_2329,In_1554,In_1426);
and U2330 (N_2330,In_1890,In_586);
nand U2331 (N_2331,In_1358,In_1495);
xnor U2332 (N_2332,In_201,In_1924);
or U2333 (N_2333,In_891,In_1104);
or U2334 (N_2334,In_36,In_927);
and U2335 (N_2335,In_67,In_758);
xnor U2336 (N_2336,In_194,In_1021);
and U2337 (N_2337,In_1607,In_1218);
and U2338 (N_2338,In_1571,In_1286);
nand U2339 (N_2339,In_955,In_969);
xor U2340 (N_2340,In_957,In_1506);
nor U2341 (N_2341,In_996,In_154);
or U2342 (N_2342,In_1913,In_1220);
xnor U2343 (N_2343,In_1458,In_1115);
nand U2344 (N_2344,In_1967,In_80);
nor U2345 (N_2345,In_1464,In_779);
nand U2346 (N_2346,In_772,In_851);
and U2347 (N_2347,In_1393,In_1213);
or U2348 (N_2348,In_1929,In_1254);
xor U2349 (N_2349,In_1671,In_1871);
xor U2350 (N_2350,In_1778,In_542);
or U2351 (N_2351,In_837,In_1750);
xnor U2352 (N_2352,In_737,In_1650);
or U2353 (N_2353,In_127,In_1988);
nor U2354 (N_2354,In_1042,In_1890);
nand U2355 (N_2355,In_1196,In_1724);
nand U2356 (N_2356,In_1149,In_669);
or U2357 (N_2357,In_1530,In_516);
or U2358 (N_2358,In_1983,In_254);
or U2359 (N_2359,In_1179,In_497);
or U2360 (N_2360,In_1464,In_182);
nor U2361 (N_2361,In_795,In_585);
nor U2362 (N_2362,In_222,In_873);
and U2363 (N_2363,In_1088,In_350);
and U2364 (N_2364,In_569,In_366);
nor U2365 (N_2365,In_1379,In_936);
or U2366 (N_2366,In_586,In_1588);
or U2367 (N_2367,In_1605,In_461);
or U2368 (N_2368,In_1559,In_1695);
or U2369 (N_2369,In_1247,In_1326);
or U2370 (N_2370,In_910,In_1984);
and U2371 (N_2371,In_1486,In_39);
xor U2372 (N_2372,In_966,In_1425);
and U2373 (N_2373,In_523,In_1888);
xnor U2374 (N_2374,In_1652,In_325);
nand U2375 (N_2375,In_1474,In_960);
nor U2376 (N_2376,In_1359,In_1586);
or U2377 (N_2377,In_305,In_1022);
nand U2378 (N_2378,In_956,In_380);
or U2379 (N_2379,In_1831,In_1988);
or U2380 (N_2380,In_675,In_1798);
xor U2381 (N_2381,In_616,In_1698);
nor U2382 (N_2382,In_1967,In_693);
xor U2383 (N_2383,In_1129,In_743);
nand U2384 (N_2384,In_804,In_558);
nand U2385 (N_2385,In_1996,In_1329);
and U2386 (N_2386,In_210,In_1995);
or U2387 (N_2387,In_1105,In_774);
nand U2388 (N_2388,In_907,In_698);
nor U2389 (N_2389,In_307,In_1382);
xor U2390 (N_2390,In_535,In_243);
nand U2391 (N_2391,In_1692,In_951);
or U2392 (N_2392,In_374,In_810);
nand U2393 (N_2393,In_660,In_135);
or U2394 (N_2394,In_149,In_477);
or U2395 (N_2395,In_1579,In_261);
and U2396 (N_2396,In_1294,In_1711);
nor U2397 (N_2397,In_682,In_240);
xor U2398 (N_2398,In_283,In_16);
and U2399 (N_2399,In_1312,In_344);
xor U2400 (N_2400,In_1197,In_1952);
nor U2401 (N_2401,In_315,In_1064);
xnor U2402 (N_2402,In_315,In_1358);
and U2403 (N_2403,In_1517,In_1220);
or U2404 (N_2404,In_1204,In_1261);
nor U2405 (N_2405,In_1216,In_230);
nor U2406 (N_2406,In_851,In_956);
or U2407 (N_2407,In_1904,In_86);
nor U2408 (N_2408,In_1182,In_1111);
and U2409 (N_2409,In_1859,In_806);
and U2410 (N_2410,In_1180,In_112);
or U2411 (N_2411,In_297,In_868);
or U2412 (N_2412,In_1575,In_55);
or U2413 (N_2413,In_459,In_189);
xor U2414 (N_2414,In_1297,In_1331);
xnor U2415 (N_2415,In_1115,In_1620);
or U2416 (N_2416,In_822,In_1660);
or U2417 (N_2417,In_1315,In_1859);
nor U2418 (N_2418,In_1553,In_1451);
and U2419 (N_2419,In_1970,In_502);
xnor U2420 (N_2420,In_218,In_1806);
nor U2421 (N_2421,In_479,In_509);
and U2422 (N_2422,In_1760,In_1362);
xnor U2423 (N_2423,In_466,In_1203);
xnor U2424 (N_2424,In_89,In_1716);
and U2425 (N_2425,In_145,In_255);
nor U2426 (N_2426,In_188,In_410);
or U2427 (N_2427,In_1336,In_769);
or U2428 (N_2428,In_1472,In_832);
nor U2429 (N_2429,In_382,In_1925);
xnor U2430 (N_2430,In_1441,In_755);
xor U2431 (N_2431,In_812,In_61);
or U2432 (N_2432,In_356,In_942);
and U2433 (N_2433,In_1842,In_1411);
nand U2434 (N_2434,In_26,In_1426);
or U2435 (N_2435,In_84,In_140);
or U2436 (N_2436,In_285,In_1605);
nand U2437 (N_2437,In_1880,In_1363);
nand U2438 (N_2438,In_1579,In_1078);
nand U2439 (N_2439,In_1292,In_1838);
and U2440 (N_2440,In_1415,In_1745);
and U2441 (N_2441,In_1927,In_1348);
nand U2442 (N_2442,In_106,In_1660);
or U2443 (N_2443,In_695,In_1064);
and U2444 (N_2444,In_14,In_516);
nand U2445 (N_2445,In_1660,In_610);
or U2446 (N_2446,In_992,In_20);
xor U2447 (N_2447,In_831,In_1996);
nand U2448 (N_2448,In_1723,In_396);
xnor U2449 (N_2449,In_457,In_1400);
nand U2450 (N_2450,In_1733,In_1134);
and U2451 (N_2451,In_1642,In_1906);
nor U2452 (N_2452,In_1992,In_225);
nor U2453 (N_2453,In_1152,In_977);
xor U2454 (N_2454,In_497,In_547);
nand U2455 (N_2455,In_1602,In_860);
nand U2456 (N_2456,In_464,In_1726);
xor U2457 (N_2457,In_165,In_1766);
nand U2458 (N_2458,In_1698,In_271);
nand U2459 (N_2459,In_1228,In_546);
nor U2460 (N_2460,In_1001,In_1787);
or U2461 (N_2461,In_996,In_808);
nand U2462 (N_2462,In_226,In_1222);
nand U2463 (N_2463,In_710,In_1073);
nor U2464 (N_2464,In_1934,In_1305);
xnor U2465 (N_2465,In_420,In_1563);
or U2466 (N_2466,In_1268,In_1926);
nand U2467 (N_2467,In_536,In_728);
xnor U2468 (N_2468,In_436,In_203);
nand U2469 (N_2469,In_827,In_905);
or U2470 (N_2470,In_1227,In_1359);
nor U2471 (N_2471,In_733,In_1065);
or U2472 (N_2472,In_406,In_768);
nor U2473 (N_2473,In_237,In_808);
and U2474 (N_2474,In_932,In_1070);
nor U2475 (N_2475,In_1793,In_1178);
xnor U2476 (N_2476,In_1779,In_266);
and U2477 (N_2477,In_1614,In_1016);
and U2478 (N_2478,In_849,In_220);
or U2479 (N_2479,In_1718,In_1588);
nor U2480 (N_2480,In_880,In_1871);
or U2481 (N_2481,In_132,In_860);
nor U2482 (N_2482,In_1867,In_463);
nor U2483 (N_2483,In_837,In_1041);
nand U2484 (N_2484,In_19,In_584);
xnor U2485 (N_2485,In_978,In_1814);
nand U2486 (N_2486,In_1617,In_1781);
or U2487 (N_2487,In_342,In_971);
nand U2488 (N_2488,In_1402,In_474);
and U2489 (N_2489,In_983,In_147);
nand U2490 (N_2490,In_776,In_607);
xor U2491 (N_2491,In_1029,In_489);
or U2492 (N_2492,In_851,In_469);
nor U2493 (N_2493,In_29,In_538);
nor U2494 (N_2494,In_1338,In_891);
or U2495 (N_2495,In_1028,In_1754);
or U2496 (N_2496,In_1113,In_1860);
nand U2497 (N_2497,In_1624,In_1438);
nand U2498 (N_2498,In_1802,In_751);
nand U2499 (N_2499,In_754,In_301);
and U2500 (N_2500,In_577,In_1249);
xnor U2501 (N_2501,In_1028,In_37);
xnor U2502 (N_2502,In_393,In_1783);
and U2503 (N_2503,In_405,In_914);
and U2504 (N_2504,In_1383,In_1884);
nor U2505 (N_2505,In_9,In_1110);
nand U2506 (N_2506,In_1662,In_957);
nor U2507 (N_2507,In_440,In_368);
nor U2508 (N_2508,In_36,In_1796);
nor U2509 (N_2509,In_1460,In_1921);
or U2510 (N_2510,In_1300,In_36);
xor U2511 (N_2511,In_1078,In_716);
and U2512 (N_2512,In_732,In_615);
nor U2513 (N_2513,In_894,In_1252);
or U2514 (N_2514,In_359,In_1712);
nand U2515 (N_2515,In_486,In_1818);
nor U2516 (N_2516,In_1563,In_910);
nand U2517 (N_2517,In_515,In_927);
nor U2518 (N_2518,In_1592,In_20);
or U2519 (N_2519,In_627,In_1602);
xor U2520 (N_2520,In_1381,In_634);
xor U2521 (N_2521,In_560,In_471);
nand U2522 (N_2522,In_681,In_1850);
and U2523 (N_2523,In_1787,In_1736);
nor U2524 (N_2524,In_48,In_1764);
or U2525 (N_2525,In_1278,In_1441);
nor U2526 (N_2526,In_1448,In_1111);
xor U2527 (N_2527,In_1021,In_389);
or U2528 (N_2528,In_784,In_1093);
nand U2529 (N_2529,In_159,In_723);
or U2530 (N_2530,In_112,In_1074);
and U2531 (N_2531,In_1583,In_1913);
nand U2532 (N_2532,In_601,In_807);
nand U2533 (N_2533,In_20,In_1328);
nor U2534 (N_2534,In_629,In_1940);
nand U2535 (N_2535,In_378,In_151);
xnor U2536 (N_2536,In_282,In_1171);
or U2537 (N_2537,In_1774,In_464);
nand U2538 (N_2538,In_408,In_1031);
nor U2539 (N_2539,In_583,In_96);
or U2540 (N_2540,In_267,In_590);
nor U2541 (N_2541,In_276,In_85);
or U2542 (N_2542,In_235,In_1269);
xor U2543 (N_2543,In_1558,In_1564);
and U2544 (N_2544,In_1601,In_779);
xor U2545 (N_2545,In_857,In_519);
or U2546 (N_2546,In_845,In_1874);
or U2547 (N_2547,In_533,In_1242);
nand U2548 (N_2548,In_136,In_1982);
nor U2549 (N_2549,In_152,In_1125);
or U2550 (N_2550,In_936,In_649);
or U2551 (N_2551,In_1464,In_1258);
nand U2552 (N_2552,In_1675,In_135);
nor U2553 (N_2553,In_786,In_442);
xnor U2554 (N_2554,In_1160,In_550);
or U2555 (N_2555,In_1998,In_1023);
and U2556 (N_2556,In_889,In_1387);
or U2557 (N_2557,In_700,In_720);
and U2558 (N_2558,In_229,In_1600);
or U2559 (N_2559,In_1723,In_917);
or U2560 (N_2560,In_1262,In_1370);
xor U2561 (N_2561,In_231,In_515);
and U2562 (N_2562,In_741,In_330);
xor U2563 (N_2563,In_1,In_1157);
nor U2564 (N_2564,In_1128,In_436);
nor U2565 (N_2565,In_880,In_879);
nand U2566 (N_2566,In_1468,In_697);
nor U2567 (N_2567,In_971,In_871);
nor U2568 (N_2568,In_1538,In_1991);
or U2569 (N_2569,In_371,In_341);
nor U2570 (N_2570,In_721,In_1433);
nand U2571 (N_2571,In_979,In_1549);
and U2572 (N_2572,In_1939,In_454);
xor U2573 (N_2573,In_297,In_765);
or U2574 (N_2574,In_956,In_1284);
nand U2575 (N_2575,In_422,In_506);
or U2576 (N_2576,In_942,In_957);
and U2577 (N_2577,In_682,In_1418);
or U2578 (N_2578,In_1515,In_600);
xor U2579 (N_2579,In_1026,In_109);
nand U2580 (N_2580,In_94,In_1635);
nand U2581 (N_2581,In_1014,In_1789);
nand U2582 (N_2582,In_1106,In_910);
nor U2583 (N_2583,In_1966,In_38);
nor U2584 (N_2584,In_1971,In_1436);
and U2585 (N_2585,In_336,In_743);
nand U2586 (N_2586,In_1218,In_585);
nand U2587 (N_2587,In_1294,In_171);
xor U2588 (N_2588,In_1966,In_1395);
and U2589 (N_2589,In_1335,In_1502);
xnor U2590 (N_2590,In_421,In_61);
and U2591 (N_2591,In_1718,In_608);
or U2592 (N_2592,In_1621,In_1019);
nor U2593 (N_2593,In_1352,In_1271);
or U2594 (N_2594,In_1612,In_887);
or U2595 (N_2595,In_1496,In_1361);
xnor U2596 (N_2596,In_1852,In_550);
nand U2597 (N_2597,In_1132,In_941);
nor U2598 (N_2598,In_793,In_648);
xor U2599 (N_2599,In_749,In_1093);
nand U2600 (N_2600,In_102,In_1716);
nand U2601 (N_2601,In_427,In_746);
nand U2602 (N_2602,In_1199,In_1784);
nor U2603 (N_2603,In_1756,In_1621);
and U2604 (N_2604,In_584,In_855);
nor U2605 (N_2605,In_600,In_1941);
or U2606 (N_2606,In_184,In_70);
nor U2607 (N_2607,In_1375,In_1756);
and U2608 (N_2608,In_1808,In_1836);
or U2609 (N_2609,In_475,In_727);
or U2610 (N_2610,In_1234,In_889);
nand U2611 (N_2611,In_217,In_1901);
nor U2612 (N_2612,In_591,In_1743);
xnor U2613 (N_2613,In_829,In_1679);
or U2614 (N_2614,In_1701,In_1502);
and U2615 (N_2615,In_984,In_592);
nand U2616 (N_2616,In_502,In_821);
xor U2617 (N_2617,In_392,In_141);
nor U2618 (N_2618,In_308,In_1956);
nand U2619 (N_2619,In_1550,In_178);
nand U2620 (N_2620,In_1502,In_1141);
nor U2621 (N_2621,In_1813,In_49);
and U2622 (N_2622,In_163,In_816);
and U2623 (N_2623,In_729,In_744);
or U2624 (N_2624,In_805,In_583);
xnor U2625 (N_2625,In_815,In_1312);
nor U2626 (N_2626,In_463,In_45);
nor U2627 (N_2627,In_219,In_400);
xnor U2628 (N_2628,In_821,In_498);
nand U2629 (N_2629,In_87,In_1900);
nor U2630 (N_2630,In_1278,In_702);
and U2631 (N_2631,In_669,In_1774);
or U2632 (N_2632,In_780,In_1251);
and U2633 (N_2633,In_1542,In_181);
xor U2634 (N_2634,In_1186,In_935);
nand U2635 (N_2635,In_570,In_1690);
nand U2636 (N_2636,In_1601,In_1036);
nor U2637 (N_2637,In_1240,In_623);
xor U2638 (N_2638,In_289,In_1947);
and U2639 (N_2639,In_719,In_128);
xor U2640 (N_2640,In_1666,In_1824);
nand U2641 (N_2641,In_608,In_1438);
or U2642 (N_2642,In_26,In_1869);
and U2643 (N_2643,In_1814,In_971);
xnor U2644 (N_2644,In_222,In_836);
or U2645 (N_2645,In_1191,In_767);
xor U2646 (N_2646,In_1447,In_946);
xor U2647 (N_2647,In_84,In_365);
nand U2648 (N_2648,In_1447,In_266);
and U2649 (N_2649,In_1289,In_458);
nand U2650 (N_2650,In_91,In_1814);
nand U2651 (N_2651,In_615,In_827);
xnor U2652 (N_2652,In_984,In_203);
and U2653 (N_2653,In_478,In_28);
nor U2654 (N_2654,In_770,In_1124);
xor U2655 (N_2655,In_102,In_1620);
nand U2656 (N_2656,In_747,In_815);
nand U2657 (N_2657,In_1628,In_1402);
or U2658 (N_2658,In_1707,In_919);
nor U2659 (N_2659,In_234,In_1665);
xnor U2660 (N_2660,In_1286,In_69);
xor U2661 (N_2661,In_989,In_186);
nor U2662 (N_2662,In_1799,In_174);
nand U2663 (N_2663,In_280,In_1824);
or U2664 (N_2664,In_486,In_1406);
and U2665 (N_2665,In_279,In_443);
nor U2666 (N_2666,In_1468,In_1661);
nor U2667 (N_2667,In_1946,In_111);
xor U2668 (N_2668,In_1724,In_515);
and U2669 (N_2669,In_1838,In_1221);
and U2670 (N_2670,In_1356,In_1380);
xor U2671 (N_2671,In_663,In_802);
nand U2672 (N_2672,In_438,In_1109);
and U2673 (N_2673,In_166,In_68);
xor U2674 (N_2674,In_463,In_1514);
and U2675 (N_2675,In_134,In_317);
and U2676 (N_2676,In_562,In_1538);
and U2677 (N_2677,In_732,In_1333);
and U2678 (N_2678,In_1646,In_1668);
or U2679 (N_2679,In_1312,In_1654);
nand U2680 (N_2680,In_646,In_1380);
nand U2681 (N_2681,In_1528,In_951);
nand U2682 (N_2682,In_1211,In_1105);
xor U2683 (N_2683,In_36,In_1688);
nor U2684 (N_2684,In_1528,In_207);
nand U2685 (N_2685,In_1790,In_1160);
xnor U2686 (N_2686,In_1168,In_1109);
and U2687 (N_2687,In_1465,In_150);
nand U2688 (N_2688,In_398,In_8);
or U2689 (N_2689,In_1134,In_1436);
or U2690 (N_2690,In_1179,In_449);
xnor U2691 (N_2691,In_1173,In_1569);
and U2692 (N_2692,In_1791,In_1403);
nand U2693 (N_2693,In_1307,In_1432);
or U2694 (N_2694,In_155,In_1318);
or U2695 (N_2695,In_1930,In_164);
xnor U2696 (N_2696,In_1259,In_183);
nor U2697 (N_2697,In_1581,In_465);
or U2698 (N_2698,In_1427,In_1453);
nor U2699 (N_2699,In_549,In_191);
nor U2700 (N_2700,In_1413,In_1351);
nor U2701 (N_2701,In_990,In_1031);
nand U2702 (N_2702,In_1098,In_1371);
and U2703 (N_2703,In_461,In_1236);
nor U2704 (N_2704,In_1481,In_1645);
xnor U2705 (N_2705,In_1252,In_1504);
nor U2706 (N_2706,In_1794,In_39);
or U2707 (N_2707,In_1529,In_235);
nor U2708 (N_2708,In_1106,In_1032);
or U2709 (N_2709,In_1293,In_1188);
nor U2710 (N_2710,In_1811,In_638);
nand U2711 (N_2711,In_718,In_122);
or U2712 (N_2712,In_419,In_252);
xor U2713 (N_2713,In_1580,In_1183);
nand U2714 (N_2714,In_1276,In_77);
xor U2715 (N_2715,In_1470,In_433);
xnor U2716 (N_2716,In_57,In_1903);
or U2717 (N_2717,In_1292,In_1342);
nor U2718 (N_2718,In_53,In_1551);
nor U2719 (N_2719,In_983,In_583);
xor U2720 (N_2720,In_384,In_442);
nand U2721 (N_2721,In_306,In_1427);
or U2722 (N_2722,In_316,In_506);
xnor U2723 (N_2723,In_1840,In_587);
and U2724 (N_2724,In_1100,In_1213);
or U2725 (N_2725,In_1787,In_1071);
nor U2726 (N_2726,In_1977,In_342);
xor U2727 (N_2727,In_1977,In_300);
nor U2728 (N_2728,In_1202,In_108);
xnor U2729 (N_2729,In_1806,In_1248);
xor U2730 (N_2730,In_1994,In_1586);
or U2731 (N_2731,In_560,In_670);
or U2732 (N_2732,In_8,In_180);
or U2733 (N_2733,In_1251,In_1559);
and U2734 (N_2734,In_962,In_1748);
nand U2735 (N_2735,In_329,In_939);
nand U2736 (N_2736,In_596,In_1504);
xnor U2737 (N_2737,In_528,In_1580);
or U2738 (N_2738,In_1409,In_1274);
and U2739 (N_2739,In_592,In_893);
or U2740 (N_2740,In_1086,In_1766);
xor U2741 (N_2741,In_1499,In_1352);
and U2742 (N_2742,In_467,In_932);
nand U2743 (N_2743,In_1469,In_1495);
or U2744 (N_2744,In_1835,In_1209);
nand U2745 (N_2745,In_939,In_149);
nor U2746 (N_2746,In_1835,In_1849);
or U2747 (N_2747,In_223,In_1426);
xnor U2748 (N_2748,In_766,In_1420);
or U2749 (N_2749,In_139,In_454);
and U2750 (N_2750,In_456,In_117);
nor U2751 (N_2751,In_1212,In_1875);
nor U2752 (N_2752,In_5,In_812);
xnor U2753 (N_2753,In_339,In_572);
and U2754 (N_2754,In_1331,In_1492);
xnor U2755 (N_2755,In_305,In_435);
and U2756 (N_2756,In_1867,In_1195);
nor U2757 (N_2757,In_1090,In_74);
nand U2758 (N_2758,In_1312,In_8);
nand U2759 (N_2759,In_1145,In_197);
or U2760 (N_2760,In_741,In_22);
xnor U2761 (N_2761,In_1619,In_1197);
nor U2762 (N_2762,In_1785,In_1634);
and U2763 (N_2763,In_140,In_511);
xor U2764 (N_2764,In_1099,In_912);
or U2765 (N_2765,In_1023,In_1186);
nor U2766 (N_2766,In_1482,In_1123);
xor U2767 (N_2767,In_855,In_739);
nand U2768 (N_2768,In_1767,In_1579);
and U2769 (N_2769,In_1305,In_1219);
xnor U2770 (N_2770,In_1238,In_476);
nand U2771 (N_2771,In_513,In_331);
nor U2772 (N_2772,In_746,In_1594);
or U2773 (N_2773,In_361,In_1017);
xnor U2774 (N_2774,In_1317,In_700);
or U2775 (N_2775,In_1822,In_1356);
xor U2776 (N_2776,In_1450,In_1000);
nand U2777 (N_2777,In_1498,In_1817);
nand U2778 (N_2778,In_1248,In_574);
xor U2779 (N_2779,In_789,In_606);
and U2780 (N_2780,In_346,In_1212);
and U2781 (N_2781,In_625,In_321);
nand U2782 (N_2782,In_16,In_1375);
nand U2783 (N_2783,In_419,In_630);
and U2784 (N_2784,In_542,In_1761);
nand U2785 (N_2785,In_1103,In_54);
and U2786 (N_2786,In_401,In_628);
or U2787 (N_2787,In_300,In_1455);
nor U2788 (N_2788,In_1039,In_986);
xor U2789 (N_2789,In_1390,In_276);
nor U2790 (N_2790,In_828,In_1054);
nor U2791 (N_2791,In_1824,In_749);
xnor U2792 (N_2792,In_780,In_821);
nand U2793 (N_2793,In_1723,In_1863);
nand U2794 (N_2794,In_705,In_1445);
nor U2795 (N_2795,In_1178,In_1573);
and U2796 (N_2796,In_1875,In_526);
and U2797 (N_2797,In_1191,In_999);
and U2798 (N_2798,In_635,In_586);
or U2799 (N_2799,In_1315,In_1045);
and U2800 (N_2800,In_23,In_1747);
xnor U2801 (N_2801,In_738,In_418);
and U2802 (N_2802,In_48,In_1928);
nand U2803 (N_2803,In_1303,In_1888);
nand U2804 (N_2804,In_479,In_217);
and U2805 (N_2805,In_1728,In_401);
nand U2806 (N_2806,In_302,In_681);
xnor U2807 (N_2807,In_575,In_1502);
xnor U2808 (N_2808,In_1136,In_1483);
xnor U2809 (N_2809,In_1989,In_1590);
nor U2810 (N_2810,In_1642,In_760);
and U2811 (N_2811,In_1123,In_99);
and U2812 (N_2812,In_1928,In_1530);
or U2813 (N_2813,In_1455,In_1679);
or U2814 (N_2814,In_315,In_230);
or U2815 (N_2815,In_225,In_957);
or U2816 (N_2816,In_120,In_489);
xnor U2817 (N_2817,In_1028,In_1986);
or U2818 (N_2818,In_617,In_83);
xnor U2819 (N_2819,In_1671,In_1395);
xor U2820 (N_2820,In_1026,In_1375);
and U2821 (N_2821,In_222,In_1519);
and U2822 (N_2822,In_873,In_279);
and U2823 (N_2823,In_1292,In_1493);
and U2824 (N_2824,In_149,In_733);
xnor U2825 (N_2825,In_36,In_1);
nor U2826 (N_2826,In_371,In_991);
nor U2827 (N_2827,In_1475,In_413);
nor U2828 (N_2828,In_1192,In_1742);
nor U2829 (N_2829,In_1440,In_448);
or U2830 (N_2830,In_772,In_1945);
or U2831 (N_2831,In_1470,In_1150);
or U2832 (N_2832,In_826,In_1434);
nor U2833 (N_2833,In_312,In_848);
nor U2834 (N_2834,In_1758,In_1749);
nor U2835 (N_2835,In_1230,In_1733);
or U2836 (N_2836,In_1159,In_115);
nand U2837 (N_2837,In_621,In_1397);
xnor U2838 (N_2838,In_819,In_71);
xnor U2839 (N_2839,In_1109,In_577);
and U2840 (N_2840,In_1935,In_594);
and U2841 (N_2841,In_483,In_1930);
xor U2842 (N_2842,In_1184,In_714);
or U2843 (N_2843,In_1362,In_1815);
nand U2844 (N_2844,In_1031,In_164);
xnor U2845 (N_2845,In_1056,In_926);
and U2846 (N_2846,In_1604,In_1281);
nand U2847 (N_2847,In_178,In_1841);
nor U2848 (N_2848,In_832,In_1174);
nor U2849 (N_2849,In_685,In_262);
nand U2850 (N_2850,In_1360,In_1372);
and U2851 (N_2851,In_1975,In_1056);
nand U2852 (N_2852,In_1707,In_1357);
nand U2853 (N_2853,In_78,In_1497);
nand U2854 (N_2854,In_1586,In_334);
nand U2855 (N_2855,In_1923,In_6);
xnor U2856 (N_2856,In_1408,In_161);
nand U2857 (N_2857,In_817,In_800);
or U2858 (N_2858,In_1533,In_12);
nor U2859 (N_2859,In_134,In_1658);
nand U2860 (N_2860,In_46,In_12);
nand U2861 (N_2861,In_202,In_1071);
nand U2862 (N_2862,In_1356,In_319);
xnor U2863 (N_2863,In_1384,In_1927);
nor U2864 (N_2864,In_270,In_1845);
nand U2865 (N_2865,In_1853,In_437);
xnor U2866 (N_2866,In_1282,In_1367);
nor U2867 (N_2867,In_1909,In_1608);
or U2868 (N_2868,In_590,In_506);
or U2869 (N_2869,In_333,In_1136);
nor U2870 (N_2870,In_638,In_816);
or U2871 (N_2871,In_1870,In_1628);
xor U2872 (N_2872,In_1146,In_1117);
nor U2873 (N_2873,In_582,In_178);
and U2874 (N_2874,In_1150,In_458);
nor U2875 (N_2875,In_993,In_393);
xor U2876 (N_2876,In_707,In_666);
nand U2877 (N_2877,In_47,In_23);
or U2878 (N_2878,In_1455,In_994);
nor U2879 (N_2879,In_1885,In_62);
or U2880 (N_2880,In_204,In_17);
and U2881 (N_2881,In_1315,In_158);
and U2882 (N_2882,In_743,In_1672);
or U2883 (N_2883,In_1247,In_1748);
xnor U2884 (N_2884,In_353,In_1643);
xor U2885 (N_2885,In_135,In_1014);
nand U2886 (N_2886,In_376,In_802);
nor U2887 (N_2887,In_605,In_1355);
xnor U2888 (N_2888,In_1646,In_1301);
xnor U2889 (N_2889,In_1303,In_1508);
and U2890 (N_2890,In_73,In_325);
or U2891 (N_2891,In_504,In_690);
or U2892 (N_2892,In_193,In_1169);
and U2893 (N_2893,In_788,In_1740);
nand U2894 (N_2894,In_978,In_1474);
and U2895 (N_2895,In_716,In_225);
xor U2896 (N_2896,In_1900,In_120);
nor U2897 (N_2897,In_1730,In_1261);
and U2898 (N_2898,In_150,In_133);
and U2899 (N_2899,In_72,In_1393);
or U2900 (N_2900,In_1884,In_983);
nand U2901 (N_2901,In_1746,In_1684);
nand U2902 (N_2902,In_86,In_1046);
or U2903 (N_2903,In_930,In_776);
nand U2904 (N_2904,In_1355,In_1442);
and U2905 (N_2905,In_1722,In_1978);
and U2906 (N_2906,In_1438,In_281);
xnor U2907 (N_2907,In_724,In_432);
nand U2908 (N_2908,In_1097,In_397);
nor U2909 (N_2909,In_1585,In_1439);
and U2910 (N_2910,In_834,In_1371);
and U2911 (N_2911,In_1700,In_0);
and U2912 (N_2912,In_1912,In_230);
and U2913 (N_2913,In_676,In_1336);
nor U2914 (N_2914,In_1490,In_1657);
and U2915 (N_2915,In_1094,In_121);
xnor U2916 (N_2916,In_1659,In_35);
or U2917 (N_2917,In_373,In_395);
nand U2918 (N_2918,In_690,In_375);
or U2919 (N_2919,In_1002,In_832);
or U2920 (N_2920,In_1423,In_906);
nand U2921 (N_2921,In_486,In_1185);
xnor U2922 (N_2922,In_393,In_1199);
and U2923 (N_2923,In_1039,In_849);
xor U2924 (N_2924,In_1918,In_1687);
xnor U2925 (N_2925,In_570,In_1917);
or U2926 (N_2926,In_493,In_1757);
or U2927 (N_2927,In_1363,In_273);
nor U2928 (N_2928,In_1145,In_1869);
nand U2929 (N_2929,In_346,In_1837);
nor U2930 (N_2930,In_1741,In_295);
nor U2931 (N_2931,In_596,In_872);
or U2932 (N_2932,In_1614,In_1271);
nand U2933 (N_2933,In_1523,In_218);
or U2934 (N_2934,In_37,In_1603);
nand U2935 (N_2935,In_654,In_861);
nor U2936 (N_2936,In_1883,In_1630);
xor U2937 (N_2937,In_58,In_334);
and U2938 (N_2938,In_172,In_1751);
nand U2939 (N_2939,In_952,In_1068);
or U2940 (N_2940,In_1237,In_590);
nand U2941 (N_2941,In_399,In_1692);
and U2942 (N_2942,In_1164,In_1655);
and U2943 (N_2943,In_570,In_912);
xor U2944 (N_2944,In_1170,In_558);
or U2945 (N_2945,In_1928,In_1211);
and U2946 (N_2946,In_1447,In_1149);
nor U2947 (N_2947,In_1255,In_938);
nand U2948 (N_2948,In_231,In_800);
and U2949 (N_2949,In_1361,In_854);
nor U2950 (N_2950,In_610,In_1042);
or U2951 (N_2951,In_1816,In_1538);
and U2952 (N_2952,In_0,In_75);
and U2953 (N_2953,In_912,In_1154);
nand U2954 (N_2954,In_912,In_1919);
xor U2955 (N_2955,In_771,In_407);
xor U2956 (N_2956,In_164,In_1257);
or U2957 (N_2957,In_1157,In_708);
or U2958 (N_2958,In_1812,In_847);
xor U2959 (N_2959,In_631,In_568);
or U2960 (N_2960,In_1560,In_1259);
nor U2961 (N_2961,In_532,In_433);
nor U2962 (N_2962,In_55,In_1657);
nand U2963 (N_2963,In_198,In_1317);
nor U2964 (N_2964,In_1067,In_1397);
or U2965 (N_2965,In_249,In_1743);
nor U2966 (N_2966,In_1334,In_1446);
and U2967 (N_2967,In_1405,In_1713);
nor U2968 (N_2968,In_1890,In_60);
nand U2969 (N_2969,In_498,In_1564);
or U2970 (N_2970,In_1944,In_1615);
and U2971 (N_2971,In_1881,In_1126);
and U2972 (N_2972,In_1508,In_222);
xnor U2973 (N_2973,In_74,In_605);
or U2974 (N_2974,In_517,In_1104);
and U2975 (N_2975,In_576,In_63);
xor U2976 (N_2976,In_1096,In_1012);
and U2977 (N_2977,In_250,In_1087);
nor U2978 (N_2978,In_350,In_1179);
xor U2979 (N_2979,In_1534,In_601);
nand U2980 (N_2980,In_1314,In_69);
xor U2981 (N_2981,In_119,In_545);
xnor U2982 (N_2982,In_1035,In_1090);
or U2983 (N_2983,In_1760,In_1575);
xor U2984 (N_2984,In_1317,In_1280);
or U2985 (N_2985,In_1876,In_168);
or U2986 (N_2986,In_459,In_1529);
nor U2987 (N_2987,In_1446,In_1367);
nand U2988 (N_2988,In_1942,In_273);
or U2989 (N_2989,In_1678,In_1083);
xnor U2990 (N_2990,In_1047,In_433);
or U2991 (N_2991,In_1677,In_1933);
xnor U2992 (N_2992,In_1924,In_813);
xor U2993 (N_2993,In_388,In_1575);
nand U2994 (N_2994,In_1704,In_1451);
nand U2995 (N_2995,In_302,In_1219);
or U2996 (N_2996,In_813,In_905);
nand U2997 (N_2997,In_381,In_1347);
xor U2998 (N_2998,In_268,In_1875);
and U2999 (N_2999,In_1558,In_492);
nor U3000 (N_3000,In_1,In_1034);
nand U3001 (N_3001,In_1249,In_1519);
nand U3002 (N_3002,In_1232,In_491);
xor U3003 (N_3003,In_1549,In_1615);
nand U3004 (N_3004,In_1757,In_376);
or U3005 (N_3005,In_1843,In_1410);
nand U3006 (N_3006,In_138,In_1589);
or U3007 (N_3007,In_414,In_1438);
xnor U3008 (N_3008,In_90,In_983);
nand U3009 (N_3009,In_123,In_857);
nand U3010 (N_3010,In_724,In_1592);
nor U3011 (N_3011,In_412,In_1297);
nand U3012 (N_3012,In_183,In_191);
and U3013 (N_3013,In_1001,In_1754);
xnor U3014 (N_3014,In_496,In_952);
xnor U3015 (N_3015,In_816,In_1891);
xnor U3016 (N_3016,In_395,In_1479);
nand U3017 (N_3017,In_1482,In_1236);
and U3018 (N_3018,In_241,In_119);
or U3019 (N_3019,In_410,In_57);
nand U3020 (N_3020,In_543,In_78);
nor U3021 (N_3021,In_1078,In_1985);
xor U3022 (N_3022,In_1108,In_504);
and U3023 (N_3023,In_1264,In_681);
or U3024 (N_3024,In_1586,In_336);
or U3025 (N_3025,In_1250,In_684);
nor U3026 (N_3026,In_1829,In_648);
xor U3027 (N_3027,In_92,In_1235);
nand U3028 (N_3028,In_683,In_1808);
nor U3029 (N_3029,In_1909,In_1925);
nor U3030 (N_3030,In_1135,In_1435);
nand U3031 (N_3031,In_1603,In_1542);
and U3032 (N_3032,In_652,In_210);
or U3033 (N_3033,In_897,In_44);
xor U3034 (N_3034,In_1831,In_1562);
nor U3035 (N_3035,In_1045,In_877);
xnor U3036 (N_3036,In_870,In_1877);
nor U3037 (N_3037,In_1469,In_235);
nand U3038 (N_3038,In_955,In_1030);
xor U3039 (N_3039,In_1288,In_1280);
nor U3040 (N_3040,In_477,In_773);
xnor U3041 (N_3041,In_180,In_161);
and U3042 (N_3042,In_1475,In_787);
or U3043 (N_3043,In_1726,In_1021);
nor U3044 (N_3044,In_359,In_209);
nand U3045 (N_3045,In_123,In_423);
or U3046 (N_3046,In_941,In_861);
nor U3047 (N_3047,In_1182,In_1365);
or U3048 (N_3048,In_1575,In_621);
nor U3049 (N_3049,In_1754,In_256);
nor U3050 (N_3050,In_1439,In_1405);
nand U3051 (N_3051,In_692,In_79);
or U3052 (N_3052,In_686,In_1395);
nor U3053 (N_3053,In_312,In_889);
nor U3054 (N_3054,In_1954,In_103);
xor U3055 (N_3055,In_247,In_795);
nand U3056 (N_3056,In_1115,In_751);
or U3057 (N_3057,In_1698,In_1150);
nand U3058 (N_3058,In_1470,In_1167);
nand U3059 (N_3059,In_1257,In_647);
nor U3060 (N_3060,In_110,In_1428);
nor U3061 (N_3061,In_315,In_287);
and U3062 (N_3062,In_1894,In_966);
nor U3063 (N_3063,In_3,In_1458);
nor U3064 (N_3064,In_891,In_1667);
or U3065 (N_3065,In_1387,In_142);
xor U3066 (N_3066,In_751,In_1581);
nand U3067 (N_3067,In_649,In_1963);
or U3068 (N_3068,In_1,In_176);
xor U3069 (N_3069,In_922,In_904);
xnor U3070 (N_3070,In_332,In_897);
and U3071 (N_3071,In_281,In_390);
xnor U3072 (N_3072,In_1524,In_1001);
xnor U3073 (N_3073,In_979,In_454);
nor U3074 (N_3074,In_634,In_1654);
xnor U3075 (N_3075,In_1331,In_945);
nor U3076 (N_3076,In_1384,In_150);
or U3077 (N_3077,In_376,In_870);
and U3078 (N_3078,In_30,In_1500);
or U3079 (N_3079,In_914,In_954);
nand U3080 (N_3080,In_1583,In_1179);
nor U3081 (N_3081,In_119,In_727);
and U3082 (N_3082,In_549,In_49);
xor U3083 (N_3083,In_44,In_781);
nor U3084 (N_3084,In_1062,In_1733);
nand U3085 (N_3085,In_76,In_219);
xor U3086 (N_3086,In_593,In_1988);
nand U3087 (N_3087,In_422,In_1415);
or U3088 (N_3088,In_1478,In_964);
and U3089 (N_3089,In_1049,In_1604);
nand U3090 (N_3090,In_1645,In_1188);
and U3091 (N_3091,In_10,In_51);
or U3092 (N_3092,In_185,In_1089);
and U3093 (N_3093,In_1650,In_1564);
and U3094 (N_3094,In_141,In_1457);
or U3095 (N_3095,In_952,In_737);
and U3096 (N_3096,In_1848,In_1967);
and U3097 (N_3097,In_327,In_84);
and U3098 (N_3098,In_889,In_1766);
nand U3099 (N_3099,In_130,In_1443);
or U3100 (N_3100,In_1926,In_1975);
nand U3101 (N_3101,In_1887,In_410);
nand U3102 (N_3102,In_1781,In_1339);
nor U3103 (N_3103,In_1249,In_1769);
nand U3104 (N_3104,In_1536,In_763);
nand U3105 (N_3105,In_648,In_775);
or U3106 (N_3106,In_1558,In_223);
and U3107 (N_3107,In_1151,In_1537);
or U3108 (N_3108,In_744,In_1147);
nand U3109 (N_3109,In_1486,In_10);
or U3110 (N_3110,In_1804,In_303);
nand U3111 (N_3111,In_136,In_360);
or U3112 (N_3112,In_870,In_829);
nor U3113 (N_3113,In_1516,In_1824);
xnor U3114 (N_3114,In_483,In_1664);
and U3115 (N_3115,In_960,In_320);
or U3116 (N_3116,In_240,In_1426);
and U3117 (N_3117,In_1089,In_979);
xnor U3118 (N_3118,In_547,In_67);
xor U3119 (N_3119,In_371,In_1490);
nor U3120 (N_3120,In_45,In_1004);
nand U3121 (N_3121,In_362,In_264);
and U3122 (N_3122,In_825,In_1828);
nor U3123 (N_3123,In_448,In_1693);
nand U3124 (N_3124,In_685,In_1979);
nor U3125 (N_3125,In_389,In_783);
or U3126 (N_3126,In_255,In_1359);
and U3127 (N_3127,In_1727,In_1241);
xnor U3128 (N_3128,In_566,In_714);
and U3129 (N_3129,In_1375,In_1611);
or U3130 (N_3130,In_1373,In_791);
xor U3131 (N_3131,In_844,In_1428);
or U3132 (N_3132,In_1367,In_1921);
and U3133 (N_3133,In_1433,In_1984);
and U3134 (N_3134,In_25,In_804);
and U3135 (N_3135,In_500,In_1834);
nor U3136 (N_3136,In_552,In_1763);
nand U3137 (N_3137,In_712,In_1249);
nor U3138 (N_3138,In_479,In_787);
xor U3139 (N_3139,In_139,In_1209);
nand U3140 (N_3140,In_348,In_460);
xor U3141 (N_3141,In_930,In_277);
or U3142 (N_3142,In_1456,In_655);
or U3143 (N_3143,In_707,In_1448);
xor U3144 (N_3144,In_280,In_1285);
xnor U3145 (N_3145,In_953,In_1299);
xnor U3146 (N_3146,In_195,In_1323);
and U3147 (N_3147,In_1963,In_1581);
xnor U3148 (N_3148,In_924,In_357);
xnor U3149 (N_3149,In_1046,In_1739);
or U3150 (N_3150,In_1911,In_108);
xor U3151 (N_3151,In_1865,In_1907);
or U3152 (N_3152,In_29,In_1446);
xor U3153 (N_3153,In_1647,In_1877);
xor U3154 (N_3154,In_575,In_328);
nand U3155 (N_3155,In_196,In_1155);
and U3156 (N_3156,In_1162,In_645);
or U3157 (N_3157,In_1797,In_415);
and U3158 (N_3158,In_1692,In_1264);
nand U3159 (N_3159,In_892,In_831);
xor U3160 (N_3160,In_1705,In_71);
or U3161 (N_3161,In_149,In_1192);
and U3162 (N_3162,In_1169,In_1446);
and U3163 (N_3163,In_730,In_420);
xor U3164 (N_3164,In_787,In_73);
and U3165 (N_3165,In_950,In_594);
nand U3166 (N_3166,In_1280,In_632);
nor U3167 (N_3167,In_355,In_1511);
nand U3168 (N_3168,In_317,In_1557);
xor U3169 (N_3169,In_1171,In_1778);
xor U3170 (N_3170,In_1337,In_1454);
and U3171 (N_3171,In_1401,In_1819);
nor U3172 (N_3172,In_391,In_784);
or U3173 (N_3173,In_225,In_952);
nand U3174 (N_3174,In_612,In_1810);
and U3175 (N_3175,In_745,In_332);
xor U3176 (N_3176,In_654,In_1293);
xnor U3177 (N_3177,In_658,In_54);
xnor U3178 (N_3178,In_1221,In_191);
and U3179 (N_3179,In_936,In_1212);
xnor U3180 (N_3180,In_359,In_857);
and U3181 (N_3181,In_782,In_139);
and U3182 (N_3182,In_543,In_1932);
nor U3183 (N_3183,In_54,In_689);
nor U3184 (N_3184,In_1632,In_201);
nor U3185 (N_3185,In_824,In_1004);
and U3186 (N_3186,In_1529,In_1839);
nand U3187 (N_3187,In_29,In_464);
and U3188 (N_3188,In_721,In_117);
and U3189 (N_3189,In_776,In_1932);
or U3190 (N_3190,In_880,In_1835);
and U3191 (N_3191,In_1683,In_589);
nor U3192 (N_3192,In_883,In_1937);
and U3193 (N_3193,In_1275,In_1733);
nor U3194 (N_3194,In_1116,In_1197);
and U3195 (N_3195,In_801,In_479);
or U3196 (N_3196,In_447,In_1623);
or U3197 (N_3197,In_482,In_1999);
nor U3198 (N_3198,In_1176,In_1858);
nand U3199 (N_3199,In_869,In_43);
xor U3200 (N_3200,In_628,In_1739);
xnor U3201 (N_3201,In_1829,In_166);
and U3202 (N_3202,In_1715,In_330);
nand U3203 (N_3203,In_743,In_1011);
and U3204 (N_3204,In_422,In_1656);
or U3205 (N_3205,In_1199,In_1556);
and U3206 (N_3206,In_1179,In_934);
nand U3207 (N_3207,In_52,In_651);
nor U3208 (N_3208,In_895,In_1871);
or U3209 (N_3209,In_347,In_240);
and U3210 (N_3210,In_798,In_1572);
nor U3211 (N_3211,In_1121,In_1065);
nor U3212 (N_3212,In_1477,In_820);
xor U3213 (N_3213,In_919,In_338);
and U3214 (N_3214,In_201,In_189);
and U3215 (N_3215,In_594,In_1994);
and U3216 (N_3216,In_74,In_1363);
xor U3217 (N_3217,In_1970,In_581);
or U3218 (N_3218,In_832,In_1458);
nand U3219 (N_3219,In_1571,In_1244);
or U3220 (N_3220,In_1083,In_1880);
nor U3221 (N_3221,In_630,In_1250);
nand U3222 (N_3222,In_1895,In_1967);
xnor U3223 (N_3223,In_564,In_537);
nand U3224 (N_3224,In_305,In_1192);
and U3225 (N_3225,In_146,In_1179);
or U3226 (N_3226,In_1885,In_1456);
and U3227 (N_3227,In_1294,In_1461);
and U3228 (N_3228,In_1214,In_1630);
nand U3229 (N_3229,In_1210,In_905);
and U3230 (N_3230,In_512,In_748);
and U3231 (N_3231,In_54,In_1053);
xnor U3232 (N_3232,In_933,In_1229);
nor U3233 (N_3233,In_1147,In_640);
xor U3234 (N_3234,In_532,In_1771);
and U3235 (N_3235,In_1252,In_530);
xnor U3236 (N_3236,In_1901,In_1344);
nor U3237 (N_3237,In_1170,In_92);
and U3238 (N_3238,In_608,In_255);
or U3239 (N_3239,In_1858,In_787);
and U3240 (N_3240,In_883,In_1385);
nand U3241 (N_3241,In_993,In_280);
and U3242 (N_3242,In_270,In_1491);
or U3243 (N_3243,In_1220,In_1211);
nand U3244 (N_3244,In_1578,In_623);
nand U3245 (N_3245,In_724,In_223);
or U3246 (N_3246,In_1641,In_839);
nor U3247 (N_3247,In_1703,In_906);
and U3248 (N_3248,In_841,In_211);
nand U3249 (N_3249,In_1431,In_736);
xnor U3250 (N_3250,In_611,In_408);
nor U3251 (N_3251,In_325,In_1075);
and U3252 (N_3252,In_742,In_1597);
or U3253 (N_3253,In_1215,In_1593);
xor U3254 (N_3254,In_707,In_1877);
nand U3255 (N_3255,In_1056,In_335);
nor U3256 (N_3256,In_588,In_1366);
xor U3257 (N_3257,In_439,In_1875);
and U3258 (N_3258,In_1694,In_659);
xnor U3259 (N_3259,In_173,In_1215);
and U3260 (N_3260,In_1213,In_1307);
xnor U3261 (N_3261,In_8,In_1743);
or U3262 (N_3262,In_448,In_149);
xnor U3263 (N_3263,In_1381,In_728);
nand U3264 (N_3264,In_929,In_372);
xor U3265 (N_3265,In_1546,In_45);
nor U3266 (N_3266,In_85,In_1877);
nand U3267 (N_3267,In_882,In_1759);
and U3268 (N_3268,In_1959,In_1302);
nand U3269 (N_3269,In_795,In_161);
xnor U3270 (N_3270,In_1337,In_445);
xnor U3271 (N_3271,In_721,In_1216);
nand U3272 (N_3272,In_187,In_327);
nand U3273 (N_3273,In_448,In_35);
nor U3274 (N_3274,In_360,In_1247);
nand U3275 (N_3275,In_638,In_1166);
and U3276 (N_3276,In_954,In_750);
nand U3277 (N_3277,In_1500,In_673);
nand U3278 (N_3278,In_361,In_1343);
and U3279 (N_3279,In_1991,In_421);
nand U3280 (N_3280,In_1918,In_1333);
or U3281 (N_3281,In_1316,In_410);
xor U3282 (N_3282,In_1433,In_254);
and U3283 (N_3283,In_1250,In_1614);
xnor U3284 (N_3284,In_647,In_318);
and U3285 (N_3285,In_1199,In_254);
nor U3286 (N_3286,In_571,In_884);
or U3287 (N_3287,In_328,In_1993);
xnor U3288 (N_3288,In_819,In_1998);
or U3289 (N_3289,In_661,In_850);
xor U3290 (N_3290,In_1957,In_407);
xor U3291 (N_3291,In_376,In_1686);
nor U3292 (N_3292,In_214,In_1017);
and U3293 (N_3293,In_106,In_379);
and U3294 (N_3294,In_421,In_1466);
nand U3295 (N_3295,In_1749,In_329);
or U3296 (N_3296,In_476,In_741);
nor U3297 (N_3297,In_165,In_1285);
and U3298 (N_3298,In_631,In_677);
nand U3299 (N_3299,In_332,In_1163);
xor U3300 (N_3300,In_1890,In_760);
nor U3301 (N_3301,In_1492,In_1129);
and U3302 (N_3302,In_911,In_1584);
xnor U3303 (N_3303,In_951,In_1491);
nor U3304 (N_3304,In_1912,In_1022);
nor U3305 (N_3305,In_450,In_979);
nor U3306 (N_3306,In_605,In_570);
or U3307 (N_3307,In_1138,In_44);
or U3308 (N_3308,In_1651,In_153);
nand U3309 (N_3309,In_1920,In_1275);
nor U3310 (N_3310,In_1650,In_378);
nor U3311 (N_3311,In_607,In_1391);
nand U3312 (N_3312,In_1555,In_1162);
nor U3313 (N_3313,In_527,In_809);
or U3314 (N_3314,In_1708,In_1080);
nand U3315 (N_3315,In_339,In_1028);
or U3316 (N_3316,In_239,In_831);
nand U3317 (N_3317,In_56,In_546);
or U3318 (N_3318,In_315,In_1934);
nand U3319 (N_3319,In_875,In_1677);
xnor U3320 (N_3320,In_774,In_631);
nor U3321 (N_3321,In_1714,In_699);
and U3322 (N_3322,In_1761,In_110);
nor U3323 (N_3323,In_1443,In_1585);
nor U3324 (N_3324,In_1840,In_1819);
nor U3325 (N_3325,In_1691,In_1386);
nand U3326 (N_3326,In_1310,In_1481);
nor U3327 (N_3327,In_1814,In_1725);
nand U3328 (N_3328,In_1101,In_523);
nand U3329 (N_3329,In_1942,In_1691);
nand U3330 (N_3330,In_176,In_568);
xor U3331 (N_3331,In_1676,In_1976);
nor U3332 (N_3332,In_119,In_1365);
and U3333 (N_3333,In_824,In_267);
or U3334 (N_3334,In_1428,In_1042);
nand U3335 (N_3335,In_1600,In_90);
nand U3336 (N_3336,In_25,In_1699);
nor U3337 (N_3337,In_1860,In_144);
nand U3338 (N_3338,In_1678,In_1487);
nor U3339 (N_3339,In_1004,In_1146);
or U3340 (N_3340,In_952,In_1424);
nor U3341 (N_3341,In_669,In_1659);
or U3342 (N_3342,In_408,In_651);
xor U3343 (N_3343,In_1246,In_1388);
or U3344 (N_3344,In_442,In_1704);
or U3345 (N_3345,In_861,In_398);
nand U3346 (N_3346,In_181,In_1958);
or U3347 (N_3347,In_1994,In_1781);
and U3348 (N_3348,In_178,In_1408);
nand U3349 (N_3349,In_1381,In_525);
nand U3350 (N_3350,In_1528,In_276);
or U3351 (N_3351,In_1459,In_1072);
and U3352 (N_3352,In_275,In_222);
nor U3353 (N_3353,In_28,In_379);
xor U3354 (N_3354,In_374,In_724);
xor U3355 (N_3355,In_1820,In_546);
or U3356 (N_3356,In_537,In_71);
or U3357 (N_3357,In_389,In_344);
and U3358 (N_3358,In_27,In_1722);
xor U3359 (N_3359,In_1896,In_256);
or U3360 (N_3360,In_1186,In_1993);
nand U3361 (N_3361,In_1776,In_1035);
nand U3362 (N_3362,In_272,In_1436);
nor U3363 (N_3363,In_1745,In_1801);
nand U3364 (N_3364,In_1003,In_599);
nand U3365 (N_3365,In_716,In_93);
or U3366 (N_3366,In_1512,In_968);
nor U3367 (N_3367,In_516,In_541);
nand U3368 (N_3368,In_412,In_127);
nand U3369 (N_3369,In_252,In_85);
or U3370 (N_3370,In_1331,In_1483);
or U3371 (N_3371,In_1679,In_549);
xor U3372 (N_3372,In_521,In_49);
nand U3373 (N_3373,In_108,In_1898);
nand U3374 (N_3374,In_357,In_1568);
nor U3375 (N_3375,In_1170,In_46);
and U3376 (N_3376,In_1372,In_529);
xnor U3377 (N_3377,In_513,In_1243);
xnor U3378 (N_3378,In_1003,In_402);
nor U3379 (N_3379,In_1191,In_1017);
nand U3380 (N_3380,In_61,In_1482);
and U3381 (N_3381,In_1107,In_240);
xnor U3382 (N_3382,In_1056,In_860);
or U3383 (N_3383,In_297,In_477);
and U3384 (N_3384,In_1772,In_1234);
nor U3385 (N_3385,In_1236,In_1724);
xnor U3386 (N_3386,In_997,In_1815);
nand U3387 (N_3387,In_1677,In_409);
and U3388 (N_3388,In_621,In_1064);
and U3389 (N_3389,In_302,In_1525);
xnor U3390 (N_3390,In_914,In_1811);
or U3391 (N_3391,In_607,In_385);
nand U3392 (N_3392,In_1112,In_1185);
and U3393 (N_3393,In_1529,In_1939);
and U3394 (N_3394,In_1380,In_340);
and U3395 (N_3395,In_1501,In_1478);
nor U3396 (N_3396,In_1291,In_1236);
nand U3397 (N_3397,In_1753,In_123);
nand U3398 (N_3398,In_131,In_479);
or U3399 (N_3399,In_1423,In_1962);
or U3400 (N_3400,In_1616,In_1934);
nand U3401 (N_3401,In_915,In_1716);
or U3402 (N_3402,In_693,In_199);
and U3403 (N_3403,In_1971,In_1437);
xnor U3404 (N_3404,In_1475,In_370);
nor U3405 (N_3405,In_983,In_1703);
xnor U3406 (N_3406,In_1437,In_1528);
nand U3407 (N_3407,In_1672,In_1928);
nor U3408 (N_3408,In_1596,In_1245);
nand U3409 (N_3409,In_1388,In_1364);
and U3410 (N_3410,In_1566,In_1575);
nor U3411 (N_3411,In_84,In_48);
nand U3412 (N_3412,In_1937,In_336);
xor U3413 (N_3413,In_1010,In_969);
xor U3414 (N_3414,In_856,In_977);
and U3415 (N_3415,In_1,In_326);
nand U3416 (N_3416,In_1319,In_750);
nor U3417 (N_3417,In_1732,In_476);
nor U3418 (N_3418,In_1901,In_805);
nor U3419 (N_3419,In_511,In_1023);
xor U3420 (N_3420,In_1450,In_1027);
nand U3421 (N_3421,In_604,In_1669);
xor U3422 (N_3422,In_958,In_378);
nand U3423 (N_3423,In_603,In_1882);
or U3424 (N_3424,In_1183,In_1171);
or U3425 (N_3425,In_862,In_1317);
nand U3426 (N_3426,In_1795,In_396);
and U3427 (N_3427,In_977,In_883);
nand U3428 (N_3428,In_290,In_1749);
and U3429 (N_3429,In_754,In_1835);
xor U3430 (N_3430,In_451,In_87);
or U3431 (N_3431,In_291,In_260);
or U3432 (N_3432,In_127,In_1615);
or U3433 (N_3433,In_1848,In_1643);
xor U3434 (N_3434,In_1468,In_1184);
nand U3435 (N_3435,In_756,In_519);
nor U3436 (N_3436,In_1911,In_976);
nor U3437 (N_3437,In_1346,In_1396);
or U3438 (N_3438,In_1089,In_1768);
and U3439 (N_3439,In_1028,In_1252);
or U3440 (N_3440,In_1647,In_229);
or U3441 (N_3441,In_1494,In_1146);
nand U3442 (N_3442,In_318,In_1074);
xnor U3443 (N_3443,In_1411,In_91);
nand U3444 (N_3444,In_1310,In_698);
nor U3445 (N_3445,In_1116,In_1799);
xnor U3446 (N_3446,In_848,In_959);
or U3447 (N_3447,In_836,In_1146);
nor U3448 (N_3448,In_1472,In_242);
xnor U3449 (N_3449,In_264,In_1580);
nand U3450 (N_3450,In_1802,In_158);
and U3451 (N_3451,In_953,In_1554);
xor U3452 (N_3452,In_162,In_1521);
and U3453 (N_3453,In_1064,In_1339);
and U3454 (N_3454,In_1611,In_777);
nor U3455 (N_3455,In_943,In_1580);
and U3456 (N_3456,In_1524,In_839);
and U3457 (N_3457,In_1557,In_138);
or U3458 (N_3458,In_1499,In_258);
or U3459 (N_3459,In_331,In_1030);
xor U3460 (N_3460,In_1875,In_1072);
xnor U3461 (N_3461,In_1358,In_1872);
nand U3462 (N_3462,In_1921,In_778);
nand U3463 (N_3463,In_1062,In_528);
or U3464 (N_3464,In_151,In_980);
and U3465 (N_3465,In_1918,In_54);
or U3466 (N_3466,In_1782,In_1241);
nand U3467 (N_3467,In_1820,In_1076);
nor U3468 (N_3468,In_1661,In_815);
nand U3469 (N_3469,In_157,In_788);
nor U3470 (N_3470,In_1182,In_116);
nand U3471 (N_3471,In_1563,In_1009);
nand U3472 (N_3472,In_630,In_174);
and U3473 (N_3473,In_402,In_118);
and U3474 (N_3474,In_193,In_1127);
and U3475 (N_3475,In_467,In_523);
xnor U3476 (N_3476,In_889,In_130);
xnor U3477 (N_3477,In_1773,In_1897);
nand U3478 (N_3478,In_721,In_9);
nand U3479 (N_3479,In_158,In_207);
or U3480 (N_3480,In_1021,In_1447);
nand U3481 (N_3481,In_1070,In_1760);
nand U3482 (N_3482,In_678,In_1260);
nor U3483 (N_3483,In_631,In_996);
and U3484 (N_3484,In_1345,In_594);
or U3485 (N_3485,In_1875,In_333);
nor U3486 (N_3486,In_1052,In_1172);
nor U3487 (N_3487,In_224,In_1498);
xor U3488 (N_3488,In_1911,In_252);
xnor U3489 (N_3489,In_1253,In_1881);
and U3490 (N_3490,In_281,In_540);
nand U3491 (N_3491,In_1632,In_1917);
and U3492 (N_3492,In_269,In_549);
or U3493 (N_3493,In_1885,In_1624);
nor U3494 (N_3494,In_1940,In_1261);
and U3495 (N_3495,In_235,In_1765);
nor U3496 (N_3496,In_1857,In_1165);
nand U3497 (N_3497,In_1387,In_1832);
or U3498 (N_3498,In_1007,In_1384);
nor U3499 (N_3499,In_1723,In_1829);
nor U3500 (N_3500,In_1622,In_1611);
or U3501 (N_3501,In_1311,In_377);
nor U3502 (N_3502,In_451,In_1378);
xnor U3503 (N_3503,In_816,In_425);
and U3504 (N_3504,In_1296,In_367);
nand U3505 (N_3505,In_721,In_1944);
and U3506 (N_3506,In_1873,In_1896);
nand U3507 (N_3507,In_796,In_1402);
nand U3508 (N_3508,In_1851,In_443);
nor U3509 (N_3509,In_886,In_1684);
nand U3510 (N_3510,In_347,In_760);
nor U3511 (N_3511,In_1815,In_154);
nor U3512 (N_3512,In_525,In_573);
nand U3513 (N_3513,In_854,In_1598);
nand U3514 (N_3514,In_159,In_1768);
nand U3515 (N_3515,In_568,In_562);
and U3516 (N_3516,In_1084,In_612);
nand U3517 (N_3517,In_50,In_1512);
nor U3518 (N_3518,In_1922,In_954);
xor U3519 (N_3519,In_227,In_1266);
xnor U3520 (N_3520,In_996,In_1799);
nor U3521 (N_3521,In_1269,In_1042);
xnor U3522 (N_3522,In_1856,In_709);
nor U3523 (N_3523,In_189,In_1480);
xor U3524 (N_3524,In_135,In_1410);
xor U3525 (N_3525,In_190,In_1069);
and U3526 (N_3526,In_1601,In_320);
and U3527 (N_3527,In_1691,In_1141);
xnor U3528 (N_3528,In_214,In_1839);
nand U3529 (N_3529,In_1345,In_1778);
xnor U3530 (N_3530,In_850,In_1647);
nand U3531 (N_3531,In_600,In_1708);
xor U3532 (N_3532,In_36,In_309);
xor U3533 (N_3533,In_601,In_681);
or U3534 (N_3534,In_1900,In_868);
nor U3535 (N_3535,In_1338,In_0);
or U3536 (N_3536,In_1560,In_1705);
nand U3537 (N_3537,In_786,In_1213);
nor U3538 (N_3538,In_437,In_1478);
nand U3539 (N_3539,In_1117,In_266);
xnor U3540 (N_3540,In_49,In_1001);
nand U3541 (N_3541,In_1493,In_1439);
nand U3542 (N_3542,In_485,In_1031);
xor U3543 (N_3543,In_1261,In_1370);
or U3544 (N_3544,In_1360,In_973);
nor U3545 (N_3545,In_449,In_1664);
nor U3546 (N_3546,In_787,In_700);
nor U3547 (N_3547,In_1186,In_235);
or U3548 (N_3548,In_1851,In_148);
xnor U3549 (N_3549,In_826,In_778);
or U3550 (N_3550,In_745,In_1044);
or U3551 (N_3551,In_215,In_315);
nor U3552 (N_3552,In_1760,In_562);
or U3553 (N_3553,In_1153,In_1548);
nand U3554 (N_3554,In_1154,In_866);
or U3555 (N_3555,In_348,In_1668);
xor U3556 (N_3556,In_1193,In_1918);
nand U3557 (N_3557,In_1421,In_152);
and U3558 (N_3558,In_159,In_1973);
xnor U3559 (N_3559,In_1974,In_308);
xnor U3560 (N_3560,In_130,In_1626);
nand U3561 (N_3561,In_431,In_930);
nand U3562 (N_3562,In_1264,In_1599);
xnor U3563 (N_3563,In_888,In_755);
or U3564 (N_3564,In_555,In_733);
and U3565 (N_3565,In_1165,In_1463);
and U3566 (N_3566,In_1749,In_180);
xnor U3567 (N_3567,In_574,In_1163);
xnor U3568 (N_3568,In_1271,In_1306);
nand U3569 (N_3569,In_750,In_1509);
and U3570 (N_3570,In_302,In_1603);
or U3571 (N_3571,In_565,In_1460);
or U3572 (N_3572,In_1667,In_1700);
nor U3573 (N_3573,In_1163,In_685);
or U3574 (N_3574,In_1216,In_1979);
and U3575 (N_3575,In_1352,In_659);
nor U3576 (N_3576,In_1828,In_848);
nand U3577 (N_3577,In_57,In_1240);
nand U3578 (N_3578,In_1986,In_803);
and U3579 (N_3579,In_1550,In_813);
nand U3580 (N_3580,In_201,In_87);
or U3581 (N_3581,In_1908,In_1691);
or U3582 (N_3582,In_933,In_314);
xor U3583 (N_3583,In_1842,In_938);
or U3584 (N_3584,In_1624,In_659);
xor U3585 (N_3585,In_755,In_1870);
nor U3586 (N_3586,In_158,In_993);
nor U3587 (N_3587,In_1199,In_1049);
nor U3588 (N_3588,In_1403,In_750);
and U3589 (N_3589,In_1949,In_757);
nand U3590 (N_3590,In_911,In_749);
and U3591 (N_3591,In_676,In_1705);
and U3592 (N_3592,In_1094,In_1671);
or U3593 (N_3593,In_1496,In_1308);
and U3594 (N_3594,In_332,In_1952);
nor U3595 (N_3595,In_909,In_739);
nor U3596 (N_3596,In_1855,In_1446);
and U3597 (N_3597,In_1224,In_659);
xor U3598 (N_3598,In_1408,In_1635);
nand U3599 (N_3599,In_290,In_996);
xor U3600 (N_3600,In_1166,In_1659);
or U3601 (N_3601,In_924,In_1468);
and U3602 (N_3602,In_1179,In_1586);
xnor U3603 (N_3603,In_1190,In_1280);
nor U3604 (N_3604,In_519,In_1961);
or U3605 (N_3605,In_438,In_1016);
xnor U3606 (N_3606,In_1615,In_285);
nor U3607 (N_3607,In_411,In_386);
nor U3608 (N_3608,In_757,In_1724);
nor U3609 (N_3609,In_1236,In_1562);
nand U3610 (N_3610,In_107,In_1803);
xor U3611 (N_3611,In_1751,In_357);
and U3612 (N_3612,In_1241,In_375);
nor U3613 (N_3613,In_454,In_596);
and U3614 (N_3614,In_1502,In_1602);
nor U3615 (N_3615,In_835,In_1293);
nor U3616 (N_3616,In_1027,In_672);
xnor U3617 (N_3617,In_930,In_1217);
xnor U3618 (N_3618,In_862,In_1670);
and U3619 (N_3619,In_92,In_51);
xor U3620 (N_3620,In_770,In_1402);
and U3621 (N_3621,In_964,In_91);
and U3622 (N_3622,In_465,In_126);
and U3623 (N_3623,In_1211,In_1199);
and U3624 (N_3624,In_1078,In_1518);
or U3625 (N_3625,In_590,In_1698);
and U3626 (N_3626,In_804,In_781);
nor U3627 (N_3627,In_867,In_370);
xnor U3628 (N_3628,In_1905,In_955);
nand U3629 (N_3629,In_835,In_1021);
and U3630 (N_3630,In_827,In_1530);
and U3631 (N_3631,In_840,In_97);
xor U3632 (N_3632,In_1091,In_55);
or U3633 (N_3633,In_1551,In_1547);
nand U3634 (N_3634,In_105,In_620);
xnor U3635 (N_3635,In_664,In_1842);
nand U3636 (N_3636,In_1850,In_61);
or U3637 (N_3637,In_326,In_1517);
or U3638 (N_3638,In_404,In_565);
nand U3639 (N_3639,In_541,In_953);
or U3640 (N_3640,In_10,In_490);
nor U3641 (N_3641,In_597,In_724);
nor U3642 (N_3642,In_307,In_1656);
xnor U3643 (N_3643,In_7,In_1091);
xnor U3644 (N_3644,In_1915,In_1405);
nand U3645 (N_3645,In_1345,In_207);
nor U3646 (N_3646,In_1568,In_1123);
nand U3647 (N_3647,In_1509,In_616);
nor U3648 (N_3648,In_1622,In_267);
or U3649 (N_3649,In_1759,In_609);
nor U3650 (N_3650,In_1466,In_1610);
nor U3651 (N_3651,In_655,In_601);
nor U3652 (N_3652,In_1596,In_631);
or U3653 (N_3653,In_1343,In_1949);
xor U3654 (N_3654,In_1307,In_1158);
xor U3655 (N_3655,In_1939,In_531);
nor U3656 (N_3656,In_731,In_474);
xor U3657 (N_3657,In_15,In_562);
or U3658 (N_3658,In_656,In_729);
nand U3659 (N_3659,In_1517,In_1416);
xor U3660 (N_3660,In_1383,In_832);
xnor U3661 (N_3661,In_1074,In_1914);
nand U3662 (N_3662,In_1095,In_394);
nand U3663 (N_3663,In_18,In_1643);
xnor U3664 (N_3664,In_1486,In_225);
xnor U3665 (N_3665,In_1311,In_37);
nor U3666 (N_3666,In_1281,In_1380);
and U3667 (N_3667,In_1293,In_20);
nor U3668 (N_3668,In_1218,In_1961);
xnor U3669 (N_3669,In_1087,In_953);
or U3670 (N_3670,In_615,In_216);
or U3671 (N_3671,In_1146,In_686);
nand U3672 (N_3672,In_701,In_619);
xor U3673 (N_3673,In_1781,In_1309);
and U3674 (N_3674,In_1166,In_54);
xor U3675 (N_3675,In_1899,In_1016);
nand U3676 (N_3676,In_25,In_140);
xor U3677 (N_3677,In_107,In_1814);
or U3678 (N_3678,In_913,In_1672);
nor U3679 (N_3679,In_1195,In_33);
or U3680 (N_3680,In_1099,In_1850);
nor U3681 (N_3681,In_1852,In_171);
xor U3682 (N_3682,In_727,In_774);
xnor U3683 (N_3683,In_160,In_19);
or U3684 (N_3684,In_303,In_156);
or U3685 (N_3685,In_1033,In_899);
xnor U3686 (N_3686,In_385,In_1058);
or U3687 (N_3687,In_247,In_1097);
nor U3688 (N_3688,In_1778,In_158);
xnor U3689 (N_3689,In_1295,In_1788);
and U3690 (N_3690,In_893,In_797);
nor U3691 (N_3691,In_1733,In_709);
nand U3692 (N_3692,In_1603,In_1832);
and U3693 (N_3693,In_1128,In_1977);
or U3694 (N_3694,In_963,In_1276);
and U3695 (N_3695,In_1113,In_1717);
or U3696 (N_3696,In_247,In_471);
xor U3697 (N_3697,In_909,In_251);
and U3698 (N_3698,In_806,In_169);
or U3699 (N_3699,In_377,In_857);
or U3700 (N_3700,In_1266,In_694);
or U3701 (N_3701,In_1692,In_260);
nand U3702 (N_3702,In_1195,In_1921);
nor U3703 (N_3703,In_808,In_368);
xnor U3704 (N_3704,In_982,In_1740);
nor U3705 (N_3705,In_1548,In_1034);
xor U3706 (N_3706,In_1152,In_785);
nand U3707 (N_3707,In_1460,In_411);
nor U3708 (N_3708,In_1527,In_1724);
nor U3709 (N_3709,In_560,In_1889);
or U3710 (N_3710,In_1839,In_32);
nor U3711 (N_3711,In_463,In_1767);
xnor U3712 (N_3712,In_508,In_92);
nand U3713 (N_3713,In_931,In_1973);
and U3714 (N_3714,In_391,In_633);
nand U3715 (N_3715,In_261,In_1649);
nor U3716 (N_3716,In_1042,In_267);
nor U3717 (N_3717,In_389,In_317);
or U3718 (N_3718,In_32,In_103);
nand U3719 (N_3719,In_996,In_1167);
and U3720 (N_3720,In_586,In_1096);
xor U3721 (N_3721,In_39,In_325);
or U3722 (N_3722,In_737,In_1136);
xor U3723 (N_3723,In_12,In_1512);
and U3724 (N_3724,In_93,In_1296);
nand U3725 (N_3725,In_412,In_1137);
or U3726 (N_3726,In_50,In_172);
xor U3727 (N_3727,In_1418,In_1136);
or U3728 (N_3728,In_50,In_395);
nand U3729 (N_3729,In_1194,In_846);
xnor U3730 (N_3730,In_1353,In_1757);
nand U3731 (N_3731,In_1943,In_1907);
or U3732 (N_3732,In_1536,In_1482);
and U3733 (N_3733,In_628,In_1744);
and U3734 (N_3734,In_1190,In_1163);
and U3735 (N_3735,In_533,In_315);
nand U3736 (N_3736,In_437,In_267);
nand U3737 (N_3737,In_1577,In_1990);
and U3738 (N_3738,In_899,In_1953);
xor U3739 (N_3739,In_719,In_251);
xor U3740 (N_3740,In_1797,In_633);
and U3741 (N_3741,In_774,In_1583);
or U3742 (N_3742,In_1688,In_1262);
nand U3743 (N_3743,In_1130,In_1406);
and U3744 (N_3744,In_1401,In_1039);
or U3745 (N_3745,In_1059,In_973);
xor U3746 (N_3746,In_847,In_1507);
nand U3747 (N_3747,In_1139,In_1734);
nand U3748 (N_3748,In_1165,In_145);
xnor U3749 (N_3749,In_1229,In_1112);
or U3750 (N_3750,In_712,In_1796);
nand U3751 (N_3751,In_985,In_1379);
xnor U3752 (N_3752,In_1586,In_660);
and U3753 (N_3753,In_1060,In_469);
nand U3754 (N_3754,In_1433,In_1730);
or U3755 (N_3755,In_399,In_233);
xnor U3756 (N_3756,In_886,In_66);
xnor U3757 (N_3757,In_1127,In_1209);
nor U3758 (N_3758,In_235,In_355);
nand U3759 (N_3759,In_842,In_1795);
nand U3760 (N_3760,In_794,In_28);
nand U3761 (N_3761,In_969,In_1236);
xnor U3762 (N_3762,In_1189,In_707);
nand U3763 (N_3763,In_463,In_116);
or U3764 (N_3764,In_297,In_1418);
and U3765 (N_3765,In_908,In_902);
and U3766 (N_3766,In_1060,In_1686);
nor U3767 (N_3767,In_1984,In_940);
or U3768 (N_3768,In_660,In_948);
or U3769 (N_3769,In_1532,In_133);
xor U3770 (N_3770,In_25,In_1246);
and U3771 (N_3771,In_427,In_1309);
nor U3772 (N_3772,In_778,In_999);
nor U3773 (N_3773,In_672,In_491);
and U3774 (N_3774,In_1211,In_1975);
nand U3775 (N_3775,In_857,In_1229);
nor U3776 (N_3776,In_1954,In_202);
xnor U3777 (N_3777,In_10,In_224);
and U3778 (N_3778,In_751,In_701);
nand U3779 (N_3779,In_1115,In_1566);
and U3780 (N_3780,In_1768,In_1593);
xnor U3781 (N_3781,In_646,In_1885);
or U3782 (N_3782,In_987,In_766);
nor U3783 (N_3783,In_1957,In_1898);
and U3784 (N_3784,In_1531,In_514);
nor U3785 (N_3785,In_884,In_359);
nand U3786 (N_3786,In_409,In_7);
and U3787 (N_3787,In_382,In_1009);
or U3788 (N_3788,In_117,In_756);
nor U3789 (N_3789,In_894,In_85);
or U3790 (N_3790,In_1618,In_627);
or U3791 (N_3791,In_1180,In_296);
nor U3792 (N_3792,In_784,In_383);
or U3793 (N_3793,In_937,In_1415);
nand U3794 (N_3794,In_1194,In_1998);
nor U3795 (N_3795,In_807,In_120);
or U3796 (N_3796,In_1500,In_1668);
and U3797 (N_3797,In_1645,In_1199);
nand U3798 (N_3798,In_1443,In_1584);
xor U3799 (N_3799,In_181,In_1637);
and U3800 (N_3800,In_441,In_393);
xnor U3801 (N_3801,In_85,In_499);
and U3802 (N_3802,In_146,In_1590);
xnor U3803 (N_3803,In_1741,In_1596);
nand U3804 (N_3804,In_1135,In_1751);
or U3805 (N_3805,In_1656,In_1814);
or U3806 (N_3806,In_686,In_1920);
nand U3807 (N_3807,In_1499,In_1582);
and U3808 (N_3808,In_1840,In_821);
xor U3809 (N_3809,In_748,In_1074);
or U3810 (N_3810,In_283,In_106);
nor U3811 (N_3811,In_650,In_1819);
nand U3812 (N_3812,In_1319,In_1076);
nor U3813 (N_3813,In_1537,In_1772);
or U3814 (N_3814,In_667,In_653);
nand U3815 (N_3815,In_37,In_650);
xnor U3816 (N_3816,In_230,In_247);
and U3817 (N_3817,In_1438,In_1476);
xnor U3818 (N_3818,In_316,In_1608);
nand U3819 (N_3819,In_1231,In_1793);
nand U3820 (N_3820,In_338,In_1884);
xor U3821 (N_3821,In_1000,In_1531);
nand U3822 (N_3822,In_1515,In_1310);
and U3823 (N_3823,In_93,In_1021);
and U3824 (N_3824,In_980,In_1494);
and U3825 (N_3825,In_1971,In_1826);
and U3826 (N_3826,In_137,In_658);
nand U3827 (N_3827,In_66,In_1865);
and U3828 (N_3828,In_1824,In_194);
xor U3829 (N_3829,In_575,In_1882);
xor U3830 (N_3830,In_1420,In_1178);
nor U3831 (N_3831,In_828,In_1667);
or U3832 (N_3832,In_586,In_236);
or U3833 (N_3833,In_590,In_58);
or U3834 (N_3834,In_1837,In_283);
and U3835 (N_3835,In_353,In_1157);
nor U3836 (N_3836,In_571,In_961);
nor U3837 (N_3837,In_1574,In_610);
nand U3838 (N_3838,In_952,In_190);
nor U3839 (N_3839,In_916,In_469);
xnor U3840 (N_3840,In_1821,In_1713);
xnor U3841 (N_3841,In_66,In_1466);
nor U3842 (N_3842,In_942,In_1424);
nand U3843 (N_3843,In_652,In_257);
xnor U3844 (N_3844,In_434,In_383);
nand U3845 (N_3845,In_1224,In_709);
or U3846 (N_3846,In_150,In_1711);
nor U3847 (N_3847,In_541,In_131);
and U3848 (N_3848,In_941,In_1412);
nor U3849 (N_3849,In_672,In_629);
or U3850 (N_3850,In_1597,In_686);
nor U3851 (N_3851,In_1472,In_26);
nand U3852 (N_3852,In_1799,In_127);
nor U3853 (N_3853,In_1093,In_1336);
or U3854 (N_3854,In_1378,In_737);
and U3855 (N_3855,In_154,In_1926);
nor U3856 (N_3856,In_709,In_1674);
or U3857 (N_3857,In_1844,In_1545);
or U3858 (N_3858,In_79,In_1912);
xor U3859 (N_3859,In_1920,In_858);
xor U3860 (N_3860,In_618,In_1519);
or U3861 (N_3861,In_1876,In_338);
and U3862 (N_3862,In_1006,In_954);
nor U3863 (N_3863,In_1296,In_849);
and U3864 (N_3864,In_1768,In_1431);
nor U3865 (N_3865,In_1124,In_1139);
xnor U3866 (N_3866,In_9,In_1509);
or U3867 (N_3867,In_1089,In_1);
nand U3868 (N_3868,In_1328,In_364);
and U3869 (N_3869,In_1998,In_73);
nor U3870 (N_3870,In_1947,In_1939);
nand U3871 (N_3871,In_1949,In_1193);
nand U3872 (N_3872,In_649,In_215);
nand U3873 (N_3873,In_595,In_1064);
nand U3874 (N_3874,In_1682,In_1357);
xor U3875 (N_3875,In_486,In_1404);
or U3876 (N_3876,In_894,In_1967);
xor U3877 (N_3877,In_1629,In_1988);
xnor U3878 (N_3878,In_1030,In_732);
nand U3879 (N_3879,In_387,In_445);
nand U3880 (N_3880,In_1819,In_544);
nand U3881 (N_3881,In_1404,In_1389);
and U3882 (N_3882,In_871,In_1735);
and U3883 (N_3883,In_14,In_582);
xor U3884 (N_3884,In_920,In_1031);
nor U3885 (N_3885,In_936,In_1614);
nand U3886 (N_3886,In_411,In_192);
xor U3887 (N_3887,In_988,In_1135);
and U3888 (N_3888,In_549,In_177);
and U3889 (N_3889,In_1040,In_1811);
or U3890 (N_3890,In_435,In_1504);
nor U3891 (N_3891,In_177,In_1993);
nand U3892 (N_3892,In_244,In_800);
and U3893 (N_3893,In_411,In_1944);
nand U3894 (N_3894,In_623,In_875);
or U3895 (N_3895,In_1015,In_885);
nand U3896 (N_3896,In_180,In_1058);
nand U3897 (N_3897,In_1205,In_1621);
nand U3898 (N_3898,In_882,In_1040);
and U3899 (N_3899,In_1007,In_859);
or U3900 (N_3900,In_488,In_636);
or U3901 (N_3901,In_1776,In_371);
or U3902 (N_3902,In_1321,In_1386);
or U3903 (N_3903,In_1527,In_1024);
nand U3904 (N_3904,In_1548,In_89);
nand U3905 (N_3905,In_1467,In_262);
nand U3906 (N_3906,In_588,In_1101);
and U3907 (N_3907,In_1875,In_611);
and U3908 (N_3908,In_1702,In_548);
or U3909 (N_3909,In_1992,In_1374);
or U3910 (N_3910,In_596,In_377);
nor U3911 (N_3911,In_1277,In_393);
or U3912 (N_3912,In_1705,In_991);
and U3913 (N_3913,In_1260,In_1177);
nand U3914 (N_3914,In_1494,In_176);
or U3915 (N_3915,In_683,In_988);
nor U3916 (N_3916,In_1732,In_325);
nand U3917 (N_3917,In_1989,In_236);
nor U3918 (N_3918,In_980,In_1760);
nand U3919 (N_3919,In_420,In_1211);
nand U3920 (N_3920,In_881,In_811);
or U3921 (N_3921,In_1810,In_929);
nand U3922 (N_3922,In_106,In_1486);
xnor U3923 (N_3923,In_1469,In_1806);
nand U3924 (N_3924,In_1883,In_4);
nor U3925 (N_3925,In_760,In_352);
xor U3926 (N_3926,In_1011,In_551);
and U3927 (N_3927,In_888,In_357);
or U3928 (N_3928,In_1067,In_1142);
and U3929 (N_3929,In_1051,In_1539);
or U3930 (N_3930,In_1442,In_1850);
nand U3931 (N_3931,In_419,In_1181);
and U3932 (N_3932,In_1060,In_602);
nand U3933 (N_3933,In_945,In_1837);
nand U3934 (N_3934,In_399,In_1199);
nand U3935 (N_3935,In_252,In_1119);
or U3936 (N_3936,In_1877,In_1872);
or U3937 (N_3937,In_124,In_1005);
xor U3938 (N_3938,In_1882,In_851);
xnor U3939 (N_3939,In_318,In_1354);
nand U3940 (N_3940,In_1081,In_911);
and U3941 (N_3941,In_537,In_352);
or U3942 (N_3942,In_931,In_903);
or U3943 (N_3943,In_523,In_1009);
or U3944 (N_3944,In_216,In_1770);
nand U3945 (N_3945,In_1323,In_1740);
and U3946 (N_3946,In_1738,In_1102);
or U3947 (N_3947,In_389,In_373);
nor U3948 (N_3948,In_1004,In_1573);
or U3949 (N_3949,In_26,In_1330);
or U3950 (N_3950,In_1457,In_368);
and U3951 (N_3951,In_368,In_1649);
xor U3952 (N_3952,In_1836,In_776);
and U3953 (N_3953,In_810,In_1683);
and U3954 (N_3954,In_1480,In_1307);
nor U3955 (N_3955,In_620,In_101);
xnor U3956 (N_3956,In_1123,In_1090);
and U3957 (N_3957,In_1508,In_617);
nor U3958 (N_3958,In_1221,In_446);
xor U3959 (N_3959,In_1499,In_789);
nor U3960 (N_3960,In_1232,In_1006);
and U3961 (N_3961,In_769,In_1413);
and U3962 (N_3962,In_1961,In_1709);
nor U3963 (N_3963,In_855,In_1758);
nand U3964 (N_3964,In_81,In_264);
xnor U3965 (N_3965,In_1074,In_529);
nand U3966 (N_3966,In_1018,In_794);
nor U3967 (N_3967,In_374,In_994);
nand U3968 (N_3968,In_147,In_1225);
nor U3969 (N_3969,In_1363,In_811);
nand U3970 (N_3970,In_434,In_857);
and U3971 (N_3971,In_673,In_1240);
xor U3972 (N_3972,In_1207,In_776);
nand U3973 (N_3973,In_1336,In_1816);
xor U3974 (N_3974,In_1704,In_1226);
and U3975 (N_3975,In_702,In_1643);
nand U3976 (N_3976,In_644,In_689);
nand U3977 (N_3977,In_1137,In_1399);
xnor U3978 (N_3978,In_488,In_1178);
or U3979 (N_3979,In_772,In_1238);
nand U3980 (N_3980,In_655,In_737);
nor U3981 (N_3981,In_219,In_461);
or U3982 (N_3982,In_1695,In_875);
or U3983 (N_3983,In_1018,In_1121);
xnor U3984 (N_3984,In_645,In_570);
nor U3985 (N_3985,In_438,In_345);
nor U3986 (N_3986,In_125,In_1490);
xor U3987 (N_3987,In_152,In_1059);
xnor U3988 (N_3988,In_870,In_1002);
nand U3989 (N_3989,In_223,In_1125);
xnor U3990 (N_3990,In_810,In_1511);
and U3991 (N_3991,In_1735,In_382);
and U3992 (N_3992,In_1351,In_781);
nor U3993 (N_3993,In_1089,In_326);
and U3994 (N_3994,In_1660,In_826);
xor U3995 (N_3995,In_575,In_232);
nand U3996 (N_3996,In_836,In_841);
and U3997 (N_3997,In_204,In_1560);
and U3998 (N_3998,In_1346,In_878);
and U3999 (N_3999,In_3,In_1406);
xnor U4000 (N_4000,N_3023,N_1281);
or U4001 (N_4001,N_2952,N_913);
or U4002 (N_4002,N_3444,N_970);
nor U4003 (N_4003,N_95,N_3824);
or U4004 (N_4004,N_3475,N_73);
xor U4005 (N_4005,N_1805,N_2708);
xnor U4006 (N_4006,N_882,N_2801);
or U4007 (N_4007,N_2895,N_3188);
nor U4008 (N_4008,N_2403,N_3976);
nor U4009 (N_4009,N_647,N_2618);
xnor U4010 (N_4010,N_3116,N_1750);
nand U4011 (N_4011,N_220,N_1225);
nand U4012 (N_4012,N_126,N_847);
or U4013 (N_4013,N_1504,N_3187);
or U4014 (N_4014,N_34,N_3120);
xnor U4015 (N_4015,N_4,N_3590);
or U4016 (N_4016,N_1407,N_544);
or U4017 (N_4017,N_1951,N_3496);
nand U4018 (N_4018,N_1467,N_3529);
nand U4019 (N_4019,N_3431,N_1239);
nand U4020 (N_4020,N_2941,N_1617);
xor U4021 (N_4021,N_370,N_3509);
nor U4022 (N_4022,N_2164,N_3884);
or U4023 (N_4023,N_21,N_3858);
nor U4024 (N_4024,N_2770,N_56);
nand U4025 (N_4025,N_3576,N_1672);
nand U4026 (N_4026,N_2898,N_2358);
nand U4027 (N_4027,N_3546,N_1860);
nor U4028 (N_4028,N_3470,N_2589);
nor U4029 (N_4029,N_2319,N_2094);
or U4030 (N_4030,N_3071,N_3512);
nor U4031 (N_4031,N_908,N_2191);
or U4032 (N_4032,N_2310,N_2957);
or U4033 (N_4033,N_2900,N_805);
nor U4034 (N_4034,N_162,N_525);
or U4035 (N_4035,N_201,N_3243);
nand U4036 (N_4036,N_792,N_164);
nor U4037 (N_4037,N_1279,N_3629);
and U4038 (N_4038,N_2307,N_2679);
and U4039 (N_4039,N_1027,N_31);
or U4040 (N_4040,N_2919,N_1587);
or U4041 (N_4041,N_1775,N_2486);
nand U4042 (N_4042,N_920,N_502);
nand U4043 (N_4043,N_3753,N_1479);
or U4044 (N_4044,N_2045,N_341);
nor U4045 (N_4045,N_33,N_3506);
and U4046 (N_4046,N_1584,N_1622);
nand U4047 (N_4047,N_3485,N_497);
nor U4048 (N_4048,N_864,N_541);
and U4049 (N_4049,N_1194,N_535);
or U4050 (N_4050,N_415,N_3736);
or U4051 (N_4051,N_3683,N_866);
xor U4052 (N_4052,N_476,N_2217);
or U4053 (N_4053,N_2138,N_3096);
xor U4054 (N_4054,N_1289,N_3796);
nand U4055 (N_4055,N_3272,N_3015);
and U4056 (N_4056,N_918,N_1862);
and U4057 (N_4057,N_3534,N_2264);
nand U4058 (N_4058,N_1261,N_3981);
nand U4059 (N_4059,N_1947,N_270);
nand U4060 (N_4060,N_246,N_799);
and U4061 (N_4061,N_3893,N_3494);
or U4062 (N_4062,N_3920,N_2093);
nand U4063 (N_4063,N_3806,N_937);
xor U4064 (N_4064,N_2354,N_1842);
nor U4065 (N_4065,N_2864,N_3702);
and U4066 (N_4066,N_396,N_3403);
nor U4067 (N_4067,N_2567,N_3548);
or U4068 (N_4068,N_1403,N_2577);
xor U4069 (N_4069,N_1123,N_2306);
nand U4070 (N_4070,N_2800,N_2650);
or U4071 (N_4071,N_3533,N_3793);
nand U4072 (N_4072,N_3021,N_668);
nor U4073 (N_4073,N_2112,N_406);
nor U4074 (N_4074,N_1188,N_3507);
nand U4075 (N_4075,N_3776,N_3360);
nand U4076 (N_4076,N_3693,N_3684);
or U4077 (N_4077,N_3678,N_1374);
nand U4078 (N_4078,N_2980,N_1573);
xor U4079 (N_4079,N_3751,N_3337);
nor U4080 (N_4080,N_1868,N_2869);
nand U4081 (N_4081,N_1711,N_3685);
nor U4082 (N_4082,N_3038,N_1925);
and U4083 (N_4083,N_218,N_2498);
or U4084 (N_4084,N_815,N_955);
or U4085 (N_4085,N_1898,N_2436);
and U4086 (N_4086,N_1344,N_1994);
xnor U4087 (N_4087,N_2953,N_1393);
xor U4088 (N_4088,N_372,N_921);
and U4089 (N_4089,N_971,N_1782);
nand U4090 (N_4090,N_631,N_1710);
nor U4091 (N_4091,N_2202,N_1468);
nand U4092 (N_4092,N_2735,N_2853);
or U4093 (N_4093,N_249,N_3962);
nor U4094 (N_4094,N_2846,N_1424);
and U4095 (N_4095,N_1899,N_2553);
nor U4096 (N_4096,N_1248,N_3564);
nor U4097 (N_4097,N_707,N_1462);
nor U4098 (N_4098,N_3321,N_3316);
or U4099 (N_4099,N_3923,N_3906);
and U4100 (N_4100,N_3450,N_2825);
nand U4101 (N_4101,N_3220,N_2361);
or U4102 (N_4102,N_2224,N_1223);
nor U4103 (N_4103,N_2756,N_1278);
xnor U4104 (N_4104,N_1777,N_3457);
or U4105 (N_4105,N_1618,N_2990);
xnor U4106 (N_4106,N_2,N_771);
or U4107 (N_4107,N_3274,N_3613);
and U4108 (N_4108,N_204,N_992);
xor U4109 (N_4109,N_1574,N_2611);
nor U4110 (N_4110,N_3675,N_2249);
and U4111 (N_4111,N_1316,N_3643);
nor U4112 (N_4112,N_1724,N_1355);
xor U4113 (N_4113,N_836,N_2592);
xnor U4114 (N_4114,N_858,N_738);
or U4115 (N_4115,N_3549,N_616);
xnor U4116 (N_4116,N_3789,N_1816);
and U4117 (N_4117,N_1492,N_2017);
and U4118 (N_4118,N_3260,N_1695);
and U4119 (N_4119,N_2487,N_1077);
xor U4120 (N_4120,N_2186,N_3612);
nor U4121 (N_4121,N_2771,N_2451);
or U4122 (N_4122,N_935,N_2473);
nand U4123 (N_4123,N_3184,N_2751);
or U4124 (N_4124,N_834,N_3451);
xnor U4125 (N_4125,N_1890,N_290);
or U4126 (N_4126,N_1160,N_1713);
or U4127 (N_4127,N_2190,N_3869);
or U4128 (N_4128,N_491,N_548);
nor U4129 (N_4129,N_2137,N_3039);
nor U4130 (N_4130,N_2839,N_589);
xor U4131 (N_4131,N_3910,N_1290);
or U4132 (N_4132,N_3126,N_152);
or U4133 (N_4133,N_1082,N_781);
xor U4134 (N_4134,N_915,N_1485);
xnor U4135 (N_4135,N_1737,N_3861);
or U4136 (N_4136,N_678,N_710);
nand U4137 (N_4137,N_1146,N_3498);
and U4138 (N_4138,N_1671,N_3086);
or U4139 (N_4139,N_365,N_2344);
nor U4140 (N_4140,N_2485,N_1444);
nor U4141 (N_4141,N_354,N_3449);
and U4142 (N_4142,N_2764,N_2605);
nor U4143 (N_4143,N_596,N_1885);
nand U4144 (N_4144,N_1092,N_2244);
nor U4145 (N_4145,N_1981,N_1634);
and U4146 (N_4146,N_330,N_1635);
and U4147 (N_4147,N_459,N_3010);
and U4148 (N_4148,N_227,N_2871);
xnor U4149 (N_4149,N_1426,N_3939);
xnor U4150 (N_4150,N_2969,N_376);
xor U4151 (N_4151,N_1208,N_3222);
or U4152 (N_4152,N_2144,N_1230);
nand U4153 (N_4153,N_1073,N_195);
and U4154 (N_4154,N_3924,N_3456);
nand U4155 (N_4155,N_482,N_437);
and U4156 (N_4156,N_508,N_3179);
and U4157 (N_4157,N_3617,N_465);
xnor U4158 (N_4158,N_2755,N_1387);
xor U4159 (N_4159,N_3281,N_2608);
nand U4160 (N_4160,N_665,N_2377);
xor U4161 (N_4161,N_730,N_3836);
and U4162 (N_4162,N_1464,N_1756);
nor U4163 (N_4163,N_1833,N_927);
xor U4164 (N_4164,N_2099,N_747);
or U4165 (N_4165,N_2215,N_3302);
xor U4166 (N_4166,N_948,N_280);
xnor U4167 (N_4167,N_2599,N_2302);
and U4168 (N_4168,N_3294,N_2011);
xor U4169 (N_4169,N_884,N_1997);
nand U4170 (N_4170,N_3365,N_2899);
or U4171 (N_4171,N_1484,N_111);
nand U4172 (N_4172,N_3659,N_2375);
and U4173 (N_4173,N_3523,N_2822);
nand U4174 (N_4174,N_3959,N_456);
nand U4175 (N_4175,N_1743,N_2496);
nor U4176 (N_4176,N_1832,N_2247);
nand U4177 (N_4177,N_1720,N_307);
xor U4178 (N_4178,N_3041,N_3415);
nor U4179 (N_4179,N_1345,N_1528);
nor U4180 (N_4180,N_1633,N_2643);
nor U4181 (N_4181,N_368,N_2297);
nor U4182 (N_4182,N_3845,N_1268);
nand U4183 (N_4183,N_573,N_1619);
and U4184 (N_4184,N_2033,N_2142);
nor U4185 (N_4185,N_2598,N_976);
or U4186 (N_4186,N_2987,N_440);
nand U4187 (N_4187,N_1326,N_2397);
and U4188 (N_4188,N_2564,N_3905);
nand U4189 (N_4189,N_718,N_2471);
nand U4190 (N_4190,N_2006,N_1338);
nor U4191 (N_4191,N_375,N_3263);
or U4192 (N_4192,N_3606,N_1181);
xnor U4193 (N_4193,N_3467,N_473);
or U4194 (N_4194,N_3600,N_2578);
and U4195 (N_4195,N_523,N_2656);
nor U4196 (N_4196,N_2418,N_1417);
nor U4197 (N_4197,N_3825,N_1849);
nand U4198 (N_4198,N_3952,N_3524);
nor U4199 (N_4199,N_568,N_1150);
or U4200 (N_4200,N_1299,N_2863);
nand U4201 (N_4201,N_3358,N_3816);
or U4202 (N_4202,N_1740,N_680);
xor U4203 (N_4203,N_591,N_1983);
or U4204 (N_4204,N_18,N_943);
or U4205 (N_4205,N_3327,N_3515);
xor U4206 (N_4206,N_3503,N_166);
xnor U4207 (N_4207,N_1570,N_3110);
xnor U4208 (N_4208,N_1480,N_874);
nand U4209 (N_4209,N_3822,N_3723);
or U4210 (N_4210,N_416,N_3938);
nor U4211 (N_4211,N_392,N_3622);
or U4212 (N_4212,N_2360,N_1565);
or U4213 (N_4213,N_426,N_2075);
or U4214 (N_4214,N_2688,N_3244);
xnor U4215 (N_4215,N_2491,N_2661);
and U4216 (N_4216,N_2676,N_1663);
nor U4217 (N_4217,N_1309,N_2862);
xor U4218 (N_4218,N_1943,N_1844);
or U4219 (N_4219,N_2887,N_2013);
nor U4220 (N_4220,N_2586,N_1677);
nand U4221 (N_4221,N_277,N_3649);
nand U4222 (N_4222,N_1478,N_2012);
xor U4223 (N_4223,N_2736,N_959);
and U4224 (N_4224,N_3504,N_1033);
xnor U4225 (N_4225,N_2162,N_3602);
and U4226 (N_4226,N_658,N_438);
nand U4227 (N_4227,N_956,N_2734);
xnor U4228 (N_4228,N_1975,N_261);
xnor U4229 (N_4229,N_2235,N_2762);
and U4230 (N_4230,N_2628,N_2369);
nor U4231 (N_4231,N_694,N_1946);
nand U4232 (N_4232,N_511,N_1763);
xnor U4233 (N_4233,N_505,N_1283);
nand U4234 (N_4234,N_1390,N_1297);
nand U4235 (N_4235,N_3551,N_2313);
and U4236 (N_4236,N_1076,N_2902);
or U4237 (N_4237,N_952,N_688);
nand U4238 (N_4238,N_3291,N_474);
or U4239 (N_4239,N_3625,N_540);
xor U4240 (N_4240,N_1138,N_3781);
nor U4241 (N_4241,N_2081,N_1689);
or U4242 (N_4242,N_788,N_3757);
nor U4243 (N_4243,N_1116,N_225);
nand U4244 (N_4244,N_1219,N_37);
nand U4245 (N_4245,N_3248,N_234);
nand U4246 (N_4246,N_1628,N_3348);
nand U4247 (N_4247,N_2936,N_253);
nand U4248 (N_4248,N_3441,N_3607);
nor U4249 (N_4249,N_2285,N_760);
nor U4250 (N_4250,N_1031,N_916);
or U4251 (N_4251,N_2972,N_1674);
xor U4252 (N_4252,N_1159,N_1402);
and U4253 (N_4253,N_853,N_3968);
or U4254 (N_4254,N_711,N_3306);
xor U4255 (N_4255,N_627,N_1568);
xor U4256 (N_4256,N_1666,N_993);
nor U4257 (N_4257,N_2866,N_3577);
and U4258 (N_4258,N_973,N_3091);
nand U4259 (N_4259,N_845,N_3267);
nor U4260 (N_4260,N_554,N_1255);
or U4261 (N_4261,N_332,N_3763);
or U4262 (N_4262,N_1836,N_3278);
xnor U4263 (N_4263,N_708,N_278);
xnor U4264 (N_4264,N_2289,N_1643);
and U4265 (N_4265,N_1662,N_2644);
nor U4266 (N_4266,N_401,N_910);
nand U4267 (N_4267,N_1420,N_1771);
xor U4268 (N_4268,N_77,N_1825);
or U4269 (N_4269,N_320,N_2018);
xor U4270 (N_4270,N_2410,N_1115);
nand U4271 (N_4271,N_1460,N_563);
xor U4272 (N_4272,N_3668,N_3801);
or U4273 (N_4273,N_3090,N_20);
nor U4274 (N_4274,N_531,N_1175);
and U4275 (N_4275,N_1329,N_495);
xor U4276 (N_4276,N_1973,N_789);
or U4277 (N_4277,N_3212,N_1629);
nand U4278 (N_4278,N_1614,N_3364);
and U4279 (N_4279,N_184,N_3644);
nor U4280 (N_4280,N_2897,N_44);
or U4281 (N_4281,N_2114,N_351);
nor U4282 (N_4282,N_2096,N_3676);
nand U4283 (N_4283,N_1598,N_264);
nand U4284 (N_4284,N_3448,N_488);
or U4285 (N_4285,N_2229,N_2245);
and U4286 (N_4286,N_3854,N_2110);
nand U4287 (N_4287,N_3129,N_3565);
xor U4288 (N_4288,N_1386,N_3235);
nor U4289 (N_4289,N_2696,N_1398);
xor U4290 (N_4290,N_3987,N_1829);
or U4291 (N_4291,N_3759,N_1843);
or U4292 (N_4292,N_2423,N_1045);
or U4293 (N_4293,N_2893,N_1960);
or U4294 (N_4294,N_765,N_3252);
or U4295 (N_4295,N_1024,N_527);
or U4296 (N_4296,N_2063,N_499);
nor U4297 (N_4297,N_3588,N_802);
xor U4298 (N_4298,N_2200,N_1220);
nor U4299 (N_4299,N_1957,N_2753);
and U4300 (N_4300,N_475,N_3902);
xnor U4301 (N_4301,N_2205,N_782);
nor U4302 (N_4302,N_859,N_2689);
nor U4303 (N_4303,N_2083,N_776);
nor U4304 (N_4304,N_41,N_26);
xor U4305 (N_4305,N_1922,N_298);
or U4306 (N_4306,N_3308,N_127);
or U4307 (N_4307,N_2341,N_1394);
or U4308 (N_4308,N_3626,N_2007);
xnor U4309 (N_4309,N_569,N_1526);
xnor U4310 (N_4310,N_388,N_2729);
nand U4311 (N_4311,N_3866,N_1515);
xnor U4312 (N_4312,N_912,N_3724);
xnor U4313 (N_4313,N_294,N_385);
nand U4314 (N_4314,N_2796,N_186);
xor U4315 (N_4315,N_1902,N_562);
nand U4316 (N_4316,N_3257,N_1800);
nand U4317 (N_4317,N_2185,N_504);
nand U4318 (N_4318,N_529,N_3390);
nand U4319 (N_4319,N_1105,N_93);
xor U4320 (N_4320,N_232,N_3557);
or U4321 (N_4321,N_2971,N_3961);
or U4322 (N_4322,N_2118,N_2444);
or U4323 (N_4323,N_3885,N_2010);
xnor U4324 (N_4324,N_871,N_2746);
nor U4325 (N_4325,N_672,N_2167);
or U4326 (N_4326,N_1164,N_1243);
or U4327 (N_4327,N_763,N_395);
and U4328 (N_4328,N_1717,N_2930);
xor U4329 (N_4329,N_693,N_2973);
nand U4330 (N_4330,N_2353,N_2653);
or U4331 (N_4331,N_870,N_3249);
nor U4332 (N_4332,N_1380,N_1524);
or U4333 (N_4333,N_2402,N_2311);
nor U4334 (N_4334,N_599,N_2945);
xnor U4335 (N_4335,N_808,N_2911);
xnor U4336 (N_4336,N_216,N_720);
or U4337 (N_4337,N_3933,N_2937);
and U4338 (N_4338,N_2488,N_1419);
nor U4339 (N_4339,N_2068,N_1995);
nand U4340 (N_4340,N_2576,N_3057);
nand U4341 (N_4341,N_192,N_594);
or U4342 (N_4342,N_1486,N_1483);
nor U4343 (N_4343,N_3640,N_2482);
xor U4344 (N_4344,N_825,N_3677);
xnor U4345 (N_4345,N_1974,N_2615);
xnor U4346 (N_4346,N_315,N_1755);
xor U4347 (N_4347,N_2808,N_2391);
xnor U4348 (N_4348,N_1228,N_1335);
and U4349 (N_4349,N_297,N_10);
and U4350 (N_4350,N_609,N_1752);
nor U4351 (N_4351,N_1648,N_3554);
nor U4352 (N_4352,N_2121,N_830);
nor U4353 (N_4353,N_2398,N_2681);
and U4354 (N_4354,N_3881,N_3133);
and U4355 (N_4355,N_1804,N_986);
or U4356 (N_4356,N_2909,N_1719);
and U4357 (N_4357,N_942,N_3024);
nor U4358 (N_4358,N_2888,N_480);
and U4359 (N_4359,N_1507,N_2935);
or U4360 (N_4360,N_773,N_2819);
and U4361 (N_4361,N_1636,N_1915);
nor U4362 (N_4362,N_173,N_997);
nand U4363 (N_4363,N_3849,N_3349);
nor U4364 (N_4364,N_3972,N_1976);
or U4365 (N_4365,N_284,N_3208);
xor U4366 (N_4366,N_1348,N_1064);
or U4367 (N_4367,N_3234,N_3592);
or U4368 (N_4368,N_1411,N_1137);
and U4369 (N_4369,N_3639,N_1611);
xnor U4370 (N_4370,N_50,N_222);
and U4371 (N_4371,N_1182,N_610);
and U4372 (N_4372,N_724,N_1000);
or U4373 (N_4373,N_3713,N_2145);
xnor U4374 (N_4374,N_2085,N_2886);
xor U4375 (N_4375,N_2654,N_1513);
nor U4376 (N_4376,N_3755,N_3383);
xor U4377 (N_4377,N_102,N_1012);
nor U4378 (N_4378,N_3814,N_3988);
and U4379 (N_4379,N_1798,N_2721);
nand U4380 (N_4380,N_78,N_2526);
nor U4381 (N_4381,N_2194,N_1726);
nand U4382 (N_4382,N_9,N_1530);
xor U4383 (N_4383,N_3690,N_1416);
nand U4384 (N_4384,N_2505,N_798);
xor U4385 (N_4385,N_831,N_2804);
xor U4386 (N_4386,N_3058,N_2959);
and U4387 (N_4387,N_287,N_2981);
and U4388 (N_4388,N_1207,N_2772);
and U4389 (N_4389,N_140,N_3971);
xor U4390 (N_4390,N_160,N_2443);
nor U4391 (N_4391,N_3773,N_1108);
or U4392 (N_4392,N_311,N_3811);
nand U4393 (N_4393,N_2533,N_1660);
nor U4394 (N_4394,N_1971,N_1776);
nor U4395 (N_4395,N_2831,N_3199);
nor U4396 (N_4396,N_786,N_2292);
nand U4397 (N_4397,N_1015,N_2627);
xnor U4398 (N_4398,N_2633,N_457);
xnor U4399 (N_4399,N_2793,N_2748);
or U4400 (N_4400,N_2466,N_3191);
and U4401 (N_4401,N_313,N_1315);
xor U4402 (N_4402,N_1632,N_1809);
and U4403 (N_4403,N_1746,N_3001);
nor U4404 (N_4404,N_3810,N_468);
nand U4405 (N_4405,N_3452,N_2697);
nand U4406 (N_4406,N_1692,N_1494);
xnor U4407 (N_4407,N_1149,N_2064);
and U4408 (N_4408,N_2457,N_3236);
nand U4409 (N_4409,N_2580,N_3397);
nor U4410 (N_4410,N_2960,N_2701);
or U4411 (N_4411,N_2216,N_1291);
and U4412 (N_4412,N_3673,N_946);
or U4413 (N_4413,N_2231,N_3786);
nor U4414 (N_4414,N_3632,N_2690);
or U4415 (N_4415,N_318,N_2431);
and U4416 (N_4416,N_2780,N_3157);
or U4417 (N_4417,N_3935,N_2738);
and U4418 (N_4418,N_1556,N_1491);
xor U4419 (N_4419,N_1133,N_1933);
xor U4420 (N_4420,N_1023,N_3273);
and U4421 (N_4421,N_3510,N_2976);
or U4422 (N_4422,N_3570,N_3293);
and U4423 (N_4423,N_2784,N_461);
nand U4424 (N_4424,N_2835,N_861);
and U4425 (N_4425,N_1053,N_3730);
or U4426 (N_4426,N_3508,N_2035);
nor U4427 (N_4427,N_3237,N_1806);
nor U4428 (N_4428,N_2115,N_1900);
xor U4429 (N_4429,N_3746,N_2623);
or U4430 (N_4430,N_750,N_2521);
nor U4431 (N_4431,N_1373,N_549);
or U4432 (N_4432,N_143,N_3547);
xor U4433 (N_4433,N_3522,N_3221);
nor U4434 (N_4434,N_1979,N_2108);
or U4435 (N_4435,N_2910,N_1909);
nand U4436 (N_4436,N_2585,N_2761);
nand U4437 (N_4437,N_3813,N_757);
or U4438 (N_4438,N_3653,N_1233);
nor U4439 (N_4439,N_3595,N_2299);
or U4440 (N_4440,N_953,N_1826);
nor U4441 (N_4441,N_231,N_2940);
nor U4442 (N_4442,N_863,N_2587);
xor U4443 (N_4443,N_2896,N_3050);
nor U4444 (N_4444,N_2868,N_2401);
or U4445 (N_4445,N_2885,N_2683);
and U4446 (N_4446,N_2539,N_1381);
and U4447 (N_4447,N_2345,N_151);
or U4448 (N_4448,N_1729,N_3253);
nor U4449 (N_4449,N_3404,N_1131);
and U4450 (N_4450,N_1376,N_2253);
nand U4451 (N_4451,N_3658,N_2575);
xnor U4452 (N_4452,N_1203,N_1014);
nor U4453 (N_4453,N_2464,N_2206);
nand U4454 (N_4454,N_2320,N_2130);
xor U4455 (N_4455,N_3324,N_1287);
and U4456 (N_4456,N_206,N_342);
or U4457 (N_4457,N_2693,N_1429);
and U4458 (N_4458,N_3284,N_2504);
nand U4459 (N_4459,N_3492,N_613);
and U4460 (N_4460,N_2616,N_1964);
and U4461 (N_4461,N_2750,N_1953);
nor U4462 (N_4462,N_3648,N_1705);
nand U4463 (N_4463,N_3165,N_2924);
or U4464 (N_4464,N_876,N_2991);
nor U4465 (N_4465,N_2022,N_1594);
nor U4466 (N_4466,N_1699,N_3768);
nor U4467 (N_4467,N_2610,N_1452);
xnor U4468 (N_4468,N_1349,N_2023);
nor U4469 (N_4469,N_3550,N_816);
or U4470 (N_4470,N_3687,N_3876);
and U4471 (N_4471,N_112,N_3998);
and U4472 (N_4472,N_3213,N_1401);
or U4473 (N_4473,N_1231,N_2889);
nand U4474 (N_4474,N_3473,N_263);
nand U4475 (N_4475,N_1659,N_713);
and U4476 (N_4476,N_657,N_2844);
and U4477 (N_4477,N_700,N_2270);
xnor U4478 (N_4478,N_2706,N_1437);
nor U4479 (N_4479,N_3282,N_2393);
nor U4480 (N_4480,N_2026,N_2707);
xnor U4481 (N_4481,N_1582,N_1496);
nand U4482 (N_4482,N_1317,N_1272);
or U4483 (N_4483,N_110,N_3800);
or U4484 (N_4484,N_3720,N_3647);
nand U4485 (N_4485,N_2579,N_560);
and U4486 (N_4486,N_3717,N_2284);
xnor U4487 (N_4487,N_2597,N_174);
and U4488 (N_4488,N_2630,N_3931);
xor U4489 (N_4489,N_1210,N_2055);
nand U4490 (N_4490,N_2407,N_829);
nor U4491 (N_4491,N_3040,N_303);
xnor U4492 (N_4492,N_2970,N_2645);
and U4493 (N_4493,N_1180,N_827);
nand U4494 (N_4494,N_1924,N_2333);
and U4495 (N_4495,N_593,N_486);
xor U4496 (N_4496,N_3335,N_3525);
or U4497 (N_4497,N_3121,N_1642);
nand U4498 (N_4498,N_3105,N_571);
or U4499 (N_4499,N_1564,N_1110);
or U4500 (N_4500,N_1371,N_2478);
or U4501 (N_4501,N_3788,N_3582);
xor U4502 (N_4502,N_3589,N_382);
nor U4503 (N_4503,N_479,N_2845);
xnor U4504 (N_4504,N_642,N_1880);
and U4505 (N_4505,N_62,N_1709);
nand U4506 (N_4506,N_2716,N_1578);
and U4507 (N_4507,N_841,N_3352);
and U4508 (N_4508,N_1512,N_405);
nand U4509 (N_4509,N_939,N_75);
and U4510 (N_4510,N_739,N_1436);
xnor U4511 (N_4511,N_2648,N_3064);
and U4512 (N_4512,N_3268,N_3478);
xnor U4513 (N_4513,N_3447,N_1227);
xor U4514 (N_4514,N_1969,N_821);
and U4515 (N_4515,N_3181,N_1382);
and U4516 (N_4516,N_3967,N_3775);
and U4517 (N_4517,N_2983,N_1414);
or U4518 (N_4518,N_2283,N_3598);
nand U4519 (N_4519,N_1550,N_2104);
or U4520 (N_4520,N_412,N_97);
nor U4521 (N_4521,N_3476,N_3505);
nand U4522 (N_4522,N_3715,N_1448);
nor U4523 (N_4523,N_229,N_2038);
or U4524 (N_4524,N_2421,N_304);
or U4525 (N_4525,N_2454,N_702);
nand U4526 (N_4526,N_1758,N_2056);
or U4527 (N_4527,N_1120,N_2754);
nor U4528 (N_4528,N_1872,N_3226);
nand U4529 (N_4529,N_2877,N_2140);
or U4530 (N_4530,N_3738,N_87);
nand U4531 (N_4531,N_1883,N_17);
or U4532 (N_4532,N_439,N_2776);
xnor U4533 (N_4533,N_310,N_621);
or U4534 (N_4534,N_2084,N_1089);
xor U4535 (N_4535,N_2327,N_2647);
nor U4536 (N_4536,N_1410,N_444);
and U4537 (N_4537,N_1029,N_445);
nor U4538 (N_4538,N_3742,N_417);
nand U4539 (N_4539,N_1135,N_2204);
nand U4540 (N_4540,N_2066,N_3699);
xnor U4541 (N_4541,N_2717,N_2014);
nand U4542 (N_4542,N_1802,N_3883);
and U4543 (N_4543,N_2040,N_620);
nor U4544 (N_4544,N_3331,N_1575);
and U4545 (N_4545,N_3180,N_54);
and U4546 (N_4546,N_2400,N_1679);
and U4547 (N_4547,N_178,N_3318);
nand U4548 (N_4548,N_1546,N_470);
and U4549 (N_4549,N_3454,N_3667);
xor U4550 (N_4550,N_2483,N_1232);
or U4551 (N_4551,N_1409,N_1132);
xor U4552 (N_4552,N_3210,N_2078);
nor U4553 (N_4553,N_2034,N_1347);
nor U4554 (N_4554,N_12,N_767);
xnor U4555 (N_4555,N_2422,N_2370);
nor U4556 (N_4556,N_1537,N_3163);
or U4557 (N_4557,N_3892,N_1122);
and U4558 (N_4558,N_2170,N_1375);
nand U4559 (N_4559,N_1519,N_1070);
nor U4560 (N_4560,N_2057,N_814);
nand U4561 (N_4561,N_3037,N_3238);
or U4562 (N_4562,N_2903,N_2348);
xnor U4563 (N_4563,N_3139,N_3879);
and U4564 (N_4564,N_3936,N_3873);
xnor U4565 (N_4565,N_2543,N_1787);
xor U4566 (N_4566,N_3727,N_2020);
or U4567 (N_4567,N_1229,N_35);
nand U4568 (N_4568,N_3309,N_3488);
and U4569 (N_4569,N_1897,N_1655);
and U4570 (N_4570,N_3423,N_2159);
xor U4571 (N_4571,N_3154,N_1905);
xnor U4572 (N_4572,N_134,N_1544);
and U4573 (N_4573,N_1647,N_1966);
nand U4574 (N_4574,N_1047,N_2143);
xor U4575 (N_4575,N_2542,N_3843);
or U4576 (N_4576,N_746,N_2614);
nand U4577 (N_4577,N_1783,N_3927);
nor U4578 (N_4578,N_2540,N_2472);
or U4579 (N_4579,N_1050,N_2126);
and U4580 (N_4580,N_2519,N_1903);
and U4581 (N_4581,N_2467,N_2453);
nand U4582 (N_4582,N_588,N_3563);
xor U4583 (N_4583,N_3756,N_3127);
and U4584 (N_4584,N_3880,N_3095);
and U4585 (N_4585,N_3314,N_2856);
nand U4586 (N_4586,N_300,N_2830);
xnor U4587 (N_4587,N_3279,N_3292);
nand U4588 (N_4588,N_817,N_1236);
nand U4589 (N_4589,N_1238,N_325);
and U4590 (N_4590,N_2399,N_1352);
and U4591 (N_4591,N_2925,N_3597);
nand U4592 (N_4592,N_1497,N_877);
xnor U4593 (N_4593,N_936,N_3679);
xnor U4594 (N_4594,N_1621,N_1521);
xor U4595 (N_4595,N_434,N_1010);
nand U4596 (N_4596,N_2946,N_1658);
nor U4597 (N_4597,N_450,N_196);
and U4598 (N_4598,N_451,N_3074);
nor U4599 (N_4599,N_1147,N_3044);
and U4600 (N_4600,N_1189,N_2415);
nor U4601 (N_4601,N_1780,N_3144);
xnor U4602 (N_4602,N_533,N_2290);
or U4603 (N_4603,N_349,N_3148);
nand U4604 (N_4604,N_1697,N_2184);
xor U4605 (N_4605,N_2827,N_2203);
or U4606 (N_4606,N_2221,N_1245);
and U4607 (N_4607,N_3299,N_2922);
and U4608 (N_4608,N_3792,N_1784);
and U4609 (N_4609,N_1036,N_1930);
nand U4610 (N_4610,N_3513,N_3559);
xnor U4611 (N_4611,N_3614,N_175);
xor U4612 (N_4612,N_214,N_1368);
and U4613 (N_4613,N_2635,N_27);
nor U4614 (N_4614,N_251,N_630);
nand U4615 (N_4615,N_2807,N_509);
or U4616 (N_4616,N_2069,N_2537);
nor U4617 (N_4617,N_3764,N_3633);
and U4618 (N_4618,N_43,N_3578);
and U4619 (N_4619,N_2476,N_1989);
nand U4620 (N_4620,N_2912,N_3377);
xor U4621 (N_4621,N_1177,N_1701);
nand U4622 (N_4622,N_2914,N_3735);
and U4623 (N_4623,N_1781,N_1169);
or U4624 (N_4624,N_2420,N_1079);
nand U4625 (N_4625,N_536,N_3914);
and U4626 (N_4626,N_3288,N_1532);
nor U4627 (N_4627,N_213,N_938);
and U4628 (N_4628,N_949,N_506);
nor U4629 (N_4629,N_1367,N_1435);
and U4630 (N_4630,N_2649,N_3138);
nor U4631 (N_4631,N_89,N_2213);
and U4632 (N_4632,N_2165,N_2658);
nand U4633 (N_4633,N_1102,N_1912);
or U4634 (N_4634,N_274,N_2282);
nor U4635 (N_4635,N_3501,N_1961);
nor U4636 (N_4636,N_2406,N_242);
or U4637 (N_4637,N_72,N_3201);
xnor U4638 (N_4638,N_1422,N_2923);
nand U4639 (N_4639,N_267,N_189);
nor U4640 (N_4640,N_22,N_2365);
xnor U4641 (N_4641,N_2833,N_2328);
nand U4642 (N_4642,N_326,N_3953);
nand U4643 (N_4643,N_3894,N_266);
nor U4644 (N_4644,N_513,N_557);
nand U4645 (N_4645,N_1857,N_2974);
and U4646 (N_4646,N_3966,N_1919);
or U4647 (N_4647,N_2872,N_1725);
nand U4648 (N_4648,N_1886,N_3895);
or U4649 (N_4649,N_2666,N_3198);
nand U4650 (N_4650,N_3872,N_380);
nand U4651 (N_4651,N_122,N_1412);
nand U4652 (N_4652,N_696,N_2192);
nor U4653 (N_4653,N_91,N_1837);
and U4654 (N_4654,N_1602,N_207);
nand U4655 (N_4655,N_2461,N_3323);
nand U4656 (N_4656,N_431,N_45);
nor U4657 (N_4657,N_3432,N_1962);
xnor U4658 (N_4658,N_364,N_1482);
nor U4659 (N_4659,N_3493,N_682);
or U4660 (N_4660,N_2607,N_576);
nor U4661 (N_4661,N_1580,N_65);
and U4662 (N_4662,N_1968,N_990);
or U4663 (N_4663,N_583,N_2316);
and U4664 (N_4664,N_510,N_3153);
and U4665 (N_4665,N_1209,N_3749);
nor U4666 (N_4666,N_2515,N_914);
nand U4667 (N_4667,N_3651,N_2865);
and U4668 (N_4668,N_3897,N_3944);
or U4669 (N_4669,N_2089,N_2698);
nand U4670 (N_4670,N_329,N_2368);
and U4671 (N_4671,N_3338,N_180);
nand U4672 (N_4672,N_1986,N_237);
or U4673 (N_4673,N_926,N_2481);
or U4674 (N_4674,N_1221,N_3584);
nor U4675 (N_4675,N_397,N_1341);
and U4676 (N_4676,N_907,N_194);
nor U4677 (N_4677,N_1038,N_1500);
xor U4678 (N_4678,N_1514,N_2363);
xnor U4679 (N_4679,N_2612,N_1850);
or U4680 (N_4680,N_1222,N_469);
or U4681 (N_4681,N_1509,N_1163);
nand U4682 (N_4682,N_1723,N_3251);
nand U4683 (N_4683,N_848,N_3002);
or U4684 (N_4684,N_2702,N_3012);
nand U4685 (N_4685,N_3013,N_3922);
or U4686 (N_4686,N_1682,N_1608);
or U4687 (N_4687,N_2685,N_2274);
nand U4688 (N_4688,N_3808,N_3985);
and U4689 (N_4689,N_2506,N_2783);
nand U4690 (N_4690,N_3874,N_3917);
xor U4691 (N_4691,N_1554,N_608);
nor U4692 (N_4692,N_3964,N_2210);
and U4693 (N_4693,N_2392,N_2331);
nor U4694 (N_4694,N_1797,N_754);
or U4695 (N_4695,N_1342,N_3994);
or U4696 (N_4696,N_3461,N_626);
xnor U4697 (N_4697,N_3712,N_1404);
and U4698 (N_4698,N_1817,N_520);
xor U4699 (N_4699,N_1799,N_3117);
and U4700 (N_4700,N_363,N_3043);
nand U4701 (N_4701,N_1008,N_3631);
nor U4702 (N_4702,N_2582,N_3169);
and U4703 (N_4703,N_2220,N_1835);
and U4704 (N_4704,N_2549,N_994);
nand U4705 (N_4705,N_2052,N_3558);
nor U4706 (N_4706,N_295,N_159);
xnor U4707 (N_4707,N_3830,N_1988);
and U4708 (N_4708,N_2269,N_706);
and U4709 (N_4709,N_2424,N_1296);
or U4710 (N_4710,N_359,N_1035);
nor U4711 (N_4711,N_3011,N_1708);
nor U4712 (N_4712,N_2792,N_2309);
or U4713 (N_4713,N_3479,N_995);
or U4714 (N_4714,N_1593,N_1086);
and U4715 (N_4715,N_1728,N_2982);
or U4716 (N_4716,N_3426,N_1310);
xnor U4717 (N_4717,N_3232,N_128);
nor U4718 (N_4718,N_645,N_3921);
nand U4719 (N_4719,N_567,N_3100);
nor U4720 (N_4720,N_2558,N_51);
and U4721 (N_4721,N_3356,N_3051);
nor U4722 (N_4722,N_3307,N_1455);
xnor U4723 (N_4723,N_3280,N_1469);
nor U4724 (N_4724,N_106,N_1848);
xnor U4725 (N_4725,N_2155,N_2222);
or U4726 (N_4726,N_2025,N_3216);
nand U4727 (N_4727,N_1875,N_3124);
nand U4728 (N_4728,N_3490,N_1668);
and U4729 (N_4729,N_2809,N_3254);
and U4730 (N_4730,N_2356,N_2870);
nor U4731 (N_4731,N_3097,N_1827);
xor U4732 (N_4732,N_1249,N_1665);
nor U4733 (N_4733,N_2257,N_1286);
or U4734 (N_4734,N_2258,N_1901);
or U4735 (N_4735,N_2637,N_2890);
nor U4736 (N_4736,N_1277,N_3016);
nand U4737 (N_4737,N_366,N_1273);
nor U4738 (N_4738,N_977,N_689);
nand U4739 (N_4739,N_137,N_2291);
and U4740 (N_4740,N_1214,N_25);
and U4741 (N_4741,N_794,N_3857);
xnor U4742 (N_4742,N_2300,N_2458);
or U4743 (N_4743,N_1906,N_1104);
xor U4744 (N_4744,N_981,N_1044);
and U4745 (N_4745,N_998,N_2039);
and U4746 (N_4746,N_323,N_1768);
xnor U4747 (N_4747,N_2469,N_2594);
or U4748 (N_4748,N_751,N_481);
xnor U4749 (N_4749,N_893,N_1876);
nand U4750 (N_4750,N_1395,N_2076);
xor U4751 (N_4751,N_3141,N_3535);
or U4752 (N_4752,N_1434,N_288);
xnor U4753 (N_4753,N_519,N_1877);
and U4754 (N_4754,N_745,N_3085);
nor U4755 (N_4755,N_3223,N_3459);
and U4756 (N_4756,N_265,N_2321);
nand U4757 (N_4757,N_2449,N_2175);
or U4758 (N_4758,N_3839,N_104);
nand U4759 (N_4759,N_2559,N_32);
nor U4760 (N_4760,N_3954,N_570);
xor U4761 (N_4761,N_1751,N_612);
nor U4762 (N_4762,N_3471,N_3692);
nand U4763 (N_4763,N_2296,N_3500);
nor U4764 (N_4764,N_2484,N_574);
and U4765 (N_4765,N_3787,N_2061);
xnor U4766 (N_4766,N_3663,N_1114);
xor U4767 (N_4767,N_1428,N_1865);
nand U4768 (N_4768,N_331,N_2916);
xnor U4769 (N_4769,N_116,N_135);
nor U4770 (N_4770,N_3204,N_2799);
and U4771 (N_4771,N_1361,N_3744);
nor U4772 (N_4772,N_2152,N_64);
nor U4773 (N_4773,N_1993,N_374);
xor U4774 (N_4774,N_2122,N_2117);
and U4775 (N_4775,N_3560,N_1151);
or U4776 (N_4776,N_1489,N_2816);
or U4777 (N_4777,N_3093,N_1866);
and U4778 (N_4778,N_3783,N_3974);
xor U4779 (N_4779,N_308,N_3929);
nor U4780 (N_4780,N_521,N_967);
xnor U4781 (N_4781,N_2905,N_2875);
or U4782 (N_4782,N_2439,N_756);
or U4783 (N_4783,N_1304,N_3852);
nor U4784 (N_4784,N_1423,N_1558);
nand U4785 (N_4785,N_584,N_1557);
nor U4786 (N_4786,N_305,N_146);
and U4787 (N_4787,N_1950,N_478);
nor U4788 (N_4788,N_447,N_2050);
or U4789 (N_4789,N_1377,N_339);
or U4790 (N_4790,N_321,N_3363);
nand U4791 (N_4791,N_3006,N_3075);
and U4792 (N_4792,N_2355,N_2913);
and U4793 (N_4793,N_224,N_2318);
nand U4794 (N_4794,N_2416,N_2016);
and U4795 (N_4795,N_203,N_3545);
xor U4796 (N_4796,N_2534,N_1891);
and U4797 (N_4797,N_649,N_2759);
nor U4798 (N_4798,N_1421,N_71);
xor U4799 (N_4799,N_124,N_2625);
and U4800 (N_4800,N_3194,N_3132);
and U4801 (N_4801,N_595,N_3708);
nand U4802 (N_4802,N_2984,N_1911);
xor U4803 (N_4803,N_983,N_1028);
and U4804 (N_4804,N_2171,N_3947);
or U4805 (N_4805,N_407,N_2000);
or U4806 (N_4806,N_806,N_3934);
xnor U4807 (N_4807,N_3666,N_2634);
nand U4808 (N_4808,N_335,N_896);
and U4809 (N_4809,N_3820,N_3729);
or U4810 (N_4810,N_1140,N_972);
and U4811 (N_4811,N_843,N_3686);
or U4812 (N_4812,N_3850,N_577);
nand U4813 (N_4813,N_3680,N_3721);
nand U4814 (N_4814,N_3691,N_157);
nand U4815 (N_4815,N_250,N_3645);
and U4816 (N_4816,N_3380,N_3207);
nor U4817 (N_4817,N_356,N_664);
nand U4818 (N_4818,N_837,N_737);
nor U4819 (N_4819,N_1458,N_555);
or U4820 (N_4820,N_666,N_3464);
and U4821 (N_4821,N_723,N_3150);
xor U4822 (N_4822,N_2841,N_975);
or U4823 (N_4823,N_3726,N_553);
xor U4824 (N_4824,N_3999,N_2385);
nand U4825 (N_4825,N_3396,N_906);
or U4826 (N_4826,N_1284,N_1295);
and U4827 (N_4827,N_641,N_1142);
or U4828 (N_4828,N_822,N_1603);
and U4829 (N_4829,N_1605,N_3135);
and U4830 (N_4830,N_1794,N_851);
nand U4831 (N_4831,N_2752,N_878);
or U4832 (N_4832,N_3160,N_3804);
and U4833 (N_4833,N_1184,N_3081);
or U4834 (N_4834,N_3018,N_3700);
and U4835 (N_4835,N_353,N_5);
and U4836 (N_4836,N_2760,N_887);
and U4837 (N_4837,N_501,N_2596);
nand U4838 (N_4838,N_2277,N_2060);
xnor U4839 (N_4839,N_2077,N_1935);
xor U4840 (N_4840,N_3552,N_343);
nand U4841 (N_4841,N_1945,N_3530);
and U4842 (N_4842,N_2268,N_1795);
and U4843 (N_4843,N_1148,N_1360);
nand U4844 (N_4844,N_3532,N_333);
or U4845 (N_4845,N_3076,N_3630);
xor U4846 (N_4846,N_3519,N_2267);
xnor U4847 (N_4847,N_167,N_1785);
xnor U4848 (N_4848,N_3382,N_1257);
xor U4849 (N_4849,N_1936,N_1954);
or U4850 (N_4850,N_2329,N_748);
nor U4851 (N_4851,N_1218,N_2272);
or U4852 (N_4852,N_2758,N_2259);
nor U4853 (N_4853,N_2087,N_1576);
and U4854 (N_4854,N_3960,N_1118);
xnor U4855 (N_4855,N_534,N_1440);
and U4856 (N_4856,N_3615,N_639);
and U4857 (N_4857,N_1263,N_2003);
nand U4858 (N_4858,N_546,N_800);
xnor U4859 (N_4859,N_726,N_1956);
or U4860 (N_4860,N_3445,N_3088);
xnor U4861 (N_4861,N_766,N_1275);
and U4862 (N_4862,N_1980,N_1921);
nand U4863 (N_4863,N_3847,N_3605);
nand U4864 (N_4864,N_3305,N_2334);
nand U4865 (N_4865,N_1651,N_3731);
nand U4866 (N_4866,N_1109,N_1653);
nand U4867 (N_4867,N_1818,N_3368);
nor U4868 (N_4868,N_1441,N_2532);
nand U4869 (N_4869,N_2359,N_3803);
nand U4870 (N_4870,N_714,N_2591);
and U4871 (N_4871,N_1681,N_3020);
xor U4872 (N_4872,N_3669,N_165);
xor U4873 (N_4873,N_1516,N_2166);
nor U4874 (N_4874,N_42,N_2417);
nand U4875 (N_4875,N_886,N_259);
nand U4876 (N_4876,N_1153,N_1372);
xor U4877 (N_4877,N_1730,N_3152);
xor U4878 (N_4878,N_964,N_276);
nor U4879 (N_4879,N_3030,N_3242);
or U4880 (N_4880,N_2657,N_40);
xor U4881 (N_4881,N_2852,N_2892);
xnor U4882 (N_4882,N_3082,N_1917);
nor U4883 (N_4883,N_778,N_1669);
nand U4884 (N_4884,N_255,N_2405);
xor U4885 (N_4885,N_2709,N_2246);
nor U4886 (N_4886,N_671,N_787);
xnor U4887 (N_4887,N_2636,N_3246);
nand U4888 (N_4888,N_1433,N_3863);
nand U4889 (N_4889,N_3772,N_291);
nor U4890 (N_4890,N_1447,N_795);
or U4891 (N_4891,N_3205,N_628);
and U4892 (N_4892,N_2499,N_1271);
nor U4893 (N_4893,N_2675,N_3567);
nor U4894 (N_4894,N_1314,N_846);
or U4895 (N_4895,N_3269,N_1301);
and U4896 (N_4896,N_3728,N_3209);
or U4897 (N_4897,N_1714,N_241);
or U4898 (N_4898,N_3167,N_1215);
and U4899 (N_4899,N_3695,N_2394);
and U4900 (N_4900,N_2015,N_962);
nor U4901 (N_4901,N_669,N_1415);
nor U4902 (N_4902,N_3398,N_2198);
or U4903 (N_4903,N_1425,N_1165);
xnor U4904 (N_4904,N_1718,N_793);
xor U4905 (N_4905,N_233,N_2720);
or U4906 (N_4906,N_729,N_3531);
or U4907 (N_4907,N_3128,N_389);
nand U4908 (N_4908,N_632,N_489);
and U4909 (N_4909,N_951,N_1224);
nand U4910 (N_4910,N_2456,N_1680);
xnor U4911 (N_4911,N_1620,N_2455);
xor U4912 (N_4912,N_322,N_176);
nand U4913 (N_4913,N_338,N_2552);
nand U4914 (N_4914,N_328,N_3511);
xnor U4915 (N_4915,N_1432,N_1363);
and U4916 (N_4916,N_3419,N_2640);
xor U4917 (N_4917,N_2523,N_2929);
xor U4918 (N_4918,N_1379,N_2497);
nand U4919 (N_4919,N_892,N_2381);
nor U4920 (N_4920,N_463,N_3575);
nor U4921 (N_4921,N_367,N_1408);
and U4922 (N_4922,N_2501,N_3620);
nand U4923 (N_4923,N_3901,N_775);
xor U4924 (N_4924,N_3975,N_3026);
nor U4925 (N_4925,N_2781,N_779);
xnor U4926 (N_4926,N_1830,N_2775);
nand U4927 (N_4927,N_603,N_2642);
or U4928 (N_4928,N_1332,N_2766);
nor U4929 (N_4929,N_2250,N_804);
nand U4930 (N_4930,N_3357,N_3697);
xnor U4931 (N_4931,N_443,N_3948);
or U4932 (N_4932,N_170,N_1533);
and U4933 (N_4933,N_2281,N_1626);
and U4934 (N_4934,N_791,N_1199);
xnor U4935 (N_4935,N_275,N_2251);
nor U4936 (N_4936,N_2447,N_1938);
xnor U4937 (N_4937,N_698,N_2349);
or U4938 (N_4938,N_487,N_1982);
xnor U4939 (N_4939,N_575,N_1853);
and U4940 (N_4940,N_3932,N_1502);
nand U4941 (N_4941,N_15,N_1200);
or U4942 (N_4942,N_1586,N_1990);
and U4943 (N_4943,N_552,N_3435);
xor U4944 (N_4944,N_530,N_2146);
xor U4945 (N_4945,N_716,N_537);
nand U4946 (N_4946,N_3146,N_347);
nor U4947 (N_4947,N_1745,N_812);
and U4948 (N_4948,N_3518,N_3619);
xnor U4949 (N_4949,N_543,N_2074);
or U4950 (N_4950,N_1878,N_1869);
and U4951 (N_4951,N_985,N_3797);
nand U4952 (N_4952,N_2396,N_2278);
xnor U4953 (N_4953,N_721,N_247);
nand U4954 (N_4954,N_2133,N_2961);
xor U4955 (N_4955,N_2855,N_2670);
nor U4956 (N_4956,N_3634,N_3186);
nor U4957 (N_4957,N_272,N_2823);
xnor U4958 (N_4958,N_14,N_1613);
or U4959 (N_4959,N_2100,N_19);
or U4960 (N_4960,N_3301,N_236);
xnor U4961 (N_4961,N_2574,N_3940);
nand U4962 (N_4962,N_1126,N_243);
or U4963 (N_4963,N_3233,N_3069);
xnor U4964 (N_4964,N_3573,N_2655);
nand U4965 (N_4965,N_3627,N_850);
xor U4966 (N_4966,N_1192,N_1471);
nor U4967 (N_4967,N_897,N_1560);
nand U4968 (N_4968,N_963,N_2873);
nand U4969 (N_4969,N_2109,N_3270);
or U4970 (N_4970,N_1454,N_435);
xnor U4971 (N_4971,N_2357,N_3108);
nor U4972 (N_4972,N_3172,N_2951);
nand U4973 (N_4973,N_483,N_2445);
xor U4974 (N_4974,N_1056,N_3672);
xor U4975 (N_4975,N_418,N_699);
nand U4976 (N_4976,N_3170,N_1529);
nand U4977 (N_4977,N_2743,N_3637);
or U4978 (N_4978,N_1551,N_561);
and U4979 (N_4979,N_1265,N_1923);
nor U4980 (N_4980,N_133,N_3303);
and U4981 (N_4981,N_823,N_1093);
nor U4982 (N_4982,N_3285,N_3412);
xor U4983 (N_4983,N_3798,N_3109);
or U4984 (N_4984,N_2638,N_82);
xor U4985 (N_4985,N_3098,N_2832);
xnor U4986 (N_4986,N_2883,N_258);
or U4987 (N_4987,N_1041,N_3827);
xor U4988 (N_4988,N_644,N_840);
nand U4989 (N_4989,N_3118,N_2373);
nand U4990 (N_4990,N_3474,N_230);
xnor U4991 (N_4991,N_3553,N_1855);
nand U4992 (N_4992,N_3624,N_3402);
xor U4993 (N_4993,N_1269,N_3174);
nor U4994 (N_4994,N_1327,N_1563);
or U4995 (N_4995,N_929,N_614);
nor U4996 (N_4996,N_3835,N_3374);
xnor U4997 (N_4997,N_1226,N_2188);
or U4998 (N_4998,N_969,N_1001);
nand U4999 (N_4999,N_2065,N_602);
or U5000 (N_5000,N_1623,N_1955);
and U5001 (N_5001,N_3063,N_114);
xor U5002 (N_5002,N_2749,N_419);
nand U5003 (N_5003,N_60,N_2646);
nor U5004 (N_5004,N_2965,N_3739);
nand U5005 (N_5005,N_1840,N_188);
xnor U5006 (N_5006,N_515,N_1350);
nor U5007 (N_5007,N_1094,N_2490);
and U5008 (N_5008,N_3818,N_1418);
or U5009 (N_5009,N_585,N_317);
nand U5010 (N_5010,N_235,N_158);
nand U5011 (N_5011,N_1808,N_1734);
or U5012 (N_5012,N_1517,N_3460);
nor U5013 (N_5013,N_941,N_1601);
nor U5014 (N_5014,N_153,N_2241);
xor U5015 (N_5015,N_2196,N_432);
and U5016 (N_5016,N_2684,N_3844);
and U5017 (N_5017,N_777,N_3541);
nor U5018 (N_5018,N_1450,N_3909);
nor U5019 (N_5019,N_559,N_2252);
nand U5020 (N_5020,N_3860,N_2882);
and U5021 (N_5021,N_2128,N_1274);
or U5022 (N_5022,N_2260,N_1453);
or U5023 (N_5023,N_1884,N_358);
nor U5024 (N_5024,N_2158,N_2622);
or U5025 (N_5025,N_1940,N_2502);
xor U5026 (N_5026,N_3083,N_2180);
and U5027 (N_5027,N_1384,N_2699);
xnor U5028 (N_5028,N_3418,N_704);
or U5029 (N_5029,N_2120,N_683);
nor U5030 (N_5030,N_2325,N_2092);
and U5031 (N_5031,N_212,N_905);
nand U5032 (N_5032,N_402,N_1488);
xor U5033 (N_5033,N_3031,N_826);
and U5034 (N_5034,N_1892,N_3543);
nand U5035 (N_5035,N_2849,N_1977);
or U5036 (N_5036,N_3277,N_2802);
nor U5037 (N_5037,N_932,N_3171);
and U5038 (N_5038,N_2452,N_1927);
and U5039 (N_5039,N_2797,N_2097);
or U5040 (N_5040,N_138,N_1684);
or U5041 (N_5041,N_67,N_378);
or U5042 (N_5042,N_1839,N_3984);
and U5043 (N_5043,N_1870,N_1091);
xor U5044 (N_5044,N_2412,N_2566);
nor U5045 (N_5045,N_1527,N_1313);
or U5046 (N_5046,N_2837,N_1863);
nand U5047 (N_5047,N_1895,N_1354);
nand U5048 (N_5048,N_3908,N_3636);
nor U5049 (N_5049,N_3943,N_2147);
and U5050 (N_5050,N_3750,N_1847);
and U5051 (N_5051,N_2347,N_2495);
nand U5052 (N_5052,N_1235,N_319);
and U5053 (N_5053,N_1127,N_3855);
or U5054 (N_5054,N_735,N_1185);
xnor U5055 (N_5055,N_659,N_2340);
or U5056 (N_5056,N_123,N_744);
nand U5057 (N_5057,N_2374,N_1242);
and U5058 (N_5058,N_1518,N_2101);
nor U5059 (N_5059,N_835,N_2463);
xor U5060 (N_5060,N_1545,N_1244);
nor U5061 (N_5061,N_3385,N_1097);
nor U5062 (N_5062,N_2226,N_1095);
nand U5063 (N_5063,N_3889,N_3089);
nand U5064 (N_5064,N_3899,N_1675);
nor U5065 (N_5065,N_1125,N_2547);
xnor U5066 (N_5066,N_410,N_1828);
and U5067 (N_5067,N_1088,N_954);
nand U5068 (N_5068,N_1548,N_774);
xor U5069 (N_5069,N_1106,N_136);
xnor U5070 (N_5070,N_1461,N_3609);
and U5071 (N_5071,N_2604,N_1770);
xnor U5072 (N_5072,N_2955,N_2978);
or U5073 (N_5073,N_1049,N_2314);
and U5074 (N_5074,N_3871,N_99);
or U5075 (N_5075,N_466,N_2994);
and U5076 (N_5076,N_3752,N_3149);
nor U5077 (N_5077,N_3574,N_3983);
xor U5078 (N_5078,N_801,N_539);
or U5079 (N_5079,N_3189,N_3422);
nor U5080 (N_5080,N_3949,N_3661);
or U5081 (N_5081,N_344,N_2024);
or U5082 (N_5082,N_2854,N_1258);
xnor U5083 (N_5083,N_2438,N_1970);
and U5084 (N_5084,N_709,N_2053);
nand U5085 (N_5085,N_1926,N_695);
xnor U5086 (N_5086,N_2019,N_2103);
nand U5087 (N_5087,N_1282,N_373);
and U5088 (N_5088,N_880,N_1152);
or U5089 (N_5089,N_1908,N_2435);
xor U5090 (N_5090,N_350,N_1736);
nand U5091 (N_5091,N_2826,N_1813);
xor U5092 (N_5092,N_2419,N_399);
and U5093 (N_5093,N_2535,N_3711);
or U5094 (N_5094,N_3200,N_2330);
or U5095 (N_5095,N_3566,N_1638);
nand U5096 (N_5096,N_2243,N_2156);
nand U5097 (N_5097,N_92,N_103);
and U5098 (N_5098,N_391,N_3178);
and U5099 (N_5099,N_3297,N_3134);
or U5100 (N_5100,N_455,N_512);
and U5101 (N_5101,N_2728,N_2135);
nand U5102 (N_5102,N_1716,N_3514);
xor U5103 (N_5103,N_3113,N_1538);
xor U5104 (N_5104,N_3453,N_1786);
nor U5105 (N_5105,N_3218,N_3344);
or U5106 (N_5106,N_2583,N_1366);
nand U5107 (N_5107,N_2765,N_1676);
and U5108 (N_5108,N_1744,N_3991);
nor U5109 (N_5109,N_2169,N_2032);
nand U5110 (N_5110,N_3593,N_1003);
and U5111 (N_5111,N_1362,N_384);
nand U5112 (N_5112,N_3214,N_3521);
and U5113 (N_5113,N_2516,N_889);
nor U5114 (N_5114,N_582,N_3147);
or U5115 (N_5115,N_1657,N_3650);
and U5116 (N_5116,N_1353,N_717);
or U5117 (N_5117,N_3401,N_3054);
xnor U5118 (N_5118,N_625,N_1539);
nand U5119 (N_5119,N_3891,N_2715);
and U5120 (N_5120,N_2915,N_2686);
and U5121 (N_5121,N_2301,N_2624);
and U5122 (N_5122,N_2172,N_163);
nand U5123 (N_5123,N_1952,N_3068);
nand U5124 (N_5124,N_2428,N_3250);
or U5125 (N_5125,N_3989,N_572);
nand U5126 (N_5126,N_556,N_2768);
and U5127 (N_5127,N_2219,N_3778);
or U5128 (N_5128,N_587,N_1357);
and U5129 (N_5129,N_448,N_839);
nor U5130 (N_5130,N_2737,N_2857);
or U5131 (N_5131,N_141,N_1254);
nand U5132 (N_5132,N_336,N_1446);
nand U5133 (N_5133,N_1427,N_3815);
nand U5134 (N_5134,N_551,N_3616);
xor U5135 (N_5135,N_3311,N_3969);
nand U5136 (N_5136,N_772,N_1059);
and U5137 (N_5137,N_1640,N_1211);
nand U5138 (N_5138,N_842,N_1549);
or U5139 (N_5139,N_902,N_1340);
and U5140 (N_5140,N_2814,N_1294);
xor U5141 (N_5141,N_1060,N_2388);
or U5142 (N_5142,N_2233,N_922);
xor U5143 (N_5143,N_1874,N_2323);
nor U5144 (N_5144,N_3604,N_2986);
nor U5145 (N_5145,N_2091,N_1639);
and U5146 (N_5146,N_2593,N_2880);
or U5147 (N_5147,N_2999,N_120);
nor U5148 (N_5148,N_2778,N_252);
or U5149 (N_5149,N_1399,N_2304);
or U5150 (N_5150,N_144,N_3709);
nand U5151 (N_5151,N_3164,N_1234);
xor U5152 (N_5152,N_52,N_2312);
nor U5153 (N_5153,N_1871,N_1702);
nor U5154 (N_5154,N_2450,N_961);
nand U5155 (N_5155,N_179,N_2674);
or U5156 (N_5156,N_1823,N_2028);
nor U5157 (N_5157,N_2174,N_2798);
nor U5158 (N_5158,N_3782,N_1325);
nor U5159 (N_5159,N_3539,N_0);
nand U5160 (N_5160,N_1046,N_607);
or U5161 (N_5161,N_3340,N_3125);
and U5162 (N_5162,N_2362,N_909);
or U5163 (N_5163,N_2733,N_2884);
nor U5164 (N_5164,N_2280,N_2107);
nand U5165 (N_5165,N_3092,N_3287);
or U5166 (N_5166,N_2950,N_1585);
or U5167 (N_5167,N_881,N_865);
and U5168 (N_5168,N_1778,N_492);
and U5169 (N_5169,N_3084,N_340);
nor U5170 (N_5170,N_3099,N_2390);
nand U5171 (N_5171,N_3480,N_1443);
and U5172 (N_5172,N_3489,N_1764);
xnor U5173 (N_5173,N_2080,N_3950);
xnor U5174 (N_5174,N_3466,N_958);
or U5175 (N_5175,N_2931,N_3409);
xnor U5176 (N_5176,N_1761,N_2906);
nand U5177 (N_5177,N_2788,N_3992);
nand U5178 (N_5178,N_869,N_3714);
nand U5179 (N_5179,N_125,N_226);
xor U5180 (N_5180,N_2928,N_2710);
nor U5181 (N_5181,N_1615,N_3414);
xnor U5182 (N_5182,N_1067,N_1773);
and U5183 (N_5183,N_3045,N_3973);
and U5184 (N_5184,N_1942,N_3848);
and U5185 (N_5185,N_507,N_142);
and U5186 (N_5186,N_2668,N_813);
and U5187 (N_5187,N_61,N_369);
nor U5188 (N_5188,N_547,N_611);
nand U5189 (N_5189,N_1760,N_3166);
nor U5190 (N_5190,N_1948,N_282);
xnor U5191 (N_5191,N_2565,N_1978);
or U5192 (N_5192,N_2425,N_223);
or U5193 (N_5193,N_1591,N_1534);
nor U5194 (N_5194,N_1365,N_108);
or U5195 (N_5195,N_719,N_3376);
and U5196 (N_5196,N_1996,N_411);
and U5197 (N_5197,N_2255,N_2207);
xor U5198 (N_5198,N_314,N_1083);
nor U5199 (N_5199,N_1246,N_2197);
or U5200 (N_5200,N_414,N_2095);
xor U5201 (N_5201,N_2286,N_442);
or U5202 (N_5202,N_2964,N_3725);
nand U5203 (N_5203,N_2460,N_2047);
xor U5204 (N_5204,N_2288,N_1656);
and U5205 (N_5205,N_2652,N_3);
nor U5206 (N_5206,N_2201,N_1812);
and U5207 (N_5207,N_2315,N_3407);
nand U5208 (N_5208,N_59,N_3217);
nor U5209 (N_5209,N_1793,N_3611);
and U5210 (N_5210,N_1262,N_1588);
nor U5211 (N_5211,N_3387,N_2503);
and U5212 (N_5212,N_2305,N_1320);
nand U5213 (N_5213,N_3319,N_1166);
nand U5214 (N_5214,N_2111,N_1928);
or U5215 (N_5215,N_228,N_260);
nand U5216 (N_5216,N_1498,N_3197);
nor U5217 (N_5217,N_1385,N_2161);
xnor U5218 (N_5218,N_462,N_1493);
xnor U5219 (N_5219,N_312,N_1606);
nor U5220 (N_5220,N_1319,N_2556);
nor U5221 (N_5221,N_80,N_420);
xnor U5222 (N_5222,N_400,N_1334);
xnor U5223 (N_5223,N_1774,N_769);
xnor U5224 (N_5224,N_86,N_3289);
xnor U5225 (N_5225,N_3055,N_768);
xnor U5226 (N_5226,N_302,N_3182);
and U5227 (N_5227,N_1704,N_2861);
and U5228 (N_5228,N_2508,N_1339);
nand U5229 (N_5229,N_1914,N_3837);
nor U5230 (N_5230,N_1178,N_526);
nor U5231 (N_5231,N_13,N_2254);
nor U5232 (N_5232,N_2212,N_1103);
or U5233 (N_5233,N_3536,N_2376);
xor U5234 (N_5234,N_2536,N_383);
nor U5235 (N_5235,N_403,N_3336);
and U5236 (N_5236,N_1336,N_268);
or U5237 (N_5237,N_452,N_1757);
xor U5238 (N_5238,N_3660,N_2086);
or U5239 (N_5239,N_3670,N_2462);
xor U5240 (N_5240,N_660,N_1101);
and U5241 (N_5241,N_2641,N_3047);
or U5242 (N_5242,N_3192,N_924);
or U5243 (N_5243,N_1501,N_3946);
and U5244 (N_5244,N_3103,N_3603);
and U5245 (N_5245,N_3351,N_2001);
and U5246 (N_5246,N_1413,N_2947);
or U5247 (N_5247,N_3048,N_155);
and U5248 (N_5248,N_2954,N_2672);
or U5249 (N_5249,N_2119,N_199);
or U5250 (N_5250,N_76,N_98);
or U5251 (N_5251,N_2230,N_3741);
and U5252 (N_5252,N_1631,N_3990);
or U5253 (N_5253,N_433,N_2836);
nor U5254 (N_5254,N_1963,N_1260);
and U5255 (N_5255,N_3864,N_3469);
xnor U5256 (N_5256,N_524,N_3599);
nor U5257 (N_5257,N_48,N_1197);
nor U5258 (N_5258,N_3119,N_2632);
nand U5259 (N_5259,N_2921,N_1685);
or U5260 (N_5260,N_2541,N_3261);
and U5261 (N_5261,N_875,N_3594);
or U5262 (N_5262,N_1156,N_3762);
and U5263 (N_5263,N_1157,N_3151);
nor U5264 (N_5264,N_1765,N_1559);
and U5265 (N_5265,N_3413,N_3332);
xor U5266 (N_5266,N_3779,N_2512);
xor U5267 (N_5267,N_485,N_1176);
nor U5268 (N_5268,N_1590,N_856);
or U5269 (N_5269,N_3621,N_3003);
xnor U5270 (N_5270,N_1690,N_656);
nand U5271 (N_5271,N_1397,N_1967);
nand U5272 (N_5272,N_3439,N_3907);
or U5273 (N_5273,N_2105,N_1019);
nand U5274 (N_5274,N_2009,N_3286);
and U5275 (N_5275,N_70,N_1846);
nand U5276 (N_5276,N_3036,N_650);
nor U5277 (N_5277,N_2153,N_183);
nand U5278 (N_5278,N_3219,N_2673);
nor U5279 (N_5279,N_3925,N_3572);
and U5280 (N_5280,N_423,N_209);
nor U5281 (N_5281,N_2695,N_758);
nor U5282 (N_5282,N_1307,N_3517);
or U5283 (N_5283,N_3361,N_3046);
nor U5284 (N_5284,N_2182,N_3161);
nor U5285 (N_5285,N_3227,N_3131);
and U5286 (N_5286,N_3635,N_749);
nand U5287 (N_5287,N_345,N_244);
and U5288 (N_5288,N_2303,N_169);
or U5289 (N_5289,N_1139,N_1481);
nand U5290 (N_5290,N_1251,N_3491);
nand U5291 (N_5291,N_1916,N_1396);
nand U5292 (N_5292,N_3173,N_618);
and U5293 (N_5293,N_1889,N_2123);
xor U5294 (N_5294,N_1063,N_3993);
xnor U5295 (N_5295,N_1694,N_3898);
and U5296 (N_5296,N_3329,N_3791);
nand U5297 (N_5297,N_2544,N_1624);
nor U5298 (N_5298,N_2602,N_3391);
or U5299 (N_5299,N_2294,N_2308);
or U5300 (N_5300,N_2027,N_899);
xor U5301 (N_5301,N_2881,N_2525);
nand U5302 (N_5302,N_1854,N_619);
nor U5303 (N_5303,N_3239,N_3433);
and U5304 (N_5304,N_1113,N_803);
nor U5305 (N_5305,N_1068,N_581);
nand U5306 (N_5306,N_2665,N_430);
nand U5307 (N_5307,N_2225,N_728);
and U5308 (N_5308,N_1312,N_2606);
or U5309 (N_5309,N_1431,N_2429);
xor U5310 (N_5310,N_3339,N_686);
or U5311 (N_5311,N_1043,N_2295);
nand U5312 (N_5312,N_2433,N_2550);
and U5313 (N_5313,N_873,N_3203);
nor U5314 (N_5314,N_377,N_3758);
and U5315 (N_5315,N_1861,N_361);
nor U5316 (N_5316,N_1553,N_755);
nor U5317 (N_5317,N_982,N_580);
nand U5318 (N_5318,N_3265,N_2154);
nor U5319 (N_5319,N_3982,N_1664);
or U5320 (N_5320,N_979,N_1667);
nor U5321 (N_5321,N_2187,N_1749);
nor U5322 (N_5322,N_3458,N_3123);
xor U5323 (N_5323,N_3913,N_3928);
and U5324 (N_5324,N_1474,N_3628);
xnor U5325 (N_5325,N_3231,N_944);
nor U5326 (N_5326,N_1168,N_1098);
nand U5327 (N_5327,N_1597,N_3516);
xnor U5328 (N_5328,N_999,N_1748);
nor U5329 (N_5329,N_2767,N_1815);
or U5330 (N_5330,N_3838,N_3389);
nor U5331 (N_5331,N_1991,N_522);
and U5332 (N_5332,N_1072,N_514);
nor U5333 (N_5333,N_3941,N_2939);
or U5334 (N_5334,N_2568,N_679);
xnor U5335 (N_5335,N_3823,N_245);
nor U5336 (N_5336,N_652,N_1025);
or U5337 (N_5337,N_327,N_3399);
or U5338 (N_5338,N_3034,N_3162);
xor U5339 (N_5339,N_2189,N_3211);
nand U5340 (N_5340,N_1250,N_156);
nor U5341 (N_5341,N_2601,N_2958);
nor U5342 (N_5342,N_2555,N_3842);
and U5343 (N_5343,N_3703,N_2448);
and U5344 (N_5344,N_1627,N_1145);
xnor U5345 (N_5345,N_1018,N_1739);
nand U5346 (N_5346,N_3878,N_785);
and U5347 (N_5347,N_2997,N_1090);
and U5348 (N_5348,N_2046,N_1753);
or U5349 (N_5349,N_762,N_1463);
nor U5350 (N_5350,N_890,N_3425);
xor U5351 (N_5351,N_3367,N_1984);
and U5352 (N_5352,N_732,N_3185);
nand U5353 (N_5353,N_2531,N_83);
xor U5354 (N_5354,N_2005,N_1535);
nor U5355 (N_5355,N_3106,N_852);
and U5356 (N_5356,N_2993,N_3472);
nand U5357 (N_5357,N_3664,N_2584);
nor U5358 (N_5358,N_1510,N_3195);
nand U5359 (N_5359,N_3029,N_2477);
xor U5360 (N_5360,N_3245,N_3032);
and U5361 (N_5361,N_2790,N_3919);
nor U5362 (N_5362,N_810,N_2379);
xor U5363 (N_5363,N_1747,N_3061);
nand U5364 (N_5364,N_2275,N_3865);
nor U5365 (N_5365,N_692,N_3562);
or U5366 (N_5366,N_3350,N_3455);
nor U5367 (N_5367,N_1061,N_2432);
nand U5368 (N_5368,N_966,N_1117);
or U5369 (N_5369,N_1678,N_398);
or U5370 (N_5370,N_2989,N_3137);
nand U5371 (N_5371,N_3326,N_113);
nor U5372 (N_5372,N_177,N_285);
nor U5373 (N_5373,N_3834,N_1612);
or U5374 (N_5374,N_2346,N_2132);
nor U5375 (N_5375,N_2513,N_96);
xor U5376 (N_5376,N_2043,N_1499);
nor U5377 (N_5377,N_2139,N_2178);
nor U5378 (N_5378,N_1466,N_3346);
nand U5379 (N_5379,N_1607,N_2072);
nand U5380 (N_5380,N_2795,N_2727);
nand U5381 (N_5381,N_2116,N_2054);
xnor U5382 (N_5382,N_2530,N_3882);
or U5383 (N_5383,N_1652,N_2413);
and U5384 (N_5384,N_3072,N_833);
or U5385 (N_5385,N_2850,N_1522);
or U5386 (N_5386,N_2181,N_2507);
xor U5387 (N_5387,N_2967,N_1333);
nor U5388 (N_5388,N_2590,N_1920);
nand U5389 (N_5389,N_2037,N_215);
and U5390 (N_5390,N_1506,N_1369);
xor U5391 (N_5391,N_2273,N_3155);
xor U5392 (N_5392,N_1796,N_55);
nand U5393 (N_5393,N_496,N_2193);
and U5394 (N_5394,N_2465,N_3322);
nand U5395 (N_5395,N_1266,N_917);
or U5396 (N_5396,N_752,N_3190);
or U5397 (N_5397,N_2378,N_1321);
xnor U5398 (N_5398,N_532,N_2667);
xor U5399 (N_5399,N_1790,N_2745);
and U5400 (N_5400,N_1581,N_2518);
and U5401 (N_5401,N_1107,N_1733);
and U5402 (N_5402,N_3143,N_3979);
nand U5403 (N_5403,N_1547,N_862);
nor U5404 (N_5404,N_3440,N_1293);
nand U5405 (N_5405,N_947,N_796);
nor U5406 (N_5406,N_883,N_2726);
nand U5407 (N_5407,N_2177,N_854);
and U5408 (N_5408,N_705,N_2474);
xor U5409 (N_5409,N_2364,N_3937);
nand U5410 (N_5410,N_919,N_1167);
nor U5411 (N_5411,N_1071,N_28);
and U5412 (N_5412,N_3904,N_712);
nand U5413 (N_5413,N_107,N_1006);
or U5414 (N_5414,N_2524,N_1566);
nor U5415 (N_5415,N_2811,N_269);
or U5416 (N_5416,N_3310,N_3978);
or U5417 (N_5417,N_3394,N_2002);
xor U5418 (N_5418,N_2298,N_3215);
and U5419 (N_5419,N_3229,N_3300);
nand U5420 (N_5420,N_3392,N_3304);
nand U5421 (N_5421,N_1625,N_494);
nand U5422 (N_5422,N_2468,N_888);
or U5423 (N_5423,N_2847,N_1378);
and U5424 (N_5424,N_2279,N_1009);
and U5425 (N_5425,N_1075,N_3526);
and U5426 (N_5426,N_1579,N_8);
nand U5427 (N_5427,N_181,N_3875);
or U5428 (N_5428,N_1080,N_2350);
nor U5429 (N_5429,N_3328,N_518);
and U5430 (N_5430,N_615,N_2113);
and U5431 (N_5431,N_2520,N_1005);
nor U5432 (N_5432,N_3104,N_1569);
and U5433 (N_5433,N_2995,N_1561);
nand U5434 (N_5434,N_617,N_421);
xor U5435 (N_5435,N_903,N_1992);
xor U5436 (N_5436,N_3373,N_1351);
nor U5437 (N_5437,N_2102,N_674);
xnor U5438 (N_5438,N_3995,N_2440);
nand U5439 (N_5439,N_2773,N_633);
and U5440 (N_5440,N_1637,N_1691);
and U5441 (N_5441,N_1052,N_1328);
and U5442 (N_5442,N_2942,N_493);
nor U5443 (N_5443,N_66,N_3502);
xor U5444 (N_5444,N_2125,N_2336);
xor U5445 (N_5445,N_2687,N_1841);
nand U5446 (N_5446,N_3770,N_2239);
xor U5447 (N_5447,N_2395,N_1856);
nand U5448 (N_5448,N_1654,N_109);
and U5449 (N_5449,N_940,N_2500);
xor U5450 (N_5450,N_3295,N_2262);
or U5451 (N_5451,N_453,N_2660);
or U5452 (N_5452,N_371,N_503);
and U5453 (N_5453,N_687,N_1143);
or U5454 (N_5454,N_2774,N_2098);
or U5455 (N_5455,N_211,N_2256);
nor U5456 (N_5456,N_2894,N_2287);
xnor U5457 (N_5457,N_90,N_3740);
nor U5458 (N_5458,N_3704,N_38);
xor U5459 (N_5459,N_53,N_819);
nor U5460 (N_5460,N_1252,N_784);
nor U5461 (N_5461,N_753,N_1011);
nand U5462 (N_5462,N_2528,N_1630);
xnor U5463 (N_5463,N_1822,N_1324);
xor U5464 (N_5464,N_1300,N_3145);
xor U5465 (N_5465,N_637,N_256);
and U5466 (N_5466,N_662,N_2129);
xor U5467 (N_5467,N_47,N_1949);
nand U5468 (N_5468,N_2242,N_2527);
nor U5469 (N_5469,N_895,N_1814);
nor U5470 (N_5470,N_289,N_3014);
and U5471 (N_5471,N_2840,N_101);
nand U5472 (N_5472,N_538,N_2366);
xor U5473 (N_5473,N_467,N_1040);
xnor U5474 (N_5474,N_667,N_2427);
xnor U5475 (N_5475,N_1616,N_3468);
nor U5476 (N_5476,N_7,N_629);
xor U5477 (N_5477,N_85,N_1477);
and U5478 (N_5478,N_81,N_703);
or U5479 (N_5479,N_3652,N_1959);
or U5480 (N_5480,N_3140,N_3315);
xor U5481 (N_5481,N_202,N_219);
xor U5482 (N_5482,N_1834,N_1811);
and U5483 (N_5483,N_1383,N_1449);
nor U5484 (N_5484,N_2041,N_2860);
nand U5485 (N_5485,N_3330,N_352);
and U5486 (N_5486,N_3583,N_2088);
nor U5487 (N_5487,N_2920,N_2722);
xnor U5488 (N_5488,N_324,N_3483);
nor U5489 (N_5489,N_1715,N_1542);
nor U5490 (N_5490,N_58,N_3785);
or U5491 (N_5491,N_3900,N_3122);
xnor U5492 (N_5492,N_2371,N_3259);
xor U5493 (N_5493,N_3886,N_3896);
and U5494 (N_5494,N_550,N_3463);
and U5495 (N_5495,N_3027,N_1789);
nor U5496 (N_5496,N_3062,N_3381);
and U5497 (N_5497,N_2051,N_3369);
nand U5498 (N_5498,N_1520,N_2639);
and U5499 (N_5499,N_2149,N_1128);
or U5500 (N_5500,N_1661,N_2571);
xor U5501 (N_5501,N_2437,N_348);
or U5502 (N_5502,N_2663,N_3794);
and U5503 (N_5503,N_2058,N_1767);
and U5504 (N_5504,N_3264,N_1735);
or U5505 (N_5505,N_2714,N_1456);
nor U5506 (N_5506,N_566,N_1706);
nand U5507 (N_5507,N_460,N_1859);
xnor U5508 (N_5508,N_3706,N_3442);
nand U5509 (N_5509,N_651,N_2828);
or U5510 (N_5510,N_2442,N_3266);
nand U5511 (N_5511,N_79,N_2548);
and U5512 (N_5512,N_1134,N_770);
nand U5513 (N_5513,N_3005,N_2446);
xnor U5514 (N_5514,N_601,N_2237);
nand U5515 (N_5515,N_1259,N_293);
nand U5516 (N_5516,N_3698,N_3437);
nand U5517 (N_5517,N_2569,N_117);
nand U5518 (N_5518,N_780,N_498);
xor U5519 (N_5519,N_3320,N_1965);
xnor U5520 (N_5520,N_3087,N_240);
xor U5521 (N_5521,N_458,N_1589);
nor U5522 (N_5522,N_1190,N_1972);
or U5523 (N_5523,N_205,N_1712);
or U5524 (N_5524,N_3202,N_663);
or U5525 (N_5525,N_3049,N_606);
nand U5526 (N_5526,N_2560,N_2918);
and U5527 (N_5527,N_2240,N_1022);
or U5528 (N_5528,N_697,N_3945);
and U5529 (N_5529,N_1649,N_2271);
or U5530 (N_5530,N_2510,N_622);
nor U5531 (N_5531,N_2963,N_1934);
and U5532 (N_5532,N_2820,N_1337);
nor U5533 (N_5533,N_200,N_2785);
nand U5534 (N_5534,N_1002,N_2763);
or U5535 (N_5535,N_1051,N_2563);
nand U5536 (N_5536,N_2704,N_3230);
and U5537 (N_5537,N_172,N_3028);
and U5538 (N_5538,N_3481,N_1894);
or U5539 (N_5539,N_740,N_29);
nor U5540 (N_5540,N_63,N_653);
or U5541 (N_5541,N_1769,N_3681);
xor U5542 (N_5542,N_1457,N_2090);
nand U5543 (N_5543,N_1087,N_2529);
nor U5544 (N_5544,N_193,N_3774);
and U5545 (N_5545,N_2938,N_3890);
and U5546 (N_5546,N_743,N_1193);
nor U5547 (N_5547,N_634,N_1913);
nor U5548 (N_5548,N_3520,N_1129);
or U5549 (N_5549,N_1186,N_1732);
nor U5550 (N_5550,N_1567,N_1803);
nand U5551 (N_5551,N_1356,N_429);
or U5552 (N_5552,N_1144,N_1592);
nor U5553 (N_5553,N_3206,N_68);
nor U5554 (N_5554,N_3283,N_2150);
xor U5555 (N_5555,N_3388,N_1596);
nor U5556 (N_5556,N_855,N_3766);
nor U5557 (N_5557,N_2561,N_2956);
nor U5558 (N_5558,N_1406,N_3065);
nand U5559 (N_5559,N_148,N_24);
or U5560 (N_5560,N_3378,N_3748);
and U5561 (N_5561,N_2926,N_197);
nor U5562 (N_5562,N_3411,N_2036);
nand U5563 (N_5563,N_1158,N_2332);
nor U5564 (N_5564,N_390,N_381);
nor U5565 (N_5565,N_2742,N_2740);
and U5566 (N_5566,N_182,N_2694);
nand U5567 (N_5567,N_1030,N_844);
xnor U5568 (N_5568,N_2572,N_1673);
and U5569 (N_5569,N_3754,N_1171);
or U5570 (N_5570,N_161,N_30);
and U5571 (N_5571,N_2441,N_477);
xnor U5572 (N_5572,N_545,N_3366);
or U5573 (N_5573,N_1042,N_925);
nand U5574 (N_5574,N_1907,N_3654);
nor U5575 (N_5575,N_891,N_1931);
nand U5576 (N_5576,N_1893,N_1610);
or U5577 (N_5577,N_2824,N_3856);
and U5578 (N_5578,N_3298,N_3406);
nand U5579 (N_5579,N_1392,N_1688);
and U5580 (N_5580,N_1154,N_3042);
and U5581 (N_5581,N_262,N_1187);
xnor U5582 (N_5582,N_2163,N_3262);
xor U5583 (N_5583,N_2867,N_3156);
and U5584 (N_5584,N_2794,N_945);
or U5585 (N_5585,N_783,N_3537);
nor U5586 (N_5586,N_208,N_734);
xor U5587 (N_5587,N_2949,N_1562);
or U5588 (N_5588,N_3970,N_3079);
nor U5589 (N_5589,N_187,N_3393);
or U5590 (N_5590,N_3416,N_2209);
and U5591 (N_5591,N_2494,N_221);
xnor U5592 (N_5592,N_3362,N_3826);
nand U5593 (N_5593,N_2030,N_1078);
or U5594 (N_5594,N_2621,N_3767);
nand U5595 (N_5595,N_3325,N_3379);
and U5596 (N_5596,N_1358,N_3111);
and U5597 (N_5597,N_2409,N_3710);
and U5598 (N_5598,N_2724,N_3078);
nor U5599 (N_5599,N_516,N_3341);
nand U5600 (N_5600,N_2489,N_3996);
or U5601 (N_5601,N_3912,N_422);
nor U5602 (N_5602,N_3809,N_2777);
nand U5603 (N_5603,N_1065,N_132);
or U5604 (N_5604,N_36,N_2769);
and U5605 (N_5605,N_824,N_2382);
or U5606 (N_5606,N_2426,N_1240);
or U5607 (N_5607,N_1609,N_1298);
and U5608 (N_5608,N_3142,N_149);
and U5609 (N_5609,N_3642,N_675);
or U5610 (N_5610,N_1958,N_3241);
nand U5611 (N_5611,N_337,N_722);
nand U5612 (N_5612,N_1824,N_316);
nor U5613 (N_5613,N_3384,N_3060);
nor U5614 (N_5614,N_731,N_761);
and U5615 (N_5615,N_2351,N_105);
nand U5616 (N_5616,N_2731,N_1998);
xor U5617 (N_5617,N_2821,N_565);
and U5618 (N_5618,N_2812,N_2070);
xnor U5619 (N_5619,N_3601,N_3841);
xor U5620 (N_5620,N_3429,N_3671);
nor U5621 (N_5621,N_1741,N_2414);
and U5622 (N_5622,N_1302,N_2907);
xor U5623 (N_5623,N_1476,N_3591);
or U5624 (N_5624,N_2141,N_996);
and U5625 (N_5625,N_3997,N_1851);
nand U5626 (N_5626,N_1696,N_2339);
nand U5627 (N_5627,N_3585,N_1016);
nor U5628 (N_5628,N_2265,N_3258);
nand U5629 (N_5629,N_3747,N_2459);
xnor U5630 (N_5630,N_1766,N_257);
xor U5631 (N_5631,N_3833,N_2404);
nor U5632 (N_5632,N_3019,N_3052);
or U5633 (N_5633,N_1599,N_1195);
xor U5634 (N_5634,N_2700,N_3484);
xor U5635 (N_5635,N_2948,N_3312);
xnor U5636 (N_5636,N_1445,N_1021);
or U5637 (N_5637,N_3965,N_472);
and U5638 (N_5638,N_984,N_3581);
xnor U5639 (N_5639,N_1359,N_1470);
xor U5640 (N_5640,N_3528,N_425);
nand U5641 (N_5641,N_2789,N_790);
xor U5642 (N_5642,N_1703,N_2136);
xnor U5643 (N_5643,N_1465,N_1810);
and U5644 (N_5644,N_3586,N_931);
nor U5645 (N_5645,N_1944,N_2603);
nor U5646 (N_5646,N_3107,N_3159);
or U5647 (N_5647,N_3313,N_2779);
nor U5648 (N_5648,N_3465,N_1267);
and U5649 (N_5649,N_6,N_3877);
nand U5650 (N_5650,N_1887,N_1389);
and U5651 (N_5651,N_3859,N_3408);
or U5652 (N_5652,N_1683,N_2492);
xor U5653 (N_5653,N_1288,N_2730);
or U5654 (N_5654,N_1204,N_1057);
or U5655 (N_5655,N_3436,N_3482);
and U5656 (N_5656,N_1896,N_900);
nor U5657 (N_5657,N_3569,N_558);
or U5658 (N_5658,N_725,N_3225);
and U5659 (N_5659,N_3022,N_3158);
nor U5660 (N_5660,N_2480,N_2173);
nor U5661 (N_5661,N_3035,N_2124);
nor U5662 (N_5662,N_3868,N_2059);
xnor U5663 (N_5663,N_1738,N_1904);
nor U5664 (N_5664,N_1918,N_3555);
or U5665 (N_5665,N_1459,N_2943);
nor U5666 (N_5666,N_1525,N_69);
or U5667 (N_5667,N_2843,N_3395);
and U5668 (N_5668,N_3443,N_1112);
or U5669 (N_5669,N_3275,N_1552);
xnor U5670 (N_5670,N_3682,N_564);
nand U5671 (N_5671,N_3853,N_3102);
and U5672 (N_5672,N_1852,N_764);
or U5673 (N_5673,N_1439,N_3375);
and U5674 (N_5674,N_1888,N_3623);
nor U5675 (N_5675,N_1276,N_2195);
xnor U5676 (N_5676,N_820,N_950);
xnor U5677 (N_5677,N_1216,N_1330);
nor U5678 (N_5678,N_1318,N_1881);
and U5679 (N_5679,N_2551,N_2904);
nor U5680 (N_5680,N_3462,N_1292);
xnor U5681 (N_5681,N_2276,N_1343);
xor U5682 (N_5682,N_741,N_2134);
and U5683 (N_5683,N_2739,N_2384);
nor U5684 (N_5684,N_597,N_2732);
nand U5685 (N_5685,N_3760,N_3009);
xor U5686 (N_5686,N_1084,N_1693);
nor U5687 (N_5687,N_3193,N_3354);
xnor U5688 (N_5688,N_1311,N_1831);
xnor U5689 (N_5689,N_1237,N_299);
nor U5690 (N_5690,N_691,N_3716);
and U5691 (N_5691,N_1987,N_306);
nand U5692 (N_5692,N_500,N_1);
nand U5693 (N_5693,N_2975,N_1508);
nand U5694 (N_5694,N_2338,N_3115);
or U5695 (N_5695,N_88,N_1305);
nand U5696 (N_5696,N_3618,N_3271);
nor U5697 (N_5697,N_3812,N_3737);
and U5698 (N_5698,N_661,N_1451);
or U5699 (N_5699,N_3101,N_1066);
nor U5700 (N_5700,N_1700,N_16);
nand U5701 (N_5701,N_3918,N_1707);
nor U5702 (N_5702,N_1670,N_3977);
and U5703 (N_5703,N_393,N_3177);
xor U5704 (N_5704,N_2998,N_894);
xor U5705 (N_5705,N_2842,N_1111);
nor U5706 (N_5706,N_2343,N_1644);
and U5707 (N_5707,N_2168,N_3112);
nor U5708 (N_5708,N_2874,N_3347);
or U5709 (N_5709,N_3771,N_860);
nand U5710 (N_5710,N_1405,N_1388);
nor U5711 (N_5711,N_3674,N_3769);
nand U5712 (N_5712,N_579,N_901);
nand U5713 (N_5713,N_3255,N_3495);
nor U5714 (N_5714,N_129,N_1721);
nand U5715 (N_5715,N_3638,N_3438);
xor U5716 (N_5716,N_3094,N_3080);
nand U5717 (N_5717,N_2838,N_427);
and U5718 (N_5718,N_424,N_1364);
nor U5719 (N_5719,N_484,N_1062);
xor U5720 (N_5720,N_191,N_346);
and U5721 (N_5721,N_360,N_2719);
and U5722 (N_5722,N_2554,N_2713);
or U5723 (N_5723,N_3696,N_1646);
and U5724 (N_5724,N_3228,N_131);
xnor U5725 (N_5725,N_1645,N_2021);
xor U5726 (N_5726,N_3017,N_1754);
nand U5727 (N_5727,N_1792,N_2723);
nor U5728 (N_5728,N_928,N_1346);
nor U5729 (N_5729,N_1541,N_590);
and U5730 (N_5730,N_2859,N_1174);
nor U5731 (N_5731,N_2677,N_2335);
nand U5732 (N_5732,N_3795,N_2342);
nor U5733 (N_5733,N_2470,N_960);
nand U5734 (N_5734,N_646,N_248);
or U5735 (N_5735,N_121,N_2127);
nor U5736 (N_5736,N_811,N_2741);
nand U5737 (N_5737,N_3956,N_1490);
xnor U5738 (N_5738,N_911,N_2324);
nand U5739 (N_5739,N_334,N_3867);
nand U5740 (N_5740,N_3707,N_2383);
xnor U5741 (N_5741,N_809,N_2545);
xnor U5742 (N_5742,N_2293,N_185);
nor U5743 (N_5743,N_673,N_643);
nor U5744 (N_5744,N_454,N_3371);
and U5745 (N_5745,N_3059,N_1069);
nor U5746 (N_5746,N_1280,N_968);
or U5747 (N_5747,N_3821,N_2326);
nand U5748 (N_5748,N_1081,N_838);
nand U5749 (N_5749,N_685,N_623);
and U5750 (N_5750,N_1577,N_3641);
nand U5751 (N_5751,N_2977,N_2806);
xor U5752 (N_5752,N_2234,N_957);
nand U5753 (N_5753,N_3846,N_2996);
nand U5754 (N_5754,N_2858,N_1473);
xor U5755 (N_5755,N_1323,N_1020);
nor U5756 (N_5756,N_2044,N_1788);
xor U5757 (N_5757,N_2818,N_74);
and U5758 (N_5758,N_2718,N_3915);
and U5759 (N_5759,N_3345,N_2692);
nand U5760 (N_5760,N_387,N_2992);
or U5761 (N_5761,N_210,N_3542);
xor U5762 (N_5762,N_2179,N_3688);
or U5763 (N_5763,N_3887,N_3662);
nor U5764 (N_5764,N_1303,N_1583);
xnor U5765 (N_5765,N_2813,N_2029);
xor U5766 (N_5766,N_2876,N_150);
xor U5767 (N_5767,N_1985,N_3077);
or U5768 (N_5768,N_2322,N_1124);
or U5769 (N_5769,N_1791,N_2609);
nand U5770 (N_5770,N_1523,N_2062);
and U5771 (N_5771,N_2042,N_2386);
xnor U5772 (N_5772,N_3568,N_1731);
xor U5773 (N_5773,N_1845,N_598);
and U5774 (N_5774,N_408,N_3580);
xor U5775 (N_5775,N_2522,N_3176);
nand U5776 (N_5776,N_3168,N_3930);
and U5777 (N_5777,N_3719,N_1253);
and U5778 (N_5778,N_1196,N_987);
nor U5779 (N_5779,N_2817,N_436);
or U5780 (N_5780,N_2232,N_2538);
nor U5781 (N_5781,N_273,N_2966);
or U5782 (N_5782,N_441,N_2600);
nor U5783 (N_5783,N_2791,N_3817);
xnor U5784 (N_5784,N_100,N_2157);
nor U5785 (N_5785,N_2834,N_1400);
nand U5786 (N_5786,N_3247,N_1820);
nand U5787 (N_5787,N_3777,N_3957);
and U5788 (N_5788,N_3556,N_1285);
and U5789 (N_5789,N_1322,N_2372);
and U5790 (N_5790,N_2711,N_3743);
nor U5791 (N_5791,N_362,N_857);
xor U5792 (N_5792,N_828,N_624);
and U5793 (N_5793,N_677,N_2509);
or U5794 (N_5794,N_3819,N_2183);
or U5795 (N_5795,N_517,N_94);
or U5796 (N_5796,N_1241,N_1179);
xor U5797 (N_5797,N_1882,N_2662);
and U5798 (N_5798,N_2049,N_2236);
nand U5799 (N_5799,N_3386,N_1442);
xor U5800 (N_5800,N_1600,N_1034);
xnor U5801 (N_5801,N_2387,N_3355);
nand U5802 (N_5802,N_2848,N_2514);
xor U5803 (N_5803,N_3527,N_2067);
nor U5804 (N_5804,N_3903,N_279);
nand U5805 (N_5805,N_2803,N_2176);
nand U5806 (N_5806,N_2160,N_3807);
or U5807 (N_5807,N_2934,N_3334);
xor U5808 (N_5808,N_3732,N_1256);
nor U5809 (N_5809,N_2744,N_2248);
nor U5810 (N_5810,N_394,N_3802);
and U5811 (N_5811,N_2266,N_965);
nand U5812 (N_5812,N_3831,N_3420);
xnor U5813 (N_5813,N_3916,N_301);
xnor U5814 (N_5814,N_3372,N_3587);
xnor U5815 (N_5815,N_3007,N_115);
and U5816 (N_5816,N_3784,N_1779);
nand U5817 (N_5817,N_638,N_1727);
nand U5818 (N_5818,N_3487,N_684);
and U5819 (N_5819,N_271,N_1821);
nor U5820 (N_5820,N_168,N_2829);
or U5821 (N_5821,N_2747,N_3073);
nor U5822 (N_5822,N_1155,N_217);
or U5823 (N_5823,N_3963,N_2475);
and U5824 (N_5824,N_3828,N_3342);
and U5825 (N_5825,N_1130,N_84);
and U5826 (N_5826,N_3070,N_2944);
or U5827 (N_5827,N_1595,N_1212);
or U5828 (N_5828,N_1032,N_898);
nor U5829 (N_5829,N_2430,N_2479);
and U5830 (N_5830,N_3888,N_2810);
xor U5831 (N_5831,N_1017,N_1074);
and U5832 (N_5832,N_655,N_2680);
nand U5833 (N_5833,N_2573,N_3056);
and U5834 (N_5834,N_974,N_3790);
and U5835 (N_5835,N_1819,N_3477);
and U5836 (N_5836,N_3734,N_3424);
xor U5837 (N_5837,N_1838,N_2570);
nor U5838 (N_5838,N_1879,N_3986);
nor U5839 (N_5839,N_923,N_2851);
nor U5840 (N_5840,N_3066,N_1759);
nand U5841 (N_5841,N_586,N_239);
and U5842 (N_5842,N_1247,N_636);
or U5843 (N_5843,N_3610,N_292);
xnor U5844 (N_5844,N_604,N_2581);
xor U5845 (N_5845,N_3579,N_3656);
nor U5846 (N_5846,N_1937,N_1306);
or U5847 (N_5847,N_409,N_3290);
nor U5848 (N_5848,N_3955,N_3224);
nand U5849 (N_5849,N_3733,N_1999);
nand U5850 (N_5850,N_2588,N_2004);
nand U5851 (N_5851,N_3951,N_2411);
nor U5852 (N_5852,N_832,N_3430);
xor U5853 (N_5853,N_2151,N_3499);
and U5854 (N_5854,N_1495,N_2493);
nand U5855 (N_5855,N_3832,N_2682);
nor U5856 (N_5856,N_2557,N_3694);
or U5857 (N_5857,N_1929,N_2988);
or U5858 (N_5858,N_1430,N_2678);
xor U5859 (N_5859,N_449,N_654);
nor U5860 (N_5860,N_733,N_1055);
nor U5861 (N_5861,N_1013,N_1201);
xnor U5862 (N_5862,N_2620,N_2878);
or U5863 (N_5863,N_3421,N_2979);
and U5864 (N_5864,N_1503,N_1141);
or U5865 (N_5865,N_3446,N_933);
or U5866 (N_5866,N_1555,N_1206);
and U5867 (N_5867,N_2933,N_872);
xor U5868 (N_5868,N_3130,N_3655);
nor U5869 (N_5869,N_2705,N_355);
nor U5870 (N_5870,N_2659,N_3761);
and U5871 (N_5871,N_2238,N_2408);
xnor U5872 (N_5872,N_2712,N_1858);
nor U5873 (N_5873,N_1722,N_2048);
xor U5874 (N_5874,N_1505,N_3183);
nand U5875 (N_5875,N_3400,N_130);
and U5876 (N_5876,N_2629,N_147);
nand U5877 (N_5877,N_118,N_2786);
xor U5878 (N_5878,N_1048,N_2927);
nor U5879 (N_5879,N_2962,N_3175);
or U5880 (N_5880,N_3370,N_2082);
xor U5881 (N_5881,N_868,N_2671);
or U5882 (N_5882,N_3196,N_3428);
nand U5883 (N_5883,N_3359,N_3561);
and U5884 (N_5884,N_2263,N_1270);
and U5885 (N_5885,N_978,N_3870);
xor U5886 (N_5886,N_1121,N_3067);
xnor U5887 (N_5887,N_2669,N_404);
or U5888 (N_5888,N_3353,N_2223);
nor U5889 (N_5889,N_2211,N_139);
nor U5890 (N_5890,N_988,N_446);
xor U5891 (N_5891,N_1162,N_904);
nand U5892 (N_5892,N_736,N_3256);
or U5893 (N_5893,N_3343,N_1571);
and U5894 (N_5894,N_2782,N_1698);
and U5895 (N_5895,N_3805,N_2619);
or U5896 (N_5896,N_605,N_1004);
and U5897 (N_5897,N_3434,N_3718);
or U5898 (N_5898,N_1531,N_357);
nor U5899 (N_5899,N_1213,N_198);
xor U5900 (N_5900,N_1572,N_592);
xor U5901 (N_5901,N_3486,N_1191);
xor U5902 (N_5902,N_379,N_238);
and U5903 (N_5903,N_3722,N_281);
xor U5904 (N_5904,N_2595,N_1511);
nand U5905 (N_5905,N_2725,N_2787);
xor U5906 (N_5906,N_119,N_1037);
or U5907 (N_5907,N_3596,N_2617);
nor U5908 (N_5908,N_2317,N_1170);
or U5909 (N_5909,N_1308,N_2691);
nor U5910 (N_5910,N_1472,N_3646);
xnor U5911 (N_5911,N_1172,N_648);
nand U5912 (N_5912,N_3829,N_3780);
or U5913 (N_5913,N_1536,N_1438);
nor U5914 (N_5914,N_797,N_3000);
and U5915 (N_5915,N_2651,N_3004);
nor U5916 (N_5916,N_1641,N_3799);
and U5917 (N_5917,N_3276,N_1604);
and U5918 (N_5918,N_3417,N_3926);
xnor U5919 (N_5919,N_2968,N_1687);
and U5920 (N_5920,N_818,N_286);
and U5921 (N_5921,N_3114,N_2613);
or U5922 (N_5922,N_1099,N_528);
xnor U5923 (N_5923,N_3705,N_2352);
nand U5924 (N_5924,N_2106,N_1161);
nor U5925 (N_5925,N_2757,N_49);
xnor U5926 (N_5926,N_2131,N_1742);
nand U5927 (N_5927,N_2985,N_3410);
and U5928 (N_5928,N_1487,N_2380);
or U5929 (N_5929,N_3571,N_2071);
or U5930 (N_5930,N_759,N_2337);
nor U5931 (N_5931,N_1331,N_2517);
xor U5932 (N_5932,N_3544,N_39);
xnor U5933 (N_5933,N_885,N_1941);
or U5934 (N_5934,N_1202,N_542);
xnor U5935 (N_5935,N_3025,N_2891);
or U5936 (N_5936,N_3497,N_1217);
xnor U5937 (N_5937,N_57,N_2079);
or U5938 (N_5938,N_2901,N_670);
nand U5939 (N_5939,N_2148,N_1085);
nand U5940 (N_5940,N_2908,N_1540);
nor U5941 (N_5941,N_1864,N_1026);
or U5942 (N_5942,N_2815,N_2631);
and U5943 (N_5943,N_3053,N_254);
or U5944 (N_5944,N_991,N_849);
nor U5945 (N_5945,N_1543,N_2879);
xnor U5946 (N_5946,N_2389,N_1039);
xor U5947 (N_5947,N_1370,N_1910);
or U5948 (N_5948,N_1932,N_2562);
xnor U5949 (N_5949,N_1391,N_930);
nand U5950 (N_5950,N_2199,N_867);
nor U5951 (N_5951,N_742,N_676);
xor U5952 (N_5952,N_1264,N_1650);
or U5953 (N_5953,N_635,N_46);
and U5954 (N_5954,N_3333,N_190);
xor U5955 (N_5955,N_3942,N_681);
nor U5956 (N_5956,N_1867,N_3980);
and U5957 (N_5957,N_1807,N_2367);
nand U5958 (N_5958,N_3538,N_715);
and U5959 (N_5959,N_2917,N_1100);
nand U5960 (N_5960,N_1873,N_3765);
nand U5961 (N_5961,N_3427,N_1054);
or U5962 (N_5962,N_2073,N_1772);
or U5963 (N_5963,N_2546,N_3405);
xor U5964 (N_5964,N_600,N_464);
xor U5965 (N_5965,N_1096,N_2434);
nand U5966 (N_5966,N_2664,N_727);
and U5967 (N_5967,N_3665,N_701);
or U5968 (N_5968,N_3851,N_3862);
or U5969 (N_5969,N_3689,N_2228);
nand U5970 (N_5970,N_980,N_3296);
xor U5971 (N_5971,N_1198,N_690);
nor U5972 (N_5972,N_3701,N_1762);
xor U5973 (N_5973,N_1801,N_296);
and U5974 (N_5974,N_309,N_989);
nor U5975 (N_5975,N_3136,N_1058);
and U5976 (N_5976,N_3540,N_640);
nand U5977 (N_5977,N_2703,N_471);
and U5978 (N_5978,N_145,N_2208);
nand U5979 (N_5979,N_11,N_3608);
or U5980 (N_5980,N_2214,N_3033);
or U5981 (N_5981,N_1183,N_3840);
xnor U5982 (N_5982,N_3657,N_3911);
nor U5983 (N_5983,N_2626,N_23);
nand U5984 (N_5984,N_2008,N_1686);
nand U5985 (N_5985,N_3008,N_1475);
and U5986 (N_5986,N_3317,N_428);
nor U5987 (N_5987,N_1939,N_879);
nand U5988 (N_5988,N_578,N_154);
nand U5989 (N_5989,N_1136,N_934);
and U5990 (N_5990,N_1119,N_2511);
nor U5991 (N_5991,N_171,N_386);
or U5992 (N_5992,N_1173,N_3745);
and U5993 (N_5993,N_2932,N_2218);
xor U5994 (N_5994,N_2031,N_1205);
or U5995 (N_5995,N_283,N_413);
nand U5996 (N_5996,N_2261,N_807);
nor U5997 (N_5997,N_2805,N_3958);
or U5998 (N_5998,N_2227,N_490);
or U5999 (N_5999,N_1007,N_3240);
or U6000 (N_6000,N_416,N_1897);
nor U6001 (N_6001,N_1099,N_3186);
and U6002 (N_6002,N_3530,N_2648);
and U6003 (N_6003,N_3430,N_3875);
and U6004 (N_6004,N_2300,N_1969);
or U6005 (N_6005,N_3704,N_1224);
nor U6006 (N_6006,N_1164,N_979);
xnor U6007 (N_6007,N_3707,N_3477);
xnor U6008 (N_6008,N_1473,N_216);
and U6009 (N_6009,N_3052,N_672);
and U6010 (N_6010,N_3888,N_2539);
and U6011 (N_6011,N_1597,N_1277);
and U6012 (N_6012,N_2844,N_3386);
or U6013 (N_6013,N_3499,N_3840);
and U6014 (N_6014,N_1796,N_1605);
nor U6015 (N_6015,N_3895,N_3237);
nor U6016 (N_6016,N_463,N_1592);
or U6017 (N_6017,N_3007,N_1335);
xor U6018 (N_6018,N_2066,N_2655);
and U6019 (N_6019,N_529,N_1855);
xor U6020 (N_6020,N_580,N_380);
nand U6021 (N_6021,N_3296,N_1225);
or U6022 (N_6022,N_1408,N_2781);
nor U6023 (N_6023,N_465,N_2976);
xor U6024 (N_6024,N_3071,N_1057);
nor U6025 (N_6025,N_2240,N_2736);
and U6026 (N_6026,N_9,N_891);
nand U6027 (N_6027,N_3399,N_3702);
and U6028 (N_6028,N_188,N_659);
or U6029 (N_6029,N_3371,N_3713);
nand U6030 (N_6030,N_2589,N_2723);
and U6031 (N_6031,N_1604,N_595);
xnor U6032 (N_6032,N_137,N_2517);
and U6033 (N_6033,N_591,N_23);
nand U6034 (N_6034,N_2558,N_3575);
nand U6035 (N_6035,N_2219,N_584);
xnor U6036 (N_6036,N_665,N_3490);
and U6037 (N_6037,N_1819,N_890);
nor U6038 (N_6038,N_2699,N_1654);
xnor U6039 (N_6039,N_1272,N_450);
nand U6040 (N_6040,N_922,N_3673);
and U6041 (N_6041,N_2563,N_1408);
nor U6042 (N_6042,N_529,N_1016);
and U6043 (N_6043,N_3654,N_1484);
and U6044 (N_6044,N_2955,N_1307);
xnor U6045 (N_6045,N_2276,N_1757);
xor U6046 (N_6046,N_2826,N_2808);
or U6047 (N_6047,N_1446,N_2549);
or U6048 (N_6048,N_3383,N_1766);
and U6049 (N_6049,N_2226,N_791);
nand U6050 (N_6050,N_1025,N_1336);
nor U6051 (N_6051,N_599,N_2373);
or U6052 (N_6052,N_1159,N_1648);
or U6053 (N_6053,N_1258,N_692);
nand U6054 (N_6054,N_3310,N_2666);
or U6055 (N_6055,N_2389,N_3797);
or U6056 (N_6056,N_533,N_776);
nand U6057 (N_6057,N_3717,N_978);
nor U6058 (N_6058,N_684,N_2068);
or U6059 (N_6059,N_2827,N_2578);
and U6060 (N_6060,N_44,N_2650);
or U6061 (N_6061,N_3018,N_1630);
xnor U6062 (N_6062,N_2684,N_1376);
and U6063 (N_6063,N_881,N_3749);
nand U6064 (N_6064,N_1595,N_2975);
or U6065 (N_6065,N_3848,N_350);
or U6066 (N_6066,N_3132,N_1818);
xor U6067 (N_6067,N_2696,N_1092);
nand U6068 (N_6068,N_3834,N_618);
nand U6069 (N_6069,N_3954,N_3579);
nand U6070 (N_6070,N_2940,N_3800);
nand U6071 (N_6071,N_100,N_2825);
nor U6072 (N_6072,N_1372,N_1222);
nand U6073 (N_6073,N_777,N_1674);
nor U6074 (N_6074,N_3838,N_151);
and U6075 (N_6075,N_786,N_3656);
and U6076 (N_6076,N_2404,N_965);
and U6077 (N_6077,N_2896,N_158);
or U6078 (N_6078,N_3352,N_1034);
or U6079 (N_6079,N_1115,N_3085);
xnor U6080 (N_6080,N_1509,N_2779);
or U6081 (N_6081,N_683,N_998);
nor U6082 (N_6082,N_722,N_3228);
xor U6083 (N_6083,N_3203,N_115);
nor U6084 (N_6084,N_1941,N_2780);
or U6085 (N_6085,N_23,N_505);
and U6086 (N_6086,N_3994,N_3792);
or U6087 (N_6087,N_3833,N_2039);
or U6088 (N_6088,N_1879,N_1853);
nor U6089 (N_6089,N_2973,N_3855);
nand U6090 (N_6090,N_3202,N_3334);
and U6091 (N_6091,N_108,N_3508);
nor U6092 (N_6092,N_907,N_2407);
nor U6093 (N_6093,N_2427,N_2850);
nor U6094 (N_6094,N_1982,N_2975);
and U6095 (N_6095,N_155,N_3660);
or U6096 (N_6096,N_1335,N_1701);
and U6097 (N_6097,N_1930,N_2907);
nor U6098 (N_6098,N_117,N_2083);
nor U6099 (N_6099,N_1441,N_2655);
and U6100 (N_6100,N_1814,N_811);
nor U6101 (N_6101,N_2788,N_1011);
or U6102 (N_6102,N_3370,N_92);
nor U6103 (N_6103,N_3843,N_2447);
nor U6104 (N_6104,N_3318,N_1900);
xnor U6105 (N_6105,N_1518,N_3400);
nand U6106 (N_6106,N_1573,N_2923);
nand U6107 (N_6107,N_3877,N_2098);
nor U6108 (N_6108,N_1874,N_2158);
and U6109 (N_6109,N_297,N_2149);
nor U6110 (N_6110,N_3396,N_2029);
xor U6111 (N_6111,N_2292,N_970);
xnor U6112 (N_6112,N_3863,N_2672);
nor U6113 (N_6113,N_3879,N_51);
nand U6114 (N_6114,N_721,N_2345);
nor U6115 (N_6115,N_390,N_1658);
nand U6116 (N_6116,N_3388,N_797);
xor U6117 (N_6117,N_2768,N_1975);
and U6118 (N_6118,N_2709,N_3286);
nand U6119 (N_6119,N_3569,N_2419);
or U6120 (N_6120,N_2903,N_1913);
nor U6121 (N_6121,N_1673,N_689);
or U6122 (N_6122,N_2246,N_2223);
or U6123 (N_6123,N_3533,N_3465);
nor U6124 (N_6124,N_2086,N_988);
and U6125 (N_6125,N_1906,N_2121);
nand U6126 (N_6126,N_3534,N_3686);
nand U6127 (N_6127,N_1757,N_955);
or U6128 (N_6128,N_3581,N_3733);
nor U6129 (N_6129,N_2655,N_2272);
or U6130 (N_6130,N_2630,N_1871);
nand U6131 (N_6131,N_1638,N_649);
xnor U6132 (N_6132,N_1679,N_2399);
and U6133 (N_6133,N_474,N_472);
or U6134 (N_6134,N_2577,N_2511);
or U6135 (N_6135,N_1817,N_3782);
or U6136 (N_6136,N_2025,N_2587);
nand U6137 (N_6137,N_1068,N_2699);
nand U6138 (N_6138,N_75,N_3081);
xor U6139 (N_6139,N_606,N_2385);
nand U6140 (N_6140,N_2143,N_3942);
and U6141 (N_6141,N_2588,N_1989);
and U6142 (N_6142,N_1635,N_1163);
nand U6143 (N_6143,N_167,N_3387);
nor U6144 (N_6144,N_340,N_3816);
nor U6145 (N_6145,N_3473,N_3823);
nand U6146 (N_6146,N_3139,N_313);
xor U6147 (N_6147,N_2544,N_1114);
or U6148 (N_6148,N_3671,N_2807);
nand U6149 (N_6149,N_1678,N_168);
and U6150 (N_6150,N_3241,N_1790);
or U6151 (N_6151,N_563,N_1011);
nor U6152 (N_6152,N_204,N_1366);
nor U6153 (N_6153,N_3186,N_1113);
xor U6154 (N_6154,N_1896,N_610);
nor U6155 (N_6155,N_3284,N_2212);
xnor U6156 (N_6156,N_2208,N_3991);
or U6157 (N_6157,N_284,N_2436);
nand U6158 (N_6158,N_758,N_949);
xor U6159 (N_6159,N_2124,N_3682);
nor U6160 (N_6160,N_3932,N_410);
nand U6161 (N_6161,N_2814,N_3021);
nand U6162 (N_6162,N_1120,N_973);
nand U6163 (N_6163,N_2243,N_1961);
and U6164 (N_6164,N_672,N_347);
and U6165 (N_6165,N_3428,N_2676);
nand U6166 (N_6166,N_503,N_2656);
xnor U6167 (N_6167,N_3107,N_2115);
and U6168 (N_6168,N_3953,N_1278);
and U6169 (N_6169,N_298,N_2758);
and U6170 (N_6170,N_3732,N_2216);
nor U6171 (N_6171,N_3964,N_1797);
or U6172 (N_6172,N_705,N_3643);
xor U6173 (N_6173,N_3466,N_141);
xor U6174 (N_6174,N_3328,N_1655);
or U6175 (N_6175,N_1794,N_3922);
xnor U6176 (N_6176,N_2539,N_546);
and U6177 (N_6177,N_1349,N_3726);
nand U6178 (N_6178,N_1179,N_37);
nor U6179 (N_6179,N_3795,N_1478);
or U6180 (N_6180,N_1109,N_737);
and U6181 (N_6181,N_2487,N_3327);
or U6182 (N_6182,N_3190,N_61);
or U6183 (N_6183,N_1333,N_3433);
or U6184 (N_6184,N_3902,N_124);
xnor U6185 (N_6185,N_1338,N_2053);
and U6186 (N_6186,N_3871,N_1076);
nor U6187 (N_6187,N_3030,N_2136);
nand U6188 (N_6188,N_2396,N_1884);
and U6189 (N_6189,N_2387,N_104);
nand U6190 (N_6190,N_3375,N_1018);
nor U6191 (N_6191,N_1240,N_2807);
nand U6192 (N_6192,N_1618,N_1587);
nor U6193 (N_6193,N_1109,N_2831);
and U6194 (N_6194,N_2246,N_181);
nand U6195 (N_6195,N_3506,N_3170);
nor U6196 (N_6196,N_1494,N_2506);
and U6197 (N_6197,N_2522,N_1658);
nand U6198 (N_6198,N_1390,N_3661);
xnor U6199 (N_6199,N_3791,N_2905);
nand U6200 (N_6200,N_1925,N_3090);
nand U6201 (N_6201,N_963,N_2052);
and U6202 (N_6202,N_3299,N_423);
nand U6203 (N_6203,N_2490,N_1365);
nor U6204 (N_6204,N_3138,N_801);
nand U6205 (N_6205,N_3157,N_2352);
or U6206 (N_6206,N_1594,N_1239);
and U6207 (N_6207,N_3185,N_1483);
nor U6208 (N_6208,N_1596,N_1194);
or U6209 (N_6209,N_2672,N_3636);
nor U6210 (N_6210,N_1432,N_3924);
or U6211 (N_6211,N_1237,N_282);
and U6212 (N_6212,N_1229,N_994);
nor U6213 (N_6213,N_1846,N_2510);
xnor U6214 (N_6214,N_1059,N_2091);
nor U6215 (N_6215,N_3460,N_292);
and U6216 (N_6216,N_2793,N_971);
or U6217 (N_6217,N_3003,N_3401);
nor U6218 (N_6218,N_2811,N_928);
nor U6219 (N_6219,N_3637,N_3709);
or U6220 (N_6220,N_342,N_2394);
and U6221 (N_6221,N_1437,N_423);
xnor U6222 (N_6222,N_2917,N_1638);
nor U6223 (N_6223,N_1686,N_2009);
xor U6224 (N_6224,N_1235,N_3454);
nor U6225 (N_6225,N_2713,N_419);
nand U6226 (N_6226,N_501,N_2645);
and U6227 (N_6227,N_3759,N_2423);
xnor U6228 (N_6228,N_1019,N_3567);
or U6229 (N_6229,N_3426,N_525);
and U6230 (N_6230,N_670,N_983);
nand U6231 (N_6231,N_3817,N_3005);
nand U6232 (N_6232,N_3290,N_46);
or U6233 (N_6233,N_3201,N_2394);
nand U6234 (N_6234,N_1941,N_3063);
or U6235 (N_6235,N_2074,N_3627);
nor U6236 (N_6236,N_468,N_3305);
nor U6237 (N_6237,N_1255,N_1074);
or U6238 (N_6238,N_2344,N_2800);
and U6239 (N_6239,N_2208,N_3143);
nor U6240 (N_6240,N_3938,N_689);
nor U6241 (N_6241,N_3736,N_3976);
nor U6242 (N_6242,N_2426,N_3599);
xnor U6243 (N_6243,N_795,N_170);
and U6244 (N_6244,N_2640,N_342);
nand U6245 (N_6245,N_3241,N_256);
or U6246 (N_6246,N_3147,N_1841);
or U6247 (N_6247,N_1341,N_2076);
xnor U6248 (N_6248,N_3098,N_3283);
nor U6249 (N_6249,N_1353,N_1487);
xor U6250 (N_6250,N_289,N_400);
or U6251 (N_6251,N_3780,N_2502);
or U6252 (N_6252,N_3770,N_3289);
xor U6253 (N_6253,N_1353,N_1075);
nor U6254 (N_6254,N_2413,N_521);
or U6255 (N_6255,N_2392,N_1745);
or U6256 (N_6256,N_2701,N_1548);
or U6257 (N_6257,N_3961,N_2030);
nor U6258 (N_6258,N_2244,N_2120);
or U6259 (N_6259,N_1782,N_3146);
and U6260 (N_6260,N_993,N_2976);
nor U6261 (N_6261,N_1113,N_1368);
nor U6262 (N_6262,N_2384,N_920);
and U6263 (N_6263,N_407,N_3007);
nand U6264 (N_6264,N_2144,N_3653);
and U6265 (N_6265,N_1662,N_893);
xnor U6266 (N_6266,N_3620,N_2078);
nor U6267 (N_6267,N_3466,N_2270);
nor U6268 (N_6268,N_3640,N_2891);
xnor U6269 (N_6269,N_1736,N_2081);
nand U6270 (N_6270,N_2959,N_3868);
nand U6271 (N_6271,N_1661,N_2472);
or U6272 (N_6272,N_2459,N_2540);
or U6273 (N_6273,N_956,N_996);
and U6274 (N_6274,N_339,N_2126);
nand U6275 (N_6275,N_3292,N_2321);
nand U6276 (N_6276,N_1502,N_1393);
or U6277 (N_6277,N_448,N_1451);
nand U6278 (N_6278,N_120,N_1026);
xor U6279 (N_6279,N_1061,N_3982);
nor U6280 (N_6280,N_166,N_2129);
or U6281 (N_6281,N_762,N_3202);
and U6282 (N_6282,N_1501,N_2961);
nand U6283 (N_6283,N_2247,N_832);
and U6284 (N_6284,N_591,N_380);
or U6285 (N_6285,N_3776,N_927);
or U6286 (N_6286,N_2093,N_1975);
or U6287 (N_6287,N_1372,N_1364);
xnor U6288 (N_6288,N_3796,N_188);
nor U6289 (N_6289,N_2957,N_2649);
and U6290 (N_6290,N_2275,N_2741);
nor U6291 (N_6291,N_2423,N_639);
nand U6292 (N_6292,N_2608,N_138);
nor U6293 (N_6293,N_425,N_146);
nand U6294 (N_6294,N_3461,N_3213);
or U6295 (N_6295,N_2210,N_1181);
nor U6296 (N_6296,N_2625,N_3341);
or U6297 (N_6297,N_648,N_2312);
xor U6298 (N_6298,N_132,N_3046);
xor U6299 (N_6299,N_2919,N_539);
nor U6300 (N_6300,N_1187,N_3645);
nand U6301 (N_6301,N_1001,N_324);
nor U6302 (N_6302,N_1326,N_1386);
xnor U6303 (N_6303,N_3600,N_2790);
xor U6304 (N_6304,N_3251,N_3351);
xnor U6305 (N_6305,N_552,N_31);
nor U6306 (N_6306,N_2519,N_2736);
and U6307 (N_6307,N_2357,N_1067);
nor U6308 (N_6308,N_1488,N_2435);
nor U6309 (N_6309,N_2685,N_744);
nand U6310 (N_6310,N_641,N_3613);
xor U6311 (N_6311,N_3722,N_3828);
nor U6312 (N_6312,N_910,N_3342);
nor U6313 (N_6313,N_1275,N_709);
nand U6314 (N_6314,N_2307,N_3277);
nor U6315 (N_6315,N_3104,N_1594);
nor U6316 (N_6316,N_2877,N_2249);
xor U6317 (N_6317,N_2111,N_2736);
nor U6318 (N_6318,N_1510,N_2162);
or U6319 (N_6319,N_1033,N_3163);
xnor U6320 (N_6320,N_1297,N_1859);
nand U6321 (N_6321,N_27,N_720);
and U6322 (N_6322,N_353,N_1702);
nand U6323 (N_6323,N_1933,N_1669);
and U6324 (N_6324,N_1966,N_3655);
nand U6325 (N_6325,N_2672,N_3536);
nand U6326 (N_6326,N_598,N_1041);
and U6327 (N_6327,N_1898,N_3195);
xor U6328 (N_6328,N_2495,N_2907);
or U6329 (N_6329,N_3205,N_460);
or U6330 (N_6330,N_2779,N_2528);
xor U6331 (N_6331,N_438,N_1692);
and U6332 (N_6332,N_3009,N_3257);
nand U6333 (N_6333,N_2297,N_962);
nand U6334 (N_6334,N_3374,N_3940);
xnor U6335 (N_6335,N_2656,N_2740);
nor U6336 (N_6336,N_1442,N_314);
or U6337 (N_6337,N_1200,N_1834);
nand U6338 (N_6338,N_3200,N_111);
or U6339 (N_6339,N_1390,N_2234);
nand U6340 (N_6340,N_631,N_1191);
nand U6341 (N_6341,N_693,N_840);
nand U6342 (N_6342,N_3710,N_700);
and U6343 (N_6343,N_2558,N_851);
xnor U6344 (N_6344,N_677,N_2278);
nor U6345 (N_6345,N_1446,N_574);
and U6346 (N_6346,N_2031,N_2597);
and U6347 (N_6347,N_1401,N_1026);
or U6348 (N_6348,N_3472,N_759);
or U6349 (N_6349,N_455,N_451);
or U6350 (N_6350,N_1003,N_2170);
nor U6351 (N_6351,N_2055,N_3755);
nor U6352 (N_6352,N_1609,N_46);
and U6353 (N_6353,N_3859,N_1106);
xor U6354 (N_6354,N_2854,N_348);
or U6355 (N_6355,N_532,N_2198);
nor U6356 (N_6356,N_543,N_793);
nand U6357 (N_6357,N_481,N_2490);
xor U6358 (N_6358,N_3837,N_1470);
nand U6359 (N_6359,N_2862,N_2434);
or U6360 (N_6360,N_3499,N_3695);
and U6361 (N_6361,N_2439,N_1435);
xnor U6362 (N_6362,N_979,N_648);
nand U6363 (N_6363,N_3228,N_1149);
xnor U6364 (N_6364,N_336,N_2524);
or U6365 (N_6365,N_3897,N_3524);
or U6366 (N_6366,N_3202,N_2215);
or U6367 (N_6367,N_1875,N_2025);
nand U6368 (N_6368,N_51,N_538);
and U6369 (N_6369,N_3329,N_3695);
and U6370 (N_6370,N_1579,N_3050);
and U6371 (N_6371,N_1397,N_3858);
nand U6372 (N_6372,N_2592,N_2526);
xnor U6373 (N_6373,N_3058,N_1794);
and U6374 (N_6374,N_759,N_1315);
xnor U6375 (N_6375,N_1899,N_2318);
or U6376 (N_6376,N_3915,N_2020);
nand U6377 (N_6377,N_744,N_114);
nand U6378 (N_6378,N_3199,N_3890);
xnor U6379 (N_6379,N_977,N_2568);
and U6380 (N_6380,N_1265,N_820);
nand U6381 (N_6381,N_1529,N_3996);
xnor U6382 (N_6382,N_2423,N_1031);
and U6383 (N_6383,N_3017,N_3771);
nor U6384 (N_6384,N_3845,N_3796);
xor U6385 (N_6385,N_3598,N_728);
xnor U6386 (N_6386,N_3780,N_404);
xnor U6387 (N_6387,N_1628,N_1985);
and U6388 (N_6388,N_134,N_3500);
and U6389 (N_6389,N_1870,N_3742);
nor U6390 (N_6390,N_507,N_1058);
xnor U6391 (N_6391,N_3517,N_3983);
nand U6392 (N_6392,N_1031,N_1959);
nand U6393 (N_6393,N_2244,N_3743);
and U6394 (N_6394,N_2867,N_997);
or U6395 (N_6395,N_3958,N_327);
nand U6396 (N_6396,N_2236,N_1236);
and U6397 (N_6397,N_2276,N_2785);
xor U6398 (N_6398,N_578,N_2129);
nand U6399 (N_6399,N_2673,N_3819);
xnor U6400 (N_6400,N_1691,N_2382);
nor U6401 (N_6401,N_1611,N_15);
nand U6402 (N_6402,N_3841,N_3590);
xor U6403 (N_6403,N_1219,N_1782);
or U6404 (N_6404,N_3145,N_1009);
nand U6405 (N_6405,N_3737,N_1192);
or U6406 (N_6406,N_3539,N_3793);
nor U6407 (N_6407,N_2864,N_1969);
nand U6408 (N_6408,N_893,N_2652);
nor U6409 (N_6409,N_3422,N_496);
nand U6410 (N_6410,N_3009,N_340);
or U6411 (N_6411,N_3098,N_412);
nand U6412 (N_6412,N_2196,N_1213);
nor U6413 (N_6413,N_921,N_2733);
nand U6414 (N_6414,N_2072,N_2423);
nand U6415 (N_6415,N_3850,N_3183);
and U6416 (N_6416,N_1825,N_3516);
nor U6417 (N_6417,N_1372,N_210);
or U6418 (N_6418,N_2452,N_744);
or U6419 (N_6419,N_338,N_2951);
xor U6420 (N_6420,N_1227,N_3568);
nand U6421 (N_6421,N_1527,N_811);
nor U6422 (N_6422,N_151,N_1849);
nand U6423 (N_6423,N_571,N_1622);
xor U6424 (N_6424,N_772,N_3314);
and U6425 (N_6425,N_3345,N_1200);
nand U6426 (N_6426,N_2395,N_1606);
nor U6427 (N_6427,N_1886,N_3781);
xnor U6428 (N_6428,N_3640,N_87);
xor U6429 (N_6429,N_1918,N_736);
or U6430 (N_6430,N_1456,N_237);
or U6431 (N_6431,N_3058,N_1689);
nor U6432 (N_6432,N_1082,N_18);
xor U6433 (N_6433,N_2477,N_94);
and U6434 (N_6434,N_3855,N_635);
nor U6435 (N_6435,N_3260,N_3018);
and U6436 (N_6436,N_781,N_2260);
xor U6437 (N_6437,N_2326,N_3197);
nand U6438 (N_6438,N_3896,N_1903);
xor U6439 (N_6439,N_35,N_2116);
or U6440 (N_6440,N_1325,N_532);
xor U6441 (N_6441,N_3436,N_1982);
and U6442 (N_6442,N_3213,N_3321);
and U6443 (N_6443,N_3304,N_234);
nand U6444 (N_6444,N_3527,N_3290);
nand U6445 (N_6445,N_864,N_832);
nor U6446 (N_6446,N_631,N_979);
nor U6447 (N_6447,N_1288,N_1116);
nand U6448 (N_6448,N_1116,N_965);
nand U6449 (N_6449,N_100,N_1883);
and U6450 (N_6450,N_3522,N_3577);
nor U6451 (N_6451,N_1243,N_3343);
nand U6452 (N_6452,N_3046,N_2119);
nor U6453 (N_6453,N_1447,N_2504);
and U6454 (N_6454,N_117,N_3325);
nor U6455 (N_6455,N_862,N_1948);
and U6456 (N_6456,N_2872,N_2762);
and U6457 (N_6457,N_2716,N_3957);
xor U6458 (N_6458,N_2709,N_3915);
nor U6459 (N_6459,N_2090,N_1986);
and U6460 (N_6460,N_2791,N_2445);
and U6461 (N_6461,N_3230,N_3488);
or U6462 (N_6462,N_262,N_539);
or U6463 (N_6463,N_2141,N_1486);
or U6464 (N_6464,N_2600,N_2147);
nor U6465 (N_6465,N_1183,N_702);
and U6466 (N_6466,N_1047,N_1406);
nand U6467 (N_6467,N_3126,N_2996);
xnor U6468 (N_6468,N_3028,N_3825);
xor U6469 (N_6469,N_616,N_3539);
nand U6470 (N_6470,N_1885,N_759);
or U6471 (N_6471,N_249,N_659);
xnor U6472 (N_6472,N_1289,N_1592);
xnor U6473 (N_6473,N_1238,N_2690);
nor U6474 (N_6474,N_3379,N_105);
nor U6475 (N_6475,N_3216,N_331);
nor U6476 (N_6476,N_546,N_1224);
and U6477 (N_6477,N_2095,N_1654);
nor U6478 (N_6478,N_2561,N_3074);
and U6479 (N_6479,N_668,N_1933);
xnor U6480 (N_6480,N_2101,N_2842);
xor U6481 (N_6481,N_3684,N_238);
xor U6482 (N_6482,N_2892,N_2871);
and U6483 (N_6483,N_2573,N_2809);
xor U6484 (N_6484,N_2748,N_1897);
xnor U6485 (N_6485,N_1787,N_2354);
or U6486 (N_6486,N_3356,N_1975);
nand U6487 (N_6487,N_639,N_1431);
xnor U6488 (N_6488,N_1272,N_798);
nor U6489 (N_6489,N_3030,N_277);
or U6490 (N_6490,N_927,N_3005);
nor U6491 (N_6491,N_2753,N_1043);
and U6492 (N_6492,N_3647,N_166);
or U6493 (N_6493,N_2854,N_2406);
nor U6494 (N_6494,N_1515,N_127);
and U6495 (N_6495,N_758,N_803);
nor U6496 (N_6496,N_3581,N_2159);
and U6497 (N_6497,N_1437,N_2622);
or U6498 (N_6498,N_2991,N_120);
nor U6499 (N_6499,N_357,N_324);
nor U6500 (N_6500,N_2685,N_1273);
xor U6501 (N_6501,N_2960,N_3711);
nand U6502 (N_6502,N_701,N_2008);
xnor U6503 (N_6503,N_576,N_476);
nor U6504 (N_6504,N_3438,N_1405);
nor U6505 (N_6505,N_2540,N_3990);
or U6506 (N_6506,N_2332,N_2181);
or U6507 (N_6507,N_2715,N_1891);
or U6508 (N_6508,N_494,N_508);
nor U6509 (N_6509,N_357,N_2760);
and U6510 (N_6510,N_11,N_3680);
and U6511 (N_6511,N_1616,N_730);
nor U6512 (N_6512,N_1903,N_2155);
and U6513 (N_6513,N_2189,N_959);
nor U6514 (N_6514,N_3903,N_3941);
nand U6515 (N_6515,N_139,N_2534);
nor U6516 (N_6516,N_2682,N_2511);
nor U6517 (N_6517,N_1867,N_1272);
nor U6518 (N_6518,N_1600,N_2931);
and U6519 (N_6519,N_1173,N_3515);
or U6520 (N_6520,N_976,N_3881);
xor U6521 (N_6521,N_600,N_1687);
xor U6522 (N_6522,N_374,N_3812);
xnor U6523 (N_6523,N_3507,N_603);
and U6524 (N_6524,N_2100,N_3576);
or U6525 (N_6525,N_3679,N_871);
nand U6526 (N_6526,N_3849,N_3403);
xnor U6527 (N_6527,N_2726,N_3235);
nor U6528 (N_6528,N_686,N_715);
and U6529 (N_6529,N_1634,N_404);
or U6530 (N_6530,N_540,N_1533);
nor U6531 (N_6531,N_1219,N_2016);
or U6532 (N_6532,N_2063,N_357);
nor U6533 (N_6533,N_1623,N_3730);
and U6534 (N_6534,N_1174,N_2103);
nand U6535 (N_6535,N_3747,N_2277);
nor U6536 (N_6536,N_1245,N_952);
and U6537 (N_6537,N_3285,N_693);
nor U6538 (N_6538,N_3593,N_1692);
xnor U6539 (N_6539,N_2931,N_1604);
and U6540 (N_6540,N_2421,N_2449);
xnor U6541 (N_6541,N_429,N_2521);
nor U6542 (N_6542,N_2136,N_3468);
or U6543 (N_6543,N_3847,N_3038);
xnor U6544 (N_6544,N_2310,N_3498);
or U6545 (N_6545,N_463,N_1719);
nand U6546 (N_6546,N_1170,N_1619);
nand U6547 (N_6547,N_2790,N_3929);
and U6548 (N_6548,N_454,N_2645);
and U6549 (N_6549,N_2180,N_1589);
and U6550 (N_6550,N_2323,N_3190);
or U6551 (N_6551,N_137,N_2812);
xnor U6552 (N_6552,N_1596,N_1294);
nor U6553 (N_6553,N_2815,N_905);
or U6554 (N_6554,N_3870,N_3338);
nor U6555 (N_6555,N_1447,N_2383);
nand U6556 (N_6556,N_2235,N_1970);
and U6557 (N_6557,N_490,N_1421);
nand U6558 (N_6558,N_590,N_743);
nand U6559 (N_6559,N_2428,N_3872);
or U6560 (N_6560,N_725,N_1271);
and U6561 (N_6561,N_3868,N_962);
xnor U6562 (N_6562,N_710,N_3548);
xor U6563 (N_6563,N_1203,N_698);
nor U6564 (N_6564,N_2135,N_759);
nand U6565 (N_6565,N_595,N_3395);
or U6566 (N_6566,N_285,N_1923);
and U6567 (N_6567,N_2436,N_2863);
and U6568 (N_6568,N_2592,N_3759);
nor U6569 (N_6569,N_2157,N_1953);
and U6570 (N_6570,N_3742,N_909);
xnor U6571 (N_6571,N_2874,N_3395);
nand U6572 (N_6572,N_1186,N_669);
xnor U6573 (N_6573,N_1485,N_1781);
nor U6574 (N_6574,N_1334,N_478);
nor U6575 (N_6575,N_2368,N_587);
and U6576 (N_6576,N_487,N_3582);
nand U6577 (N_6577,N_2605,N_271);
nand U6578 (N_6578,N_2755,N_3654);
nand U6579 (N_6579,N_1889,N_668);
xor U6580 (N_6580,N_1897,N_2936);
nand U6581 (N_6581,N_553,N_714);
nand U6582 (N_6582,N_2463,N_2507);
or U6583 (N_6583,N_3396,N_3400);
nor U6584 (N_6584,N_1699,N_1245);
or U6585 (N_6585,N_2308,N_3182);
nand U6586 (N_6586,N_2214,N_1965);
nand U6587 (N_6587,N_3986,N_3759);
nor U6588 (N_6588,N_318,N_2266);
and U6589 (N_6589,N_192,N_49);
nand U6590 (N_6590,N_322,N_303);
nand U6591 (N_6591,N_215,N_201);
xor U6592 (N_6592,N_3358,N_1419);
nand U6593 (N_6593,N_1966,N_913);
xor U6594 (N_6594,N_3844,N_3791);
or U6595 (N_6595,N_1632,N_188);
xnor U6596 (N_6596,N_594,N_1668);
nor U6597 (N_6597,N_2207,N_2109);
and U6598 (N_6598,N_2733,N_979);
nor U6599 (N_6599,N_2927,N_3594);
xor U6600 (N_6600,N_3615,N_2663);
nor U6601 (N_6601,N_961,N_1576);
and U6602 (N_6602,N_1419,N_3774);
nand U6603 (N_6603,N_533,N_2687);
or U6604 (N_6604,N_2268,N_1761);
and U6605 (N_6605,N_2090,N_2493);
xnor U6606 (N_6606,N_3501,N_138);
xor U6607 (N_6607,N_1238,N_1107);
and U6608 (N_6608,N_2294,N_766);
and U6609 (N_6609,N_529,N_3626);
nand U6610 (N_6610,N_697,N_1124);
nor U6611 (N_6611,N_1865,N_737);
and U6612 (N_6612,N_2038,N_3132);
and U6613 (N_6613,N_2950,N_2692);
or U6614 (N_6614,N_2161,N_983);
nor U6615 (N_6615,N_2386,N_432);
xor U6616 (N_6616,N_2915,N_103);
nand U6617 (N_6617,N_241,N_394);
or U6618 (N_6618,N_1873,N_2262);
nor U6619 (N_6619,N_277,N_2510);
xnor U6620 (N_6620,N_1579,N_1948);
nand U6621 (N_6621,N_2613,N_2839);
nor U6622 (N_6622,N_3130,N_1167);
nand U6623 (N_6623,N_2266,N_1737);
xor U6624 (N_6624,N_454,N_2896);
or U6625 (N_6625,N_2885,N_2454);
nand U6626 (N_6626,N_1706,N_1046);
nand U6627 (N_6627,N_3619,N_1298);
or U6628 (N_6628,N_3800,N_540);
and U6629 (N_6629,N_2738,N_3031);
xnor U6630 (N_6630,N_368,N_258);
or U6631 (N_6631,N_1292,N_1925);
or U6632 (N_6632,N_2157,N_3138);
and U6633 (N_6633,N_3199,N_672);
or U6634 (N_6634,N_1432,N_672);
and U6635 (N_6635,N_1338,N_1997);
or U6636 (N_6636,N_1596,N_1779);
and U6637 (N_6637,N_470,N_2959);
nor U6638 (N_6638,N_1813,N_383);
nor U6639 (N_6639,N_1523,N_2919);
nand U6640 (N_6640,N_2743,N_1828);
nand U6641 (N_6641,N_3943,N_1891);
or U6642 (N_6642,N_3518,N_192);
xnor U6643 (N_6643,N_3301,N_1364);
nor U6644 (N_6644,N_2339,N_625);
or U6645 (N_6645,N_3160,N_699);
xor U6646 (N_6646,N_1879,N_896);
or U6647 (N_6647,N_1542,N_1308);
xnor U6648 (N_6648,N_38,N_367);
nand U6649 (N_6649,N_2127,N_3087);
nor U6650 (N_6650,N_2789,N_1450);
xor U6651 (N_6651,N_2979,N_2105);
and U6652 (N_6652,N_1342,N_1880);
nor U6653 (N_6653,N_2196,N_3563);
xor U6654 (N_6654,N_3493,N_3164);
and U6655 (N_6655,N_1231,N_468);
nand U6656 (N_6656,N_3930,N_3519);
and U6657 (N_6657,N_2603,N_3734);
nor U6658 (N_6658,N_16,N_2624);
xnor U6659 (N_6659,N_2485,N_975);
nor U6660 (N_6660,N_2000,N_1333);
and U6661 (N_6661,N_3764,N_2710);
or U6662 (N_6662,N_2157,N_2608);
nand U6663 (N_6663,N_1221,N_218);
nor U6664 (N_6664,N_3478,N_3529);
nor U6665 (N_6665,N_215,N_2593);
or U6666 (N_6666,N_238,N_1155);
nor U6667 (N_6667,N_968,N_2988);
or U6668 (N_6668,N_3411,N_3775);
xnor U6669 (N_6669,N_2530,N_1893);
nand U6670 (N_6670,N_1020,N_816);
nor U6671 (N_6671,N_1478,N_3682);
or U6672 (N_6672,N_2878,N_3665);
nand U6673 (N_6673,N_308,N_3274);
xor U6674 (N_6674,N_1822,N_294);
xor U6675 (N_6675,N_1943,N_697);
and U6676 (N_6676,N_873,N_3195);
nor U6677 (N_6677,N_3679,N_1287);
and U6678 (N_6678,N_1892,N_2868);
and U6679 (N_6679,N_3254,N_2197);
xor U6680 (N_6680,N_2996,N_1503);
nand U6681 (N_6681,N_690,N_2383);
and U6682 (N_6682,N_3445,N_1552);
and U6683 (N_6683,N_2535,N_3313);
nor U6684 (N_6684,N_2858,N_232);
or U6685 (N_6685,N_1525,N_2158);
nor U6686 (N_6686,N_2045,N_3567);
nor U6687 (N_6687,N_692,N_1784);
xnor U6688 (N_6688,N_3482,N_3217);
xnor U6689 (N_6689,N_1193,N_3829);
xnor U6690 (N_6690,N_967,N_1045);
or U6691 (N_6691,N_3449,N_3060);
nor U6692 (N_6692,N_3172,N_326);
xnor U6693 (N_6693,N_2364,N_1841);
or U6694 (N_6694,N_3677,N_3034);
nand U6695 (N_6695,N_1567,N_630);
or U6696 (N_6696,N_270,N_2323);
and U6697 (N_6697,N_2505,N_3659);
and U6698 (N_6698,N_887,N_2483);
and U6699 (N_6699,N_457,N_1135);
and U6700 (N_6700,N_335,N_1380);
xnor U6701 (N_6701,N_2825,N_930);
or U6702 (N_6702,N_1310,N_2380);
nand U6703 (N_6703,N_2453,N_2218);
xor U6704 (N_6704,N_1044,N_3785);
nor U6705 (N_6705,N_3075,N_2456);
nor U6706 (N_6706,N_1944,N_3334);
and U6707 (N_6707,N_1512,N_4);
nand U6708 (N_6708,N_453,N_3627);
xnor U6709 (N_6709,N_1434,N_2409);
and U6710 (N_6710,N_2321,N_3826);
nand U6711 (N_6711,N_93,N_1633);
or U6712 (N_6712,N_2841,N_318);
nor U6713 (N_6713,N_2915,N_2599);
nand U6714 (N_6714,N_3548,N_190);
nor U6715 (N_6715,N_3658,N_2527);
xnor U6716 (N_6716,N_1687,N_3912);
or U6717 (N_6717,N_860,N_2917);
or U6718 (N_6718,N_2477,N_2325);
nor U6719 (N_6719,N_1936,N_1595);
nor U6720 (N_6720,N_3894,N_3461);
xnor U6721 (N_6721,N_667,N_3063);
or U6722 (N_6722,N_388,N_1458);
nand U6723 (N_6723,N_586,N_1611);
nor U6724 (N_6724,N_2332,N_2180);
or U6725 (N_6725,N_811,N_767);
nor U6726 (N_6726,N_3378,N_3606);
or U6727 (N_6727,N_2242,N_3353);
nand U6728 (N_6728,N_2999,N_751);
xnor U6729 (N_6729,N_2501,N_1532);
and U6730 (N_6730,N_337,N_665);
nand U6731 (N_6731,N_775,N_585);
xnor U6732 (N_6732,N_1946,N_1838);
xor U6733 (N_6733,N_1238,N_2380);
or U6734 (N_6734,N_2315,N_3824);
xor U6735 (N_6735,N_3256,N_3308);
nand U6736 (N_6736,N_2562,N_1323);
and U6737 (N_6737,N_1316,N_3717);
and U6738 (N_6738,N_2704,N_3681);
nand U6739 (N_6739,N_3432,N_3567);
nand U6740 (N_6740,N_33,N_191);
nor U6741 (N_6741,N_3062,N_2932);
xor U6742 (N_6742,N_407,N_839);
nand U6743 (N_6743,N_459,N_2538);
nand U6744 (N_6744,N_3520,N_2596);
nand U6745 (N_6745,N_1400,N_3823);
and U6746 (N_6746,N_2094,N_2500);
nor U6747 (N_6747,N_60,N_1986);
or U6748 (N_6748,N_2253,N_996);
and U6749 (N_6749,N_2327,N_103);
xnor U6750 (N_6750,N_799,N_2559);
or U6751 (N_6751,N_2466,N_996);
nand U6752 (N_6752,N_2117,N_695);
nand U6753 (N_6753,N_3623,N_1991);
or U6754 (N_6754,N_680,N_757);
nor U6755 (N_6755,N_854,N_1816);
nand U6756 (N_6756,N_3186,N_1031);
nand U6757 (N_6757,N_3862,N_3463);
or U6758 (N_6758,N_1420,N_2994);
nand U6759 (N_6759,N_1716,N_327);
nand U6760 (N_6760,N_1505,N_320);
xnor U6761 (N_6761,N_3773,N_639);
nor U6762 (N_6762,N_126,N_643);
or U6763 (N_6763,N_1001,N_2033);
xor U6764 (N_6764,N_1030,N_1235);
and U6765 (N_6765,N_2610,N_216);
nand U6766 (N_6766,N_3904,N_1708);
xnor U6767 (N_6767,N_2096,N_3572);
xnor U6768 (N_6768,N_551,N_1829);
or U6769 (N_6769,N_2360,N_2670);
nand U6770 (N_6770,N_2103,N_2837);
xnor U6771 (N_6771,N_2108,N_1482);
nand U6772 (N_6772,N_3414,N_3635);
nor U6773 (N_6773,N_373,N_952);
and U6774 (N_6774,N_1740,N_1424);
nor U6775 (N_6775,N_3764,N_269);
nand U6776 (N_6776,N_936,N_76);
and U6777 (N_6777,N_568,N_3879);
nor U6778 (N_6778,N_2545,N_3304);
and U6779 (N_6779,N_1477,N_1697);
nand U6780 (N_6780,N_2489,N_316);
nor U6781 (N_6781,N_3402,N_3885);
and U6782 (N_6782,N_1667,N_463);
xnor U6783 (N_6783,N_2518,N_1165);
nand U6784 (N_6784,N_1732,N_3112);
nor U6785 (N_6785,N_1184,N_1846);
nand U6786 (N_6786,N_3986,N_2232);
and U6787 (N_6787,N_342,N_1206);
and U6788 (N_6788,N_95,N_570);
or U6789 (N_6789,N_237,N_1);
and U6790 (N_6790,N_532,N_1097);
and U6791 (N_6791,N_554,N_1397);
nor U6792 (N_6792,N_53,N_1513);
nand U6793 (N_6793,N_3055,N_2662);
nand U6794 (N_6794,N_2150,N_804);
xor U6795 (N_6795,N_2679,N_2879);
xnor U6796 (N_6796,N_1550,N_1138);
and U6797 (N_6797,N_1072,N_3039);
and U6798 (N_6798,N_887,N_3944);
xnor U6799 (N_6799,N_3195,N_1450);
or U6800 (N_6800,N_857,N_1330);
nand U6801 (N_6801,N_1098,N_814);
or U6802 (N_6802,N_2591,N_1347);
nor U6803 (N_6803,N_3131,N_911);
nor U6804 (N_6804,N_1493,N_1893);
nor U6805 (N_6805,N_3394,N_3416);
or U6806 (N_6806,N_942,N_2204);
and U6807 (N_6807,N_982,N_2387);
nand U6808 (N_6808,N_2627,N_2497);
nand U6809 (N_6809,N_2819,N_3709);
nor U6810 (N_6810,N_1766,N_3897);
or U6811 (N_6811,N_2779,N_1545);
xnor U6812 (N_6812,N_3676,N_1157);
nor U6813 (N_6813,N_3328,N_1436);
nor U6814 (N_6814,N_846,N_3820);
or U6815 (N_6815,N_274,N_3372);
and U6816 (N_6816,N_3298,N_1753);
nand U6817 (N_6817,N_2920,N_3113);
xor U6818 (N_6818,N_3464,N_2807);
or U6819 (N_6819,N_550,N_3842);
nor U6820 (N_6820,N_3146,N_934);
nor U6821 (N_6821,N_2251,N_660);
nor U6822 (N_6822,N_3964,N_1778);
nand U6823 (N_6823,N_1979,N_2837);
nand U6824 (N_6824,N_1650,N_3057);
nand U6825 (N_6825,N_3394,N_1886);
xnor U6826 (N_6826,N_295,N_1258);
or U6827 (N_6827,N_3555,N_3155);
or U6828 (N_6828,N_1917,N_3852);
xnor U6829 (N_6829,N_3605,N_3081);
nor U6830 (N_6830,N_153,N_2619);
xnor U6831 (N_6831,N_2319,N_2524);
nor U6832 (N_6832,N_1559,N_3512);
or U6833 (N_6833,N_3344,N_2971);
nor U6834 (N_6834,N_2063,N_1118);
nand U6835 (N_6835,N_2265,N_1970);
and U6836 (N_6836,N_129,N_2101);
nand U6837 (N_6837,N_42,N_3786);
and U6838 (N_6838,N_2854,N_1916);
nor U6839 (N_6839,N_3260,N_3298);
or U6840 (N_6840,N_3247,N_2598);
nand U6841 (N_6841,N_485,N_1075);
and U6842 (N_6842,N_956,N_1203);
and U6843 (N_6843,N_2669,N_951);
or U6844 (N_6844,N_2388,N_1947);
nor U6845 (N_6845,N_3130,N_1000);
nor U6846 (N_6846,N_1260,N_648);
and U6847 (N_6847,N_2107,N_362);
and U6848 (N_6848,N_2155,N_102);
or U6849 (N_6849,N_2600,N_414);
xnor U6850 (N_6850,N_1940,N_1620);
nor U6851 (N_6851,N_2483,N_1628);
nand U6852 (N_6852,N_2527,N_1907);
nor U6853 (N_6853,N_303,N_3105);
and U6854 (N_6854,N_2702,N_3415);
nand U6855 (N_6855,N_1755,N_3718);
xnor U6856 (N_6856,N_372,N_2040);
nand U6857 (N_6857,N_3080,N_1064);
xnor U6858 (N_6858,N_3393,N_3732);
or U6859 (N_6859,N_499,N_1954);
nor U6860 (N_6860,N_3221,N_1778);
xor U6861 (N_6861,N_170,N_222);
or U6862 (N_6862,N_802,N_3699);
and U6863 (N_6863,N_1083,N_3136);
nand U6864 (N_6864,N_695,N_3026);
nor U6865 (N_6865,N_2564,N_3648);
xnor U6866 (N_6866,N_3261,N_2245);
or U6867 (N_6867,N_3686,N_691);
nand U6868 (N_6868,N_1731,N_196);
or U6869 (N_6869,N_386,N_1393);
nor U6870 (N_6870,N_2425,N_1785);
and U6871 (N_6871,N_365,N_929);
or U6872 (N_6872,N_534,N_1926);
nand U6873 (N_6873,N_1960,N_98);
and U6874 (N_6874,N_2071,N_2761);
nor U6875 (N_6875,N_465,N_3902);
nor U6876 (N_6876,N_2195,N_572);
xor U6877 (N_6877,N_279,N_3915);
nand U6878 (N_6878,N_3048,N_2914);
xnor U6879 (N_6879,N_2950,N_2882);
nand U6880 (N_6880,N_1083,N_876);
xor U6881 (N_6881,N_2560,N_560);
nand U6882 (N_6882,N_843,N_2395);
nor U6883 (N_6883,N_2232,N_3909);
nand U6884 (N_6884,N_1878,N_2404);
xor U6885 (N_6885,N_1188,N_1640);
or U6886 (N_6886,N_323,N_1671);
nand U6887 (N_6887,N_2782,N_2542);
nand U6888 (N_6888,N_3685,N_3430);
nand U6889 (N_6889,N_3646,N_1432);
xor U6890 (N_6890,N_3265,N_2945);
nand U6891 (N_6891,N_3029,N_3953);
nand U6892 (N_6892,N_2046,N_1478);
xnor U6893 (N_6893,N_734,N_3896);
and U6894 (N_6894,N_3289,N_442);
or U6895 (N_6895,N_1778,N_1676);
nand U6896 (N_6896,N_1786,N_734);
or U6897 (N_6897,N_3140,N_2339);
nand U6898 (N_6898,N_950,N_2521);
xnor U6899 (N_6899,N_3239,N_178);
nand U6900 (N_6900,N_3466,N_2757);
xnor U6901 (N_6901,N_305,N_3740);
nand U6902 (N_6902,N_3520,N_2147);
xor U6903 (N_6903,N_230,N_2383);
nor U6904 (N_6904,N_2761,N_2950);
nand U6905 (N_6905,N_493,N_1585);
and U6906 (N_6906,N_3970,N_3810);
and U6907 (N_6907,N_2510,N_2629);
xor U6908 (N_6908,N_580,N_1843);
nand U6909 (N_6909,N_3408,N_3594);
and U6910 (N_6910,N_2012,N_1931);
nand U6911 (N_6911,N_1695,N_360);
nand U6912 (N_6912,N_1469,N_1444);
or U6913 (N_6913,N_1406,N_107);
xor U6914 (N_6914,N_2083,N_1895);
xnor U6915 (N_6915,N_1778,N_1827);
or U6916 (N_6916,N_2320,N_1269);
nor U6917 (N_6917,N_400,N_1845);
or U6918 (N_6918,N_534,N_848);
nand U6919 (N_6919,N_1038,N_2618);
and U6920 (N_6920,N_1689,N_1745);
and U6921 (N_6921,N_3834,N_977);
nor U6922 (N_6922,N_532,N_195);
and U6923 (N_6923,N_3753,N_981);
xor U6924 (N_6924,N_2575,N_3633);
or U6925 (N_6925,N_949,N_3807);
and U6926 (N_6926,N_2474,N_2813);
xnor U6927 (N_6927,N_3706,N_3761);
nand U6928 (N_6928,N_1451,N_1875);
nand U6929 (N_6929,N_3668,N_2998);
nor U6930 (N_6930,N_781,N_2180);
or U6931 (N_6931,N_3552,N_853);
xnor U6932 (N_6932,N_3368,N_2918);
xnor U6933 (N_6933,N_1987,N_2583);
nor U6934 (N_6934,N_3282,N_552);
and U6935 (N_6935,N_631,N_1867);
or U6936 (N_6936,N_244,N_2031);
and U6937 (N_6937,N_1971,N_995);
xnor U6938 (N_6938,N_2956,N_2471);
nor U6939 (N_6939,N_2738,N_746);
nand U6940 (N_6940,N_3283,N_3440);
nor U6941 (N_6941,N_1114,N_2088);
or U6942 (N_6942,N_3961,N_3640);
xnor U6943 (N_6943,N_1785,N_122);
and U6944 (N_6944,N_940,N_525);
xnor U6945 (N_6945,N_1085,N_2816);
nand U6946 (N_6946,N_2655,N_1263);
nor U6947 (N_6947,N_3905,N_3376);
nand U6948 (N_6948,N_664,N_2654);
nor U6949 (N_6949,N_3769,N_2491);
nand U6950 (N_6950,N_3863,N_3461);
xor U6951 (N_6951,N_2506,N_2767);
nor U6952 (N_6952,N_2099,N_2772);
and U6953 (N_6953,N_1222,N_704);
xnor U6954 (N_6954,N_3170,N_2692);
nor U6955 (N_6955,N_3642,N_1491);
nand U6956 (N_6956,N_646,N_2494);
nor U6957 (N_6957,N_2647,N_211);
or U6958 (N_6958,N_3137,N_1769);
xor U6959 (N_6959,N_2368,N_68);
nor U6960 (N_6960,N_2921,N_1382);
nor U6961 (N_6961,N_3632,N_2112);
nor U6962 (N_6962,N_3054,N_2223);
nor U6963 (N_6963,N_3037,N_3415);
nand U6964 (N_6964,N_3719,N_2171);
and U6965 (N_6965,N_3458,N_1549);
nand U6966 (N_6966,N_380,N_13);
nor U6967 (N_6967,N_528,N_1107);
and U6968 (N_6968,N_3916,N_1387);
xor U6969 (N_6969,N_1758,N_619);
or U6970 (N_6970,N_1116,N_2942);
nor U6971 (N_6971,N_1321,N_2381);
nor U6972 (N_6972,N_3305,N_2352);
nand U6973 (N_6973,N_2336,N_186);
nor U6974 (N_6974,N_1772,N_3361);
and U6975 (N_6975,N_3425,N_86);
or U6976 (N_6976,N_2741,N_3510);
and U6977 (N_6977,N_1806,N_467);
nor U6978 (N_6978,N_2783,N_1641);
xnor U6979 (N_6979,N_2229,N_3286);
nand U6980 (N_6980,N_3550,N_394);
nor U6981 (N_6981,N_2463,N_594);
xor U6982 (N_6982,N_1416,N_1548);
xor U6983 (N_6983,N_3414,N_1256);
xor U6984 (N_6984,N_171,N_2976);
and U6985 (N_6985,N_2686,N_3585);
nor U6986 (N_6986,N_3018,N_2264);
xnor U6987 (N_6987,N_736,N_2037);
and U6988 (N_6988,N_1946,N_1548);
xor U6989 (N_6989,N_2717,N_3154);
nand U6990 (N_6990,N_2161,N_3975);
and U6991 (N_6991,N_2288,N_3803);
nor U6992 (N_6992,N_2391,N_2782);
nor U6993 (N_6993,N_732,N_172);
xnor U6994 (N_6994,N_2569,N_2085);
and U6995 (N_6995,N_1834,N_1098);
and U6996 (N_6996,N_593,N_179);
nand U6997 (N_6997,N_1674,N_2152);
nor U6998 (N_6998,N_1249,N_3655);
xnor U6999 (N_6999,N_2741,N_3215);
xnor U7000 (N_7000,N_1933,N_424);
nor U7001 (N_7001,N_2783,N_1199);
and U7002 (N_7002,N_3428,N_3038);
nor U7003 (N_7003,N_3189,N_1273);
or U7004 (N_7004,N_653,N_1383);
and U7005 (N_7005,N_2308,N_2988);
nor U7006 (N_7006,N_3603,N_605);
and U7007 (N_7007,N_1737,N_3045);
or U7008 (N_7008,N_2226,N_2343);
nand U7009 (N_7009,N_2087,N_324);
or U7010 (N_7010,N_1751,N_3282);
xor U7011 (N_7011,N_2653,N_1094);
xor U7012 (N_7012,N_3973,N_3566);
nor U7013 (N_7013,N_3825,N_3519);
or U7014 (N_7014,N_1477,N_2199);
and U7015 (N_7015,N_2104,N_2819);
and U7016 (N_7016,N_507,N_3465);
and U7017 (N_7017,N_2584,N_3141);
xor U7018 (N_7018,N_3957,N_1661);
nor U7019 (N_7019,N_264,N_41);
nor U7020 (N_7020,N_851,N_88);
or U7021 (N_7021,N_2143,N_1996);
nand U7022 (N_7022,N_3764,N_469);
nor U7023 (N_7023,N_2204,N_3662);
or U7024 (N_7024,N_3485,N_1226);
nand U7025 (N_7025,N_606,N_1330);
xnor U7026 (N_7026,N_1736,N_1285);
and U7027 (N_7027,N_2379,N_223);
nor U7028 (N_7028,N_1928,N_2298);
nor U7029 (N_7029,N_410,N_2487);
and U7030 (N_7030,N_1150,N_3144);
nand U7031 (N_7031,N_1091,N_3450);
nand U7032 (N_7032,N_2749,N_2840);
xor U7033 (N_7033,N_2303,N_906);
or U7034 (N_7034,N_732,N_677);
xor U7035 (N_7035,N_710,N_3835);
nor U7036 (N_7036,N_1416,N_3773);
nand U7037 (N_7037,N_3887,N_3290);
nand U7038 (N_7038,N_314,N_2237);
xor U7039 (N_7039,N_3162,N_593);
and U7040 (N_7040,N_2604,N_2086);
nor U7041 (N_7041,N_1826,N_574);
xor U7042 (N_7042,N_1488,N_3484);
or U7043 (N_7043,N_415,N_1349);
xor U7044 (N_7044,N_108,N_2603);
and U7045 (N_7045,N_1595,N_2595);
nor U7046 (N_7046,N_534,N_3798);
nand U7047 (N_7047,N_3623,N_3811);
nand U7048 (N_7048,N_1794,N_1135);
xnor U7049 (N_7049,N_1003,N_1480);
and U7050 (N_7050,N_572,N_866);
and U7051 (N_7051,N_423,N_2881);
nor U7052 (N_7052,N_2119,N_3040);
nand U7053 (N_7053,N_3969,N_3665);
xor U7054 (N_7054,N_2357,N_2345);
xor U7055 (N_7055,N_1527,N_528);
xor U7056 (N_7056,N_3400,N_3067);
xnor U7057 (N_7057,N_2076,N_3939);
and U7058 (N_7058,N_2764,N_3505);
nand U7059 (N_7059,N_2044,N_137);
or U7060 (N_7060,N_195,N_75);
xnor U7061 (N_7061,N_213,N_1496);
nand U7062 (N_7062,N_1558,N_264);
nand U7063 (N_7063,N_3711,N_821);
xor U7064 (N_7064,N_1280,N_3833);
xnor U7065 (N_7065,N_2603,N_2436);
xor U7066 (N_7066,N_74,N_2910);
nand U7067 (N_7067,N_536,N_2017);
nand U7068 (N_7068,N_2681,N_2873);
xor U7069 (N_7069,N_1362,N_60);
nor U7070 (N_7070,N_2612,N_2390);
nor U7071 (N_7071,N_2064,N_1803);
or U7072 (N_7072,N_58,N_1013);
nand U7073 (N_7073,N_3692,N_1837);
and U7074 (N_7074,N_3087,N_1901);
nor U7075 (N_7075,N_127,N_749);
nand U7076 (N_7076,N_2794,N_3820);
or U7077 (N_7077,N_3819,N_2907);
xnor U7078 (N_7078,N_3439,N_1011);
or U7079 (N_7079,N_3664,N_2474);
nor U7080 (N_7080,N_2442,N_1114);
nand U7081 (N_7081,N_420,N_3530);
and U7082 (N_7082,N_1244,N_937);
xnor U7083 (N_7083,N_746,N_1809);
xor U7084 (N_7084,N_1890,N_1869);
nor U7085 (N_7085,N_3884,N_2397);
nor U7086 (N_7086,N_2490,N_1315);
nand U7087 (N_7087,N_2026,N_3121);
or U7088 (N_7088,N_3685,N_2891);
or U7089 (N_7089,N_691,N_3824);
xnor U7090 (N_7090,N_412,N_498);
xor U7091 (N_7091,N_1431,N_153);
xor U7092 (N_7092,N_2491,N_2824);
xnor U7093 (N_7093,N_941,N_2801);
or U7094 (N_7094,N_835,N_1659);
and U7095 (N_7095,N_1369,N_1800);
nor U7096 (N_7096,N_2260,N_876);
and U7097 (N_7097,N_2298,N_215);
nand U7098 (N_7098,N_1493,N_1575);
nor U7099 (N_7099,N_2605,N_2455);
and U7100 (N_7100,N_1249,N_3253);
xor U7101 (N_7101,N_1771,N_194);
nand U7102 (N_7102,N_3701,N_3870);
and U7103 (N_7103,N_650,N_2623);
or U7104 (N_7104,N_3003,N_880);
or U7105 (N_7105,N_3501,N_3116);
and U7106 (N_7106,N_2918,N_1991);
nand U7107 (N_7107,N_3726,N_27);
or U7108 (N_7108,N_114,N_2674);
or U7109 (N_7109,N_2054,N_3367);
nand U7110 (N_7110,N_1070,N_3655);
nor U7111 (N_7111,N_1833,N_810);
nor U7112 (N_7112,N_1625,N_990);
and U7113 (N_7113,N_3015,N_2816);
xor U7114 (N_7114,N_1888,N_2124);
or U7115 (N_7115,N_3827,N_3996);
xor U7116 (N_7116,N_2124,N_1132);
nor U7117 (N_7117,N_1783,N_1743);
nand U7118 (N_7118,N_3192,N_3563);
nand U7119 (N_7119,N_1402,N_261);
and U7120 (N_7120,N_624,N_156);
xor U7121 (N_7121,N_2672,N_780);
nor U7122 (N_7122,N_3698,N_2235);
nor U7123 (N_7123,N_232,N_645);
nor U7124 (N_7124,N_1495,N_761);
nor U7125 (N_7125,N_1168,N_1414);
and U7126 (N_7126,N_3322,N_57);
and U7127 (N_7127,N_1998,N_3383);
or U7128 (N_7128,N_124,N_2429);
and U7129 (N_7129,N_3683,N_2739);
nand U7130 (N_7130,N_3643,N_688);
nor U7131 (N_7131,N_2760,N_3643);
and U7132 (N_7132,N_3595,N_3934);
and U7133 (N_7133,N_38,N_1247);
xor U7134 (N_7134,N_3159,N_1486);
or U7135 (N_7135,N_3,N_2944);
nor U7136 (N_7136,N_1501,N_2903);
nand U7137 (N_7137,N_3508,N_1446);
xnor U7138 (N_7138,N_2472,N_605);
nand U7139 (N_7139,N_3575,N_2113);
and U7140 (N_7140,N_1667,N_60);
or U7141 (N_7141,N_1115,N_2504);
xnor U7142 (N_7142,N_2080,N_3642);
nor U7143 (N_7143,N_2222,N_898);
nor U7144 (N_7144,N_323,N_2322);
or U7145 (N_7145,N_2888,N_1824);
xor U7146 (N_7146,N_3690,N_2538);
nor U7147 (N_7147,N_1053,N_2129);
nor U7148 (N_7148,N_12,N_2129);
nand U7149 (N_7149,N_2617,N_2698);
xor U7150 (N_7150,N_2270,N_1725);
and U7151 (N_7151,N_3731,N_252);
nor U7152 (N_7152,N_1369,N_596);
or U7153 (N_7153,N_2035,N_3092);
nand U7154 (N_7154,N_3889,N_939);
xor U7155 (N_7155,N_3125,N_16);
xnor U7156 (N_7156,N_720,N_316);
xnor U7157 (N_7157,N_2428,N_693);
xor U7158 (N_7158,N_2984,N_3383);
nand U7159 (N_7159,N_2168,N_1103);
or U7160 (N_7160,N_2164,N_1210);
and U7161 (N_7161,N_1804,N_403);
and U7162 (N_7162,N_3327,N_576);
nand U7163 (N_7163,N_2497,N_1576);
xor U7164 (N_7164,N_1516,N_862);
and U7165 (N_7165,N_1917,N_2664);
nor U7166 (N_7166,N_785,N_547);
xor U7167 (N_7167,N_3659,N_951);
and U7168 (N_7168,N_141,N_1363);
nor U7169 (N_7169,N_1333,N_3474);
and U7170 (N_7170,N_3455,N_3609);
xnor U7171 (N_7171,N_2847,N_3801);
and U7172 (N_7172,N_1324,N_2338);
nor U7173 (N_7173,N_3838,N_1829);
nor U7174 (N_7174,N_3,N_1155);
and U7175 (N_7175,N_3400,N_330);
nand U7176 (N_7176,N_3030,N_1631);
xor U7177 (N_7177,N_736,N_681);
or U7178 (N_7178,N_3143,N_884);
xnor U7179 (N_7179,N_1942,N_1037);
nor U7180 (N_7180,N_1949,N_1401);
xnor U7181 (N_7181,N_1081,N_3861);
xnor U7182 (N_7182,N_3346,N_686);
and U7183 (N_7183,N_2496,N_3656);
or U7184 (N_7184,N_75,N_261);
and U7185 (N_7185,N_966,N_1409);
nor U7186 (N_7186,N_3171,N_1790);
xnor U7187 (N_7187,N_1972,N_1593);
or U7188 (N_7188,N_3990,N_1258);
or U7189 (N_7189,N_3178,N_1000);
nand U7190 (N_7190,N_1903,N_3893);
nor U7191 (N_7191,N_1828,N_6);
nor U7192 (N_7192,N_570,N_3135);
and U7193 (N_7193,N_3529,N_126);
nand U7194 (N_7194,N_1529,N_1937);
and U7195 (N_7195,N_2600,N_3899);
and U7196 (N_7196,N_1091,N_2122);
or U7197 (N_7197,N_3783,N_296);
or U7198 (N_7198,N_3921,N_426);
nand U7199 (N_7199,N_639,N_3756);
nand U7200 (N_7200,N_3685,N_1421);
or U7201 (N_7201,N_1835,N_1289);
nand U7202 (N_7202,N_3413,N_1662);
nor U7203 (N_7203,N_454,N_2809);
xor U7204 (N_7204,N_1448,N_2789);
nand U7205 (N_7205,N_758,N_1837);
and U7206 (N_7206,N_125,N_2302);
nor U7207 (N_7207,N_437,N_3670);
and U7208 (N_7208,N_3645,N_727);
nor U7209 (N_7209,N_3911,N_1260);
nor U7210 (N_7210,N_1730,N_921);
xor U7211 (N_7211,N_3361,N_2493);
and U7212 (N_7212,N_1206,N_409);
nor U7213 (N_7213,N_3248,N_2863);
nand U7214 (N_7214,N_392,N_2499);
nand U7215 (N_7215,N_3859,N_583);
nor U7216 (N_7216,N_3945,N_999);
nor U7217 (N_7217,N_3217,N_2137);
nand U7218 (N_7218,N_883,N_600);
xnor U7219 (N_7219,N_807,N_3563);
nor U7220 (N_7220,N_3223,N_3715);
xnor U7221 (N_7221,N_3386,N_3549);
nand U7222 (N_7222,N_1760,N_180);
and U7223 (N_7223,N_513,N_2765);
nand U7224 (N_7224,N_806,N_203);
nand U7225 (N_7225,N_1036,N_1877);
nor U7226 (N_7226,N_1397,N_686);
nor U7227 (N_7227,N_3323,N_3214);
nor U7228 (N_7228,N_1201,N_381);
nand U7229 (N_7229,N_1742,N_2073);
xnor U7230 (N_7230,N_278,N_659);
xnor U7231 (N_7231,N_2966,N_2869);
xnor U7232 (N_7232,N_85,N_737);
nand U7233 (N_7233,N_3961,N_3816);
xnor U7234 (N_7234,N_1690,N_1762);
or U7235 (N_7235,N_958,N_1355);
or U7236 (N_7236,N_807,N_1241);
nor U7237 (N_7237,N_1554,N_2427);
or U7238 (N_7238,N_330,N_2617);
xnor U7239 (N_7239,N_58,N_1621);
nand U7240 (N_7240,N_1106,N_2502);
nand U7241 (N_7241,N_36,N_3268);
xnor U7242 (N_7242,N_3790,N_1773);
nand U7243 (N_7243,N_1424,N_703);
or U7244 (N_7244,N_300,N_3889);
xnor U7245 (N_7245,N_2869,N_1930);
xnor U7246 (N_7246,N_2440,N_1654);
nor U7247 (N_7247,N_2795,N_1060);
xor U7248 (N_7248,N_283,N_2588);
nand U7249 (N_7249,N_2536,N_2921);
nor U7250 (N_7250,N_2200,N_3915);
or U7251 (N_7251,N_951,N_473);
and U7252 (N_7252,N_2633,N_3348);
nand U7253 (N_7253,N_367,N_1021);
nor U7254 (N_7254,N_2132,N_896);
or U7255 (N_7255,N_2076,N_28);
xnor U7256 (N_7256,N_3981,N_1051);
and U7257 (N_7257,N_1364,N_896);
and U7258 (N_7258,N_2971,N_414);
nand U7259 (N_7259,N_1264,N_303);
nand U7260 (N_7260,N_3106,N_3966);
or U7261 (N_7261,N_669,N_2330);
or U7262 (N_7262,N_3121,N_2701);
nor U7263 (N_7263,N_1092,N_818);
nor U7264 (N_7264,N_1520,N_2987);
nor U7265 (N_7265,N_942,N_448);
or U7266 (N_7266,N_2103,N_372);
xnor U7267 (N_7267,N_2447,N_1578);
nor U7268 (N_7268,N_1465,N_3665);
and U7269 (N_7269,N_3846,N_2896);
or U7270 (N_7270,N_3104,N_2719);
and U7271 (N_7271,N_2383,N_2268);
nand U7272 (N_7272,N_1170,N_978);
and U7273 (N_7273,N_2140,N_162);
nand U7274 (N_7274,N_3371,N_102);
nand U7275 (N_7275,N_579,N_3490);
and U7276 (N_7276,N_60,N_1614);
nor U7277 (N_7277,N_3682,N_3071);
nor U7278 (N_7278,N_3535,N_423);
nor U7279 (N_7279,N_3895,N_2103);
or U7280 (N_7280,N_508,N_374);
or U7281 (N_7281,N_826,N_415);
xnor U7282 (N_7282,N_25,N_3963);
or U7283 (N_7283,N_3155,N_1532);
xnor U7284 (N_7284,N_1596,N_3699);
or U7285 (N_7285,N_3666,N_1448);
nand U7286 (N_7286,N_3143,N_878);
and U7287 (N_7287,N_443,N_458);
and U7288 (N_7288,N_3182,N_851);
xor U7289 (N_7289,N_277,N_1441);
or U7290 (N_7290,N_521,N_3744);
nor U7291 (N_7291,N_207,N_827);
xor U7292 (N_7292,N_2987,N_2786);
xnor U7293 (N_7293,N_482,N_2262);
nand U7294 (N_7294,N_3732,N_3319);
and U7295 (N_7295,N_1867,N_2921);
nor U7296 (N_7296,N_1818,N_2724);
and U7297 (N_7297,N_3805,N_3974);
nor U7298 (N_7298,N_3058,N_2757);
and U7299 (N_7299,N_2645,N_3569);
or U7300 (N_7300,N_799,N_2501);
xor U7301 (N_7301,N_2739,N_75);
and U7302 (N_7302,N_2985,N_2069);
and U7303 (N_7303,N_2575,N_861);
nor U7304 (N_7304,N_1049,N_1764);
nor U7305 (N_7305,N_2095,N_3885);
and U7306 (N_7306,N_3132,N_2511);
nand U7307 (N_7307,N_1453,N_3081);
nor U7308 (N_7308,N_15,N_2489);
nor U7309 (N_7309,N_486,N_719);
or U7310 (N_7310,N_3113,N_2585);
nand U7311 (N_7311,N_2658,N_3036);
nand U7312 (N_7312,N_1340,N_2383);
nand U7313 (N_7313,N_3074,N_3564);
or U7314 (N_7314,N_3286,N_2315);
and U7315 (N_7315,N_165,N_288);
nor U7316 (N_7316,N_547,N_1307);
nand U7317 (N_7317,N_583,N_1209);
xor U7318 (N_7318,N_2174,N_2387);
or U7319 (N_7319,N_3907,N_1723);
nand U7320 (N_7320,N_1977,N_1704);
xnor U7321 (N_7321,N_1794,N_3159);
or U7322 (N_7322,N_2164,N_3261);
and U7323 (N_7323,N_2008,N_2957);
xor U7324 (N_7324,N_2147,N_3059);
nor U7325 (N_7325,N_2984,N_3227);
nand U7326 (N_7326,N_3845,N_174);
and U7327 (N_7327,N_2001,N_2880);
nand U7328 (N_7328,N_1727,N_3092);
nor U7329 (N_7329,N_3699,N_790);
or U7330 (N_7330,N_2685,N_3203);
and U7331 (N_7331,N_1325,N_3371);
nor U7332 (N_7332,N_1786,N_482);
xor U7333 (N_7333,N_1833,N_2972);
and U7334 (N_7334,N_1591,N_122);
and U7335 (N_7335,N_2629,N_1131);
and U7336 (N_7336,N_2581,N_3308);
xor U7337 (N_7337,N_708,N_203);
or U7338 (N_7338,N_1029,N_1817);
xnor U7339 (N_7339,N_364,N_1293);
xnor U7340 (N_7340,N_594,N_450);
xor U7341 (N_7341,N_1314,N_2294);
xnor U7342 (N_7342,N_3812,N_2141);
xnor U7343 (N_7343,N_204,N_3684);
nor U7344 (N_7344,N_3957,N_3537);
nand U7345 (N_7345,N_926,N_1306);
xnor U7346 (N_7346,N_3306,N_313);
and U7347 (N_7347,N_11,N_910);
and U7348 (N_7348,N_3887,N_3461);
and U7349 (N_7349,N_808,N_1725);
xor U7350 (N_7350,N_2603,N_305);
and U7351 (N_7351,N_3973,N_1362);
or U7352 (N_7352,N_3639,N_1051);
and U7353 (N_7353,N_841,N_123);
or U7354 (N_7354,N_873,N_1362);
and U7355 (N_7355,N_3256,N_1341);
xor U7356 (N_7356,N_2446,N_2156);
or U7357 (N_7357,N_523,N_2149);
or U7358 (N_7358,N_3487,N_449);
xnor U7359 (N_7359,N_3773,N_1336);
and U7360 (N_7360,N_2832,N_1688);
xor U7361 (N_7361,N_2251,N_3443);
xor U7362 (N_7362,N_804,N_1874);
nor U7363 (N_7363,N_1834,N_1262);
nand U7364 (N_7364,N_2712,N_2669);
nor U7365 (N_7365,N_2454,N_479);
or U7366 (N_7366,N_3557,N_798);
or U7367 (N_7367,N_1392,N_345);
and U7368 (N_7368,N_1855,N_3942);
xnor U7369 (N_7369,N_26,N_1215);
nor U7370 (N_7370,N_3270,N_2166);
nand U7371 (N_7371,N_1456,N_1659);
nor U7372 (N_7372,N_2652,N_1014);
nor U7373 (N_7373,N_1527,N_2374);
or U7374 (N_7374,N_1435,N_1419);
nand U7375 (N_7375,N_1159,N_362);
and U7376 (N_7376,N_3245,N_1881);
xnor U7377 (N_7377,N_936,N_398);
and U7378 (N_7378,N_2292,N_3844);
and U7379 (N_7379,N_913,N_2634);
and U7380 (N_7380,N_2070,N_207);
nor U7381 (N_7381,N_2772,N_1897);
nor U7382 (N_7382,N_614,N_273);
nor U7383 (N_7383,N_3792,N_135);
nor U7384 (N_7384,N_221,N_1357);
xor U7385 (N_7385,N_2829,N_751);
xor U7386 (N_7386,N_2445,N_939);
xnor U7387 (N_7387,N_3818,N_3042);
and U7388 (N_7388,N_661,N_2228);
nor U7389 (N_7389,N_70,N_592);
nand U7390 (N_7390,N_2973,N_2012);
and U7391 (N_7391,N_1863,N_3480);
xor U7392 (N_7392,N_319,N_2790);
xnor U7393 (N_7393,N_1322,N_1358);
and U7394 (N_7394,N_933,N_2438);
nor U7395 (N_7395,N_3738,N_449);
nor U7396 (N_7396,N_1876,N_1301);
xor U7397 (N_7397,N_2831,N_1822);
nand U7398 (N_7398,N_2127,N_2217);
nor U7399 (N_7399,N_952,N_1089);
and U7400 (N_7400,N_3843,N_3907);
and U7401 (N_7401,N_1292,N_3675);
nand U7402 (N_7402,N_1454,N_3109);
nand U7403 (N_7403,N_55,N_1962);
or U7404 (N_7404,N_3473,N_1035);
nand U7405 (N_7405,N_2605,N_3337);
xor U7406 (N_7406,N_565,N_2225);
and U7407 (N_7407,N_2537,N_1310);
and U7408 (N_7408,N_3273,N_3783);
xor U7409 (N_7409,N_2120,N_788);
nor U7410 (N_7410,N_3475,N_3088);
nor U7411 (N_7411,N_2333,N_2676);
nand U7412 (N_7412,N_313,N_1881);
xor U7413 (N_7413,N_162,N_3674);
nand U7414 (N_7414,N_3865,N_3941);
nor U7415 (N_7415,N_2126,N_1849);
and U7416 (N_7416,N_112,N_2865);
or U7417 (N_7417,N_1095,N_190);
xnor U7418 (N_7418,N_681,N_3346);
or U7419 (N_7419,N_802,N_2247);
nand U7420 (N_7420,N_114,N_1652);
or U7421 (N_7421,N_3110,N_2700);
and U7422 (N_7422,N_1240,N_3749);
and U7423 (N_7423,N_976,N_275);
nand U7424 (N_7424,N_950,N_538);
xor U7425 (N_7425,N_2966,N_2381);
and U7426 (N_7426,N_1018,N_159);
nor U7427 (N_7427,N_1694,N_849);
and U7428 (N_7428,N_2089,N_937);
nor U7429 (N_7429,N_3346,N_1420);
and U7430 (N_7430,N_1851,N_3030);
nand U7431 (N_7431,N_1479,N_307);
or U7432 (N_7432,N_611,N_2917);
nand U7433 (N_7433,N_675,N_2961);
or U7434 (N_7434,N_2327,N_1017);
xnor U7435 (N_7435,N_196,N_2905);
xor U7436 (N_7436,N_2893,N_1384);
or U7437 (N_7437,N_2232,N_1571);
nand U7438 (N_7438,N_3275,N_1506);
and U7439 (N_7439,N_236,N_1762);
nor U7440 (N_7440,N_1505,N_1179);
and U7441 (N_7441,N_668,N_859);
or U7442 (N_7442,N_3964,N_3366);
xnor U7443 (N_7443,N_2442,N_3210);
or U7444 (N_7444,N_3742,N_697);
nand U7445 (N_7445,N_2165,N_3334);
xnor U7446 (N_7446,N_2675,N_1746);
nor U7447 (N_7447,N_1511,N_846);
nor U7448 (N_7448,N_3744,N_1885);
xnor U7449 (N_7449,N_1711,N_2451);
xnor U7450 (N_7450,N_3135,N_517);
xor U7451 (N_7451,N_725,N_995);
and U7452 (N_7452,N_1179,N_3892);
nand U7453 (N_7453,N_3339,N_1063);
xnor U7454 (N_7454,N_452,N_1882);
nor U7455 (N_7455,N_369,N_1420);
or U7456 (N_7456,N_3810,N_526);
nand U7457 (N_7457,N_572,N_1938);
and U7458 (N_7458,N_3001,N_1347);
and U7459 (N_7459,N_3584,N_587);
nor U7460 (N_7460,N_497,N_2476);
or U7461 (N_7461,N_855,N_2918);
and U7462 (N_7462,N_147,N_2015);
xor U7463 (N_7463,N_1447,N_2505);
nand U7464 (N_7464,N_1847,N_650);
or U7465 (N_7465,N_3366,N_2914);
and U7466 (N_7466,N_2518,N_469);
and U7467 (N_7467,N_1728,N_1583);
or U7468 (N_7468,N_1319,N_3189);
nor U7469 (N_7469,N_392,N_230);
nand U7470 (N_7470,N_493,N_1911);
nand U7471 (N_7471,N_252,N_1324);
nand U7472 (N_7472,N_2501,N_1424);
xor U7473 (N_7473,N_3592,N_2318);
or U7474 (N_7474,N_3340,N_479);
nand U7475 (N_7475,N_3455,N_117);
xor U7476 (N_7476,N_1654,N_2420);
and U7477 (N_7477,N_3251,N_701);
and U7478 (N_7478,N_2211,N_2835);
and U7479 (N_7479,N_256,N_1996);
nand U7480 (N_7480,N_473,N_1150);
and U7481 (N_7481,N_397,N_3067);
nor U7482 (N_7482,N_3333,N_2952);
or U7483 (N_7483,N_774,N_77);
nor U7484 (N_7484,N_765,N_2040);
nand U7485 (N_7485,N_2125,N_3755);
and U7486 (N_7486,N_3989,N_288);
nand U7487 (N_7487,N_1175,N_1925);
or U7488 (N_7488,N_3259,N_2062);
and U7489 (N_7489,N_1163,N_12);
xnor U7490 (N_7490,N_2822,N_2926);
nand U7491 (N_7491,N_2141,N_1117);
and U7492 (N_7492,N_1369,N_1921);
and U7493 (N_7493,N_1847,N_762);
nor U7494 (N_7494,N_323,N_3250);
and U7495 (N_7495,N_2415,N_1807);
nor U7496 (N_7496,N_1685,N_1561);
nor U7497 (N_7497,N_2913,N_1618);
and U7498 (N_7498,N_3330,N_1578);
and U7499 (N_7499,N_3241,N_432);
nor U7500 (N_7500,N_3568,N_1892);
nor U7501 (N_7501,N_48,N_788);
or U7502 (N_7502,N_3827,N_752);
and U7503 (N_7503,N_3733,N_288);
nor U7504 (N_7504,N_2793,N_3750);
xnor U7505 (N_7505,N_2856,N_3714);
xnor U7506 (N_7506,N_2157,N_631);
and U7507 (N_7507,N_3461,N_919);
and U7508 (N_7508,N_20,N_678);
or U7509 (N_7509,N_1323,N_3879);
nand U7510 (N_7510,N_1655,N_1169);
nand U7511 (N_7511,N_2300,N_2970);
nor U7512 (N_7512,N_1038,N_3375);
xor U7513 (N_7513,N_2717,N_1695);
nand U7514 (N_7514,N_3481,N_1641);
xor U7515 (N_7515,N_2822,N_3080);
and U7516 (N_7516,N_3133,N_3617);
xnor U7517 (N_7517,N_1258,N_3382);
and U7518 (N_7518,N_3617,N_2962);
xor U7519 (N_7519,N_135,N_2494);
xor U7520 (N_7520,N_3830,N_6);
xor U7521 (N_7521,N_1538,N_1213);
nand U7522 (N_7522,N_3374,N_2211);
xnor U7523 (N_7523,N_1996,N_3778);
xnor U7524 (N_7524,N_97,N_663);
nand U7525 (N_7525,N_1136,N_1732);
and U7526 (N_7526,N_1673,N_196);
and U7527 (N_7527,N_3813,N_856);
or U7528 (N_7528,N_942,N_2246);
nand U7529 (N_7529,N_1601,N_610);
and U7530 (N_7530,N_1563,N_2618);
xor U7531 (N_7531,N_3750,N_3502);
or U7532 (N_7532,N_464,N_1073);
nand U7533 (N_7533,N_2612,N_3699);
or U7534 (N_7534,N_1142,N_2985);
or U7535 (N_7535,N_2028,N_1863);
xor U7536 (N_7536,N_2062,N_2350);
xnor U7537 (N_7537,N_2574,N_1245);
xor U7538 (N_7538,N_2712,N_384);
xnor U7539 (N_7539,N_579,N_178);
nor U7540 (N_7540,N_3705,N_1457);
nand U7541 (N_7541,N_2734,N_1068);
nor U7542 (N_7542,N_2179,N_849);
nand U7543 (N_7543,N_407,N_1311);
nand U7544 (N_7544,N_3865,N_3154);
nand U7545 (N_7545,N_2570,N_1500);
or U7546 (N_7546,N_1276,N_2798);
or U7547 (N_7547,N_1359,N_3985);
and U7548 (N_7548,N_3424,N_3574);
xnor U7549 (N_7549,N_399,N_3590);
and U7550 (N_7550,N_1579,N_2677);
and U7551 (N_7551,N_2832,N_3204);
or U7552 (N_7552,N_1920,N_2785);
nor U7553 (N_7553,N_559,N_2770);
xor U7554 (N_7554,N_2827,N_3422);
xnor U7555 (N_7555,N_1570,N_842);
nor U7556 (N_7556,N_1391,N_1991);
or U7557 (N_7557,N_205,N_1856);
or U7558 (N_7558,N_1420,N_2599);
xnor U7559 (N_7559,N_3524,N_3262);
xnor U7560 (N_7560,N_997,N_2378);
and U7561 (N_7561,N_400,N_2410);
or U7562 (N_7562,N_2984,N_2595);
and U7563 (N_7563,N_174,N_717);
xnor U7564 (N_7564,N_253,N_2023);
or U7565 (N_7565,N_1394,N_3553);
or U7566 (N_7566,N_228,N_3926);
nand U7567 (N_7567,N_2671,N_2073);
xnor U7568 (N_7568,N_2612,N_2578);
nand U7569 (N_7569,N_3055,N_1794);
xnor U7570 (N_7570,N_1042,N_892);
nand U7571 (N_7571,N_1773,N_2853);
or U7572 (N_7572,N_3328,N_1335);
nand U7573 (N_7573,N_3686,N_1649);
xnor U7574 (N_7574,N_1103,N_15);
nor U7575 (N_7575,N_1367,N_475);
and U7576 (N_7576,N_2361,N_638);
xnor U7577 (N_7577,N_1013,N_3304);
and U7578 (N_7578,N_3019,N_2473);
nand U7579 (N_7579,N_239,N_1224);
xor U7580 (N_7580,N_3171,N_133);
nand U7581 (N_7581,N_714,N_3592);
or U7582 (N_7582,N_532,N_1258);
nand U7583 (N_7583,N_2007,N_3572);
and U7584 (N_7584,N_744,N_2074);
or U7585 (N_7585,N_3499,N_625);
nor U7586 (N_7586,N_240,N_2826);
nand U7587 (N_7587,N_3279,N_3775);
and U7588 (N_7588,N_2747,N_3324);
and U7589 (N_7589,N_934,N_1544);
and U7590 (N_7590,N_1714,N_338);
or U7591 (N_7591,N_3137,N_2878);
xor U7592 (N_7592,N_2540,N_1235);
nor U7593 (N_7593,N_2627,N_2614);
xnor U7594 (N_7594,N_3746,N_320);
xnor U7595 (N_7595,N_3308,N_1059);
nor U7596 (N_7596,N_841,N_1216);
and U7597 (N_7597,N_3200,N_1697);
nand U7598 (N_7598,N_3582,N_3089);
xor U7599 (N_7599,N_1455,N_1469);
nor U7600 (N_7600,N_2785,N_884);
or U7601 (N_7601,N_2946,N_3338);
and U7602 (N_7602,N_3957,N_999);
and U7603 (N_7603,N_393,N_3629);
nand U7604 (N_7604,N_3003,N_3040);
xnor U7605 (N_7605,N_2086,N_1486);
nor U7606 (N_7606,N_511,N_2143);
nor U7607 (N_7607,N_2432,N_895);
or U7608 (N_7608,N_1110,N_3048);
or U7609 (N_7609,N_1969,N_179);
or U7610 (N_7610,N_372,N_3445);
nor U7611 (N_7611,N_2114,N_1334);
xnor U7612 (N_7612,N_93,N_3026);
nor U7613 (N_7613,N_3637,N_1219);
xor U7614 (N_7614,N_3323,N_3004);
nor U7615 (N_7615,N_2146,N_2596);
or U7616 (N_7616,N_2057,N_2007);
nand U7617 (N_7617,N_1623,N_3793);
or U7618 (N_7618,N_498,N_808);
nand U7619 (N_7619,N_2604,N_376);
or U7620 (N_7620,N_3071,N_1098);
nand U7621 (N_7621,N_891,N_955);
xnor U7622 (N_7622,N_2344,N_1741);
nand U7623 (N_7623,N_2118,N_491);
and U7624 (N_7624,N_3582,N_386);
xor U7625 (N_7625,N_54,N_2821);
nor U7626 (N_7626,N_986,N_3615);
nor U7627 (N_7627,N_529,N_3541);
xnor U7628 (N_7628,N_3837,N_3886);
nor U7629 (N_7629,N_1911,N_3648);
nand U7630 (N_7630,N_2361,N_2686);
xnor U7631 (N_7631,N_3786,N_3905);
and U7632 (N_7632,N_1951,N_195);
xnor U7633 (N_7633,N_2965,N_2119);
xor U7634 (N_7634,N_2942,N_1611);
nand U7635 (N_7635,N_2295,N_3931);
and U7636 (N_7636,N_1629,N_1468);
xnor U7637 (N_7637,N_879,N_3209);
and U7638 (N_7638,N_3641,N_2917);
xnor U7639 (N_7639,N_1649,N_46);
nor U7640 (N_7640,N_1143,N_3313);
nand U7641 (N_7641,N_2218,N_3901);
xnor U7642 (N_7642,N_1025,N_413);
nor U7643 (N_7643,N_1315,N_1917);
nor U7644 (N_7644,N_1941,N_3990);
xor U7645 (N_7645,N_485,N_1707);
nand U7646 (N_7646,N_2498,N_2469);
nor U7647 (N_7647,N_757,N_2763);
nor U7648 (N_7648,N_1716,N_1266);
xor U7649 (N_7649,N_502,N_1595);
nand U7650 (N_7650,N_2030,N_1764);
xor U7651 (N_7651,N_525,N_1713);
nand U7652 (N_7652,N_2613,N_2127);
or U7653 (N_7653,N_631,N_2037);
nor U7654 (N_7654,N_2812,N_2436);
nor U7655 (N_7655,N_2230,N_223);
nand U7656 (N_7656,N_1414,N_2694);
nand U7657 (N_7657,N_2377,N_2722);
or U7658 (N_7658,N_555,N_2358);
nand U7659 (N_7659,N_2862,N_1098);
and U7660 (N_7660,N_3292,N_3980);
or U7661 (N_7661,N_3135,N_535);
xor U7662 (N_7662,N_3202,N_3995);
or U7663 (N_7663,N_983,N_2306);
xnor U7664 (N_7664,N_238,N_2395);
and U7665 (N_7665,N_1346,N_2308);
nand U7666 (N_7666,N_3041,N_3443);
nand U7667 (N_7667,N_1438,N_1561);
nor U7668 (N_7668,N_3686,N_556);
nand U7669 (N_7669,N_2596,N_2024);
nor U7670 (N_7670,N_2201,N_615);
nand U7671 (N_7671,N_3382,N_172);
nor U7672 (N_7672,N_3890,N_691);
nand U7673 (N_7673,N_132,N_1003);
and U7674 (N_7674,N_612,N_1623);
and U7675 (N_7675,N_2292,N_1002);
xnor U7676 (N_7676,N_1135,N_730);
xor U7677 (N_7677,N_1038,N_1885);
nor U7678 (N_7678,N_2470,N_1009);
and U7679 (N_7679,N_1595,N_3239);
xnor U7680 (N_7680,N_576,N_1086);
nor U7681 (N_7681,N_3858,N_1147);
xnor U7682 (N_7682,N_3919,N_187);
nand U7683 (N_7683,N_2392,N_2480);
or U7684 (N_7684,N_3325,N_2118);
and U7685 (N_7685,N_2829,N_2108);
nor U7686 (N_7686,N_1308,N_339);
nor U7687 (N_7687,N_1421,N_3009);
nor U7688 (N_7688,N_2462,N_3642);
and U7689 (N_7689,N_3148,N_1336);
and U7690 (N_7690,N_125,N_2252);
xnor U7691 (N_7691,N_299,N_1443);
nor U7692 (N_7692,N_1315,N_2778);
and U7693 (N_7693,N_3550,N_3852);
and U7694 (N_7694,N_3666,N_562);
and U7695 (N_7695,N_127,N_2191);
nand U7696 (N_7696,N_179,N_1439);
and U7697 (N_7697,N_3218,N_1721);
or U7698 (N_7698,N_783,N_1957);
xor U7699 (N_7699,N_1440,N_3340);
or U7700 (N_7700,N_200,N_2911);
nand U7701 (N_7701,N_1637,N_740);
and U7702 (N_7702,N_832,N_3174);
and U7703 (N_7703,N_3769,N_1968);
or U7704 (N_7704,N_1093,N_3649);
or U7705 (N_7705,N_2940,N_3646);
and U7706 (N_7706,N_2655,N_1665);
and U7707 (N_7707,N_3040,N_1133);
and U7708 (N_7708,N_939,N_2685);
nand U7709 (N_7709,N_366,N_101);
nand U7710 (N_7710,N_985,N_2317);
xor U7711 (N_7711,N_1478,N_3183);
and U7712 (N_7712,N_3298,N_2029);
and U7713 (N_7713,N_1494,N_3734);
xor U7714 (N_7714,N_3309,N_403);
and U7715 (N_7715,N_658,N_3268);
and U7716 (N_7716,N_2367,N_1758);
xor U7717 (N_7717,N_1757,N_1043);
nor U7718 (N_7718,N_3127,N_2716);
xnor U7719 (N_7719,N_2255,N_1806);
or U7720 (N_7720,N_1098,N_2824);
and U7721 (N_7721,N_758,N_15);
nor U7722 (N_7722,N_2492,N_260);
or U7723 (N_7723,N_3508,N_2864);
and U7724 (N_7724,N_2982,N_1367);
nor U7725 (N_7725,N_1565,N_2214);
xor U7726 (N_7726,N_57,N_1922);
and U7727 (N_7727,N_3002,N_3369);
and U7728 (N_7728,N_3449,N_1532);
or U7729 (N_7729,N_1150,N_1967);
xnor U7730 (N_7730,N_3332,N_1);
and U7731 (N_7731,N_3133,N_2124);
nor U7732 (N_7732,N_2804,N_2819);
xnor U7733 (N_7733,N_942,N_3120);
nor U7734 (N_7734,N_1506,N_3446);
and U7735 (N_7735,N_1236,N_1307);
nand U7736 (N_7736,N_1142,N_3338);
xor U7737 (N_7737,N_2946,N_3857);
nor U7738 (N_7738,N_30,N_1137);
or U7739 (N_7739,N_80,N_1744);
and U7740 (N_7740,N_1307,N_2784);
or U7741 (N_7741,N_651,N_3694);
and U7742 (N_7742,N_2827,N_3774);
or U7743 (N_7743,N_1864,N_509);
or U7744 (N_7744,N_1727,N_3070);
nand U7745 (N_7745,N_321,N_174);
xnor U7746 (N_7746,N_3006,N_3866);
nor U7747 (N_7747,N_1238,N_2800);
and U7748 (N_7748,N_1166,N_602);
or U7749 (N_7749,N_1700,N_2581);
nand U7750 (N_7750,N_3333,N_1345);
xor U7751 (N_7751,N_158,N_281);
nor U7752 (N_7752,N_3148,N_1536);
or U7753 (N_7753,N_1606,N_1387);
nor U7754 (N_7754,N_839,N_504);
nand U7755 (N_7755,N_2291,N_3102);
nand U7756 (N_7756,N_168,N_85);
nand U7757 (N_7757,N_144,N_3984);
or U7758 (N_7758,N_2281,N_535);
nor U7759 (N_7759,N_367,N_23);
nor U7760 (N_7760,N_1110,N_806);
or U7761 (N_7761,N_3164,N_1444);
and U7762 (N_7762,N_2362,N_571);
xnor U7763 (N_7763,N_1272,N_2019);
nand U7764 (N_7764,N_3796,N_2068);
or U7765 (N_7765,N_174,N_1458);
nand U7766 (N_7766,N_2083,N_1573);
and U7767 (N_7767,N_897,N_1008);
or U7768 (N_7768,N_1502,N_3808);
nor U7769 (N_7769,N_2758,N_1075);
and U7770 (N_7770,N_605,N_1702);
or U7771 (N_7771,N_3089,N_2149);
nand U7772 (N_7772,N_802,N_2771);
or U7773 (N_7773,N_1786,N_1095);
and U7774 (N_7774,N_531,N_1391);
nor U7775 (N_7775,N_2676,N_636);
and U7776 (N_7776,N_1680,N_2562);
and U7777 (N_7777,N_501,N_1956);
xnor U7778 (N_7778,N_1650,N_707);
nor U7779 (N_7779,N_1431,N_2202);
or U7780 (N_7780,N_2989,N_2395);
nand U7781 (N_7781,N_1073,N_1061);
and U7782 (N_7782,N_1598,N_289);
or U7783 (N_7783,N_3067,N_3076);
or U7784 (N_7784,N_659,N_1385);
nor U7785 (N_7785,N_2325,N_362);
xor U7786 (N_7786,N_3539,N_1545);
nand U7787 (N_7787,N_3220,N_117);
or U7788 (N_7788,N_3556,N_310);
nor U7789 (N_7789,N_996,N_679);
and U7790 (N_7790,N_1413,N_374);
and U7791 (N_7791,N_154,N_1043);
or U7792 (N_7792,N_2043,N_416);
and U7793 (N_7793,N_2389,N_60);
nand U7794 (N_7794,N_223,N_3385);
and U7795 (N_7795,N_491,N_2434);
and U7796 (N_7796,N_2097,N_3247);
nor U7797 (N_7797,N_1933,N_2781);
and U7798 (N_7798,N_1032,N_1529);
or U7799 (N_7799,N_1987,N_1638);
nor U7800 (N_7800,N_3668,N_3739);
or U7801 (N_7801,N_2277,N_147);
and U7802 (N_7802,N_2210,N_1341);
and U7803 (N_7803,N_2769,N_3906);
xor U7804 (N_7804,N_3424,N_3455);
xnor U7805 (N_7805,N_2190,N_1623);
and U7806 (N_7806,N_1215,N_609);
and U7807 (N_7807,N_765,N_1429);
or U7808 (N_7808,N_3626,N_3456);
nor U7809 (N_7809,N_1641,N_3621);
nand U7810 (N_7810,N_802,N_3788);
and U7811 (N_7811,N_1637,N_2321);
nand U7812 (N_7812,N_3119,N_1786);
nor U7813 (N_7813,N_2794,N_3795);
and U7814 (N_7814,N_2294,N_588);
xor U7815 (N_7815,N_1798,N_2150);
nor U7816 (N_7816,N_1132,N_2885);
xnor U7817 (N_7817,N_2832,N_1835);
nand U7818 (N_7818,N_3863,N_1966);
or U7819 (N_7819,N_1154,N_2806);
and U7820 (N_7820,N_2992,N_3511);
or U7821 (N_7821,N_3852,N_2141);
and U7822 (N_7822,N_1554,N_3519);
xnor U7823 (N_7823,N_1834,N_1014);
and U7824 (N_7824,N_2514,N_1791);
and U7825 (N_7825,N_2231,N_727);
nand U7826 (N_7826,N_75,N_1231);
nor U7827 (N_7827,N_2683,N_3287);
nand U7828 (N_7828,N_266,N_1807);
or U7829 (N_7829,N_3660,N_1318);
or U7830 (N_7830,N_2044,N_3255);
and U7831 (N_7831,N_1658,N_2631);
nand U7832 (N_7832,N_1564,N_1952);
xnor U7833 (N_7833,N_1470,N_1843);
nor U7834 (N_7834,N_2416,N_826);
and U7835 (N_7835,N_2772,N_1746);
xor U7836 (N_7836,N_1566,N_2914);
nor U7837 (N_7837,N_524,N_1543);
xor U7838 (N_7838,N_2249,N_2828);
and U7839 (N_7839,N_3228,N_2441);
nor U7840 (N_7840,N_723,N_3812);
nor U7841 (N_7841,N_3660,N_223);
nand U7842 (N_7842,N_3465,N_425);
nor U7843 (N_7843,N_3502,N_2500);
nand U7844 (N_7844,N_2877,N_1352);
xor U7845 (N_7845,N_3541,N_2936);
nor U7846 (N_7846,N_2526,N_2683);
and U7847 (N_7847,N_854,N_1312);
xnor U7848 (N_7848,N_413,N_149);
or U7849 (N_7849,N_1360,N_1990);
xnor U7850 (N_7850,N_863,N_2961);
and U7851 (N_7851,N_2295,N_1055);
xnor U7852 (N_7852,N_208,N_2513);
or U7853 (N_7853,N_886,N_3043);
nor U7854 (N_7854,N_277,N_1059);
xor U7855 (N_7855,N_3963,N_3017);
and U7856 (N_7856,N_276,N_3385);
nand U7857 (N_7857,N_514,N_3566);
and U7858 (N_7858,N_1532,N_407);
and U7859 (N_7859,N_1805,N_26);
and U7860 (N_7860,N_398,N_2032);
nand U7861 (N_7861,N_2933,N_1171);
nor U7862 (N_7862,N_837,N_1624);
nor U7863 (N_7863,N_1830,N_3733);
and U7864 (N_7864,N_2167,N_3092);
xnor U7865 (N_7865,N_3651,N_317);
and U7866 (N_7866,N_3814,N_1583);
or U7867 (N_7867,N_2586,N_1806);
nand U7868 (N_7868,N_912,N_2428);
nand U7869 (N_7869,N_586,N_1441);
nand U7870 (N_7870,N_2466,N_1104);
xor U7871 (N_7871,N_3907,N_1501);
nor U7872 (N_7872,N_1320,N_2327);
or U7873 (N_7873,N_3015,N_3409);
xor U7874 (N_7874,N_3040,N_2389);
nor U7875 (N_7875,N_3284,N_3184);
xor U7876 (N_7876,N_122,N_1526);
xnor U7877 (N_7877,N_2393,N_1725);
nor U7878 (N_7878,N_734,N_930);
xor U7879 (N_7879,N_545,N_2267);
and U7880 (N_7880,N_815,N_3632);
xor U7881 (N_7881,N_2113,N_619);
or U7882 (N_7882,N_3072,N_1514);
and U7883 (N_7883,N_1656,N_2416);
nor U7884 (N_7884,N_1296,N_367);
xnor U7885 (N_7885,N_1804,N_1943);
and U7886 (N_7886,N_3117,N_1792);
nor U7887 (N_7887,N_1457,N_1756);
or U7888 (N_7888,N_2621,N_1498);
or U7889 (N_7889,N_3516,N_3696);
xor U7890 (N_7890,N_3739,N_748);
or U7891 (N_7891,N_2553,N_3478);
or U7892 (N_7892,N_3812,N_2042);
xnor U7893 (N_7893,N_949,N_3880);
or U7894 (N_7894,N_3898,N_3920);
and U7895 (N_7895,N_3834,N_1426);
xor U7896 (N_7896,N_2909,N_3540);
and U7897 (N_7897,N_2120,N_3726);
or U7898 (N_7898,N_2183,N_2901);
and U7899 (N_7899,N_2201,N_1629);
nand U7900 (N_7900,N_628,N_101);
and U7901 (N_7901,N_2474,N_1267);
and U7902 (N_7902,N_368,N_2468);
xor U7903 (N_7903,N_946,N_1672);
nor U7904 (N_7904,N_3276,N_2589);
nor U7905 (N_7905,N_3518,N_370);
nor U7906 (N_7906,N_1066,N_2561);
or U7907 (N_7907,N_1052,N_1334);
xor U7908 (N_7908,N_3155,N_379);
xnor U7909 (N_7909,N_2247,N_3757);
nor U7910 (N_7910,N_1871,N_1298);
xnor U7911 (N_7911,N_1369,N_3380);
xor U7912 (N_7912,N_437,N_3016);
or U7913 (N_7913,N_618,N_216);
nand U7914 (N_7914,N_2934,N_3083);
or U7915 (N_7915,N_1302,N_2501);
or U7916 (N_7916,N_3796,N_3679);
or U7917 (N_7917,N_2802,N_1070);
xor U7918 (N_7918,N_719,N_3760);
xnor U7919 (N_7919,N_3113,N_3375);
xnor U7920 (N_7920,N_1550,N_945);
nand U7921 (N_7921,N_2604,N_2295);
or U7922 (N_7922,N_12,N_1266);
nor U7923 (N_7923,N_1243,N_2422);
xnor U7924 (N_7924,N_116,N_2602);
nand U7925 (N_7925,N_57,N_1141);
nor U7926 (N_7926,N_3492,N_217);
or U7927 (N_7927,N_1118,N_3693);
or U7928 (N_7928,N_1606,N_1448);
nor U7929 (N_7929,N_3489,N_3519);
nor U7930 (N_7930,N_1650,N_868);
nand U7931 (N_7931,N_3935,N_2828);
nand U7932 (N_7932,N_2899,N_1136);
or U7933 (N_7933,N_263,N_257);
nor U7934 (N_7934,N_2785,N_2369);
nor U7935 (N_7935,N_1093,N_3117);
and U7936 (N_7936,N_636,N_1655);
nor U7937 (N_7937,N_156,N_573);
or U7938 (N_7938,N_2116,N_1325);
nand U7939 (N_7939,N_1800,N_1914);
nand U7940 (N_7940,N_959,N_2788);
nand U7941 (N_7941,N_2500,N_3042);
and U7942 (N_7942,N_3798,N_3684);
and U7943 (N_7943,N_2913,N_1497);
nor U7944 (N_7944,N_2133,N_412);
xor U7945 (N_7945,N_2202,N_2132);
nor U7946 (N_7946,N_2131,N_3861);
or U7947 (N_7947,N_68,N_3603);
nand U7948 (N_7948,N_3532,N_1683);
and U7949 (N_7949,N_2674,N_1618);
nand U7950 (N_7950,N_3483,N_3963);
nand U7951 (N_7951,N_789,N_3632);
xor U7952 (N_7952,N_2826,N_510);
nor U7953 (N_7953,N_518,N_3361);
xnor U7954 (N_7954,N_2816,N_1699);
or U7955 (N_7955,N_945,N_3661);
or U7956 (N_7956,N_2881,N_2840);
nor U7957 (N_7957,N_930,N_3529);
nor U7958 (N_7958,N_2593,N_3433);
nor U7959 (N_7959,N_390,N_1878);
or U7960 (N_7960,N_822,N_1872);
nor U7961 (N_7961,N_477,N_2236);
or U7962 (N_7962,N_1457,N_3412);
or U7963 (N_7963,N_1670,N_932);
xnor U7964 (N_7964,N_1633,N_1794);
nor U7965 (N_7965,N_2729,N_1655);
and U7966 (N_7966,N_1219,N_937);
nor U7967 (N_7967,N_3781,N_2611);
nand U7968 (N_7968,N_3894,N_1462);
and U7969 (N_7969,N_295,N_1631);
nor U7970 (N_7970,N_447,N_1794);
xor U7971 (N_7971,N_3402,N_3811);
nor U7972 (N_7972,N_3865,N_1062);
or U7973 (N_7973,N_486,N_1394);
nor U7974 (N_7974,N_724,N_1363);
nand U7975 (N_7975,N_2456,N_2317);
or U7976 (N_7976,N_616,N_1724);
nand U7977 (N_7977,N_1981,N_2014);
and U7978 (N_7978,N_1990,N_2642);
nor U7979 (N_7979,N_555,N_2309);
or U7980 (N_7980,N_1037,N_2172);
xor U7981 (N_7981,N_3957,N_2286);
or U7982 (N_7982,N_3889,N_1267);
nand U7983 (N_7983,N_1746,N_17);
or U7984 (N_7984,N_3352,N_1543);
or U7985 (N_7985,N_1540,N_2581);
and U7986 (N_7986,N_1721,N_482);
xnor U7987 (N_7987,N_3592,N_3755);
nand U7988 (N_7988,N_1706,N_3019);
nor U7989 (N_7989,N_2111,N_1812);
and U7990 (N_7990,N_3150,N_1655);
xor U7991 (N_7991,N_2125,N_1057);
nor U7992 (N_7992,N_2069,N_775);
and U7993 (N_7993,N_2305,N_2081);
xor U7994 (N_7994,N_2307,N_465);
or U7995 (N_7995,N_484,N_13);
or U7996 (N_7996,N_2268,N_2613);
or U7997 (N_7997,N_2174,N_2580);
nor U7998 (N_7998,N_3731,N_2980);
xnor U7999 (N_7999,N_1650,N_109);
or U8000 (N_8000,N_7972,N_6115);
or U8001 (N_8001,N_6116,N_4259);
nor U8002 (N_8002,N_5532,N_7200);
or U8003 (N_8003,N_6831,N_4010);
xor U8004 (N_8004,N_4368,N_5142);
nand U8005 (N_8005,N_7121,N_7273);
xor U8006 (N_8006,N_5274,N_5345);
and U8007 (N_8007,N_5346,N_4646);
nor U8008 (N_8008,N_4763,N_4280);
nor U8009 (N_8009,N_4121,N_5954);
and U8010 (N_8010,N_7058,N_7777);
nor U8011 (N_8011,N_5609,N_6486);
xnor U8012 (N_8012,N_6938,N_7441);
nor U8013 (N_8013,N_6921,N_4752);
and U8014 (N_8014,N_6806,N_7349);
or U8015 (N_8015,N_6519,N_4045);
or U8016 (N_8016,N_5572,N_5215);
xor U8017 (N_8017,N_4793,N_6452);
nor U8018 (N_8018,N_6492,N_6850);
and U8019 (N_8019,N_6458,N_5703);
nor U8020 (N_8020,N_4746,N_4900);
nand U8021 (N_8021,N_7959,N_5307);
and U8022 (N_8022,N_7849,N_7380);
or U8023 (N_8023,N_7540,N_7427);
nand U8024 (N_8024,N_7597,N_5071);
or U8025 (N_8025,N_6509,N_4326);
nand U8026 (N_8026,N_4817,N_7585);
xor U8027 (N_8027,N_6852,N_7339);
and U8028 (N_8028,N_6587,N_6530);
and U8029 (N_8029,N_5129,N_5798);
or U8030 (N_8030,N_6232,N_5728);
nor U8031 (N_8031,N_4771,N_5131);
nand U8032 (N_8032,N_6319,N_5746);
xor U8033 (N_8033,N_6657,N_6900);
xor U8034 (N_8034,N_5789,N_4507);
nor U8035 (N_8035,N_7825,N_6197);
xnor U8036 (N_8036,N_5693,N_7493);
nor U8037 (N_8037,N_4457,N_5642);
and U8038 (N_8038,N_4761,N_5682);
and U8039 (N_8039,N_7030,N_6017);
nor U8040 (N_8040,N_4574,N_7341);
xnor U8041 (N_8041,N_6479,N_5784);
or U8042 (N_8042,N_4160,N_7128);
or U8043 (N_8043,N_7438,N_4783);
and U8044 (N_8044,N_4464,N_4286);
and U8045 (N_8045,N_6392,N_4289);
nor U8046 (N_8046,N_6340,N_7244);
nor U8047 (N_8047,N_5687,N_7281);
and U8048 (N_8048,N_7345,N_4973);
and U8049 (N_8049,N_5880,N_6954);
and U8050 (N_8050,N_6923,N_7462);
nor U8051 (N_8051,N_5821,N_4364);
nand U8052 (N_8052,N_6150,N_5648);
nand U8053 (N_8053,N_4926,N_6446);
or U8054 (N_8054,N_6095,N_5725);
nor U8055 (N_8055,N_6717,N_5440);
nor U8056 (N_8056,N_5390,N_6864);
and U8057 (N_8057,N_5741,N_5143);
and U8058 (N_8058,N_4437,N_4653);
xnor U8059 (N_8059,N_6905,N_4596);
xnor U8060 (N_8060,N_5067,N_4307);
nand U8061 (N_8061,N_7584,N_5810);
nor U8062 (N_8062,N_5596,N_6907);
xnor U8063 (N_8063,N_6410,N_5571);
xnor U8064 (N_8064,N_4863,N_7769);
and U8065 (N_8065,N_6192,N_4684);
nor U8066 (N_8066,N_6825,N_4529);
nand U8067 (N_8067,N_5975,N_4099);
nand U8068 (N_8068,N_5502,N_5630);
and U8069 (N_8069,N_7787,N_5433);
or U8070 (N_8070,N_7811,N_5212);
nand U8071 (N_8071,N_4113,N_7876);
nand U8072 (N_8072,N_5152,N_4577);
and U8073 (N_8073,N_5267,N_7402);
xnor U8074 (N_8074,N_4236,N_7791);
xor U8075 (N_8075,N_5236,N_7542);
or U8076 (N_8076,N_5177,N_4439);
and U8077 (N_8077,N_6840,N_4395);
xor U8078 (N_8078,N_4903,N_7446);
xnor U8079 (N_8079,N_4321,N_7251);
nor U8080 (N_8080,N_5968,N_5332);
and U8081 (N_8081,N_6306,N_4481);
or U8082 (N_8082,N_5047,N_7978);
or U8083 (N_8083,N_6484,N_5251);
or U8084 (N_8084,N_5545,N_6573);
and U8085 (N_8085,N_5221,N_4417);
nor U8086 (N_8086,N_6201,N_6108);
and U8087 (N_8087,N_4140,N_7471);
xor U8088 (N_8088,N_7831,N_6843);
or U8089 (N_8089,N_6280,N_6353);
or U8090 (N_8090,N_6637,N_5624);
and U8091 (N_8091,N_7956,N_6447);
nor U8092 (N_8092,N_6389,N_7814);
and U8093 (N_8093,N_7027,N_4887);
xnor U8094 (N_8094,N_4150,N_5158);
and U8095 (N_8095,N_4130,N_6733);
nand U8096 (N_8096,N_6832,N_5631);
or U8097 (N_8097,N_7476,N_5181);
xor U8098 (N_8098,N_6231,N_7217);
nor U8099 (N_8099,N_4453,N_4965);
nand U8100 (N_8100,N_6415,N_5356);
or U8101 (N_8101,N_7442,N_4060);
nor U8102 (N_8102,N_6411,N_6222);
or U8103 (N_8103,N_5232,N_7136);
nand U8104 (N_8104,N_4301,N_7155);
or U8105 (N_8105,N_7119,N_4686);
xor U8106 (N_8106,N_7163,N_5457);
or U8107 (N_8107,N_6638,N_5077);
nand U8108 (N_8108,N_5781,N_5583);
nand U8109 (N_8109,N_6589,N_4054);
nand U8110 (N_8110,N_4100,N_7731);
and U8111 (N_8111,N_4818,N_4153);
nor U8112 (N_8112,N_6588,N_6069);
or U8113 (N_8113,N_5992,N_5841);
and U8114 (N_8114,N_5849,N_7113);
or U8115 (N_8115,N_5877,N_7756);
nand U8116 (N_8116,N_4908,N_6749);
nor U8117 (N_8117,N_7412,N_4294);
nor U8118 (N_8118,N_5618,N_4603);
or U8119 (N_8119,N_5833,N_5589);
nand U8120 (N_8120,N_6844,N_4943);
and U8121 (N_8121,N_5445,N_4008);
and U8122 (N_8122,N_6024,N_5522);
nand U8123 (N_8123,N_4252,N_5770);
nor U8124 (N_8124,N_7134,N_7377);
nor U8125 (N_8125,N_6285,N_5593);
nor U8126 (N_8126,N_7929,N_4024);
nor U8127 (N_8127,N_7424,N_7620);
and U8128 (N_8128,N_6960,N_7302);
or U8129 (N_8129,N_6799,N_7818);
nor U8130 (N_8130,N_5973,N_5504);
or U8131 (N_8131,N_6033,N_4508);
xnor U8132 (N_8132,N_5917,N_6976);
nand U8133 (N_8133,N_6372,N_5956);
xor U8134 (N_8134,N_6742,N_7259);
xor U8135 (N_8135,N_6768,N_7866);
nand U8136 (N_8136,N_7591,N_6370);
and U8137 (N_8137,N_4569,N_4261);
nand U8138 (N_8138,N_6283,N_7779);
or U8139 (N_8139,N_7486,N_7741);
or U8140 (N_8140,N_6300,N_7903);
or U8141 (N_8141,N_4142,N_4914);
and U8142 (N_8142,N_4734,N_5452);
nor U8143 (N_8143,N_5949,N_4629);
or U8144 (N_8144,N_5681,N_5766);
and U8145 (N_8145,N_5892,N_6350);
nor U8146 (N_8146,N_5520,N_7029);
or U8147 (N_8147,N_7391,N_6711);
nor U8148 (N_8148,N_6896,N_4857);
xor U8149 (N_8149,N_4512,N_6523);
and U8150 (N_8150,N_7108,N_4046);
xor U8151 (N_8151,N_4338,N_6999);
nand U8152 (N_8152,N_6225,N_7025);
nand U8153 (N_8153,N_5004,N_6234);
and U8154 (N_8154,N_4423,N_5438);
and U8155 (N_8155,N_7690,N_7783);
nor U8156 (N_8156,N_6553,N_4936);
nor U8157 (N_8157,N_4541,N_6145);
or U8158 (N_8158,N_4001,N_5016);
or U8159 (N_8159,N_5429,N_7644);
and U8160 (N_8160,N_5931,N_7503);
or U8161 (N_8161,N_6035,N_4249);
or U8162 (N_8162,N_7291,N_5406);
and U8163 (N_8163,N_5832,N_4617);
xor U8164 (N_8164,N_6104,N_7011);
and U8165 (N_8165,N_4768,N_7336);
and U8166 (N_8166,N_7957,N_6468);
nand U8167 (N_8167,N_5434,N_7537);
and U8168 (N_8168,N_6027,N_6105);
and U8169 (N_8169,N_4122,N_5393);
nor U8170 (N_8170,N_5455,N_4089);
and U8171 (N_8171,N_7406,N_5339);
or U8172 (N_8172,N_6379,N_7186);
or U8173 (N_8173,N_7781,N_4604);
or U8174 (N_8174,N_6781,N_4285);
nor U8175 (N_8175,N_4036,N_5573);
xnor U8176 (N_8176,N_4733,N_7374);
xnor U8177 (N_8177,N_6329,N_5189);
nand U8178 (N_8178,N_5132,N_6561);
or U8179 (N_8179,N_5320,N_7151);
and U8180 (N_8180,N_6489,N_7545);
nor U8181 (N_8181,N_7039,N_4867);
or U8182 (N_8182,N_4103,N_6253);
and U8183 (N_8183,N_6526,N_6810);
or U8184 (N_8184,N_7786,N_4850);
and U8185 (N_8185,N_4282,N_6867);
and U8186 (N_8186,N_5400,N_6546);
or U8187 (N_8187,N_4503,N_6780);
or U8188 (N_8188,N_4590,N_7735);
xor U8189 (N_8189,N_7421,N_7041);
or U8190 (N_8190,N_7198,N_7352);
or U8191 (N_8191,N_6516,N_6124);
nor U8192 (N_8192,N_7160,N_6119);
or U8193 (N_8193,N_7414,N_6310);
xor U8194 (N_8194,N_7373,N_5620);
nor U8195 (N_8195,N_7586,N_7673);
xor U8196 (N_8196,N_7677,N_5924);
nand U8197 (N_8197,N_7546,N_4151);
or U8198 (N_8198,N_5122,N_6178);
or U8199 (N_8199,N_7371,N_7082);
or U8200 (N_8200,N_5051,N_4764);
nand U8201 (N_8201,N_6953,N_7533);
and U8202 (N_8202,N_6368,N_6224);
xor U8203 (N_8203,N_7055,N_4921);
xnor U8204 (N_8204,N_4689,N_5021);
nand U8205 (N_8205,N_5603,N_7216);
nand U8206 (N_8206,N_4788,N_5235);
or U8207 (N_8207,N_7842,N_5480);
and U8208 (N_8208,N_4969,N_5328);
and U8209 (N_8209,N_7975,N_7116);
or U8210 (N_8210,N_6209,N_7447);
nand U8211 (N_8211,N_7073,N_4056);
nand U8212 (N_8212,N_7892,N_5319);
nand U8213 (N_8213,N_7871,N_4674);
xnor U8214 (N_8214,N_4913,N_4377);
xor U8215 (N_8215,N_4199,N_7942);
and U8216 (N_8216,N_5028,N_7449);
nor U8217 (N_8217,N_5918,N_7782);
xor U8218 (N_8218,N_7299,N_5903);
xor U8219 (N_8219,N_4539,N_6747);
nor U8220 (N_8220,N_5425,N_5905);
nor U8221 (N_8221,N_6592,N_7410);
nand U8222 (N_8222,N_4071,N_4846);
or U8223 (N_8223,N_7579,N_7875);
nor U8224 (N_8224,N_4677,N_5488);
or U8225 (N_8225,N_6743,N_6063);
and U8226 (N_8226,N_4749,N_6268);
nand U8227 (N_8227,N_4586,N_7289);
or U8228 (N_8228,N_7453,N_5660);
nor U8229 (N_8229,N_7606,N_7989);
and U8230 (N_8230,N_4820,N_5932);
nor U8231 (N_8231,N_7425,N_6291);
and U8232 (N_8232,N_5684,N_4981);
nand U8233 (N_8233,N_4494,N_5839);
nand U8234 (N_8234,N_7515,N_4979);
nand U8235 (N_8235,N_7626,N_5500);
and U8236 (N_8236,N_6414,N_4405);
nand U8237 (N_8237,N_5991,N_6481);
nor U8238 (N_8238,N_7538,N_5835);
nor U8239 (N_8239,N_5173,N_4651);
and U8240 (N_8240,N_6880,N_7277);
nand U8241 (N_8241,N_5707,N_4032);
and U8242 (N_8242,N_4525,N_7665);
nand U8243 (N_8243,N_6435,N_6522);
or U8244 (N_8244,N_4474,N_6075);
xor U8245 (N_8245,N_5848,N_6918);
xnor U8246 (N_8246,N_4889,N_7201);
xnor U8247 (N_8247,N_7640,N_5120);
nor U8248 (N_8248,N_5613,N_7845);
xnor U8249 (N_8249,N_6818,N_5617);
and U8250 (N_8250,N_4445,N_5058);
or U8251 (N_8251,N_7258,N_4354);
xnor U8252 (N_8252,N_7149,N_6514);
nor U8253 (N_8253,N_6330,N_7398);
and U8254 (N_8254,N_7635,N_6791);
nand U8255 (N_8255,N_5408,N_5822);
nand U8256 (N_8256,N_7433,N_4762);
xor U8257 (N_8257,N_4069,N_6014);
xor U8258 (N_8258,N_6972,N_6482);
xor U8259 (N_8259,N_7387,N_6162);
nor U8260 (N_8260,N_5785,N_6821);
nor U8261 (N_8261,N_5426,N_4263);
nand U8262 (N_8262,N_5538,N_4080);
or U8263 (N_8263,N_5579,N_7897);
xnor U8264 (N_8264,N_6412,N_7834);
xnor U8265 (N_8265,N_5601,N_5009);
nand U8266 (N_8266,N_5288,N_5556);
xor U8267 (N_8267,N_6985,N_5898);
and U8268 (N_8268,N_6641,N_4849);
and U8269 (N_8269,N_4030,N_5159);
xnor U8270 (N_8270,N_7556,N_5279);
and U8271 (N_8271,N_7622,N_5943);
nor U8272 (N_8272,N_7507,N_5167);
and U8273 (N_8273,N_4666,N_4509);
or U8274 (N_8274,N_7315,N_5263);
or U8275 (N_8275,N_4422,N_6143);
and U8276 (N_8276,N_4007,N_4801);
and U8277 (N_8277,N_4182,N_7148);
or U8278 (N_8278,N_4465,N_4819);
nor U8279 (N_8279,N_6057,N_4862);
xor U8280 (N_8280,N_7378,N_5727);
and U8281 (N_8281,N_6670,N_4860);
nand U8282 (N_8282,N_7824,N_6173);
or U8283 (N_8283,N_5972,N_4083);
nor U8284 (N_8284,N_5735,N_7409);
nand U8285 (N_8285,N_6451,N_5614);
and U8286 (N_8286,N_4934,N_7212);
or U8287 (N_8287,N_4014,N_6689);
nor U8288 (N_8288,N_5678,N_7706);
xnor U8289 (N_8289,N_5192,N_5729);
xnor U8290 (N_8290,N_4126,N_5944);
nor U8291 (N_8291,N_6182,N_6345);
xor U8292 (N_8292,N_5361,N_5214);
nand U8293 (N_8293,N_5371,N_7571);
or U8294 (N_8294,N_6673,N_6328);
nand U8295 (N_8295,N_6092,N_5790);
xor U8296 (N_8296,N_4524,N_5378);
xnor U8297 (N_8297,N_6973,N_6076);
nand U8298 (N_8298,N_6763,N_6387);
and U8299 (N_8299,N_4949,N_6236);
xor U8300 (N_8300,N_6512,N_6691);
nor U8301 (N_8301,N_5534,N_4984);
nand U8302 (N_8302,N_6333,N_6109);
and U8303 (N_8303,N_4196,N_6501);
nor U8304 (N_8304,N_7682,N_6679);
or U8305 (N_8305,N_4436,N_5278);
xor U8306 (N_8306,N_4971,N_5829);
nand U8307 (N_8307,N_7712,N_7093);
or U8308 (N_8308,N_5064,N_7309);
and U8309 (N_8309,N_4154,N_5777);
nor U8310 (N_8310,N_6254,N_6888);
nand U8311 (N_8311,N_6245,N_5906);
or U8312 (N_8312,N_4661,N_4805);
xor U8313 (N_8313,N_7179,N_5019);
nand U8314 (N_8314,N_7778,N_6440);
xor U8315 (N_8315,N_6674,N_4622);
nor U8316 (N_8316,N_4476,N_6740);
nor U8317 (N_8317,N_6029,N_6114);
or U8318 (N_8318,N_7539,N_5476);
xor U8319 (N_8319,N_7060,N_7973);
and U8320 (N_8320,N_4327,N_7437);
and U8321 (N_8321,N_4898,N_6241);
nand U8322 (N_8322,N_5169,N_4162);
nor U8323 (N_8323,N_5403,N_7173);
or U8324 (N_8324,N_4115,N_5331);
xor U8325 (N_8325,N_6626,N_4579);
nor U8326 (N_8326,N_5748,N_6127);
nor U8327 (N_8327,N_7311,N_6585);
and U8328 (N_8328,N_4425,N_5373);
and U8329 (N_8329,N_6302,N_5869);
nand U8330 (N_8330,N_7314,N_4528);
nor U8331 (N_8331,N_6559,N_7182);
xor U8332 (N_8332,N_5258,N_4206);
xor U8333 (N_8333,N_4462,N_5791);
and U8334 (N_8334,N_5204,N_4595);
or U8335 (N_8335,N_5422,N_5894);
or U8336 (N_8336,N_7900,N_4773);
and U8337 (N_8337,N_4379,N_5333);
nor U8338 (N_8338,N_5138,N_7111);
and U8339 (N_8339,N_7066,N_6431);
and U8340 (N_8340,N_5076,N_7685);
nand U8341 (N_8341,N_6614,N_5118);
and U8342 (N_8342,N_7254,N_5888);
nor U8343 (N_8343,N_7492,N_4953);
and U8344 (N_8344,N_6337,N_4102);
nor U8345 (N_8345,N_7805,N_4255);
nand U8346 (N_8346,N_5222,N_5807);
nor U8347 (N_8347,N_4493,N_4156);
or U8348 (N_8348,N_4808,N_6226);
and U8349 (N_8349,N_4132,N_4696);
or U8350 (N_8350,N_7724,N_5397);
xor U8351 (N_8351,N_7249,N_6453);
nand U8352 (N_8352,N_5809,N_4811);
and U8353 (N_8353,N_4550,N_6212);
nor U8354 (N_8354,N_6243,N_6590);
and U8355 (N_8355,N_5301,N_4697);
xnor U8356 (N_8356,N_6261,N_7906);
nor U8357 (N_8357,N_7560,N_5605);
nand U8358 (N_8358,N_6160,N_5535);
and U8359 (N_8359,N_5084,N_7553);
and U8360 (N_8360,N_6534,N_6753);
nor U8361 (N_8361,N_7949,N_4444);
nand U8362 (N_8362,N_7890,N_7918);
xnor U8363 (N_8363,N_7607,N_5419);
xnor U8364 (N_8364,N_7870,N_6217);
xnor U8365 (N_8365,N_6043,N_5537);
or U8366 (N_8366,N_6205,N_4692);
or U8367 (N_8367,N_6338,N_4598);
or U8368 (N_8368,N_6906,N_6537);
nor U8369 (N_8369,N_6195,N_6172);
xor U8370 (N_8370,N_7867,N_5228);
xor U8371 (N_8371,N_5878,N_7841);
nor U8372 (N_8372,N_6346,N_7970);
xor U8373 (N_8373,N_7687,N_7850);
nand U8374 (N_8374,N_4238,N_7480);
nand U8375 (N_8375,N_6438,N_4429);
and U8376 (N_8376,N_6012,N_5874);
nor U8377 (N_8377,N_6547,N_4918);
nand U8378 (N_8378,N_7836,N_5471);
or U8379 (N_8379,N_5424,N_7645);
or U8380 (N_8380,N_6581,N_4948);
nor U8381 (N_8381,N_4399,N_6171);
nand U8382 (N_8382,N_5806,N_6286);
xor U8383 (N_8383,N_5141,N_6752);
nor U8384 (N_8384,N_4513,N_5135);
and U8385 (N_8385,N_5865,N_6480);
nand U8386 (N_8386,N_4033,N_4624);
nand U8387 (N_8387,N_6180,N_7617);
nor U8388 (N_8388,N_4682,N_5945);
xor U8389 (N_8389,N_4837,N_6085);
xor U8390 (N_8390,N_7381,N_6951);
nor U8391 (N_8391,N_7721,N_4068);
and U8392 (N_8392,N_5310,N_5939);
nand U8393 (N_8393,N_7512,N_6878);
or U8394 (N_8394,N_6500,N_6658);
xnor U8395 (N_8395,N_5704,N_7326);
xor U8396 (N_8396,N_5449,N_7843);
and U8397 (N_8397,N_4814,N_6958);
xnor U8398 (N_8398,N_6683,N_4640);
and U8399 (N_8399,N_4770,N_7117);
or U8400 (N_8400,N_6642,N_4726);
nor U8401 (N_8401,N_5745,N_4005);
and U8402 (N_8402,N_4879,N_4253);
or U8403 (N_8403,N_7941,N_5290);
or U8404 (N_8404,N_6493,N_6255);
nor U8405 (N_8405,N_5011,N_6409);
or U8406 (N_8406,N_5753,N_6282);
nor U8407 (N_8407,N_4662,N_6750);
nand U8408 (N_8408,N_7650,N_6513);
nand U8409 (N_8409,N_5376,N_5626);
xnor U8410 (N_8410,N_7231,N_4145);
and U8411 (N_8411,N_7250,N_7931);
and U8412 (N_8412,N_7361,N_5762);
and U8413 (N_8413,N_7693,N_6853);
xnor U8414 (N_8414,N_7388,N_4028);
or U8415 (N_8415,N_7203,N_6964);
nand U8416 (N_8416,N_4856,N_6375);
nand U8417 (N_8417,N_7698,N_4844);
xnor U8418 (N_8418,N_6230,N_7594);
and U8419 (N_8419,N_4092,N_7142);
nor U8420 (N_8420,N_5099,N_4039);
xnor U8421 (N_8421,N_4774,N_7547);
xnor U8422 (N_8422,N_5533,N_4610);
xor U8423 (N_8423,N_7994,N_7317);
and U8424 (N_8424,N_6246,N_7821);
or U8425 (N_8425,N_4521,N_7732);
or U8426 (N_8426,N_7206,N_5778);
nand U8427 (N_8427,N_7202,N_5531);
and U8428 (N_8428,N_7395,N_4670);
or U8429 (N_8429,N_7404,N_6083);
or U8430 (N_8430,N_4631,N_7616);
nand U8431 (N_8431,N_4348,N_5073);
nand U8432 (N_8432,N_4553,N_6779);
nand U8433 (N_8433,N_4487,N_7432);
or U8434 (N_8434,N_6093,N_4357);
and U8435 (N_8435,N_5742,N_7686);
nor U8436 (N_8436,N_7312,N_4821);
xnor U8437 (N_8437,N_7977,N_5847);
or U8438 (N_8438,N_5767,N_5088);
or U8439 (N_8439,N_7104,N_5639);
nor U8440 (N_8440,N_6814,N_4968);
nor U8441 (N_8441,N_7764,N_7132);
nand U8442 (N_8442,N_6214,N_7268);
or U8443 (N_8443,N_7467,N_5997);
or U8444 (N_8444,N_6407,N_5386);
and U8445 (N_8445,N_6380,N_5416);
nor U8446 (N_8446,N_7727,N_5827);
and U8447 (N_8447,N_5763,N_6727);
or U8448 (N_8448,N_6672,N_6931);
or U8449 (N_8449,N_5870,N_5292);
and U8450 (N_8450,N_7282,N_4623);
nand U8451 (N_8451,N_4823,N_7565);
nand U8452 (N_8452,N_6869,N_4906);
or U8453 (N_8453,N_5559,N_5362);
and U8454 (N_8454,N_4390,N_5552);
and U8455 (N_8455,N_4840,N_5428);
nand U8456 (N_8456,N_7382,N_6003);
and U8457 (N_8457,N_7411,N_7733);
nor U8458 (N_8458,N_5649,N_7710);
nor U8459 (N_8459,N_4011,N_7051);
nand U8460 (N_8460,N_7917,N_5868);
nor U8461 (N_8461,N_5166,N_6998);
or U8462 (N_8462,N_6366,N_7487);
and U8463 (N_8463,N_4125,N_5792);
or U8464 (N_8464,N_6894,N_7817);
and U8465 (N_8465,N_4681,N_6073);
nor U8466 (N_8466,N_4738,N_4048);
nand U8467 (N_8467,N_4530,N_7376);
nand U8468 (N_8468,N_5486,N_7046);
nand U8469 (N_8469,N_4139,N_5038);
nor U8470 (N_8470,N_5760,N_4580);
and U8471 (N_8471,N_6895,N_5585);
xor U8472 (N_8472,N_4871,N_6707);
or U8473 (N_8473,N_5780,N_7468);
or U8474 (N_8474,N_4352,N_5128);
xnor U8475 (N_8475,N_6097,N_7350);
or U8476 (N_8476,N_6554,N_5417);
xor U8477 (N_8477,N_5414,N_7236);
or U8478 (N_8478,N_5484,N_4096);
nand U8479 (N_8479,N_7789,N_4950);
and U8480 (N_8480,N_4776,N_7482);
xnor U8481 (N_8481,N_4363,N_6648);
xnor U8482 (N_8482,N_6422,N_5160);
and U8483 (N_8483,N_7475,N_6576);
nand U8484 (N_8484,N_6483,N_4185);
and U8485 (N_8485,N_4884,N_5238);
nor U8486 (N_8486,N_6577,N_5358);
xnor U8487 (N_8487,N_7122,N_7318);
or U8488 (N_8488,N_5505,N_4495);
nor U8489 (N_8489,N_4594,N_5719);
or U8490 (N_8490,N_4643,N_5819);
nor U8491 (N_8491,N_5330,N_5316);
xnor U8492 (N_8492,N_7489,N_4314);
and U8493 (N_8493,N_7924,N_7103);
or U8494 (N_8494,N_5637,N_7508);
xnor U8495 (N_8495,N_7985,N_5580);
or U8496 (N_8496,N_4518,N_6675);
nor U8497 (N_8497,N_6548,N_4878);
and U8498 (N_8498,N_5269,N_4556);
and U8499 (N_8499,N_7045,N_4864);
xnor U8500 (N_8500,N_4748,N_4777);
nand U8501 (N_8501,N_4227,N_5712);
xnor U8502 (N_8502,N_7750,N_5271);
nor U8503 (N_8503,N_4346,N_5861);
or U8504 (N_8504,N_4833,N_4380);
or U8505 (N_8505,N_7099,N_4313);
nand U8506 (N_8506,N_6847,N_6312);
nand U8507 (N_8507,N_6059,N_7759);
xor U8508 (N_8508,N_5999,N_4794);
nor U8509 (N_8509,N_5942,N_7050);
nor U8510 (N_8510,N_7450,N_6332);
nand U8511 (N_8511,N_6992,N_4165);
nor U8512 (N_8512,N_4345,N_5494);
and U8513 (N_8513,N_4737,N_4567);
and U8514 (N_8514,N_4319,N_6485);
nor U8515 (N_8515,N_4297,N_4627);
and U8516 (N_8516,N_6315,N_7510);
xor U8517 (N_8517,N_4831,N_7997);
xnor U8518 (N_8518,N_6430,N_5926);
xor U8519 (N_8519,N_4107,N_4739);
nor U8520 (N_8520,N_4866,N_7192);
nor U8521 (N_8521,N_6861,N_6690);
and U8522 (N_8522,N_5396,N_6425);
nor U8523 (N_8523,N_6732,N_4891);
and U8524 (N_8524,N_5658,N_5920);
and U8525 (N_8525,N_4460,N_5199);
xnor U8526 (N_8526,N_4907,N_6620);
and U8527 (N_8527,N_4625,N_5680);
nor U8528 (N_8528,N_4939,N_5048);
nor U8529 (N_8529,N_5380,N_5495);
and U8530 (N_8530,N_7573,N_7047);
or U8531 (N_8531,N_5294,N_7551);
and U8532 (N_8532,N_7499,N_7766);
or U8533 (N_8533,N_7223,N_5957);
nand U8534 (N_8534,N_6816,N_5800);
nor U8535 (N_8535,N_4719,N_6363);
nor U8536 (N_8536,N_4491,N_5280);
and U8537 (N_8537,N_6597,N_4786);
nor U8538 (N_8538,N_5871,N_4458);
and U8539 (N_8539,N_4540,N_7008);
or U8540 (N_8540,N_5757,N_7528);
nand U8541 (N_8541,N_5340,N_5750);
and U8542 (N_8542,N_5953,N_7355);
nor U8543 (N_8543,N_5739,N_5659);
xor U8544 (N_8544,N_6562,N_6314);
nor U8545 (N_8545,N_4432,N_7456);
nor U8546 (N_8546,N_6859,N_5402);
xnor U8547 (N_8547,N_7955,N_4482);
xnor U8548 (N_8548,N_7745,N_5555);
and U8549 (N_8549,N_5831,N_7776);
nand U8550 (N_8550,N_7734,N_4229);
and U8551 (N_8551,N_4633,N_5989);
and U8552 (N_8552,N_4469,N_4335);
xor U8553 (N_8553,N_7514,N_4418);
nand U8554 (N_8554,N_4257,N_6174);
nand U8555 (N_8555,N_5628,N_4073);
nand U8556 (N_8556,N_4834,N_5211);
and U8557 (N_8557,N_4652,N_7775);
nor U8558 (N_8558,N_6937,N_6705);
or U8559 (N_8559,N_6714,N_4626);
nand U8560 (N_8560,N_4146,N_4291);
nor U8561 (N_8561,N_4951,N_4003);
and U8562 (N_8562,N_5042,N_5565);
nand U8563 (N_8563,N_4510,N_6560);
xor U8564 (N_8564,N_7641,N_6185);
and U8565 (N_8565,N_5284,N_5706);
or U8566 (N_8566,N_4351,N_5384);
and U8567 (N_8567,N_5577,N_5454);
xnor U8568 (N_8568,N_6018,N_5276);
nor U8569 (N_8569,N_5523,N_4163);
nand U8570 (N_8570,N_6549,N_6406);
nor U8571 (N_8571,N_7102,N_4742);
and U8572 (N_8572,N_4408,N_4964);
nor U8573 (N_8573,N_7637,N_5851);
and U8574 (N_8574,N_6542,N_4720);
nor U8575 (N_8575,N_4273,N_6759);
xnor U8576 (N_8576,N_6729,N_5769);
or U8577 (N_8577,N_4784,N_4987);
and U8578 (N_8578,N_4589,N_5096);
and U8579 (N_8579,N_5788,N_4159);
nand U8580 (N_8580,N_5253,N_5001);
or U8581 (N_8581,N_4672,N_7070);
nor U8582 (N_8582,N_7241,N_5150);
and U8583 (N_8583,N_6849,N_7338);
and U8584 (N_8584,N_7696,N_4004);
and U8585 (N_8585,N_5879,N_7463);
nor U8586 (N_8586,N_7298,N_6404);
and U8587 (N_8587,N_6848,N_7288);
nor U8588 (N_8588,N_4079,N_5959);
nand U8589 (N_8589,N_5635,N_6872);
nand U8590 (N_8590,N_4702,N_4767);
and U8591 (N_8591,N_7502,N_5843);
nor U8592 (N_8592,N_5489,N_5306);
or U8593 (N_8593,N_7519,N_5043);
and U8594 (N_8594,N_5015,N_5491);
and U8595 (N_8595,N_4061,N_4038);
xnor U8596 (N_8596,N_6106,N_7566);
and U8597 (N_8597,N_5799,N_7144);
xnor U8598 (N_8598,N_7129,N_6860);
nor U8599 (N_8599,N_7383,N_5701);
or U8600 (N_8600,N_6772,N_7948);
and U8601 (N_8601,N_6044,N_6434);
nand U8602 (N_8602,N_4358,N_4880);
xnor U8603 (N_8603,N_7943,N_7295);
xor U8604 (N_8604,N_5582,N_4260);
and U8605 (N_8605,N_6833,N_6146);
xnor U8606 (N_8606,N_4452,N_7003);
nand U8607 (N_8607,N_4195,N_5950);
nor U8608 (N_8608,N_6439,N_4403);
nand U8609 (N_8609,N_4299,N_5566);
xor U8610 (N_8610,N_7257,N_4466);
and U8611 (N_8611,N_6868,N_4727);
xor U8612 (N_8612,N_5544,N_4328);
and U8613 (N_8613,N_5890,N_5551);
or U8614 (N_8614,N_4991,N_7146);
nor U8615 (N_8615,N_7497,N_7094);
and U8616 (N_8616,N_6601,N_4367);
nand U8617 (N_8617,N_7334,N_5541);
xnor U8618 (N_8618,N_7195,N_7276);
and U8619 (N_8619,N_6491,N_5529);
or U8620 (N_8620,N_5387,N_5343);
nor U8621 (N_8621,N_4281,N_4179);
nor U8622 (N_8622,N_4781,N_4201);
xor U8623 (N_8623,N_4268,N_4074);
xor U8624 (N_8624,N_4695,N_4219);
nand U8625 (N_8625,N_4087,N_6038);
and U8626 (N_8626,N_7652,N_6432);
nor U8627 (N_8627,N_5960,N_5065);
nand U8628 (N_8628,N_6813,N_7052);
xor U8629 (N_8629,N_4371,N_6563);
and U8630 (N_8630,N_4359,N_6357);
nand U8631 (N_8631,N_5720,N_4051);
and U8632 (N_8632,N_7321,N_6710);
nand U8633 (N_8633,N_7407,N_4873);
xnor U8634 (N_8634,N_7713,N_6339);
and U8635 (N_8635,N_4724,N_4826);
and U8636 (N_8636,N_4999,N_6238);
xor U8637 (N_8637,N_7272,N_7629);
xor U8638 (N_8638,N_5933,N_7472);
xnor U8639 (N_8639,N_5512,N_4416);
nand U8640 (N_8640,N_4955,N_5647);
nand U8641 (N_8641,N_5722,N_6277);
xor U8642 (N_8642,N_6094,N_7840);
xnor U8643 (N_8643,N_6713,N_6567);
nor U8644 (N_8644,N_6600,N_4366);
xor U8645 (N_8645,N_7246,N_5030);
nor U8646 (N_8646,N_7961,N_6256);
or U8647 (N_8647,N_5003,N_6902);
or U8648 (N_8648,N_4447,N_7436);
or U8649 (N_8649,N_5549,N_4757);
nor U8650 (N_8650,N_4571,N_6536);
xnor U8651 (N_8651,N_7718,N_7305);
nand U8652 (N_8652,N_5264,N_7904);
nand U8653 (N_8653,N_7197,N_4435);
nand U8654 (N_8654,N_6071,N_4854);
or U8655 (N_8655,N_7813,N_5367);
nand U8656 (N_8656,N_7634,N_4128);
and U8657 (N_8657,N_7147,N_5510);
nor U8658 (N_8658,N_4736,N_4233);
or U8659 (N_8659,N_6072,N_5059);
and U8660 (N_8660,N_7061,N_6360);
nor U8661 (N_8661,N_6541,N_7385);
nor U8662 (N_8662,N_7920,N_4551);
nand U8663 (N_8663,N_4728,N_7224);
nor U8664 (N_8664,N_4802,N_4218);
nor U8665 (N_8665,N_6531,N_7788);
nand U8666 (N_8666,N_5109,N_6639);
or U8667 (N_8667,N_7426,N_6060);
or U8668 (N_8668,N_6025,N_6386);
xor U8669 (N_8669,N_7853,N_7043);
nor U8670 (N_8670,N_4461,N_6963);
or U8671 (N_8671,N_6148,N_6800);
nor U8672 (N_8672,N_4300,N_6099);
nor U8673 (N_8673,N_5952,N_5104);
nor U8674 (N_8674,N_5130,N_5665);
nor U8675 (N_8675,N_6510,N_6757);
nor U8676 (N_8676,N_6249,N_6532);
or U8677 (N_8677,N_7242,N_4810);
nor U8678 (N_8678,N_4790,N_5176);
or U8679 (N_8679,N_7225,N_6262);
xnor U8680 (N_8680,N_7676,N_5080);
and U8681 (N_8681,N_5242,N_5272);
nor U8682 (N_8682,N_4772,N_5268);
nor U8683 (N_8683,N_7452,N_6219);
nor U8684 (N_8684,N_6702,N_6565);
and U8685 (N_8685,N_4954,N_7575);
nand U8686 (N_8686,N_7264,N_5699);
and U8687 (N_8687,N_5830,N_5977);
and U8688 (N_8688,N_4189,N_7681);
xnor U8689 (N_8689,N_7988,N_5364);
xnor U8690 (N_8690,N_5955,N_5415);
and U8691 (N_8691,N_7987,N_4138);
nand U8692 (N_8692,N_7568,N_6628);
and U8693 (N_8693,N_6260,N_5147);
xnor U8694 (N_8694,N_5289,N_7666);
and U8695 (N_8695,N_5733,N_4133);
nand U8696 (N_8696,N_7928,N_4053);
nor U8697 (N_8697,N_5496,N_7348);
nor U8698 (N_8698,N_7852,N_7632);
xnor U8699 (N_8699,N_4207,N_4334);
nand U8700 (N_8700,N_5646,N_6026);
or U8701 (N_8701,N_5599,N_7598);
and U8702 (N_8702,N_4387,N_4210);
nand U8703 (N_8703,N_7806,N_6009);
xor U8704 (N_8704,N_7974,N_4989);
or U8705 (N_8705,N_5041,N_7614);
nand U8706 (N_8706,N_6369,N_7833);
and U8707 (N_8707,N_4754,N_5156);
nand U8708 (N_8708,N_7754,N_6267);
or U8709 (N_8709,N_6916,N_7075);
xor U8710 (N_8710,N_6013,N_7697);
or U8711 (N_8711,N_4339,N_4016);
nand U8712 (N_8712,N_7026,N_6857);
nand U8713 (N_8713,N_5479,N_6465);
nor U8714 (N_8714,N_6054,N_7561);
nor U8715 (N_8715,N_6804,N_5082);
and U8716 (N_8716,N_4478,N_6946);
xnor U8717 (N_8717,N_6719,N_5857);
and U8718 (N_8718,N_4022,N_7613);
nand U8719 (N_8719,N_6504,N_5721);
and U8720 (N_8720,N_6870,N_6289);
xnor U8721 (N_8721,N_6615,N_4838);
or U8722 (N_8722,N_4373,N_4178);
xnor U8723 (N_8723,N_6052,N_6975);
and U8724 (N_8724,N_6602,N_5442);
nand U8725 (N_8725,N_4824,N_4853);
and U8726 (N_8726,N_6477,N_6000);
xor U8727 (N_8727,N_5468,N_6687);
nor U8728 (N_8728,N_4077,N_7587);
nor U8729 (N_8729,N_4332,N_5163);
nand U8730 (N_8730,N_6792,N_5470);
and U8731 (N_8731,N_4922,N_4193);
nor U8732 (N_8732,N_7835,N_4645);
or U8733 (N_8733,N_7368,N_5695);
nand U8734 (N_8734,N_7984,N_4707);
nor U8735 (N_8735,N_5540,N_5747);
xor U8736 (N_8736,N_4058,N_5094);
nand U8737 (N_8737,N_7098,N_6420);
nand U8738 (N_8738,N_7534,N_7137);
nor U8739 (N_8739,N_5629,N_5348);
nand U8740 (N_8740,N_7222,N_7651);
and U8741 (N_8741,N_5190,N_7408);
xnor U8742 (N_8742,N_4375,N_5187);
nor U8743 (N_8743,N_5350,N_4546);
nor U8744 (N_8744,N_6188,N_6771);
and U8745 (N_8745,N_6331,N_7164);
nor U8746 (N_8746,N_5431,N_5550);
and U8747 (N_8747,N_7874,N_4740);
nand U8748 (N_8748,N_4975,N_5341);
or U8749 (N_8749,N_7602,N_7214);
xnor U8750 (N_8750,N_7028,N_7396);
nand U8751 (N_8751,N_4455,N_7705);
and U8752 (N_8752,N_5916,N_7319);
and U8753 (N_8753,N_6004,N_7112);
or U8754 (N_8754,N_6656,N_7909);
nand U8755 (N_8755,N_5490,N_5446);
or U8756 (N_8756,N_7347,N_5186);
and U8757 (N_8757,N_7877,N_6616);
and U8758 (N_8758,N_5247,N_5909);
or U8759 (N_8759,N_5095,N_4192);
nand U8760 (N_8760,N_5401,N_5194);
and U8761 (N_8761,N_5074,N_6227);
or U8762 (N_8762,N_7523,N_4209);
or U8763 (N_8763,N_4075,N_4632);
xor U8764 (N_8764,N_5149,N_5574);
nor U8765 (N_8765,N_5964,N_7496);
xor U8766 (N_8766,N_5309,N_6031);
nand U8767 (N_8767,N_5666,N_5698);
nand U8768 (N_8768,N_4269,N_6889);
or U8769 (N_8769,N_6845,N_7765);
and U8770 (N_8770,N_5893,N_4519);
or U8771 (N_8771,N_4655,N_4224);
or U8772 (N_8772,N_6866,N_4688);
xnor U8773 (N_8773,N_6962,N_6264);
nand U8774 (N_8774,N_7726,N_6275);
or U8775 (N_8775,N_5499,N_5007);
and U8776 (N_8776,N_4657,N_6700);
or U8777 (N_8777,N_4944,N_4886);
nand U8778 (N_8778,N_4349,N_4374);
xor U8779 (N_8779,N_4713,N_4822);
nor U8780 (N_8780,N_5255,N_7921);
xor U8781 (N_8781,N_5102,N_4607);
nor U8782 (N_8782,N_5126,N_4996);
xnor U8783 (N_8783,N_7976,N_7701);
nand U8784 (N_8784,N_7991,N_7770);
nand U8785 (N_8785,N_5022,N_6274);
or U8786 (N_8786,N_5846,N_5394);
and U8787 (N_8787,N_7580,N_7552);
and U8788 (N_8788,N_6997,N_5243);
and U8789 (N_8789,N_5363,N_7807);
xor U8790 (N_8790,N_5040,N_4526);
nor U8791 (N_8791,N_7185,N_4490);
or U8792 (N_8792,N_6391,N_6478);
nor U8793 (N_8793,N_7287,N_7695);
nor U8794 (N_8794,N_6540,N_7086);
xnor U8795 (N_8795,N_5370,N_6873);
nor U8796 (N_8796,N_6764,N_7278);
nor U8797 (N_8797,N_5899,N_5518);
or U8798 (N_8798,N_5196,N_5157);
and U8799 (N_8799,N_7359,N_6296);
nor U8800 (N_8800,N_7979,N_6163);
or U8801 (N_8801,N_5453,N_6745);
nand U8802 (N_8802,N_7068,N_4155);
nand U8803 (N_8803,N_6834,N_6604);
xor U8804 (N_8804,N_7544,N_7969);
or U8805 (N_8805,N_7459,N_5420);
nor U8806 (N_8806,N_6910,N_6726);
or U8807 (N_8807,N_5718,N_7369);
nor U8808 (N_8808,N_5413,N_4500);
nand U8809 (N_8809,N_6882,N_4111);
nor U8810 (N_8810,N_7458,N_5776);
nor U8811 (N_8811,N_7667,N_5165);
or U8812 (N_8812,N_4769,N_5590);
or U8813 (N_8813,N_7430,N_7760);
or U8814 (N_8814,N_7394,N_4205);
nand U8815 (N_8815,N_5842,N_5312);
nand U8816 (N_8816,N_7416,N_5575);
or U8817 (N_8817,N_6395,N_6736);
nand U8818 (N_8818,N_6318,N_5210);
and U8819 (N_8819,N_6394,N_7945);
or U8820 (N_8820,N_4892,N_4573);
nand U8821 (N_8821,N_4803,N_7501);
nand U8822 (N_8822,N_7367,N_7280);
xnor U8823 (N_8823,N_6881,N_6239);
nand U8824 (N_8824,N_7596,N_7772);
and U8825 (N_8825,N_7190,N_6704);
xnor U8826 (N_8826,N_7996,N_7797);
nand U8827 (N_8827,N_4941,N_5927);
or U8828 (N_8828,N_4029,N_6661);
xnor U8829 (N_8829,N_4705,N_4475);
or U8830 (N_8830,N_5245,N_5653);
nor U8831 (N_8831,N_7101,N_6293);
or U8832 (N_8832,N_7882,N_4221);
and U8833 (N_8833,N_6001,N_7608);
xor U8834 (N_8834,N_6457,N_5297);
xor U8835 (N_8835,N_6950,N_4843);
xnor U8836 (N_8836,N_7191,N_7729);
and U8837 (N_8837,N_6049,N_4861);
nor U8838 (N_8838,N_5473,N_4109);
xor U8839 (N_8839,N_6098,N_5127);
or U8840 (N_8840,N_6778,N_4483);
nor U8841 (N_8841,N_5325,N_4414);
or U8842 (N_8842,N_7153,N_5709);
and U8843 (N_8843,N_4020,N_4897);
nor U8844 (N_8844,N_6237,N_6100);
nor U8845 (N_8845,N_4599,N_5930);
and U8846 (N_8846,N_4082,N_7260);
xor U8847 (N_8847,N_4434,N_6987);
nand U8848 (N_8848,N_6139,N_6662);
xor U8849 (N_8849,N_4568,N_4064);
or U8850 (N_8850,N_7196,N_7124);
and U8851 (N_8851,N_5825,N_6824);
or U8852 (N_8852,N_7166,N_5225);
nor U8853 (N_8853,N_6258,N_6064);
and U8854 (N_8854,N_5281,N_5570);
xnor U8855 (N_8855,N_7513,N_7823);
nand U8856 (N_8856,N_6203,N_4591);
nor U8857 (N_8857,N_6417,N_5023);
nor U8858 (N_8858,N_4040,N_7018);
or U8859 (N_8859,N_4059,N_5482);
or U8860 (N_8860,N_6159,N_6367);
xor U8861 (N_8861,N_4127,N_7680);
and U8862 (N_8862,N_5090,N_4527);
xnor U8863 (N_8863,N_7563,N_6944);
and U8864 (N_8864,N_6462,N_7630);
and U8865 (N_8865,N_7504,N_4894);
and U8866 (N_8866,N_7106,N_7554);
and U8867 (N_8867,N_5661,N_4468);
nor U8868 (N_8868,N_6475,N_7951);
xor U8869 (N_8869,N_4638,N_5114);
and U8870 (N_8870,N_7576,N_5481);
xor U8871 (N_8871,N_6659,N_6444);
and U8872 (N_8872,N_5702,N_6487);
nor U8873 (N_8873,N_4741,N_5435);
xor U8874 (N_8874,N_6879,N_6157);
or U8875 (N_8875,N_6045,N_6494);
and U8876 (N_8876,N_4441,N_6079);
or U8877 (N_8877,N_4882,N_7485);
nor U8878 (N_8878,N_6041,N_6908);
nand U8879 (N_8879,N_5257,N_7744);
nand U8880 (N_8880,N_4310,N_5717);
nand U8881 (N_8881,N_5093,N_7572);
xor U8882 (N_8882,N_6011,N_6361);
or U8883 (N_8883,N_5111,N_5322);
or U8884 (N_8884,N_6966,N_5070);
nor U8885 (N_8885,N_6161,N_5811);
nor U8886 (N_8886,N_6968,N_6647);
nand U8887 (N_8887,N_6826,N_6917);
xor U8888 (N_8888,N_5285,N_7638);
and U8889 (N_8889,N_7627,N_4830);
nor U8890 (N_8890,N_5560,N_4890);
xor U8891 (N_8891,N_6584,N_5056);
xor U8892 (N_8892,N_7656,N_5398);
xor U8893 (N_8893,N_6979,N_5947);
or U8894 (N_8894,N_5239,N_4129);
nand U8895 (N_8895,N_6718,N_6077);
nand U8896 (N_8896,N_6943,N_7455);
nor U8897 (N_8897,N_6456,N_6785);
and U8898 (N_8898,N_5864,N_5828);
and U8899 (N_8899,N_4909,N_6955);
nand U8900 (N_8900,N_4945,N_4656);
nand U8901 (N_8901,N_4967,N_5881);
and U8902 (N_8902,N_6047,N_6884);
nor U8903 (N_8903,N_6218,N_5086);
nor U8904 (N_8904,N_6582,N_6272);
or U8905 (N_8905,N_5774,N_7323);
nand U8906 (N_8906,N_5671,N_5794);
xor U8907 (N_8907,N_6575,N_6754);
xor U8908 (N_8908,N_7530,N_6067);
nor U8909 (N_8909,N_7982,N_6508);
nor U8910 (N_8910,N_7992,N_5318);
xor U8911 (N_8911,N_4232,N_4497);
or U8912 (N_8912,N_4472,N_5010);
nand U8913 (N_8913,N_5336,N_7327);
xnor U8914 (N_8914,N_6206,N_7708);
nand U8915 (N_8915,N_7663,N_6942);
xnor U8916 (N_8916,N_6930,N_5226);
xnor U8917 (N_8917,N_5388,N_4424);
nor U8918 (N_8918,N_5463,N_6460);
or U8919 (N_8919,N_7854,N_6805);
nor U8920 (N_8920,N_5636,N_7465);
nand U8921 (N_8921,N_6716,N_4078);
nor U8922 (N_8922,N_5994,N_4176);
or U8923 (N_8923,N_7157,N_4584);
and U8924 (N_8924,N_6819,N_7518);
nor U8925 (N_8925,N_7054,N_4295);
nor U8926 (N_8926,N_5664,N_5081);
nor U8927 (N_8927,N_5850,N_4614);
nand U8928 (N_8928,N_4729,N_4683);
nand U8929 (N_8929,N_5304,N_5405);
and U8930 (N_8930,N_4386,N_7156);
nor U8931 (N_8931,N_6915,N_7839);
xnor U8932 (N_8932,N_5731,N_7154);
or U8933 (N_8933,N_6087,N_4049);
nand U8934 (N_8934,N_7418,N_4164);
and U8935 (N_8935,N_4315,N_7080);
nand U8936 (N_8936,N_7832,N_6154);
nand U8937 (N_8937,N_6952,N_5385);
xor U8938 (N_8938,N_5548,N_7859);
nand U8939 (N_8939,N_7922,N_6823);
or U8940 (N_8940,N_7474,N_7810);
and U8941 (N_8941,N_5524,N_5853);
nand U8942 (N_8942,N_5134,N_4203);
nor U8943 (N_8943,N_6595,N_5123);
xor U8944 (N_8944,N_4501,N_6359);
nor U8945 (N_8945,N_5327,N_7059);
nand U8946 (N_8946,N_6798,N_4438);
or U8947 (N_8947,N_4874,N_5293);
and U8948 (N_8948,N_4093,N_6887);
and U8949 (N_8949,N_6746,N_4549);
xor U8950 (N_8950,N_5818,N_4533);
nand U8951 (N_8951,N_4636,N_5752);
and U8952 (N_8952,N_5690,N_4480);
and U8953 (N_8953,N_4166,N_6603);
nand U8954 (N_8954,N_7033,N_5514);
nand U8955 (N_8955,N_6039,N_7133);
xnor U8956 (N_8956,N_4852,N_6470);
or U8957 (N_8957,N_4718,N_4026);
and U8958 (N_8958,N_4559,N_4402);
xnor U8959 (N_8959,N_5816,N_7654);
xnor U8960 (N_8960,N_4583,N_4241);
nand U8961 (N_8961,N_7592,N_5600);
or U8962 (N_8962,N_4184,N_6594);
or U8963 (N_8963,N_4383,N_6802);
nand U8964 (N_8964,N_5887,N_5813);
xor U8965 (N_8965,N_4148,N_4267);
and U8966 (N_8966,N_5317,N_7550);
nor U8967 (N_8967,N_4063,N_6912);
and U8968 (N_8968,N_6686,N_7329);
and U8969 (N_8969,N_7590,N_5795);
nor U8970 (N_8970,N_6397,N_5513);
nor U8971 (N_8971,N_5277,N_7934);
or U8972 (N_8972,N_4311,N_4406);
or U8973 (N_8973,N_6741,N_4756);
nor U8974 (N_8974,N_4169,N_6418);
xnor U8975 (N_8975,N_5014,N_5911);
and U8976 (N_8976,N_4714,N_5458);
nor U8977 (N_8977,N_6934,N_4023);
nor U8978 (N_8978,N_6220,N_6803);
xnor U8979 (N_8979,N_5133,N_7885);
nor U8980 (N_8980,N_6605,N_6552);
or U8981 (N_8981,N_5965,N_6898);
nand U8982 (N_8982,N_6544,N_7443);
nor U8983 (N_8983,N_7230,N_7484);
nor U8984 (N_8984,N_4194,N_6539);
or U8985 (N_8985,N_5961,N_4186);
xnor U8986 (N_8986,N_7199,N_7393);
and U8987 (N_8987,N_6619,N_5501);
or U8988 (N_8988,N_7506,N_4234);
or U8989 (N_8989,N_5754,N_6737);
nor U8990 (N_8990,N_5802,N_6187);
nor U8991 (N_8991,N_5657,N_5516);
nor U8992 (N_8992,N_7531,N_6735);
nand U8993 (N_8993,N_7858,N_5467);
nand U8994 (N_8994,N_5797,N_6455);
or U8995 (N_8995,N_6762,N_5112);
or U8996 (N_8996,N_4613,N_6211);
and U8997 (N_8997,N_4701,N_7965);
nand U8998 (N_8998,N_7095,N_5592);
and U8999 (N_8999,N_7076,N_7228);
nand U9000 (N_9000,N_4735,N_5025);
and U9001 (N_9001,N_7847,N_5808);
nor U9002 (N_9002,N_4881,N_5775);
nor U9003 (N_9003,N_4095,N_7234);
nor U9004 (N_9004,N_5528,N_4993);
nand U9005 (N_9005,N_5044,N_7748);
nand U9006 (N_9006,N_7187,N_4928);
nand U9007 (N_9007,N_5498,N_6617);
nor U9008 (N_9008,N_4198,N_7403);
nand U9009 (N_9009,N_6070,N_7653);
nand U9010 (N_9010,N_5672,N_4994);
xnor U9011 (N_9011,N_5732,N_5714);
nor U9012 (N_9012,N_5539,N_5652);
nand U9013 (N_9013,N_5303,N_6307);
xor U9014 (N_9014,N_6935,N_6257);
xor U9015 (N_9015,N_6699,N_6273);
or U9016 (N_9016,N_6967,N_6671);
xor U9017 (N_9017,N_5667,N_7891);
or U9018 (N_9018,N_4101,N_5213);
nand U9019 (N_9019,N_4202,N_5683);
nand U9020 (N_9020,N_7963,N_4393);
and U9021 (N_9021,N_6933,N_4572);
nand U9022 (N_9022,N_6053,N_5436);
xor U9023 (N_9023,N_7535,N_6789);
nor U9024 (N_9024,N_6533,N_6362);
nand U9025 (N_9025,N_4911,N_7183);
nand U9026 (N_9026,N_5670,N_6820);
xnor U9027 (N_9027,N_6684,N_6939);
and U9028 (N_9028,N_6466,N_4809);
or U9029 (N_9029,N_6215,N_6876);
or U9030 (N_9030,N_5103,N_7007);
xnor U9031 (N_9031,N_6538,N_5198);
xnor U9032 (N_9032,N_7266,N_6278);
nor U9033 (N_9033,N_7822,N_4065);
and U9034 (N_9034,N_5354,N_5066);
and U9035 (N_9035,N_7601,N_5858);
and U9036 (N_9036,N_4340,N_5078);
or U9037 (N_9037,N_5308,N_4963);
xnor U9038 (N_9038,N_5561,N_6189);
and U9039 (N_9039,N_5772,N_4717);
nor U9040 (N_9040,N_6551,N_4516);
nor U9041 (N_9041,N_6334,N_6680);
nor U9042 (N_9042,N_5241,N_4904);
or U9043 (N_9043,N_7844,N_5761);
xnor U9044 (N_9044,N_7354,N_7032);
nand U9045 (N_9045,N_7658,N_5115);
xnor U9046 (N_9046,N_4356,N_5979);
or U9047 (N_9047,N_7802,N_6995);
or U9048 (N_9048,N_7077,N_4715);
nor U9049 (N_9049,N_7524,N_5430);
nor U9050 (N_9050,N_5632,N_6767);
and U9051 (N_9051,N_7703,N_4899);
nor U9052 (N_9052,N_4247,N_5153);
nor U9053 (N_9053,N_5368,N_5723);
and U9054 (N_9054,N_7364,N_4985);
xnor U9055 (N_9055,N_6932,N_5674);
and U9056 (N_9056,N_4404,N_7647);
and U9057 (N_9057,N_7846,N_5355);
or U9058 (N_9058,N_6202,N_7574);
xor U9059 (N_9059,N_4242,N_5352);
and U9060 (N_9060,N_4961,N_4245);
nand U9061 (N_9061,N_7263,N_4034);
and U9062 (N_9062,N_6751,N_5404);
nor U9063 (N_9063,N_5377,N_7660);
nand U9064 (N_9064,N_7328,N_5908);
and U9065 (N_9065,N_6517,N_5324);
nor U9066 (N_9066,N_5033,N_6660);
nor U9067 (N_9067,N_6893,N_7356);
and U9068 (N_9068,N_7603,N_7274);
xnor U9069 (N_9069,N_7386,N_5223);
nand U9070 (N_9070,N_5738,N_5602);
xnor U9071 (N_9071,N_7362,N_5759);
xor U9072 (N_9072,N_5820,N_5606);
and U9073 (N_9073,N_5493,N_5527);
nand U9074 (N_9074,N_7953,N_5969);
xor U9075 (N_9075,N_4977,N_7088);
and U9076 (N_9076,N_5995,N_5526);
nor U9077 (N_9077,N_7761,N_4489);
nand U9078 (N_9078,N_7999,N_7527);
nor U9079 (N_9079,N_6665,N_6006);
xor U9080 (N_9080,N_7252,N_6472);
and U9081 (N_9081,N_6429,N_6290);
nand U9082 (N_9082,N_4585,N_7588);
nor U9083 (N_9083,N_4277,N_5013);
xor U9084 (N_9084,N_4035,N_4330);
nand U9085 (N_9085,N_6204,N_5768);
xor U9086 (N_9086,N_6121,N_5910);
nor U9087 (N_9087,N_7100,N_4308);
and U9088 (N_9088,N_7351,N_5338);
and U9089 (N_9089,N_6940,N_7000);
xor U9090 (N_9090,N_4916,N_5347);
or U9091 (N_9091,N_5202,N_7946);
nor U9092 (N_9092,N_6388,N_7020);
xnor U9093 (N_9093,N_7239,N_7429);
xor U9094 (N_9094,N_5940,N_4070);
nand U9095 (N_9095,N_7564,N_7063);
nand U9096 (N_9096,N_4935,N_5451);
or U9097 (N_9097,N_6040,N_7930);
xor U9098 (N_9098,N_6356,N_5576);
nor U9099 (N_9099,N_5530,N_6364);
or U9100 (N_9100,N_6048,N_7010);
nor U9101 (N_9101,N_4498,N_7017);
or U9102 (N_9102,N_5922,N_5359);
xnor U9103 (N_9103,N_5483,N_7469);
nor U9104 (N_9104,N_6142,N_7420);
xor U9105 (N_9105,N_7646,N_6488);
nand U9106 (N_9106,N_4215,N_7722);
nand U9107 (N_9107,N_6168,N_4396);
and U9108 (N_9108,N_7912,N_4216);
nor U9109 (N_9109,N_5688,N_4391);
or U9110 (N_9110,N_4105,N_4650);
nor U9111 (N_9111,N_6496,N_7505);
and U9112 (N_9112,N_6766,N_7078);
and U9113 (N_9113,N_7886,N_6983);
or U9114 (N_9114,N_5907,N_6287);
nor U9115 (N_9115,N_7773,N_4828);
or U9116 (N_9116,N_7332,N_4047);
nor U9117 (N_9117,N_5946,N_4256);
xor U9118 (N_9118,N_5963,N_4350);
nor U9119 (N_9119,N_6636,N_6593);
nor U9120 (N_9120,N_4804,N_7998);
or U9121 (N_9121,N_7589,N_5587);
or U9122 (N_9122,N_5543,N_6507);
or U9123 (N_9123,N_7445,N_5383);
nor U9124 (N_9124,N_5349,N_7618);
and U9125 (N_9125,N_7643,N_7838);
and U9126 (N_9126,N_5389,N_6107);
nor U9127 (N_9127,N_5921,N_5478);
nor U9128 (N_9128,N_4620,N_4431);
nand U9129 (N_9129,N_6155,N_7784);
and U9130 (N_9130,N_4384,N_4982);
or U9131 (N_9131,N_6897,N_6010);
and U9132 (N_9132,N_4937,N_6811);
xnor U9133 (N_9133,N_6579,N_7019);
nor U9134 (N_9134,N_7375,N_6126);
and U9135 (N_9135,N_5117,N_7700);
or U9136 (N_9136,N_5634,N_7555);
nand U9137 (N_9137,N_5008,N_7152);
nor U9138 (N_9138,N_4118,N_5554);
nor U9139 (N_9139,N_6770,N_7611);
and U9140 (N_9140,N_6571,N_4780);
nand U9141 (N_9141,N_7400,N_4088);
nand U9142 (N_9142,N_6865,N_5914);
nand U9143 (N_9143,N_6374,N_7461);
or U9144 (N_9144,N_6056,N_5020);
nand U9145 (N_9145,N_7049,N_4564);
nor U9146 (N_9146,N_6066,N_4392);
nor U9147 (N_9147,N_7110,N_4542);
or U9148 (N_9148,N_5756,N_7440);
or U9149 (N_9149,N_5970,N_7933);
xor U9150 (N_9150,N_5063,N_7013);
nand U9151 (N_9151,N_4108,N_7873);
xor U9152 (N_9152,N_5814,N_4663);
nor U9153 (N_9153,N_7899,N_6783);
nor U9154 (N_9154,N_6281,N_7862);
and U9155 (N_9155,N_6961,N_4730);
and U9156 (N_9156,N_6784,N_4114);
or U9157 (N_9157,N_6696,N_5391);
nand U9158 (N_9158,N_7127,N_6120);
nor U9159 (N_9159,N_5443,N_5146);
nand U9160 (N_9160,N_6090,N_7939);
or U9161 (N_9161,N_6839,N_5689);
nand U9162 (N_9162,N_7520,N_6316);
and U9163 (N_9163,N_6682,N_6348);
or U9164 (N_9164,N_6807,N_7074);
or U9165 (N_9165,N_7171,N_4394);
and U9166 (N_9166,N_7990,N_5224);
or U9167 (N_9167,N_4353,N_7758);
and U9168 (N_9168,N_6463,N_5113);
nor U9169 (N_9169,N_7902,N_7751);
xor U9170 (N_9170,N_4592,N_4208);
xnor U9171 (N_9171,N_7925,N_5170);
or U9172 (N_9172,N_5335,N_7473);
nand U9173 (N_9173,N_6653,N_5487);
and U9174 (N_9174,N_7307,N_4137);
nor U9175 (N_9175,N_5503,N_5854);
nor U9176 (N_9176,N_6974,N_5201);
nand U9177 (N_9177,N_7297,N_6427);
nand U9178 (N_9178,N_5993,N_7623);
nor U9179 (N_9179,N_6685,N_4017);
nand U9180 (N_9180,N_4543,N_4796);
and U9181 (N_9181,N_6613,N_4976);
xor U9182 (N_9182,N_5216,N_5787);
and U9183 (N_9183,N_6354,N_4865);
and U9184 (N_9184,N_4433,N_5012);
or U9185 (N_9185,N_6574,N_7865);
or U9186 (N_9186,N_6796,N_7699);
or U9187 (N_9187,N_6028,N_4912);
xor U9188 (N_9188,N_5779,N_6309);
nand U9189 (N_9189,N_7636,N_4868);
nor U9190 (N_9190,N_5586,N_6936);
nand U9191 (N_9191,N_6676,N_6474);
nor U9192 (N_9192,N_7803,N_5983);
or U9193 (N_9193,N_7419,N_7439);
nor U9194 (N_9194,N_5783,N_4230);
xnor U9195 (N_9195,N_4923,N_5755);
xnor U9196 (N_9196,N_5427,N_4443);
or U9197 (N_9197,N_6005,N_6461);
nand U9198 (N_9198,N_4223,N_6152);
nand U9199 (N_9199,N_6051,N_7967);
xor U9200 (N_9200,N_4243,N_4806);
or U9201 (N_9201,N_5410,N_4798);
and U9202 (N_9202,N_6244,N_7220);
xor U9203 (N_9203,N_4605,N_6088);
or U9204 (N_9204,N_4988,N_7194);
xnor U9205 (N_9205,N_6138,N_5296);
and U9206 (N_9206,N_6454,N_6949);
or U9207 (N_9207,N_6122,N_4616);
and U9208 (N_9208,N_5154,N_5000);
and U9209 (N_9209,N_6198,N_6986);
xor U9210 (N_9210,N_6977,N_5584);
nand U9211 (N_9211,N_6351,N_7209);
xor U9212 (N_9212,N_7757,N_7662);
or U9213 (N_9213,N_6276,N_4200);
or U9214 (N_9214,N_6812,N_5105);
nor U9215 (N_9215,N_6858,N_7397);
nor U9216 (N_9216,N_7683,N_6808);
nand U9217 (N_9217,N_7958,N_4015);
xnor U9218 (N_9218,N_7541,N_4751);
nand U9219 (N_9219,N_4293,N_4602);
and U9220 (N_9220,N_5805,N_4411);
nand U9221 (N_9221,N_5594,N_6184);
xnor U9222 (N_9222,N_6786,N_6842);
or U9223 (N_9223,N_4709,N_4492);
nor U9224 (N_9224,N_5654,N_7084);
nand U9225 (N_9225,N_6922,N_6557);
nand U9226 (N_9226,N_7605,N_6165);
nand U9227 (N_9227,N_4006,N_4331);
nand U9228 (N_9228,N_7800,N_7235);
nand U9229 (N_9229,N_7174,N_6758);
xor U9230 (N_9230,N_4547,N_4685);
nand U9231 (N_9231,N_5017,N_6957);
and U9232 (N_9232,N_7279,N_5581);
xor U9233 (N_9233,N_7444,N_5633);
xnor U9234 (N_9234,N_6401,N_5260);
nand U9235 (N_9235,N_4789,N_5938);
and U9236 (N_9236,N_5087,N_7451);
and U9237 (N_9237,N_4002,N_7292);
or U9238 (N_9238,N_4212,N_6730);
nand U9239 (N_9239,N_6141,N_7316);
xor U9240 (N_9240,N_7161,N_4097);
and U9241 (N_9241,N_6566,N_6511);
or U9242 (N_9242,N_5897,N_5508);
or U9243 (N_9243,N_7771,N_4306);
or U9244 (N_9244,N_4081,N_7366);
or U9245 (N_9245,N_4517,N_7204);
nand U9246 (N_9246,N_7170,N_6959);
and U9247 (N_9247,N_7237,N_7401);
or U9248 (N_9248,N_7140,N_5627);
or U9249 (N_9249,N_5444,N_6311);
xnor U9250 (N_9250,N_4836,N_7624);
nor U9251 (N_9251,N_4235,N_6611);
nor U9252 (N_9252,N_7024,N_7211);
nor U9253 (N_9253,N_6376,N_4858);
nor U9254 (N_9254,N_7684,N_5542);
nand U9255 (N_9255,N_7333,N_5329);
nor U9256 (N_9256,N_7141,N_6343);
or U9257 (N_9257,N_4427,N_4634);
xor U9258 (N_9258,N_7582,N_5145);
xor U9259 (N_9259,N_7313,N_7343);
nor U9260 (N_9260,N_5891,N_4532);
or U9261 (N_9261,N_7135,N_4246);
nand U9262 (N_9262,N_4952,N_6706);
and U9263 (N_9263,N_5060,N_5466);
nor U9264 (N_9264,N_4119,N_5546);
nor U9265 (N_9265,N_4658,N_6788);
and U9266 (N_9266,N_6317,N_7256);
and U9267 (N_9267,N_4642,N_6755);
or U9268 (N_9268,N_7768,N_7213);
or U9269 (N_9269,N_5815,N_4382);
xnor U9270 (N_9270,N_7670,N_4608);
xnor U9271 (N_9271,N_5840,N_7536);
and U9272 (N_9272,N_6408,N_5557);
or U9273 (N_9273,N_5962,N_5875);
nor U9274 (N_9274,N_6065,N_6352);
or U9275 (N_9275,N_4226,N_5162);
or U9276 (N_9276,N_7995,N_5344);
xor U9277 (N_9277,N_4347,N_5625);
xnor U9278 (N_9278,N_7322,N_4704);
xnor U9279 (N_9279,N_7290,N_6635);
nor U9280 (N_9280,N_6292,N_5450);
nand U9281 (N_9281,N_5250,N_7615);
or U9282 (N_9282,N_7829,N_4690);
or U9283 (N_9283,N_6913,N_7285);
nor U9284 (N_9284,N_4407,N_4917);
and U9285 (N_9285,N_6233,N_5337);
nor U9286 (N_9286,N_7578,N_6701);
or U9287 (N_9287,N_4535,N_7749);
and U9288 (N_9288,N_5651,N_5507);
nor U9289 (N_9289,N_7855,N_6326);
xnor U9290 (N_9290,N_4807,N_6096);
or U9291 (N_9291,N_4560,N_5615);
xnor U9292 (N_9292,N_7340,N_4732);
nand U9293 (N_9293,N_7631,N_6271);
and U9294 (N_9294,N_5121,N_6543);
nor U9295 (N_9295,N_7901,N_5282);
xnor U9296 (N_9296,N_5817,N_7324);
nor U9297 (N_9297,N_4919,N_6550);
and U9298 (N_9298,N_6400,N_4409);
and U9299 (N_9299,N_5031,N_5553);
nor U9300 (N_9300,N_5622,N_7888);
xor U9301 (N_9301,N_5353,N_6608);
and U9302 (N_9302,N_4298,N_6336);
and U9303 (N_9303,N_4986,N_4698);
nor U9304 (N_9304,N_6240,N_6419);
or U9305 (N_9305,N_4086,N_7457);
xor U9306 (N_9306,N_7392,N_4855);
nor U9307 (N_9307,N_6994,N_5039);
nor U9308 (N_9308,N_4628,N_4659);
nor U9309 (N_9309,N_7139,N_6022);
nand U9310 (N_9310,N_4635,N_6723);
nor U9311 (N_9311,N_7072,N_5796);
nor U9312 (N_9312,N_7860,N_7177);
or U9313 (N_9313,N_5597,N_5036);
nor U9314 (N_9314,N_4136,N_6815);
xnor U9315 (N_9315,N_4870,N_4938);
nand U9316 (N_9316,N_4117,N_4009);
nand U9317 (N_9317,N_6618,N_7370);
nor U9318 (N_9318,N_4451,N_6166);
and U9319 (N_9319,N_7678,N_6862);
xor U9320 (N_9320,N_4463,N_7522);
nor U9321 (N_9321,N_7529,N_7600);
or U9322 (N_9322,N_5155,N_6622);
and U9323 (N_9323,N_7267,N_7123);
nor U9324 (N_9324,N_5936,N_4721);
and U9325 (N_9325,N_7460,N_5562);
xnor U9326 (N_9326,N_5027,N_7178);
nand U9327 (N_9327,N_4276,N_4362);
nor U9328 (N_9328,N_5191,N_5286);
nor U9329 (N_9329,N_5262,N_7887);
and U9330 (N_9330,N_4664,N_6591);
and U9331 (N_9331,N_6855,N_4266);
or U9332 (N_9332,N_6709,N_5925);
xor U9333 (N_9333,N_7739,N_4254);
or U9334 (N_9334,N_7238,N_6301);
nand U9335 (N_9335,N_6797,N_6982);
xnor U9336 (N_9336,N_7828,N_7717);
nand U9337 (N_9337,N_4859,N_6344);
and U9338 (N_9338,N_6062,N_7331);
nand U9339 (N_9339,N_4706,N_5941);
or U9340 (N_9340,N_7964,N_4534);
nand U9341 (N_9341,N_4290,N_6520);
and U9342 (N_9342,N_5089,N_4910);
nor U9343 (N_9343,N_6091,N_5935);
nor U9344 (N_9344,N_4320,N_6449);
and U9345 (N_9345,N_5092,N_5098);
nand U9346 (N_9346,N_6978,N_7950);
xnor U9347 (N_9347,N_7812,N_4747);
and U9348 (N_9348,N_7405,N_4369);
and U9349 (N_9349,N_4522,N_7815);
xor U9350 (N_9350,N_5650,N_6288);
and U9351 (N_9351,N_4496,N_6469);
nor U9352 (N_9352,N_4959,N_5275);
xnor U9353 (N_9353,N_7434,N_5673);
xnor U9354 (N_9354,N_6250,N_4929);
and U9355 (N_9355,N_6666,N_6086);
nand U9356 (N_9356,N_4449,N_5447);
nand U9357 (N_9357,N_6681,N_5692);
nand U9358 (N_9358,N_7294,N_5607);
and U9359 (N_9359,N_6556,N_5381);
and U9360 (N_9360,N_5261,N_7002);
nand U9361 (N_9361,N_7826,N_5448);
xnor U9362 (N_9362,N_5598,N_5220);
nor U9363 (N_9363,N_6782,N_6625);
and U9364 (N_9364,N_6208,N_5883);
or U9365 (N_9365,N_5357,N_4237);
xnor U9366 (N_9366,N_7162,N_6190);
nand U9367 (N_9367,N_7709,N_6654);
xnor U9368 (N_9368,N_5083,N_7937);
nand U9369 (N_9369,N_7325,N_4947);
nand U9370 (N_9370,N_5998,N_4037);
or U9371 (N_9371,N_6265,N_7628);
nor U9372 (N_9372,N_6295,N_7714);
xnor U9373 (N_9373,N_5209,N_4211);
or U9374 (N_9374,N_5119,N_5195);
nor U9375 (N_9375,N_4085,N_5697);
nor U9376 (N_9376,N_7927,N_5291);
or U9377 (N_9377,N_4181,N_7905);
nor U9378 (N_9378,N_6871,N_6630);
xnor U9379 (N_9379,N_6196,N_7908);
nand U9380 (N_9380,N_6919,N_6269);
xnor U9381 (N_9381,N_6437,N_6569);
nand U9382 (N_9382,N_5360,N_4177);
nor U9383 (N_9383,N_5311,N_4012);
or U9384 (N_9384,N_6186,N_5321);
or U9385 (N_9385,N_7067,N_6643);
or U9386 (N_9386,N_5736,N_7181);
xor U9387 (N_9387,N_4563,N_4170);
xnor U9388 (N_9388,N_4141,N_5233);
and U9389 (N_9389,N_4552,N_5032);
nor U9390 (N_9390,N_6891,N_6996);
xnor U9391 (N_9391,N_7346,N_4576);
xor U9392 (N_9392,N_5171,N_5161);
xor U9393 (N_9393,N_7488,N_4618);
xnor U9394 (N_9394,N_7431,N_6693);
or U9395 (N_9395,N_5985,N_4970);
and U9396 (N_9396,N_6299,N_6945);
or U9397 (N_9397,N_4570,N_6927);
nor U9398 (N_9398,N_5313,N_6123);
and U9399 (N_9399,N_5200,N_7827);
nor U9400 (N_9400,N_4333,N_4992);
nand U9401 (N_9401,N_6134,N_6393);
and U9402 (N_9402,N_5342,N_6760);
and U9403 (N_9403,N_6156,N_5231);
nor U9404 (N_9404,N_5859,N_4283);
or U9405 (N_9405,N_4302,N_5676);
and U9406 (N_9406,N_7932,N_7062);
nor U9407 (N_9407,N_5299,N_4875);
xnor U9408 (N_9408,N_4318,N_5967);
nor U9409 (N_9409,N_6827,N_7511);
and U9410 (N_9410,N_7753,N_6505);
xnor U9411 (N_9411,N_4264,N_5675);
nor U9412 (N_9412,N_6692,N_5148);
or U9413 (N_9413,N_5421,N_5860);
nor U9414 (N_9414,N_6448,N_4470);
nand U9415 (N_9415,N_4389,N_7881);
nor U9416 (N_9416,N_4940,N_5616);
or U9417 (N_9417,N_4609,N_4180);
and U9418 (N_9418,N_4502,N_6042);
xnor U9419 (N_9419,N_6984,N_4385);
and U9420 (N_9420,N_7923,N_4699);
nor U9421 (N_9421,N_5726,N_7261);
xor U9422 (N_9422,N_5249,N_5283);
nor U9423 (N_9423,N_7168,N_4168);
or U9424 (N_9424,N_7240,N_6756);
nand U9425 (N_9425,N_4785,N_4410);
nor U9426 (N_9426,N_7894,N_7138);
nand U9427 (N_9427,N_7498,N_4057);
or U9428 (N_9428,N_5974,N_7926);
nor U9429 (N_9429,N_6739,N_7752);
nand U9430 (N_9430,N_5751,N_4171);
nor U9431 (N_9431,N_7150,N_4341);
xnor U9432 (N_9432,N_6270,N_7034);
xnor U9433 (N_9433,N_4578,N_4687);
nor U9434 (N_9434,N_6384,N_7938);
nand U9435 (N_9435,N_6424,N_4927);
xor U9436 (N_9436,N_5547,N_5485);
nand U9437 (N_9437,N_6137,N_7532);
nor U9438 (N_9438,N_4143,N_6506);
nor U9439 (N_9439,N_7464,N_7172);
nand U9440 (N_9440,N_7720,N_6221);
xnor U9441 (N_9441,N_6324,N_6708);
nand U9442 (N_9442,N_4084,N_6499);
xnor U9443 (N_9443,N_5536,N_7688);
xor U9444 (N_9444,N_7935,N_7916);
nor U9445 (N_9445,N_5990,N_4755);
xor U9446 (N_9446,N_7861,N_7208);
and U9447 (N_9447,N_7557,N_4760);
nand U9448 (N_9448,N_4419,N_6207);
and U9449 (N_9449,N_6298,N_7023);
and U9450 (N_9450,N_7306,N_7986);
nand U9451 (N_9451,N_5934,N_7483);
nor U9452 (N_9452,N_7262,N_7763);
nand U9453 (N_9453,N_5867,N_5655);
nand U9454 (N_9454,N_5412,N_5107);
nand U9455 (N_9455,N_6920,N_5168);
nor U9456 (N_9456,N_7570,N_7158);
and U9457 (N_9457,N_6036,N_4581);
xnor U9458 (N_9458,N_6564,N_4505);
nor U9459 (N_9459,N_6761,N_5694);
nand U9460 (N_9460,N_6183,N_6304);
nand U9461 (N_9461,N_4841,N_7633);
nand U9462 (N_9462,N_7971,N_5140);
or U9463 (N_9463,N_7143,N_6473);
nand U9464 (N_9464,N_6627,N_5110);
and U9465 (N_9465,N_6381,N_4587);
xor U9466 (N_9466,N_7303,N_5183);
and U9467 (N_9467,N_4775,N_7639);
nand U9468 (N_9468,N_5256,N_4342);
or U9469 (N_9469,N_4018,N_6909);
xor U9470 (N_9470,N_5302,N_4456);
nor U9471 (N_9471,N_6667,N_5079);
nand U9472 (N_9472,N_7819,N_5517);
nor U9473 (N_9473,N_6378,N_6131);
nor U9474 (N_9474,N_5913,N_6323);
or U9475 (N_9475,N_4997,N_4600);
or U9476 (N_9476,N_6623,N_4931);
nor U9477 (N_9477,N_6652,N_5456);
nor U9478 (N_9478,N_4336,N_7005);
or U9479 (N_9479,N_6697,N_4745);
nor U9480 (N_9480,N_7478,N_4816);
nand U9481 (N_9481,N_4597,N_4459);
xnor U9482 (N_9482,N_6586,N_5734);
nand U9483 (N_9483,N_7549,N_5511);
nor U9484 (N_9484,N_5382,N_7293);
and U9485 (N_9485,N_7423,N_4262);
nand U9486 (N_9486,N_7808,N_5872);
nand U9487 (N_9487,N_4378,N_5984);
or U9488 (N_9488,N_4759,N_7893);
or U9489 (N_9489,N_4782,N_6606);
or U9490 (N_9490,N_5876,N_4019);
xnor U9491 (N_9491,N_5765,N_6181);
nor U9492 (N_9492,N_5061,N_7809);
nor U9493 (N_9493,N_5895,N_6596);
or U9494 (N_9494,N_5462,N_4144);
xor U9495 (N_9495,N_4548,N_5928);
xnor U9496 (N_9496,N_4278,N_7044);
or U9497 (N_9497,N_7913,N_5679);
nand U9498 (N_9498,N_4123,N_6377);
or U9499 (N_9499,N_6191,N_5175);
or U9500 (N_9500,N_4167,N_7165);
xor U9501 (N_9501,N_4933,N_5108);
nand U9502 (N_9502,N_5980,N_5771);
xnor U9503 (N_9503,N_6640,N_5492);
nor U9504 (N_9504,N_4675,N_6663);
xor U9505 (N_9505,N_7215,N_5515);
nor U9506 (N_9506,N_5844,N_4648);
or U9507 (N_9507,N_7330,N_5237);
nor U9508 (N_9508,N_7762,N_6175);
and U9509 (N_9509,N_7569,N_7087);
or U9510 (N_9510,N_5409,N_7031);
nor U9511 (N_9511,N_6633,N_4932);
xor U9512 (N_9512,N_6034,N_6179);
or U9513 (N_9513,N_4272,N_5472);
xor U9514 (N_9514,N_5838,N_5884);
xor U9515 (N_9515,N_5987,N_5826);
xnor U9516 (N_9516,N_7851,N_5623);
nand U9517 (N_9517,N_4270,N_7936);
or U9518 (N_9518,N_4134,N_5229);
nor U9519 (N_9519,N_7301,N_7577);
nor U9520 (N_9520,N_5136,N_4649);
nor U9521 (N_9521,N_5569,N_6213);
or U9522 (N_9522,N_6385,N_6194);
and U9523 (N_9523,N_7747,N_7689);
xor U9524 (N_9524,N_7609,N_6335);
nor U9525 (N_9525,N_4000,N_7804);
xnor U9526 (N_9526,N_4787,N_6830);
or U9527 (N_9527,N_4013,N_5461);
nand U9528 (N_9528,N_6132,N_5106);
xnor U9529 (N_9529,N_5469,N_7245);
nand U9530 (N_9530,N_6991,N_7428);
or U9531 (N_9531,N_6738,N_7907);
nor U9532 (N_9532,N_5621,N_7619);
nand U9533 (N_9533,N_5610,N_7738);
and U9534 (N_9534,N_7357,N_4027);
xor U9535 (N_9535,N_6441,N_4876);
or U9536 (N_9536,N_4660,N_7798);
or U9537 (N_9537,N_6081,N_5418);
and U9538 (N_9538,N_4175,N_4120);
nor U9539 (N_9539,N_5525,N_6023);
and U9540 (N_9540,N_6838,N_4693);
and U9541 (N_9541,N_4639,N_4813);
nor U9542 (N_9542,N_5072,N_6365);
nor U9543 (N_9543,N_4343,N_7114);
nor U9544 (N_9544,N_6216,N_6863);
and U9545 (N_9545,N_6734,N_6990);
or U9546 (N_9546,N_4799,N_5644);
nand U9547 (N_9547,N_7889,N_5786);
or U9548 (N_9548,N_6655,N_7283);
and U9549 (N_9549,N_6169,N_6128);
nand U9550 (N_9550,N_4124,N_7642);
or U9551 (N_9551,N_4067,N_6078);
nand U9552 (N_9552,N_7740,N_6459);
and U9553 (N_9553,N_7526,N_7415);
or U9554 (N_9554,N_7255,N_7275);
or U9555 (N_9555,N_5948,N_5182);
xnor U9556 (N_9556,N_5475,N_6703);
nand U9557 (N_9557,N_5369,N_4515);
nand U9558 (N_9558,N_6794,N_4538);
and U9559 (N_9559,N_5886,N_7746);
xor U9560 (N_9560,N_6177,N_6856);
and U9561 (N_9561,N_5812,N_5459);
xnor U9562 (N_9562,N_4477,N_4554);
xnor U9563 (N_9563,N_7707,N_5521);
and U9564 (N_9564,N_6941,N_6019);
and U9565 (N_9565,N_4448,N_4372);
xnor U9566 (N_9566,N_4220,N_7120);
xnor U9567 (N_9567,N_5834,N_7801);
xor U9568 (N_9568,N_4667,N_6773);
nand U9569 (N_9569,N_6669,N_7304);
nand U9570 (N_9570,N_5244,N_6877);
and U9571 (N_9571,N_7730,N_4197);
and U9572 (N_9572,N_4275,N_6247);
nor U9573 (N_9573,N_4847,N_5270);
nand U9574 (N_9574,N_5951,N_6545);
nor U9575 (N_9575,N_6664,N_4956);
nand U9576 (N_9576,N_6263,N_7335);
and U9577 (N_9577,N_6525,N_7384);
xor U9578 (N_9578,N_6828,N_7448);
nand U9579 (N_9579,N_7210,N_5180);
nand U9580 (N_9580,N_5758,N_4312);
and U9581 (N_9581,N_6136,N_7612);
or U9582 (N_9582,N_4401,N_5366);
nor U9583 (N_9583,N_7227,N_4361);
xor U9584 (N_9584,N_4031,N_5018);
or U9585 (N_9585,N_7491,N_4974);
nor U9586 (N_9586,N_4983,N_5026);
nand U9587 (N_9587,N_6503,N_5217);
or U9588 (N_9588,N_7269,N_6371);
and U9589 (N_9589,N_7360,N_5919);
or U9590 (N_9590,N_7417,N_4575);
and U9591 (N_9591,N_4930,N_5392);
nand U9592 (N_9592,N_6515,N_7742);
nor U9593 (N_9593,N_4700,N_6629);
nor U9594 (N_9594,N_4152,N_7232);
xnor U9595 (N_9595,N_7954,N_6349);
and U9596 (N_9596,N_4545,N_6223);
or U9597 (N_9597,N_4174,N_5700);
and U9598 (N_9598,N_4191,N_7981);
nor U9599 (N_9599,N_5929,N_5889);
or U9600 (N_9600,N_7308,N_4562);
or U9601 (N_9601,N_5804,N_4222);
xor U9602 (N_9602,N_7816,N_6382);
or U9603 (N_9603,N_5305,N_4920);
and U9604 (N_9604,N_7743,N_5743);
and U9605 (N_9605,N_6130,N_6118);
nor U9606 (N_9606,N_7310,N_4673);
or U9607 (N_9607,N_6795,N_5248);
xnor U9608 (N_9608,N_5638,N_5773);
and U9609 (N_9609,N_4292,N_6135);
and U9610 (N_9610,N_6901,N_5050);
and U9611 (N_9611,N_5708,N_5205);
and U9612 (N_9612,N_6695,N_6809);
nand U9613 (N_9613,N_6969,N_6403);
and U9614 (N_9614,N_5986,N_5710);
nand U9615 (N_9615,N_5465,N_4883);
nor U9616 (N_9616,N_7012,N_4960);
nand U9617 (N_9617,N_7053,N_5923);
or U9618 (N_9618,N_7085,N_6158);
nand U9619 (N_9619,N_6021,N_7671);
nand U9620 (N_9620,N_5863,N_4792);
or U9621 (N_9621,N_6775,N_5437);
nand U9622 (N_9622,N_4815,N_4654);
nand U9623 (N_9623,N_5519,N_5568);
nor U9624 (N_9624,N_4305,N_5045);
nand U9625 (N_9625,N_5764,N_7035);
nand U9626 (N_9626,N_5856,N_7983);
xnor U9627 (N_9627,N_6981,N_7479);
and U9628 (N_9628,N_6110,N_5885);
nand U9629 (N_9629,N_4400,N_5691);
xor U9630 (N_9630,N_6321,N_6715);
and U9631 (N_9631,N_7915,N_7125);
nor U9632 (N_9632,N_5207,N_7253);
xor U9633 (N_9633,N_7193,N_4606);
xor U9634 (N_9634,N_4360,N_7599);
xor U9635 (N_9635,N_4694,N_5611);
and U9636 (N_9636,N_4750,N_7792);
nor U9637 (N_9637,N_6874,N_5588);
or U9638 (N_9638,N_7895,N_7661);
or U9639 (N_9639,N_5900,N_7218);
or U9640 (N_9640,N_4072,N_7799);
nor U9641 (N_9641,N_7581,N_5982);
nor U9642 (N_9642,N_5677,N_5685);
nand U9643 (N_9643,N_4484,N_5439);
and U9644 (N_9644,N_6007,N_7344);
or U9645 (N_9645,N_4758,N_6599);
or U9646 (N_9646,N_6846,N_7648);
and U9647 (N_9647,N_4116,N_4511);
nand U9648 (N_9648,N_5234,N_6535);
nor U9649 (N_9649,N_7001,N_6080);
and U9650 (N_9650,N_6402,N_7342);
xor U9651 (N_9651,N_5197,N_4106);
nor U9652 (N_9652,N_7040,N_4877);
and U9653 (N_9653,N_5240,N_7495);
nor U9654 (N_9654,N_5395,N_7490);
xnor U9655 (N_9655,N_4467,N_5862);
and U9656 (N_9656,N_6242,N_5399);
and U9657 (N_9657,N_4214,N_6854);
xor U9658 (N_9658,N_7226,N_6327);
nand U9659 (N_9659,N_4679,N_6650);
or U9660 (N_9660,N_4561,N_5218);
and U9661 (N_9661,N_4978,N_7115);
xnor U9662 (N_9662,N_6836,N_6129);
or U9663 (N_9663,N_4303,N_7184);
nor U9664 (N_9664,N_6632,N_4050);
and U9665 (N_9665,N_7109,N_6875);
and U9666 (N_9666,N_4766,N_5174);
nor U9667 (N_9667,N_4397,N_7466);
nor U9668 (N_9668,N_6471,N_7169);
and U9669 (N_9669,N_6698,N_7848);
nand U9670 (N_9670,N_6082,N_5029);
and U9671 (N_9671,N_6442,N_6829);
and U9672 (N_9672,N_5411,N_4365);
and U9673 (N_9673,N_7107,N_7284);
xnor U9674 (N_9674,N_5902,N_5558);
and U9675 (N_9675,N_4671,N_7657);
and U9676 (N_9676,N_7167,N_4296);
nand U9677 (N_9677,N_6030,N_4557);
nor U9678 (N_9678,N_4499,N_6524);
xnor U9679 (N_9679,N_7725,N_7517);
nor U9680 (N_9680,N_6947,N_4231);
or U9681 (N_9681,N_6436,N_5645);
nor U9682 (N_9682,N_4412,N_4848);
nand U9683 (N_9683,N_7015,N_6528);
nand U9684 (N_9684,N_5823,N_7296);
nor U9685 (N_9685,N_5365,N_4800);
nor U9686 (N_9686,N_7337,N_7567);
xnor U9687 (N_9687,N_5151,N_5254);
and U9688 (N_9688,N_4090,N_7159);
or U9689 (N_9689,N_5716,N_4098);
or U9690 (N_9690,N_6248,N_6008);
or U9691 (N_9691,N_6164,N_6297);
and U9692 (N_9692,N_7097,N_7896);
or U9693 (N_9693,N_4778,N_5696);
nand U9694 (N_9694,N_4323,N_5608);
nand U9695 (N_9695,N_4479,N_5567);
nor U9696 (N_9696,N_4716,N_4388);
and U9697 (N_9697,N_7790,N_4531);
and U9698 (N_9698,N_7691,N_6068);
or U9699 (N_9699,N_6476,N_4668);
nor U9700 (N_9700,N_6924,N_6744);
nand U9701 (N_9701,N_6399,N_5730);
nor U9702 (N_9702,N_4473,N_6801);
or U9703 (N_9703,N_6649,N_5724);
and U9704 (N_9704,N_7919,N_6341);
xnor U9705 (N_9705,N_5100,N_7270);
nor U9706 (N_9706,N_4450,N_7004);
nand U9707 (N_9707,N_7604,N_6502);
or U9708 (N_9708,N_5662,N_7219);
nand U9709 (N_9709,N_7300,N_4094);
xnor U9710 (N_9710,N_5075,N_6101);
and U9711 (N_9711,N_6490,N_7247);
or U9712 (N_9712,N_5097,N_7271);
xor U9713 (N_9713,N_4173,N_4157);
or U9714 (N_9714,N_5740,N_4213);
and U9715 (N_9715,N_6851,N_6776);
xnor U9716 (N_9716,N_4370,N_6050);
nand U9717 (N_9717,N_4454,N_7516);
nor U9718 (N_9718,N_7399,N_4797);
xnor U9719 (N_9719,N_4398,N_6822);
nor U9720 (N_9720,N_6993,N_7830);
nand U9721 (N_9721,N_7543,N_4588);
or U9722 (N_9722,N_5423,N_5591);
nand U9723 (N_9723,N_6443,N_5604);
nor U9724 (N_9724,N_5715,N_4665);
nor U9725 (N_9725,N_4725,N_6645);
and U9726 (N_9726,N_7521,N_6724);
and U9727 (N_9727,N_7081,N_4832);
nor U9728 (N_9728,N_6061,N_6199);
nor U9729 (N_9729,N_5005,N_5374);
nand U9730 (N_9730,N_7056,N_4520);
nand U9731 (N_9731,N_7793,N_7176);
or U9732 (N_9732,N_6694,N_5506);
nand U9733 (N_9733,N_4504,N_7390);
and U9734 (N_9734,N_6149,N_6153);
nand U9735 (N_9735,N_6790,N_6598);
xnor U9736 (N_9736,N_4615,N_6787);
and U9737 (N_9737,N_6728,N_6396);
nand U9738 (N_9738,N_5188,N_4835);
and U9739 (N_9739,N_6748,N_7878);
or U9740 (N_9740,N_4112,N_4062);
xnor U9741 (N_9741,N_4187,N_6929);
and U9742 (N_9742,N_6911,N_4021);
nor U9743 (N_9743,N_5372,N_4743);
nand U9744 (N_9744,N_4888,N_4161);
nor U9745 (N_9745,N_6252,N_5978);
nand U9746 (N_9746,N_4316,N_6058);
xnor U9747 (N_9747,N_5315,N_4376);
or U9748 (N_9748,N_6210,N_6956);
nor U9749 (N_9749,N_4415,N_6383);
and U9750 (N_9750,N_4712,N_4413);
nor U9751 (N_9751,N_7857,N_4183);
nand U9752 (N_9752,N_6580,N_4791);
xnor U9753 (N_9753,N_6193,N_7320);
and U9754 (N_9754,N_7558,N_7675);
nor U9755 (N_9755,N_7864,N_6279);
xnor U9756 (N_9756,N_7962,N_6837);
or U9757 (N_9757,N_6433,N_6712);
or U9758 (N_9758,N_5203,N_4555);
nand U9759 (N_9759,N_7071,N_4942);
and U9760 (N_9760,N_6634,N_5124);
and U9761 (N_9761,N_6303,N_6147);
and U9762 (N_9762,N_4962,N_6102);
or U9763 (N_9763,N_5988,N_4440);
nor U9764 (N_9764,N_5006,N_4593);
xnor U9765 (N_9765,N_7672,N_6678);
xor U9766 (N_9766,N_6646,N_5323);
xnor U9767 (N_9767,N_4998,N_5882);
or U9768 (N_9768,N_6925,N_7069);
nand U9769 (N_9769,N_5460,N_4344);
nor U9770 (N_9770,N_4647,N_6325);
and U9771 (N_9771,N_7872,N_7243);
and U9772 (N_9772,N_4204,N_5643);
or U9773 (N_9773,N_6518,N_7481);
xor U9774 (N_9774,N_7655,N_5852);
and U9775 (N_9775,N_5749,N_4265);
xnor U9776 (N_9776,N_4678,N_5966);
and U9777 (N_9777,N_6883,N_6284);
or U9778 (N_9778,N_5298,N_6428);
or U9779 (N_9779,N_5866,N_6725);
nor U9780 (N_9780,N_4381,N_4795);
nor U9781 (N_9781,N_6610,N_5782);
xor U9782 (N_9782,N_6497,N_4669);
xor U9783 (N_9783,N_4611,N_5904);
xor U9784 (N_9784,N_4925,N_7856);
nor U9785 (N_9785,N_7470,N_5164);
and U9786 (N_9786,N_7180,N_4076);
or U9787 (N_9787,N_7233,N_4915);
nand U9788 (N_9788,N_4271,N_6609);
nor U9789 (N_9789,N_5208,N_6413);
and U9790 (N_9790,N_4066,N_7910);
or U9791 (N_9791,N_5915,N_7207);
or U9792 (N_9792,N_5178,N_6568);
nor U9793 (N_9793,N_4644,N_7966);
nor U9794 (N_9794,N_6970,N_4708);
xnor U9795 (N_9795,N_6125,N_6390);
xor U9796 (N_9796,N_4966,N_4471);
and U9797 (N_9797,N_4523,N_6151);
or U9798 (N_9798,N_5509,N_4172);
xnor U9799 (N_9799,N_6358,N_5037);
xor U9800 (N_9800,N_7079,N_6572);
or U9801 (N_9801,N_7796,N_4506);
and U9802 (N_9802,N_7820,N_5937);
xnor U9803 (N_9803,N_6621,N_7286);
nand U9804 (N_9804,N_4421,N_7960);
nand U9805 (N_9805,N_5300,N_6835);
xor U9806 (N_9806,N_4566,N_5227);
xor U9807 (N_9807,N_6117,N_6892);
nor U9808 (N_9808,N_4924,N_4612);
or U9809 (N_9809,N_4958,N_7780);
xor U9810 (N_9810,N_6308,N_5252);
or U9811 (N_9811,N_6084,N_7022);
and U9812 (N_9812,N_7610,N_5219);
nand U9813 (N_9813,N_6777,N_4869);
and U9814 (N_9814,N_7595,N_6037);
nor U9815 (N_9815,N_7083,N_6055);
nor U9816 (N_9816,N_7118,N_4043);
nand U9817 (N_9817,N_6677,N_6089);
and U9818 (N_9818,N_5334,N_6113);
and U9819 (N_9819,N_5259,N_5137);
nand U9820 (N_9820,N_4217,N_6774);
nand U9821 (N_9821,N_7006,N_5837);
and U9822 (N_9822,N_7091,N_6423);
or U9823 (N_9823,N_7021,N_5477);
nand U9824 (N_9824,N_4895,N_5206);
or U9825 (N_9825,N_4957,N_5803);
nor U9826 (N_9826,N_5184,N_7880);
xnor U9827 (N_9827,N_7692,N_6373);
or U9828 (N_9828,N_6570,N_6294);
xor U9829 (N_9829,N_4980,N_6885);
nand U9830 (N_9830,N_4104,N_6971);
xnor U9831 (N_9831,N_5125,N_4825);
or U9832 (N_9832,N_7774,N_4972);
xnor U9833 (N_9833,N_5668,N_4722);
nand U9834 (N_9834,N_6914,N_7130);
or U9835 (N_9835,N_5035,N_6355);
nor U9836 (N_9836,N_4946,N_5669);
and U9837 (N_9837,N_5049,N_7715);
xor U9838 (N_9838,N_4676,N_6817);
nand U9839 (N_9839,N_7014,N_7189);
nand U9840 (N_9840,N_5002,N_4905);
xor U9841 (N_9841,N_7785,N_4251);
nand U9842 (N_9842,N_6989,N_4190);
nand U9843 (N_9843,N_4188,N_6721);
and U9844 (N_9844,N_7711,N_6320);
xnor U9845 (N_9845,N_6890,N_7525);
nand U9846 (N_9846,N_6904,N_4514);
or U9847 (N_9847,N_7096,N_6259);
and U9848 (N_9848,N_6176,N_5971);
nor U9849 (N_9849,N_4845,N_4990);
xor U9850 (N_9850,N_5273,N_7911);
nand U9851 (N_9851,N_4691,N_7668);
nor U9852 (N_9852,N_7898,N_7649);
xnor U9853 (N_9853,N_6926,N_5054);
and U9854 (N_9854,N_5101,N_4279);
and U9855 (N_9855,N_4779,N_5873);
or U9856 (N_9856,N_7883,N_4147);
xnor U9857 (N_9857,N_5314,N_6251);
nor U9858 (N_9858,N_5612,N_7477);
nor U9859 (N_9859,N_7145,N_5845);
or U9860 (N_9860,N_7064,N_5958);
or U9861 (N_9861,N_7621,N_7625);
xnor U9862 (N_9862,N_7679,N_7372);
or U9863 (N_9863,N_5855,N_7358);
xor U9864 (N_9864,N_6631,N_6112);
or U9865 (N_9865,N_5663,N_6111);
nand U9866 (N_9866,N_6229,N_5801);
nor U9867 (N_9867,N_7993,N_7042);
nor U9868 (N_9868,N_5793,N_5686);
xnor U9869 (N_9869,N_6899,N_5640);
nand U9870 (N_9870,N_6322,N_4893);
or U9871 (N_9871,N_7593,N_4135);
or U9872 (N_9872,N_5172,N_7719);
or U9873 (N_9873,N_7205,N_4995);
xor U9874 (N_9874,N_4225,N_6793);
nand U9875 (N_9875,N_4901,N_6074);
and U9876 (N_9876,N_4711,N_5595);
and U9877 (N_9877,N_6416,N_6347);
and U9878 (N_9878,N_7413,N_5497);
or U9879 (N_9879,N_7365,N_5055);
nor U9880 (N_9880,N_4355,N_4446);
nor U9881 (N_9881,N_7422,N_6398);
and U9882 (N_9882,N_7559,N_7509);
xnor U9883 (N_9883,N_5996,N_4041);
nor U9884 (N_9884,N_5379,N_4765);
nand U9885 (N_9885,N_4329,N_4486);
or U9886 (N_9886,N_4258,N_6731);
nand U9887 (N_9887,N_7980,N_6046);
nor U9888 (N_9888,N_4485,N_6965);
xor U9889 (N_9889,N_4619,N_5179);
or U9890 (N_9890,N_5024,N_7952);
nor U9891 (N_9891,N_7562,N_6769);
and U9892 (N_9892,N_4288,N_6032);
and U9893 (N_9893,N_4753,N_6644);
or U9894 (N_9894,N_6002,N_5824);
or U9895 (N_9895,N_7702,N_7126);
xor U9896 (N_9896,N_4025,N_5351);
and U9897 (N_9897,N_4317,N_5705);
xor U9898 (N_9898,N_6578,N_5295);
nand U9899 (N_9899,N_4442,N_7863);
nor U9900 (N_9900,N_6948,N_6103);
or U9901 (N_9901,N_6421,N_7736);
nand U9902 (N_9902,N_4287,N_6583);
nor U9903 (N_9903,N_7016,N_7914);
nor U9904 (N_9904,N_5912,N_4637);
nand U9905 (N_9905,N_6342,N_4052);
nor U9906 (N_9906,N_7944,N_7728);
xor U9907 (N_9907,N_5656,N_5896);
and U9908 (N_9908,N_4537,N_6495);
or U9909 (N_9909,N_4723,N_5085);
or U9910 (N_9910,N_4839,N_6651);
nor U9911 (N_9911,N_4309,N_5464);
xor U9912 (N_9912,N_7248,N_4902);
and U9913 (N_9913,N_7664,N_6498);
xor U9914 (N_9914,N_5069,N_5053);
and U9915 (N_9915,N_7048,N_4228);
nand U9916 (N_9916,N_5375,N_7755);
xnor U9917 (N_9917,N_5062,N_7548);
and U9918 (N_9918,N_7009,N_5326);
or U9919 (N_9919,N_7795,N_4744);
nand U9920 (N_9920,N_6765,N_6886);
nand U9921 (N_9921,N_5737,N_5057);
xor U9922 (N_9922,N_6235,N_7947);
nor U9923 (N_9923,N_7229,N_4426);
and U9924 (N_9924,N_5287,N_5901);
or U9925 (N_9925,N_4558,N_6903);
or U9926 (N_9926,N_5563,N_5432);
nand U9927 (N_9927,N_6928,N_6016);
nor U9928 (N_9928,N_4842,N_7221);
and U9929 (N_9929,N_7065,N_4885);
nand U9930 (N_9930,N_7704,N_6722);
nor U9931 (N_9931,N_4250,N_5046);
and U9932 (N_9932,N_4149,N_7968);
nor U9933 (N_9933,N_7389,N_4641);
nor U9934 (N_9934,N_5713,N_5266);
nor U9935 (N_9935,N_7494,N_7723);
xor U9936 (N_9936,N_5744,N_4284);
nor U9937 (N_9937,N_6612,N_5144);
and U9938 (N_9938,N_4322,N_4324);
or U9939 (N_9939,N_5981,N_6140);
nor U9940 (N_9940,N_5836,N_5619);
nand U9941 (N_9941,N_7674,N_5474);
xnor U9942 (N_9942,N_4731,N_6305);
nor U9943 (N_9943,N_7092,N_6720);
nor U9944 (N_9944,N_5034,N_4158);
or U9945 (N_9945,N_5185,N_7884);
xor U9946 (N_9946,N_7105,N_6521);
or U9947 (N_9947,N_4710,N_7940);
and U9948 (N_9948,N_5641,N_6426);
and U9949 (N_9949,N_5578,N_7379);
nand U9950 (N_9950,N_5265,N_7057);
and U9951 (N_9951,N_4055,N_4872);
nor U9952 (N_9952,N_6313,N_7175);
or U9953 (N_9953,N_5052,N_5441);
nor U9954 (N_9954,N_4829,N_7188);
and U9955 (N_9955,N_6558,N_7089);
nand U9956 (N_9956,N_4244,N_7837);
nand U9957 (N_9957,N_7694,N_7716);
or U9958 (N_9958,N_6555,N_7500);
or U9959 (N_9959,N_6015,N_6200);
and U9960 (N_9960,N_6607,N_5564);
and U9961 (N_9961,N_4680,N_6980);
nand U9962 (N_9962,N_4325,N_4565);
nor U9963 (N_9963,N_4044,N_4337);
or U9964 (N_9964,N_4544,N_6266);
or U9965 (N_9965,N_7879,N_4110);
or U9966 (N_9966,N_4274,N_7669);
xor U9967 (N_9967,N_4304,N_5091);
nand U9968 (N_9968,N_4630,N_6467);
or U9969 (N_9969,N_5711,N_4621);
and U9970 (N_9970,N_7363,N_5407);
and U9971 (N_9971,N_7036,N_6527);
nand U9972 (N_9972,N_7454,N_5230);
and U9973 (N_9973,N_7767,N_6624);
nor U9974 (N_9974,N_4248,N_6841);
xor U9975 (N_9975,N_4239,N_4536);
nor U9976 (N_9976,N_6133,N_4488);
or U9977 (N_9977,N_6668,N_4240);
or U9978 (N_9978,N_6170,N_6405);
nor U9979 (N_9979,N_4827,N_4703);
nor U9980 (N_9980,N_6144,N_7583);
nand U9981 (N_9981,N_4582,N_4091);
and U9982 (N_9982,N_4428,N_6464);
and U9983 (N_9983,N_6020,N_5976);
xor U9984 (N_9984,N_7090,N_5139);
and U9985 (N_9985,N_4042,N_5116);
nor U9986 (N_9986,N_7737,N_7794);
nor U9987 (N_9987,N_5068,N_6228);
nand U9988 (N_9988,N_6445,N_4896);
and U9989 (N_9989,N_4812,N_5193);
nand U9990 (N_9990,N_7038,N_6167);
and U9991 (N_9991,N_7868,N_6450);
nor U9992 (N_9992,N_6529,N_4420);
nor U9993 (N_9993,N_6688,N_7869);
xor U9994 (N_9994,N_4131,N_7037);
xor U9995 (N_9995,N_7131,N_6988);
and U9996 (N_9996,N_7265,N_7435);
xnor U9997 (N_9997,N_7353,N_7659);
and U9998 (N_9998,N_5246,N_4851);
nor U9999 (N_9999,N_4601,N_4430);
nand U10000 (N_10000,N_7420,N_7635);
and U10001 (N_10001,N_5415,N_7125);
nand U10002 (N_10002,N_7663,N_5532);
xor U10003 (N_10003,N_5745,N_5904);
and U10004 (N_10004,N_6125,N_5237);
and U10005 (N_10005,N_5812,N_7952);
nor U10006 (N_10006,N_5416,N_4019);
nor U10007 (N_10007,N_5321,N_7581);
xnor U10008 (N_10008,N_5672,N_5743);
and U10009 (N_10009,N_7524,N_4279);
nor U10010 (N_10010,N_4161,N_4870);
and U10011 (N_10011,N_5157,N_5895);
nor U10012 (N_10012,N_5946,N_7898);
and U10013 (N_10013,N_4464,N_7762);
or U10014 (N_10014,N_4707,N_6554);
and U10015 (N_10015,N_4460,N_7609);
and U10016 (N_10016,N_6923,N_6304);
nor U10017 (N_10017,N_5718,N_7868);
nand U10018 (N_10018,N_7138,N_7820);
xor U10019 (N_10019,N_6952,N_6826);
nor U10020 (N_10020,N_5145,N_5674);
nand U10021 (N_10021,N_7461,N_4350);
or U10022 (N_10022,N_7617,N_7022);
and U10023 (N_10023,N_5736,N_5391);
nor U10024 (N_10024,N_4056,N_7184);
and U10025 (N_10025,N_4919,N_7178);
nor U10026 (N_10026,N_7744,N_6540);
or U10027 (N_10027,N_7187,N_5333);
nor U10028 (N_10028,N_6240,N_6569);
and U10029 (N_10029,N_7790,N_5848);
nor U10030 (N_10030,N_4734,N_5537);
nor U10031 (N_10031,N_6795,N_6852);
nand U10032 (N_10032,N_7205,N_4262);
and U10033 (N_10033,N_4560,N_4539);
xor U10034 (N_10034,N_7055,N_6813);
nor U10035 (N_10035,N_7792,N_6497);
nand U10036 (N_10036,N_6908,N_5551);
xor U10037 (N_10037,N_5994,N_6338);
nor U10038 (N_10038,N_7048,N_4066);
nor U10039 (N_10039,N_5231,N_4986);
nor U10040 (N_10040,N_7396,N_6175);
xnor U10041 (N_10041,N_7686,N_4582);
nand U10042 (N_10042,N_5436,N_4360);
or U10043 (N_10043,N_7346,N_6251);
xor U10044 (N_10044,N_7481,N_4636);
or U10045 (N_10045,N_4744,N_7448);
or U10046 (N_10046,N_5614,N_4073);
xnor U10047 (N_10047,N_6445,N_6048);
xor U10048 (N_10048,N_4599,N_6732);
nand U10049 (N_10049,N_4351,N_6141);
xnor U10050 (N_10050,N_4264,N_7856);
nor U10051 (N_10051,N_4112,N_6074);
and U10052 (N_10052,N_4241,N_5181);
xor U10053 (N_10053,N_5550,N_5868);
nand U10054 (N_10054,N_4536,N_5106);
nor U10055 (N_10055,N_6622,N_5289);
xnor U10056 (N_10056,N_4849,N_5038);
or U10057 (N_10057,N_4711,N_5124);
or U10058 (N_10058,N_6983,N_7487);
nand U10059 (N_10059,N_6852,N_4532);
nand U10060 (N_10060,N_6574,N_6682);
nor U10061 (N_10061,N_6325,N_5544);
and U10062 (N_10062,N_6283,N_4461);
xnor U10063 (N_10063,N_5991,N_6874);
or U10064 (N_10064,N_4398,N_5665);
nor U10065 (N_10065,N_7938,N_7870);
xor U10066 (N_10066,N_5676,N_4268);
nor U10067 (N_10067,N_6877,N_7490);
and U10068 (N_10068,N_5438,N_4225);
nor U10069 (N_10069,N_7868,N_7710);
or U10070 (N_10070,N_4930,N_5506);
or U10071 (N_10071,N_6096,N_7678);
xor U10072 (N_10072,N_7647,N_5120);
nand U10073 (N_10073,N_7900,N_5208);
and U10074 (N_10074,N_7547,N_4108);
and U10075 (N_10075,N_7589,N_4477);
and U10076 (N_10076,N_7713,N_4414);
and U10077 (N_10077,N_5774,N_7207);
nor U10078 (N_10078,N_7989,N_5484);
or U10079 (N_10079,N_4059,N_7417);
and U10080 (N_10080,N_7757,N_7323);
or U10081 (N_10081,N_4590,N_6270);
or U10082 (N_10082,N_5748,N_5977);
nor U10083 (N_10083,N_5927,N_6836);
nand U10084 (N_10084,N_7864,N_4969);
nor U10085 (N_10085,N_4831,N_6845);
nor U10086 (N_10086,N_5611,N_7721);
xor U10087 (N_10087,N_7030,N_5086);
nand U10088 (N_10088,N_4525,N_4082);
xnor U10089 (N_10089,N_7923,N_5380);
xnor U10090 (N_10090,N_6715,N_5887);
xnor U10091 (N_10091,N_4520,N_5023);
xor U10092 (N_10092,N_4016,N_4524);
nand U10093 (N_10093,N_4190,N_5246);
or U10094 (N_10094,N_5203,N_6511);
and U10095 (N_10095,N_7474,N_7465);
and U10096 (N_10096,N_4726,N_7585);
and U10097 (N_10097,N_6253,N_4735);
nor U10098 (N_10098,N_7226,N_4780);
or U10099 (N_10099,N_5787,N_7949);
xnor U10100 (N_10100,N_7721,N_5009);
xor U10101 (N_10101,N_6366,N_4325);
and U10102 (N_10102,N_7454,N_4528);
nand U10103 (N_10103,N_4390,N_5363);
nand U10104 (N_10104,N_5503,N_4998);
nand U10105 (N_10105,N_6128,N_7452);
or U10106 (N_10106,N_7539,N_7800);
and U10107 (N_10107,N_5309,N_4286);
and U10108 (N_10108,N_4091,N_7811);
nand U10109 (N_10109,N_6003,N_7544);
nand U10110 (N_10110,N_7619,N_4996);
xor U10111 (N_10111,N_7742,N_4648);
nand U10112 (N_10112,N_6016,N_7419);
or U10113 (N_10113,N_6279,N_7406);
nand U10114 (N_10114,N_7577,N_4602);
nor U10115 (N_10115,N_5443,N_5477);
and U10116 (N_10116,N_6985,N_4948);
or U10117 (N_10117,N_5405,N_4301);
nand U10118 (N_10118,N_4836,N_6086);
xor U10119 (N_10119,N_4605,N_6769);
xnor U10120 (N_10120,N_4361,N_7602);
nand U10121 (N_10121,N_6967,N_7615);
nand U10122 (N_10122,N_6243,N_4350);
or U10123 (N_10123,N_5564,N_4898);
xnor U10124 (N_10124,N_4341,N_6776);
nand U10125 (N_10125,N_4525,N_4651);
and U10126 (N_10126,N_5053,N_7095);
nor U10127 (N_10127,N_4490,N_4507);
and U10128 (N_10128,N_6034,N_4049);
or U10129 (N_10129,N_6534,N_4728);
nor U10130 (N_10130,N_5113,N_4314);
or U10131 (N_10131,N_4055,N_6938);
nor U10132 (N_10132,N_6498,N_5805);
or U10133 (N_10133,N_5988,N_7790);
or U10134 (N_10134,N_4709,N_6672);
xor U10135 (N_10135,N_6207,N_7217);
or U10136 (N_10136,N_7226,N_5990);
xor U10137 (N_10137,N_5526,N_6062);
xnor U10138 (N_10138,N_7013,N_7918);
and U10139 (N_10139,N_7097,N_6141);
nor U10140 (N_10140,N_4012,N_5186);
nand U10141 (N_10141,N_5069,N_4539);
or U10142 (N_10142,N_6835,N_7782);
xnor U10143 (N_10143,N_4184,N_5474);
nor U10144 (N_10144,N_7821,N_6392);
nand U10145 (N_10145,N_7358,N_5697);
and U10146 (N_10146,N_7277,N_7255);
and U10147 (N_10147,N_4339,N_5640);
nor U10148 (N_10148,N_7000,N_5085);
or U10149 (N_10149,N_4887,N_5137);
nand U10150 (N_10150,N_5833,N_5358);
or U10151 (N_10151,N_4374,N_5884);
xnor U10152 (N_10152,N_5621,N_5458);
xor U10153 (N_10153,N_4620,N_5613);
or U10154 (N_10154,N_6445,N_4448);
or U10155 (N_10155,N_5459,N_4053);
xor U10156 (N_10156,N_5290,N_6877);
nor U10157 (N_10157,N_6434,N_5099);
or U10158 (N_10158,N_7945,N_6334);
nor U10159 (N_10159,N_6696,N_7018);
nand U10160 (N_10160,N_7918,N_4300);
and U10161 (N_10161,N_5924,N_6204);
nand U10162 (N_10162,N_7591,N_5328);
xnor U10163 (N_10163,N_4336,N_5856);
nand U10164 (N_10164,N_4481,N_6170);
nor U10165 (N_10165,N_5112,N_6660);
or U10166 (N_10166,N_6106,N_5703);
nand U10167 (N_10167,N_5014,N_7351);
and U10168 (N_10168,N_5095,N_6443);
nand U10169 (N_10169,N_4693,N_4401);
xor U10170 (N_10170,N_6470,N_7740);
nand U10171 (N_10171,N_7889,N_6212);
and U10172 (N_10172,N_4784,N_6721);
and U10173 (N_10173,N_7541,N_6904);
nor U10174 (N_10174,N_7716,N_7598);
nand U10175 (N_10175,N_5900,N_4922);
xor U10176 (N_10176,N_4669,N_5596);
nand U10177 (N_10177,N_4744,N_7586);
nand U10178 (N_10178,N_4094,N_5227);
nor U10179 (N_10179,N_5931,N_4758);
and U10180 (N_10180,N_6121,N_4641);
nand U10181 (N_10181,N_5134,N_4896);
nand U10182 (N_10182,N_5825,N_6005);
and U10183 (N_10183,N_7077,N_7934);
xnor U10184 (N_10184,N_4945,N_6630);
xnor U10185 (N_10185,N_5996,N_4359);
xor U10186 (N_10186,N_6206,N_6630);
nand U10187 (N_10187,N_7671,N_6991);
nor U10188 (N_10188,N_4764,N_4378);
nor U10189 (N_10189,N_7694,N_6742);
nor U10190 (N_10190,N_7224,N_6889);
or U10191 (N_10191,N_7389,N_7789);
xnor U10192 (N_10192,N_4955,N_4766);
xnor U10193 (N_10193,N_6512,N_5044);
xnor U10194 (N_10194,N_7089,N_7948);
nor U10195 (N_10195,N_4070,N_5570);
and U10196 (N_10196,N_5576,N_7092);
nand U10197 (N_10197,N_4525,N_6824);
nor U10198 (N_10198,N_5949,N_5260);
nand U10199 (N_10199,N_7353,N_6201);
nand U10200 (N_10200,N_4090,N_6673);
or U10201 (N_10201,N_4397,N_4736);
and U10202 (N_10202,N_6439,N_7430);
or U10203 (N_10203,N_5934,N_7117);
nor U10204 (N_10204,N_5193,N_5603);
and U10205 (N_10205,N_4278,N_6105);
or U10206 (N_10206,N_5777,N_7966);
and U10207 (N_10207,N_4368,N_4371);
or U10208 (N_10208,N_4473,N_4476);
xnor U10209 (N_10209,N_4965,N_5864);
xor U10210 (N_10210,N_6652,N_6446);
and U10211 (N_10211,N_5307,N_7173);
nor U10212 (N_10212,N_4069,N_4527);
or U10213 (N_10213,N_5545,N_5620);
and U10214 (N_10214,N_7196,N_7019);
or U10215 (N_10215,N_4622,N_5735);
nand U10216 (N_10216,N_5056,N_7233);
nand U10217 (N_10217,N_5625,N_7068);
or U10218 (N_10218,N_4008,N_6785);
nand U10219 (N_10219,N_6542,N_5209);
xor U10220 (N_10220,N_4437,N_7334);
or U10221 (N_10221,N_7112,N_5896);
xnor U10222 (N_10222,N_6809,N_5274);
or U10223 (N_10223,N_6395,N_4416);
xnor U10224 (N_10224,N_6519,N_7225);
or U10225 (N_10225,N_7553,N_4266);
or U10226 (N_10226,N_4145,N_5953);
or U10227 (N_10227,N_6377,N_6789);
nand U10228 (N_10228,N_7201,N_5436);
xor U10229 (N_10229,N_7902,N_7540);
nand U10230 (N_10230,N_7431,N_6369);
xnor U10231 (N_10231,N_4913,N_5276);
xor U10232 (N_10232,N_4063,N_7163);
xnor U10233 (N_10233,N_6943,N_4638);
and U10234 (N_10234,N_6689,N_6917);
nor U10235 (N_10235,N_7895,N_7260);
nand U10236 (N_10236,N_7488,N_5373);
nand U10237 (N_10237,N_5933,N_4502);
xor U10238 (N_10238,N_6145,N_6528);
xnor U10239 (N_10239,N_7647,N_5395);
nor U10240 (N_10240,N_4926,N_5095);
nor U10241 (N_10241,N_7991,N_5875);
or U10242 (N_10242,N_7205,N_6044);
xnor U10243 (N_10243,N_4024,N_4677);
nand U10244 (N_10244,N_5500,N_4960);
nand U10245 (N_10245,N_5545,N_4579);
and U10246 (N_10246,N_4841,N_4901);
nand U10247 (N_10247,N_6944,N_5616);
nor U10248 (N_10248,N_7158,N_6454);
nor U10249 (N_10249,N_7770,N_5903);
nor U10250 (N_10250,N_7475,N_6211);
nand U10251 (N_10251,N_4841,N_5020);
nand U10252 (N_10252,N_4502,N_7793);
nand U10253 (N_10253,N_6182,N_7860);
xor U10254 (N_10254,N_5918,N_7945);
nand U10255 (N_10255,N_7809,N_6844);
xnor U10256 (N_10256,N_6446,N_4984);
and U10257 (N_10257,N_6391,N_5535);
and U10258 (N_10258,N_6403,N_4299);
xnor U10259 (N_10259,N_5972,N_5085);
or U10260 (N_10260,N_5343,N_6870);
or U10261 (N_10261,N_6217,N_5751);
and U10262 (N_10262,N_4240,N_4744);
nor U10263 (N_10263,N_7954,N_7787);
and U10264 (N_10264,N_4361,N_7160);
nor U10265 (N_10265,N_4284,N_5226);
and U10266 (N_10266,N_5377,N_7578);
xor U10267 (N_10267,N_6886,N_5549);
nand U10268 (N_10268,N_7672,N_7588);
or U10269 (N_10269,N_7598,N_4254);
nand U10270 (N_10270,N_7395,N_5435);
or U10271 (N_10271,N_5941,N_6551);
nand U10272 (N_10272,N_7656,N_5532);
or U10273 (N_10273,N_6216,N_6122);
xnor U10274 (N_10274,N_7066,N_7206);
xnor U10275 (N_10275,N_7563,N_6217);
nor U10276 (N_10276,N_7264,N_4655);
nand U10277 (N_10277,N_5848,N_6650);
nor U10278 (N_10278,N_7631,N_7388);
and U10279 (N_10279,N_4387,N_6275);
nor U10280 (N_10280,N_5196,N_5308);
and U10281 (N_10281,N_4788,N_7335);
xor U10282 (N_10282,N_5313,N_4194);
nor U10283 (N_10283,N_4875,N_7302);
or U10284 (N_10284,N_4460,N_5541);
or U10285 (N_10285,N_7297,N_4472);
and U10286 (N_10286,N_5668,N_4140);
nor U10287 (N_10287,N_6600,N_7085);
nor U10288 (N_10288,N_5366,N_4183);
xnor U10289 (N_10289,N_5965,N_7444);
or U10290 (N_10290,N_5360,N_6060);
nor U10291 (N_10291,N_7459,N_4025);
and U10292 (N_10292,N_6659,N_4317);
nand U10293 (N_10293,N_5027,N_6980);
xnor U10294 (N_10294,N_4941,N_6953);
or U10295 (N_10295,N_6434,N_5643);
nand U10296 (N_10296,N_7403,N_7852);
nor U10297 (N_10297,N_4805,N_6118);
nand U10298 (N_10298,N_7394,N_5899);
nand U10299 (N_10299,N_6776,N_6104);
nand U10300 (N_10300,N_6663,N_6749);
xor U10301 (N_10301,N_5323,N_5349);
nor U10302 (N_10302,N_4710,N_7680);
nand U10303 (N_10303,N_5796,N_6718);
xor U10304 (N_10304,N_5574,N_5651);
nor U10305 (N_10305,N_7885,N_7310);
xor U10306 (N_10306,N_5549,N_7978);
nor U10307 (N_10307,N_5051,N_5117);
nand U10308 (N_10308,N_6411,N_7608);
or U10309 (N_10309,N_4839,N_6753);
nand U10310 (N_10310,N_7760,N_4072);
and U10311 (N_10311,N_7925,N_7990);
or U10312 (N_10312,N_5602,N_5088);
xnor U10313 (N_10313,N_7457,N_7950);
nand U10314 (N_10314,N_4516,N_7519);
and U10315 (N_10315,N_4838,N_7318);
and U10316 (N_10316,N_4202,N_5571);
nand U10317 (N_10317,N_7745,N_7537);
xnor U10318 (N_10318,N_4462,N_4343);
xor U10319 (N_10319,N_7814,N_6231);
or U10320 (N_10320,N_5924,N_4474);
or U10321 (N_10321,N_5628,N_6684);
or U10322 (N_10322,N_7586,N_5693);
nand U10323 (N_10323,N_6019,N_7789);
nand U10324 (N_10324,N_5183,N_6070);
xor U10325 (N_10325,N_6910,N_6122);
or U10326 (N_10326,N_4618,N_6212);
nand U10327 (N_10327,N_5455,N_5179);
nand U10328 (N_10328,N_4340,N_4237);
xnor U10329 (N_10329,N_4063,N_7364);
and U10330 (N_10330,N_4031,N_5893);
nor U10331 (N_10331,N_7097,N_7952);
nand U10332 (N_10332,N_4119,N_4130);
and U10333 (N_10333,N_7183,N_5491);
xnor U10334 (N_10334,N_4376,N_7152);
xor U10335 (N_10335,N_4394,N_7760);
and U10336 (N_10336,N_4222,N_5502);
nor U10337 (N_10337,N_4552,N_7358);
nand U10338 (N_10338,N_4142,N_4911);
nor U10339 (N_10339,N_5388,N_6991);
and U10340 (N_10340,N_5177,N_5200);
and U10341 (N_10341,N_6621,N_6799);
and U10342 (N_10342,N_7760,N_4630);
or U10343 (N_10343,N_4823,N_7430);
and U10344 (N_10344,N_4387,N_6517);
nor U10345 (N_10345,N_6907,N_7258);
and U10346 (N_10346,N_7229,N_7617);
or U10347 (N_10347,N_5615,N_6140);
or U10348 (N_10348,N_5603,N_7621);
nand U10349 (N_10349,N_6730,N_4862);
xnor U10350 (N_10350,N_7595,N_5685);
and U10351 (N_10351,N_5137,N_4124);
nand U10352 (N_10352,N_5001,N_6133);
nand U10353 (N_10353,N_6570,N_6270);
nand U10354 (N_10354,N_6685,N_5336);
xnor U10355 (N_10355,N_4412,N_7971);
nand U10356 (N_10356,N_7006,N_6274);
or U10357 (N_10357,N_4880,N_6432);
and U10358 (N_10358,N_6602,N_7756);
nand U10359 (N_10359,N_6284,N_7484);
and U10360 (N_10360,N_4277,N_5067);
xor U10361 (N_10361,N_4643,N_7463);
nor U10362 (N_10362,N_6780,N_7314);
and U10363 (N_10363,N_6219,N_4458);
nor U10364 (N_10364,N_4265,N_5764);
nor U10365 (N_10365,N_4380,N_6816);
or U10366 (N_10366,N_5663,N_6163);
nand U10367 (N_10367,N_5489,N_5619);
nor U10368 (N_10368,N_5000,N_5040);
and U10369 (N_10369,N_4939,N_7259);
nor U10370 (N_10370,N_5687,N_6386);
and U10371 (N_10371,N_6385,N_6112);
xnor U10372 (N_10372,N_6885,N_7460);
nor U10373 (N_10373,N_5261,N_6180);
or U10374 (N_10374,N_7129,N_5929);
nor U10375 (N_10375,N_7107,N_4569);
xor U10376 (N_10376,N_5822,N_6408);
nor U10377 (N_10377,N_7780,N_4718);
nor U10378 (N_10378,N_4135,N_6715);
or U10379 (N_10379,N_7142,N_4998);
nand U10380 (N_10380,N_4685,N_5068);
xor U10381 (N_10381,N_7095,N_6802);
nor U10382 (N_10382,N_6864,N_7150);
and U10383 (N_10383,N_7821,N_5223);
and U10384 (N_10384,N_7569,N_7410);
nand U10385 (N_10385,N_5153,N_6826);
nor U10386 (N_10386,N_4645,N_7315);
xnor U10387 (N_10387,N_6904,N_4930);
nand U10388 (N_10388,N_6239,N_7036);
nand U10389 (N_10389,N_4763,N_5988);
nor U10390 (N_10390,N_6088,N_4723);
nand U10391 (N_10391,N_4644,N_6285);
and U10392 (N_10392,N_7946,N_5892);
and U10393 (N_10393,N_4385,N_4238);
and U10394 (N_10394,N_4944,N_4844);
or U10395 (N_10395,N_7165,N_4919);
xnor U10396 (N_10396,N_4437,N_4062);
or U10397 (N_10397,N_5052,N_5246);
or U10398 (N_10398,N_7661,N_5237);
or U10399 (N_10399,N_5866,N_5947);
xnor U10400 (N_10400,N_5557,N_6202);
xnor U10401 (N_10401,N_6221,N_7149);
nor U10402 (N_10402,N_4954,N_6419);
nand U10403 (N_10403,N_6566,N_6194);
or U10404 (N_10404,N_6873,N_6521);
or U10405 (N_10405,N_4080,N_5669);
or U10406 (N_10406,N_4214,N_4289);
and U10407 (N_10407,N_5205,N_7650);
and U10408 (N_10408,N_7369,N_7467);
xnor U10409 (N_10409,N_7014,N_4746);
and U10410 (N_10410,N_7400,N_5681);
nor U10411 (N_10411,N_4692,N_6915);
xor U10412 (N_10412,N_6388,N_6381);
xnor U10413 (N_10413,N_5542,N_5070);
nand U10414 (N_10414,N_7346,N_7508);
and U10415 (N_10415,N_5451,N_5882);
or U10416 (N_10416,N_4061,N_6072);
and U10417 (N_10417,N_7672,N_6977);
and U10418 (N_10418,N_4232,N_7972);
nor U10419 (N_10419,N_5694,N_4002);
xor U10420 (N_10420,N_4671,N_7074);
and U10421 (N_10421,N_4654,N_5755);
nand U10422 (N_10422,N_5630,N_7488);
and U10423 (N_10423,N_7767,N_7309);
and U10424 (N_10424,N_7599,N_7865);
nand U10425 (N_10425,N_4265,N_4295);
nand U10426 (N_10426,N_4890,N_7766);
nor U10427 (N_10427,N_4037,N_5169);
nand U10428 (N_10428,N_7195,N_7546);
or U10429 (N_10429,N_5448,N_6499);
xnor U10430 (N_10430,N_7030,N_4413);
nand U10431 (N_10431,N_6556,N_6871);
nor U10432 (N_10432,N_5447,N_6086);
or U10433 (N_10433,N_6128,N_5036);
nor U10434 (N_10434,N_5553,N_4058);
nand U10435 (N_10435,N_4403,N_4921);
nand U10436 (N_10436,N_6614,N_6602);
xnor U10437 (N_10437,N_5651,N_4600);
or U10438 (N_10438,N_5946,N_6028);
and U10439 (N_10439,N_7584,N_4843);
nand U10440 (N_10440,N_5834,N_6120);
and U10441 (N_10441,N_6111,N_7501);
xnor U10442 (N_10442,N_6946,N_5419);
and U10443 (N_10443,N_7846,N_7186);
nand U10444 (N_10444,N_7928,N_5983);
and U10445 (N_10445,N_5773,N_6872);
nor U10446 (N_10446,N_7555,N_6672);
nand U10447 (N_10447,N_6941,N_7815);
or U10448 (N_10448,N_7105,N_5761);
nand U10449 (N_10449,N_7279,N_5225);
and U10450 (N_10450,N_6542,N_7664);
nand U10451 (N_10451,N_5750,N_6204);
nand U10452 (N_10452,N_5345,N_6590);
nor U10453 (N_10453,N_6146,N_5391);
nand U10454 (N_10454,N_6737,N_7790);
or U10455 (N_10455,N_6984,N_4962);
and U10456 (N_10456,N_7979,N_5324);
nand U10457 (N_10457,N_4776,N_4004);
xnor U10458 (N_10458,N_5280,N_4123);
nor U10459 (N_10459,N_5833,N_6860);
nand U10460 (N_10460,N_6911,N_7536);
xor U10461 (N_10461,N_5508,N_5320);
nor U10462 (N_10462,N_5558,N_4677);
nand U10463 (N_10463,N_6415,N_4589);
nand U10464 (N_10464,N_6591,N_5388);
nor U10465 (N_10465,N_7068,N_7542);
nand U10466 (N_10466,N_7899,N_5393);
xnor U10467 (N_10467,N_7383,N_5368);
or U10468 (N_10468,N_5732,N_7359);
xor U10469 (N_10469,N_4614,N_7567);
and U10470 (N_10470,N_5342,N_7833);
and U10471 (N_10471,N_4914,N_5306);
and U10472 (N_10472,N_5842,N_7116);
xor U10473 (N_10473,N_6127,N_4430);
nand U10474 (N_10474,N_6220,N_7057);
nand U10475 (N_10475,N_6065,N_7112);
nand U10476 (N_10476,N_7917,N_6633);
and U10477 (N_10477,N_6874,N_5955);
xnor U10478 (N_10478,N_5822,N_7021);
nor U10479 (N_10479,N_6141,N_6547);
nor U10480 (N_10480,N_4258,N_7743);
and U10481 (N_10481,N_5491,N_6923);
nor U10482 (N_10482,N_6367,N_6486);
nand U10483 (N_10483,N_6906,N_7015);
and U10484 (N_10484,N_4676,N_6981);
nor U10485 (N_10485,N_5949,N_6901);
nor U10486 (N_10486,N_6726,N_4921);
nor U10487 (N_10487,N_6373,N_4882);
nor U10488 (N_10488,N_6477,N_4095);
nand U10489 (N_10489,N_4884,N_7020);
xnor U10490 (N_10490,N_6528,N_5669);
nand U10491 (N_10491,N_5522,N_5441);
xnor U10492 (N_10492,N_4199,N_7296);
nand U10493 (N_10493,N_6890,N_6309);
and U10494 (N_10494,N_4570,N_5036);
nor U10495 (N_10495,N_6883,N_4152);
and U10496 (N_10496,N_7509,N_7642);
or U10497 (N_10497,N_5207,N_7742);
xnor U10498 (N_10498,N_7472,N_6726);
or U10499 (N_10499,N_4060,N_5246);
nand U10500 (N_10500,N_4211,N_5402);
nor U10501 (N_10501,N_6281,N_7910);
xnor U10502 (N_10502,N_5661,N_6827);
and U10503 (N_10503,N_4398,N_7860);
nor U10504 (N_10504,N_5419,N_4289);
and U10505 (N_10505,N_7792,N_5679);
xor U10506 (N_10506,N_6170,N_5553);
or U10507 (N_10507,N_4657,N_4228);
and U10508 (N_10508,N_6167,N_6804);
nand U10509 (N_10509,N_7029,N_5041);
nand U10510 (N_10510,N_7988,N_6149);
xnor U10511 (N_10511,N_5211,N_6122);
or U10512 (N_10512,N_4549,N_6526);
nor U10513 (N_10513,N_5327,N_6582);
nor U10514 (N_10514,N_5002,N_6806);
nor U10515 (N_10515,N_5529,N_4247);
nor U10516 (N_10516,N_7770,N_6080);
or U10517 (N_10517,N_5891,N_7192);
nand U10518 (N_10518,N_4128,N_4392);
xnor U10519 (N_10519,N_6468,N_4836);
xor U10520 (N_10520,N_5097,N_7320);
or U10521 (N_10521,N_6597,N_7852);
or U10522 (N_10522,N_5963,N_5401);
xnor U10523 (N_10523,N_6991,N_5862);
nand U10524 (N_10524,N_5502,N_4075);
nand U10525 (N_10525,N_5978,N_4481);
nand U10526 (N_10526,N_6680,N_6349);
xor U10527 (N_10527,N_7155,N_6095);
or U10528 (N_10528,N_5841,N_6212);
xnor U10529 (N_10529,N_6172,N_5820);
xor U10530 (N_10530,N_7597,N_7240);
nand U10531 (N_10531,N_7155,N_7308);
nand U10532 (N_10532,N_5996,N_7919);
and U10533 (N_10533,N_7689,N_4232);
or U10534 (N_10534,N_7338,N_4843);
nor U10535 (N_10535,N_4150,N_4105);
or U10536 (N_10536,N_5008,N_7444);
nor U10537 (N_10537,N_6295,N_5405);
xor U10538 (N_10538,N_7410,N_6496);
and U10539 (N_10539,N_5526,N_7699);
nand U10540 (N_10540,N_5845,N_4664);
xor U10541 (N_10541,N_7152,N_4187);
and U10542 (N_10542,N_7516,N_7892);
and U10543 (N_10543,N_7200,N_7191);
xor U10544 (N_10544,N_6204,N_6933);
xnor U10545 (N_10545,N_4438,N_4696);
xor U10546 (N_10546,N_7023,N_4616);
nand U10547 (N_10547,N_7046,N_4256);
and U10548 (N_10548,N_4175,N_7787);
xor U10549 (N_10549,N_7026,N_4533);
or U10550 (N_10550,N_5493,N_4037);
xor U10551 (N_10551,N_7196,N_6366);
or U10552 (N_10552,N_4792,N_6837);
xnor U10553 (N_10553,N_7580,N_6250);
or U10554 (N_10554,N_7519,N_7285);
nand U10555 (N_10555,N_7448,N_6236);
nor U10556 (N_10556,N_7396,N_5825);
nor U10557 (N_10557,N_6792,N_7013);
or U10558 (N_10558,N_5803,N_7764);
or U10559 (N_10559,N_5442,N_5283);
or U10560 (N_10560,N_4157,N_5696);
or U10561 (N_10561,N_6614,N_5942);
and U10562 (N_10562,N_7422,N_7723);
or U10563 (N_10563,N_6836,N_7795);
xor U10564 (N_10564,N_7885,N_5976);
nor U10565 (N_10565,N_6430,N_4298);
xor U10566 (N_10566,N_6669,N_5940);
nor U10567 (N_10567,N_7562,N_5595);
nor U10568 (N_10568,N_6047,N_4811);
xor U10569 (N_10569,N_4349,N_5181);
or U10570 (N_10570,N_7858,N_7925);
or U10571 (N_10571,N_6613,N_4624);
or U10572 (N_10572,N_4501,N_6988);
or U10573 (N_10573,N_4459,N_7670);
and U10574 (N_10574,N_6675,N_7695);
xnor U10575 (N_10575,N_7616,N_4400);
or U10576 (N_10576,N_5419,N_5749);
xnor U10577 (N_10577,N_7780,N_6054);
and U10578 (N_10578,N_4936,N_4343);
nor U10579 (N_10579,N_6630,N_7649);
xor U10580 (N_10580,N_5311,N_5882);
nor U10581 (N_10581,N_4812,N_4837);
xnor U10582 (N_10582,N_7699,N_5243);
and U10583 (N_10583,N_5466,N_5757);
nor U10584 (N_10584,N_4021,N_5467);
and U10585 (N_10585,N_6498,N_6826);
or U10586 (N_10586,N_6567,N_5291);
xor U10587 (N_10587,N_7732,N_5190);
xor U10588 (N_10588,N_6322,N_4422);
and U10589 (N_10589,N_6694,N_4928);
and U10590 (N_10590,N_4744,N_5412);
xor U10591 (N_10591,N_4073,N_7324);
xor U10592 (N_10592,N_4597,N_5812);
nor U10593 (N_10593,N_4084,N_7971);
nor U10594 (N_10594,N_7710,N_6383);
xnor U10595 (N_10595,N_4479,N_6900);
nor U10596 (N_10596,N_6508,N_4162);
and U10597 (N_10597,N_7130,N_6725);
and U10598 (N_10598,N_4747,N_7679);
or U10599 (N_10599,N_7175,N_4071);
nor U10600 (N_10600,N_4333,N_7133);
or U10601 (N_10601,N_5100,N_6187);
nand U10602 (N_10602,N_7443,N_4354);
nand U10603 (N_10603,N_7090,N_6576);
nand U10604 (N_10604,N_5395,N_6379);
xor U10605 (N_10605,N_4529,N_4033);
nor U10606 (N_10606,N_4181,N_7832);
nand U10607 (N_10607,N_6527,N_5717);
and U10608 (N_10608,N_7793,N_7282);
xnor U10609 (N_10609,N_7736,N_6545);
xor U10610 (N_10610,N_5181,N_5188);
xor U10611 (N_10611,N_4451,N_6172);
nand U10612 (N_10612,N_7355,N_5362);
and U10613 (N_10613,N_6306,N_6373);
or U10614 (N_10614,N_5003,N_5234);
nand U10615 (N_10615,N_4065,N_7932);
nor U10616 (N_10616,N_6844,N_6612);
nand U10617 (N_10617,N_7720,N_6937);
nor U10618 (N_10618,N_4769,N_6298);
or U10619 (N_10619,N_5756,N_7261);
or U10620 (N_10620,N_5118,N_7513);
or U10621 (N_10621,N_7310,N_7592);
nand U10622 (N_10622,N_5868,N_5431);
nor U10623 (N_10623,N_4697,N_5294);
nor U10624 (N_10624,N_7091,N_7217);
nand U10625 (N_10625,N_6964,N_5670);
xnor U10626 (N_10626,N_5107,N_7481);
nand U10627 (N_10627,N_7276,N_7058);
and U10628 (N_10628,N_5831,N_7144);
nand U10629 (N_10629,N_6168,N_4292);
nor U10630 (N_10630,N_6527,N_5515);
nor U10631 (N_10631,N_7877,N_6298);
nand U10632 (N_10632,N_5913,N_6184);
or U10633 (N_10633,N_4600,N_6864);
or U10634 (N_10634,N_5945,N_4796);
xor U10635 (N_10635,N_7524,N_4843);
nor U10636 (N_10636,N_6798,N_5997);
nand U10637 (N_10637,N_4584,N_7982);
or U10638 (N_10638,N_4003,N_4676);
and U10639 (N_10639,N_7736,N_5498);
nor U10640 (N_10640,N_6641,N_5255);
xor U10641 (N_10641,N_7066,N_5286);
and U10642 (N_10642,N_5259,N_4240);
nand U10643 (N_10643,N_5170,N_4014);
nor U10644 (N_10644,N_4770,N_7056);
xnor U10645 (N_10645,N_4899,N_6269);
nor U10646 (N_10646,N_4964,N_6945);
or U10647 (N_10647,N_7932,N_6389);
and U10648 (N_10648,N_6430,N_4882);
and U10649 (N_10649,N_4190,N_6574);
xnor U10650 (N_10650,N_5791,N_5299);
xor U10651 (N_10651,N_6625,N_7162);
xnor U10652 (N_10652,N_5893,N_5007);
nand U10653 (N_10653,N_7221,N_6063);
or U10654 (N_10654,N_4537,N_6960);
xor U10655 (N_10655,N_6608,N_6346);
nand U10656 (N_10656,N_4163,N_5013);
or U10657 (N_10657,N_5981,N_7334);
nor U10658 (N_10658,N_6221,N_6563);
nand U10659 (N_10659,N_6280,N_4052);
xor U10660 (N_10660,N_6791,N_7440);
and U10661 (N_10661,N_5331,N_5342);
or U10662 (N_10662,N_7773,N_6996);
nand U10663 (N_10663,N_5763,N_6297);
or U10664 (N_10664,N_6229,N_7266);
and U10665 (N_10665,N_5802,N_6309);
or U10666 (N_10666,N_5398,N_4065);
or U10667 (N_10667,N_5131,N_7922);
nand U10668 (N_10668,N_4964,N_6117);
nor U10669 (N_10669,N_6761,N_4587);
nor U10670 (N_10670,N_4497,N_4686);
nor U10671 (N_10671,N_5769,N_5690);
nor U10672 (N_10672,N_6460,N_4093);
nor U10673 (N_10673,N_6710,N_4623);
nor U10674 (N_10674,N_7881,N_7866);
and U10675 (N_10675,N_5623,N_6719);
or U10676 (N_10676,N_7842,N_5442);
xor U10677 (N_10677,N_7536,N_5538);
xnor U10678 (N_10678,N_5543,N_5019);
xnor U10679 (N_10679,N_4997,N_6747);
nand U10680 (N_10680,N_7338,N_4331);
xor U10681 (N_10681,N_4625,N_4776);
xnor U10682 (N_10682,N_7076,N_6388);
nand U10683 (N_10683,N_7968,N_4625);
nand U10684 (N_10684,N_5014,N_5340);
and U10685 (N_10685,N_7345,N_5684);
xnor U10686 (N_10686,N_5462,N_5658);
and U10687 (N_10687,N_6711,N_7679);
nor U10688 (N_10688,N_4883,N_4464);
or U10689 (N_10689,N_6966,N_5878);
or U10690 (N_10690,N_5769,N_7879);
nand U10691 (N_10691,N_4970,N_6972);
and U10692 (N_10692,N_6979,N_6639);
nor U10693 (N_10693,N_6895,N_6163);
or U10694 (N_10694,N_6621,N_4541);
nand U10695 (N_10695,N_5620,N_5869);
xor U10696 (N_10696,N_5958,N_6787);
and U10697 (N_10697,N_5734,N_6875);
and U10698 (N_10698,N_4168,N_5409);
and U10699 (N_10699,N_7898,N_4917);
nor U10700 (N_10700,N_4135,N_4916);
xnor U10701 (N_10701,N_5734,N_7974);
xor U10702 (N_10702,N_4103,N_6959);
or U10703 (N_10703,N_5957,N_6316);
nor U10704 (N_10704,N_5243,N_6615);
nand U10705 (N_10705,N_4380,N_7972);
or U10706 (N_10706,N_6831,N_5295);
xor U10707 (N_10707,N_4942,N_4805);
and U10708 (N_10708,N_4042,N_5745);
nand U10709 (N_10709,N_4229,N_4445);
nor U10710 (N_10710,N_5916,N_4599);
xnor U10711 (N_10711,N_7973,N_7707);
or U10712 (N_10712,N_5622,N_5648);
or U10713 (N_10713,N_7313,N_6997);
nor U10714 (N_10714,N_4073,N_4877);
xnor U10715 (N_10715,N_6229,N_6590);
nand U10716 (N_10716,N_6637,N_6687);
nor U10717 (N_10717,N_7684,N_5010);
and U10718 (N_10718,N_4151,N_5609);
nand U10719 (N_10719,N_5980,N_7154);
and U10720 (N_10720,N_7115,N_5609);
nor U10721 (N_10721,N_7549,N_6021);
and U10722 (N_10722,N_6471,N_7030);
nor U10723 (N_10723,N_4658,N_7055);
xnor U10724 (N_10724,N_5358,N_6285);
nor U10725 (N_10725,N_7544,N_7014);
or U10726 (N_10726,N_6040,N_5370);
nor U10727 (N_10727,N_4019,N_4869);
nor U10728 (N_10728,N_5858,N_4446);
nand U10729 (N_10729,N_5407,N_5937);
and U10730 (N_10730,N_4415,N_4481);
or U10731 (N_10731,N_4310,N_4367);
or U10732 (N_10732,N_4372,N_4542);
nor U10733 (N_10733,N_7426,N_5235);
nor U10734 (N_10734,N_5258,N_7058);
nand U10735 (N_10735,N_7785,N_7617);
nor U10736 (N_10736,N_7257,N_4809);
and U10737 (N_10737,N_6190,N_4250);
nor U10738 (N_10738,N_5267,N_6727);
nor U10739 (N_10739,N_7383,N_7049);
or U10740 (N_10740,N_4855,N_4254);
or U10741 (N_10741,N_7871,N_5180);
or U10742 (N_10742,N_4506,N_7211);
xor U10743 (N_10743,N_7685,N_6807);
nand U10744 (N_10744,N_4380,N_6764);
nand U10745 (N_10745,N_5523,N_7641);
nand U10746 (N_10746,N_7858,N_4685);
and U10747 (N_10747,N_5258,N_5840);
xor U10748 (N_10748,N_7623,N_5125);
and U10749 (N_10749,N_5241,N_7858);
xor U10750 (N_10750,N_5948,N_5683);
nor U10751 (N_10751,N_6543,N_6913);
or U10752 (N_10752,N_6839,N_6360);
and U10753 (N_10753,N_6846,N_6831);
nor U10754 (N_10754,N_4517,N_4659);
or U10755 (N_10755,N_5312,N_5817);
or U10756 (N_10756,N_6167,N_6378);
xnor U10757 (N_10757,N_7287,N_5897);
nand U10758 (N_10758,N_7560,N_4070);
or U10759 (N_10759,N_7468,N_7508);
xor U10760 (N_10760,N_6576,N_6461);
nand U10761 (N_10761,N_4346,N_4436);
and U10762 (N_10762,N_5069,N_6541);
nand U10763 (N_10763,N_7401,N_7093);
nor U10764 (N_10764,N_4090,N_5653);
nand U10765 (N_10765,N_6279,N_6460);
nor U10766 (N_10766,N_5587,N_6992);
nor U10767 (N_10767,N_5455,N_5205);
nand U10768 (N_10768,N_5991,N_4454);
nor U10769 (N_10769,N_4901,N_5098);
nand U10770 (N_10770,N_4933,N_5254);
xnor U10771 (N_10771,N_6381,N_6321);
xor U10772 (N_10772,N_6286,N_7624);
nor U10773 (N_10773,N_5802,N_5362);
or U10774 (N_10774,N_7782,N_4325);
and U10775 (N_10775,N_6548,N_5671);
xnor U10776 (N_10776,N_6869,N_5523);
nor U10777 (N_10777,N_7352,N_5328);
xor U10778 (N_10778,N_4679,N_4486);
nand U10779 (N_10779,N_7096,N_6700);
nand U10780 (N_10780,N_7712,N_5460);
and U10781 (N_10781,N_7743,N_5514);
nand U10782 (N_10782,N_7340,N_4419);
or U10783 (N_10783,N_6933,N_5912);
or U10784 (N_10784,N_6602,N_5423);
or U10785 (N_10785,N_7776,N_5777);
nor U10786 (N_10786,N_6215,N_7615);
nor U10787 (N_10787,N_4819,N_6993);
nand U10788 (N_10788,N_6638,N_4135);
xor U10789 (N_10789,N_7895,N_7707);
or U10790 (N_10790,N_4202,N_6697);
nor U10791 (N_10791,N_5373,N_4493);
and U10792 (N_10792,N_6779,N_4781);
nand U10793 (N_10793,N_4583,N_7968);
nor U10794 (N_10794,N_6182,N_4193);
and U10795 (N_10795,N_4459,N_4455);
nand U10796 (N_10796,N_7085,N_7550);
xnor U10797 (N_10797,N_4401,N_6162);
nand U10798 (N_10798,N_4994,N_6843);
or U10799 (N_10799,N_7780,N_5080);
and U10800 (N_10800,N_4829,N_6421);
nand U10801 (N_10801,N_6816,N_6472);
and U10802 (N_10802,N_6961,N_4253);
nor U10803 (N_10803,N_7523,N_4020);
nor U10804 (N_10804,N_4957,N_4038);
nor U10805 (N_10805,N_7895,N_4918);
or U10806 (N_10806,N_5121,N_5186);
or U10807 (N_10807,N_6364,N_7097);
nand U10808 (N_10808,N_5105,N_6599);
and U10809 (N_10809,N_4135,N_4102);
or U10810 (N_10810,N_5381,N_7454);
nand U10811 (N_10811,N_4662,N_6663);
or U10812 (N_10812,N_4785,N_6099);
nor U10813 (N_10813,N_5833,N_4695);
nor U10814 (N_10814,N_6682,N_6314);
or U10815 (N_10815,N_7792,N_4437);
and U10816 (N_10816,N_4288,N_7676);
and U10817 (N_10817,N_6158,N_7433);
or U10818 (N_10818,N_4915,N_6193);
nand U10819 (N_10819,N_7523,N_5103);
and U10820 (N_10820,N_7711,N_4581);
xnor U10821 (N_10821,N_6563,N_6434);
xnor U10822 (N_10822,N_6892,N_4671);
and U10823 (N_10823,N_4629,N_6204);
nand U10824 (N_10824,N_7892,N_6546);
or U10825 (N_10825,N_4968,N_6077);
nand U10826 (N_10826,N_6404,N_7086);
xor U10827 (N_10827,N_6851,N_4448);
nor U10828 (N_10828,N_4038,N_6225);
xor U10829 (N_10829,N_5846,N_5786);
nand U10830 (N_10830,N_5390,N_4918);
nand U10831 (N_10831,N_6711,N_5959);
and U10832 (N_10832,N_4303,N_7993);
and U10833 (N_10833,N_4224,N_4134);
xnor U10834 (N_10834,N_6657,N_7236);
or U10835 (N_10835,N_5113,N_4373);
or U10836 (N_10836,N_6366,N_7550);
nor U10837 (N_10837,N_4282,N_5020);
xor U10838 (N_10838,N_7762,N_5205);
and U10839 (N_10839,N_7185,N_6142);
nand U10840 (N_10840,N_7784,N_4294);
and U10841 (N_10841,N_6466,N_4417);
or U10842 (N_10842,N_5132,N_6071);
and U10843 (N_10843,N_6037,N_7475);
xnor U10844 (N_10844,N_7071,N_4074);
xor U10845 (N_10845,N_4537,N_6265);
or U10846 (N_10846,N_5502,N_5727);
nand U10847 (N_10847,N_4819,N_5492);
nand U10848 (N_10848,N_5451,N_7804);
or U10849 (N_10849,N_7752,N_5003);
or U10850 (N_10850,N_5236,N_7324);
nor U10851 (N_10851,N_5786,N_5109);
nor U10852 (N_10852,N_7534,N_7689);
or U10853 (N_10853,N_7251,N_6803);
nor U10854 (N_10854,N_7179,N_7033);
nand U10855 (N_10855,N_5160,N_6102);
nor U10856 (N_10856,N_5639,N_4301);
and U10857 (N_10857,N_7725,N_5105);
xor U10858 (N_10858,N_6763,N_6625);
xor U10859 (N_10859,N_5032,N_4277);
and U10860 (N_10860,N_4655,N_6486);
or U10861 (N_10861,N_5505,N_4106);
or U10862 (N_10862,N_7150,N_7617);
or U10863 (N_10863,N_5060,N_7604);
nand U10864 (N_10864,N_5714,N_6937);
or U10865 (N_10865,N_6766,N_4276);
xnor U10866 (N_10866,N_5260,N_6160);
or U10867 (N_10867,N_6158,N_4571);
nand U10868 (N_10868,N_5354,N_6652);
or U10869 (N_10869,N_5258,N_6495);
xor U10870 (N_10870,N_7044,N_4371);
xnor U10871 (N_10871,N_4195,N_7685);
nand U10872 (N_10872,N_6143,N_4527);
or U10873 (N_10873,N_4988,N_7698);
xnor U10874 (N_10874,N_7437,N_7526);
xor U10875 (N_10875,N_7279,N_6802);
nor U10876 (N_10876,N_6892,N_4968);
or U10877 (N_10877,N_6110,N_7154);
nor U10878 (N_10878,N_5566,N_7336);
and U10879 (N_10879,N_5426,N_4317);
or U10880 (N_10880,N_6222,N_7780);
nor U10881 (N_10881,N_7343,N_4666);
xor U10882 (N_10882,N_6820,N_7044);
and U10883 (N_10883,N_4032,N_5473);
nor U10884 (N_10884,N_6404,N_7875);
nand U10885 (N_10885,N_6387,N_6495);
xnor U10886 (N_10886,N_6301,N_7002);
xor U10887 (N_10887,N_4275,N_4679);
nor U10888 (N_10888,N_4915,N_4939);
xor U10889 (N_10889,N_6966,N_6673);
nor U10890 (N_10890,N_4115,N_7222);
or U10891 (N_10891,N_6318,N_4742);
or U10892 (N_10892,N_4500,N_4377);
nand U10893 (N_10893,N_5111,N_5859);
and U10894 (N_10894,N_6929,N_6710);
and U10895 (N_10895,N_5928,N_5213);
and U10896 (N_10896,N_6115,N_5153);
and U10897 (N_10897,N_4827,N_4630);
xor U10898 (N_10898,N_6485,N_6054);
nor U10899 (N_10899,N_7669,N_4982);
nand U10900 (N_10900,N_5623,N_7907);
xor U10901 (N_10901,N_5542,N_7618);
nand U10902 (N_10902,N_5656,N_7793);
xor U10903 (N_10903,N_4322,N_7891);
nand U10904 (N_10904,N_4250,N_5421);
or U10905 (N_10905,N_7156,N_5933);
xnor U10906 (N_10906,N_5895,N_5981);
or U10907 (N_10907,N_4209,N_5500);
xor U10908 (N_10908,N_7091,N_7765);
xnor U10909 (N_10909,N_7810,N_7618);
or U10910 (N_10910,N_5857,N_6225);
nand U10911 (N_10911,N_6168,N_4181);
xor U10912 (N_10912,N_4900,N_5915);
or U10913 (N_10913,N_7659,N_5244);
or U10914 (N_10914,N_5855,N_4310);
or U10915 (N_10915,N_5251,N_5028);
or U10916 (N_10916,N_7836,N_4767);
or U10917 (N_10917,N_5226,N_7042);
or U10918 (N_10918,N_7576,N_6445);
and U10919 (N_10919,N_6038,N_4611);
nor U10920 (N_10920,N_7767,N_4280);
nand U10921 (N_10921,N_6600,N_5817);
or U10922 (N_10922,N_4955,N_7156);
nand U10923 (N_10923,N_4353,N_4759);
nor U10924 (N_10924,N_5630,N_6763);
and U10925 (N_10925,N_7463,N_5882);
xor U10926 (N_10926,N_4259,N_4766);
or U10927 (N_10927,N_5997,N_7355);
nor U10928 (N_10928,N_4160,N_7057);
and U10929 (N_10929,N_6633,N_5070);
nor U10930 (N_10930,N_7777,N_7584);
nand U10931 (N_10931,N_5295,N_6840);
nand U10932 (N_10932,N_4632,N_7113);
nor U10933 (N_10933,N_7770,N_5844);
xor U10934 (N_10934,N_5798,N_7858);
nand U10935 (N_10935,N_6002,N_6291);
and U10936 (N_10936,N_6396,N_4260);
or U10937 (N_10937,N_4982,N_4100);
xnor U10938 (N_10938,N_7114,N_5565);
nand U10939 (N_10939,N_6314,N_7869);
or U10940 (N_10940,N_4380,N_5149);
nor U10941 (N_10941,N_7715,N_4568);
and U10942 (N_10942,N_4717,N_7079);
and U10943 (N_10943,N_5259,N_4688);
xnor U10944 (N_10944,N_4565,N_4162);
and U10945 (N_10945,N_7888,N_4538);
nor U10946 (N_10946,N_7182,N_5819);
nand U10947 (N_10947,N_5549,N_6660);
nor U10948 (N_10948,N_6120,N_7348);
and U10949 (N_10949,N_4691,N_5532);
nor U10950 (N_10950,N_6144,N_7487);
and U10951 (N_10951,N_5674,N_6715);
and U10952 (N_10952,N_7742,N_6228);
nand U10953 (N_10953,N_7440,N_5348);
nand U10954 (N_10954,N_5269,N_6953);
and U10955 (N_10955,N_6013,N_6933);
or U10956 (N_10956,N_5085,N_5975);
nand U10957 (N_10957,N_4802,N_4592);
and U10958 (N_10958,N_5512,N_5676);
nor U10959 (N_10959,N_4587,N_4537);
xor U10960 (N_10960,N_5905,N_6391);
or U10961 (N_10961,N_4386,N_5993);
and U10962 (N_10962,N_5725,N_4751);
xnor U10963 (N_10963,N_4147,N_7541);
or U10964 (N_10964,N_5858,N_7467);
or U10965 (N_10965,N_5431,N_7825);
or U10966 (N_10966,N_4735,N_4798);
nor U10967 (N_10967,N_7452,N_5534);
and U10968 (N_10968,N_4434,N_5852);
nand U10969 (N_10969,N_6390,N_6888);
nor U10970 (N_10970,N_7518,N_4678);
and U10971 (N_10971,N_7745,N_6267);
and U10972 (N_10972,N_6695,N_5610);
and U10973 (N_10973,N_5598,N_4422);
or U10974 (N_10974,N_7550,N_5519);
and U10975 (N_10975,N_7304,N_5748);
nand U10976 (N_10976,N_5847,N_7338);
or U10977 (N_10977,N_5374,N_4405);
or U10978 (N_10978,N_7961,N_5017);
nand U10979 (N_10979,N_6449,N_6179);
and U10980 (N_10980,N_7762,N_4559);
nor U10981 (N_10981,N_6067,N_5683);
nand U10982 (N_10982,N_6937,N_6049);
nor U10983 (N_10983,N_6310,N_5738);
and U10984 (N_10984,N_6966,N_5413);
or U10985 (N_10985,N_4969,N_6318);
or U10986 (N_10986,N_6056,N_4533);
xor U10987 (N_10987,N_6246,N_6510);
nand U10988 (N_10988,N_5703,N_4017);
nor U10989 (N_10989,N_5638,N_4961);
or U10990 (N_10990,N_5704,N_5147);
xnor U10991 (N_10991,N_6961,N_7752);
or U10992 (N_10992,N_7867,N_7398);
or U10993 (N_10993,N_7479,N_4653);
nor U10994 (N_10994,N_5998,N_6714);
or U10995 (N_10995,N_4280,N_6805);
nand U10996 (N_10996,N_7910,N_6507);
and U10997 (N_10997,N_4150,N_4107);
and U10998 (N_10998,N_7098,N_5927);
and U10999 (N_10999,N_6837,N_4223);
or U11000 (N_11000,N_6607,N_7371);
or U11001 (N_11001,N_5929,N_5065);
and U11002 (N_11002,N_5914,N_5555);
and U11003 (N_11003,N_4825,N_6384);
nor U11004 (N_11004,N_6163,N_4827);
xor U11005 (N_11005,N_4746,N_6011);
xor U11006 (N_11006,N_7344,N_4834);
and U11007 (N_11007,N_5065,N_5931);
or U11008 (N_11008,N_5796,N_4915);
and U11009 (N_11009,N_4471,N_5698);
nand U11010 (N_11010,N_4584,N_7120);
or U11011 (N_11011,N_6680,N_4787);
or U11012 (N_11012,N_5737,N_5265);
nor U11013 (N_11013,N_6648,N_7932);
and U11014 (N_11014,N_4222,N_7220);
or U11015 (N_11015,N_7766,N_5124);
nand U11016 (N_11016,N_6843,N_4020);
nand U11017 (N_11017,N_5342,N_6374);
nand U11018 (N_11018,N_7753,N_7043);
xor U11019 (N_11019,N_4102,N_6386);
or U11020 (N_11020,N_7649,N_4463);
or U11021 (N_11021,N_4949,N_6811);
and U11022 (N_11022,N_7263,N_4268);
and U11023 (N_11023,N_5835,N_5501);
and U11024 (N_11024,N_7475,N_4703);
or U11025 (N_11025,N_4716,N_6463);
or U11026 (N_11026,N_7968,N_5806);
or U11027 (N_11027,N_5813,N_6528);
xor U11028 (N_11028,N_7395,N_4058);
xnor U11029 (N_11029,N_6819,N_5182);
nor U11030 (N_11030,N_4367,N_6243);
and U11031 (N_11031,N_4951,N_5055);
nor U11032 (N_11032,N_7692,N_7613);
or U11033 (N_11033,N_7610,N_4894);
and U11034 (N_11034,N_5242,N_4356);
xor U11035 (N_11035,N_7261,N_4300);
or U11036 (N_11036,N_4359,N_5859);
nand U11037 (N_11037,N_7928,N_7062);
nand U11038 (N_11038,N_4611,N_4048);
xnor U11039 (N_11039,N_6211,N_5102);
and U11040 (N_11040,N_6660,N_7532);
nand U11041 (N_11041,N_7151,N_4636);
xor U11042 (N_11042,N_5690,N_7337);
and U11043 (N_11043,N_4239,N_5280);
xor U11044 (N_11044,N_7943,N_7247);
nand U11045 (N_11045,N_7066,N_6991);
and U11046 (N_11046,N_4308,N_7026);
nand U11047 (N_11047,N_5017,N_5061);
or U11048 (N_11048,N_5190,N_6737);
nand U11049 (N_11049,N_4832,N_4649);
nor U11050 (N_11050,N_6395,N_5543);
or U11051 (N_11051,N_6644,N_7126);
xnor U11052 (N_11052,N_7637,N_5838);
xor U11053 (N_11053,N_5745,N_6488);
xor U11054 (N_11054,N_5393,N_7967);
nor U11055 (N_11055,N_4904,N_6988);
nand U11056 (N_11056,N_5887,N_4173);
xnor U11057 (N_11057,N_5195,N_6188);
or U11058 (N_11058,N_7473,N_5640);
nand U11059 (N_11059,N_4082,N_6742);
or U11060 (N_11060,N_5766,N_4405);
nor U11061 (N_11061,N_7970,N_7478);
nand U11062 (N_11062,N_6720,N_6180);
and U11063 (N_11063,N_7222,N_7152);
nor U11064 (N_11064,N_6921,N_5132);
and U11065 (N_11065,N_7863,N_4978);
nand U11066 (N_11066,N_4001,N_7064);
and U11067 (N_11067,N_6472,N_6186);
nor U11068 (N_11068,N_4029,N_7449);
and U11069 (N_11069,N_5883,N_5416);
nor U11070 (N_11070,N_6203,N_4150);
and U11071 (N_11071,N_5839,N_7655);
nor U11072 (N_11072,N_4668,N_7341);
or U11073 (N_11073,N_7619,N_6837);
and U11074 (N_11074,N_6346,N_5336);
nand U11075 (N_11075,N_6607,N_4828);
or U11076 (N_11076,N_7838,N_5931);
and U11077 (N_11077,N_4454,N_5889);
or U11078 (N_11078,N_5873,N_7430);
xnor U11079 (N_11079,N_7997,N_4058);
nand U11080 (N_11080,N_6634,N_6361);
nand U11081 (N_11081,N_5251,N_7711);
or U11082 (N_11082,N_5466,N_4570);
xor U11083 (N_11083,N_5621,N_7532);
nor U11084 (N_11084,N_5249,N_5270);
and U11085 (N_11085,N_6334,N_5241);
nor U11086 (N_11086,N_6149,N_5868);
or U11087 (N_11087,N_5723,N_7843);
nand U11088 (N_11088,N_7469,N_5659);
nand U11089 (N_11089,N_6975,N_5841);
and U11090 (N_11090,N_6025,N_7198);
nor U11091 (N_11091,N_7162,N_4767);
nand U11092 (N_11092,N_5605,N_4373);
nand U11093 (N_11093,N_5764,N_7856);
nand U11094 (N_11094,N_6493,N_5345);
or U11095 (N_11095,N_6460,N_5453);
xnor U11096 (N_11096,N_4238,N_7835);
nand U11097 (N_11097,N_5863,N_7054);
nand U11098 (N_11098,N_4518,N_7421);
or U11099 (N_11099,N_7149,N_6297);
or U11100 (N_11100,N_7791,N_4689);
xor U11101 (N_11101,N_6971,N_5921);
xnor U11102 (N_11102,N_7458,N_5489);
and U11103 (N_11103,N_7882,N_5107);
nand U11104 (N_11104,N_4493,N_7834);
and U11105 (N_11105,N_6296,N_4767);
and U11106 (N_11106,N_4291,N_4652);
nor U11107 (N_11107,N_6277,N_5517);
or U11108 (N_11108,N_7003,N_7320);
nor U11109 (N_11109,N_4986,N_7143);
nand U11110 (N_11110,N_6499,N_4608);
and U11111 (N_11111,N_4764,N_6410);
nand U11112 (N_11112,N_4946,N_6281);
nor U11113 (N_11113,N_6577,N_5174);
and U11114 (N_11114,N_4165,N_5364);
nor U11115 (N_11115,N_5062,N_6468);
and U11116 (N_11116,N_4947,N_7946);
xnor U11117 (N_11117,N_6327,N_5079);
and U11118 (N_11118,N_5383,N_7690);
xor U11119 (N_11119,N_6077,N_7961);
nand U11120 (N_11120,N_5794,N_7063);
or U11121 (N_11121,N_5465,N_4021);
xnor U11122 (N_11122,N_6464,N_4997);
nand U11123 (N_11123,N_5885,N_7918);
nor U11124 (N_11124,N_6961,N_4178);
xor U11125 (N_11125,N_5390,N_7032);
xnor U11126 (N_11126,N_7505,N_5294);
nand U11127 (N_11127,N_4572,N_6630);
xor U11128 (N_11128,N_5354,N_6894);
and U11129 (N_11129,N_6536,N_5607);
xor U11130 (N_11130,N_7587,N_4521);
xnor U11131 (N_11131,N_5343,N_5431);
nor U11132 (N_11132,N_7104,N_6743);
and U11133 (N_11133,N_6482,N_5224);
xnor U11134 (N_11134,N_7502,N_6142);
or U11135 (N_11135,N_4833,N_5186);
nor U11136 (N_11136,N_4667,N_5849);
or U11137 (N_11137,N_7748,N_7326);
or U11138 (N_11138,N_4825,N_4035);
nand U11139 (N_11139,N_4764,N_6219);
xnor U11140 (N_11140,N_4657,N_6211);
or U11141 (N_11141,N_7192,N_5935);
and U11142 (N_11142,N_4341,N_5714);
nand U11143 (N_11143,N_5132,N_6052);
xor U11144 (N_11144,N_5267,N_5788);
nand U11145 (N_11145,N_6155,N_5835);
xor U11146 (N_11146,N_4750,N_6823);
xnor U11147 (N_11147,N_6084,N_4510);
xnor U11148 (N_11148,N_5010,N_6896);
and U11149 (N_11149,N_5060,N_7698);
xor U11150 (N_11150,N_6374,N_6017);
or U11151 (N_11151,N_4130,N_5545);
nand U11152 (N_11152,N_7268,N_6601);
or U11153 (N_11153,N_7985,N_4166);
nand U11154 (N_11154,N_6653,N_4443);
nor U11155 (N_11155,N_5265,N_4568);
xnor U11156 (N_11156,N_6007,N_5226);
and U11157 (N_11157,N_4629,N_5273);
and U11158 (N_11158,N_6463,N_4618);
nor U11159 (N_11159,N_4668,N_6613);
nand U11160 (N_11160,N_6332,N_7565);
or U11161 (N_11161,N_7187,N_5226);
nor U11162 (N_11162,N_4644,N_7471);
and U11163 (N_11163,N_5545,N_5443);
or U11164 (N_11164,N_7275,N_6037);
nand U11165 (N_11165,N_4134,N_5165);
and U11166 (N_11166,N_6439,N_5305);
nor U11167 (N_11167,N_6205,N_5610);
and U11168 (N_11168,N_5081,N_5448);
or U11169 (N_11169,N_5422,N_6129);
xnor U11170 (N_11170,N_6520,N_5138);
and U11171 (N_11171,N_6232,N_5917);
nor U11172 (N_11172,N_5202,N_4975);
and U11173 (N_11173,N_6982,N_7107);
or U11174 (N_11174,N_7901,N_5345);
xor U11175 (N_11175,N_5813,N_6732);
or U11176 (N_11176,N_6422,N_4343);
nor U11177 (N_11177,N_6888,N_6265);
nor U11178 (N_11178,N_4692,N_7531);
and U11179 (N_11179,N_7683,N_6641);
nand U11180 (N_11180,N_6463,N_5349);
nand U11181 (N_11181,N_7615,N_4673);
xnor U11182 (N_11182,N_7486,N_4572);
nand U11183 (N_11183,N_4059,N_5943);
nor U11184 (N_11184,N_6580,N_4035);
xor U11185 (N_11185,N_5852,N_4687);
nor U11186 (N_11186,N_4710,N_4437);
xnor U11187 (N_11187,N_4086,N_4078);
and U11188 (N_11188,N_4346,N_4076);
xor U11189 (N_11189,N_4494,N_6461);
nand U11190 (N_11190,N_5034,N_7198);
or U11191 (N_11191,N_5656,N_4376);
nor U11192 (N_11192,N_4322,N_7110);
nor U11193 (N_11193,N_7667,N_4537);
xnor U11194 (N_11194,N_6816,N_7881);
and U11195 (N_11195,N_4669,N_5856);
or U11196 (N_11196,N_4562,N_4439);
xnor U11197 (N_11197,N_6808,N_4273);
nand U11198 (N_11198,N_6307,N_5371);
xor U11199 (N_11199,N_6264,N_6467);
xor U11200 (N_11200,N_4067,N_5506);
or U11201 (N_11201,N_6742,N_4219);
nor U11202 (N_11202,N_7674,N_5643);
and U11203 (N_11203,N_7837,N_6124);
nor U11204 (N_11204,N_4809,N_6772);
and U11205 (N_11205,N_6353,N_6696);
or U11206 (N_11206,N_4616,N_6777);
or U11207 (N_11207,N_5500,N_6456);
nand U11208 (N_11208,N_7801,N_4197);
and U11209 (N_11209,N_4478,N_7889);
xor U11210 (N_11210,N_6697,N_4994);
or U11211 (N_11211,N_5908,N_6929);
and U11212 (N_11212,N_4323,N_7566);
or U11213 (N_11213,N_4830,N_7246);
or U11214 (N_11214,N_5932,N_5292);
nor U11215 (N_11215,N_7726,N_6139);
nand U11216 (N_11216,N_5490,N_6504);
and U11217 (N_11217,N_6491,N_4713);
nor U11218 (N_11218,N_6581,N_5660);
and U11219 (N_11219,N_6727,N_4659);
or U11220 (N_11220,N_6203,N_5513);
xnor U11221 (N_11221,N_6673,N_6680);
xor U11222 (N_11222,N_7486,N_6802);
or U11223 (N_11223,N_6235,N_4091);
nand U11224 (N_11224,N_7887,N_7576);
nor U11225 (N_11225,N_7238,N_6028);
and U11226 (N_11226,N_5429,N_7239);
and U11227 (N_11227,N_4096,N_4267);
and U11228 (N_11228,N_4212,N_5148);
nor U11229 (N_11229,N_6069,N_4369);
or U11230 (N_11230,N_4330,N_4747);
and U11231 (N_11231,N_6117,N_4058);
and U11232 (N_11232,N_6085,N_4698);
or U11233 (N_11233,N_5062,N_7493);
and U11234 (N_11234,N_7419,N_5847);
nor U11235 (N_11235,N_6869,N_7587);
nand U11236 (N_11236,N_7709,N_7935);
and U11237 (N_11237,N_4623,N_5239);
nor U11238 (N_11238,N_5733,N_7369);
nor U11239 (N_11239,N_5810,N_7985);
or U11240 (N_11240,N_7726,N_6191);
or U11241 (N_11241,N_7489,N_4215);
nand U11242 (N_11242,N_5472,N_4461);
nand U11243 (N_11243,N_5455,N_4020);
nor U11244 (N_11244,N_6612,N_6462);
xor U11245 (N_11245,N_4950,N_5365);
and U11246 (N_11246,N_7293,N_4105);
or U11247 (N_11247,N_7681,N_4993);
or U11248 (N_11248,N_7345,N_4080);
nor U11249 (N_11249,N_4712,N_5351);
nor U11250 (N_11250,N_7854,N_7476);
or U11251 (N_11251,N_4911,N_6618);
or U11252 (N_11252,N_7967,N_4539);
nand U11253 (N_11253,N_5354,N_7542);
or U11254 (N_11254,N_5634,N_5017);
xnor U11255 (N_11255,N_6024,N_5112);
or U11256 (N_11256,N_5425,N_7112);
nand U11257 (N_11257,N_4223,N_4739);
nand U11258 (N_11258,N_4425,N_6986);
xnor U11259 (N_11259,N_7165,N_7509);
and U11260 (N_11260,N_7477,N_6585);
nand U11261 (N_11261,N_5803,N_6600);
xnor U11262 (N_11262,N_7898,N_4324);
xor U11263 (N_11263,N_6489,N_7724);
and U11264 (N_11264,N_7501,N_6164);
and U11265 (N_11265,N_4752,N_5778);
nor U11266 (N_11266,N_6291,N_5619);
nand U11267 (N_11267,N_5854,N_7989);
and U11268 (N_11268,N_6166,N_4601);
xnor U11269 (N_11269,N_7240,N_7176);
xnor U11270 (N_11270,N_4034,N_7182);
xor U11271 (N_11271,N_7307,N_6145);
and U11272 (N_11272,N_4988,N_5677);
nor U11273 (N_11273,N_6736,N_4207);
xnor U11274 (N_11274,N_7018,N_5394);
or U11275 (N_11275,N_4691,N_4217);
and U11276 (N_11276,N_4333,N_6355);
xor U11277 (N_11277,N_4569,N_4683);
nor U11278 (N_11278,N_5164,N_5768);
and U11279 (N_11279,N_6194,N_4590);
and U11280 (N_11280,N_7013,N_7581);
nor U11281 (N_11281,N_4654,N_4147);
and U11282 (N_11282,N_4935,N_5522);
xor U11283 (N_11283,N_6360,N_7173);
nor U11284 (N_11284,N_4203,N_7946);
nor U11285 (N_11285,N_7818,N_6488);
or U11286 (N_11286,N_5962,N_6117);
nor U11287 (N_11287,N_7604,N_7026);
xor U11288 (N_11288,N_5454,N_6065);
nand U11289 (N_11289,N_4842,N_5508);
or U11290 (N_11290,N_5503,N_7417);
or U11291 (N_11291,N_7858,N_7864);
nand U11292 (N_11292,N_4056,N_4447);
nor U11293 (N_11293,N_5445,N_6502);
nor U11294 (N_11294,N_4012,N_5423);
nor U11295 (N_11295,N_4406,N_7144);
nor U11296 (N_11296,N_7706,N_6868);
xor U11297 (N_11297,N_4184,N_7773);
or U11298 (N_11298,N_7431,N_5468);
xor U11299 (N_11299,N_6657,N_7862);
nand U11300 (N_11300,N_7838,N_5147);
and U11301 (N_11301,N_6223,N_7960);
xnor U11302 (N_11302,N_7733,N_6413);
xor U11303 (N_11303,N_7704,N_7592);
nor U11304 (N_11304,N_6907,N_5484);
or U11305 (N_11305,N_5059,N_6881);
xor U11306 (N_11306,N_6325,N_5276);
nand U11307 (N_11307,N_7402,N_6198);
nand U11308 (N_11308,N_5850,N_6290);
or U11309 (N_11309,N_6066,N_7178);
and U11310 (N_11310,N_5891,N_6927);
and U11311 (N_11311,N_5367,N_6033);
nor U11312 (N_11312,N_5997,N_6021);
or U11313 (N_11313,N_4266,N_4904);
xor U11314 (N_11314,N_5932,N_6514);
or U11315 (N_11315,N_5230,N_6770);
nand U11316 (N_11316,N_4431,N_6383);
nor U11317 (N_11317,N_5333,N_7327);
or U11318 (N_11318,N_5146,N_6564);
and U11319 (N_11319,N_5328,N_4693);
xnor U11320 (N_11320,N_4280,N_6972);
nand U11321 (N_11321,N_7886,N_4266);
nor U11322 (N_11322,N_7463,N_4215);
nor U11323 (N_11323,N_7332,N_5903);
and U11324 (N_11324,N_4567,N_4558);
nand U11325 (N_11325,N_5377,N_6203);
and U11326 (N_11326,N_7937,N_4787);
and U11327 (N_11327,N_6227,N_7880);
or U11328 (N_11328,N_4825,N_6115);
or U11329 (N_11329,N_6824,N_6098);
or U11330 (N_11330,N_7437,N_5617);
nand U11331 (N_11331,N_6463,N_6359);
or U11332 (N_11332,N_5792,N_6402);
nand U11333 (N_11333,N_7048,N_5422);
and U11334 (N_11334,N_5844,N_7841);
xnor U11335 (N_11335,N_5902,N_7533);
or U11336 (N_11336,N_7026,N_4859);
and U11337 (N_11337,N_5016,N_7533);
or U11338 (N_11338,N_4986,N_5354);
nor U11339 (N_11339,N_5859,N_4582);
or U11340 (N_11340,N_6292,N_7483);
or U11341 (N_11341,N_5977,N_5732);
nand U11342 (N_11342,N_4902,N_5225);
nor U11343 (N_11343,N_5900,N_5914);
nand U11344 (N_11344,N_6343,N_6165);
nor U11345 (N_11345,N_4105,N_4052);
xnor U11346 (N_11346,N_5391,N_5280);
xnor U11347 (N_11347,N_5547,N_5555);
nor U11348 (N_11348,N_6341,N_5019);
or U11349 (N_11349,N_7358,N_4091);
and U11350 (N_11350,N_6484,N_6392);
nor U11351 (N_11351,N_7747,N_4324);
and U11352 (N_11352,N_7808,N_6793);
or U11353 (N_11353,N_7459,N_7099);
nor U11354 (N_11354,N_7189,N_5964);
and U11355 (N_11355,N_4128,N_7932);
and U11356 (N_11356,N_7385,N_6475);
xor U11357 (N_11357,N_4692,N_6974);
nor U11358 (N_11358,N_4718,N_5766);
nor U11359 (N_11359,N_4106,N_5290);
xnor U11360 (N_11360,N_7429,N_4739);
nand U11361 (N_11361,N_7842,N_4899);
nor U11362 (N_11362,N_5931,N_5295);
nor U11363 (N_11363,N_4783,N_7554);
nor U11364 (N_11364,N_5432,N_7048);
nand U11365 (N_11365,N_4498,N_4365);
nor U11366 (N_11366,N_4822,N_7354);
nand U11367 (N_11367,N_6669,N_6328);
nor U11368 (N_11368,N_7411,N_7471);
and U11369 (N_11369,N_5235,N_5016);
nand U11370 (N_11370,N_5348,N_6244);
xnor U11371 (N_11371,N_5148,N_5257);
nand U11372 (N_11372,N_5112,N_5776);
and U11373 (N_11373,N_6644,N_7746);
nand U11374 (N_11374,N_6762,N_4880);
or U11375 (N_11375,N_6382,N_4681);
nor U11376 (N_11376,N_4206,N_6663);
or U11377 (N_11377,N_5077,N_4059);
xor U11378 (N_11378,N_7645,N_6007);
and U11379 (N_11379,N_6709,N_6531);
and U11380 (N_11380,N_5539,N_6324);
or U11381 (N_11381,N_4198,N_7934);
xnor U11382 (N_11382,N_6681,N_6243);
or U11383 (N_11383,N_7412,N_5757);
xnor U11384 (N_11384,N_7040,N_6450);
nand U11385 (N_11385,N_7160,N_5798);
and U11386 (N_11386,N_6619,N_6810);
or U11387 (N_11387,N_7669,N_6175);
and U11388 (N_11388,N_6788,N_5585);
xnor U11389 (N_11389,N_5390,N_7373);
or U11390 (N_11390,N_6334,N_4340);
and U11391 (N_11391,N_7765,N_7600);
nor U11392 (N_11392,N_6512,N_6160);
nor U11393 (N_11393,N_7438,N_5986);
xnor U11394 (N_11394,N_4739,N_4166);
xnor U11395 (N_11395,N_4847,N_4516);
or U11396 (N_11396,N_7499,N_4787);
xnor U11397 (N_11397,N_6486,N_7566);
and U11398 (N_11398,N_4021,N_7797);
xnor U11399 (N_11399,N_4786,N_4113);
nor U11400 (N_11400,N_4875,N_5382);
xor U11401 (N_11401,N_7579,N_7111);
nor U11402 (N_11402,N_7073,N_7772);
and U11403 (N_11403,N_4565,N_5128);
nand U11404 (N_11404,N_7478,N_6774);
and U11405 (N_11405,N_5773,N_6005);
xnor U11406 (N_11406,N_7272,N_7883);
xnor U11407 (N_11407,N_6909,N_5844);
nand U11408 (N_11408,N_7756,N_6760);
nand U11409 (N_11409,N_7558,N_4222);
or U11410 (N_11410,N_6333,N_7818);
nor U11411 (N_11411,N_4785,N_5200);
nor U11412 (N_11412,N_6008,N_5145);
or U11413 (N_11413,N_4636,N_5305);
or U11414 (N_11414,N_7577,N_6566);
and U11415 (N_11415,N_7545,N_5737);
nor U11416 (N_11416,N_5702,N_5058);
xnor U11417 (N_11417,N_7388,N_6128);
xor U11418 (N_11418,N_4862,N_7969);
xnor U11419 (N_11419,N_4415,N_7874);
xor U11420 (N_11420,N_7321,N_5830);
nand U11421 (N_11421,N_6039,N_5363);
or U11422 (N_11422,N_7749,N_7935);
nor U11423 (N_11423,N_7940,N_5182);
nor U11424 (N_11424,N_7289,N_4671);
xor U11425 (N_11425,N_5628,N_5183);
or U11426 (N_11426,N_4512,N_5369);
nand U11427 (N_11427,N_7840,N_7772);
nor U11428 (N_11428,N_7160,N_7464);
or U11429 (N_11429,N_5189,N_4720);
nor U11430 (N_11430,N_7384,N_5168);
nor U11431 (N_11431,N_7264,N_7420);
nor U11432 (N_11432,N_5618,N_4739);
and U11433 (N_11433,N_7737,N_4796);
xor U11434 (N_11434,N_4049,N_5987);
nand U11435 (N_11435,N_5478,N_5860);
nand U11436 (N_11436,N_4701,N_4322);
xnor U11437 (N_11437,N_5993,N_4803);
and U11438 (N_11438,N_5280,N_4554);
and U11439 (N_11439,N_4863,N_6448);
or U11440 (N_11440,N_5095,N_6492);
and U11441 (N_11441,N_7875,N_6378);
and U11442 (N_11442,N_6227,N_7405);
nand U11443 (N_11443,N_6346,N_6392);
and U11444 (N_11444,N_4323,N_5095);
nor U11445 (N_11445,N_4020,N_6606);
nand U11446 (N_11446,N_5492,N_7828);
xor U11447 (N_11447,N_7529,N_7308);
or U11448 (N_11448,N_6669,N_5640);
or U11449 (N_11449,N_4535,N_4556);
nor U11450 (N_11450,N_6951,N_4650);
nor U11451 (N_11451,N_4229,N_6105);
xnor U11452 (N_11452,N_5235,N_6824);
or U11453 (N_11453,N_4317,N_7217);
nand U11454 (N_11454,N_6601,N_7981);
nand U11455 (N_11455,N_6720,N_7339);
and U11456 (N_11456,N_5277,N_5336);
nand U11457 (N_11457,N_5929,N_5726);
or U11458 (N_11458,N_7014,N_5083);
nand U11459 (N_11459,N_7149,N_7117);
xnor U11460 (N_11460,N_7736,N_4545);
nor U11461 (N_11461,N_5507,N_6958);
xor U11462 (N_11462,N_5825,N_7889);
or U11463 (N_11463,N_6695,N_6526);
nand U11464 (N_11464,N_5232,N_6750);
nor U11465 (N_11465,N_7051,N_5787);
nand U11466 (N_11466,N_4165,N_6659);
nand U11467 (N_11467,N_6540,N_6054);
nand U11468 (N_11468,N_4342,N_4491);
nor U11469 (N_11469,N_7536,N_7025);
xor U11470 (N_11470,N_5675,N_4201);
nor U11471 (N_11471,N_6727,N_4889);
and U11472 (N_11472,N_6428,N_7226);
and U11473 (N_11473,N_4425,N_7657);
nand U11474 (N_11474,N_7444,N_5638);
nand U11475 (N_11475,N_6938,N_4370);
nand U11476 (N_11476,N_6743,N_7092);
xor U11477 (N_11477,N_7163,N_4558);
or U11478 (N_11478,N_5707,N_7610);
and U11479 (N_11479,N_6138,N_4794);
nor U11480 (N_11480,N_5306,N_7150);
nor U11481 (N_11481,N_5663,N_5144);
or U11482 (N_11482,N_6413,N_7594);
nand U11483 (N_11483,N_5813,N_7057);
nor U11484 (N_11484,N_5385,N_5652);
or U11485 (N_11485,N_6712,N_7029);
nand U11486 (N_11486,N_5888,N_6203);
and U11487 (N_11487,N_5296,N_6941);
and U11488 (N_11488,N_4830,N_5961);
and U11489 (N_11489,N_5541,N_5772);
nor U11490 (N_11490,N_4279,N_7472);
and U11491 (N_11491,N_7962,N_6111);
or U11492 (N_11492,N_6737,N_4958);
nand U11493 (N_11493,N_4557,N_4419);
nand U11494 (N_11494,N_5793,N_5117);
and U11495 (N_11495,N_6934,N_7984);
or U11496 (N_11496,N_6772,N_5878);
xor U11497 (N_11497,N_5495,N_7649);
nor U11498 (N_11498,N_4070,N_7536);
nand U11499 (N_11499,N_4193,N_7516);
and U11500 (N_11500,N_5594,N_4084);
and U11501 (N_11501,N_6508,N_4214);
nand U11502 (N_11502,N_5219,N_5083);
xnor U11503 (N_11503,N_4889,N_5037);
xnor U11504 (N_11504,N_6801,N_4474);
and U11505 (N_11505,N_6894,N_7092);
nand U11506 (N_11506,N_4863,N_7714);
or U11507 (N_11507,N_4478,N_7812);
and U11508 (N_11508,N_7955,N_7357);
nand U11509 (N_11509,N_5018,N_7466);
nor U11510 (N_11510,N_6950,N_5206);
and U11511 (N_11511,N_5099,N_7132);
xnor U11512 (N_11512,N_5380,N_7676);
xnor U11513 (N_11513,N_5482,N_6376);
and U11514 (N_11514,N_5129,N_5182);
nand U11515 (N_11515,N_5704,N_4633);
or U11516 (N_11516,N_6988,N_7162);
or U11517 (N_11517,N_5872,N_6928);
or U11518 (N_11518,N_5612,N_4242);
and U11519 (N_11519,N_4170,N_5739);
and U11520 (N_11520,N_5986,N_7230);
nand U11521 (N_11521,N_4990,N_4463);
and U11522 (N_11522,N_5496,N_6722);
nor U11523 (N_11523,N_4886,N_5870);
xor U11524 (N_11524,N_5440,N_4548);
nand U11525 (N_11525,N_5706,N_7672);
xor U11526 (N_11526,N_5400,N_4685);
nor U11527 (N_11527,N_7600,N_6521);
xnor U11528 (N_11528,N_4977,N_6543);
nand U11529 (N_11529,N_6341,N_6380);
or U11530 (N_11530,N_7269,N_7000);
xnor U11531 (N_11531,N_4081,N_5204);
xor U11532 (N_11532,N_7107,N_4591);
nor U11533 (N_11533,N_6832,N_4413);
nand U11534 (N_11534,N_7433,N_4791);
or U11535 (N_11535,N_7172,N_5721);
and U11536 (N_11536,N_5958,N_4556);
nand U11537 (N_11537,N_4241,N_5098);
or U11538 (N_11538,N_5670,N_4454);
nand U11539 (N_11539,N_7043,N_4220);
or U11540 (N_11540,N_7466,N_7882);
xnor U11541 (N_11541,N_7436,N_5156);
xor U11542 (N_11542,N_4216,N_5186);
and U11543 (N_11543,N_5446,N_7568);
nor U11544 (N_11544,N_7303,N_5535);
and U11545 (N_11545,N_5207,N_7900);
and U11546 (N_11546,N_5296,N_5870);
or U11547 (N_11547,N_4935,N_4404);
nand U11548 (N_11548,N_5918,N_6378);
nand U11549 (N_11549,N_5317,N_4128);
and U11550 (N_11550,N_5556,N_5433);
and U11551 (N_11551,N_4185,N_7831);
nor U11552 (N_11552,N_5342,N_7630);
nand U11553 (N_11553,N_5686,N_5048);
and U11554 (N_11554,N_5999,N_7564);
nor U11555 (N_11555,N_5072,N_6915);
or U11556 (N_11556,N_7068,N_5883);
and U11557 (N_11557,N_4190,N_6985);
nor U11558 (N_11558,N_5059,N_6201);
and U11559 (N_11559,N_6941,N_7354);
nor U11560 (N_11560,N_7502,N_6069);
xor U11561 (N_11561,N_7181,N_5761);
or U11562 (N_11562,N_5876,N_4622);
nor U11563 (N_11563,N_4450,N_7049);
nor U11564 (N_11564,N_5172,N_4518);
nor U11565 (N_11565,N_5728,N_5625);
and U11566 (N_11566,N_5200,N_4048);
nor U11567 (N_11567,N_6057,N_5603);
nand U11568 (N_11568,N_6926,N_5860);
or U11569 (N_11569,N_6648,N_5493);
nor U11570 (N_11570,N_5655,N_5803);
nand U11571 (N_11571,N_6029,N_6880);
nor U11572 (N_11572,N_4600,N_7432);
nand U11573 (N_11573,N_4173,N_4484);
xnor U11574 (N_11574,N_5884,N_5374);
xor U11575 (N_11575,N_5681,N_4836);
nor U11576 (N_11576,N_5109,N_4657);
nor U11577 (N_11577,N_6915,N_7597);
and U11578 (N_11578,N_5802,N_7896);
nor U11579 (N_11579,N_4778,N_6232);
xnor U11580 (N_11580,N_6800,N_7046);
and U11581 (N_11581,N_4855,N_6822);
nor U11582 (N_11582,N_5486,N_5308);
or U11583 (N_11583,N_4304,N_7268);
xnor U11584 (N_11584,N_4778,N_5656);
nand U11585 (N_11585,N_5297,N_6939);
or U11586 (N_11586,N_4390,N_6476);
nor U11587 (N_11587,N_5090,N_4137);
xnor U11588 (N_11588,N_5693,N_5100);
nand U11589 (N_11589,N_5073,N_4954);
nand U11590 (N_11590,N_7120,N_5516);
nor U11591 (N_11591,N_5319,N_6467);
or U11592 (N_11592,N_4946,N_5486);
nor U11593 (N_11593,N_5490,N_5571);
or U11594 (N_11594,N_5577,N_5721);
nand U11595 (N_11595,N_7125,N_6441);
nand U11596 (N_11596,N_6442,N_6509);
nor U11597 (N_11597,N_4749,N_4211);
xor U11598 (N_11598,N_7854,N_4736);
or U11599 (N_11599,N_4934,N_7156);
nand U11600 (N_11600,N_5365,N_6279);
and U11601 (N_11601,N_6894,N_4255);
and U11602 (N_11602,N_5455,N_4719);
nor U11603 (N_11603,N_6146,N_6821);
or U11604 (N_11604,N_6386,N_4471);
nor U11605 (N_11605,N_4773,N_6159);
nor U11606 (N_11606,N_6228,N_7025);
xnor U11607 (N_11607,N_5507,N_5992);
xnor U11608 (N_11608,N_5906,N_7760);
nand U11609 (N_11609,N_7810,N_6397);
xnor U11610 (N_11610,N_4733,N_7292);
nand U11611 (N_11611,N_7849,N_4160);
or U11612 (N_11612,N_4827,N_5052);
nor U11613 (N_11613,N_4809,N_6581);
xnor U11614 (N_11614,N_6725,N_4614);
nor U11615 (N_11615,N_6475,N_7237);
nand U11616 (N_11616,N_4085,N_6073);
nand U11617 (N_11617,N_6392,N_5321);
nor U11618 (N_11618,N_6360,N_7518);
xor U11619 (N_11619,N_4289,N_5678);
nor U11620 (N_11620,N_4054,N_6860);
or U11621 (N_11621,N_4746,N_5386);
nor U11622 (N_11622,N_7211,N_7881);
xnor U11623 (N_11623,N_7210,N_5373);
xnor U11624 (N_11624,N_6022,N_4658);
nor U11625 (N_11625,N_7100,N_6422);
and U11626 (N_11626,N_7564,N_7997);
nand U11627 (N_11627,N_5278,N_5701);
or U11628 (N_11628,N_7204,N_6467);
and U11629 (N_11629,N_6632,N_4639);
xnor U11630 (N_11630,N_6572,N_4670);
nand U11631 (N_11631,N_7659,N_5098);
and U11632 (N_11632,N_5366,N_4444);
nor U11633 (N_11633,N_6256,N_6747);
xor U11634 (N_11634,N_6571,N_7526);
nand U11635 (N_11635,N_4671,N_7986);
nor U11636 (N_11636,N_6889,N_5832);
xnor U11637 (N_11637,N_4313,N_7366);
nand U11638 (N_11638,N_4724,N_7650);
nand U11639 (N_11639,N_5781,N_6855);
nor U11640 (N_11640,N_5300,N_5083);
nand U11641 (N_11641,N_4631,N_6534);
xor U11642 (N_11642,N_6087,N_6947);
nor U11643 (N_11643,N_7730,N_4855);
xor U11644 (N_11644,N_7175,N_5874);
or U11645 (N_11645,N_7234,N_4131);
and U11646 (N_11646,N_6805,N_7951);
xnor U11647 (N_11647,N_4259,N_6998);
or U11648 (N_11648,N_4540,N_5899);
or U11649 (N_11649,N_4525,N_4352);
nand U11650 (N_11650,N_4511,N_7372);
or U11651 (N_11651,N_4574,N_4705);
xor U11652 (N_11652,N_7389,N_6358);
and U11653 (N_11653,N_6763,N_4361);
and U11654 (N_11654,N_6662,N_7865);
nor U11655 (N_11655,N_6175,N_7554);
and U11656 (N_11656,N_4852,N_7673);
nor U11657 (N_11657,N_4537,N_7461);
xor U11658 (N_11658,N_5535,N_6878);
or U11659 (N_11659,N_7551,N_6916);
or U11660 (N_11660,N_6983,N_4180);
xnor U11661 (N_11661,N_4936,N_7742);
or U11662 (N_11662,N_6046,N_7273);
nand U11663 (N_11663,N_7441,N_5043);
or U11664 (N_11664,N_4073,N_7738);
and U11665 (N_11665,N_7400,N_7519);
nor U11666 (N_11666,N_6519,N_4999);
or U11667 (N_11667,N_6987,N_6268);
xor U11668 (N_11668,N_4118,N_6597);
nand U11669 (N_11669,N_4772,N_6008);
xnor U11670 (N_11670,N_7696,N_6478);
nand U11671 (N_11671,N_5402,N_7479);
nand U11672 (N_11672,N_6778,N_6388);
xor U11673 (N_11673,N_6552,N_4471);
nor U11674 (N_11674,N_6334,N_5496);
nor U11675 (N_11675,N_6431,N_6328);
nor U11676 (N_11676,N_4298,N_4464);
nor U11677 (N_11677,N_6936,N_7547);
and U11678 (N_11678,N_5519,N_6883);
and U11679 (N_11679,N_7349,N_5126);
and U11680 (N_11680,N_6472,N_6660);
nand U11681 (N_11681,N_5122,N_7067);
and U11682 (N_11682,N_6305,N_7806);
or U11683 (N_11683,N_4080,N_5839);
and U11684 (N_11684,N_5075,N_5779);
or U11685 (N_11685,N_4731,N_6548);
or U11686 (N_11686,N_4252,N_5335);
or U11687 (N_11687,N_5415,N_5258);
and U11688 (N_11688,N_5692,N_7364);
nor U11689 (N_11689,N_5738,N_5401);
or U11690 (N_11690,N_5828,N_5735);
nand U11691 (N_11691,N_7590,N_5671);
nand U11692 (N_11692,N_4369,N_6938);
xnor U11693 (N_11693,N_4319,N_6930);
nand U11694 (N_11694,N_5527,N_6637);
and U11695 (N_11695,N_6870,N_4742);
xnor U11696 (N_11696,N_6988,N_5327);
nor U11697 (N_11697,N_5653,N_7515);
xnor U11698 (N_11698,N_6453,N_7335);
and U11699 (N_11699,N_6480,N_7980);
xor U11700 (N_11700,N_7194,N_7964);
nor U11701 (N_11701,N_4076,N_4510);
nor U11702 (N_11702,N_6517,N_4699);
nor U11703 (N_11703,N_7205,N_5527);
nand U11704 (N_11704,N_6712,N_4645);
and U11705 (N_11705,N_7004,N_6505);
and U11706 (N_11706,N_5617,N_6578);
nand U11707 (N_11707,N_7990,N_6853);
nand U11708 (N_11708,N_7325,N_6597);
and U11709 (N_11709,N_7282,N_5370);
xor U11710 (N_11710,N_7117,N_7942);
or U11711 (N_11711,N_7553,N_7249);
and U11712 (N_11712,N_4598,N_4229);
xnor U11713 (N_11713,N_5005,N_7651);
and U11714 (N_11714,N_4047,N_7281);
nand U11715 (N_11715,N_5096,N_6175);
or U11716 (N_11716,N_6862,N_5361);
or U11717 (N_11717,N_6483,N_6572);
and U11718 (N_11718,N_4607,N_6750);
and U11719 (N_11719,N_7782,N_4464);
xor U11720 (N_11720,N_7051,N_5304);
xnor U11721 (N_11721,N_4207,N_7145);
nor U11722 (N_11722,N_5677,N_4151);
and U11723 (N_11723,N_5919,N_5032);
nor U11724 (N_11724,N_5333,N_5797);
xnor U11725 (N_11725,N_4601,N_7667);
nand U11726 (N_11726,N_4239,N_6162);
xnor U11727 (N_11727,N_7750,N_6670);
nor U11728 (N_11728,N_5939,N_4292);
xnor U11729 (N_11729,N_4770,N_5053);
nor U11730 (N_11730,N_7656,N_5211);
nor U11731 (N_11731,N_5013,N_7938);
and U11732 (N_11732,N_7640,N_6336);
nor U11733 (N_11733,N_7032,N_5331);
nand U11734 (N_11734,N_4428,N_6026);
and U11735 (N_11735,N_4455,N_4515);
nand U11736 (N_11736,N_5931,N_4300);
xor U11737 (N_11737,N_7473,N_4376);
nor U11738 (N_11738,N_6296,N_5413);
nor U11739 (N_11739,N_4221,N_6925);
or U11740 (N_11740,N_6956,N_6600);
or U11741 (N_11741,N_7078,N_4512);
nand U11742 (N_11742,N_5066,N_5867);
and U11743 (N_11743,N_5147,N_5656);
or U11744 (N_11744,N_7230,N_7926);
xor U11745 (N_11745,N_7146,N_7860);
or U11746 (N_11746,N_7790,N_5096);
and U11747 (N_11747,N_5774,N_4530);
or U11748 (N_11748,N_7028,N_6719);
xnor U11749 (N_11749,N_4824,N_5772);
nand U11750 (N_11750,N_5530,N_5386);
xnor U11751 (N_11751,N_5520,N_4235);
xnor U11752 (N_11752,N_7222,N_6746);
xor U11753 (N_11753,N_7074,N_7534);
xor U11754 (N_11754,N_4146,N_6246);
nor U11755 (N_11755,N_6421,N_6796);
nor U11756 (N_11756,N_4992,N_4980);
and U11757 (N_11757,N_6439,N_7826);
or U11758 (N_11758,N_5787,N_7765);
xor U11759 (N_11759,N_6141,N_7077);
xnor U11760 (N_11760,N_4384,N_6878);
or U11761 (N_11761,N_4685,N_5176);
xor U11762 (N_11762,N_4805,N_5749);
xnor U11763 (N_11763,N_5571,N_6856);
and U11764 (N_11764,N_6512,N_4515);
xor U11765 (N_11765,N_4355,N_4735);
and U11766 (N_11766,N_4023,N_7045);
and U11767 (N_11767,N_4934,N_4758);
nand U11768 (N_11768,N_5609,N_7833);
xnor U11769 (N_11769,N_5912,N_4344);
xor U11770 (N_11770,N_5323,N_4726);
and U11771 (N_11771,N_5204,N_7744);
nor U11772 (N_11772,N_5313,N_4833);
or U11773 (N_11773,N_4138,N_5617);
xor U11774 (N_11774,N_6799,N_4312);
or U11775 (N_11775,N_6196,N_6474);
nor U11776 (N_11776,N_4535,N_7495);
nand U11777 (N_11777,N_4698,N_7485);
or U11778 (N_11778,N_5822,N_5016);
or U11779 (N_11779,N_5208,N_5843);
and U11780 (N_11780,N_6895,N_6585);
nor U11781 (N_11781,N_7368,N_6676);
or U11782 (N_11782,N_4776,N_7844);
xor U11783 (N_11783,N_4570,N_4905);
nand U11784 (N_11784,N_7202,N_4395);
and U11785 (N_11785,N_5765,N_6712);
nand U11786 (N_11786,N_6914,N_5467);
or U11787 (N_11787,N_4616,N_5770);
nand U11788 (N_11788,N_5981,N_5885);
and U11789 (N_11789,N_7529,N_6567);
and U11790 (N_11790,N_5233,N_5968);
nand U11791 (N_11791,N_4270,N_5309);
and U11792 (N_11792,N_6483,N_5233);
nand U11793 (N_11793,N_5384,N_4735);
xnor U11794 (N_11794,N_5247,N_5220);
nand U11795 (N_11795,N_6825,N_5390);
nand U11796 (N_11796,N_5839,N_6253);
or U11797 (N_11797,N_5951,N_6693);
xnor U11798 (N_11798,N_4520,N_4726);
and U11799 (N_11799,N_4909,N_5164);
or U11800 (N_11800,N_4728,N_5366);
or U11801 (N_11801,N_6826,N_7938);
nor U11802 (N_11802,N_7408,N_6315);
or U11803 (N_11803,N_4687,N_4751);
or U11804 (N_11804,N_4273,N_6294);
nand U11805 (N_11805,N_7903,N_4076);
and U11806 (N_11806,N_7406,N_5100);
and U11807 (N_11807,N_7740,N_4431);
xnor U11808 (N_11808,N_7076,N_7820);
nand U11809 (N_11809,N_7675,N_5872);
nand U11810 (N_11810,N_6559,N_4462);
nand U11811 (N_11811,N_5152,N_6618);
nand U11812 (N_11812,N_4701,N_7041);
and U11813 (N_11813,N_6734,N_4667);
nor U11814 (N_11814,N_7247,N_7298);
nor U11815 (N_11815,N_5766,N_6726);
xnor U11816 (N_11816,N_5638,N_7824);
nand U11817 (N_11817,N_7245,N_5129);
or U11818 (N_11818,N_5468,N_7909);
nor U11819 (N_11819,N_6901,N_6113);
nor U11820 (N_11820,N_6942,N_6833);
or U11821 (N_11821,N_7910,N_6562);
and U11822 (N_11822,N_7116,N_4202);
nand U11823 (N_11823,N_7909,N_4131);
and U11824 (N_11824,N_4373,N_7021);
nand U11825 (N_11825,N_6185,N_6194);
and U11826 (N_11826,N_7943,N_7043);
or U11827 (N_11827,N_5309,N_6568);
nand U11828 (N_11828,N_7097,N_7316);
nor U11829 (N_11829,N_7915,N_6853);
xor U11830 (N_11830,N_5343,N_4404);
nand U11831 (N_11831,N_7430,N_7247);
and U11832 (N_11832,N_7667,N_7580);
nand U11833 (N_11833,N_7333,N_6412);
nor U11834 (N_11834,N_4031,N_5915);
or U11835 (N_11835,N_6582,N_5236);
nand U11836 (N_11836,N_7088,N_7922);
xnor U11837 (N_11837,N_6324,N_5398);
xnor U11838 (N_11838,N_7949,N_4334);
and U11839 (N_11839,N_7746,N_4827);
nor U11840 (N_11840,N_4087,N_4667);
nor U11841 (N_11841,N_7374,N_7042);
or U11842 (N_11842,N_4661,N_7572);
nor U11843 (N_11843,N_5556,N_7122);
xor U11844 (N_11844,N_6976,N_5126);
and U11845 (N_11845,N_5192,N_5594);
nor U11846 (N_11846,N_6246,N_4593);
nor U11847 (N_11847,N_6750,N_7247);
xnor U11848 (N_11848,N_5563,N_7770);
nor U11849 (N_11849,N_4120,N_4826);
nand U11850 (N_11850,N_5435,N_6346);
xnor U11851 (N_11851,N_6450,N_4227);
and U11852 (N_11852,N_7283,N_5237);
xor U11853 (N_11853,N_4936,N_7769);
xnor U11854 (N_11854,N_7602,N_7834);
xnor U11855 (N_11855,N_5620,N_6907);
xor U11856 (N_11856,N_7292,N_5028);
and U11857 (N_11857,N_5555,N_5539);
xor U11858 (N_11858,N_7032,N_5443);
nor U11859 (N_11859,N_6522,N_6541);
nor U11860 (N_11860,N_6986,N_6602);
and U11861 (N_11861,N_5784,N_6768);
xor U11862 (N_11862,N_4434,N_4276);
xnor U11863 (N_11863,N_6487,N_4069);
xnor U11864 (N_11864,N_4790,N_5621);
nor U11865 (N_11865,N_4452,N_7464);
nor U11866 (N_11866,N_4010,N_4365);
xnor U11867 (N_11867,N_7995,N_4116);
nand U11868 (N_11868,N_5260,N_7094);
nand U11869 (N_11869,N_6068,N_5125);
xor U11870 (N_11870,N_6846,N_7308);
nand U11871 (N_11871,N_5863,N_4089);
and U11872 (N_11872,N_7166,N_4142);
nand U11873 (N_11873,N_5531,N_7237);
nand U11874 (N_11874,N_4156,N_4323);
nand U11875 (N_11875,N_5357,N_6719);
xor U11876 (N_11876,N_4179,N_6826);
and U11877 (N_11877,N_5574,N_5309);
xnor U11878 (N_11878,N_4776,N_6337);
nor U11879 (N_11879,N_7390,N_7406);
nor U11880 (N_11880,N_4064,N_5956);
nand U11881 (N_11881,N_6241,N_6007);
and U11882 (N_11882,N_5619,N_7103);
nor U11883 (N_11883,N_7755,N_4099);
and U11884 (N_11884,N_5911,N_4439);
or U11885 (N_11885,N_7404,N_7346);
or U11886 (N_11886,N_6276,N_6488);
nor U11887 (N_11887,N_5622,N_4802);
and U11888 (N_11888,N_4803,N_6737);
and U11889 (N_11889,N_6992,N_5180);
nand U11890 (N_11890,N_5782,N_5296);
nand U11891 (N_11891,N_7739,N_6856);
nor U11892 (N_11892,N_6799,N_7866);
and U11893 (N_11893,N_7086,N_6948);
nand U11894 (N_11894,N_4030,N_5481);
or U11895 (N_11895,N_6786,N_4712);
and U11896 (N_11896,N_7054,N_5572);
xor U11897 (N_11897,N_5844,N_4978);
nand U11898 (N_11898,N_4154,N_4480);
and U11899 (N_11899,N_5257,N_5633);
nor U11900 (N_11900,N_5880,N_7498);
nand U11901 (N_11901,N_7301,N_7414);
or U11902 (N_11902,N_7466,N_4112);
nand U11903 (N_11903,N_4771,N_6552);
or U11904 (N_11904,N_6171,N_5941);
nand U11905 (N_11905,N_4187,N_7106);
nor U11906 (N_11906,N_6366,N_5291);
or U11907 (N_11907,N_7255,N_6003);
nor U11908 (N_11908,N_4182,N_6536);
nor U11909 (N_11909,N_4179,N_6249);
nor U11910 (N_11910,N_4613,N_6458);
or U11911 (N_11911,N_7015,N_6004);
nand U11912 (N_11912,N_6703,N_6519);
or U11913 (N_11913,N_4091,N_7037);
and U11914 (N_11914,N_4204,N_5550);
nor U11915 (N_11915,N_6158,N_6833);
nand U11916 (N_11916,N_4984,N_4309);
or U11917 (N_11917,N_6015,N_4808);
nor U11918 (N_11918,N_6629,N_4904);
nor U11919 (N_11919,N_5913,N_5411);
nor U11920 (N_11920,N_7480,N_6002);
nor U11921 (N_11921,N_5781,N_7046);
and U11922 (N_11922,N_6540,N_5442);
or U11923 (N_11923,N_7943,N_5397);
or U11924 (N_11924,N_6150,N_5285);
or U11925 (N_11925,N_4518,N_4661);
or U11926 (N_11926,N_6135,N_7595);
nor U11927 (N_11927,N_5006,N_4400);
and U11928 (N_11928,N_7180,N_6271);
nand U11929 (N_11929,N_5044,N_5858);
and U11930 (N_11930,N_7188,N_6149);
nand U11931 (N_11931,N_4095,N_5686);
xnor U11932 (N_11932,N_4296,N_7523);
and U11933 (N_11933,N_4369,N_5907);
or U11934 (N_11934,N_4367,N_4066);
xnor U11935 (N_11935,N_5479,N_7867);
nor U11936 (N_11936,N_4029,N_4302);
nand U11937 (N_11937,N_5112,N_5275);
nor U11938 (N_11938,N_4525,N_5154);
or U11939 (N_11939,N_4622,N_5158);
or U11940 (N_11940,N_7117,N_5106);
xnor U11941 (N_11941,N_5683,N_4617);
or U11942 (N_11942,N_6266,N_7180);
nand U11943 (N_11943,N_6744,N_6099);
and U11944 (N_11944,N_7736,N_7402);
or U11945 (N_11945,N_4941,N_5753);
and U11946 (N_11946,N_7635,N_6673);
nand U11947 (N_11947,N_4011,N_5709);
nor U11948 (N_11948,N_5703,N_7787);
xnor U11949 (N_11949,N_6896,N_7585);
or U11950 (N_11950,N_7191,N_6895);
xnor U11951 (N_11951,N_6477,N_6501);
nor U11952 (N_11952,N_7429,N_6944);
xnor U11953 (N_11953,N_5408,N_6594);
xnor U11954 (N_11954,N_4818,N_7058);
nor U11955 (N_11955,N_7727,N_6998);
nand U11956 (N_11956,N_7443,N_4871);
xnor U11957 (N_11957,N_7579,N_4255);
nand U11958 (N_11958,N_7707,N_4720);
nand U11959 (N_11959,N_6005,N_6220);
and U11960 (N_11960,N_7390,N_7018);
or U11961 (N_11961,N_5807,N_5588);
and U11962 (N_11962,N_5598,N_5234);
or U11963 (N_11963,N_7443,N_5587);
xnor U11964 (N_11964,N_6378,N_4903);
nor U11965 (N_11965,N_4692,N_5072);
nor U11966 (N_11966,N_6809,N_5726);
nand U11967 (N_11967,N_4426,N_7650);
xor U11968 (N_11968,N_7680,N_4962);
nand U11969 (N_11969,N_7419,N_4367);
or U11970 (N_11970,N_4558,N_5115);
or U11971 (N_11971,N_5432,N_4713);
or U11972 (N_11972,N_6499,N_5240);
nor U11973 (N_11973,N_7648,N_7064);
nor U11974 (N_11974,N_4268,N_4865);
nor U11975 (N_11975,N_5314,N_6998);
nor U11976 (N_11976,N_6264,N_4596);
nor U11977 (N_11977,N_7846,N_7485);
or U11978 (N_11978,N_5496,N_5663);
or U11979 (N_11979,N_7774,N_5151);
xnor U11980 (N_11980,N_7201,N_4883);
nand U11981 (N_11981,N_7058,N_4333);
or U11982 (N_11982,N_7733,N_7677);
xor U11983 (N_11983,N_5154,N_7430);
or U11984 (N_11984,N_5233,N_4433);
nand U11985 (N_11985,N_7093,N_7879);
and U11986 (N_11986,N_7306,N_5888);
xnor U11987 (N_11987,N_7602,N_5821);
nor U11988 (N_11988,N_4000,N_4248);
nor U11989 (N_11989,N_6578,N_6202);
and U11990 (N_11990,N_5222,N_4770);
nand U11991 (N_11991,N_5287,N_7843);
or U11992 (N_11992,N_5478,N_4960);
and U11993 (N_11993,N_4870,N_6083);
nor U11994 (N_11994,N_6922,N_7752);
or U11995 (N_11995,N_4072,N_6999);
nand U11996 (N_11996,N_4243,N_5226);
and U11997 (N_11997,N_4484,N_5413);
nand U11998 (N_11998,N_7940,N_7011);
and U11999 (N_11999,N_4623,N_7241);
nand U12000 (N_12000,N_10486,N_9295);
and U12001 (N_12001,N_9754,N_11060);
xor U12002 (N_12002,N_11792,N_9127);
xnor U12003 (N_12003,N_11575,N_9411);
nor U12004 (N_12004,N_8833,N_11755);
and U12005 (N_12005,N_10694,N_8778);
or U12006 (N_12006,N_10847,N_10987);
nor U12007 (N_12007,N_8714,N_11611);
and U12008 (N_12008,N_11508,N_11906);
nand U12009 (N_12009,N_10134,N_8489);
or U12010 (N_12010,N_8061,N_9773);
and U12011 (N_12011,N_10647,N_8491);
and U12012 (N_12012,N_10151,N_9720);
nand U12013 (N_12013,N_10029,N_11351);
or U12014 (N_12014,N_10051,N_9925);
and U12015 (N_12015,N_10042,N_11429);
nand U12016 (N_12016,N_8595,N_8636);
xor U12017 (N_12017,N_11426,N_8469);
nand U12018 (N_12018,N_10299,N_9362);
or U12019 (N_12019,N_9821,N_8933);
and U12020 (N_12020,N_8720,N_9971);
nor U12021 (N_12021,N_8166,N_11223);
xnor U12022 (N_12022,N_11872,N_11115);
nand U12023 (N_12023,N_8065,N_10104);
xnor U12024 (N_12024,N_9332,N_10329);
nand U12025 (N_12025,N_11978,N_10210);
and U12026 (N_12026,N_11838,N_8251);
and U12027 (N_12027,N_10657,N_8687);
xor U12028 (N_12028,N_9740,N_8060);
xnor U12029 (N_12029,N_10611,N_8135);
xnor U12030 (N_12030,N_10538,N_10452);
and U12031 (N_12031,N_8516,N_11803);
and U12032 (N_12032,N_9782,N_9824);
xor U12033 (N_12033,N_10767,N_8399);
xnor U12034 (N_12034,N_8622,N_11393);
nand U12035 (N_12035,N_11328,N_9827);
or U12036 (N_12036,N_10145,N_11262);
nor U12037 (N_12037,N_11034,N_11680);
nor U12038 (N_12038,N_11686,N_8233);
or U12039 (N_12039,N_9230,N_9822);
xnor U12040 (N_12040,N_8498,N_10478);
or U12041 (N_12041,N_10750,N_8019);
or U12042 (N_12042,N_9231,N_8904);
nor U12043 (N_12043,N_8403,N_8855);
xnor U12044 (N_12044,N_8841,N_11135);
or U12045 (N_12045,N_10566,N_11161);
nor U12046 (N_12046,N_9061,N_9285);
nand U12047 (N_12047,N_11902,N_11323);
and U12048 (N_12048,N_8635,N_9932);
nand U12049 (N_12049,N_8675,N_11372);
xnor U12050 (N_12050,N_8400,N_11530);
and U12051 (N_12051,N_8144,N_9811);
nand U12052 (N_12052,N_8999,N_10221);
and U12053 (N_12053,N_8073,N_10991);
and U12054 (N_12054,N_8996,N_8850);
and U12055 (N_12055,N_10512,N_8390);
and U12056 (N_12056,N_10632,N_8112);
and U12057 (N_12057,N_9785,N_9561);
nor U12058 (N_12058,N_8197,N_9923);
xor U12059 (N_12059,N_10460,N_10803);
xor U12060 (N_12060,N_8467,N_8838);
nor U12061 (N_12061,N_8965,N_8790);
nand U12062 (N_12062,N_9918,N_9469);
nor U12063 (N_12063,N_9137,N_10619);
nand U12064 (N_12064,N_10164,N_10077);
xor U12065 (N_12065,N_11360,N_10624);
nand U12066 (N_12066,N_11618,N_8523);
xnor U12067 (N_12067,N_10124,N_11566);
nor U12068 (N_12068,N_8101,N_8685);
or U12069 (N_12069,N_9978,N_11016);
nor U12070 (N_12070,N_10895,N_11664);
xnor U12071 (N_12071,N_10935,N_11668);
or U12072 (N_12072,N_8653,N_8842);
xor U12073 (N_12073,N_9000,N_10644);
nand U12074 (N_12074,N_9956,N_8416);
xor U12075 (N_12075,N_11364,N_8995);
nor U12076 (N_12076,N_10214,N_10296);
xnor U12077 (N_12077,N_11879,N_10807);
and U12078 (N_12078,N_11207,N_11312);
and U12079 (N_12079,N_11859,N_11158);
nor U12080 (N_12080,N_9883,N_8663);
or U12081 (N_12081,N_9074,N_11639);
xnor U12082 (N_12082,N_11469,N_10114);
xor U12083 (N_12083,N_8918,N_11368);
nand U12084 (N_12084,N_11754,N_9857);
xor U12085 (N_12085,N_9632,N_11220);
nor U12086 (N_12086,N_11685,N_10468);
nand U12087 (N_12087,N_10626,N_11319);
and U12088 (N_12088,N_11967,N_11747);
nand U12089 (N_12089,N_10359,N_11259);
nand U12090 (N_12090,N_9993,N_9988);
or U12091 (N_12091,N_8555,N_9123);
xnor U12092 (N_12092,N_11420,N_11850);
and U12093 (N_12093,N_9159,N_8621);
or U12094 (N_12094,N_8844,N_11586);
nor U12095 (N_12095,N_11828,N_11149);
nor U12096 (N_12096,N_8591,N_9083);
and U12097 (N_12097,N_8753,N_10614);
xnor U12098 (N_12098,N_10977,N_11102);
nand U12099 (N_12099,N_9305,N_8564);
or U12100 (N_12100,N_11973,N_8449);
or U12101 (N_12101,N_10113,N_9693);
nor U12102 (N_12102,N_10787,N_8150);
nor U12103 (N_12103,N_9766,N_9394);
xnor U12104 (N_12104,N_10976,N_9809);
and U12105 (N_12105,N_11403,N_11235);
xnor U12106 (N_12106,N_11009,N_9535);
or U12107 (N_12107,N_8590,N_9952);
or U12108 (N_12108,N_9694,N_10382);
xor U12109 (N_12109,N_11539,N_10660);
nor U12110 (N_12110,N_9313,N_11271);
or U12111 (N_12111,N_9338,N_11209);
or U12112 (N_12112,N_8039,N_9086);
and U12113 (N_12113,N_11437,N_9171);
or U12114 (N_12114,N_11272,N_10068);
xor U12115 (N_12115,N_8447,N_8815);
xor U12116 (N_12116,N_9335,N_8345);
nand U12117 (N_12117,N_8473,N_8169);
xnor U12118 (N_12118,N_8199,N_8957);
and U12119 (N_12119,N_9975,N_11627);
nor U12120 (N_12120,N_8160,N_9448);
or U12121 (N_12121,N_10870,N_11784);
xor U12122 (N_12122,N_8897,N_11518);
xnor U12123 (N_12123,N_11538,N_11399);
or U12124 (N_12124,N_9807,N_10677);
xor U12125 (N_12125,N_11369,N_8533);
nor U12126 (N_12126,N_9708,N_8470);
or U12127 (N_12127,N_8421,N_8003);
or U12128 (N_12128,N_11637,N_11713);
nand U12129 (N_12129,N_11951,N_8984);
nand U12130 (N_12130,N_9985,N_10695);
or U12131 (N_12131,N_11744,N_8149);
nor U12132 (N_12132,N_9314,N_11252);
or U12133 (N_12133,N_9840,N_8924);
and U12134 (N_12134,N_11735,N_10656);
and U12135 (N_12135,N_9899,N_9795);
nand U12136 (N_12136,N_9436,N_11712);
xnor U12137 (N_12137,N_11365,N_8091);
nor U12138 (N_12138,N_10858,N_8802);
xor U12139 (N_12139,N_11127,N_10148);
and U12140 (N_12140,N_11204,N_11848);
xnor U12141 (N_12141,N_8366,N_8292);
and U12142 (N_12142,N_10588,N_10251);
nand U12143 (N_12143,N_9960,N_9351);
or U12144 (N_12144,N_11563,N_10048);
or U12145 (N_12145,N_8810,N_9623);
and U12146 (N_12146,N_8701,N_10852);
and U12147 (N_12147,N_9427,N_10794);
nand U12148 (N_12148,N_10314,N_11985);
and U12149 (N_12149,N_10628,N_11245);
and U12150 (N_12150,N_8515,N_10992);
and U12151 (N_12151,N_8444,N_11417);
or U12152 (N_12152,N_8066,N_10000);
xnor U12153 (N_12153,N_8293,N_9750);
nand U12154 (N_12154,N_11044,N_11653);
and U12155 (N_12155,N_11750,N_9024);
or U12156 (N_12156,N_8938,N_9103);
or U12157 (N_12157,N_10899,N_10203);
xnor U12158 (N_12158,N_11845,N_11304);
xor U12159 (N_12159,N_11793,N_11844);
nor U12160 (N_12160,N_8982,N_8228);
nor U12161 (N_12161,N_9528,N_8495);
xnor U12162 (N_12162,N_11876,N_11242);
nand U12163 (N_12163,N_8089,N_11684);
nand U12164 (N_12164,N_8313,N_9611);
and U12165 (N_12165,N_8243,N_11296);
and U12166 (N_12166,N_10594,N_8905);
nand U12167 (N_12167,N_9915,N_8626);
or U12168 (N_12168,N_11382,N_11960);
nor U12169 (N_12169,N_11352,N_8425);
xnor U12170 (N_12170,N_8227,N_8528);
and U12171 (N_12171,N_11896,N_10336);
nor U12172 (N_12172,N_11214,N_10881);
nand U12173 (N_12173,N_8979,N_11631);
or U12174 (N_12174,N_8411,N_11086);
and U12175 (N_12175,N_10401,N_11534);
or U12176 (N_12176,N_10685,N_9896);
or U12177 (N_12177,N_8623,N_8038);
and U12178 (N_12178,N_8868,N_9633);
nor U12179 (N_12179,N_8071,N_10716);
xnor U12180 (N_12180,N_8886,N_11385);
nor U12181 (N_12181,N_10204,N_10244);
nor U12182 (N_12182,N_8634,N_11533);
nand U12183 (N_12183,N_11432,N_10076);
nor U12184 (N_12184,N_9431,N_9062);
or U12185 (N_12185,N_11672,N_9386);
or U12186 (N_12186,N_9280,N_11972);
and U12187 (N_12187,N_9742,N_8602);
nand U12188 (N_12188,N_9818,N_8225);
nand U12189 (N_12189,N_8121,N_11455);
or U12190 (N_12190,N_11742,N_10256);
or U12191 (N_12191,N_10437,N_9038);
and U12192 (N_12192,N_8884,N_10617);
nor U12193 (N_12193,N_11461,N_11035);
and U12194 (N_12194,N_8364,N_10868);
nand U12195 (N_12195,N_9713,N_11472);
nand U12196 (N_12196,N_9626,N_8682);
xnor U12197 (N_12197,N_10719,N_9381);
xor U12198 (N_12198,N_8238,N_9449);
or U12199 (N_12199,N_9525,N_11094);
xnor U12200 (N_12200,N_11769,N_8812);
and U12201 (N_12201,N_8485,N_11689);
xnor U12202 (N_12202,N_10489,N_9120);
nand U12203 (N_12203,N_11552,N_9410);
nor U12204 (N_12204,N_11356,N_8154);
or U12205 (N_12205,N_9892,N_8214);
nor U12206 (N_12206,N_8354,N_11305);
nor U12207 (N_12207,N_8269,N_8102);
xnor U12208 (N_12208,N_9666,N_8876);
xor U12209 (N_12209,N_11887,N_11333);
nor U12210 (N_12210,N_11760,N_8240);
nor U12211 (N_12211,N_8723,N_9251);
nand U12212 (N_12212,N_11334,N_8341);
or U12213 (N_12213,N_11775,N_10763);
nand U12214 (N_12214,N_8804,N_10817);
nor U12215 (N_12215,N_8156,N_11613);
or U12216 (N_12216,N_11782,N_11173);
and U12217 (N_12217,N_9030,N_9319);
nor U12218 (N_12218,N_11743,N_8417);
and U12219 (N_12219,N_8779,N_10737);
and U12220 (N_12220,N_9378,N_10914);
nor U12221 (N_12221,N_11337,N_10886);
nand U12222 (N_12222,N_11453,N_10348);
nor U12223 (N_12223,N_9894,N_11979);
nor U12224 (N_12224,N_8527,N_9711);
nor U12225 (N_12225,N_9185,N_8207);
nor U12226 (N_12226,N_8330,N_11598);
nand U12227 (N_12227,N_10430,N_11059);
nand U12228 (N_12228,N_10843,N_9584);
or U12229 (N_12229,N_11075,N_8552);
nand U12230 (N_12230,N_10574,N_8005);
nand U12231 (N_12231,N_9279,N_9329);
xnor U12232 (N_12232,N_10412,N_8806);
nor U12233 (N_12233,N_10383,N_11055);
and U12234 (N_12234,N_11907,N_11936);
or U12235 (N_12235,N_8603,N_11033);
and U12236 (N_12236,N_8586,N_11988);
or U12237 (N_12237,N_10150,N_8923);
nand U12238 (N_12238,N_9092,N_10971);
or U12239 (N_12239,N_9296,N_9908);
nor U12240 (N_12240,N_8404,N_9169);
or U12241 (N_12241,N_8617,N_10319);
or U12242 (N_12242,N_10264,N_9580);
nor U12243 (N_12243,N_9897,N_8029);
and U12244 (N_12244,N_8284,N_9530);
nand U12245 (N_12245,N_10679,N_10398);
or U12246 (N_12246,N_8879,N_11602);
or U12247 (N_12247,N_10089,N_10200);
and U12248 (N_12248,N_8111,N_9593);
nor U12249 (N_12249,N_11152,N_8832);
or U12250 (N_12250,N_11609,N_10833);
xnor U12251 (N_12251,N_8713,N_8215);
or U12252 (N_12252,N_8769,N_9316);
or U12253 (N_12253,N_8670,N_11662);
xor U12254 (N_12254,N_8624,N_10438);
and U12255 (N_12255,N_8948,N_10072);
xor U12256 (N_12256,N_10321,N_11159);
nor U12257 (N_12257,N_11180,N_9508);
and U12258 (N_12258,N_8711,N_10819);
xnor U12259 (N_12259,N_10826,N_10380);
nand U12260 (N_12260,N_10427,N_8993);
and U12261 (N_12261,N_9813,N_9532);
and U12262 (N_12262,N_9933,N_8182);
xnor U12263 (N_12263,N_9346,N_10111);
xor U12264 (N_12264,N_11338,N_9376);
nand U12265 (N_12265,N_10050,N_10127);
xnor U12266 (N_12266,N_9138,N_11423);
xor U12267 (N_12267,N_10715,N_9459);
nor U12268 (N_12268,N_9273,N_8695);
or U12269 (N_12269,N_9458,N_8631);
nand U12270 (N_12270,N_8335,N_11700);
xor U12271 (N_12271,N_8654,N_10394);
nor U12272 (N_12272,N_11343,N_11422);
or U12273 (N_12273,N_8749,N_8070);
xor U12274 (N_12274,N_10254,N_10934);
or U12275 (N_12275,N_10567,N_8232);
and U12276 (N_12276,N_9465,N_11787);
nor U12277 (N_12277,N_8348,N_8762);
or U12278 (N_12278,N_11720,N_8656);
and U12279 (N_12279,N_9499,N_11506);
nand U12280 (N_12280,N_10900,N_10302);
nand U12281 (N_12281,N_11039,N_11504);
and U12282 (N_12282,N_9423,N_8170);
xnor U12283 (N_12283,N_11258,N_10268);
and U12284 (N_12284,N_10549,N_10506);
nand U12285 (N_12285,N_11625,N_11568);
and U12286 (N_12286,N_11977,N_8519);
nand U12287 (N_12287,N_10109,N_11435);
nor U12288 (N_12288,N_8322,N_10183);
nand U12289 (N_12289,N_9622,N_10691);
and U12290 (N_12290,N_10283,N_11624);
nor U12291 (N_12291,N_9311,N_11064);
nand U12292 (N_12292,N_10032,N_8488);
or U12293 (N_12293,N_11778,N_11541);
xnor U12294 (N_12294,N_8852,N_8194);
and U12295 (N_12295,N_11468,N_8480);
nand U12296 (N_12296,N_8807,N_9594);
nor U12297 (N_12297,N_11766,N_8543);
and U12298 (N_12298,N_10056,N_11080);
and U12299 (N_12299,N_11647,N_8766);
xnor U12300 (N_12300,N_8601,N_8683);
or U12301 (N_12301,N_9865,N_8800);
nor U12302 (N_12302,N_9921,N_10101);
and U12303 (N_12303,N_10045,N_10206);
nor U12304 (N_12304,N_8817,N_11120);
nor U12305 (N_12305,N_10673,N_9064);
nand U12306 (N_12306,N_8064,N_8556);
xor U12307 (N_12307,N_9603,N_11719);
and U12308 (N_12308,N_9578,N_11724);
and U12309 (N_12309,N_11234,N_11615);
nand U12310 (N_12310,N_10376,N_11137);
and U12311 (N_12311,N_11567,N_8704);
xnor U12312 (N_12312,N_11141,N_8420);
xnor U12313 (N_12313,N_8037,N_11354);
nand U12314 (N_12314,N_11721,N_8406);
nor U12315 (N_12315,N_11903,N_9849);
or U12316 (N_12316,N_8946,N_8945);
xor U12317 (N_12317,N_11546,N_8895);
and U12318 (N_12318,N_8192,N_8090);
nand U12319 (N_12319,N_9791,N_8718);
xor U12320 (N_12320,N_10196,N_8497);
or U12321 (N_12321,N_11544,N_11826);
or U12322 (N_12322,N_11537,N_11893);
or U12323 (N_12323,N_10809,N_10562);
nand U12324 (N_12324,N_11666,N_11431);
nor U12325 (N_12325,N_10553,N_9806);
or U12326 (N_12326,N_11248,N_8853);
nor U12327 (N_12327,N_11677,N_9704);
or U12328 (N_12328,N_8566,N_11278);
nor U12329 (N_12329,N_8964,N_10587);
nand U12330 (N_12330,N_9384,N_8963);
xnor U12331 (N_12331,N_10088,N_11197);
or U12332 (N_12332,N_10026,N_10022);
xnor U12333 (N_12333,N_8319,N_11361);
nand U12334 (N_12334,N_11324,N_9100);
or U12335 (N_12335,N_8051,N_10525);
or U12336 (N_12336,N_11881,N_11147);
nand U12337 (N_12337,N_10205,N_9223);
nor U12338 (N_12338,N_11083,N_9730);
or U12339 (N_12339,N_8575,N_11679);
and U12340 (N_12340,N_11938,N_11731);
and U12341 (N_12341,N_9728,N_10238);
xnor U12342 (N_12342,N_8068,N_10707);
or U12343 (N_12343,N_8840,N_11722);
and U12344 (N_12344,N_11641,N_10721);
or U12345 (N_12345,N_9589,N_8347);
or U12346 (N_12346,N_11971,N_11692);
nand U12347 (N_12347,N_10568,N_8678);
xor U12348 (N_12348,N_11867,N_9571);
and U12349 (N_12349,N_10778,N_10988);
and U12350 (N_12350,N_9228,N_8477);
xor U12351 (N_12351,N_11471,N_10651);
or U12352 (N_12352,N_10516,N_8268);
xnor U12353 (N_12353,N_11975,N_10573);
nor U12354 (N_12354,N_8652,N_9526);
nor U12355 (N_12355,N_11619,N_11433);
or U12356 (N_12356,N_11196,N_10649);
and U12357 (N_12357,N_10704,N_9003);
or U12358 (N_12358,N_11154,N_8981);
nand U12359 (N_12359,N_10297,N_9113);
or U12360 (N_12360,N_9540,N_8805);
nor U12361 (N_12361,N_8605,N_9333);
xnor U12362 (N_12362,N_10600,N_11911);
and U12363 (N_12363,N_10927,N_11134);
and U12364 (N_12364,N_9205,N_9710);
xor U12365 (N_12365,N_9702,N_10073);
and U12366 (N_12366,N_9267,N_9174);
nand U12367 (N_12367,N_11790,N_9390);
xor U12368 (N_12368,N_10755,N_11184);
nand U12369 (N_12369,N_11600,N_9581);
nor U12370 (N_12370,N_9035,N_10867);
nor U12371 (N_12371,N_9013,N_8304);
nor U12372 (N_12372,N_8359,N_10931);
or U12373 (N_12373,N_10292,N_10240);
xnor U12374 (N_12374,N_8357,N_11583);
and U12375 (N_12375,N_9276,N_10173);
nand U12376 (N_12376,N_9794,N_8715);
and U12377 (N_12377,N_11999,N_11189);
or U12378 (N_12378,N_11163,N_8198);
or U12379 (N_12379,N_11373,N_8930);
and U12380 (N_12380,N_11551,N_11560);
nand U12381 (N_12381,N_10890,N_8889);
nor U12382 (N_12382,N_9480,N_8503);
and U12383 (N_12383,N_9999,N_8901);
and U12384 (N_12384,N_11132,N_9027);
or U12385 (N_12385,N_11610,N_8024);
xnor U12386 (N_12386,N_11481,N_8862);
and U12387 (N_12387,N_10255,N_11375);
nor U12388 (N_12388,N_8740,N_11236);
nand U12389 (N_12389,N_9845,N_9793);
nor U12390 (N_12390,N_9732,N_8735);
and U12391 (N_12391,N_11962,N_9995);
and U12392 (N_12392,N_8151,N_9360);
nor U12393 (N_12393,N_8450,N_8791);
and U12394 (N_12394,N_9825,N_10492);
nor U12395 (N_12395,N_11047,N_10597);
or U12396 (N_12396,N_10764,N_10693);
nand U12397 (N_12397,N_10207,N_10869);
nor U12398 (N_12398,N_10970,N_11465);
and U12399 (N_12399,N_10317,N_11652);
nand U12400 (N_12400,N_10387,N_9916);
nand U12401 (N_12401,N_11202,N_11557);
nor U12402 (N_12402,N_10179,N_9033);
nand U12403 (N_12403,N_9667,N_10634);
and U12404 (N_12404,N_8526,N_8312);
and U12405 (N_12405,N_9778,N_10313);
xor U12406 (N_12406,N_11952,N_9422);
nand U12407 (N_12407,N_8052,N_8321);
or U12408 (N_12408,N_11108,N_9037);
xor U12409 (N_12409,N_10702,N_9789);
and U12410 (N_12410,N_9986,N_11063);
nand U12411 (N_12411,N_10547,N_8258);
nor U12412 (N_12412,N_10655,N_11340);
xnor U12413 (N_12413,N_11010,N_11443);
xor U12414 (N_12414,N_9587,N_9922);
nand U12415 (N_12415,N_11190,N_11029);
nand U12416 (N_12416,N_9810,N_9537);
xor U12417 (N_12417,N_11263,N_8205);
nand U12418 (N_12418,N_8922,N_8985);
nand U12419 (N_12419,N_8544,N_11933);
or U12420 (N_12420,N_9025,N_9592);
nand U12421 (N_12421,N_9853,N_8970);
nand U12422 (N_12422,N_8463,N_10783);
xnor U12423 (N_12423,N_8794,N_11756);
or U12424 (N_12424,N_8576,N_11232);
nor U12425 (N_12425,N_8476,N_10324);
nor U12426 (N_12426,N_8742,N_8496);
and U12427 (N_12427,N_8158,N_10269);
and U12428 (N_12428,N_9719,N_8725);
nor U12429 (N_12429,N_11847,N_10410);
or U12430 (N_12430,N_11909,N_10137);
and U12431 (N_12431,N_8422,N_10342);
xor U12432 (N_12432,N_9884,N_8407);
xnor U12433 (N_12433,N_9392,N_8758);
or U12434 (N_12434,N_9218,N_10305);
xnor U12435 (N_12435,N_9399,N_8655);
nor U12436 (N_12436,N_10237,N_8989);
nor U12437 (N_12437,N_11384,N_9082);
and U12438 (N_12438,N_8373,N_11941);
xnor U12439 (N_12439,N_10316,N_9124);
nand U12440 (N_12440,N_9429,N_10245);
nor U12441 (N_12441,N_11852,N_9557);
nand U12442 (N_12442,N_10772,N_8282);
or U12443 (N_12443,N_10175,N_10580);
nor U12444 (N_12444,N_11717,N_9400);
or U12445 (N_12445,N_10084,N_8569);
xor U12446 (N_12446,N_9637,N_9681);
and U12447 (N_12447,N_8380,N_10092);
nand U12448 (N_12448,N_9753,N_9536);
nor U12449 (N_12449,N_10864,N_10170);
nor U12450 (N_12450,N_10793,N_8415);
and U12451 (N_12451,N_10945,N_10328);
or U12452 (N_12452,N_10020,N_8317);
or U12453 (N_12453,N_11707,N_11066);
nand U12454 (N_12454,N_11379,N_9647);
or U12455 (N_12455,N_11581,N_9520);
nand U12456 (N_12456,N_9767,N_10820);
xor U12457 (N_12457,N_10083,N_11993);
or U12458 (N_12458,N_10766,N_11317);
and U12459 (N_12459,N_9900,N_11483);
nor U12460 (N_12460,N_8696,N_8358);
nand U12461 (N_12461,N_11122,N_11839);
xnor U12462 (N_12462,N_8370,N_8218);
xor U12463 (N_12463,N_11485,N_8332);
xnor U12464 (N_12464,N_9690,N_9457);
and U12465 (N_12465,N_10711,N_10855);
and U12466 (N_12466,N_8176,N_9182);
xnor U12467 (N_12467,N_11400,N_11133);
nand U12468 (N_12468,N_11545,N_8303);
xnor U12469 (N_12469,N_9856,N_8055);
or U12470 (N_12470,N_10469,N_11331);
nand U12471 (N_12471,N_10335,N_9072);
or U12472 (N_12472,N_9168,N_10675);
nand U12473 (N_12473,N_9109,N_8222);
xnor U12474 (N_12474,N_11843,N_9725);
nor U12475 (N_12475,N_11771,N_8427);
or U12476 (N_12476,N_11968,N_10683);
nand U12477 (N_12477,N_10643,N_9541);
nor U12478 (N_12478,N_10922,N_10005);
or U12479 (N_12479,N_9406,N_9848);
or U12480 (N_12480,N_9248,N_8860);
xor U12481 (N_12481,N_8123,N_10075);
nor U12482 (N_12482,N_10454,N_8223);
and U12483 (N_12483,N_10968,N_9660);
nor U12484 (N_12484,N_11145,N_8035);
and U12485 (N_12485,N_8761,N_9391);
and U12486 (N_12486,N_8436,N_9984);
nor U12487 (N_12487,N_9761,N_11148);
nor U12488 (N_12488,N_9680,N_8919);
nand U12489 (N_12489,N_8372,N_10768);
xor U12490 (N_12490,N_9359,N_11621);
xnor U12491 (N_12491,N_11057,N_9885);
and U12492 (N_12492,N_10239,N_9602);
or U12493 (N_12493,N_9994,N_11654);
or U12494 (N_12494,N_11899,N_10872);
xnor U12495 (N_12495,N_9101,N_8186);
xnor U12496 (N_12496,N_10105,N_10246);
nand U12497 (N_12497,N_10197,N_8075);
or U12498 (N_12498,N_11620,N_10749);
nor U12499 (N_12499,N_11617,N_9902);
or U12500 (N_12500,N_9017,N_10458);
nand U12501 (N_12501,N_9253,N_11162);
and U12502 (N_12502,N_10474,N_8201);
xnor U12503 (N_12503,N_11438,N_8729);
and U12504 (N_12504,N_11576,N_8961);
nor U12505 (N_12505,N_9403,N_9613);
or U12506 (N_12506,N_9692,N_10609);
or U12507 (N_12507,N_11298,N_9158);
nand U12508 (N_12508,N_10877,N_9322);
nand U12509 (N_12509,N_11723,N_10668);
and U12510 (N_12510,N_11030,N_9860);
xnor U12511 (N_12511,N_9321,N_11591);
nand U12512 (N_12512,N_10692,N_10709);
nor U12513 (N_12513,N_11470,N_10701);
and U12514 (N_12514,N_9555,N_10873);
xor U12515 (N_12515,N_9347,N_11124);
nand U12516 (N_12516,N_10080,N_10365);
nand U12517 (N_12517,N_9365,N_11413);
xnor U12518 (N_12518,N_10208,N_9277);
and U12519 (N_12519,N_9595,N_8187);
and U12520 (N_12520,N_9928,N_10323);
xnor U12521 (N_12521,N_8677,N_10355);
nor U12522 (N_12522,N_8632,N_10569);
nand U12523 (N_12523,N_8693,N_11231);
xor U12524 (N_12524,N_11300,N_9832);
nand U12525 (N_12525,N_10937,N_11737);
nand U12526 (N_12526,N_9619,N_9706);
nor U12527 (N_12527,N_11153,N_10194);
nand U12528 (N_12528,N_9598,N_8974);
or U12529 (N_12529,N_10790,N_11728);
nand U12530 (N_12530,N_11752,N_8589);
nor U12531 (N_12531,N_8826,N_8152);
nand U12532 (N_12532,N_11498,N_10747);
nand U12533 (N_12533,N_8958,N_11980);
nor U12534 (N_12534,N_11405,N_11346);
nand U12535 (N_12535,N_8139,N_10161);
and U12536 (N_12536,N_10714,N_11556);
or U12537 (N_12537,N_11604,N_8582);
or U12538 (N_12538,N_10360,N_10663);
nand U12539 (N_12539,N_11812,N_11386);
nor U12540 (N_12540,N_9664,N_10054);
or U12541 (N_12541,N_11897,N_11846);
xnor U12542 (N_12542,N_9797,N_8874);
xor U12543 (N_12543,N_10878,N_10825);
nand U12544 (N_12544,N_8661,N_10658);
nand U12545 (N_12545,N_10120,N_11114);
and U12546 (N_12546,N_8746,N_9377);
or U12547 (N_12547,N_11517,N_8615);
xnor U12548 (N_12548,N_10505,N_9746);
nor U12549 (N_12549,N_10172,N_9585);
and U12550 (N_12550,N_10182,N_11448);
xor U12551 (N_12551,N_9968,N_10061);
or U12552 (N_12552,N_9393,N_11306);
or U12553 (N_12553,N_10907,N_11446);
nand U12554 (N_12554,N_11415,N_10774);
xor U12555 (N_12555,N_9320,N_8706);
nand U12556 (N_12556,N_8609,N_8517);
nand U12557 (N_12557,N_9575,N_8820);
and U12558 (N_12558,N_8445,N_9247);
or U12559 (N_12559,N_10738,N_8988);
xor U12560 (N_12560,N_10728,N_9250);
and U12561 (N_12561,N_8062,N_9938);
nor U12562 (N_12562,N_11491,N_9868);
nand U12563 (N_12563,N_9831,N_11525);
xnor U12564 (N_12564,N_10964,N_8834);
nor U12565 (N_12565,N_11901,N_9076);
or U12566 (N_12566,N_10470,N_9190);
nand U12567 (N_12567,N_9770,N_8752);
nor U12568 (N_12568,N_10304,N_11182);
nand U12569 (N_12569,N_10641,N_10635);
xor U12570 (N_12570,N_8045,N_8865);
and U12571 (N_12571,N_8505,N_9287);
xor U12572 (N_12572,N_11486,N_11165);
xor U12573 (N_12573,N_8026,N_11274);
and U12574 (N_12574,N_11428,N_10333);
nand U12575 (N_12575,N_10834,N_8600);
and U12576 (N_12576,N_8242,N_10112);
or U12577 (N_12577,N_9880,N_11878);
xor U12578 (N_12578,N_10717,N_9997);
or U12579 (N_12579,N_10053,N_9864);
xnor U12580 (N_12580,N_10443,N_9662);
xnor U12581 (N_12581,N_10924,N_11592);
and U12582 (N_12582,N_10584,N_11487);
and U12583 (N_12583,N_10144,N_8795);
xor U12584 (N_12584,N_11194,N_11579);
or U12585 (N_12585,N_9395,N_10910);
or U12586 (N_12586,N_8353,N_9010);
or U12587 (N_12587,N_9208,N_8103);
xnor U12588 (N_12588,N_9430,N_11763);
or U12589 (N_12589,N_11215,N_8108);
nor U12590 (N_12590,N_9042,N_8881);
nor U12591 (N_12591,N_8162,N_10653);
xor U12592 (N_12592,N_8368,N_9291);
or U12593 (N_12593,N_11820,N_8520);
nand U12594 (N_12594,N_10422,N_10533);
or U12595 (N_12595,N_11806,N_9172);
and U12596 (N_12596,N_8314,N_9189);
or U12597 (N_12597,N_10479,N_8927);
nand U12598 (N_12598,N_9866,N_10542);
xor U12599 (N_12599,N_11674,N_9309);
xor U12600 (N_12600,N_10284,N_9197);
or U12601 (N_12601,N_11005,N_8883);
nor U12602 (N_12602,N_9191,N_11228);
nor U12603 (N_12603,N_10842,N_9886);
and U12604 (N_12604,N_11661,N_8960);
or U12605 (N_12605,N_11799,N_11418);
nor U12606 (N_12606,N_8069,N_10229);
and U12607 (N_12607,N_10110,N_11589);
or U12608 (N_12608,N_10374,N_9389);
nand U12609 (N_12609,N_10429,N_8393);
or U12610 (N_12610,N_9128,N_10928);
or U12611 (N_12611,N_9015,N_9252);
nand U12612 (N_12612,N_8522,N_10485);
and U12613 (N_12613,N_8630,N_10142);
xor U12614 (N_12614,N_9246,N_11705);
and U12615 (N_12615,N_9130,N_11053);
xnor U12616 (N_12616,N_9198,N_11345);
or U12617 (N_12617,N_11380,N_9207);
nor U12618 (N_12618,N_9563,N_9743);
nand U12619 (N_12619,N_11014,N_8098);
and U12620 (N_12620,N_8266,N_9841);
and U12621 (N_12621,N_11396,N_9605);
nor U12622 (N_12622,N_9370,N_9088);
nor U12623 (N_12623,N_10350,N_8259);
and U12624 (N_12624,N_9616,N_9302);
nand U12625 (N_12625,N_10467,N_8819);
nand U12626 (N_12626,N_8466,N_11739);
xnor U12627 (N_12627,N_11482,N_9047);
xor U12628 (N_12628,N_10232,N_10493);
nand U12629 (N_12629,N_11270,N_8639);
nor U12630 (N_12630,N_9511,N_11004);
xor U12631 (N_12631,N_11489,N_11326);
or U12632 (N_12632,N_11942,N_11953);
nor U12633 (N_12633,N_10720,N_11050);
nor U12634 (N_12634,N_8598,N_11176);
xor U12635 (N_12635,N_11265,N_10300);
and U12636 (N_12636,N_11217,N_10638);
xor U12637 (N_12637,N_11836,N_8885);
or U12638 (N_12638,N_11175,N_11956);
nor U12639 (N_12639,N_9876,N_10781);
xnor U12640 (N_12640,N_8221,N_11411);
xnor U12641 (N_12641,N_10500,N_9946);
nor U12642 (N_12642,N_8046,N_8684);
nand U12643 (N_12643,N_10499,N_10098);
xor U12644 (N_12644,N_10322,N_9747);
xnor U12645 (N_12645,N_11996,N_11097);
or U12646 (N_12646,N_11244,N_8699);
and U12647 (N_12647,N_10497,N_10372);
or U12648 (N_12648,N_9361,N_9917);
nand U12649 (N_12649,N_11753,N_11377);
nand U12650 (N_12650,N_8383,N_9278);
nand U12651 (N_12651,N_10689,N_11529);
or U12652 (N_12652,N_8990,N_10598);
or U12653 (N_12653,N_9031,N_11822);
nor U12654 (N_12654,N_11330,N_8195);
nor U12655 (N_12655,N_8086,N_9714);
or U12656 (N_12656,N_10381,N_9052);
nand U12657 (N_12657,N_10276,N_10126);
xnor U12658 (N_12658,N_11578,N_10059);
and U12659 (N_12659,N_10532,N_10259);
nor U12660 (N_12660,N_10769,N_10920);
xor U12661 (N_12661,N_8869,N_9787);
xor U12662 (N_12662,N_8487,N_11054);
and U12663 (N_12663,N_8129,N_8759);
nand U12664 (N_12664,N_10442,N_10997);
nand U12665 (N_12665,N_11842,N_11570);
nand U12666 (N_12666,N_10217,N_8140);
and U12667 (N_12667,N_11247,N_9345);
nand U12668 (N_12668,N_11067,N_8570);
xor U12669 (N_12669,N_9407,N_8471);
and U12670 (N_12670,N_11995,N_10713);
and U12671 (N_12671,N_11089,N_11535);
xor U12672 (N_12672,N_8327,N_8703);
xor U12673 (N_12673,N_8917,N_11796);
or U12674 (N_12674,N_10631,N_9646);
and U12675 (N_12675,N_9944,N_9142);
and U12676 (N_12676,N_11288,N_9648);
and U12677 (N_12677,N_9135,N_11006);
nand U12678 (N_12678,N_10058,N_9259);
xor U12679 (N_12679,N_10223,N_10610);
nand U12680 (N_12680,N_11816,N_8365);
xor U12681 (N_12681,N_8934,N_9586);
nand U12682 (N_12682,N_8584,N_9254);
and U12683 (N_12683,N_11841,N_11745);
xor U12684 (N_12684,N_9485,N_9951);
xnor U12685 (N_12685,N_11976,N_8835);
xor U12686 (N_12686,N_9550,N_10247);
and U12687 (N_12687,N_8780,N_9227);
or U12688 (N_12688,N_11531,N_11947);
nand U12689 (N_12689,N_8648,N_11320);
or U12690 (N_12690,N_9105,N_9566);
or U12691 (N_12691,N_10583,N_9166);
and U12692 (N_12692,N_9504,N_8732);
xnor U12693 (N_12693,N_10267,N_9745);
nand U12694 (N_12694,N_9548,N_8234);
nand U12695 (N_12695,N_9687,N_10243);
xor U12696 (N_12696,N_10565,N_8827);
nor U12697 (N_12697,N_11521,N_10307);
and U12698 (N_12698,N_9873,N_9122);
and U12699 (N_12699,N_9863,N_8264);
and U12700 (N_12700,N_11548,N_9119);
nor U12701 (N_12701,N_8565,N_10887);
xor U12702 (N_12702,N_8773,N_8510);
xor U12703 (N_12703,N_11681,N_8125);
nor U12704 (N_12704,N_10535,N_11629);
or U12705 (N_12705,N_10212,N_9910);
nor U12706 (N_12706,N_9981,N_10132);
nor U12707 (N_12707,N_9601,N_8118);
or U12708 (N_12708,N_8305,N_11930);
xor U12709 (N_12709,N_9089,N_11187);
or U12710 (N_12710,N_8702,N_10162);
xnor U12711 (N_12711,N_9979,N_8754);
xor U12712 (N_12712,N_9569,N_8694);
nand U12713 (N_12713,N_10974,N_10520);
and U12714 (N_12714,N_10613,N_11018);
and U12715 (N_12715,N_9972,N_10403);
nand U12716 (N_12716,N_9736,N_11948);
nor U12717 (N_12717,N_8535,N_10501);
nand U12718 (N_12718,N_10969,N_11238);
nand U12719 (N_12719,N_9415,N_10057);
and U12720 (N_12720,N_8512,N_8968);
xor U12721 (N_12721,N_11606,N_9420);
nand U12722 (N_12722,N_10659,N_9869);
nand U12723 (N_12723,N_8482,N_10289);
and U12724 (N_12724,N_8439,N_8032);
and U12725 (N_12725,N_11221,N_10046);
nor U12726 (N_12726,N_8311,N_8597);
nor U12727 (N_12727,N_11751,N_8451);
nor U12728 (N_12728,N_9163,N_11359);
nand U12729 (N_12729,N_10923,N_9147);
xnor U12730 (N_12730,N_11031,N_9355);
and U12731 (N_12731,N_9658,N_10178);
and U12732 (N_12732,N_8921,N_8698);
or U12733 (N_12733,N_8915,N_8942);
xnor U12734 (N_12734,N_8360,N_8916);
and U12735 (N_12735,N_11023,N_8388);
nand U12736 (N_12736,N_10531,N_11110);
nand U12737 (N_12737,N_8287,N_8574);
and U12738 (N_12738,N_9552,N_10352);
and U12739 (N_12739,N_10522,N_9628);
and U12740 (N_12740,N_8627,N_10191);
nand U12741 (N_12741,N_8343,N_11507);
or U12742 (N_12742,N_10028,N_11922);
nand U12743 (N_12743,N_9644,N_8438);
nor U12744 (N_12744,N_10473,N_9492);
or U12745 (N_12745,N_10851,N_10414);
nand U12746 (N_12746,N_11857,N_8596);
or U12747 (N_12747,N_11068,N_8339);
or U12748 (N_12748,N_10616,N_8502);
and U12749 (N_12749,N_9851,N_8900);
and U12750 (N_12750,N_8208,N_9201);
nand U12751 (N_12751,N_11167,N_10883);
xnor U12752 (N_12752,N_10282,N_9513);
or U12753 (N_12753,N_10160,N_8642);
xnor U12754 (N_12754,N_9518,N_9294);
nor U12755 (N_12755,N_8458,N_10889);
xnor U12756 (N_12756,N_8730,N_10235);
and U12757 (N_12757,N_9094,N_11797);
or U12758 (N_12758,N_8031,N_10761);
or U12759 (N_12759,N_8418,N_11358);
and U12760 (N_12760,N_9272,N_8736);
and U12761 (N_12761,N_11098,N_8295);
nand U12762 (N_12762,N_10963,N_10687);
nand U12763 (N_12763,N_10027,N_8787);
nor U12764 (N_12764,N_11725,N_11107);
and U12765 (N_12765,N_9855,N_10786);
xor U12766 (N_12766,N_11282,N_8457);
or U12767 (N_12767,N_11397,N_8953);
xor U12768 (N_12768,N_11253,N_8454);
nand U12769 (N_12769,N_9502,N_9051);
or U12770 (N_12770,N_9668,N_11366);
and U12771 (N_12771,N_9939,N_11254);
or U12772 (N_12772,N_9405,N_9924);
xor U12773 (N_12773,N_11036,N_10391);
and U12774 (N_12774,N_8285,N_11950);
and U12775 (N_12775,N_11439,N_9695);
nand U12776 (N_12776,N_9665,N_8018);
xnor U12777 (N_12777,N_8494,N_10388);
and U12778 (N_12778,N_9912,N_8536);
or U12779 (N_12779,N_8011,N_10407);
nand U12780 (N_12780,N_10652,N_9590);
xnor U12781 (N_12781,N_8153,N_8157);
nand U12782 (N_12782,N_8878,N_10016);
and U12783 (N_12783,N_10163,N_9036);
or U12784 (N_12784,N_10220,N_9192);
xnor U12785 (N_12785,N_10257,N_10278);
nand U12786 (N_12786,N_9591,N_11917);
or U12787 (N_12787,N_11703,N_8551);
and U12788 (N_12788,N_11772,N_10417);
nor U12789 (N_12789,N_8681,N_9258);
xnor U12790 (N_12790,N_9698,N_11601);
xor U12791 (N_12791,N_9104,N_10985);
or U12792 (N_12792,N_10498,N_9424);
nand U12793 (N_12793,N_10961,N_9534);
xor U12794 (N_12794,N_10067,N_11349);
xnor U12795 (N_12795,N_10832,N_11032);
nor U12796 (N_12796,N_10033,N_10960);
nand U12797 (N_12797,N_8047,N_10275);
nor U12798 (N_12798,N_8063,N_11791);
or U12799 (N_12799,N_8181,N_9959);
nor U12800 (N_12800,N_9482,N_9402);
or U12801 (N_12801,N_9936,N_10815);
nand U12802 (N_12802,N_8017,N_11283);
or U12803 (N_12803,N_11553,N_8532);
and U12804 (N_12804,N_11440,N_11889);
nand U12805 (N_12805,N_8310,N_10202);
or U12806 (N_12806,N_10791,N_8413);
and U12807 (N_12807,N_8508,N_9839);
xnor U12808 (N_12808,N_9288,N_10125);
and U12809 (N_12809,N_8541,N_11761);
and U12810 (N_12810,N_11526,N_9629);
or U12811 (N_12811,N_10599,N_11093);
xnor U12812 (N_12812,N_11193,N_9098);
and U12813 (N_12813,N_11561,N_10537);
xor U12814 (N_12814,N_10413,N_8328);
and U12815 (N_12815,N_9636,N_9739);
nor U12816 (N_12816,N_9419,N_9020);
and U12817 (N_12817,N_9240,N_8468);
xnor U12818 (N_12818,N_9093,N_11201);
xor U12819 (N_12819,N_8932,N_9816);
and U12820 (N_12820,N_11676,N_11022);
or U12821 (N_12821,N_11286,N_11675);
xor U12822 (N_12822,N_9249,N_11370);
xnor U12823 (N_12823,N_10370,N_10069);
or U12824 (N_12824,N_9336,N_10735);
and U12825 (N_12825,N_10262,N_8530);
and U12826 (N_12826,N_8803,N_10451);
and U12827 (N_12827,N_11225,N_11118);
and U12828 (N_12828,N_9131,N_8168);
or U12829 (N_12829,N_9149,N_11109);
nor U12830 (N_12830,N_9022,N_9312);
and U12831 (N_12831,N_10559,N_9023);
and U12832 (N_12832,N_8442,N_11877);
nor U12833 (N_12833,N_11898,N_11645);
or U12834 (N_12834,N_8326,N_8931);
xnor U12835 (N_12835,N_11227,N_9211);
and U12836 (N_12836,N_11801,N_8175);
nor U12837 (N_12837,N_10258,N_8254);
or U12838 (N_12838,N_10344,N_11456);
and U12839 (N_12839,N_9339,N_9388);
and U12840 (N_12840,N_8712,N_8581);
and U12841 (N_12841,N_10690,N_11946);
or U12842 (N_12842,N_8475,N_9139);
or U12843 (N_12843,N_10272,N_11290);
xor U12844 (N_12844,N_11572,N_10463);
nor U12845 (N_12845,N_11087,N_11587);
nand U12846 (N_12846,N_11640,N_8346);
nor U12847 (N_12847,N_8010,N_11302);
nand U12848 (N_12848,N_9963,N_11211);
and U12849 (N_12849,N_9931,N_9516);
and U12850 (N_12850,N_11191,N_11042);
nand U12851 (N_12851,N_11213,N_9677);
xnor U12852 (N_12852,N_11702,N_10921);
xnor U12853 (N_12853,N_11216,N_8405);
nand U12854 (N_12854,N_10039,N_10896);
and U12855 (N_12855,N_10871,N_8837);
and U12856 (N_12856,N_11805,N_11940);
nand U12857 (N_12857,N_8030,N_11934);
nand U12858 (N_12858,N_10780,N_10545);
or U12859 (N_12859,N_8824,N_11090);
or U12860 (N_12860,N_11457,N_8509);
nand U12861 (N_12861,N_9763,N_10508);
or U12862 (N_12862,N_10894,N_11085);
and U12863 (N_12863,N_8548,N_8799);
and U12864 (N_12864,N_9045,N_11628);
or U12865 (N_12865,N_10676,N_9107);
or U12866 (N_12866,N_8550,N_11856);
nor U12867 (N_12867,N_8361,N_11091);
nor U12868 (N_12868,N_10595,N_10570);
xnor U12869 (N_12869,N_9491,N_10139);
nor U12870 (N_12870,N_10338,N_10367);
and U12871 (N_12871,N_8320,N_9751);
nor U12872 (N_12872,N_10959,N_10177);
nand U12873 (N_12873,N_10457,N_9369);
xnor U12874 (N_12874,N_9156,N_11851);
or U12875 (N_12875,N_9779,N_9224);
xor U12876 (N_12876,N_9735,N_11890);
xor U12877 (N_12877,N_11974,N_9799);
xor U12878 (N_12878,N_11749,N_8747);
nand U12879 (N_12879,N_9261,N_8342);
xor U12880 (N_12880,N_9435,N_10312);
and U12881 (N_12881,N_10742,N_9477);
nand U12882 (N_12882,N_8929,N_11635);
xor U12883 (N_12883,N_11131,N_9955);
xnor U12884 (N_12884,N_9179,N_10030);
nand U12885 (N_12885,N_11151,N_10854);
nand U12886 (N_12886,N_9914,N_8106);
xor U12887 (N_12887,N_8757,N_10724);
nor U12888 (N_12888,N_8183,N_11061);
xor U12889 (N_12889,N_9948,N_9904);
nor U12890 (N_12890,N_9947,N_9738);
xnor U12891 (N_12891,N_10373,N_8907);
nor U12892 (N_12892,N_10555,N_8200);
and U12893 (N_12893,N_10930,N_11502);
xor U12894 (N_12894,N_9756,N_8906);
xor U12895 (N_12895,N_11071,N_8355);
nand U12896 (N_12896,N_10445,N_9385);
nand U12897 (N_12897,N_9489,N_8854);
and U12898 (N_12898,N_8846,N_10729);
or U12899 (N_12899,N_11817,N_10919);
nand U12900 (N_12900,N_10122,N_11450);
nand U12901 (N_12901,N_11734,N_9941);
nand U12902 (N_12902,N_10082,N_8908);
or U12903 (N_12903,N_10629,N_10184);
and U12904 (N_12904,N_11865,N_10157);
nor U12905 (N_12905,N_9244,N_8583);
nor U12906 (N_12906,N_11821,N_10751);
nand U12907 (N_12907,N_8847,N_10186);
and U12908 (N_12908,N_9510,N_10827);
nand U12909 (N_12909,N_9463,N_10816);
nor U12910 (N_12910,N_9078,N_11303);
nor U12911 (N_12911,N_8781,N_10734);
and U12912 (N_12912,N_8376,N_9723);
xnor U12913 (N_12913,N_9187,N_9209);
nor U12914 (N_12914,N_10710,N_11121);
and U12915 (N_12915,N_9111,N_10529);
xor U12916 (N_12916,N_10236,N_9432);
nand U12917 (N_12917,N_8235,N_9468);
nand U12918 (N_12918,N_9049,N_11958);
nand U12919 (N_12919,N_11585,N_11168);
or U12920 (N_12920,N_9519,N_11143);
xnor U12921 (N_12921,N_8273,N_11169);
and U12922 (N_12922,N_8830,N_11308);
and U12923 (N_12923,N_9447,N_11595);
xnor U12924 (N_12924,N_9396,N_10354);
or U12925 (N_12925,N_9217,N_11926);
nand U12926 (N_12926,N_8278,N_8001);
nand U12927 (N_12927,N_9462,N_9160);
xnor U12928 (N_12928,N_9497,N_11882);
nand U12929 (N_12929,N_8912,N_11875);
and U12930 (N_12930,N_8894,N_9683);
or U12931 (N_12931,N_10853,N_8668);
or U12932 (N_12932,N_9417,N_11347);
or U12933 (N_12933,N_9193,N_9949);
nor U12934 (N_12934,N_10266,N_8020);
or U12935 (N_12935,N_8577,N_10060);
nor U12936 (N_12936,N_11701,N_8148);
nor U12937 (N_12937,N_10678,N_9133);
nor U12938 (N_12938,N_11565,N_10697);
nand U12939 (N_12939,N_9837,N_8283);
nand U12940 (N_12940,N_11381,N_10436);
nor U12941 (N_12941,N_10025,N_8899);
xor U12942 (N_12942,N_10477,N_9715);
xor U12943 (N_12943,N_11353,N_8914);
nand U12944 (N_12944,N_8947,N_11919);
nand U12945 (N_12945,N_8481,N_8816);
nor U12946 (N_12946,N_8788,N_10754);
nor U12947 (N_12947,N_9297,N_9890);
xor U12948 (N_12948,N_8072,N_9814);
and U12949 (N_12949,N_8499,N_8553);
or U12950 (N_12950,N_11757,N_10006);
and U12951 (N_12951,N_8525,N_8297);
or U12952 (N_12952,N_8858,N_8744);
or U12953 (N_12953,N_11224,N_9819);
xor U12954 (N_12954,N_11831,N_8377);
nand U12955 (N_12955,N_11970,N_11494);
xor U12956 (N_12956,N_9588,N_11657);
xnor U12957 (N_12957,N_9676,N_10408);
nand U12958 (N_12958,N_8136,N_8460);
nor U12959 (N_12959,N_9058,N_10129);
nor U12960 (N_12960,N_10765,N_9188);
xor U12961 (N_12961,N_8143,N_8056);
nor U12962 (N_12962,N_11650,N_10265);
xnor U12963 (N_12963,N_8851,N_9115);
nor U12964 (N_12964,N_10024,N_10723);
nand U12965 (N_12965,N_10848,N_9262);
nand U12966 (N_12966,N_11321,N_11656);
nand U12967 (N_12967,N_10674,N_9654);
xnor U12968 (N_12968,N_8811,N_8686);
nand U12969 (N_12969,N_10514,N_9998);
and U12970 (N_12970,N_10226,N_10201);
and U12971 (N_12971,N_10366,N_8674);
xnor U12972 (N_12972,N_8697,N_10131);
xnor U12973 (N_12973,N_11780,N_10171);
or U12974 (N_12974,N_8665,N_10671);
xnor U12975 (N_12975,N_10231,N_11255);
xnor U12976 (N_12976,N_11622,N_8443);
xnor U12977 (N_12977,N_11011,N_11773);
or U12978 (N_12978,N_9293,N_8859);
nor U12979 (N_12979,N_9790,N_10193);
xor U12980 (N_12980,N_10402,N_8558);
nor U12981 (N_12981,N_10250,N_11669);
or U12982 (N_12982,N_8448,N_10982);
nor U12983 (N_12983,N_8220,N_8771);
nand U12984 (N_12984,N_9467,N_10100);
nor U12985 (N_12985,N_8367,N_8256);
and U12986 (N_12986,N_10218,N_11101);
and U12987 (N_12987,N_11607,N_10770);
nor U12988 (N_12988,N_10539,N_8048);
nor U12989 (N_12989,N_8954,N_11699);
or U12990 (N_12990,N_11275,N_10490);
and U12991 (N_12991,N_11070,N_8709);
xor U12992 (N_12992,N_10805,N_9784);
or U12993 (N_12993,N_9509,N_10698);
or U12994 (N_12994,N_11043,N_9464);
nand U12995 (N_12995,N_9167,N_9212);
nor U12996 (N_12996,N_10875,N_10431);
nor U12997 (N_12997,N_8972,N_9281);
xor U12998 (N_12998,N_8267,N_11445);
nor U12999 (N_12999,N_8325,N_9712);
nand U13000 (N_13000,N_10472,N_10571);
and U13001 (N_13001,N_9239,N_8015);
nor U13002 (N_13002,N_8716,N_9974);
nor U13003 (N_13003,N_11954,N_11913);
and U13004 (N_13004,N_9691,N_11748);
or U13005 (N_13005,N_8432,N_8707);
nor U13006 (N_13006,N_8434,N_8006);
xor U13007 (N_13007,N_8119,N_10818);
xor U13008 (N_13008,N_8433,N_8875);
or U13009 (N_13009,N_11350,N_8856);
and U13010 (N_13010,N_10014,N_11452);
nor U13011 (N_13011,N_11869,N_9838);
or U13012 (N_13012,N_9046,N_8350);
or U13013 (N_13013,N_8428,N_9538);
nand U13014 (N_13014,N_11874,N_8633);
nor U13015 (N_13015,N_9803,N_11648);
or U13016 (N_13016,N_9517,N_9669);
xor U13017 (N_13017,N_8733,N_9741);
xnor U13018 (N_13018,N_11218,N_11931);
nor U13019 (N_13019,N_9473,N_9373);
nor U13020 (N_13020,N_10209,N_9141);
xnor U13021 (N_13021,N_10601,N_9069);
or U13022 (N_13022,N_8629,N_8349);
nor U13023 (N_13023,N_8518,N_11663);
and U13024 (N_13024,N_11998,N_9498);
nor U13025 (N_13025,N_10981,N_11612);
nand U13026 (N_13026,N_9292,N_11119);
nand U13027 (N_13027,N_10944,N_10849);
or U13028 (N_13028,N_10263,N_11955);
and U13029 (N_13029,N_11708,N_9755);
nor U13030 (N_13030,N_8387,N_9655);
or U13031 (N_13031,N_9340,N_9847);
nor U13032 (N_13032,N_9727,N_8100);
nor U13033 (N_13033,N_10189,N_11488);
xor U13034 (N_13034,N_11840,N_9673);
and U13035 (N_13035,N_8774,N_11113);
and U13036 (N_13036,N_10511,N_9439);
or U13037 (N_13037,N_10953,N_10154);
xnor U13038 (N_13038,N_9114,N_8540);
and U13039 (N_13039,N_10844,N_11233);
and U13040 (N_13040,N_10762,N_8049);
xnor U13041 (N_13041,N_9206,N_11528);
and U13042 (N_13042,N_11419,N_10812);
and U13043 (N_13043,N_8892,N_11632);
xnor U13044 (N_13044,N_9146,N_8316);
or U13045 (N_13045,N_8986,N_11520);
and U13046 (N_13046,N_8077,N_11710);
or U13047 (N_13047,N_9153,N_11833);
and U13048 (N_13048,N_9846,N_10782);
nor U13049 (N_13049,N_11532,N_10309);
nor U13050 (N_13050,N_8538,N_10940);
xor U13051 (N_13051,N_8237,N_8296);
and U13052 (N_13052,N_9815,N_9317);
and U13053 (N_13053,N_10828,N_9213);
nand U13054 (N_13054,N_8226,N_10517);
nor U13055 (N_13055,N_10423,N_11925);
or U13056 (N_13056,N_10736,N_8426);
nand U13057 (N_13057,N_8114,N_8567);
or U13058 (N_13058,N_11299,N_8647);
nor U13059 (N_13059,N_9183,N_8033);
nand U13060 (N_13060,N_10215,N_9342);
nor U13061 (N_13061,N_8845,N_11293);
xnor U13062 (N_13062,N_8760,N_9478);
nand U13063 (N_13063,N_9913,N_9505);
and U13064 (N_13064,N_8177,N_9445);
and U13065 (N_13065,N_11698,N_11827);
nand U13066 (N_13066,N_11982,N_9372);
and U13067 (N_13067,N_11559,N_9151);
or U13068 (N_13068,N_11479,N_11542);
nand U13069 (N_13069,N_9597,N_8028);
and U13070 (N_13070,N_11726,N_11571);
nand U13071 (N_13071,N_11019,N_8542);
and U13072 (N_13072,N_9893,N_8389);
xor U13073 (N_13073,N_8657,N_10361);
nor U13074 (N_13074,N_8823,N_9330);
or U13075 (N_13075,N_9625,N_8813);
and U13076 (N_13076,N_10918,N_10386);
nor U13077 (N_13077,N_11523,N_9007);
or U13078 (N_13078,N_11767,N_10949);
nor U13079 (N_13079,N_9895,N_8849);
or U13080 (N_13080,N_11363,N_10228);
nand U13081 (N_13081,N_9675,N_10185);
or U13082 (N_13082,N_11401,N_8040);
xnor U13083 (N_13083,N_11424,N_8374);
nand U13084 (N_13084,N_10043,N_8561);
or U13085 (N_13085,N_8618,N_9570);
nor U13086 (N_13086,N_11626,N_9688);
or U13087 (N_13087,N_9178,N_10932);
or U13088 (N_13088,N_9398,N_9129);
nor U13089 (N_13089,N_11687,N_11441);
nand U13090 (N_13090,N_8279,N_11316);
nor U13091 (N_13091,N_9071,N_9861);
or U13092 (N_13092,N_10009,N_11863);
nor U13093 (N_13093,N_9006,N_11125);
nand U13094 (N_13094,N_8949,N_10311);
and U13095 (N_13095,N_10788,N_8545);
nand U13096 (N_13096,N_11260,N_10277);
or U13097 (N_13097,N_10503,N_9408);
or U13098 (N_13098,N_8453,N_9018);
nor U13099 (N_13099,N_10739,N_11144);
nand U13100 (N_13100,N_10234,N_9764);
or U13101 (N_13101,N_11870,N_9783);
or U13102 (N_13102,N_8738,N_9685);
xnor U13103 (N_13103,N_9070,N_11853);
xnor U13104 (N_13104,N_8236,N_10001);
and U13105 (N_13105,N_9148,N_10070);
xnor U13106 (N_13106,N_9872,N_8396);
nand U13107 (N_13107,N_9649,N_9126);
nand U13108 (N_13108,N_11335,N_11313);
nand U13109 (N_13109,N_11957,N_11510);
nor U13110 (N_13110,N_10623,N_9907);
or U13111 (N_13111,N_11688,N_11577);
nor U13112 (N_13112,N_10480,N_11910);
nor U13113 (N_13113,N_9699,N_10983);
nand U13114 (N_13114,N_11709,N_11478);
xnor U13115 (N_13115,N_10074,N_9483);
nor U13116 (N_13116,N_9762,N_8423);
or U13117 (N_13117,N_11183,N_9854);
or U13118 (N_13118,N_11341,N_8245);
xor U13119 (N_13119,N_8700,N_10099);
nor U13120 (N_13120,N_11549,N_8902);
or U13121 (N_13121,N_11020,N_11923);
and U13122 (N_13122,N_10863,N_10285);
xnor U13123 (N_13123,N_10128,N_10705);
nand U13124 (N_13124,N_11398,N_9382);
xor U13125 (N_13125,N_8362,N_11342);
or U13126 (N_13126,N_9029,N_11287);
xor U13127 (N_13127,N_10290,N_9850);
or U13128 (N_13128,N_10622,N_10384);
nor U13129 (N_13129,N_11540,N_10681);
nand U13130 (N_13130,N_8104,N_9323);
nand U13131 (N_13131,N_11284,N_8230);
and U13132 (N_13132,N_11311,N_10563);
nor U13133 (N_13133,N_8755,N_8419);
nand U13134 (N_13134,N_10397,N_9674);
nor U13135 (N_13135,N_9726,N_10446);
and U13136 (N_13136,N_11069,N_9651);
nor U13137 (N_13137,N_8592,N_11503);
nor U13138 (N_13138,N_10320,N_8705);
nor U13139 (N_13139,N_11495,N_11394);
or U13140 (N_13140,N_11166,N_9195);
nor U13141 (N_13141,N_10906,N_10012);
nor U13142 (N_13142,N_8424,N_9349);
and U13143 (N_13143,N_8531,N_9418);
xor U13144 (N_13144,N_8190,N_8814);
or U13145 (N_13145,N_10994,N_8016);
nor U13146 (N_13146,N_10063,N_8863);
xnor U13147 (N_13147,N_9833,N_10840);
xnor U13148 (N_13148,N_10115,N_10252);
xor U13149 (N_13149,N_10368,N_8562);
and U13150 (N_13150,N_9495,N_8137);
and U13151 (N_13151,N_9315,N_11501);
and U13152 (N_13152,N_10279,N_10837);
xor U13153 (N_13153,N_10990,N_10465);
nand U13154 (N_13154,N_9919,N_9961);
and U13155 (N_13155,N_9990,N_8708);
xnor U13156 (N_13156,N_11206,N_11100);
and U13157 (N_13157,N_11558,N_11718);
nand U13158 (N_13158,N_10411,N_9503);
nand U13159 (N_13159,N_9479,N_9679);
nand U13160 (N_13160,N_8966,N_9980);
and U13161 (N_13161,N_9175,N_11944);
and U13162 (N_13162,N_10509,N_10481);
nand U13163 (N_13163,N_11830,N_8004);
nor U13164 (N_13164,N_9019,N_9522);
and U13165 (N_13165,N_8625,N_11593);
nand U13166 (N_13166,N_8903,N_11855);
or U13167 (N_13167,N_8133,N_11146);
or U13168 (N_13168,N_11730,N_11388);
xor U13169 (N_13169,N_9812,N_9290);
nand U13170 (N_13170,N_11667,N_8260);
or U13171 (N_13171,N_10802,N_11058);
or U13172 (N_13172,N_10666,N_9533);
xnor U13173 (N_13173,N_8117,N_11854);
nand U13174 (N_13174,N_9021,N_10699);
nor U13175 (N_13175,N_9733,N_8262);
nand U13176 (N_13176,N_9554,N_8928);
nand U13177 (N_13177,N_11434,N_10592);
or U13178 (N_13178,N_9055,N_9494);
nor U13179 (N_13179,N_10581,N_11264);
nor U13180 (N_13180,N_11390,N_8777);
and U13181 (N_13181,N_9573,N_8076);
nand U13182 (N_13182,N_8171,N_9829);
xor U13183 (N_13183,N_11580,N_10606);
nand U13184 (N_13184,N_10119,N_9926);
nand U13185 (N_13185,N_9243,N_11513);
or U13186 (N_13186,N_9717,N_11785);
nand U13187 (N_13187,N_8164,N_8616);
or U13188 (N_13188,N_9460,N_8765);
and U13189 (N_13189,N_10966,N_11912);
xor U13190 (N_13190,N_11673,N_9256);
nand U13191 (N_13191,N_9367,N_9325);
and U13192 (N_13192,N_9871,N_10395);
xnor U13193 (N_13193,N_10420,N_8023);
nand U13194 (N_13194,N_10835,N_8252);
nand U13195 (N_13195,N_9911,N_10456);
nor U13196 (N_13196,N_11339,N_10813);
nand U13197 (N_13197,N_9091,N_8913);
or U13198 (N_13198,N_10461,N_9366);
xor U13199 (N_13199,N_8455,N_9004);
nand U13200 (N_13200,N_11096,N_10722);
nor U13201 (N_13201,N_10425,N_8401);
or U13202 (N_13202,N_11037,N_9672);
and U13203 (N_13203,N_9927,N_8126);
xor U13204 (N_13204,N_10334,N_9453);
nand U13205 (N_13205,N_8937,N_8204);
nand U13206 (N_13206,N_9450,N_10295);
nor U13207 (N_13207,N_10636,N_11142);
or U13208 (N_13208,N_11808,N_8880);
nor U13209 (N_13209,N_8767,N_8808);
or U13210 (N_13210,N_11603,N_8379);
xnor U13211 (N_13211,N_9930,N_8009);
and U13212 (N_13212,N_10866,N_10515);
and U13213 (N_13213,N_11864,N_8437);
and U13214 (N_13214,N_9363,N_8058);
and U13215 (N_13215,N_9102,N_11765);
nand U13216 (N_13216,N_8506,N_8087);
and U13217 (N_13217,N_11387,N_10017);
or U13218 (N_13218,N_11496,N_10684);
xnor U13219 (N_13219,N_9881,N_8783);
or U13220 (N_13220,N_9043,N_9067);
xor U13221 (N_13221,N_8142,N_8501);
nand U13222 (N_13222,N_9638,N_10947);
nor U13223 (N_13223,N_9729,N_11052);
and U13224 (N_13224,N_10996,N_10484);
nor U13225 (N_13225,N_11155,N_11008);
xnor U13226 (N_13226,N_11466,N_10390);
xnor U13227 (N_13227,N_8641,N_8386);
nor U13228 (N_13228,N_9906,N_8789);
and U13229 (N_13229,N_8768,N_11246);
nor U13230 (N_13230,N_11860,N_10330);
nand U13231 (N_13231,N_8307,N_8673);
or U13232 (N_13232,N_11076,N_9544);
and U13233 (N_13233,N_11021,N_8839);
and U13234 (N_13234,N_11040,N_8378);
and U13235 (N_13235,N_10586,N_10346);
nor U13236 (N_13236,N_11200,N_10884);
xor U13237 (N_13237,N_11395,N_11547);
xnor U13238 (N_13238,N_10308,N_9652);
nand U13239 (N_13239,N_9737,N_9232);
xor U13240 (N_13240,N_9765,N_9144);
nor U13241 (N_13241,N_10798,N_9624);
nand U13242 (N_13242,N_11297,N_10912);
or U13243 (N_13243,N_9060,N_9079);
and U13244 (N_13244,N_9909,N_11389);
nor U13245 (N_13245,N_9531,N_11642);
nand U13246 (N_13246,N_10011,N_8392);
xor U13247 (N_13247,N_8870,N_11776);
and U13248 (N_13248,N_9099,N_11914);
nor U13249 (N_13249,N_9992,N_11802);
nor U13250 (N_13250,N_8027,N_9270);
xor U13251 (N_13251,N_10806,N_9757);
or U13252 (N_13252,N_8593,N_8280);
or U13253 (N_13253,N_8211,N_10686);
or U13254 (N_13254,N_8384,N_9132);
nor U13255 (N_13255,N_9375,N_8025);
or U13256 (N_13256,N_8352,N_8721);
and U13257 (N_13257,N_8082,N_8521);
xor U13258 (N_13258,N_10286,N_10118);
xor U13259 (N_13259,N_11695,N_11715);
nand U13260 (N_13260,N_11929,N_8271);
nor U13261 (N_13261,N_11140,N_8772);
and U13262 (N_13262,N_9887,N_10095);
nor U13263 (N_13263,N_9170,N_11819);
and U13264 (N_13264,N_10141,N_8557);
or U13265 (N_13265,N_10444,N_9461);
or U13266 (N_13266,N_11279,N_9703);
xnor U13267 (N_13267,N_9878,N_10349);
xnor U13268 (N_13268,N_9820,N_8578);
nor U13269 (N_13269,N_10040,N_8628);
nand U13270 (N_13270,N_10861,N_11123);
nor U13271 (N_13271,N_8315,N_11770);
nor U13272 (N_13272,N_9327,N_10369);
nand U13273 (N_13273,N_10948,N_8679);
or U13274 (N_13274,N_10637,N_10168);
nor U13275 (N_13275,N_8391,N_10358);
or U13276 (N_13276,N_10967,N_9774);
or U13277 (N_13277,N_10560,N_9800);
and U13278 (N_13278,N_11682,N_9627);
xnor U13279 (N_13279,N_10913,N_10808);
nor U13280 (N_13280,N_10487,N_9236);
or U13281 (N_13281,N_8825,N_11804);
nor U13282 (N_13282,N_9958,N_10158);
or U13283 (N_13283,N_8872,N_9444);
xor U13284 (N_13284,N_10748,N_10090);
xnor U13285 (N_13285,N_10989,N_10688);
xor U13286 (N_13286,N_10669,N_10303);
or U13287 (N_13287,N_11965,N_8882);
or U13288 (N_13288,N_8660,N_8763);
nor U13289 (N_13289,N_10015,N_10708);
nand U13290 (N_13290,N_10593,N_8128);
or U13291 (N_13291,N_9734,N_11795);
or U13292 (N_13292,N_10449,N_9298);
and U13293 (N_13293,N_10618,N_9802);
nor U13294 (N_13294,N_10356,N_10612);
nor U13295 (N_13295,N_8671,N_11177);
xnor U13296 (N_13296,N_9641,N_10602);
xor U13297 (N_13297,N_11918,N_9371);
xor U13298 (N_13298,N_9709,N_10811);
or U13299 (N_13299,N_10712,N_11357);
xor U13300 (N_13300,N_10310,N_9707);
or U13301 (N_13301,N_11188,N_10557);
nand U13302 (N_13302,N_8848,N_8649);
nand U13303 (N_13303,N_9830,N_11716);
nor U13304 (N_13304,N_11266,N_9063);
or U13305 (N_13305,N_8751,N_9523);
nand U13306 (N_13306,N_8012,N_11814);
and U13307 (N_13307,N_11741,N_10530);
xnor U13308 (N_13308,N_8507,N_9476);
and U13309 (N_13309,N_10087,N_9177);
xnor U13310 (N_13310,N_10980,N_10925);
nand U13311 (N_13311,N_9805,N_11126);
or U13312 (N_13312,N_9760,N_8299);
nand U13313 (N_13313,N_11310,N_11277);
nand U13314 (N_13314,N_8750,N_9608);
nor U13315 (N_13315,N_11490,N_9659);
nor U13316 (N_13316,N_11690,N_9154);
or U13317 (N_13317,N_10406,N_8888);
xor U13318 (N_13318,N_11990,N_8094);
nor U13319 (N_13319,N_9433,N_10558);
and U13320 (N_13320,N_10094,N_11249);
or U13321 (N_13321,N_10261,N_8951);
or U13322 (N_13322,N_8821,N_10379);
or U13323 (N_13323,N_10291,N_10326);
and U13324 (N_13324,N_10943,N_8272);
xnor U13325 (N_13325,N_9804,N_9265);
or U13326 (N_13326,N_11056,N_10519);
and U13327 (N_13327,N_8261,N_10952);
nor U13328 (N_13328,N_9121,N_10149);
nand U13329 (N_13329,N_9300,N_8524);
and U13330 (N_13330,N_11185,N_11623);
nor U13331 (N_13331,N_8662,N_11781);
xnor U13332 (N_13332,N_10156,N_8053);
and U13333 (N_13333,N_9318,N_9040);
and U13334 (N_13334,N_9556,N_9826);
xnor U13335 (N_13335,N_8690,N_9301);
and U13336 (N_13336,N_10915,N_10633);
and U13337 (N_13337,N_11409,N_11811);
and U13338 (N_13338,N_11986,N_11130);
and U13339 (N_13339,N_11516,N_9073);
nor U13340 (N_13340,N_11861,N_9882);
and U13341 (N_13341,N_11966,N_10744);
or U13342 (N_13342,N_9842,N_9176);
and U13343 (N_13343,N_11002,N_8034);
nor U13344 (N_13344,N_10325,N_9640);
and U13345 (N_13345,N_11473,N_10253);
xor U13346 (N_13346,N_10190,N_8318);
nand U13347 (N_13347,N_11049,N_9835);
or U13348 (N_13348,N_8120,N_9241);
or U13349 (N_13349,N_9870,N_11691);
nand U13350 (N_13350,N_11268,N_11459);
and U13351 (N_13351,N_11738,N_8831);
and U13352 (N_13352,N_10680,N_11160);
xnor U13353 (N_13353,N_8398,N_11943);
xnor U13354 (N_13354,N_10850,N_9421);
or U13355 (N_13355,N_10003,N_9470);
nor U13356 (N_13356,N_11908,N_11764);
xnor U13357 (N_13357,N_8132,N_11095);
xor U13358 (N_13358,N_10455,N_9542);
nor U13359 (N_13359,N_9234,N_8277);
and U13360 (N_13360,N_9650,N_10044);
nor U13361 (N_13361,N_10576,N_8952);
or U13362 (N_13362,N_11883,N_8414);
xnor U13363 (N_13363,N_9977,N_10270);
nand U13364 (N_13364,N_9989,N_10353);
nand U13365 (N_13365,N_11813,N_8155);
or U13366 (N_13366,N_8969,N_8224);
and U13367 (N_13367,N_8493,N_10670);
or U13368 (N_13368,N_10357,N_8873);
or U13369 (N_13369,N_8294,N_8385);
or U13370 (N_13370,N_8057,N_10188);
nand U13371 (N_13371,N_9090,N_11462);
and U13372 (N_13372,N_8441,N_11128);
xor U13373 (N_13373,N_8130,N_11480);
nor U13374 (N_13374,N_10273,N_11594);
nand U13375 (N_13375,N_10035,N_9284);
or U13376 (N_13376,N_8146,N_11322);
or U13377 (N_13377,N_8898,N_11746);
nor U13378 (N_13378,N_8529,N_11138);
xnor U13379 (N_13379,N_8998,N_9005);
nand U13380 (N_13380,N_8764,N_8324);
and U13381 (N_13381,N_11427,N_10824);
and U13382 (N_13382,N_9041,N_9401);
and U13383 (N_13383,N_9014,N_9614);
nand U13384 (N_13384,N_8940,N_8775);
or U13385 (N_13385,N_9642,N_9057);
xnor U13386 (N_13386,N_9220,N_10862);
and U13387 (N_13387,N_9310,N_8289);
xor U13388 (N_13388,N_8044,N_10079);
xor U13389 (N_13389,N_8680,N_8429);
nor U13390 (N_13390,N_11905,N_8138);
nor U13391 (N_13391,N_9266,N_10199);
or U13392 (N_13392,N_9032,N_9180);
nor U13393 (N_13393,N_10758,N_10954);
nand U13394 (N_13394,N_10475,N_10972);
nand U13395 (N_13395,N_9053,N_10917);
or U13396 (N_13396,N_11590,N_11442);
nand U13397 (N_13397,N_9452,N_8115);
nand U13398 (N_13398,N_8095,N_8043);
or U13399 (N_13399,N_10450,N_10880);
or U13400 (N_13400,N_11554,N_9271);
xnor U13401 (N_13401,N_10756,N_11292);
nor U13402 (N_13402,N_9724,N_10726);
nand U13403 (N_13403,N_11569,N_11222);
nor U13404 (N_13404,N_8691,N_8809);
or U13405 (N_13405,N_8081,N_11759);
nor U13406 (N_13406,N_10013,N_10415);
and U13407 (N_13407,N_9515,N_11762);
xnor U13408 (N_13408,N_10730,N_11655);
nor U13409 (N_13409,N_10347,N_9143);
nor U13410 (N_13410,N_11013,N_8580);
xor U13411 (N_13411,N_10439,N_10998);
or U13412 (N_13412,N_8054,N_9524);
nand U13413 (N_13413,N_11659,N_10893);
and U13414 (N_13414,N_9008,N_9487);
and U13415 (N_13415,N_11658,N_8866);
nor U13416 (N_13416,N_9161,N_8572);
nor U13417 (N_13417,N_8344,N_9684);
or U13418 (N_13418,N_9097,N_9639);
nor U13419 (N_13419,N_11129,N_8643);
nor U13420 (N_13420,N_9653,N_8909);
nor U13421 (N_13421,N_9155,N_10176);
or U13422 (N_13422,N_10049,N_9222);
nand U13423 (N_13423,N_11493,N_8213);
and U13424 (N_13424,N_10789,N_11256);
or U13425 (N_13425,N_10393,N_11007);
xor U13426 (N_13426,N_10645,N_11444);
nand U13427 (N_13427,N_8975,N_11891);
xor U13428 (N_13428,N_9568,N_10526);
or U13429 (N_13429,N_8007,N_11447);
or U13430 (N_13430,N_9034,N_10978);
or U13431 (N_13431,N_9199,N_11768);
and U13432 (N_13432,N_11285,N_9817);
nand U13433 (N_13433,N_10002,N_8537);
nor U13434 (N_13434,N_11961,N_9607);
and U13435 (N_13435,N_10062,N_8203);
or U13436 (N_13436,N_10343,N_10433);
xor U13437 (N_13437,N_9255,N_11186);
nand U13438 (N_13438,N_11818,N_8107);
nor U13439 (N_13439,N_11697,N_9009);
nor U13440 (N_13440,N_11584,N_11301);
and U13441 (N_13441,N_9903,N_8836);
nand U13442 (N_13442,N_8022,N_9514);
and U13443 (N_13443,N_9567,N_9268);
xor U13444 (N_13444,N_9196,N_8644);
nand U13445 (N_13445,N_9471,N_10860);
nand U13446 (N_13446,N_8131,N_10775);
nor U13447 (N_13447,N_11325,N_10010);
or U13448 (N_13448,N_8604,N_9412);
nor U13449 (N_13449,N_11404,N_11062);
xor U13450 (N_13450,N_11251,N_11212);
nand U13451 (N_13451,N_9404,N_9488);
nand U13452 (N_13452,N_9891,N_10136);
and U13453 (N_13453,N_8792,N_8588);
or U13454 (N_13454,N_8867,N_11573);
and U13455 (N_13455,N_8619,N_11048);
nor U13456 (N_13456,N_9075,N_10564);
and U13457 (N_13457,N_8323,N_8994);
nor U13458 (N_13458,N_11024,N_8724);
xnor U13459 (N_13459,N_9551,N_8612);
or U13460 (N_13460,N_9454,N_10630);
or U13461 (N_13461,N_10732,N_9202);
or U13462 (N_13462,N_9583,N_8306);
nand U13463 (N_13463,N_10955,N_8539);
xor U13464 (N_13464,N_9718,N_9777);
and U13465 (N_13465,N_8955,N_9440);
xor U13466 (N_13466,N_10143,N_11269);
nor U13467 (N_13467,N_11406,N_10287);
and U13468 (N_13468,N_10052,N_9983);
nor U13469 (N_13469,N_10575,N_8877);
nand U13470 (N_13470,N_8871,N_8579);
nor U13471 (N_13471,N_10453,N_10521);
nor U13472 (N_13472,N_9954,N_10939);
nand U13473 (N_13473,N_11849,N_10108);
and U13474 (N_13474,N_10216,N_11605);
xnor U13475 (N_13475,N_8599,N_8608);
nand U13476 (N_13476,N_11616,N_11636);
or U13477 (N_13477,N_9348,N_8640);
and U13478 (N_13478,N_8300,N_11065);
or U13479 (N_13479,N_8786,N_10476);
nand U13480 (N_13480,N_9173,N_9225);
xor U13481 (N_13481,N_9257,N_11706);
nor U13482 (N_13482,N_10541,N_11307);
and U13483 (N_13483,N_11106,N_10159);
and U13484 (N_13484,N_9701,N_8351);
or U13485 (N_13485,N_8861,N_8270);
and U13486 (N_13486,N_10879,N_11959);
and U13487 (N_13487,N_10797,N_9242);
and U13488 (N_13488,N_8381,N_10037);
nand U13489 (N_13489,N_9957,N_8956);
nor U13490 (N_13490,N_11807,N_11082);
xnor U13491 (N_13491,N_10941,N_8546);
nand U13492 (N_13492,N_9582,N_10975);
and U13493 (N_13493,N_11714,N_11866);
xnor U13494 (N_13494,N_11992,N_8962);
or U13495 (N_13495,N_11809,N_10135);
xor U13496 (N_13496,N_10225,N_8239);
nand U13497 (N_13497,N_8464,N_9560);
xnor U13498 (N_13498,N_10242,N_9671);
nand U13499 (N_13499,N_11475,N_8620);
xor U13500 (N_13500,N_11241,N_11454);
nor U13501 (N_13501,N_11499,N_11900);
or U13502 (N_13502,N_10933,N_9758);
and U13503 (N_13503,N_9165,N_10364);
and U13504 (N_13504,N_8079,N_10187);
nand U13505 (N_13505,N_10362,N_9780);
and U13506 (N_13506,N_8645,N_10169);
nand U13507 (N_13507,N_10785,N_9943);
nand U13508 (N_13508,N_9973,N_9428);
and U13509 (N_13509,N_8511,N_9048);
nand U13510 (N_13510,N_8276,N_10432);
nand U13511 (N_13511,N_8163,N_11378);
nor U13512 (N_13512,N_11937,N_8188);
xnor U13513 (N_13513,N_8229,N_8210);
nand U13514 (N_13514,N_8549,N_10318);
nand U13515 (N_13515,N_11693,N_10662);
nand U13516 (N_13516,N_11250,N_9506);
nor U13517 (N_13517,N_9689,N_10023);
or U13518 (N_13518,N_8338,N_8435);
nand U13519 (N_13519,N_10339,N_9920);
nor U13520 (N_13520,N_10378,N_8976);
nor U13521 (N_13521,N_11412,N_9547);
xor U13522 (N_13522,N_10036,N_11003);
nor U13523 (N_13523,N_10799,N_8189);
nor U13524 (N_13524,N_10909,N_8594);
and U13525 (N_13525,N_9200,N_8105);
nand U13526 (N_13526,N_10731,N_10471);
xor U13527 (N_13527,N_11945,N_9716);
xnor U13528 (N_13528,N_9630,N_8573);
and U13529 (N_13529,N_10779,N_8000);
or U13530 (N_13530,N_10399,N_9572);
and U13531 (N_13531,N_11824,N_8793);
nand U13532 (N_13532,N_11991,N_9493);
or U13533 (N_13533,N_8465,N_8196);
or U13534 (N_13534,N_11240,N_8263);
and U13535 (N_13535,N_8193,N_8461);
and U13536 (N_13536,N_11458,N_10696);
nor U13537 (N_13537,N_8944,N_9350);
xor U13538 (N_13538,N_9788,N_10435);
or U13539 (N_13539,N_8896,N_10942);
nand U13540 (N_13540,N_10892,N_8302);
xor U13541 (N_13541,N_11467,N_10034);
nand U13542 (N_13542,N_10682,N_8864);
nor U13543 (N_13543,N_11327,N_9001);
xor U13544 (N_13544,N_11451,N_9615);
nand U13545 (N_13545,N_9237,N_11179);
nor U13546 (N_13546,N_10227,N_8739);
nor U13547 (N_13547,N_9466,N_10293);
nor U13548 (N_13548,N_9413,N_10546);
xor U13549 (N_13549,N_11634,N_11644);
or U13550 (N_13550,N_9549,N_8036);
or U13551 (N_13551,N_8088,N_9962);
or U13552 (N_13552,N_10664,N_10757);
and U13553 (N_13553,N_11994,N_8067);
xor U13554 (N_13554,N_11711,N_9216);
or U13555 (N_13555,N_10153,N_11543);
nand U13556 (N_13556,N_10513,N_8676);
nand U13557 (N_13557,N_8336,N_9275);
or U13558 (N_13558,N_10986,N_9357);
nand U13559 (N_13559,N_10773,N_10752);
nor U13560 (N_13560,N_8891,N_10746);
nand U13561 (N_13561,N_10140,N_9834);
or U13562 (N_13562,N_11392,N_9289);
or U13563 (N_13563,N_8737,N_8801);
xor U13564 (N_13564,N_9670,N_8585);
nand U13565 (N_13565,N_10795,N_9387);
or U13566 (N_13566,N_11104,N_11430);
nand U13567 (N_13567,N_9054,N_9600);
or U13568 (N_13568,N_9307,N_8554);
nand U13569 (N_13569,N_10488,N_9663);
nor U13570 (N_13570,N_8409,N_10888);
xor U13571 (N_13571,N_8080,N_11774);
and U13572 (N_13572,N_10792,N_8637);
nor U13573 (N_13573,N_8571,N_8059);
and U13574 (N_13574,N_10351,N_8822);
and U13575 (N_13575,N_9443,N_11678);
or U13576 (N_13576,N_11916,N_8394);
or U13577 (N_13577,N_10979,N_8843);
nor U13578 (N_13578,N_9776,N_11779);
xnor U13579 (N_13579,N_11492,N_9862);
and U13580 (N_13580,N_11514,N_8050);
nand U13581 (N_13581,N_9356,N_10665);
and U13582 (N_13582,N_8127,N_10340);
and U13583 (N_13583,N_10116,N_10577);
or U13584 (N_13584,N_11500,N_9066);
xor U13585 (N_13585,N_9828,N_11449);
or U13586 (N_13586,N_10958,N_11599);
and U13587 (N_13587,N_10038,N_9970);
nand U13588 (N_13588,N_8726,N_8828);
xnor U13589 (N_13589,N_11825,N_11219);
or U13590 (N_13590,N_10745,N_10874);
and U13591 (N_13591,N_9967,N_11596);
and U13592 (N_13592,N_11111,N_10091);
xor U13593 (N_13593,N_10831,N_9945);
or U13594 (N_13594,N_10345,N_8084);
nor U13595 (N_13595,N_10496,N_10572);
nand U13596 (N_13596,N_9233,N_9705);
xor U13597 (N_13597,N_9935,N_9697);
or U13598 (N_13598,N_10155,N_10725);
or U13599 (N_13599,N_10804,N_10627);
or U13600 (N_13600,N_10440,N_10615);
xnor U13601 (N_13601,N_11789,N_8650);
and U13602 (N_13602,N_10181,N_11112);
or U13603 (N_13603,N_9106,N_10081);
xnor U13604 (N_13604,N_11696,N_11315);
and U13605 (N_13605,N_9836,N_9438);
or U13606 (N_13606,N_11181,N_10544);
xor U13607 (N_13607,N_8479,N_9039);
and U13608 (N_13608,N_11237,N_10409);
nor U13609 (N_13609,N_8782,N_8369);
nand U13610 (N_13610,N_8784,N_8097);
or U13611 (N_13611,N_11170,N_11630);
or U13612 (N_13612,N_11329,N_10306);
and U13613 (N_13613,N_9352,N_10315);
nand U13614 (N_13614,N_8440,N_9437);
or U13615 (N_13615,N_10891,N_10718);
or U13616 (N_13616,N_11582,N_8490);
nor U13617 (N_13617,N_10591,N_10180);
or U13618 (N_13618,N_9341,N_8291);
or U13619 (N_13619,N_9125,N_11092);
or U13620 (N_13620,N_10784,N_10621);
nand U13621 (N_13621,N_11174,N_8950);
nor U13622 (N_13622,N_9011,N_10796);
and U13623 (N_13623,N_9512,N_8514);
and U13624 (N_13624,N_9215,N_9901);
nor U13625 (N_13625,N_11407,N_9874);
nor U13626 (N_13626,N_10166,N_9617);
nand U13627 (N_13627,N_10823,N_11588);
xnor U13628 (N_13628,N_8692,N_11015);
nor U13629 (N_13629,N_10419,N_11555);
or U13630 (N_13630,N_8939,N_8244);
or U13631 (N_13631,N_8408,N_9028);
nor U13632 (N_13632,N_9801,N_8041);
xor U13633 (N_13633,N_8340,N_8829);
nand U13634 (N_13634,N_9879,N_10491);
or U13635 (N_13635,N_9087,N_9472);
and U13636 (N_13636,N_10810,N_9354);
xor U13637 (N_13637,N_11740,N_10540);
nand U13638 (N_13638,N_10579,N_9117);
or U13639 (N_13639,N_8248,N_8382);
and U13640 (N_13640,N_10097,N_8246);
or U13641 (N_13641,N_11963,N_10608);
nor U13642 (N_13642,N_9609,N_11072);
xor U13643 (N_13643,N_10836,N_10911);
or U13644 (N_13644,N_8331,N_11536);
nand U13645 (N_13645,N_8334,N_9306);
and U13646 (N_13646,N_8478,N_8308);
and U13647 (N_13647,N_9337,N_8042);
and U13648 (N_13648,N_10494,N_11815);
nand U13649 (N_13649,N_10536,N_9844);
nand U13650 (N_13650,N_10504,N_8500);
xor U13651 (N_13651,N_10534,N_10047);
nor U13652 (N_13652,N_9326,N_10331);
or U13653 (N_13653,N_9539,N_11987);
nor U13654 (N_13654,N_9775,N_11800);
and U13655 (N_13655,N_9085,N_10703);
or U13656 (N_13656,N_10152,N_8093);
nand U13657 (N_13657,N_11027,N_8410);
or U13658 (N_13658,N_9194,N_11832);
and U13659 (N_13659,N_11374,N_11638);
nor U13660 (N_13660,N_8920,N_8216);
xor U13661 (N_13661,N_10800,N_8301);
and U13662 (N_13662,N_11886,N_11088);
or U13663 (N_13663,N_11291,N_9486);
or U13664 (N_13664,N_10700,N_8002);
or U13665 (N_13665,N_9686,N_9434);
nand U13666 (N_13666,N_8959,N_9564);
nand U13667 (N_13667,N_10093,N_10241);
nor U13668 (N_13668,N_8474,N_10904);
xor U13669 (N_13669,N_8659,N_8887);
or U13670 (N_13670,N_10962,N_9500);
nand U13671 (N_13671,N_9136,N_11336);
xnor U13672 (N_13672,N_10192,N_8167);
or U13673 (N_13673,N_11694,N_8651);
nor U13674 (N_13674,N_8180,N_8206);
xor U13675 (N_13675,N_10377,N_10464);
nand U13676 (N_13676,N_8756,N_9898);
nor U13677 (N_13677,N_8172,N_10274);
nand U13678 (N_13678,N_11798,N_9081);
nand U13679 (N_13679,N_10363,N_11810);
and U13680 (N_13680,N_11524,N_9264);
nor U13681 (N_13681,N_10466,N_10561);
nor U13682 (N_13682,N_10841,N_9982);
nor U13683 (N_13683,N_10174,N_11935);
nor U13684 (N_13684,N_9238,N_9455);
or U13685 (N_13685,N_9364,N_10776);
or U13686 (N_13686,N_10830,N_8179);
nor U13687 (N_13687,N_9543,N_8275);
or U13688 (N_13688,N_11198,N_11073);
or U13689 (N_13689,N_8375,N_11178);
or U13690 (N_13690,N_9269,N_9656);
nand U13691 (N_13691,N_8356,N_10640);
nor U13692 (N_13692,N_8290,N_8217);
nand U13693 (N_13693,N_10392,N_10434);
or U13694 (N_13694,N_10524,N_11646);
and U13695 (N_13695,N_10064,N_10956);
nand U13696 (N_13696,N_10441,N_8219);
or U13697 (N_13697,N_8770,N_11837);
or U13698 (N_13698,N_10133,N_8980);
nor U13699 (N_13699,N_10167,N_9334);
xor U13700 (N_13700,N_9546,N_10482);
nor U13701 (N_13701,N_10337,N_8991);
nand U13702 (N_13702,N_11550,N_8173);
nor U13703 (N_13703,N_10066,N_10859);
or U13704 (N_13704,N_10727,N_10447);
nand U13705 (N_13705,N_8748,N_10230);
nor U13706 (N_13706,N_9425,N_11294);
nand U13707 (N_13707,N_10902,N_11038);
xor U13708 (N_13708,N_9145,N_9527);
nor U13709 (N_13709,N_10222,N_11318);
nor U13710 (N_13710,N_8973,N_10620);
xnor U13711 (N_13711,N_10903,N_8563);
nor U13712 (N_13712,N_8911,N_10916);
nand U13713 (N_13713,N_10706,N_10195);
nor U13714 (N_13714,N_9965,N_11660);
and U13715 (N_13715,N_10071,N_10603);
xnor U13716 (N_13716,N_8231,N_9164);
xnor U13717 (N_13717,N_10882,N_9749);
nor U13718 (N_13718,N_11736,N_8893);
nor U13719 (N_13719,N_11367,N_8013);
nor U13720 (N_13720,N_10138,N_8431);
xor U13721 (N_13721,N_9950,N_10743);
xnor U13722 (N_13722,N_9080,N_8085);
xor U13723 (N_13723,N_9940,N_11871);
or U13724 (N_13724,N_8669,N_11273);
nor U13725 (N_13725,N_9877,N_11868);
or U13726 (N_13726,N_9596,N_8459);
nand U13727 (N_13727,N_9964,N_8935);
xor U13728 (N_13728,N_9150,N_10078);
nor U13729 (N_13729,N_8412,N_9181);
nand U13730 (N_13730,N_10523,N_10130);
nor U13731 (N_13731,N_9576,N_8717);
or U13732 (N_13732,N_8745,N_11527);
or U13733 (N_13733,N_10589,N_10897);
xnor U13734 (N_13734,N_11964,N_8402);
or U13735 (N_13735,N_10288,N_10951);
nor U13736 (N_13736,N_8483,N_8910);
nand U13737 (N_13737,N_8255,N_11519);
and U13738 (N_13738,N_8967,N_11671);
or U13739 (N_13739,N_11243,N_11476);
or U13740 (N_13740,N_10424,N_9110);
xor U13741 (N_13741,N_8250,N_8161);
nor U13742 (N_13742,N_10973,N_9769);
xnor U13743 (N_13743,N_11777,N_9118);
nand U13744 (N_13744,N_9722,N_10839);
and U13745 (N_13745,N_10846,N_10845);
xor U13746 (N_13746,N_9002,N_11192);
or U13747 (N_13747,N_9661,N_8134);
nor U13748 (N_13748,N_9226,N_10396);
and U13749 (N_13749,N_11084,N_11408);
and U13750 (N_13750,N_11195,N_10604);
or U13751 (N_13751,N_10211,N_8249);
and U13752 (N_13752,N_8337,N_10908);
xor U13753 (N_13753,N_8587,N_9635);
xor U13754 (N_13754,N_10672,N_8971);
nor U13755 (N_13755,N_9966,N_11079);
nor U13756 (N_13756,N_11794,N_9016);
nor U13757 (N_13757,N_8333,N_11116);
xor U13758 (N_13758,N_11045,N_8992);
xnor U13759 (N_13759,N_8452,N_8247);
or U13760 (N_13760,N_10213,N_11261);
or U13761 (N_13761,N_10551,N_9792);
xnor U13762 (N_13762,N_11665,N_8309);
xor U13763 (N_13763,N_9620,N_11205);
nor U13764 (N_13764,N_9484,N_8092);
and U13765 (N_13765,N_11289,N_10646);
xor U13766 (N_13766,N_9991,N_8286);
nor U13767 (N_13767,N_8672,N_8987);
xnor U13768 (N_13768,N_10648,N_11727);
or U13769 (N_13769,N_10607,N_10642);
xnor U13770 (N_13770,N_9383,N_9496);
nor U13771 (N_13771,N_9558,N_9798);
and U13772 (N_13772,N_10753,N_8078);
or U13773 (N_13773,N_9772,N_11383);
nor U13774 (N_13774,N_9286,N_11164);
or U13775 (N_13775,N_8559,N_10103);
and U13776 (N_13776,N_11969,N_11150);
and U13777 (N_13777,N_8147,N_11051);
xor U13778 (N_13778,N_8116,N_11421);
and U13779 (N_13779,N_11460,N_9219);
or U13780 (N_13780,N_11295,N_8857);
nor U13781 (N_13781,N_11614,N_9545);
or U13782 (N_13782,N_11574,N_9606);
nand U13783 (N_13783,N_10405,N_9700);
nor U13784 (N_13784,N_10165,N_9012);
and U13785 (N_13785,N_11788,N_11117);
nor U13786 (N_13786,N_11997,N_11309);
or U13787 (N_13787,N_9942,N_11229);
or U13788 (N_13788,N_10224,N_8014);
nor U13789 (N_13789,N_10219,N_8492);
nand U13790 (N_13790,N_10106,N_8446);
or U13791 (N_13791,N_11410,N_8731);
xor U13792 (N_13792,N_11932,N_11920);
nand U13793 (N_13793,N_11425,N_10117);
xnor U13794 (N_13794,N_11894,N_9441);
xnor U13795 (N_13795,N_10856,N_8008);
and U13796 (N_13796,N_9604,N_11017);
xnor U13797 (N_13797,N_11512,N_10993);
nor U13798 (N_13798,N_8926,N_10004);
nor U13799 (N_13799,N_11416,N_11344);
xor U13800 (N_13800,N_9475,N_9574);
xor U13801 (N_13801,N_11477,N_9565);
and U13802 (N_13802,N_11862,N_9618);
nand U13803 (N_13803,N_11927,N_9521);
nand U13804 (N_13804,N_9507,N_10371);
and U13805 (N_13805,N_11704,N_10548);
or U13806 (N_13806,N_11509,N_10857);
nand U13807 (N_13807,N_8472,N_8560);
nand U13808 (N_13808,N_10404,N_9976);
and U13809 (N_13809,N_11564,N_9937);
xnor U13810 (N_13810,N_8925,N_9559);
xnor U13811 (N_13811,N_8646,N_8504);
nor U13812 (N_13812,N_9645,N_8610);
or U13813 (N_13813,N_9823,N_8722);
xor U13814 (N_13814,N_10582,N_10055);
nor U13815 (N_13815,N_9260,N_10829);
and U13816 (N_13816,N_8281,N_8978);
or U13817 (N_13817,N_9621,N_11077);
or U13818 (N_13818,N_8165,N_11729);
nor U13819 (N_13819,N_10590,N_11915);
nand U13820 (N_13820,N_8212,N_10585);
and U13821 (N_13821,N_10008,N_9162);
xnor U13822 (N_13822,N_10007,N_11025);
xor U13823 (N_13823,N_8099,N_8329);
and U13824 (N_13824,N_10552,N_11081);
xnor U13825 (N_13825,N_8611,N_10528);
xor U13826 (N_13826,N_9050,N_9634);
and U13827 (N_13827,N_10385,N_8257);
nor U13828 (N_13828,N_11314,N_9744);
or U13829 (N_13829,N_9657,N_11026);
or U13830 (N_13830,N_11436,N_10605);
and U13831 (N_13831,N_10865,N_11157);
xnor U13832 (N_13832,N_10821,N_8997);
xor U13833 (N_13833,N_10929,N_11463);
or U13834 (N_13834,N_9380,N_8124);
and U13835 (N_13835,N_10518,N_9026);
nor U13836 (N_13836,N_8977,N_8430);
and U13837 (N_13837,N_9996,N_10984);
and U13838 (N_13838,N_11041,N_9221);
and U13839 (N_13839,N_9116,N_11786);
nor U13840 (N_13840,N_10760,N_8395);
and U13841 (N_13841,N_9229,N_9553);
nand U13842 (N_13842,N_8265,N_10938);
or U13843 (N_13843,N_8613,N_10021);
xor U13844 (N_13844,N_10740,N_10041);
nand U13845 (N_13845,N_8941,N_9358);
and U13846 (N_13846,N_8776,N_10426);
xor U13847 (N_13847,N_10650,N_8298);
nand U13848 (N_13848,N_10233,N_8096);
nor U13849 (N_13849,N_9474,N_11939);
or U13850 (N_13850,N_11267,N_10654);
xnor U13851 (N_13851,N_11984,N_11732);
xnor U13852 (N_13852,N_11892,N_11884);
and U13853 (N_13853,N_11391,N_10483);
nor U13854 (N_13854,N_8534,N_8462);
xor U13855 (N_13855,N_11172,N_8943);
or U13856 (N_13856,N_9152,N_11484);
and U13857 (N_13857,N_9577,N_8688);
nor U13858 (N_13858,N_9562,N_9696);
xnor U13859 (N_13859,N_8568,N_10822);
and U13860 (N_13860,N_11895,N_11505);
nor U13861 (N_13861,N_10375,N_9771);
nand U13862 (N_13862,N_10271,N_8614);
nor U13863 (N_13863,N_8728,N_10260);
or U13864 (N_13864,N_11028,N_11511);
or U13865 (N_13865,N_9324,N_8513);
xor U13866 (N_13866,N_11888,N_9245);
and U13867 (N_13867,N_8083,N_9752);
or U13868 (N_13868,N_9044,N_8456);
or U13869 (N_13869,N_9084,N_8710);
xor U13870 (N_13870,N_8484,N_11276);
nand U13871 (N_13871,N_11171,N_9867);
xnor U13872 (N_13872,N_10901,N_10018);
or U13873 (N_13873,N_11880,N_10527);
or U13874 (N_13874,N_11099,N_10147);
nor U13875 (N_13875,N_10946,N_11371);
and U13876 (N_13876,N_8145,N_9456);
or U13877 (N_13877,N_11362,N_10667);
xnor U13878 (N_13878,N_10123,N_10065);
xnor U13879 (N_13879,N_11497,N_8727);
nor U13880 (N_13880,N_10327,N_10281);
xnor U13881 (N_13881,N_9748,N_9186);
and U13882 (N_13882,N_11348,N_11156);
or U13883 (N_13883,N_11683,N_8666);
xor U13884 (N_13884,N_9303,N_11949);
or U13885 (N_13885,N_11376,N_11414);
or U13886 (N_13886,N_9112,N_8936);
and U13887 (N_13887,N_11139,N_10248);
nand U13888 (N_13888,N_11199,N_9843);
nand U13889 (N_13889,N_8202,N_9490);
nor U13890 (N_13890,N_9768,N_11835);
nor U13891 (N_13891,N_10759,N_9328);
xnor U13892 (N_13892,N_10578,N_9056);
nand U13893 (N_13893,N_9203,N_11858);
and U13894 (N_13894,N_11103,N_8486);
xor U13895 (N_13895,N_11281,N_10741);
nor U13896 (N_13896,N_10298,N_8209);
or U13897 (N_13897,N_11924,N_8743);
nor U13898 (N_13898,N_10416,N_8174);
nand U13899 (N_13899,N_8741,N_8689);
nor U13900 (N_13900,N_10801,N_9134);
and U13901 (N_13901,N_10400,N_9374);
nor U13902 (N_13902,N_10085,N_9077);
nor U13903 (N_13903,N_10341,N_10510);
nor U13904 (N_13904,N_9643,N_8797);
or U13905 (N_13905,N_11078,N_10543);
xnor U13906 (N_13906,N_9953,N_10294);
xnor U13907 (N_13907,N_10096,N_8734);
nand U13908 (N_13908,N_9808,N_10019);
or U13909 (N_13909,N_9731,N_10280);
and U13910 (N_13910,N_9481,N_8113);
nor U13911 (N_13911,N_9235,N_11651);
and U13912 (N_13912,N_9529,N_9631);
and U13913 (N_13913,N_9934,N_8638);
nand U13914 (N_13914,N_10107,N_9610);
or U13915 (N_13915,N_9299,N_9065);
nand U13916 (N_13916,N_8371,N_9969);
xnor U13917 (N_13917,N_8184,N_8110);
and U13918 (N_13918,N_8547,N_10121);
nand U13919 (N_13919,N_9368,N_11355);
or U13920 (N_13920,N_10965,N_11904);
nand U13921 (N_13921,N_11758,N_9282);
and U13922 (N_13922,N_9414,N_9442);
xnor U13923 (N_13923,N_9858,N_9987);
nand U13924 (N_13924,N_9409,N_9344);
xnor U13925 (N_13925,N_11643,N_10957);
nor U13926 (N_13926,N_8122,N_11608);
xor U13927 (N_13927,N_11873,N_9781);
xor U13928 (N_13928,N_11921,N_8818);
or U13929 (N_13929,N_11464,N_9796);
xnor U13930 (N_13930,N_10926,N_11834);
xnor U13931 (N_13931,N_11046,N_10198);
or U13932 (N_13932,N_10459,N_10876);
nor U13933 (N_13933,N_11203,N_11000);
nor U13934 (N_13934,N_8109,N_10661);
or U13935 (N_13935,N_9140,N_9682);
or U13936 (N_13936,N_8159,N_8785);
and U13937 (N_13937,N_8288,N_9304);
nor U13938 (N_13938,N_10777,N_11928);
and U13939 (N_13939,N_10462,N_10554);
nor U13940 (N_13940,N_10596,N_11239);
or U13941 (N_13941,N_9875,N_11981);
nor U13942 (N_13942,N_10556,N_9308);
nand U13943 (N_13943,N_8241,N_11515);
or U13944 (N_13944,N_9446,N_10885);
nand U13945 (N_13945,N_10905,N_8890);
or U13946 (N_13946,N_11670,N_10550);
and U13947 (N_13947,N_9451,N_10995);
or U13948 (N_13948,N_10625,N_11649);
or U13949 (N_13949,N_8658,N_9889);
or U13950 (N_13950,N_11597,N_9204);
and U13951 (N_13951,N_8185,N_9501);
or U13952 (N_13952,N_10428,N_9343);
and U13953 (N_13953,N_9096,N_9859);
and U13954 (N_13954,N_11280,N_9210);
nor U13955 (N_13955,N_10332,N_10814);
nor U13956 (N_13956,N_11210,N_9068);
xor U13957 (N_13957,N_9599,N_10771);
and U13958 (N_13958,N_9274,N_11823);
nand U13959 (N_13959,N_11074,N_10898);
and U13960 (N_13960,N_10950,N_10301);
and U13961 (N_13961,N_9095,N_11983);
or U13962 (N_13962,N_8021,N_9426);
xnor U13963 (N_13963,N_9888,N_8719);
and U13964 (N_13964,N_9157,N_11522);
nor U13965 (N_13965,N_9184,N_11633);
xor U13966 (N_13966,N_8397,N_11562);
and U13967 (N_13967,N_8607,N_9905);
and U13968 (N_13968,N_8667,N_8363);
nand U13969 (N_13969,N_9353,N_11208);
or U13970 (N_13970,N_9721,N_11733);
or U13971 (N_13971,N_9579,N_9786);
nor U13972 (N_13972,N_9263,N_10102);
nand U13973 (N_13973,N_9059,N_8141);
nor U13974 (N_13974,N_8983,N_9416);
nand U13975 (N_13975,N_11474,N_10936);
and U13976 (N_13976,N_9331,N_8178);
or U13977 (N_13977,N_10999,N_10733);
xor U13978 (N_13978,N_8074,N_10507);
nor U13979 (N_13979,N_11829,N_10838);
and U13980 (N_13980,N_10639,N_9929);
or U13981 (N_13981,N_8253,N_8191);
nor U13982 (N_13982,N_8796,N_10418);
nor U13983 (N_13983,N_11783,N_9852);
and U13984 (N_13984,N_9108,N_9612);
nand U13985 (N_13985,N_10495,N_9379);
xnor U13986 (N_13986,N_10146,N_11105);
nor U13987 (N_13987,N_11012,N_11257);
nor U13988 (N_13988,N_10031,N_9759);
nand U13989 (N_13989,N_10421,N_11332);
nor U13990 (N_13990,N_11885,N_10086);
or U13991 (N_13991,N_8664,N_9678);
xnor U13992 (N_13992,N_8606,N_11230);
nor U13993 (N_13993,N_11136,N_10249);
nand U13994 (N_13994,N_11989,N_9397);
xor U13995 (N_13995,N_11402,N_9283);
nor U13996 (N_13996,N_10502,N_10448);
nor U13997 (N_13997,N_11226,N_8274);
nor U13998 (N_13998,N_9214,N_8798);
nor U13999 (N_13999,N_11001,N_10389);
or U14000 (N_14000,N_11859,N_11010);
nand U14001 (N_14001,N_11926,N_11847);
nor U14002 (N_14002,N_10230,N_9584);
nand U14003 (N_14003,N_10301,N_8426);
xnor U14004 (N_14004,N_9027,N_9082);
and U14005 (N_14005,N_11899,N_10363);
nand U14006 (N_14006,N_11823,N_10310);
and U14007 (N_14007,N_11229,N_10249);
or U14008 (N_14008,N_9258,N_8411);
xor U14009 (N_14009,N_8001,N_10920);
xnor U14010 (N_14010,N_9807,N_11235);
or U14011 (N_14011,N_8318,N_8676);
nand U14012 (N_14012,N_10385,N_11682);
or U14013 (N_14013,N_9136,N_11636);
and U14014 (N_14014,N_9336,N_8269);
and U14015 (N_14015,N_9862,N_10659);
xor U14016 (N_14016,N_8843,N_9107);
nand U14017 (N_14017,N_9028,N_9726);
nor U14018 (N_14018,N_10305,N_11776);
nand U14019 (N_14019,N_11801,N_10711);
nor U14020 (N_14020,N_10009,N_8735);
or U14021 (N_14021,N_9057,N_10312);
nor U14022 (N_14022,N_9654,N_8816);
nand U14023 (N_14023,N_9617,N_11388);
nand U14024 (N_14024,N_11103,N_10552);
and U14025 (N_14025,N_8237,N_11249);
xnor U14026 (N_14026,N_10846,N_11458);
xnor U14027 (N_14027,N_9118,N_10011);
or U14028 (N_14028,N_10627,N_8367);
nor U14029 (N_14029,N_8977,N_10789);
nand U14030 (N_14030,N_8606,N_8823);
xnor U14031 (N_14031,N_8148,N_9486);
nand U14032 (N_14032,N_8455,N_11962);
and U14033 (N_14033,N_9420,N_10511);
xor U14034 (N_14034,N_8769,N_10698);
nor U14035 (N_14035,N_8227,N_8685);
or U14036 (N_14036,N_9240,N_11672);
and U14037 (N_14037,N_9278,N_10878);
or U14038 (N_14038,N_10436,N_9647);
or U14039 (N_14039,N_11964,N_8839);
nor U14040 (N_14040,N_9645,N_8603);
and U14041 (N_14041,N_9084,N_8311);
nor U14042 (N_14042,N_8331,N_8349);
xnor U14043 (N_14043,N_9379,N_10535);
and U14044 (N_14044,N_10595,N_9889);
nor U14045 (N_14045,N_8466,N_11304);
and U14046 (N_14046,N_9181,N_8591);
nor U14047 (N_14047,N_8744,N_10068);
xnor U14048 (N_14048,N_9667,N_10765);
and U14049 (N_14049,N_8729,N_8293);
nor U14050 (N_14050,N_10258,N_10988);
nand U14051 (N_14051,N_9853,N_10303);
xnor U14052 (N_14052,N_10128,N_8521);
or U14053 (N_14053,N_8510,N_10676);
nand U14054 (N_14054,N_8461,N_9832);
xor U14055 (N_14055,N_9217,N_10144);
nor U14056 (N_14056,N_9073,N_11252);
and U14057 (N_14057,N_10835,N_10834);
nand U14058 (N_14058,N_9246,N_11419);
or U14059 (N_14059,N_8951,N_11139);
nand U14060 (N_14060,N_9442,N_11423);
nand U14061 (N_14061,N_8345,N_10085);
nor U14062 (N_14062,N_11199,N_11241);
nand U14063 (N_14063,N_8423,N_8775);
or U14064 (N_14064,N_8925,N_9190);
nor U14065 (N_14065,N_11082,N_9642);
xor U14066 (N_14066,N_11144,N_10431);
or U14067 (N_14067,N_8731,N_11284);
nor U14068 (N_14068,N_11577,N_11494);
nand U14069 (N_14069,N_10037,N_8534);
or U14070 (N_14070,N_10211,N_8440);
and U14071 (N_14071,N_8658,N_9497);
xnor U14072 (N_14072,N_10159,N_8327);
nand U14073 (N_14073,N_8918,N_8881);
or U14074 (N_14074,N_9216,N_11361);
nor U14075 (N_14075,N_11467,N_11488);
or U14076 (N_14076,N_10071,N_8401);
or U14077 (N_14077,N_9790,N_10338);
and U14078 (N_14078,N_8358,N_9232);
nand U14079 (N_14079,N_11007,N_8721);
xor U14080 (N_14080,N_10549,N_8089);
or U14081 (N_14081,N_10606,N_11179);
nor U14082 (N_14082,N_11320,N_11024);
and U14083 (N_14083,N_9542,N_8876);
nand U14084 (N_14084,N_11879,N_8865);
xnor U14085 (N_14085,N_11877,N_9059);
and U14086 (N_14086,N_10720,N_11988);
and U14087 (N_14087,N_9571,N_8816);
nor U14088 (N_14088,N_11424,N_8393);
xor U14089 (N_14089,N_11508,N_10047);
nand U14090 (N_14090,N_8910,N_10761);
nand U14091 (N_14091,N_11138,N_11238);
nand U14092 (N_14092,N_10526,N_9192);
and U14093 (N_14093,N_11704,N_8283);
or U14094 (N_14094,N_11852,N_9905);
nand U14095 (N_14095,N_11366,N_11951);
and U14096 (N_14096,N_8191,N_8036);
xor U14097 (N_14097,N_11731,N_10254);
or U14098 (N_14098,N_8800,N_8342);
nand U14099 (N_14099,N_8294,N_8644);
or U14100 (N_14100,N_10754,N_10549);
or U14101 (N_14101,N_11901,N_10835);
nor U14102 (N_14102,N_11069,N_9910);
nor U14103 (N_14103,N_11500,N_10493);
nor U14104 (N_14104,N_10028,N_9577);
or U14105 (N_14105,N_9925,N_8187);
and U14106 (N_14106,N_11900,N_9116);
nor U14107 (N_14107,N_8854,N_8034);
or U14108 (N_14108,N_9497,N_10523);
nand U14109 (N_14109,N_10180,N_9139);
nor U14110 (N_14110,N_9340,N_9787);
xor U14111 (N_14111,N_8955,N_11579);
nand U14112 (N_14112,N_8108,N_9603);
and U14113 (N_14113,N_8818,N_11266);
and U14114 (N_14114,N_8369,N_9155);
and U14115 (N_14115,N_9993,N_11619);
xnor U14116 (N_14116,N_11622,N_9076);
nor U14117 (N_14117,N_11116,N_8525);
xor U14118 (N_14118,N_11878,N_10516);
nand U14119 (N_14119,N_8256,N_11355);
or U14120 (N_14120,N_11703,N_11126);
nand U14121 (N_14121,N_9096,N_8971);
nor U14122 (N_14122,N_11296,N_11482);
xor U14123 (N_14123,N_11555,N_9881);
nor U14124 (N_14124,N_10906,N_11877);
nor U14125 (N_14125,N_9495,N_9923);
xnor U14126 (N_14126,N_11175,N_11770);
xnor U14127 (N_14127,N_9143,N_11425);
or U14128 (N_14128,N_8208,N_10099);
nor U14129 (N_14129,N_8803,N_8761);
nor U14130 (N_14130,N_9974,N_8810);
or U14131 (N_14131,N_11194,N_10494);
and U14132 (N_14132,N_9391,N_11907);
nor U14133 (N_14133,N_11986,N_11200);
xor U14134 (N_14134,N_11916,N_8159);
xnor U14135 (N_14135,N_11111,N_9678);
nand U14136 (N_14136,N_9598,N_10844);
xor U14137 (N_14137,N_8891,N_10008);
and U14138 (N_14138,N_8245,N_11978);
and U14139 (N_14139,N_10904,N_11492);
and U14140 (N_14140,N_9418,N_11763);
nor U14141 (N_14141,N_9887,N_9918);
xor U14142 (N_14142,N_10694,N_11938);
nor U14143 (N_14143,N_8551,N_8425);
nand U14144 (N_14144,N_9429,N_11789);
nor U14145 (N_14145,N_11441,N_10985);
nor U14146 (N_14146,N_9486,N_10828);
and U14147 (N_14147,N_9511,N_11869);
and U14148 (N_14148,N_11422,N_9214);
and U14149 (N_14149,N_10172,N_9253);
and U14150 (N_14150,N_10007,N_8207);
nor U14151 (N_14151,N_8473,N_9716);
nor U14152 (N_14152,N_10239,N_10050);
xnor U14153 (N_14153,N_10296,N_10083);
or U14154 (N_14154,N_9178,N_9250);
nor U14155 (N_14155,N_10459,N_10117);
xnor U14156 (N_14156,N_8057,N_9255);
or U14157 (N_14157,N_11132,N_8406);
or U14158 (N_14158,N_8376,N_10137);
nand U14159 (N_14159,N_11101,N_8596);
or U14160 (N_14160,N_11365,N_8662);
and U14161 (N_14161,N_11055,N_10026);
nand U14162 (N_14162,N_10575,N_10464);
or U14163 (N_14163,N_11055,N_8272);
nand U14164 (N_14164,N_10301,N_9406);
nand U14165 (N_14165,N_8224,N_10965);
xnor U14166 (N_14166,N_8751,N_11117);
xnor U14167 (N_14167,N_8046,N_8393);
nor U14168 (N_14168,N_11905,N_11675);
xor U14169 (N_14169,N_10574,N_10759);
or U14170 (N_14170,N_8665,N_8732);
nand U14171 (N_14171,N_10499,N_10940);
nand U14172 (N_14172,N_10204,N_9215);
xor U14173 (N_14173,N_9894,N_10845);
xor U14174 (N_14174,N_8423,N_10750);
and U14175 (N_14175,N_9907,N_11731);
nor U14176 (N_14176,N_11361,N_11891);
xor U14177 (N_14177,N_8865,N_9635);
xnor U14178 (N_14178,N_8163,N_9211);
or U14179 (N_14179,N_8784,N_10503);
nand U14180 (N_14180,N_11194,N_10482);
xnor U14181 (N_14181,N_8015,N_10320);
and U14182 (N_14182,N_11414,N_9187);
or U14183 (N_14183,N_9080,N_10679);
nor U14184 (N_14184,N_10949,N_8655);
nor U14185 (N_14185,N_8294,N_11032);
or U14186 (N_14186,N_11037,N_9833);
nand U14187 (N_14187,N_9131,N_10636);
xnor U14188 (N_14188,N_11602,N_8937);
nand U14189 (N_14189,N_11430,N_10684);
nand U14190 (N_14190,N_10231,N_10081);
nor U14191 (N_14191,N_9720,N_9151);
nor U14192 (N_14192,N_8839,N_10194);
or U14193 (N_14193,N_10834,N_11051);
and U14194 (N_14194,N_8394,N_8977);
or U14195 (N_14195,N_11578,N_11328);
nor U14196 (N_14196,N_11078,N_9500);
xnor U14197 (N_14197,N_11417,N_8770);
and U14198 (N_14198,N_9448,N_11601);
nor U14199 (N_14199,N_10236,N_11399);
nor U14200 (N_14200,N_11752,N_11822);
or U14201 (N_14201,N_8801,N_11578);
or U14202 (N_14202,N_11742,N_11970);
or U14203 (N_14203,N_8548,N_10227);
nor U14204 (N_14204,N_9812,N_10254);
and U14205 (N_14205,N_10304,N_10236);
or U14206 (N_14206,N_8332,N_10905);
nand U14207 (N_14207,N_9817,N_10763);
nor U14208 (N_14208,N_11241,N_10627);
nor U14209 (N_14209,N_9554,N_8346);
nand U14210 (N_14210,N_10276,N_10357);
and U14211 (N_14211,N_10090,N_11745);
xor U14212 (N_14212,N_11094,N_8425);
and U14213 (N_14213,N_9559,N_8155);
xnor U14214 (N_14214,N_8539,N_10186);
and U14215 (N_14215,N_11092,N_10518);
and U14216 (N_14216,N_9745,N_9724);
and U14217 (N_14217,N_9925,N_9066);
nand U14218 (N_14218,N_8886,N_9616);
nand U14219 (N_14219,N_9485,N_8063);
and U14220 (N_14220,N_11721,N_10754);
nand U14221 (N_14221,N_11422,N_10623);
nand U14222 (N_14222,N_8242,N_8447);
and U14223 (N_14223,N_8775,N_9471);
nand U14224 (N_14224,N_10002,N_11481);
or U14225 (N_14225,N_10567,N_11194);
and U14226 (N_14226,N_11191,N_11144);
nor U14227 (N_14227,N_9684,N_10052);
or U14228 (N_14228,N_9416,N_10769);
xor U14229 (N_14229,N_11061,N_11901);
or U14230 (N_14230,N_11700,N_8287);
and U14231 (N_14231,N_9367,N_8893);
nor U14232 (N_14232,N_11901,N_10707);
nor U14233 (N_14233,N_10928,N_9039);
and U14234 (N_14234,N_11104,N_8875);
and U14235 (N_14235,N_8278,N_8995);
or U14236 (N_14236,N_10846,N_11590);
and U14237 (N_14237,N_11115,N_8234);
nor U14238 (N_14238,N_8768,N_9721);
and U14239 (N_14239,N_9164,N_8211);
and U14240 (N_14240,N_9688,N_9428);
nand U14241 (N_14241,N_10314,N_8785);
nor U14242 (N_14242,N_11061,N_8838);
xnor U14243 (N_14243,N_11677,N_9896);
xnor U14244 (N_14244,N_9178,N_11723);
or U14245 (N_14245,N_8819,N_10111);
nand U14246 (N_14246,N_10237,N_9455);
xor U14247 (N_14247,N_11163,N_8033);
nand U14248 (N_14248,N_10977,N_9525);
and U14249 (N_14249,N_8167,N_11319);
and U14250 (N_14250,N_9260,N_9018);
or U14251 (N_14251,N_11160,N_11911);
xnor U14252 (N_14252,N_11423,N_8429);
or U14253 (N_14253,N_8836,N_10897);
nand U14254 (N_14254,N_10442,N_11087);
or U14255 (N_14255,N_9717,N_11460);
xnor U14256 (N_14256,N_10056,N_8654);
nor U14257 (N_14257,N_9322,N_9298);
or U14258 (N_14258,N_10777,N_10371);
or U14259 (N_14259,N_10811,N_8227);
xnor U14260 (N_14260,N_9979,N_10132);
or U14261 (N_14261,N_9431,N_10365);
nand U14262 (N_14262,N_10643,N_8439);
nor U14263 (N_14263,N_8598,N_9197);
or U14264 (N_14264,N_10143,N_10673);
xnor U14265 (N_14265,N_11937,N_9429);
and U14266 (N_14266,N_10624,N_11276);
or U14267 (N_14267,N_9692,N_11866);
xor U14268 (N_14268,N_10399,N_11790);
xnor U14269 (N_14269,N_8937,N_11191);
xnor U14270 (N_14270,N_9656,N_11268);
or U14271 (N_14271,N_8215,N_10713);
or U14272 (N_14272,N_10540,N_8748);
or U14273 (N_14273,N_8349,N_11722);
and U14274 (N_14274,N_11645,N_11015);
or U14275 (N_14275,N_9406,N_8933);
nand U14276 (N_14276,N_11138,N_8487);
nor U14277 (N_14277,N_8663,N_10020);
nand U14278 (N_14278,N_10716,N_11126);
xnor U14279 (N_14279,N_11768,N_10909);
nand U14280 (N_14280,N_10265,N_11185);
nor U14281 (N_14281,N_11804,N_8649);
nor U14282 (N_14282,N_11463,N_8360);
nand U14283 (N_14283,N_10813,N_11462);
nand U14284 (N_14284,N_11582,N_10757);
xor U14285 (N_14285,N_9291,N_11696);
and U14286 (N_14286,N_8867,N_11127);
nand U14287 (N_14287,N_9975,N_9135);
and U14288 (N_14288,N_10071,N_8389);
or U14289 (N_14289,N_8338,N_8634);
and U14290 (N_14290,N_11714,N_8673);
nor U14291 (N_14291,N_11799,N_11992);
xor U14292 (N_14292,N_10266,N_8464);
nand U14293 (N_14293,N_8463,N_10352);
or U14294 (N_14294,N_9571,N_8946);
nand U14295 (N_14295,N_9343,N_10567);
and U14296 (N_14296,N_11553,N_11122);
or U14297 (N_14297,N_9400,N_8046);
and U14298 (N_14298,N_11625,N_9606);
xor U14299 (N_14299,N_8375,N_8740);
and U14300 (N_14300,N_8164,N_11559);
and U14301 (N_14301,N_8226,N_11981);
xnor U14302 (N_14302,N_8581,N_8619);
xor U14303 (N_14303,N_9069,N_9281);
nor U14304 (N_14304,N_10763,N_9959);
xor U14305 (N_14305,N_10292,N_8273);
or U14306 (N_14306,N_8200,N_11063);
or U14307 (N_14307,N_11520,N_9333);
nor U14308 (N_14308,N_10598,N_10036);
or U14309 (N_14309,N_11039,N_10052);
or U14310 (N_14310,N_8341,N_11732);
nor U14311 (N_14311,N_8021,N_9864);
and U14312 (N_14312,N_10315,N_11769);
and U14313 (N_14313,N_11595,N_10750);
and U14314 (N_14314,N_8436,N_8738);
and U14315 (N_14315,N_10049,N_10833);
and U14316 (N_14316,N_10081,N_8126);
xnor U14317 (N_14317,N_9441,N_11342);
and U14318 (N_14318,N_11977,N_8783);
and U14319 (N_14319,N_9709,N_8350);
xor U14320 (N_14320,N_9938,N_11227);
or U14321 (N_14321,N_9195,N_9647);
or U14322 (N_14322,N_9699,N_8074);
or U14323 (N_14323,N_9570,N_11850);
and U14324 (N_14324,N_9477,N_8797);
nand U14325 (N_14325,N_11941,N_10291);
xnor U14326 (N_14326,N_10576,N_8968);
xor U14327 (N_14327,N_8838,N_9160);
nor U14328 (N_14328,N_11580,N_9944);
xor U14329 (N_14329,N_11225,N_8468);
or U14330 (N_14330,N_8875,N_8425);
or U14331 (N_14331,N_11071,N_8586);
or U14332 (N_14332,N_10520,N_9309);
xnor U14333 (N_14333,N_10490,N_8214);
nand U14334 (N_14334,N_11133,N_9970);
or U14335 (N_14335,N_11661,N_9522);
nand U14336 (N_14336,N_10256,N_11406);
or U14337 (N_14337,N_8257,N_9972);
nor U14338 (N_14338,N_8964,N_8034);
xor U14339 (N_14339,N_8115,N_9064);
or U14340 (N_14340,N_8579,N_10265);
xor U14341 (N_14341,N_11460,N_11411);
nor U14342 (N_14342,N_10481,N_11336);
or U14343 (N_14343,N_8617,N_10695);
nor U14344 (N_14344,N_8704,N_11879);
nor U14345 (N_14345,N_11000,N_8452);
nand U14346 (N_14346,N_8822,N_11305);
nor U14347 (N_14347,N_11914,N_11182);
nor U14348 (N_14348,N_8851,N_10481);
and U14349 (N_14349,N_9321,N_8486);
or U14350 (N_14350,N_9101,N_11713);
or U14351 (N_14351,N_11840,N_8313);
or U14352 (N_14352,N_9374,N_9818);
nand U14353 (N_14353,N_10069,N_10641);
nand U14354 (N_14354,N_10020,N_10373);
and U14355 (N_14355,N_10455,N_11558);
xnor U14356 (N_14356,N_11163,N_9060);
and U14357 (N_14357,N_11484,N_11929);
xnor U14358 (N_14358,N_10528,N_9547);
xor U14359 (N_14359,N_9158,N_9220);
nand U14360 (N_14360,N_10865,N_8579);
and U14361 (N_14361,N_9907,N_10573);
xnor U14362 (N_14362,N_10673,N_8349);
and U14363 (N_14363,N_8025,N_8369);
xnor U14364 (N_14364,N_10069,N_10203);
xnor U14365 (N_14365,N_11843,N_8745);
nand U14366 (N_14366,N_8046,N_11120);
and U14367 (N_14367,N_8191,N_8635);
nand U14368 (N_14368,N_9674,N_10905);
or U14369 (N_14369,N_8839,N_10900);
nor U14370 (N_14370,N_9251,N_10751);
and U14371 (N_14371,N_9150,N_11055);
nor U14372 (N_14372,N_8616,N_11559);
nand U14373 (N_14373,N_11271,N_10130);
and U14374 (N_14374,N_9864,N_8750);
nand U14375 (N_14375,N_9252,N_10147);
xor U14376 (N_14376,N_11183,N_11809);
and U14377 (N_14377,N_8578,N_8544);
nand U14378 (N_14378,N_9753,N_8154);
nor U14379 (N_14379,N_11745,N_8956);
nand U14380 (N_14380,N_11765,N_8093);
nand U14381 (N_14381,N_8637,N_8438);
and U14382 (N_14382,N_10238,N_8515);
or U14383 (N_14383,N_10674,N_11951);
nand U14384 (N_14384,N_11266,N_11484);
nand U14385 (N_14385,N_9013,N_8509);
and U14386 (N_14386,N_11564,N_10837);
or U14387 (N_14387,N_10918,N_9673);
or U14388 (N_14388,N_11727,N_11590);
or U14389 (N_14389,N_11815,N_11173);
or U14390 (N_14390,N_11213,N_8747);
or U14391 (N_14391,N_10547,N_9913);
nor U14392 (N_14392,N_8710,N_11691);
and U14393 (N_14393,N_11873,N_9290);
and U14394 (N_14394,N_8586,N_10607);
xor U14395 (N_14395,N_8965,N_11830);
nand U14396 (N_14396,N_10513,N_11176);
xor U14397 (N_14397,N_9689,N_11838);
nand U14398 (N_14398,N_11078,N_11751);
and U14399 (N_14399,N_11384,N_11876);
nor U14400 (N_14400,N_9777,N_8654);
or U14401 (N_14401,N_11647,N_10290);
or U14402 (N_14402,N_9644,N_11615);
nor U14403 (N_14403,N_8485,N_8362);
and U14404 (N_14404,N_8218,N_10589);
nand U14405 (N_14405,N_9419,N_11460);
xor U14406 (N_14406,N_10503,N_11724);
nand U14407 (N_14407,N_10197,N_11766);
xnor U14408 (N_14408,N_11756,N_11841);
nor U14409 (N_14409,N_10344,N_8972);
nor U14410 (N_14410,N_8343,N_10667);
and U14411 (N_14411,N_9432,N_10324);
nand U14412 (N_14412,N_10250,N_10336);
xnor U14413 (N_14413,N_11289,N_11998);
or U14414 (N_14414,N_10706,N_8987);
nor U14415 (N_14415,N_9073,N_11223);
nor U14416 (N_14416,N_9894,N_9993);
xor U14417 (N_14417,N_11726,N_10111);
nor U14418 (N_14418,N_9085,N_11149);
nand U14419 (N_14419,N_9069,N_11032);
nor U14420 (N_14420,N_9717,N_9599);
nor U14421 (N_14421,N_8352,N_10278);
xnor U14422 (N_14422,N_11904,N_9920);
xnor U14423 (N_14423,N_11750,N_9575);
nand U14424 (N_14424,N_8643,N_8476);
nand U14425 (N_14425,N_11381,N_10323);
nor U14426 (N_14426,N_9252,N_10563);
or U14427 (N_14427,N_11775,N_9141);
nand U14428 (N_14428,N_11324,N_9975);
xor U14429 (N_14429,N_10810,N_10239);
and U14430 (N_14430,N_11107,N_8513);
nand U14431 (N_14431,N_9353,N_11560);
xnor U14432 (N_14432,N_8121,N_9199);
nand U14433 (N_14433,N_10282,N_10130);
nand U14434 (N_14434,N_11664,N_8584);
xor U14435 (N_14435,N_10609,N_10165);
and U14436 (N_14436,N_9274,N_9096);
and U14437 (N_14437,N_8372,N_9951);
xor U14438 (N_14438,N_9024,N_10444);
nand U14439 (N_14439,N_11590,N_9309);
or U14440 (N_14440,N_11995,N_8353);
or U14441 (N_14441,N_9623,N_8156);
and U14442 (N_14442,N_10203,N_11948);
nor U14443 (N_14443,N_10216,N_8592);
or U14444 (N_14444,N_9602,N_9643);
nor U14445 (N_14445,N_9948,N_8634);
xnor U14446 (N_14446,N_11242,N_11968);
nand U14447 (N_14447,N_11538,N_10369);
and U14448 (N_14448,N_11085,N_9222);
or U14449 (N_14449,N_8848,N_11700);
nand U14450 (N_14450,N_8102,N_11284);
nand U14451 (N_14451,N_9089,N_9393);
nor U14452 (N_14452,N_11297,N_11534);
or U14453 (N_14453,N_11220,N_11905);
nand U14454 (N_14454,N_10812,N_8031);
nand U14455 (N_14455,N_11334,N_10320);
and U14456 (N_14456,N_11617,N_11060);
nor U14457 (N_14457,N_9933,N_9120);
nor U14458 (N_14458,N_10935,N_8481);
and U14459 (N_14459,N_9794,N_9524);
nor U14460 (N_14460,N_11032,N_10571);
and U14461 (N_14461,N_8465,N_9146);
xnor U14462 (N_14462,N_8357,N_11343);
nand U14463 (N_14463,N_9417,N_8027);
and U14464 (N_14464,N_9190,N_10014);
nand U14465 (N_14465,N_9336,N_9738);
nor U14466 (N_14466,N_8736,N_10829);
xnor U14467 (N_14467,N_8480,N_8457);
or U14468 (N_14468,N_9715,N_9926);
xnor U14469 (N_14469,N_10343,N_8613);
and U14470 (N_14470,N_10168,N_11706);
xnor U14471 (N_14471,N_9011,N_11600);
or U14472 (N_14472,N_9005,N_11399);
xor U14473 (N_14473,N_9197,N_11370);
nand U14474 (N_14474,N_9469,N_8440);
xnor U14475 (N_14475,N_10901,N_8502);
and U14476 (N_14476,N_11657,N_9279);
or U14477 (N_14477,N_8038,N_8249);
and U14478 (N_14478,N_11297,N_10790);
and U14479 (N_14479,N_10344,N_9801);
nor U14480 (N_14480,N_8962,N_8780);
nand U14481 (N_14481,N_8202,N_11271);
and U14482 (N_14482,N_9400,N_8261);
nand U14483 (N_14483,N_11651,N_10961);
and U14484 (N_14484,N_8412,N_11590);
xnor U14485 (N_14485,N_11978,N_9216);
or U14486 (N_14486,N_11425,N_8077);
xnor U14487 (N_14487,N_8379,N_11221);
or U14488 (N_14488,N_8703,N_11903);
nand U14489 (N_14489,N_11408,N_9707);
or U14490 (N_14490,N_9366,N_9102);
xnor U14491 (N_14491,N_11147,N_9372);
xor U14492 (N_14492,N_9304,N_11671);
or U14493 (N_14493,N_8476,N_11883);
xor U14494 (N_14494,N_8251,N_8213);
and U14495 (N_14495,N_8882,N_10564);
nor U14496 (N_14496,N_8392,N_10956);
nor U14497 (N_14497,N_11022,N_9911);
and U14498 (N_14498,N_11003,N_11796);
xor U14499 (N_14499,N_11609,N_8473);
nand U14500 (N_14500,N_9224,N_9821);
xnor U14501 (N_14501,N_11570,N_8046);
nor U14502 (N_14502,N_11873,N_9928);
nand U14503 (N_14503,N_11184,N_11618);
and U14504 (N_14504,N_11842,N_8969);
or U14505 (N_14505,N_11561,N_8396);
nor U14506 (N_14506,N_10244,N_8368);
and U14507 (N_14507,N_9609,N_10477);
nor U14508 (N_14508,N_10416,N_11994);
or U14509 (N_14509,N_10229,N_11536);
nor U14510 (N_14510,N_11654,N_10468);
or U14511 (N_14511,N_10749,N_8387);
nor U14512 (N_14512,N_9309,N_11363);
and U14513 (N_14513,N_11199,N_9415);
nand U14514 (N_14514,N_10987,N_11096);
nor U14515 (N_14515,N_9585,N_8364);
or U14516 (N_14516,N_8157,N_11679);
nor U14517 (N_14517,N_8273,N_9630);
or U14518 (N_14518,N_8289,N_8585);
and U14519 (N_14519,N_8589,N_10091);
nor U14520 (N_14520,N_10543,N_11517);
xnor U14521 (N_14521,N_10335,N_8256);
nand U14522 (N_14522,N_10086,N_9155);
xor U14523 (N_14523,N_8047,N_8853);
or U14524 (N_14524,N_11092,N_10350);
nor U14525 (N_14525,N_10854,N_11138);
and U14526 (N_14526,N_11249,N_10354);
xor U14527 (N_14527,N_9938,N_11589);
xnor U14528 (N_14528,N_8670,N_11745);
or U14529 (N_14529,N_9180,N_10995);
and U14530 (N_14530,N_10906,N_11282);
xor U14531 (N_14531,N_8165,N_11396);
nand U14532 (N_14532,N_9761,N_10903);
nand U14533 (N_14533,N_8850,N_9398);
xor U14534 (N_14534,N_11064,N_9390);
nand U14535 (N_14535,N_10428,N_10213);
or U14536 (N_14536,N_9475,N_10660);
and U14537 (N_14537,N_9920,N_10679);
xnor U14538 (N_14538,N_9123,N_9006);
xor U14539 (N_14539,N_9065,N_9297);
and U14540 (N_14540,N_9370,N_10164);
xnor U14541 (N_14541,N_10457,N_8203);
nand U14542 (N_14542,N_10086,N_11058);
and U14543 (N_14543,N_9379,N_11619);
or U14544 (N_14544,N_10997,N_9635);
and U14545 (N_14545,N_10187,N_10071);
xor U14546 (N_14546,N_9348,N_9042);
nor U14547 (N_14547,N_9721,N_8789);
nand U14548 (N_14548,N_9942,N_9514);
or U14549 (N_14549,N_10425,N_11165);
and U14550 (N_14550,N_11620,N_8391);
and U14551 (N_14551,N_11909,N_10840);
nand U14552 (N_14552,N_8009,N_8657);
nor U14553 (N_14553,N_11077,N_8649);
or U14554 (N_14554,N_9201,N_8116);
nand U14555 (N_14555,N_8868,N_8073);
xor U14556 (N_14556,N_10447,N_8192);
or U14557 (N_14557,N_8810,N_11512);
and U14558 (N_14558,N_11739,N_11905);
nand U14559 (N_14559,N_10854,N_11062);
nor U14560 (N_14560,N_11214,N_11726);
nor U14561 (N_14561,N_11897,N_10540);
or U14562 (N_14562,N_11007,N_9389);
or U14563 (N_14563,N_8927,N_8177);
nor U14564 (N_14564,N_10119,N_11940);
xor U14565 (N_14565,N_8945,N_11995);
xor U14566 (N_14566,N_9788,N_8356);
or U14567 (N_14567,N_10460,N_10872);
and U14568 (N_14568,N_10492,N_8573);
nand U14569 (N_14569,N_11092,N_8948);
nand U14570 (N_14570,N_10907,N_10722);
and U14571 (N_14571,N_8563,N_10261);
nor U14572 (N_14572,N_11422,N_8703);
nand U14573 (N_14573,N_11405,N_11483);
nand U14574 (N_14574,N_11835,N_9649);
nor U14575 (N_14575,N_9443,N_10773);
or U14576 (N_14576,N_11710,N_9046);
nor U14577 (N_14577,N_11358,N_11140);
and U14578 (N_14578,N_9171,N_11484);
nor U14579 (N_14579,N_10055,N_9831);
or U14580 (N_14580,N_11552,N_9486);
and U14581 (N_14581,N_9595,N_10312);
nand U14582 (N_14582,N_11150,N_9393);
nor U14583 (N_14583,N_11159,N_11535);
nor U14584 (N_14584,N_8333,N_8646);
nand U14585 (N_14585,N_11459,N_10071);
nor U14586 (N_14586,N_11981,N_10705);
nand U14587 (N_14587,N_8297,N_11229);
xnor U14588 (N_14588,N_11219,N_9364);
nor U14589 (N_14589,N_8741,N_8020);
nor U14590 (N_14590,N_11847,N_8394);
xnor U14591 (N_14591,N_11591,N_8966);
and U14592 (N_14592,N_11116,N_9695);
nor U14593 (N_14593,N_11477,N_9053);
xnor U14594 (N_14594,N_10006,N_8912);
xor U14595 (N_14595,N_11211,N_11646);
and U14596 (N_14596,N_10491,N_8213);
nand U14597 (N_14597,N_9567,N_11545);
nand U14598 (N_14598,N_11788,N_9640);
and U14599 (N_14599,N_9142,N_9451);
nor U14600 (N_14600,N_10178,N_10583);
nand U14601 (N_14601,N_8223,N_11165);
and U14602 (N_14602,N_8305,N_11128);
and U14603 (N_14603,N_11516,N_9450);
or U14604 (N_14604,N_11416,N_10855);
xor U14605 (N_14605,N_9079,N_10568);
and U14606 (N_14606,N_8674,N_11035);
or U14607 (N_14607,N_8452,N_10580);
xor U14608 (N_14608,N_10410,N_8821);
or U14609 (N_14609,N_8681,N_11975);
xnor U14610 (N_14610,N_8536,N_8914);
nand U14611 (N_14611,N_11149,N_10939);
nand U14612 (N_14612,N_8648,N_11825);
nor U14613 (N_14613,N_10860,N_11853);
or U14614 (N_14614,N_8296,N_9187);
or U14615 (N_14615,N_8685,N_8426);
and U14616 (N_14616,N_8997,N_9452);
and U14617 (N_14617,N_8659,N_10028);
nand U14618 (N_14618,N_8141,N_10347);
or U14619 (N_14619,N_11613,N_8134);
or U14620 (N_14620,N_8633,N_11644);
nand U14621 (N_14621,N_9002,N_8187);
xnor U14622 (N_14622,N_8380,N_10379);
nand U14623 (N_14623,N_10423,N_11586);
and U14624 (N_14624,N_9560,N_11357);
nand U14625 (N_14625,N_9114,N_9045);
xor U14626 (N_14626,N_9456,N_9432);
nor U14627 (N_14627,N_11144,N_10688);
nor U14628 (N_14628,N_11696,N_9569);
or U14629 (N_14629,N_8160,N_11030);
and U14630 (N_14630,N_10908,N_10565);
xor U14631 (N_14631,N_9495,N_8470);
nor U14632 (N_14632,N_10292,N_9777);
and U14633 (N_14633,N_11945,N_10722);
xor U14634 (N_14634,N_10303,N_10547);
nand U14635 (N_14635,N_9614,N_9387);
xor U14636 (N_14636,N_9968,N_8814);
xnor U14637 (N_14637,N_8158,N_9081);
nand U14638 (N_14638,N_10427,N_10675);
nand U14639 (N_14639,N_9207,N_10193);
or U14640 (N_14640,N_9390,N_10085);
nor U14641 (N_14641,N_8356,N_11503);
nor U14642 (N_14642,N_9098,N_8111);
or U14643 (N_14643,N_9137,N_10905);
and U14644 (N_14644,N_8118,N_11126);
or U14645 (N_14645,N_11380,N_10375);
nor U14646 (N_14646,N_10558,N_10225);
or U14647 (N_14647,N_9446,N_11331);
and U14648 (N_14648,N_8408,N_8440);
and U14649 (N_14649,N_10810,N_8090);
xor U14650 (N_14650,N_9751,N_9272);
and U14651 (N_14651,N_8985,N_9629);
nand U14652 (N_14652,N_11050,N_10989);
nand U14653 (N_14653,N_8037,N_11306);
or U14654 (N_14654,N_8509,N_10825);
nor U14655 (N_14655,N_9828,N_9093);
nand U14656 (N_14656,N_10175,N_9467);
or U14657 (N_14657,N_10376,N_10196);
and U14658 (N_14658,N_10660,N_11342);
xor U14659 (N_14659,N_10083,N_11288);
and U14660 (N_14660,N_8640,N_11083);
nor U14661 (N_14661,N_11857,N_8594);
xor U14662 (N_14662,N_10849,N_8893);
nand U14663 (N_14663,N_9273,N_11883);
nand U14664 (N_14664,N_9466,N_9449);
xor U14665 (N_14665,N_10331,N_9618);
nor U14666 (N_14666,N_8074,N_9648);
nand U14667 (N_14667,N_9716,N_9878);
nor U14668 (N_14668,N_10436,N_9628);
or U14669 (N_14669,N_11427,N_10194);
xor U14670 (N_14670,N_11305,N_8778);
or U14671 (N_14671,N_10952,N_9922);
and U14672 (N_14672,N_11404,N_8405);
nand U14673 (N_14673,N_9601,N_8601);
nor U14674 (N_14674,N_9203,N_11051);
or U14675 (N_14675,N_10501,N_9950);
and U14676 (N_14676,N_9114,N_10960);
and U14677 (N_14677,N_9278,N_9760);
xnor U14678 (N_14678,N_11024,N_11957);
nand U14679 (N_14679,N_11848,N_11603);
or U14680 (N_14680,N_9078,N_9585);
and U14681 (N_14681,N_9836,N_8280);
nand U14682 (N_14682,N_10445,N_9388);
nor U14683 (N_14683,N_10442,N_8963);
xor U14684 (N_14684,N_9952,N_9868);
and U14685 (N_14685,N_10622,N_9848);
nand U14686 (N_14686,N_8047,N_11710);
xnor U14687 (N_14687,N_10683,N_11023);
nand U14688 (N_14688,N_9319,N_10674);
nand U14689 (N_14689,N_9236,N_11599);
nor U14690 (N_14690,N_8534,N_9950);
nor U14691 (N_14691,N_9548,N_9288);
nor U14692 (N_14692,N_10572,N_8796);
xnor U14693 (N_14693,N_8052,N_9053);
xnor U14694 (N_14694,N_10325,N_11888);
or U14695 (N_14695,N_9059,N_9653);
nand U14696 (N_14696,N_8482,N_11812);
nand U14697 (N_14697,N_10552,N_11709);
nand U14698 (N_14698,N_9956,N_11285);
and U14699 (N_14699,N_10556,N_11320);
or U14700 (N_14700,N_10370,N_9662);
nor U14701 (N_14701,N_10612,N_10932);
or U14702 (N_14702,N_8767,N_9131);
or U14703 (N_14703,N_9089,N_9130);
and U14704 (N_14704,N_8972,N_8137);
and U14705 (N_14705,N_9993,N_9933);
nand U14706 (N_14706,N_10569,N_9646);
nand U14707 (N_14707,N_10909,N_10232);
xor U14708 (N_14708,N_10160,N_8695);
xnor U14709 (N_14709,N_8930,N_11260);
nand U14710 (N_14710,N_8272,N_11653);
and U14711 (N_14711,N_8263,N_9878);
xor U14712 (N_14712,N_8106,N_9274);
xor U14713 (N_14713,N_8728,N_8223);
nand U14714 (N_14714,N_11485,N_10363);
xor U14715 (N_14715,N_9222,N_11803);
and U14716 (N_14716,N_8362,N_11493);
or U14717 (N_14717,N_10910,N_8688);
nand U14718 (N_14718,N_11916,N_10323);
or U14719 (N_14719,N_8827,N_11591);
xor U14720 (N_14720,N_11162,N_9939);
nor U14721 (N_14721,N_8668,N_10267);
nand U14722 (N_14722,N_8258,N_11094);
xnor U14723 (N_14723,N_11704,N_9164);
nand U14724 (N_14724,N_11698,N_11772);
nor U14725 (N_14725,N_11254,N_9064);
nor U14726 (N_14726,N_10983,N_9790);
or U14727 (N_14727,N_8680,N_10794);
nand U14728 (N_14728,N_10701,N_9041);
nor U14729 (N_14729,N_9065,N_10371);
nor U14730 (N_14730,N_10493,N_11526);
or U14731 (N_14731,N_10974,N_8285);
nor U14732 (N_14732,N_10983,N_9714);
and U14733 (N_14733,N_9992,N_9894);
or U14734 (N_14734,N_11437,N_9501);
and U14735 (N_14735,N_10142,N_10096);
and U14736 (N_14736,N_9955,N_9974);
nor U14737 (N_14737,N_11297,N_8931);
or U14738 (N_14738,N_10336,N_8207);
nor U14739 (N_14739,N_9384,N_8205);
and U14740 (N_14740,N_8984,N_10344);
nand U14741 (N_14741,N_8086,N_11476);
nand U14742 (N_14742,N_10735,N_11671);
xor U14743 (N_14743,N_10322,N_10558);
nand U14744 (N_14744,N_8981,N_9898);
xor U14745 (N_14745,N_8901,N_10962);
and U14746 (N_14746,N_9031,N_9034);
and U14747 (N_14747,N_8227,N_10415);
or U14748 (N_14748,N_10636,N_8644);
nor U14749 (N_14749,N_9977,N_8063);
nor U14750 (N_14750,N_8277,N_10201);
nand U14751 (N_14751,N_8596,N_10715);
nand U14752 (N_14752,N_10193,N_8768);
xnor U14753 (N_14753,N_11217,N_10492);
nor U14754 (N_14754,N_8191,N_9916);
or U14755 (N_14755,N_8007,N_9265);
nand U14756 (N_14756,N_11929,N_8888);
nand U14757 (N_14757,N_10806,N_9701);
and U14758 (N_14758,N_9034,N_10141);
nor U14759 (N_14759,N_11124,N_8086);
nand U14760 (N_14760,N_10343,N_9255);
or U14761 (N_14761,N_8182,N_8904);
xnor U14762 (N_14762,N_9547,N_11623);
xnor U14763 (N_14763,N_9513,N_9755);
nor U14764 (N_14764,N_8008,N_10844);
nand U14765 (N_14765,N_11165,N_9199);
and U14766 (N_14766,N_10684,N_10773);
or U14767 (N_14767,N_9536,N_9439);
nand U14768 (N_14768,N_9214,N_10396);
nor U14769 (N_14769,N_10852,N_10846);
or U14770 (N_14770,N_8298,N_11227);
xnor U14771 (N_14771,N_9588,N_9075);
nand U14772 (N_14772,N_8056,N_10810);
nand U14773 (N_14773,N_11156,N_10880);
nand U14774 (N_14774,N_11232,N_11934);
or U14775 (N_14775,N_10937,N_9223);
and U14776 (N_14776,N_8118,N_8653);
nand U14777 (N_14777,N_11657,N_9554);
and U14778 (N_14778,N_9708,N_11757);
nand U14779 (N_14779,N_8251,N_8093);
or U14780 (N_14780,N_10208,N_10034);
xor U14781 (N_14781,N_9282,N_9205);
nor U14782 (N_14782,N_11717,N_9076);
or U14783 (N_14783,N_9684,N_9698);
and U14784 (N_14784,N_9174,N_10952);
or U14785 (N_14785,N_8144,N_8792);
or U14786 (N_14786,N_8176,N_10349);
nor U14787 (N_14787,N_8260,N_10210);
or U14788 (N_14788,N_11082,N_10267);
or U14789 (N_14789,N_10242,N_11703);
and U14790 (N_14790,N_10202,N_10817);
or U14791 (N_14791,N_11983,N_11248);
or U14792 (N_14792,N_9417,N_11057);
xnor U14793 (N_14793,N_10560,N_8697);
or U14794 (N_14794,N_9920,N_9355);
nand U14795 (N_14795,N_8453,N_11387);
nand U14796 (N_14796,N_10381,N_10841);
xnor U14797 (N_14797,N_9939,N_10688);
xnor U14798 (N_14798,N_10296,N_8370);
nand U14799 (N_14799,N_11752,N_9780);
xor U14800 (N_14800,N_11054,N_11635);
xor U14801 (N_14801,N_10441,N_10692);
and U14802 (N_14802,N_10110,N_10682);
or U14803 (N_14803,N_10730,N_8691);
or U14804 (N_14804,N_11833,N_10040);
xor U14805 (N_14805,N_11128,N_11978);
or U14806 (N_14806,N_11810,N_10332);
nor U14807 (N_14807,N_9557,N_11685);
or U14808 (N_14808,N_9996,N_10112);
xor U14809 (N_14809,N_11750,N_10589);
nand U14810 (N_14810,N_8292,N_9076);
and U14811 (N_14811,N_11307,N_11785);
or U14812 (N_14812,N_9806,N_10975);
nor U14813 (N_14813,N_8119,N_8570);
xor U14814 (N_14814,N_10458,N_9089);
and U14815 (N_14815,N_11393,N_9196);
or U14816 (N_14816,N_9275,N_9069);
or U14817 (N_14817,N_10762,N_8261);
nand U14818 (N_14818,N_8361,N_11734);
nand U14819 (N_14819,N_9462,N_9734);
nor U14820 (N_14820,N_8038,N_8591);
nor U14821 (N_14821,N_10727,N_9293);
nor U14822 (N_14822,N_10017,N_9302);
and U14823 (N_14823,N_8869,N_10946);
or U14824 (N_14824,N_9130,N_11209);
or U14825 (N_14825,N_9808,N_8481);
nand U14826 (N_14826,N_8907,N_9103);
xor U14827 (N_14827,N_8523,N_10138);
nor U14828 (N_14828,N_8874,N_11304);
xor U14829 (N_14829,N_11557,N_11098);
and U14830 (N_14830,N_9608,N_11693);
nor U14831 (N_14831,N_11667,N_11539);
and U14832 (N_14832,N_10245,N_11951);
and U14833 (N_14833,N_10187,N_9798);
nor U14834 (N_14834,N_8910,N_9646);
nor U14835 (N_14835,N_9462,N_11568);
and U14836 (N_14836,N_10636,N_10927);
nand U14837 (N_14837,N_10528,N_11085);
and U14838 (N_14838,N_9818,N_8110);
or U14839 (N_14839,N_8397,N_8511);
or U14840 (N_14840,N_10484,N_9377);
xnor U14841 (N_14841,N_11231,N_11742);
and U14842 (N_14842,N_10069,N_11774);
nand U14843 (N_14843,N_11010,N_8428);
xor U14844 (N_14844,N_11538,N_8018);
or U14845 (N_14845,N_10330,N_8764);
and U14846 (N_14846,N_11791,N_11113);
or U14847 (N_14847,N_8527,N_8462);
and U14848 (N_14848,N_11566,N_10296);
xor U14849 (N_14849,N_9491,N_10728);
nor U14850 (N_14850,N_11114,N_8094);
or U14851 (N_14851,N_11365,N_8797);
nor U14852 (N_14852,N_8337,N_9851);
xor U14853 (N_14853,N_8371,N_9002);
and U14854 (N_14854,N_10752,N_9165);
nor U14855 (N_14855,N_11081,N_10769);
xnor U14856 (N_14856,N_8287,N_9549);
xor U14857 (N_14857,N_9932,N_11776);
and U14858 (N_14858,N_11894,N_8682);
or U14859 (N_14859,N_9484,N_9707);
nor U14860 (N_14860,N_8309,N_8455);
nor U14861 (N_14861,N_11541,N_11189);
nor U14862 (N_14862,N_11091,N_11029);
nand U14863 (N_14863,N_8192,N_10238);
nand U14864 (N_14864,N_11846,N_8973);
or U14865 (N_14865,N_9434,N_9238);
nand U14866 (N_14866,N_8401,N_10568);
and U14867 (N_14867,N_9924,N_11371);
and U14868 (N_14868,N_11902,N_11909);
xor U14869 (N_14869,N_9146,N_11727);
or U14870 (N_14870,N_11538,N_8417);
nor U14871 (N_14871,N_9075,N_10292);
nand U14872 (N_14872,N_9487,N_9661);
xor U14873 (N_14873,N_9423,N_8308);
nor U14874 (N_14874,N_10166,N_10114);
and U14875 (N_14875,N_8995,N_10991);
or U14876 (N_14876,N_8861,N_8931);
and U14877 (N_14877,N_10477,N_9263);
nand U14878 (N_14878,N_8279,N_10462);
and U14879 (N_14879,N_9316,N_10597);
nor U14880 (N_14880,N_9333,N_8573);
nand U14881 (N_14881,N_8359,N_9441);
nor U14882 (N_14882,N_10380,N_10130);
or U14883 (N_14883,N_8553,N_9625);
nand U14884 (N_14884,N_8894,N_9900);
xor U14885 (N_14885,N_8842,N_10984);
and U14886 (N_14886,N_8846,N_8362);
xor U14887 (N_14887,N_10107,N_10497);
and U14888 (N_14888,N_11667,N_9360);
nor U14889 (N_14889,N_9619,N_10388);
or U14890 (N_14890,N_11419,N_9309);
nand U14891 (N_14891,N_9994,N_8900);
nand U14892 (N_14892,N_11670,N_9799);
xor U14893 (N_14893,N_11286,N_11437);
or U14894 (N_14894,N_10774,N_11036);
nand U14895 (N_14895,N_8718,N_11845);
or U14896 (N_14896,N_9568,N_9505);
or U14897 (N_14897,N_11413,N_10448);
xnor U14898 (N_14898,N_8831,N_8021);
or U14899 (N_14899,N_10868,N_8868);
or U14900 (N_14900,N_8776,N_9742);
nor U14901 (N_14901,N_8361,N_10450);
or U14902 (N_14902,N_9608,N_11694);
nor U14903 (N_14903,N_11502,N_8540);
nor U14904 (N_14904,N_8102,N_11633);
nor U14905 (N_14905,N_9182,N_11026);
or U14906 (N_14906,N_10690,N_10072);
nand U14907 (N_14907,N_10033,N_9339);
nor U14908 (N_14908,N_10637,N_11474);
nand U14909 (N_14909,N_9954,N_10871);
or U14910 (N_14910,N_11135,N_10221);
or U14911 (N_14911,N_8201,N_8370);
or U14912 (N_14912,N_10657,N_11026);
and U14913 (N_14913,N_8935,N_8990);
or U14914 (N_14914,N_8549,N_11347);
or U14915 (N_14915,N_9446,N_11897);
nor U14916 (N_14916,N_11169,N_9961);
and U14917 (N_14917,N_9052,N_10816);
xnor U14918 (N_14918,N_8471,N_9118);
nand U14919 (N_14919,N_9967,N_9331);
nand U14920 (N_14920,N_10508,N_11777);
nor U14921 (N_14921,N_8146,N_8195);
nand U14922 (N_14922,N_9209,N_11173);
nor U14923 (N_14923,N_8813,N_8161);
nand U14924 (N_14924,N_11552,N_11120);
and U14925 (N_14925,N_11569,N_10377);
nor U14926 (N_14926,N_11814,N_8462);
and U14927 (N_14927,N_10765,N_10011);
nand U14928 (N_14928,N_11083,N_11933);
or U14929 (N_14929,N_9197,N_11230);
nand U14930 (N_14930,N_10301,N_11581);
xnor U14931 (N_14931,N_9985,N_8524);
or U14932 (N_14932,N_11464,N_11245);
and U14933 (N_14933,N_10799,N_11975);
and U14934 (N_14934,N_10048,N_11474);
nand U14935 (N_14935,N_8768,N_8100);
or U14936 (N_14936,N_10836,N_9838);
and U14937 (N_14937,N_10854,N_9753);
and U14938 (N_14938,N_10792,N_9049);
or U14939 (N_14939,N_10205,N_11258);
nor U14940 (N_14940,N_10554,N_8999);
or U14941 (N_14941,N_11460,N_11782);
nand U14942 (N_14942,N_10492,N_11122);
or U14943 (N_14943,N_11986,N_10152);
or U14944 (N_14944,N_9619,N_11160);
or U14945 (N_14945,N_11961,N_9502);
and U14946 (N_14946,N_11899,N_10542);
nor U14947 (N_14947,N_9768,N_9088);
and U14948 (N_14948,N_8853,N_10673);
nor U14949 (N_14949,N_9052,N_9569);
and U14950 (N_14950,N_11430,N_11744);
xor U14951 (N_14951,N_11345,N_8124);
xor U14952 (N_14952,N_9002,N_9864);
and U14953 (N_14953,N_11145,N_11730);
xnor U14954 (N_14954,N_11011,N_9407);
or U14955 (N_14955,N_8667,N_9510);
xor U14956 (N_14956,N_11848,N_9862);
and U14957 (N_14957,N_8948,N_11642);
and U14958 (N_14958,N_8891,N_10247);
nand U14959 (N_14959,N_11433,N_11350);
or U14960 (N_14960,N_11836,N_11395);
and U14961 (N_14961,N_8866,N_10036);
nand U14962 (N_14962,N_10587,N_10005);
xor U14963 (N_14963,N_10020,N_9506);
xnor U14964 (N_14964,N_8920,N_11585);
xor U14965 (N_14965,N_8861,N_8587);
or U14966 (N_14966,N_8164,N_8930);
nand U14967 (N_14967,N_11128,N_9745);
and U14968 (N_14968,N_8421,N_11938);
nand U14969 (N_14969,N_9118,N_9505);
and U14970 (N_14970,N_10768,N_9189);
xor U14971 (N_14971,N_11413,N_10282);
nor U14972 (N_14972,N_10954,N_11317);
or U14973 (N_14973,N_8605,N_11620);
xor U14974 (N_14974,N_10714,N_10630);
and U14975 (N_14975,N_10696,N_11723);
and U14976 (N_14976,N_11044,N_8805);
nand U14977 (N_14977,N_8938,N_9978);
nor U14978 (N_14978,N_8373,N_11805);
or U14979 (N_14979,N_11348,N_8966);
nand U14980 (N_14980,N_11312,N_10043);
nor U14981 (N_14981,N_9540,N_11815);
nor U14982 (N_14982,N_8567,N_9471);
xnor U14983 (N_14983,N_11863,N_10853);
nand U14984 (N_14984,N_9372,N_11216);
xor U14985 (N_14985,N_10783,N_11579);
xnor U14986 (N_14986,N_9431,N_9758);
and U14987 (N_14987,N_8429,N_11085);
nand U14988 (N_14988,N_8382,N_9035);
xnor U14989 (N_14989,N_8544,N_8550);
or U14990 (N_14990,N_9165,N_9448);
nor U14991 (N_14991,N_10939,N_11313);
xor U14992 (N_14992,N_9067,N_9142);
nor U14993 (N_14993,N_8232,N_9463);
or U14994 (N_14994,N_11203,N_10359);
or U14995 (N_14995,N_8609,N_8652);
and U14996 (N_14996,N_11368,N_11116);
nor U14997 (N_14997,N_10904,N_10491);
nor U14998 (N_14998,N_8341,N_10816);
and U14999 (N_14999,N_9137,N_8324);
or U15000 (N_15000,N_9277,N_9178);
and U15001 (N_15001,N_11775,N_10498);
nand U15002 (N_15002,N_9080,N_9855);
and U15003 (N_15003,N_9469,N_11705);
nor U15004 (N_15004,N_9646,N_11357);
nand U15005 (N_15005,N_11103,N_10284);
or U15006 (N_15006,N_9310,N_10939);
nor U15007 (N_15007,N_11906,N_9662);
nand U15008 (N_15008,N_9779,N_8916);
nand U15009 (N_15009,N_10409,N_9254);
or U15010 (N_15010,N_8445,N_9792);
xnor U15011 (N_15011,N_10764,N_9362);
xor U15012 (N_15012,N_8088,N_9687);
nand U15013 (N_15013,N_11230,N_11587);
nor U15014 (N_15014,N_9893,N_11970);
nor U15015 (N_15015,N_8516,N_10310);
xor U15016 (N_15016,N_8619,N_9619);
or U15017 (N_15017,N_11848,N_9459);
and U15018 (N_15018,N_8938,N_8359);
or U15019 (N_15019,N_9911,N_11118);
nor U15020 (N_15020,N_9032,N_9279);
nor U15021 (N_15021,N_11284,N_9620);
nor U15022 (N_15022,N_9585,N_8832);
or U15023 (N_15023,N_8052,N_11324);
nor U15024 (N_15024,N_9864,N_9934);
nor U15025 (N_15025,N_11309,N_8780);
xor U15026 (N_15026,N_9588,N_11230);
xnor U15027 (N_15027,N_10033,N_11509);
nand U15028 (N_15028,N_8835,N_8905);
xor U15029 (N_15029,N_9206,N_8502);
xnor U15030 (N_15030,N_8001,N_10662);
and U15031 (N_15031,N_11248,N_10392);
nand U15032 (N_15032,N_11598,N_9521);
or U15033 (N_15033,N_11337,N_10546);
nor U15034 (N_15034,N_10078,N_9372);
and U15035 (N_15035,N_10956,N_11468);
or U15036 (N_15036,N_8614,N_9840);
xor U15037 (N_15037,N_9556,N_10773);
nor U15038 (N_15038,N_11233,N_10078);
and U15039 (N_15039,N_9688,N_11650);
nand U15040 (N_15040,N_8978,N_11111);
nor U15041 (N_15041,N_8724,N_10120);
and U15042 (N_15042,N_10520,N_11412);
nand U15043 (N_15043,N_8954,N_8529);
xor U15044 (N_15044,N_8735,N_9195);
nand U15045 (N_15045,N_10522,N_11549);
nand U15046 (N_15046,N_8101,N_8265);
nor U15047 (N_15047,N_8561,N_8062);
nor U15048 (N_15048,N_10317,N_11040);
nor U15049 (N_15049,N_9149,N_9423);
nor U15050 (N_15050,N_10120,N_11995);
or U15051 (N_15051,N_8429,N_9428);
nand U15052 (N_15052,N_11072,N_8507);
nor U15053 (N_15053,N_8950,N_9092);
nor U15054 (N_15054,N_11248,N_9619);
nor U15055 (N_15055,N_8061,N_10323);
xor U15056 (N_15056,N_10718,N_11476);
or U15057 (N_15057,N_9712,N_8127);
nand U15058 (N_15058,N_10635,N_11122);
and U15059 (N_15059,N_8551,N_10011);
and U15060 (N_15060,N_11097,N_10720);
nor U15061 (N_15061,N_9446,N_8295);
xnor U15062 (N_15062,N_8710,N_11727);
nand U15063 (N_15063,N_11058,N_11574);
xnor U15064 (N_15064,N_8328,N_9992);
nand U15065 (N_15065,N_8457,N_9904);
and U15066 (N_15066,N_11004,N_10307);
xnor U15067 (N_15067,N_9473,N_8222);
nand U15068 (N_15068,N_8941,N_11180);
nand U15069 (N_15069,N_9330,N_10402);
xor U15070 (N_15070,N_10122,N_8159);
or U15071 (N_15071,N_9119,N_10968);
or U15072 (N_15072,N_10326,N_11167);
xor U15073 (N_15073,N_8624,N_8036);
nor U15074 (N_15074,N_11978,N_8242);
nor U15075 (N_15075,N_8917,N_9709);
nor U15076 (N_15076,N_10494,N_8592);
nor U15077 (N_15077,N_11249,N_8779);
and U15078 (N_15078,N_8933,N_9868);
xnor U15079 (N_15079,N_8302,N_11940);
xnor U15080 (N_15080,N_9530,N_9459);
and U15081 (N_15081,N_8523,N_11502);
nor U15082 (N_15082,N_10934,N_10884);
nand U15083 (N_15083,N_10987,N_8173);
xor U15084 (N_15084,N_10652,N_10469);
and U15085 (N_15085,N_9868,N_9657);
or U15086 (N_15086,N_10782,N_8894);
and U15087 (N_15087,N_10849,N_8729);
nor U15088 (N_15088,N_8379,N_10556);
xnor U15089 (N_15089,N_11648,N_11864);
nor U15090 (N_15090,N_11593,N_9785);
nand U15091 (N_15091,N_8014,N_10475);
nand U15092 (N_15092,N_9057,N_9730);
or U15093 (N_15093,N_8078,N_11384);
nor U15094 (N_15094,N_8532,N_11799);
nor U15095 (N_15095,N_8590,N_11248);
nand U15096 (N_15096,N_10642,N_8760);
nor U15097 (N_15097,N_10235,N_10619);
nor U15098 (N_15098,N_9078,N_9193);
or U15099 (N_15099,N_11208,N_10186);
nand U15100 (N_15100,N_9640,N_11743);
or U15101 (N_15101,N_8402,N_11322);
and U15102 (N_15102,N_8861,N_10028);
and U15103 (N_15103,N_9471,N_8104);
nand U15104 (N_15104,N_11838,N_11699);
xnor U15105 (N_15105,N_11716,N_8535);
xor U15106 (N_15106,N_9038,N_9441);
xnor U15107 (N_15107,N_9916,N_8642);
xor U15108 (N_15108,N_11676,N_10996);
xnor U15109 (N_15109,N_9617,N_8294);
and U15110 (N_15110,N_8513,N_9542);
and U15111 (N_15111,N_9776,N_10924);
nor U15112 (N_15112,N_11311,N_9754);
nor U15113 (N_15113,N_10552,N_8326);
and U15114 (N_15114,N_9853,N_8227);
and U15115 (N_15115,N_9242,N_8350);
nor U15116 (N_15116,N_10324,N_10598);
nor U15117 (N_15117,N_8517,N_11351);
and U15118 (N_15118,N_9650,N_9580);
and U15119 (N_15119,N_10340,N_8486);
or U15120 (N_15120,N_10795,N_9056);
nor U15121 (N_15121,N_11636,N_9972);
nand U15122 (N_15122,N_11860,N_8919);
nor U15123 (N_15123,N_11882,N_11991);
nor U15124 (N_15124,N_11037,N_9206);
and U15125 (N_15125,N_11950,N_9681);
and U15126 (N_15126,N_9525,N_10062);
xnor U15127 (N_15127,N_8370,N_10137);
nand U15128 (N_15128,N_10279,N_8987);
and U15129 (N_15129,N_10504,N_9514);
nor U15130 (N_15130,N_8394,N_11895);
and U15131 (N_15131,N_8362,N_8149);
xor U15132 (N_15132,N_9335,N_9122);
and U15133 (N_15133,N_9803,N_9596);
nand U15134 (N_15134,N_8888,N_9977);
or U15135 (N_15135,N_9366,N_9817);
or U15136 (N_15136,N_8985,N_10909);
nor U15137 (N_15137,N_10326,N_8942);
nor U15138 (N_15138,N_11907,N_10943);
nand U15139 (N_15139,N_10126,N_11973);
nand U15140 (N_15140,N_9721,N_10509);
or U15141 (N_15141,N_9221,N_9138);
and U15142 (N_15142,N_9133,N_10835);
nand U15143 (N_15143,N_11881,N_9026);
and U15144 (N_15144,N_11938,N_8804);
xor U15145 (N_15145,N_10500,N_9982);
and U15146 (N_15146,N_10604,N_8129);
xnor U15147 (N_15147,N_8004,N_9670);
nand U15148 (N_15148,N_10756,N_11479);
xnor U15149 (N_15149,N_10797,N_8954);
and U15150 (N_15150,N_10619,N_11179);
nor U15151 (N_15151,N_8507,N_8004);
nand U15152 (N_15152,N_10844,N_11055);
or U15153 (N_15153,N_9031,N_10600);
nand U15154 (N_15154,N_9780,N_9083);
or U15155 (N_15155,N_9941,N_10185);
or U15156 (N_15156,N_9994,N_8356);
or U15157 (N_15157,N_11800,N_8600);
nor U15158 (N_15158,N_11285,N_8267);
and U15159 (N_15159,N_8224,N_10887);
or U15160 (N_15160,N_8551,N_11862);
nor U15161 (N_15161,N_8424,N_11343);
and U15162 (N_15162,N_9145,N_9992);
xnor U15163 (N_15163,N_9184,N_8464);
nand U15164 (N_15164,N_11277,N_8562);
nand U15165 (N_15165,N_8185,N_8353);
nand U15166 (N_15166,N_10094,N_11726);
and U15167 (N_15167,N_9493,N_8122);
and U15168 (N_15168,N_9270,N_10262);
nor U15169 (N_15169,N_8370,N_9087);
nand U15170 (N_15170,N_8345,N_10865);
or U15171 (N_15171,N_9414,N_8711);
and U15172 (N_15172,N_9079,N_11476);
nand U15173 (N_15173,N_9624,N_11233);
xnor U15174 (N_15174,N_11334,N_11534);
xnor U15175 (N_15175,N_9274,N_8660);
or U15176 (N_15176,N_9395,N_8624);
nand U15177 (N_15177,N_10160,N_8987);
or U15178 (N_15178,N_9779,N_8047);
nor U15179 (N_15179,N_11881,N_10871);
and U15180 (N_15180,N_11241,N_9529);
xor U15181 (N_15181,N_8424,N_9789);
or U15182 (N_15182,N_8395,N_11189);
nand U15183 (N_15183,N_11443,N_8754);
xor U15184 (N_15184,N_8347,N_11169);
or U15185 (N_15185,N_8271,N_8623);
and U15186 (N_15186,N_11107,N_8301);
nand U15187 (N_15187,N_8968,N_8471);
nor U15188 (N_15188,N_10821,N_10117);
xor U15189 (N_15189,N_11392,N_8340);
xor U15190 (N_15190,N_11049,N_9967);
xnor U15191 (N_15191,N_9953,N_8220);
and U15192 (N_15192,N_11776,N_10564);
nand U15193 (N_15193,N_8548,N_8141);
and U15194 (N_15194,N_8563,N_10170);
nand U15195 (N_15195,N_11641,N_10687);
nand U15196 (N_15196,N_10645,N_9923);
or U15197 (N_15197,N_8457,N_8093);
or U15198 (N_15198,N_11639,N_9726);
and U15199 (N_15199,N_8213,N_8152);
or U15200 (N_15200,N_10064,N_11722);
and U15201 (N_15201,N_9025,N_8164);
and U15202 (N_15202,N_10893,N_11226);
nand U15203 (N_15203,N_8345,N_8196);
nand U15204 (N_15204,N_11187,N_8350);
and U15205 (N_15205,N_9464,N_11677);
xor U15206 (N_15206,N_9721,N_9214);
xor U15207 (N_15207,N_8103,N_8773);
xor U15208 (N_15208,N_10093,N_8888);
xnor U15209 (N_15209,N_10723,N_8075);
xor U15210 (N_15210,N_9539,N_10341);
xor U15211 (N_15211,N_11965,N_8451);
nor U15212 (N_15212,N_11603,N_9941);
or U15213 (N_15213,N_11852,N_9331);
nand U15214 (N_15214,N_10523,N_9674);
or U15215 (N_15215,N_9180,N_9305);
nor U15216 (N_15216,N_8120,N_11792);
nor U15217 (N_15217,N_8069,N_10545);
or U15218 (N_15218,N_8782,N_9237);
xnor U15219 (N_15219,N_9607,N_8541);
or U15220 (N_15220,N_9319,N_11369);
nand U15221 (N_15221,N_11169,N_8846);
nand U15222 (N_15222,N_8746,N_8679);
or U15223 (N_15223,N_8399,N_8835);
nand U15224 (N_15224,N_9347,N_9793);
nor U15225 (N_15225,N_8440,N_9504);
or U15226 (N_15226,N_11684,N_11806);
nor U15227 (N_15227,N_11542,N_11445);
nor U15228 (N_15228,N_11463,N_10610);
and U15229 (N_15229,N_9332,N_11842);
and U15230 (N_15230,N_8981,N_10737);
or U15231 (N_15231,N_9181,N_8790);
and U15232 (N_15232,N_8546,N_9633);
xor U15233 (N_15233,N_11594,N_10436);
nand U15234 (N_15234,N_11520,N_9937);
xnor U15235 (N_15235,N_9696,N_10586);
or U15236 (N_15236,N_9250,N_11849);
nor U15237 (N_15237,N_11980,N_8154);
nor U15238 (N_15238,N_9665,N_9792);
xor U15239 (N_15239,N_9731,N_11222);
nor U15240 (N_15240,N_11469,N_9263);
nand U15241 (N_15241,N_9998,N_9419);
and U15242 (N_15242,N_9877,N_8553);
xnor U15243 (N_15243,N_9963,N_10876);
or U15244 (N_15244,N_8706,N_11862);
nor U15245 (N_15245,N_8212,N_10262);
or U15246 (N_15246,N_10974,N_8855);
xnor U15247 (N_15247,N_10327,N_9079);
nor U15248 (N_15248,N_8963,N_11950);
nand U15249 (N_15249,N_10464,N_9244);
and U15250 (N_15250,N_11371,N_10623);
xnor U15251 (N_15251,N_9404,N_10177);
or U15252 (N_15252,N_10774,N_9500);
xnor U15253 (N_15253,N_8285,N_9585);
and U15254 (N_15254,N_9358,N_9942);
xnor U15255 (N_15255,N_9688,N_11623);
xnor U15256 (N_15256,N_11031,N_10717);
nor U15257 (N_15257,N_9787,N_8085);
or U15258 (N_15258,N_9230,N_9982);
xnor U15259 (N_15259,N_9015,N_11040);
nand U15260 (N_15260,N_8692,N_9915);
or U15261 (N_15261,N_10982,N_11630);
and U15262 (N_15262,N_11967,N_8145);
nand U15263 (N_15263,N_8531,N_10590);
xnor U15264 (N_15264,N_9035,N_8139);
xnor U15265 (N_15265,N_10231,N_10970);
xor U15266 (N_15266,N_9308,N_10874);
xor U15267 (N_15267,N_11454,N_11132);
xnor U15268 (N_15268,N_9920,N_9249);
nor U15269 (N_15269,N_11596,N_11615);
nor U15270 (N_15270,N_8322,N_8435);
and U15271 (N_15271,N_8841,N_8922);
xor U15272 (N_15272,N_11853,N_8428);
xor U15273 (N_15273,N_10783,N_9941);
or U15274 (N_15274,N_11786,N_9125);
nand U15275 (N_15275,N_9076,N_8446);
nor U15276 (N_15276,N_11917,N_11169);
xnor U15277 (N_15277,N_10093,N_8550);
or U15278 (N_15278,N_8010,N_10506);
or U15279 (N_15279,N_10310,N_10120);
and U15280 (N_15280,N_8690,N_11466);
and U15281 (N_15281,N_9909,N_9088);
xor U15282 (N_15282,N_10995,N_11532);
xor U15283 (N_15283,N_10761,N_10521);
nand U15284 (N_15284,N_11316,N_8708);
nand U15285 (N_15285,N_10697,N_8128);
nand U15286 (N_15286,N_9271,N_8954);
nor U15287 (N_15287,N_11527,N_11517);
or U15288 (N_15288,N_8856,N_10485);
nor U15289 (N_15289,N_8440,N_9157);
nor U15290 (N_15290,N_11821,N_11115);
or U15291 (N_15291,N_9044,N_11787);
and U15292 (N_15292,N_10529,N_9999);
nand U15293 (N_15293,N_9926,N_8566);
nor U15294 (N_15294,N_9826,N_11601);
nor U15295 (N_15295,N_11103,N_9045);
xnor U15296 (N_15296,N_11641,N_10822);
nand U15297 (N_15297,N_10492,N_11917);
nor U15298 (N_15298,N_10546,N_8311);
xnor U15299 (N_15299,N_8913,N_11619);
nor U15300 (N_15300,N_9570,N_8806);
xnor U15301 (N_15301,N_10270,N_9696);
xnor U15302 (N_15302,N_11345,N_9283);
nand U15303 (N_15303,N_10619,N_9479);
xnor U15304 (N_15304,N_8458,N_11622);
xor U15305 (N_15305,N_9216,N_10069);
or U15306 (N_15306,N_11172,N_9803);
or U15307 (N_15307,N_10350,N_9434);
and U15308 (N_15308,N_8157,N_11919);
nor U15309 (N_15309,N_9317,N_8856);
xnor U15310 (N_15310,N_11573,N_8620);
and U15311 (N_15311,N_9542,N_9035);
xor U15312 (N_15312,N_9949,N_9077);
xor U15313 (N_15313,N_10183,N_9993);
xnor U15314 (N_15314,N_9855,N_10510);
nand U15315 (N_15315,N_10956,N_9979);
xnor U15316 (N_15316,N_8131,N_8140);
xor U15317 (N_15317,N_10846,N_9058);
or U15318 (N_15318,N_9269,N_10709);
nand U15319 (N_15319,N_8001,N_8290);
or U15320 (N_15320,N_9056,N_11751);
xnor U15321 (N_15321,N_11752,N_9218);
or U15322 (N_15322,N_8143,N_10460);
and U15323 (N_15323,N_10196,N_10119);
nand U15324 (N_15324,N_11758,N_10375);
or U15325 (N_15325,N_9117,N_10371);
xnor U15326 (N_15326,N_9678,N_9383);
nand U15327 (N_15327,N_10052,N_9054);
xor U15328 (N_15328,N_9549,N_9049);
and U15329 (N_15329,N_11757,N_10638);
nor U15330 (N_15330,N_10606,N_10974);
nor U15331 (N_15331,N_9317,N_9093);
and U15332 (N_15332,N_10093,N_10997);
nand U15333 (N_15333,N_11542,N_9541);
or U15334 (N_15334,N_8889,N_9663);
or U15335 (N_15335,N_10096,N_9795);
and U15336 (N_15336,N_9722,N_8428);
and U15337 (N_15337,N_10732,N_8361);
xor U15338 (N_15338,N_8867,N_9654);
and U15339 (N_15339,N_10066,N_8643);
xor U15340 (N_15340,N_9425,N_9377);
or U15341 (N_15341,N_10102,N_11503);
and U15342 (N_15342,N_11213,N_8450);
or U15343 (N_15343,N_11789,N_11384);
xnor U15344 (N_15344,N_10660,N_9997);
xor U15345 (N_15345,N_9228,N_8114);
or U15346 (N_15346,N_10950,N_8800);
or U15347 (N_15347,N_10908,N_9518);
and U15348 (N_15348,N_8238,N_9796);
xnor U15349 (N_15349,N_11290,N_10763);
xor U15350 (N_15350,N_11167,N_11091);
nand U15351 (N_15351,N_8806,N_11837);
xnor U15352 (N_15352,N_10664,N_10476);
xnor U15353 (N_15353,N_11637,N_9130);
nor U15354 (N_15354,N_10217,N_11266);
xnor U15355 (N_15355,N_8872,N_8722);
xnor U15356 (N_15356,N_9826,N_10324);
and U15357 (N_15357,N_8246,N_10623);
or U15358 (N_15358,N_9424,N_9677);
or U15359 (N_15359,N_9725,N_8482);
nand U15360 (N_15360,N_8577,N_8900);
nor U15361 (N_15361,N_10152,N_9794);
or U15362 (N_15362,N_11278,N_9225);
nand U15363 (N_15363,N_8829,N_10037);
and U15364 (N_15364,N_11328,N_10172);
nand U15365 (N_15365,N_8407,N_8690);
or U15366 (N_15366,N_8511,N_11417);
nor U15367 (N_15367,N_11243,N_10621);
nand U15368 (N_15368,N_9550,N_11181);
and U15369 (N_15369,N_11642,N_8161);
nand U15370 (N_15370,N_8297,N_10682);
xor U15371 (N_15371,N_8579,N_11230);
nor U15372 (N_15372,N_10165,N_10141);
nand U15373 (N_15373,N_8637,N_9800);
and U15374 (N_15374,N_8242,N_9437);
xnor U15375 (N_15375,N_11513,N_11973);
nor U15376 (N_15376,N_8833,N_11673);
and U15377 (N_15377,N_11581,N_10076);
nor U15378 (N_15378,N_10174,N_8455);
or U15379 (N_15379,N_10742,N_9831);
and U15380 (N_15380,N_11221,N_10043);
xnor U15381 (N_15381,N_8092,N_11949);
xor U15382 (N_15382,N_8316,N_11003);
and U15383 (N_15383,N_10887,N_9999);
nand U15384 (N_15384,N_11130,N_8663);
nor U15385 (N_15385,N_11406,N_10559);
xor U15386 (N_15386,N_11687,N_10555);
or U15387 (N_15387,N_10126,N_9308);
nor U15388 (N_15388,N_9688,N_9942);
nor U15389 (N_15389,N_11778,N_9851);
nand U15390 (N_15390,N_8877,N_9028);
xnor U15391 (N_15391,N_11966,N_11305);
nor U15392 (N_15392,N_11448,N_10351);
and U15393 (N_15393,N_9198,N_8446);
nor U15394 (N_15394,N_10319,N_11902);
or U15395 (N_15395,N_8861,N_8228);
or U15396 (N_15396,N_10951,N_10765);
nand U15397 (N_15397,N_9474,N_9675);
and U15398 (N_15398,N_11284,N_11296);
nor U15399 (N_15399,N_10694,N_11553);
xor U15400 (N_15400,N_9007,N_11949);
xor U15401 (N_15401,N_9044,N_8482);
nand U15402 (N_15402,N_11455,N_11727);
nand U15403 (N_15403,N_11220,N_10554);
and U15404 (N_15404,N_8248,N_8519);
and U15405 (N_15405,N_9092,N_8178);
nor U15406 (N_15406,N_8776,N_10985);
or U15407 (N_15407,N_11186,N_8929);
or U15408 (N_15408,N_11387,N_8065);
or U15409 (N_15409,N_10691,N_10375);
and U15410 (N_15410,N_8576,N_9116);
nor U15411 (N_15411,N_11376,N_9946);
xnor U15412 (N_15412,N_11151,N_9103);
nor U15413 (N_15413,N_10029,N_10004);
nand U15414 (N_15414,N_10903,N_11815);
xnor U15415 (N_15415,N_11626,N_11366);
nand U15416 (N_15416,N_8818,N_11900);
nand U15417 (N_15417,N_11709,N_11738);
xor U15418 (N_15418,N_9574,N_8904);
nor U15419 (N_15419,N_10949,N_9129);
or U15420 (N_15420,N_10874,N_8390);
or U15421 (N_15421,N_11959,N_8154);
xor U15422 (N_15422,N_10095,N_10097);
nor U15423 (N_15423,N_11859,N_8211);
xnor U15424 (N_15424,N_10491,N_9853);
and U15425 (N_15425,N_9026,N_11026);
xor U15426 (N_15426,N_9109,N_10045);
or U15427 (N_15427,N_9575,N_10601);
or U15428 (N_15428,N_11410,N_11969);
and U15429 (N_15429,N_10078,N_10863);
nor U15430 (N_15430,N_11124,N_10634);
xnor U15431 (N_15431,N_11267,N_8692);
and U15432 (N_15432,N_8777,N_9736);
and U15433 (N_15433,N_8563,N_9278);
nand U15434 (N_15434,N_8311,N_9015);
nor U15435 (N_15435,N_10360,N_8509);
and U15436 (N_15436,N_11100,N_8468);
xnor U15437 (N_15437,N_10073,N_11751);
nor U15438 (N_15438,N_9863,N_9010);
nand U15439 (N_15439,N_11514,N_9465);
xor U15440 (N_15440,N_11051,N_9481);
nor U15441 (N_15441,N_8575,N_10995);
and U15442 (N_15442,N_11241,N_8717);
and U15443 (N_15443,N_11134,N_9866);
nand U15444 (N_15444,N_10713,N_9982);
nand U15445 (N_15445,N_8521,N_10332);
or U15446 (N_15446,N_9400,N_10486);
and U15447 (N_15447,N_10211,N_9997);
or U15448 (N_15448,N_11150,N_9602);
or U15449 (N_15449,N_10864,N_9490);
nor U15450 (N_15450,N_9557,N_9428);
xnor U15451 (N_15451,N_11627,N_8109);
or U15452 (N_15452,N_10518,N_8896);
and U15453 (N_15453,N_11631,N_8268);
xor U15454 (N_15454,N_8397,N_8192);
xor U15455 (N_15455,N_10688,N_10958);
xnor U15456 (N_15456,N_9164,N_11841);
nor U15457 (N_15457,N_11024,N_9826);
nand U15458 (N_15458,N_9554,N_9497);
nor U15459 (N_15459,N_11566,N_10381);
or U15460 (N_15460,N_11390,N_8588);
xnor U15461 (N_15461,N_11917,N_11196);
nand U15462 (N_15462,N_8593,N_8504);
nor U15463 (N_15463,N_9405,N_10778);
or U15464 (N_15464,N_9429,N_11023);
or U15465 (N_15465,N_11934,N_11679);
nor U15466 (N_15466,N_10038,N_10426);
xnor U15467 (N_15467,N_8291,N_10428);
nor U15468 (N_15468,N_11029,N_8937);
or U15469 (N_15469,N_9614,N_10418);
nand U15470 (N_15470,N_8750,N_11533);
or U15471 (N_15471,N_8007,N_8307);
nand U15472 (N_15472,N_10372,N_11339);
xnor U15473 (N_15473,N_10998,N_11715);
nor U15474 (N_15474,N_9050,N_8290);
nand U15475 (N_15475,N_11473,N_8082);
xor U15476 (N_15476,N_8467,N_11759);
or U15477 (N_15477,N_10644,N_8988);
or U15478 (N_15478,N_8233,N_9840);
nand U15479 (N_15479,N_9742,N_9424);
nand U15480 (N_15480,N_11428,N_11777);
nor U15481 (N_15481,N_8006,N_8555);
xor U15482 (N_15482,N_11121,N_9403);
and U15483 (N_15483,N_9503,N_10045);
and U15484 (N_15484,N_9505,N_9762);
nor U15485 (N_15485,N_9192,N_11022);
nor U15486 (N_15486,N_8910,N_8463);
nor U15487 (N_15487,N_11739,N_10092);
and U15488 (N_15488,N_10522,N_9418);
and U15489 (N_15489,N_11922,N_9649);
or U15490 (N_15490,N_10495,N_11150);
xnor U15491 (N_15491,N_11456,N_11887);
and U15492 (N_15492,N_10785,N_9493);
xnor U15493 (N_15493,N_11708,N_9408);
and U15494 (N_15494,N_10405,N_8811);
or U15495 (N_15495,N_11014,N_11316);
or U15496 (N_15496,N_11047,N_10073);
nand U15497 (N_15497,N_9033,N_8909);
xnor U15498 (N_15498,N_9082,N_11824);
and U15499 (N_15499,N_9871,N_10551);
nor U15500 (N_15500,N_8370,N_9076);
and U15501 (N_15501,N_10835,N_8145);
xor U15502 (N_15502,N_11827,N_11778);
xnor U15503 (N_15503,N_11918,N_11210);
xnor U15504 (N_15504,N_11094,N_8091);
nor U15505 (N_15505,N_10834,N_8572);
nor U15506 (N_15506,N_10110,N_10654);
nor U15507 (N_15507,N_11257,N_10108);
or U15508 (N_15508,N_8341,N_9611);
xnor U15509 (N_15509,N_11468,N_8543);
or U15510 (N_15510,N_9178,N_10484);
xor U15511 (N_15511,N_11467,N_11278);
xor U15512 (N_15512,N_11411,N_10841);
or U15513 (N_15513,N_9842,N_11369);
xnor U15514 (N_15514,N_8088,N_9943);
xnor U15515 (N_15515,N_10309,N_9327);
and U15516 (N_15516,N_9326,N_11235);
xnor U15517 (N_15517,N_8306,N_8656);
or U15518 (N_15518,N_9166,N_10812);
and U15519 (N_15519,N_10858,N_9290);
and U15520 (N_15520,N_9457,N_11344);
nor U15521 (N_15521,N_11360,N_10889);
or U15522 (N_15522,N_8496,N_8968);
and U15523 (N_15523,N_10085,N_11496);
or U15524 (N_15524,N_9446,N_11379);
nand U15525 (N_15525,N_10889,N_11721);
xnor U15526 (N_15526,N_11969,N_8673);
or U15527 (N_15527,N_9496,N_8703);
and U15528 (N_15528,N_11862,N_9319);
and U15529 (N_15529,N_11958,N_11885);
and U15530 (N_15530,N_8850,N_11649);
nor U15531 (N_15531,N_11938,N_9039);
nor U15532 (N_15532,N_8325,N_10649);
xor U15533 (N_15533,N_8570,N_8458);
xnor U15534 (N_15534,N_9432,N_9474);
and U15535 (N_15535,N_9891,N_10940);
xnor U15536 (N_15536,N_10904,N_10640);
or U15537 (N_15537,N_11853,N_8230);
nor U15538 (N_15538,N_9172,N_11316);
and U15539 (N_15539,N_11503,N_11328);
nand U15540 (N_15540,N_11682,N_9498);
and U15541 (N_15541,N_11468,N_11061);
or U15542 (N_15542,N_11419,N_10924);
nand U15543 (N_15543,N_11016,N_9321);
or U15544 (N_15544,N_8261,N_8950);
or U15545 (N_15545,N_10509,N_10920);
or U15546 (N_15546,N_8692,N_11914);
nand U15547 (N_15547,N_11257,N_9466);
nor U15548 (N_15548,N_10300,N_10445);
and U15549 (N_15549,N_8207,N_10645);
nor U15550 (N_15550,N_9695,N_11065);
nand U15551 (N_15551,N_9105,N_11239);
nor U15552 (N_15552,N_8541,N_10910);
or U15553 (N_15553,N_11034,N_10812);
nor U15554 (N_15554,N_9278,N_11226);
xnor U15555 (N_15555,N_11772,N_8968);
or U15556 (N_15556,N_10632,N_10411);
xor U15557 (N_15557,N_11211,N_9108);
xor U15558 (N_15558,N_11553,N_8846);
xnor U15559 (N_15559,N_9346,N_8926);
xor U15560 (N_15560,N_11074,N_11769);
or U15561 (N_15561,N_9055,N_10802);
nor U15562 (N_15562,N_9546,N_9929);
nand U15563 (N_15563,N_11009,N_8854);
and U15564 (N_15564,N_9834,N_8542);
xor U15565 (N_15565,N_11737,N_8890);
xor U15566 (N_15566,N_8421,N_9053);
nor U15567 (N_15567,N_11924,N_11411);
or U15568 (N_15568,N_9637,N_11750);
and U15569 (N_15569,N_11948,N_8459);
xor U15570 (N_15570,N_10381,N_10387);
and U15571 (N_15571,N_10122,N_11715);
and U15572 (N_15572,N_10110,N_11986);
xnor U15573 (N_15573,N_11000,N_11683);
nor U15574 (N_15574,N_10240,N_9920);
or U15575 (N_15575,N_9245,N_8755);
nor U15576 (N_15576,N_9731,N_8420);
and U15577 (N_15577,N_9483,N_11221);
and U15578 (N_15578,N_9963,N_9804);
nor U15579 (N_15579,N_8442,N_10320);
or U15580 (N_15580,N_11563,N_11329);
or U15581 (N_15581,N_11968,N_11183);
and U15582 (N_15582,N_8425,N_11566);
xor U15583 (N_15583,N_11473,N_9769);
xnor U15584 (N_15584,N_8995,N_11039);
or U15585 (N_15585,N_10983,N_10287);
or U15586 (N_15586,N_10144,N_9364);
or U15587 (N_15587,N_10557,N_9383);
and U15588 (N_15588,N_11591,N_11724);
nand U15589 (N_15589,N_11862,N_9279);
nand U15590 (N_15590,N_8541,N_8462);
or U15591 (N_15591,N_9253,N_9275);
nand U15592 (N_15592,N_11651,N_8153);
nand U15593 (N_15593,N_9265,N_11029);
xor U15594 (N_15594,N_8650,N_11201);
xnor U15595 (N_15595,N_11046,N_9119);
nor U15596 (N_15596,N_9656,N_9204);
xor U15597 (N_15597,N_8175,N_10009);
nor U15598 (N_15598,N_10614,N_10975);
or U15599 (N_15599,N_11263,N_8481);
and U15600 (N_15600,N_9433,N_10450);
or U15601 (N_15601,N_9920,N_11814);
and U15602 (N_15602,N_10245,N_9006);
xnor U15603 (N_15603,N_11404,N_8387);
nand U15604 (N_15604,N_8645,N_9959);
or U15605 (N_15605,N_11158,N_10490);
nor U15606 (N_15606,N_8174,N_11584);
nor U15607 (N_15607,N_8397,N_10143);
or U15608 (N_15608,N_9248,N_8856);
nand U15609 (N_15609,N_8904,N_9002);
xor U15610 (N_15610,N_8651,N_11518);
xor U15611 (N_15611,N_9053,N_11023);
and U15612 (N_15612,N_11094,N_10891);
and U15613 (N_15613,N_8646,N_8939);
nor U15614 (N_15614,N_10456,N_11688);
xor U15615 (N_15615,N_8962,N_8483);
xnor U15616 (N_15616,N_9453,N_11519);
xnor U15617 (N_15617,N_9673,N_9281);
or U15618 (N_15618,N_8747,N_8730);
nand U15619 (N_15619,N_10709,N_9449);
nand U15620 (N_15620,N_10733,N_9719);
and U15621 (N_15621,N_11225,N_8786);
nor U15622 (N_15622,N_10383,N_10952);
and U15623 (N_15623,N_11873,N_9293);
nor U15624 (N_15624,N_11433,N_10399);
or U15625 (N_15625,N_8134,N_10525);
nor U15626 (N_15626,N_10227,N_10868);
nor U15627 (N_15627,N_10412,N_8531);
nor U15628 (N_15628,N_10951,N_10513);
or U15629 (N_15629,N_8440,N_8578);
xnor U15630 (N_15630,N_9764,N_8019);
or U15631 (N_15631,N_10826,N_11207);
or U15632 (N_15632,N_8703,N_10556);
nor U15633 (N_15633,N_9464,N_8645);
or U15634 (N_15634,N_8632,N_8314);
nor U15635 (N_15635,N_11974,N_9101);
xnor U15636 (N_15636,N_9503,N_8755);
or U15637 (N_15637,N_11228,N_8666);
nor U15638 (N_15638,N_11679,N_9244);
nor U15639 (N_15639,N_9902,N_8700);
xnor U15640 (N_15640,N_11466,N_10946);
xor U15641 (N_15641,N_11464,N_10096);
nor U15642 (N_15642,N_11910,N_9008);
xnor U15643 (N_15643,N_10480,N_11073);
nor U15644 (N_15644,N_8265,N_8177);
and U15645 (N_15645,N_8932,N_11104);
or U15646 (N_15646,N_8171,N_9855);
and U15647 (N_15647,N_8290,N_8581);
or U15648 (N_15648,N_11272,N_8976);
nor U15649 (N_15649,N_8323,N_8726);
or U15650 (N_15650,N_10625,N_10319);
and U15651 (N_15651,N_9191,N_9896);
nor U15652 (N_15652,N_11881,N_8709);
xnor U15653 (N_15653,N_11770,N_11941);
and U15654 (N_15654,N_11684,N_8530);
nor U15655 (N_15655,N_10635,N_9914);
xnor U15656 (N_15656,N_11346,N_8052);
or U15657 (N_15657,N_11460,N_9938);
xnor U15658 (N_15658,N_11837,N_10309);
or U15659 (N_15659,N_11370,N_11602);
xnor U15660 (N_15660,N_8024,N_11964);
xnor U15661 (N_15661,N_9534,N_8047);
or U15662 (N_15662,N_10077,N_11070);
nor U15663 (N_15663,N_11303,N_9506);
nand U15664 (N_15664,N_8838,N_8024);
nor U15665 (N_15665,N_11264,N_10681);
nand U15666 (N_15666,N_8716,N_9041);
xnor U15667 (N_15667,N_11745,N_11852);
or U15668 (N_15668,N_10060,N_8397);
and U15669 (N_15669,N_11649,N_9517);
nand U15670 (N_15670,N_9360,N_8082);
or U15671 (N_15671,N_11249,N_11538);
xor U15672 (N_15672,N_11182,N_9390);
and U15673 (N_15673,N_10492,N_11239);
and U15674 (N_15674,N_11105,N_11515);
and U15675 (N_15675,N_8959,N_8244);
or U15676 (N_15676,N_11719,N_10159);
nor U15677 (N_15677,N_8100,N_8110);
nand U15678 (N_15678,N_10468,N_10777);
xnor U15679 (N_15679,N_8279,N_11215);
xnor U15680 (N_15680,N_8785,N_9813);
xor U15681 (N_15681,N_9460,N_9950);
or U15682 (N_15682,N_9475,N_10707);
xnor U15683 (N_15683,N_9054,N_8563);
nor U15684 (N_15684,N_8583,N_10598);
nand U15685 (N_15685,N_10954,N_9848);
nor U15686 (N_15686,N_10863,N_11683);
nand U15687 (N_15687,N_10866,N_11372);
and U15688 (N_15688,N_8039,N_9542);
xnor U15689 (N_15689,N_11764,N_10971);
or U15690 (N_15690,N_11870,N_9001);
nor U15691 (N_15691,N_8062,N_10112);
nor U15692 (N_15692,N_10749,N_11533);
nor U15693 (N_15693,N_9242,N_9831);
xnor U15694 (N_15694,N_11740,N_9334);
and U15695 (N_15695,N_11488,N_9311);
nand U15696 (N_15696,N_10424,N_11037);
nand U15697 (N_15697,N_11257,N_8419);
and U15698 (N_15698,N_8374,N_10478);
nor U15699 (N_15699,N_9281,N_9102);
and U15700 (N_15700,N_10182,N_11541);
xnor U15701 (N_15701,N_11000,N_11590);
or U15702 (N_15702,N_11608,N_9287);
or U15703 (N_15703,N_11622,N_11021);
xnor U15704 (N_15704,N_10194,N_8808);
and U15705 (N_15705,N_8389,N_10005);
and U15706 (N_15706,N_10215,N_11995);
nor U15707 (N_15707,N_11839,N_8406);
and U15708 (N_15708,N_9328,N_9096);
or U15709 (N_15709,N_10694,N_10194);
and U15710 (N_15710,N_9654,N_11457);
xnor U15711 (N_15711,N_11409,N_9717);
nor U15712 (N_15712,N_8543,N_9259);
and U15713 (N_15713,N_11489,N_10219);
xor U15714 (N_15714,N_11479,N_11139);
nor U15715 (N_15715,N_11984,N_11796);
xor U15716 (N_15716,N_9934,N_9112);
nand U15717 (N_15717,N_11992,N_11275);
and U15718 (N_15718,N_10886,N_11271);
nor U15719 (N_15719,N_9619,N_9083);
nor U15720 (N_15720,N_10392,N_11105);
nand U15721 (N_15721,N_11022,N_9582);
and U15722 (N_15722,N_9862,N_8441);
xnor U15723 (N_15723,N_9731,N_9979);
or U15724 (N_15724,N_8093,N_10879);
and U15725 (N_15725,N_11744,N_11322);
nand U15726 (N_15726,N_11243,N_11716);
or U15727 (N_15727,N_11034,N_11491);
nor U15728 (N_15728,N_8841,N_10406);
nand U15729 (N_15729,N_9552,N_8697);
nand U15730 (N_15730,N_10555,N_8738);
xor U15731 (N_15731,N_11327,N_11081);
or U15732 (N_15732,N_11376,N_11090);
or U15733 (N_15733,N_8333,N_11487);
and U15734 (N_15734,N_9278,N_8000);
and U15735 (N_15735,N_10941,N_9959);
or U15736 (N_15736,N_9003,N_10309);
and U15737 (N_15737,N_10315,N_8189);
nand U15738 (N_15738,N_11792,N_8031);
and U15739 (N_15739,N_9256,N_10267);
and U15740 (N_15740,N_11562,N_9647);
and U15741 (N_15741,N_9562,N_10003);
and U15742 (N_15742,N_9631,N_11281);
xor U15743 (N_15743,N_8606,N_9830);
and U15744 (N_15744,N_10452,N_11178);
and U15745 (N_15745,N_9782,N_8176);
and U15746 (N_15746,N_9354,N_10596);
xnor U15747 (N_15747,N_8185,N_9592);
xnor U15748 (N_15748,N_9598,N_8002);
xor U15749 (N_15749,N_10141,N_8250);
nor U15750 (N_15750,N_9890,N_11791);
nand U15751 (N_15751,N_9531,N_11715);
xnor U15752 (N_15752,N_10304,N_11992);
nand U15753 (N_15753,N_9313,N_11735);
nor U15754 (N_15754,N_10577,N_11140);
xnor U15755 (N_15755,N_8982,N_9128);
or U15756 (N_15756,N_8213,N_9362);
nor U15757 (N_15757,N_10705,N_11677);
or U15758 (N_15758,N_10490,N_10018);
xor U15759 (N_15759,N_11601,N_11964);
and U15760 (N_15760,N_9633,N_8286);
or U15761 (N_15761,N_10015,N_11049);
nor U15762 (N_15762,N_8319,N_9264);
nor U15763 (N_15763,N_11945,N_11815);
nand U15764 (N_15764,N_9856,N_11418);
or U15765 (N_15765,N_9424,N_10883);
and U15766 (N_15766,N_11460,N_8861);
and U15767 (N_15767,N_11423,N_9040);
xnor U15768 (N_15768,N_9728,N_8931);
or U15769 (N_15769,N_9923,N_10815);
xnor U15770 (N_15770,N_9396,N_11007);
or U15771 (N_15771,N_11630,N_8601);
or U15772 (N_15772,N_10899,N_11811);
nand U15773 (N_15773,N_11444,N_8742);
xnor U15774 (N_15774,N_9527,N_11777);
nor U15775 (N_15775,N_8034,N_9847);
nor U15776 (N_15776,N_9739,N_11108);
nor U15777 (N_15777,N_8753,N_8145);
or U15778 (N_15778,N_9025,N_8072);
nand U15779 (N_15779,N_9276,N_8262);
nand U15780 (N_15780,N_8486,N_8356);
nand U15781 (N_15781,N_8528,N_10589);
or U15782 (N_15782,N_11894,N_8883);
and U15783 (N_15783,N_11289,N_8227);
and U15784 (N_15784,N_10766,N_8404);
nand U15785 (N_15785,N_11347,N_9695);
nand U15786 (N_15786,N_9745,N_8486);
or U15787 (N_15787,N_11320,N_8463);
or U15788 (N_15788,N_11521,N_10143);
xor U15789 (N_15789,N_11722,N_10929);
nor U15790 (N_15790,N_10697,N_11451);
nor U15791 (N_15791,N_11465,N_10359);
xnor U15792 (N_15792,N_10127,N_10966);
nand U15793 (N_15793,N_11458,N_10733);
or U15794 (N_15794,N_9099,N_11654);
xnor U15795 (N_15795,N_9330,N_11386);
nand U15796 (N_15796,N_8361,N_11715);
or U15797 (N_15797,N_8774,N_10051);
or U15798 (N_15798,N_9098,N_10932);
nor U15799 (N_15799,N_9984,N_8806);
and U15800 (N_15800,N_8928,N_10732);
and U15801 (N_15801,N_9954,N_10380);
nor U15802 (N_15802,N_9457,N_9184);
nand U15803 (N_15803,N_9776,N_8319);
nor U15804 (N_15804,N_10830,N_11479);
nand U15805 (N_15805,N_11680,N_10760);
and U15806 (N_15806,N_9235,N_10920);
xor U15807 (N_15807,N_10943,N_11827);
nor U15808 (N_15808,N_11752,N_10742);
nor U15809 (N_15809,N_8206,N_8532);
nor U15810 (N_15810,N_11351,N_11859);
xnor U15811 (N_15811,N_11996,N_10046);
and U15812 (N_15812,N_10024,N_10122);
nor U15813 (N_15813,N_9342,N_9459);
nand U15814 (N_15814,N_8038,N_9955);
and U15815 (N_15815,N_11942,N_10560);
nor U15816 (N_15816,N_9405,N_10718);
xnor U15817 (N_15817,N_10483,N_8546);
or U15818 (N_15818,N_10128,N_9087);
or U15819 (N_15819,N_8980,N_11420);
nor U15820 (N_15820,N_8485,N_9636);
xor U15821 (N_15821,N_8045,N_11415);
nor U15822 (N_15822,N_9443,N_10719);
nand U15823 (N_15823,N_8553,N_10836);
or U15824 (N_15824,N_10385,N_10538);
nand U15825 (N_15825,N_8471,N_8037);
nor U15826 (N_15826,N_11964,N_8228);
or U15827 (N_15827,N_10497,N_11716);
nand U15828 (N_15828,N_9152,N_9825);
nand U15829 (N_15829,N_8358,N_8065);
nand U15830 (N_15830,N_11901,N_11022);
nand U15831 (N_15831,N_9210,N_10756);
or U15832 (N_15832,N_11504,N_10677);
or U15833 (N_15833,N_8440,N_11940);
and U15834 (N_15834,N_11728,N_10678);
and U15835 (N_15835,N_10489,N_11148);
or U15836 (N_15836,N_10209,N_10944);
nor U15837 (N_15837,N_10427,N_8496);
nor U15838 (N_15838,N_8828,N_10939);
xnor U15839 (N_15839,N_9099,N_9460);
xnor U15840 (N_15840,N_9482,N_10039);
and U15841 (N_15841,N_9981,N_9999);
nor U15842 (N_15842,N_11493,N_10024);
nor U15843 (N_15843,N_9978,N_8865);
nor U15844 (N_15844,N_11630,N_10872);
or U15845 (N_15845,N_9600,N_9787);
or U15846 (N_15846,N_10245,N_9692);
xor U15847 (N_15847,N_10949,N_10270);
xor U15848 (N_15848,N_11859,N_8330);
nor U15849 (N_15849,N_8643,N_9265);
nor U15850 (N_15850,N_8783,N_9477);
nor U15851 (N_15851,N_11178,N_11638);
or U15852 (N_15852,N_11345,N_8452);
nor U15853 (N_15853,N_10171,N_11218);
nand U15854 (N_15854,N_10659,N_9461);
nand U15855 (N_15855,N_8265,N_10032);
and U15856 (N_15856,N_9422,N_10950);
xnor U15857 (N_15857,N_9240,N_8215);
nand U15858 (N_15858,N_11853,N_10019);
or U15859 (N_15859,N_10490,N_9530);
nand U15860 (N_15860,N_11346,N_10873);
nor U15861 (N_15861,N_9089,N_9652);
xnor U15862 (N_15862,N_11008,N_8782);
xnor U15863 (N_15863,N_10157,N_11386);
nand U15864 (N_15864,N_8585,N_9333);
and U15865 (N_15865,N_10250,N_8895);
nand U15866 (N_15866,N_11819,N_10157);
nor U15867 (N_15867,N_8351,N_8541);
nor U15868 (N_15868,N_9871,N_9597);
or U15869 (N_15869,N_9252,N_9485);
or U15870 (N_15870,N_9163,N_10970);
and U15871 (N_15871,N_9222,N_9062);
or U15872 (N_15872,N_9299,N_10501);
nand U15873 (N_15873,N_10337,N_10490);
xor U15874 (N_15874,N_9654,N_11875);
or U15875 (N_15875,N_11717,N_11816);
or U15876 (N_15876,N_11668,N_8809);
or U15877 (N_15877,N_8784,N_11062);
nor U15878 (N_15878,N_11497,N_11249);
or U15879 (N_15879,N_11223,N_8578);
nor U15880 (N_15880,N_8488,N_11391);
or U15881 (N_15881,N_9300,N_10657);
and U15882 (N_15882,N_9946,N_9273);
and U15883 (N_15883,N_11267,N_11528);
nand U15884 (N_15884,N_9729,N_10984);
and U15885 (N_15885,N_8063,N_9039);
xor U15886 (N_15886,N_9854,N_9985);
or U15887 (N_15887,N_10100,N_10520);
nand U15888 (N_15888,N_11831,N_10061);
and U15889 (N_15889,N_11451,N_9993);
nand U15890 (N_15890,N_9019,N_9734);
and U15891 (N_15891,N_11212,N_10242);
and U15892 (N_15892,N_11313,N_8681);
or U15893 (N_15893,N_9302,N_10230);
and U15894 (N_15894,N_10966,N_8888);
or U15895 (N_15895,N_11865,N_11719);
or U15896 (N_15896,N_11393,N_8564);
nor U15897 (N_15897,N_8761,N_10903);
and U15898 (N_15898,N_11711,N_9331);
nand U15899 (N_15899,N_9133,N_9775);
or U15900 (N_15900,N_9685,N_9280);
or U15901 (N_15901,N_11794,N_9611);
xnor U15902 (N_15902,N_8351,N_10895);
and U15903 (N_15903,N_8096,N_11594);
nand U15904 (N_15904,N_10281,N_10414);
or U15905 (N_15905,N_10233,N_11848);
and U15906 (N_15906,N_10553,N_9501);
nor U15907 (N_15907,N_9754,N_11449);
nand U15908 (N_15908,N_11205,N_8588);
and U15909 (N_15909,N_8799,N_8314);
xnor U15910 (N_15910,N_8440,N_8871);
nor U15911 (N_15911,N_9780,N_8584);
or U15912 (N_15912,N_8459,N_10688);
or U15913 (N_15913,N_11522,N_11521);
nand U15914 (N_15914,N_11278,N_8339);
and U15915 (N_15915,N_10332,N_10702);
xnor U15916 (N_15916,N_8894,N_10379);
and U15917 (N_15917,N_8409,N_11612);
xor U15918 (N_15918,N_10462,N_8609);
nand U15919 (N_15919,N_10779,N_9654);
or U15920 (N_15920,N_8264,N_8352);
or U15921 (N_15921,N_11280,N_11816);
nand U15922 (N_15922,N_8623,N_9599);
nor U15923 (N_15923,N_9933,N_11389);
xor U15924 (N_15924,N_8010,N_9838);
nand U15925 (N_15925,N_9016,N_8922);
and U15926 (N_15926,N_9686,N_8337);
nand U15927 (N_15927,N_10122,N_10103);
nand U15928 (N_15928,N_11004,N_11734);
and U15929 (N_15929,N_10461,N_8684);
nor U15930 (N_15930,N_10404,N_10210);
or U15931 (N_15931,N_11679,N_8238);
xnor U15932 (N_15932,N_9023,N_10669);
and U15933 (N_15933,N_9384,N_11639);
nor U15934 (N_15934,N_11865,N_10209);
xnor U15935 (N_15935,N_8702,N_8038);
or U15936 (N_15936,N_11890,N_8887);
nand U15937 (N_15937,N_8044,N_10327);
nor U15938 (N_15938,N_11434,N_11461);
and U15939 (N_15939,N_8683,N_8162);
or U15940 (N_15940,N_9827,N_10955);
and U15941 (N_15941,N_11612,N_11568);
xor U15942 (N_15942,N_9185,N_10416);
or U15943 (N_15943,N_11440,N_11770);
xor U15944 (N_15944,N_9384,N_10433);
and U15945 (N_15945,N_10994,N_10654);
or U15946 (N_15946,N_11431,N_11761);
nor U15947 (N_15947,N_11849,N_9710);
nand U15948 (N_15948,N_8220,N_9376);
xnor U15949 (N_15949,N_10181,N_8973);
xnor U15950 (N_15950,N_8654,N_8587);
nor U15951 (N_15951,N_9947,N_10353);
and U15952 (N_15952,N_10392,N_10612);
or U15953 (N_15953,N_10100,N_9533);
nand U15954 (N_15954,N_8636,N_8466);
nand U15955 (N_15955,N_10340,N_10817);
nand U15956 (N_15956,N_10069,N_8447);
nor U15957 (N_15957,N_11512,N_11995);
nor U15958 (N_15958,N_10970,N_9946);
or U15959 (N_15959,N_8522,N_10215);
and U15960 (N_15960,N_8894,N_11938);
xnor U15961 (N_15961,N_10644,N_9901);
nor U15962 (N_15962,N_9190,N_8670);
xor U15963 (N_15963,N_8060,N_10277);
and U15964 (N_15964,N_10202,N_8997);
nand U15965 (N_15965,N_10776,N_11572);
nor U15966 (N_15966,N_8303,N_10833);
xnor U15967 (N_15967,N_10874,N_8233);
nand U15968 (N_15968,N_11744,N_8912);
or U15969 (N_15969,N_9873,N_9448);
or U15970 (N_15970,N_8243,N_8819);
and U15971 (N_15971,N_9250,N_8791);
or U15972 (N_15972,N_9110,N_11363);
and U15973 (N_15973,N_11327,N_11948);
xnor U15974 (N_15974,N_8556,N_11946);
xnor U15975 (N_15975,N_10674,N_8848);
nand U15976 (N_15976,N_10490,N_9720);
and U15977 (N_15977,N_8688,N_11782);
nand U15978 (N_15978,N_8437,N_9596);
or U15979 (N_15979,N_10451,N_9491);
nand U15980 (N_15980,N_11241,N_8695);
nand U15981 (N_15981,N_9613,N_10769);
xor U15982 (N_15982,N_10602,N_11925);
and U15983 (N_15983,N_8224,N_10247);
and U15984 (N_15984,N_9335,N_9737);
nand U15985 (N_15985,N_9399,N_9056);
nand U15986 (N_15986,N_10441,N_9818);
nor U15987 (N_15987,N_11134,N_8911);
nand U15988 (N_15988,N_11812,N_11511);
nor U15989 (N_15989,N_9956,N_11857);
and U15990 (N_15990,N_9064,N_9264);
and U15991 (N_15991,N_10286,N_8393);
or U15992 (N_15992,N_8072,N_8486);
nand U15993 (N_15993,N_8800,N_9797);
nand U15994 (N_15994,N_10307,N_11766);
nand U15995 (N_15995,N_8548,N_10562);
or U15996 (N_15996,N_9742,N_8326);
and U15997 (N_15997,N_9966,N_8565);
and U15998 (N_15998,N_8032,N_8918);
nand U15999 (N_15999,N_11420,N_10361);
nand U16000 (N_16000,N_13722,N_13977);
or U16001 (N_16001,N_12089,N_15104);
xor U16002 (N_16002,N_12173,N_15565);
nand U16003 (N_16003,N_15933,N_12404);
nor U16004 (N_16004,N_14835,N_13062);
xnor U16005 (N_16005,N_14265,N_13139);
xnor U16006 (N_16006,N_12748,N_14410);
xnor U16007 (N_16007,N_14550,N_14307);
or U16008 (N_16008,N_14313,N_13889);
or U16009 (N_16009,N_15017,N_12854);
nand U16010 (N_16010,N_13966,N_15515);
and U16011 (N_16011,N_13668,N_12062);
nor U16012 (N_16012,N_13171,N_13572);
or U16013 (N_16013,N_15680,N_12470);
or U16014 (N_16014,N_14813,N_13375);
and U16015 (N_16015,N_14637,N_12415);
nor U16016 (N_16016,N_13614,N_14672);
nand U16017 (N_16017,N_15187,N_15156);
nand U16018 (N_16018,N_14006,N_15728);
and U16019 (N_16019,N_13731,N_12247);
and U16020 (N_16020,N_13928,N_15297);
xor U16021 (N_16021,N_13828,N_14878);
nand U16022 (N_16022,N_12432,N_15098);
nand U16023 (N_16023,N_12873,N_14953);
and U16024 (N_16024,N_13983,N_14559);
and U16025 (N_16025,N_14444,N_14485);
or U16026 (N_16026,N_12780,N_14323);
or U16027 (N_16027,N_12257,N_15776);
nand U16028 (N_16028,N_13806,N_15366);
xnor U16029 (N_16029,N_14058,N_15558);
nor U16030 (N_16030,N_13713,N_13410);
nand U16031 (N_16031,N_13687,N_15294);
or U16032 (N_16032,N_14236,N_15781);
nand U16033 (N_16033,N_15486,N_14538);
nor U16034 (N_16034,N_15578,N_15115);
or U16035 (N_16035,N_15041,N_15418);
and U16036 (N_16036,N_12944,N_12770);
nand U16037 (N_16037,N_13647,N_12816);
and U16038 (N_16038,N_12505,N_14362);
nand U16039 (N_16039,N_13753,N_14502);
or U16040 (N_16040,N_12361,N_13798);
xnor U16041 (N_16041,N_12159,N_13717);
nor U16042 (N_16042,N_15474,N_14699);
xnor U16043 (N_16043,N_13699,N_12426);
or U16044 (N_16044,N_14063,N_12813);
or U16045 (N_16045,N_15787,N_13555);
nor U16046 (N_16046,N_15038,N_13154);
or U16047 (N_16047,N_15587,N_12135);
or U16048 (N_16048,N_13786,N_15477);
nand U16049 (N_16049,N_14914,N_14949);
and U16050 (N_16050,N_14226,N_12358);
or U16051 (N_16051,N_15892,N_14503);
xor U16052 (N_16052,N_13065,N_12961);
nand U16053 (N_16053,N_12075,N_12226);
or U16054 (N_16054,N_14624,N_15072);
nor U16055 (N_16055,N_15423,N_14783);
xor U16056 (N_16056,N_13190,N_12565);
and U16057 (N_16057,N_12355,N_15989);
and U16058 (N_16058,N_14967,N_12815);
xor U16059 (N_16059,N_12641,N_14640);
nand U16060 (N_16060,N_15481,N_12604);
xnor U16061 (N_16061,N_15709,N_15824);
and U16062 (N_16062,N_15410,N_14870);
nor U16063 (N_16063,N_13101,N_14175);
xor U16064 (N_16064,N_13744,N_14218);
xor U16065 (N_16065,N_12114,N_14602);
nand U16066 (N_16066,N_14816,N_13001);
nand U16067 (N_16067,N_14588,N_14147);
nand U16068 (N_16068,N_12281,N_15930);
nor U16069 (N_16069,N_15189,N_14189);
and U16070 (N_16070,N_12365,N_13089);
nor U16071 (N_16071,N_12157,N_12841);
nor U16072 (N_16072,N_12914,N_12674);
and U16073 (N_16073,N_14324,N_15659);
nor U16074 (N_16074,N_14556,N_12821);
and U16075 (N_16075,N_13645,N_14619);
xnor U16076 (N_16076,N_12186,N_15569);
xor U16077 (N_16077,N_12289,N_12125);
xnor U16078 (N_16078,N_14670,N_13719);
xor U16079 (N_16079,N_12002,N_12935);
and U16080 (N_16080,N_15870,N_14399);
nor U16081 (N_16081,N_14231,N_13801);
nand U16082 (N_16082,N_13814,N_12338);
nand U16083 (N_16083,N_13704,N_15111);
nor U16084 (N_16084,N_15853,N_13696);
or U16085 (N_16085,N_15346,N_15538);
or U16086 (N_16086,N_13505,N_15206);
or U16087 (N_16087,N_14178,N_14979);
and U16088 (N_16088,N_14002,N_13897);
or U16089 (N_16089,N_14441,N_14309);
and U16090 (N_16090,N_13308,N_12534);
nand U16091 (N_16091,N_14613,N_15947);
xnor U16092 (N_16092,N_14150,N_13223);
nand U16093 (N_16093,N_13618,N_13938);
nand U16094 (N_16094,N_12485,N_13063);
and U16095 (N_16095,N_15161,N_14088);
nand U16096 (N_16096,N_12948,N_12497);
xor U16097 (N_16097,N_13976,N_15946);
or U16098 (N_16098,N_13491,N_12253);
and U16099 (N_16099,N_12013,N_13274);
nand U16100 (N_16100,N_13091,N_14113);
or U16101 (N_16101,N_12993,N_12046);
xnor U16102 (N_16102,N_13960,N_14331);
and U16103 (N_16103,N_12086,N_14869);
xor U16104 (N_16104,N_14257,N_12718);
xor U16105 (N_16105,N_14689,N_15829);
and U16106 (N_16106,N_12801,N_13684);
nand U16107 (N_16107,N_13901,N_12288);
nand U16108 (N_16108,N_13849,N_12467);
xor U16109 (N_16109,N_13820,N_15421);
nand U16110 (N_16110,N_15692,N_12987);
nor U16111 (N_16111,N_13815,N_12922);
xnor U16112 (N_16112,N_12618,N_15390);
or U16113 (N_16113,N_12905,N_13194);
nand U16114 (N_16114,N_14859,N_12992);
xor U16115 (N_16115,N_13840,N_13005);
or U16116 (N_16116,N_14694,N_12874);
and U16117 (N_16117,N_15371,N_13400);
nor U16118 (N_16118,N_15269,N_13835);
xnor U16119 (N_16119,N_15729,N_12439);
nor U16120 (N_16120,N_15470,N_12304);
and U16121 (N_16121,N_13356,N_13393);
nor U16122 (N_16122,N_15218,N_14888);
and U16123 (N_16123,N_14751,N_13298);
or U16124 (N_16124,N_15253,N_14668);
and U16125 (N_16125,N_12410,N_12640);
and U16126 (N_16126,N_12824,N_13403);
nand U16127 (N_16127,N_13041,N_13539);
xor U16128 (N_16128,N_13353,N_15311);
nor U16129 (N_16129,N_15670,N_14123);
nand U16130 (N_16130,N_15971,N_13252);
nor U16131 (N_16131,N_14375,N_13218);
or U16132 (N_16132,N_15281,N_14807);
nor U16133 (N_16133,N_15209,N_15237);
and U16134 (N_16134,N_15388,N_15172);
nand U16135 (N_16135,N_13965,N_15018);
nor U16136 (N_16136,N_12723,N_13258);
or U16137 (N_16137,N_12872,N_12324);
nand U16138 (N_16138,N_15998,N_15931);
nor U16139 (N_16139,N_15717,N_14373);
xnor U16140 (N_16140,N_15555,N_15282);
and U16141 (N_16141,N_14931,N_12004);
or U16142 (N_16142,N_13823,N_14061);
nand U16143 (N_16143,N_13790,N_13852);
or U16144 (N_16144,N_15148,N_14729);
and U16145 (N_16145,N_13012,N_13510);
and U16146 (N_16146,N_12556,N_15243);
nor U16147 (N_16147,N_14112,N_12176);
nand U16148 (N_16148,N_14015,N_14267);
xnor U16149 (N_16149,N_13461,N_12825);
nor U16150 (N_16150,N_12745,N_13692);
or U16151 (N_16151,N_15912,N_13818);
nand U16152 (N_16152,N_14459,N_15900);
xor U16153 (N_16153,N_12834,N_13201);
or U16154 (N_16154,N_13975,N_14627);
or U16155 (N_16155,N_15216,N_15133);
nand U16156 (N_16156,N_12945,N_13037);
or U16157 (N_16157,N_15446,N_15234);
and U16158 (N_16158,N_13902,N_14301);
or U16159 (N_16159,N_12340,N_12325);
or U16160 (N_16160,N_13459,N_14527);
or U16161 (N_16161,N_15554,N_15638);
or U16162 (N_16162,N_14449,N_12830);
xnor U16163 (N_16163,N_14174,N_14306);
or U16164 (N_16164,N_12005,N_13147);
or U16165 (N_16165,N_14037,N_15437);
xor U16166 (N_16166,N_13387,N_13413);
xor U16167 (N_16167,N_12291,N_15197);
nand U16168 (N_16168,N_12330,N_13899);
xor U16169 (N_16169,N_15419,N_12855);
or U16170 (N_16170,N_14083,N_14270);
xor U16171 (N_16171,N_12721,N_14899);
xnor U16172 (N_16172,N_13197,N_13864);
nand U16173 (N_16173,N_14078,N_13069);
or U16174 (N_16174,N_15695,N_13374);
or U16175 (N_16175,N_15322,N_14520);
nor U16176 (N_16176,N_12318,N_14902);
xor U16177 (N_16177,N_12024,N_13034);
xor U16178 (N_16178,N_13986,N_12570);
and U16179 (N_16179,N_12464,N_14514);
and U16180 (N_16180,N_12143,N_14705);
or U16181 (N_16181,N_13270,N_14885);
nand U16182 (N_16182,N_15827,N_13691);
or U16183 (N_16183,N_15043,N_12206);
or U16184 (N_16184,N_12493,N_14992);
xor U16185 (N_16185,N_13825,N_13882);
xor U16186 (N_16186,N_14724,N_14182);
nand U16187 (N_16187,N_15948,N_15888);
or U16188 (N_16188,N_13924,N_14909);
and U16189 (N_16189,N_15006,N_15014);
nand U16190 (N_16190,N_14793,N_12270);
nor U16191 (N_16191,N_12309,N_12717);
nor U16192 (N_16192,N_12805,N_13169);
nand U16193 (N_16193,N_14042,N_12583);
xnor U16194 (N_16194,N_13752,N_14455);
and U16195 (N_16195,N_13475,N_13567);
nand U16196 (N_16196,N_14688,N_13916);
nand U16197 (N_16197,N_13575,N_12042);
and U16198 (N_16198,N_13412,N_15887);
nor U16199 (N_16199,N_15633,N_15483);
nor U16200 (N_16200,N_14062,N_15743);
nor U16201 (N_16201,N_13606,N_15720);
nand U16202 (N_16202,N_14418,N_13526);
and U16203 (N_16203,N_15192,N_12906);
nand U16204 (N_16204,N_14880,N_12000);
or U16205 (N_16205,N_15866,N_15763);
nor U16206 (N_16206,N_12388,N_13275);
xor U16207 (N_16207,N_13826,N_14763);
nand U16208 (N_16208,N_15059,N_14828);
nor U16209 (N_16209,N_13803,N_14738);
nand U16210 (N_16210,N_15022,N_13980);
or U16211 (N_16211,N_14017,N_13942);
or U16212 (N_16212,N_15716,N_14634);
nor U16213 (N_16213,N_14050,N_13866);
xor U16214 (N_16214,N_14641,N_15961);
nand U16215 (N_16215,N_12681,N_13911);
nand U16216 (N_16216,N_14394,N_15178);
nand U16217 (N_16217,N_15040,N_12424);
nor U16218 (N_16218,N_13469,N_12725);
xnor U16219 (N_16219,N_15158,N_12158);
xnor U16220 (N_16220,N_13020,N_12455);
nand U16221 (N_16221,N_15517,N_12146);
and U16222 (N_16222,N_15272,N_15445);
nand U16223 (N_16223,N_13504,N_15754);
xnor U16224 (N_16224,N_12017,N_14762);
or U16225 (N_16225,N_13226,N_15263);
or U16226 (N_16226,N_13281,N_12085);
and U16227 (N_16227,N_12728,N_15087);
and U16228 (N_16228,N_14294,N_12312);
nand U16229 (N_16229,N_14060,N_15348);
xor U16230 (N_16230,N_13221,N_14489);
xnor U16231 (N_16231,N_13925,N_15976);
xnor U16232 (N_16232,N_12191,N_12994);
or U16233 (N_16233,N_14168,N_14528);
or U16234 (N_16234,N_14551,N_15983);
and U16235 (N_16235,N_15738,N_14047);
and U16236 (N_16236,N_14412,N_12831);
and U16237 (N_16237,N_12018,N_13132);
nand U16238 (N_16238,N_14454,N_14179);
nand U16239 (N_16239,N_14377,N_15898);
xnor U16240 (N_16240,N_13573,N_14658);
nand U16241 (N_16241,N_14841,N_13228);
xor U16242 (N_16242,N_14187,N_15560);
xor U16243 (N_16243,N_12925,N_15822);
nand U16244 (N_16244,N_13155,N_12224);
or U16245 (N_16245,N_15368,N_15732);
nand U16246 (N_16246,N_14234,N_15862);
xor U16247 (N_16247,N_13427,N_15747);
xnor U16248 (N_16248,N_12677,N_12675);
nor U16249 (N_16249,N_13779,N_15540);
and U16250 (N_16250,N_12055,N_14848);
nand U16251 (N_16251,N_15271,N_15190);
and U16252 (N_16252,N_15583,N_14847);
nor U16253 (N_16253,N_13198,N_15984);
and U16254 (N_16254,N_15122,N_13689);
and U16255 (N_16255,N_14838,N_13780);
nor U16256 (N_16256,N_15774,N_15492);
and U16257 (N_16257,N_12329,N_14843);
xor U16258 (N_16258,N_15413,N_15839);
nand U16259 (N_16259,N_15154,N_15547);
nand U16260 (N_16260,N_13813,N_13896);
and U16261 (N_16261,N_14702,N_15378);
nand U16262 (N_16262,N_14803,N_14214);
nor U16263 (N_16263,N_14811,N_14387);
or U16264 (N_16264,N_14928,N_14923);
nor U16265 (N_16265,N_15110,N_14163);
nand U16266 (N_16266,N_14760,N_12278);
xnor U16267 (N_16267,N_15544,N_13754);
xnor U16268 (N_16268,N_14129,N_12096);
or U16269 (N_16269,N_14114,N_15536);
and U16270 (N_16270,N_13470,N_13343);
nand U16271 (N_16271,N_13391,N_15061);
nor U16272 (N_16272,N_14476,N_13935);
xor U16273 (N_16273,N_12368,N_14831);
and U16274 (N_16274,N_14916,N_13143);
and U16275 (N_16275,N_13199,N_15454);
or U16276 (N_16276,N_15557,N_15857);
and U16277 (N_16277,N_12975,N_13629);
and U16278 (N_16278,N_15200,N_15542);
and U16279 (N_16279,N_14453,N_12030);
nand U16280 (N_16280,N_12754,N_13168);
nor U16281 (N_16281,N_12421,N_14016);
nand U16282 (N_16282,N_14706,N_13277);
nand U16283 (N_16283,N_14797,N_12938);
xnor U16284 (N_16284,N_12222,N_15600);
and U16285 (N_16285,N_13662,N_15220);
or U16286 (N_16286,N_14571,N_14090);
nand U16287 (N_16287,N_13777,N_12742);
nor U16288 (N_16288,N_14995,N_12131);
nor U16289 (N_16289,N_14385,N_15904);
nand U16290 (N_16290,N_14573,N_13732);
nor U16291 (N_16291,N_12242,N_12259);
xor U16292 (N_16292,N_12538,N_15958);
or U16293 (N_16293,N_14287,N_13487);
nor U16294 (N_16294,N_14126,N_12755);
nor U16295 (N_16295,N_12212,N_14462);
xor U16296 (N_16296,N_14443,N_14926);
or U16297 (N_16297,N_14583,N_13898);
xor U16298 (N_16298,N_15581,N_15602);
nor U16299 (N_16299,N_14767,N_15498);
and U16300 (N_16300,N_12384,N_12239);
nor U16301 (N_16301,N_13317,N_12926);
xnor U16302 (N_16302,N_12620,N_14593);
xnor U16303 (N_16303,N_14884,N_14330);
nand U16304 (N_16304,N_13110,N_15973);
or U16305 (N_16305,N_13832,N_13339);
and U16306 (N_16306,N_15279,N_14834);
xnor U16307 (N_16307,N_13758,N_12704);
xnor U16308 (N_16308,N_15066,N_15796);
nor U16309 (N_16309,N_15939,N_14321);
and U16310 (N_16310,N_15146,N_13432);
and U16311 (N_16311,N_15360,N_13426);
and U16312 (N_16312,N_13316,N_12666);
and U16313 (N_16313,N_14827,N_14285);
nand U16314 (N_16314,N_13589,N_14703);
and U16315 (N_16315,N_15980,N_14024);
or U16316 (N_16316,N_12659,N_15881);
or U16317 (N_16317,N_14603,N_12646);
xor U16318 (N_16318,N_14028,N_14326);
xor U16319 (N_16319,N_14308,N_12525);
and U16320 (N_16320,N_13466,N_12516);
or U16321 (N_16321,N_12328,N_14907);
and U16322 (N_16322,N_14130,N_12475);
or U16323 (N_16323,N_15011,N_14320);
and U16324 (N_16324,N_15710,N_15049);
nand U16325 (N_16325,N_12777,N_12586);
xor U16326 (N_16326,N_13827,N_13913);
xor U16327 (N_16327,N_13090,N_12979);
and U16328 (N_16328,N_13536,N_12150);
xor U16329 (N_16329,N_15491,N_15117);
nor U16330 (N_16330,N_15664,N_14570);
nor U16331 (N_16331,N_15576,N_13048);
and U16332 (N_16332,N_12882,N_15609);
nor U16333 (N_16333,N_12753,N_14769);
xor U16334 (N_16334,N_15396,N_12121);
nand U16335 (N_16335,N_12082,N_13013);
nor U16336 (N_16336,N_12968,N_14939);
nor U16337 (N_16337,N_15497,N_15264);
nor U16338 (N_16338,N_13763,N_13061);
xor U16339 (N_16339,N_15114,N_13544);
or U16340 (N_16340,N_15401,N_13373);
nor U16341 (N_16341,N_13655,N_14104);
nand U16342 (N_16342,N_13646,N_13157);
and U16343 (N_16343,N_14714,N_13733);
or U16344 (N_16344,N_12683,N_13566);
and U16345 (N_16345,N_15969,N_15365);
and U16346 (N_16346,N_14127,N_15439);
or U16347 (N_16347,N_15674,N_14333);
nand U16348 (N_16348,N_12901,N_15610);
or U16349 (N_16349,N_13150,N_13789);
and U16350 (N_16350,N_14122,N_15287);
nand U16351 (N_16351,N_13893,N_12795);
nor U16352 (N_16352,N_15259,N_13671);
and U16353 (N_16353,N_14351,N_15619);
nor U16354 (N_16354,N_14825,N_12936);
or U16355 (N_16355,N_13452,N_13399);
or U16356 (N_16356,N_14782,N_13576);
nand U16357 (N_16357,N_15001,N_13659);
and U16358 (N_16358,N_13049,N_12868);
or U16359 (N_16359,N_13830,N_12829);
or U16360 (N_16360,N_12773,N_15416);
nor U16361 (N_16361,N_14504,N_14988);
or U16362 (N_16362,N_14701,N_15735);
and U16363 (N_16363,N_13879,N_14601);
xor U16364 (N_16364,N_12489,N_15586);
nor U16365 (N_16365,N_13970,N_14575);
nor U16366 (N_16366,N_15910,N_13776);
nor U16367 (N_16367,N_15250,N_12769);
nor U16368 (N_16368,N_12553,N_13599);
or U16369 (N_16369,N_13102,N_14700);
or U16370 (N_16370,N_12835,N_13590);
or U16371 (N_16371,N_14761,N_13021);
and U16372 (N_16372,N_12495,N_14229);
xnor U16373 (N_16373,N_13657,N_13366);
or U16374 (N_16374,N_13266,N_15278);
nand U16375 (N_16375,N_12481,N_12602);
or U16376 (N_16376,N_14947,N_12653);
nor U16377 (N_16377,N_14020,N_15548);
and U16378 (N_16378,N_15162,N_12302);
and U16379 (N_16379,N_15952,N_13064);
nor U16380 (N_16380,N_14161,N_13774);
xor U16381 (N_16381,N_15962,N_13623);
or U16382 (N_16382,N_12663,N_15286);
nand U16383 (N_16383,N_15302,N_12272);
xor U16384 (N_16384,N_13947,N_13520);
nor U16385 (N_16385,N_14106,N_13395);
nand U16386 (N_16386,N_13148,N_14148);
xor U16387 (N_16387,N_12217,N_13341);
xor U16388 (N_16388,N_13163,N_13907);
and U16389 (N_16389,N_13128,N_14642);
or U16390 (N_16390,N_13519,N_14228);
or U16391 (N_16391,N_13680,N_12227);
and U16392 (N_16392,N_15511,N_13251);
xnor U16393 (N_16393,N_12892,N_12316);
and U16394 (N_16394,N_15164,N_14105);
nor U16395 (N_16395,N_15831,N_13730);
nand U16396 (N_16396,N_13292,N_14167);
nor U16397 (N_16397,N_12946,N_13909);
nor U16398 (N_16398,N_13097,N_13802);
nor U16399 (N_16399,N_14348,N_12295);
xnor U16400 (N_16400,N_14479,N_15714);
or U16401 (N_16401,N_13369,N_15628);
nand U16402 (N_16402,N_12271,N_15367);
and U16403 (N_16403,N_13253,N_14289);
xor U16404 (N_16404,N_14993,N_15568);
xor U16405 (N_16405,N_13950,N_13952);
nor U16406 (N_16406,N_15846,N_13113);
nand U16407 (N_16407,N_14419,N_12419);
nor U16408 (N_16408,N_15997,N_15848);
or U16409 (N_16409,N_13446,N_14456);
nand U16410 (N_16410,N_14990,N_12320);
and U16411 (N_16411,N_12094,N_12740);
and U16412 (N_16412,N_12635,N_14201);
and U16413 (N_16413,N_14662,N_12194);
nor U16414 (N_16414,N_14291,N_14927);
nor U16415 (N_16415,N_14341,N_13043);
and U16416 (N_16416,N_15813,N_15566);
nand U16417 (N_16417,N_13628,N_13074);
xor U16418 (N_16418,N_14789,N_14604);
xor U16419 (N_16419,N_14303,N_15918);
and U16420 (N_16420,N_14958,N_13917);
nor U16421 (N_16421,N_14260,N_13514);
and U16422 (N_16422,N_13014,N_12652);
nor U16423 (N_16423,N_12457,N_14810);
nand U16424 (N_16424,N_12246,N_12285);
nand U16425 (N_16425,N_13953,N_12904);
xor U16426 (N_16426,N_13152,N_12354);
or U16427 (N_16427,N_12921,N_15270);
xnor U16428 (N_16428,N_14530,N_14448);
xor U16429 (N_16429,N_13636,N_13002);
xor U16430 (N_16430,N_13245,N_15883);
xnor U16431 (N_16431,N_12336,N_15230);
nor U16432 (N_16432,N_14007,N_12654);
xor U16433 (N_16433,N_13357,N_13365);
and U16434 (N_16434,N_14707,N_13437);
xor U16435 (N_16435,N_12240,N_12452);
nand U16436 (N_16436,N_15579,N_13364);
and U16437 (N_16437,N_12308,N_13793);
xnor U16438 (N_16438,N_12373,N_15181);
or U16439 (N_16439,N_13821,N_14430);
nor U16440 (N_16440,N_12839,N_15207);
nor U16441 (N_16441,N_14259,N_15266);
xnor U16442 (N_16442,N_12183,N_14429);
xor U16443 (N_16443,N_15885,N_14258);
and U16444 (N_16444,N_13115,N_14092);
nor U16445 (N_16445,N_15212,N_12164);
or U16446 (N_16446,N_13170,N_14533);
nor U16447 (N_16447,N_15490,N_12450);
or U16448 (N_16448,N_14679,N_13421);
and U16449 (N_16449,N_12015,N_14969);
and U16450 (N_16450,N_15325,N_12326);
nor U16451 (N_16451,N_14157,N_15328);
nand U16452 (N_16452,N_12615,N_13869);
nand U16453 (N_16453,N_13552,N_12265);
nor U16454 (N_16454,N_14737,N_12864);
and U16455 (N_16455,N_12040,N_12099);
nand U16456 (N_16456,N_14293,N_12767);
nand U16457 (N_16457,N_13808,N_13883);
nand U16458 (N_16458,N_14589,N_14021);
nor U16459 (N_16459,N_12095,N_13664);
or U16460 (N_16460,N_14073,N_13868);
or U16461 (N_16461,N_12123,N_14023);
xnor U16462 (N_16462,N_13473,N_15167);
nor U16463 (N_16463,N_12954,N_13286);
and U16464 (N_16464,N_15152,N_13665);
nand U16465 (N_16465,N_12260,N_15753);
nand U16466 (N_16466,N_14963,N_15450);
nor U16467 (N_16467,N_12597,N_13990);
nand U16468 (N_16468,N_14482,N_12417);
nand U16469 (N_16469,N_15426,N_14532);
or U16470 (N_16470,N_13746,N_13345);
nor U16471 (N_16471,N_12581,N_12851);
and U16472 (N_16472,N_14547,N_12201);
nor U16473 (N_16473,N_12701,N_14590);
and U16474 (N_16474,N_13107,N_14173);
nor U16475 (N_16475,N_15730,N_12978);
xnor U16476 (N_16476,N_12826,N_13500);
and U16477 (N_16477,N_14403,N_12580);
nor U16478 (N_16478,N_13997,N_14082);
or U16479 (N_16479,N_15217,N_13431);
or U16480 (N_16480,N_12964,N_14868);
nand U16481 (N_16481,N_13705,N_12636);
or U16482 (N_16482,N_14413,N_14146);
or U16483 (N_16483,N_15075,N_13362);
or U16484 (N_16484,N_14209,N_12530);
or U16485 (N_16485,N_15356,N_12208);
and U16486 (N_16486,N_14339,N_15685);
xor U16487 (N_16487,N_14276,N_13122);
or U16488 (N_16488,N_15223,N_14788);
nand U16489 (N_16489,N_13819,N_14808);
xor U16490 (N_16490,N_12512,N_13562);
or U16491 (N_16491,N_15400,N_14465);
xor U16492 (N_16492,N_13234,N_14975);
or U16493 (N_16493,N_15712,N_13710);
nor U16494 (N_16494,N_14615,N_13644);
or U16495 (N_16495,N_13648,N_12408);
and U16496 (N_16496,N_15475,N_15341);
xnor U16497 (N_16497,N_15484,N_15045);
nand U16498 (N_16498,N_15639,N_13238);
or U16499 (N_16499,N_15847,N_12269);
xnor U16500 (N_16500,N_14460,N_14855);
nor U16501 (N_16501,N_15002,N_15711);
or U16502 (N_16502,N_13133,N_15165);
xnor U16503 (N_16503,N_15826,N_15097);
nor U16504 (N_16504,N_13036,N_15570);
or U16505 (N_16505,N_15183,N_13285);
nand U16506 (N_16506,N_14446,N_13837);
or U16507 (N_16507,N_15150,N_14644);
nand U16508 (N_16508,N_15280,N_14665);
nand U16509 (N_16509,N_13654,N_12198);
xnor U16510 (N_16510,N_13712,N_12154);
nand U16511 (N_16511,N_13631,N_14065);
nand U16512 (N_16512,N_15026,N_12381);
nand U16513 (N_16513,N_15238,N_14681);
nand U16514 (N_16514,N_13322,N_12076);
or U16515 (N_16515,N_15257,N_14610);
or U16516 (N_16516,N_13165,N_14636);
xor U16517 (N_16517,N_14137,N_14824);
xor U16518 (N_16518,N_13540,N_12889);
nand U16519 (N_16519,N_15415,N_14045);
and U16520 (N_16520,N_15179,N_13734);
and U16521 (N_16521,N_15782,N_12884);
xnor U16522 (N_16522,N_15031,N_14980);
nor U16523 (N_16523,N_15244,N_13182);
and U16524 (N_16524,N_14991,N_15873);
xnor U16525 (N_16525,N_14690,N_14781);
nor U16526 (N_16526,N_15195,N_14158);
xor U16527 (N_16527,N_14138,N_13738);
nand U16528 (N_16528,N_12682,N_12548);
or U16529 (N_16529,N_15319,N_15911);
or U16530 (N_16530,N_15101,N_14057);
or U16531 (N_16531,N_14924,N_14791);
and U16532 (N_16532,N_13846,N_14244);
xnor U16533 (N_16533,N_12713,N_13246);
or U16534 (N_16534,N_14973,N_12802);
and U16535 (N_16535,N_14865,N_15021);
xnor U16536 (N_16536,N_15742,N_12193);
nor U16537 (N_16537,N_15029,N_14632);
or U16538 (N_16538,N_13386,N_14829);
nor U16539 (N_16539,N_14833,N_12877);
xnor U16540 (N_16540,N_13914,N_12932);
nor U16541 (N_16541,N_14384,N_12971);
or U16542 (N_16542,N_14852,N_12364);
xor U16543 (N_16543,N_14160,N_15327);
and U16544 (N_16544,N_13382,N_12933);
nor U16545 (N_16545,N_15788,N_14565);
xnor U16546 (N_16546,N_13844,N_14343);
nor U16547 (N_16547,N_15621,N_13425);
and U16548 (N_16548,N_14312,N_14049);
and U16549 (N_16549,N_12607,N_14625);
nor U16550 (N_16550,N_15525,N_14211);
nand U16551 (N_16551,N_14858,N_14431);
nor U16552 (N_16552,N_13872,N_12870);
or U16553 (N_16553,N_12705,N_13532);
xnor U16554 (N_16554,N_12366,N_15830);
and U16555 (N_16555,N_12827,N_14611);
nor U16556 (N_16556,N_15724,N_13745);
nor U16557 (N_16557,N_13688,N_14223);
or U16558 (N_16558,N_14202,N_12229);
nor U16559 (N_16559,N_14739,N_12594);
xor U16560 (N_16560,N_14962,N_14569);
nor U16561 (N_16561,N_12540,N_15298);
or U16562 (N_16562,N_14420,N_12385);
nand U16563 (N_16563,N_14068,N_12202);
or U16564 (N_16564,N_15869,N_12650);
xnor U16565 (N_16565,N_12751,N_14031);
nor U16566 (N_16566,N_14523,N_15599);
or U16567 (N_16567,N_12351,N_15531);
nand U16568 (N_16568,N_14464,N_13210);
xor U16569 (N_16569,N_12077,N_15513);
and U16570 (N_16570,N_15016,N_13711);
nand U16571 (N_16571,N_15694,N_15033);
xnor U16572 (N_16572,N_13513,N_12523);
nor U16573 (N_16573,N_15089,N_14432);
nand U16574 (N_16574,N_13998,N_12036);
and U16575 (N_16575,N_12019,N_13324);
nand U16576 (N_16576,N_13811,N_13954);
or U16577 (N_16577,N_15688,N_12859);
and U16578 (N_16578,N_13658,N_12842);
and U16579 (N_16579,N_12731,N_15137);
and U16580 (N_16580,N_15701,N_15314);
nand U16581 (N_16581,N_14345,N_12915);
and U16582 (N_16582,N_14108,N_12087);
nand U16583 (N_16583,N_12596,N_12029);
nor U16584 (N_16584,N_12502,N_14595);
and U16585 (N_16585,N_12508,N_12063);
xor U16586 (N_16586,N_13415,N_15719);
or U16587 (N_16587,N_14156,N_14996);
and U16588 (N_16588,N_15915,N_12274);
nor U16589 (N_16589,N_13568,N_13242);
and U16590 (N_16590,N_12976,N_14125);
and U16591 (N_16591,N_14193,N_15047);
nand U16592 (N_16592,N_13807,N_12339);
and U16593 (N_16593,N_15646,N_15140);
nor U16594 (N_16594,N_13912,N_15096);
nand U16595 (N_16595,N_14409,N_14795);
xor U16596 (N_16596,N_14398,N_14118);
nand U16597 (N_16597,N_15361,N_13756);
or U16598 (N_16598,N_15503,N_15036);
or U16599 (N_16599,N_14004,N_15950);
nand U16600 (N_16600,N_13149,N_15383);
or U16601 (N_16601,N_14579,N_15636);
or U16602 (N_16602,N_12589,N_14250);
xnor U16603 (N_16603,N_14856,N_13805);
and U16604 (N_16604,N_12990,N_15955);
nand U16605 (N_16605,N_13202,N_15926);
nor U16606 (N_16606,N_13138,N_14806);
and U16607 (N_16607,N_14621,N_15987);
nor U16608 (N_16608,N_15797,N_14526);
nor U16609 (N_16609,N_13506,N_14915);
and U16610 (N_16610,N_15650,N_13622);
xnor U16611 (N_16611,N_12606,N_14363);
nor U16612 (N_16612,N_13280,N_14305);
xor U16613 (N_16613,N_15329,N_12436);
and U16614 (N_16614,N_14540,N_14633);
and U16615 (N_16615,N_15937,N_12392);
or U16616 (N_16616,N_13946,N_14535);
nor U16617 (N_16617,N_13894,N_13905);
xnor U16618 (N_16618,N_15995,N_13574);
nor U16619 (N_16619,N_15236,N_12106);
xnor U16620 (N_16620,N_13456,N_14117);
xor U16621 (N_16621,N_12139,N_15681);
nand U16622 (N_16622,N_14358,N_12937);
xor U16623 (N_16623,N_13055,N_14686);
or U16624 (N_16624,N_14863,N_13485);
nor U16625 (N_16625,N_13249,N_15116);
xor U16626 (N_16626,N_13371,N_13130);
nand U16627 (N_16627,N_14605,N_14994);
and U16628 (N_16628,N_14458,N_13187);
xnor U16629 (N_16629,N_15151,N_14251);
or U16630 (N_16630,N_15373,N_12856);
xnor U16631 (N_16631,N_15810,N_13455);
nand U16632 (N_16632,N_12599,N_15734);
and U16633 (N_16633,N_15449,N_14587);
nand U16634 (N_16634,N_13527,N_13367);
and U16635 (N_16635,N_14009,N_13127);
nor U16636 (N_16636,N_15828,N_15843);
and U16637 (N_16637,N_13423,N_12129);
xnor U16638 (N_16638,N_13698,N_14792);
xnor U16639 (N_16639,N_15127,N_13772);
nor U16640 (N_16640,N_14720,N_13177);
xor U16641 (N_16641,N_14381,N_14038);
nand U16642 (N_16642,N_13380,N_13507);
and U16643 (N_16643,N_14096,N_13478);
and U16644 (N_16644,N_14521,N_15109);
or U16645 (N_16645,N_13987,N_12225);
xor U16646 (N_16646,N_12422,N_13344);
nor U16647 (N_16647,N_12785,N_15509);
and U16648 (N_16648,N_14043,N_15996);
xor U16649 (N_16649,N_14591,N_14233);
or U16650 (N_16650,N_12353,N_12402);
xnor U16651 (N_16651,N_12631,N_14372);
nand U16652 (N_16652,N_12223,N_12182);
xor U16653 (N_16653,N_12022,N_14280);
and U16654 (N_16654,N_12065,N_12794);
xnor U16655 (N_16655,N_13451,N_15905);
nor U16656 (N_16656,N_14785,N_12112);
or U16657 (N_16657,N_15461,N_12584);
and U16658 (N_16658,N_14401,N_15740);
nand U16659 (N_16659,N_13847,N_15232);
or U16660 (N_16660,N_12671,N_13797);
xnor U16661 (N_16661,N_14467,N_15108);
and U16662 (N_16662,N_14194,N_14364);
nor U16663 (N_16663,N_12972,N_13273);
nand U16664 (N_16664,N_15354,N_12895);
nor U16665 (N_16665,N_13442,N_13465);
or U16666 (N_16666,N_15188,N_14752);
xnor U16667 (N_16667,N_15007,N_14205);
and U16668 (N_16668,N_14014,N_12359);
and U16669 (N_16669,N_14710,N_13268);
nor U16670 (N_16670,N_14635,N_13419);
nor U16671 (N_16671,N_13287,N_15990);
nand U16672 (N_16672,N_15034,N_12430);
nor U16673 (N_16673,N_12280,N_14555);
and U16674 (N_16674,N_12850,N_15770);
nor U16675 (N_16675,N_14745,N_15652);
nor U16676 (N_16676,N_15935,N_12546);
nand U16677 (N_16677,N_13434,N_12634);
or U16678 (N_16678,N_13222,N_15005);
nor U16679 (N_16679,N_14495,N_13433);
and U16680 (N_16680,N_15032,N_14134);
nand U16681 (N_16681,N_15803,N_14770);
xnor U16682 (N_16682,N_13207,N_13557);
nor U16683 (N_16683,N_13812,N_13092);
or U16684 (N_16684,N_12128,N_14111);
xnor U16685 (N_16685,N_14361,N_14747);
nand U16686 (N_16686,N_13581,N_15071);
xnor U16687 (N_16687,N_14415,N_13388);
nor U16688 (N_16688,N_15335,N_15441);
nand U16689 (N_16689,N_13666,N_13106);
nand U16690 (N_16690,N_15424,N_15027);
nand U16691 (N_16691,N_12561,N_15462);
nor U16692 (N_16692,N_12828,N_14470);
or U16693 (N_16693,N_14360,N_12793);
nand U16694 (N_16694,N_14253,N_15292);
xor U16695 (N_16695,N_14316,N_12369);
xnor U16696 (N_16696,N_12823,N_15015);
nand U16697 (N_16697,N_12028,N_12691);
xnor U16698 (N_16698,N_15395,N_13548);
nor U16699 (N_16699,N_13962,N_15024);
and U16700 (N_16700,N_14483,N_15725);
and U16701 (N_16701,N_14509,N_12781);
nand U16702 (N_16702,N_12349,N_14169);
nor U16703 (N_16703,N_15592,N_15376);
or U16704 (N_16704,N_14515,N_12616);
and U16705 (N_16705,N_14697,N_13495);
xnor U16706 (N_16706,N_12453,N_12434);
nand U16707 (N_16707,N_14142,N_13209);
or U16708 (N_16708,N_14136,N_15616);
and U16709 (N_16709,N_14677,N_12107);
xor U16710 (N_16710,N_13250,N_15920);
nand U16711 (N_16711,N_12910,N_12724);
xor U16712 (N_16712,N_13486,N_15103);
and U16713 (N_16713,N_13697,N_13569);
xnor U16714 (N_16714,N_14628,N_14266);
xor U16715 (N_16715,N_12097,N_15166);
xnor U16716 (N_16716,N_13650,N_12766);
nand U16717 (N_16717,N_14390,N_12010);
nor U16718 (N_16718,N_13535,N_12314);
xnor U16719 (N_16719,N_13773,N_13499);
and U16720 (N_16720,N_15529,N_14388);
or U16721 (N_16721,N_14327,N_14522);
or U16722 (N_16722,N_13585,N_13934);
nor U16723 (N_16723,N_12775,N_12649);
and U16724 (N_16724,N_12321,N_13769);
nor U16725 (N_16725,N_12820,N_13185);
nor U16726 (N_16726,N_14780,N_14772);
xnor U16727 (N_16727,N_15458,N_14353);
xnor U16728 (N_16728,N_14022,N_12624);
nor U16729 (N_16729,N_13621,N_13439);
nand U16730 (N_16730,N_14895,N_12460);
nor U16731 (N_16731,N_15175,N_15290);
nor U16732 (N_16732,N_15124,N_14820);
or U16733 (N_16733,N_13004,N_12587);
or U16734 (N_16734,N_14758,N_14243);
or U16735 (N_16735,N_14501,N_12564);
and U16736 (N_16736,N_15982,N_13766);
xor U16737 (N_16737,N_13874,N_13785);
nand U16738 (N_16738,N_12254,N_13480);
xnor U16739 (N_16739,N_13992,N_12332);
or U16740 (N_16740,N_12396,N_13625);
nor U16741 (N_16741,N_15176,N_15819);
xnor U16742 (N_16742,N_13151,N_14478);
nand U16743 (N_16743,N_13016,N_12797);
or U16744 (N_16744,N_13941,N_13449);
nand U16745 (N_16745,N_14044,N_12959);
xnor U16746 (N_16746,N_15438,N_15541);
xnor U16747 (N_16747,N_14252,N_15276);
xnor U16748 (N_16748,N_12909,N_15229);
nor U16749 (N_16749,N_12440,N_14805);
nand U16750 (N_16750,N_12899,N_13608);
nand U16751 (N_16751,N_13565,N_12983);
or U16752 (N_16752,N_13085,N_14734);
nand U16753 (N_16753,N_15632,N_15353);
or U16754 (N_16754,N_12184,N_12362);
and U16755 (N_16755,N_13079,N_13121);
xnor U16756 (N_16756,N_15841,N_15307);
or U16757 (N_16757,N_14623,N_12733);
or U16758 (N_16758,N_14506,N_13430);
nor U16759 (N_16759,N_12001,N_14984);
xnor U16760 (N_16760,N_13429,N_13921);
nor U16761 (N_16761,N_15318,N_12970);
xnor U16762 (N_16762,N_13472,N_12220);
or U16763 (N_16763,N_14790,N_13255);
nand U16764 (N_16764,N_15254,N_14510);
or U16765 (N_16765,N_14152,N_15056);
or U16766 (N_16766,N_15425,N_12255);
nand U16767 (N_16767,N_14439,N_14086);
xor U16768 (N_16768,N_12041,N_15493);
xor U16769 (N_16769,N_12844,N_14696);
or U16770 (N_16770,N_12611,N_13318);
and U16771 (N_16771,N_12442,N_13084);
nor U16772 (N_16772,N_14597,N_12473);
nand U16773 (N_16773,N_12888,N_15428);
xor U16774 (N_16774,N_13108,N_12883);
nor U16775 (N_16775,N_14121,N_15834);
nor U16776 (N_16776,N_13320,N_12617);
xor U16777 (N_16777,N_14675,N_15185);
and U16778 (N_16778,N_13017,N_13703);
or U16779 (N_16779,N_12651,N_15028);
nand U16780 (N_16780,N_15063,N_12083);
or U16781 (N_16781,N_15617,N_14823);
and U16782 (N_16782,N_14357,N_13408);
nand U16783 (N_16783,N_13624,N_14552);
xor U16784 (N_16784,N_12846,N_13233);
xor U16785 (N_16785,N_15194,N_13528);
nor U16786 (N_16786,N_12696,N_12989);
nand U16787 (N_16787,N_12490,N_15760);
nor U16788 (N_16788,N_13554,N_14171);
or U16789 (N_16789,N_15295,N_13604);
nand U16790 (N_16790,N_13381,N_14011);
nor U16791 (N_16791,N_12462,N_14941);
nor U16792 (N_16792,N_14940,N_15488);
and U16793 (N_16793,N_14765,N_14905);
nand U16794 (N_16794,N_15267,N_15863);
and U16795 (N_16795,N_12743,N_15125);
nand U16796 (N_16796,N_14746,N_14742);
nand U16797 (N_16797,N_13579,N_13760);
nand U16798 (N_16798,N_13592,N_14618);
xor U16799 (N_16799,N_15274,N_13922);
nand U16800 (N_16800,N_12261,N_13409);
nand U16801 (N_16801,N_15422,N_12009);
nor U16802 (N_16802,N_15629,N_12759);
xnor U16803 (N_16803,N_12238,N_15877);
nor U16804 (N_16804,N_14997,N_15532);
nand U16805 (N_16805,N_13136,N_15408);
nand U16806 (N_16806,N_12142,N_14901);
and U16807 (N_16807,N_14866,N_13961);
or U16808 (N_16808,N_12865,N_12494);
or U16809 (N_16809,N_14582,N_13145);
and U16810 (N_16810,N_13444,N_12737);
or U16811 (N_16811,N_12305,N_14709);
and U16812 (N_16812,N_14235,N_15086);
and U16813 (N_16813,N_12536,N_13547);
xor U16814 (N_16814,N_12020,N_12788);
and U16815 (N_16815,N_13086,N_12642);
and U16816 (N_16816,N_12047,N_14154);
xnor U16817 (N_16817,N_15715,N_14349);
nand U16818 (N_16818,N_13348,N_14716);
and U16819 (N_16819,N_13208,N_15643);
or U16820 (N_16820,N_13767,N_13162);
xnor U16821 (N_16821,N_14000,N_14913);
or U16822 (N_16822,N_15706,N_13306);
xnor U16823 (N_16823,N_14281,N_12342);
and U16824 (N_16824,N_12809,N_13981);
and U16825 (N_16825,N_15875,N_15003);
nand U16826 (N_16826,N_12177,N_15519);
and U16827 (N_16827,N_12463,N_13669);
nand U16828 (N_16828,N_12045,N_13076);
and U16829 (N_16829,N_12003,N_13718);
and U16830 (N_16830,N_14295,N_14318);
nand U16831 (N_16831,N_15757,N_13481);
nor U16832 (N_16832,N_13033,N_13193);
and U16833 (N_16833,N_13467,N_12814);
nand U16834 (N_16834,N_14774,N_13761);
or U16835 (N_16835,N_15928,N_13716);
and U16836 (N_16836,N_14204,N_14273);
xor U16837 (N_16837,N_13301,N_13764);
and U16838 (N_16838,N_15921,N_15213);
or U16839 (N_16839,N_15876,N_15794);
and U16840 (N_16840,N_12038,N_12554);
xnor U16841 (N_16841,N_12997,N_14546);
xor U16842 (N_16842,N_12287,N_12603);
or U16843 (N_16843,N_12919,N_15387);
or U16844 (N_16844,N_15008,N_12878);
nand U16845 (N_16845,N_15496,N_12786);
and U16846 (N_16846,N_15691,N_14191);
or U16847 (N_16847,N_12545,N_14976);
or U16848 (N_16848,N_13405,N_12667);
xor U16849 (N_16849,N_15703,N_12778);
nor U16850 (N_16850,N_12647,N_14951);
and U16851 (N_16851,N_13267,N_13933);
nand U16852 (N_16852,N_12148,N_14562);
nor U16853 (N_16853,N_12378,N_14687);
nand U16854 (N_16854,N_14081,N_13870);
nor U16855 (N_16855,N_13702,N_15347);
nor U16856 (N_16856,N_14026,N_15859);
nand U16857 (N_16857,N_12161,N_13404);
nand U16858 (N_16858,N_12390,N_12070);
and U16859 (N_16859,N_13355,N_12697);
xnor U16860 (N_16860,N_12412,N_14184);
nand U16861 (N_16861,N_12610,N_15064);
or U16862 (N_16862,N_14185,N_15992);
or U16863 (N_16863,N_14581,N_15198);
xor U16864 (N_16864,N_15825,N_15145);
or U16865 (N_16865,N_13792,N_14212);
xnor U16866 (N_16866,N_15420,N_13271);
xor U16867 (N_16867,N_13441,N_15612);
nand U16868 (N_16868,N_13918,N_12375);
or U16869 (N_16869,N_14982,N_12175);
xor U16870 (N_16870,N_15780,N_14727);
xor U16871 (N_16871,N_15500,N_13660);
and U16872 (N_16872,N_14153,N_13184);
xor U16873 (N_16873,N_15170,N_12374);
and U16874 (N_16874,N_12969,N_13580);
or U16875 (N_16875,N_13105,N_14368);
or U16876 (N_16876,N_13602,N_15722);
and U16877 (N_16877,N_15916,N_13060);
and U16878 (N_16878,N_14097,N_15186);
nand U16879 (N_16879,N_12614,N_12784);
nand U16880 (N_16880,N_13944,N_12335);
nand U16881 (N_16881,N_14580,N_12776);
nand U16882 (N_16882,N_15922,N_13676);
and U16883 (N_16883,N_12181,N_15896);
nor U16884 (N_16884,N_14764,N_15978);
nand U16885 (N_16885,N_14567,N_12749);
nor U16886 (N_16886,N_12196,N_15215);
nor U16887 (N_16887,N_14222,N_15504);
and U16888 (N_16888,N_13931,N_15389);
or U16889 (N_16889,N_14989,N_15572);
or U16890 (N_16890,N_15469,N_15320);
xnor U16891 (N_16891,N_14655,N_15752);
xnor U16892 (N_16892,N_13483,N_15138);
or U16893 (N_16893,N_13783,N_12952);
and U16894 (N_16894,N_12543,N_12389);
xor U16895 (N_16895,N_13176,N_13534);
and U16896 (N_16896,N_15611,N_15094);
nor U16897 (N_16897,N_13545,N_15128);
or U16898 (N_16898,N_14731,N_14354);
nor U16899 (N_16899,N_14659,N_14725);
nor U16900 (N_16900,N_12941,N_13031);
nor U16901 (N_16901,N_13936,N_12761);
or U16902 (N_16902,N_13685,N_15601);
and U16903 (N_16903,N_12703,N_15113);
nor U16904 (N_16904,N_13309,N_14374);
nand U16905 (N_16905,N_15790,N_12847);
xnor U16906 (N_16906,N_12141,N_12423);
and U16907 (N_16907,N_14428,N_14471);
xor U16908 (N_16908,N_14646,N_15631);
and U16909 (N_16909,N_12772,N_13029);
or U16910 (N_16910,N_14937,N_14719);
or U16911 (N_16911,N_13310,N_13173);
xor U16912 (N_16912,N_14030,N_15105);
or U16913 (N_16913,N_14355,N_14944);
nand U16914 (N_16914,N_12267,N_14143);
and U16915 (N_16915,N_14715,N_14445);
nor U16916 (N_16916,N_14145,N_12167);
xor U16917 (N_16917,N_13988,N_15471);
nand U16918 (N_16918,N_15690,N_13326);
xnor U16919 (N_16919,N_12861,N_15902);
and U16920 (N_16920,N_14183,N_14500);
and U16921 (N_16921,N_15308,N_15838);
or U16922 (N_16922,N_15090,N_14084);
and U16923 (N_16923,N_15673,N_12113);
xor U16924 (N_16924,N_15668,N_15802);
nand U16925 (N_16925,N_15577,N_13259);
nand U16926 (N_16926,N_13501,N_12578);
nand U16927 (N_16927,N_15897,N_12081);
or U16928 (N_16928,N_12986,N_12627);
and U16929 (N_16929,N_15874,N_13626);
nor U16930 (N_16930,N_14069,N_12263);
xor U16931 (N_16931,N_13496,N_15661);
xor U16932 (N_16932,N_13862,N_13782);
xor U16933 (N_16933,N_15671,N_14966);
nor U16934 (N_16934,N_14867,N_15012);
and U16935 (N_16935,N_12496,N_15871);
and U16936 (N_16936,N_15460,N_14784);
and U16937 (N_16937,N_12407,N_15173);
and U16938 (N_16938,N_14756,N_12284);
nand U16939 (N_16939,N_15815,N_12595);
nand U16940 (N_16940,N_15891,N_15686);
nor U16941 (N_16941,N_15432,N_13248);
and U16942 (N_16942,N_14180,N_13586);
xor U16943 (N_16943,N_15678,N_12744);
nor U16944 (N_16944,N_14684,N_15956);
xor U16945 (N_16945,N_14638,N_13677);
or U16946 (N_16946,N_15786,N_15879);
xor U16947 (N_16947,N_12379,N_15899);
nor U16948 (N_16948,N_12738,N_15649);
and U16949 (N_16949,N_13678,N_14300);
and U16950 (N_16950,N_15775,N_14423);
and U16951 (N_16951,N_14908,N_13120);
nand U16952 (N_16952,N_14718,N_13509);
and U16953 (N_16953,N_15169,N_14883);
and U16954 (N_16954,N_13164,N_12487);
nand U16955 (N_16955,N_14891,N_12943);
and U16956 (N_16956,N_12219,N_12073);
and U16957 (N_16957,N_14328,N_15769);
or U16958 (N_16958,N_15081,N_13276);
and U16959 (N_16959,N_13160,N_15351);
xor U16960 (N_16960,N_14743,N_12988);
or U16961 (N_16961,N_13653,N_13200);
nand U16962 (N_16962,N_14645,N_15487);
xnor U16963 (N_16963,N_13871,N_13630);
nor U16964 (N_16964,N_15074,N_15379);
xor U16965 (N_16965,N_13018,N_14968);
nand U16966 (N_16966,N_15523,N_15756);
xor U16967 (N_16967,N_12656,N_12562);
nor U16968 (N_16968,N_15409,N_15744);
nor U16969 (N_16969,N_12782,N_12310);
xor U16970 (N_16970,N_12840,N_12356);
nor U16971 (N_16971,N_14860,N_12050);
or U16972 (N_16972,N_13887,N_15804);
and U16973 (N_16973,N_13482,N_15476);
nand U16974 (N_16974,N_14507,N_14397);
nor U16975 (N_16975,N_13424,N_13313);
and U16976 (N_16976,N_15700,N_13402);
and U16977 (N_16977,N_15326,N_12503);
nor U16978 (N_16978,N_12057,N_13749);
nor U16979 (N_16979,N_13420,N_13284);
and U16980 (N_16980,N_12689,N_13058);
or U16981 (N_16981,N_14461,N_12625);
nand U16982 (N_16982,N_14608,N_12720);
and U16983 (N_16983,N_14930,N_12849);
and U16984 (N_16984,N_15079,N_14654);
nand U16985 (N_16985,N_12399,N_15180);
and U16986 (N_16986,N_13742,N_13642);
or U16987 (N_16987,N_12639,N_14691);
nor U16988 (N_16988,N_14003,N_15991);
or U16989 (N_16989,N_14685,N_13498);
xor U16990 (N_16990,N_15293,N_12180);
or U16991 (N_16991,N_13291,N_12266);
nor U16992 (N_16992,N_13283,N_13103);
nand U16993 (N_16993,N_14898,N_12913);
or U16994 (N_16994,N_12560,N_13715);
nor U16995 (N_16995,N_14492,N_15745);
xnor U16996 (N_16996,N_15092,N_12140);
and U16997 (N_16997,N_15448,N_12752);
nor U16998 (N_16998,N_12694,N_15772);
nor U16999 (N_16999,N_15864,N_15766);
xor U17000 (N_17000,N_12537,N_12122);
nand U17001 (N_17001,N_12228,N_12510);
and U17002 (N_17002,N_15009,N_15768);
or U17003 (N_17003,N_15852,N_15765);
nor U17004 (N_17004,N_13244,N_14652);
nor U17005 (N_17005,N_12192,N_13603);
nor U17006 (N_17006,N_15256,N_15613);
or U17007 (N_17007,N_15352,N_14664);
nand U17008 (N_17008,N_12386,N_13078);
and U17009 (N_17009,N_12195,N_13674);
xor U17010 (N_17010,N_14616,N_14768);
and U17011 (N_17011,N_15994,N_14407);
or U17012 (N_17012,N_12433,N_13272);
and U17013 (N_17013,N_13050,N_15202);
or U17014 (N_17014,N_13360,N_15660);
or U17015 (N_17015,N_12105,N_13489);
xnor U17016 (N_17016,N_14876,N_13541);
xnor U17017 (N_17017,N_14933,N_14600);
nand U17018 (N_17018,N_13098,N_15936);
nand U17019 (N_17019,N_14612,N_14484);
and U17020 (N_17020,N_15052,N_12394);
nor U17021 (N_17021,N_12500,N_13032);
or U17022 (N_17022,N_14900,N_13838);
nand U17023 (N_17023,N_15929,N_12514);
nor U17024 (N_17024,N_14376,N_12934);
nand U17025 (N_17025,N_14851,N_15573);
xnor U17026 (N_17026,N_14682,N_14110);
nand U17027 (N_17027,N_14317,N_14135);
nand U17028 (N_17028,N_15155,N_12116);
xnor U17029 (N_17029,N_15339,N_15369);
nor U17030 (N_17030,N_13166,N_12672);
nand U17031 (N_17031,N_13022,N_13615);
or U17032 (N_17032,N_15372,N_12741);
xor U17033 (N_17033,N_14451,N_14124);
and U17034 (N_17034,N_14660,N_12526);
nor U17035 (N_17035,N_15350,N_14450);
and U17036 (N_17036,N_13027,N_13007);
nand U17037 (N_17037,N_15512,N_14383);
or U17038 (N_17038,N_12574,N_15817);
or U17039 (N_17039,N_12593,N_15406);
xnor U17040 (N_17040,N_14076,N_15130);
nand U17041 (N_17041,N_15246,N_15798);
nor U17042 (N_17042,N_14920,N_13993);
or U17043 (N_17043,N_13578,N_12371);
and U17044 (N_17044,N_13923,N_14249);
and U17045 (N_17045,N_13822,N_15456);
nor U17046 (N_17046,N_14543,N_12999);
xnor U17047 (N_17047,N_15100,N_13361);
nor U17048 (N_17048,N_13957,N_14524);
nor U17049 (N_17049,N_15820,N_12277);
nand U17050 (N_17050,N_12568,N_15261);
and U17051 (N_17051,N_12327,N_15397);
nand U17052 (N_17052,N_15676,N_14286);
and U17053 (N_17053,N_13850,N_15653);
and U17054 (N_17054,N_15099,N_14297);
nor U17055 (N_17055,N_12885,N_12866);
xor U17056 (N_17056,N_13406,N_12982);
and U17057 (N_17057,N_15514,N_15472);
nor U17058 (N_17058,N_13011,N_14890);
nor U17059 (N_17059,N_15865,N_14671);
or U17060 (N_17060,N_14012,N_12832);
nor U17061 (N_17061,N_15013,N_15078);
xnor U17062 (N_17062,N_12218,N_15386);
nand U17063 (N_17063,N_15377,N_12702);
and U17064 (N_17064,N_13042,N_13290);
and U17065 (N_17065,N_13857,N_12903);
nand U17066 (N_17066,N_13315,N_14735);
nand U17067 (N_17067,N_14093,N_15893);
or U17068 (N_17068,N_12427,N_14041);
nor U17069 (N_17069,N_14299,N_13800);
or U17070 (N_17070,N_12319,N_14814);
nor U17071 (N_17071,N_13448,N_13241);
or U17072 (N_17072,N_15227,N_14728);
nor U17073 (N_17073,N_15245,N_12204);
nand U17074 (N_17074,N_14066,N_14598);
xor U17075 (N_17075,N_15836,N_13943);
xnor U17076 (N_17076,N_13971,N_15407);
nand U17077 (N_17077,N_12178,N_14626);
nor U17078 (N_17078,N_15932,N_13211);
xor U17079 (N_17079,N_13851,N_15085);
nor U17080 (N_17080,N_13885,N_13225);
xor U17081 (N_17081,N_13794,N_14493);
or U17082 (N_17082,N_12630,N_14133);
and U17083 (N_17083,N_13040,N_15459);
xor U17084 (N_17084,N_13411,N_12117);
nand U17085 (N_17085,N_15174,N_14513);
nand U17086 (N_17086,N_14188,N_13330);
or U17087 (N_17087,N_14840,N_13471);
and U17088 (N_17088,N_13333,N_14661);
nor U17089 (N_17089,N_15651,N_15679);
and U17090 (N_17090,N_13477,N_14934);
or U17091 (N_17091,N_15382,N_14822);
xnor U17092 (N_17092,N_12658,N_13046);
nor U17093 (N_17093,N_13346,N_12406);
and U17094 (N_17094,N_15135,N_15521);
or U17095 (N_17095,N_14414,N_13728);
nand U17096 (N_17096,N_14352,N_15020);
and U17097 (N_17097,N_14434,N_13261);
or U17098 (N_17098,N_14894,N_13784);
nand U17099 (N_17099,N_12484,N_14609);
nor U17100 (N_17100,N_12346,N_13627);
or U17101 (N_17101,N_15908,N_14329);
or U17102 (N_17102,N_12833,N_13314);
and U17103 (N_17103,N_15597,N_13180);
xor U17104 (N_17104,N_14648,N_13443);
xnor U17105 (N_17105,N_14576,N_14481);
xnor U17106 (N_17106,N_13112,N_12698);
and U17107 (N_17107,N_13095,N_14242);
nand U17108 (N_17108,N_15622,N_13880);
or U17109 (N_17109,N_15867,N_13295);
xor U17110 (N_17110,N_12380,N_13257);
and U17111 (N_17111,N_15023,N_12118);
xnor U17112 (N_17112,N_12902,N_15945);
xor U17113 (N_17113,N_13679,N_14197);
or U17114 (N_17114,N_13643,N_14406);
nand U17115 (N_17115,N_13299,N_13458);
nand U17116 (N_17116,N_14282,N_13053);
and U17117 (N_17117,N_13030,N_14466);
and U17118 (N_17118,N_15499,N_15733);
xnor U17119 (N_17119,N_14256,N_12690);
nor U17120 (N_17120,N_14912,N_14494);
xnor U17121 (N_17121,N_13325,N_14070);
nor U17122 (N_17122,N_14649,N_14371);
xor U17123 (N_17123,N_12974,N_12156);
nand U17124 (N_17124,N_15791,N_15321);
nand U17125 (N_17125,N_15625,N_15507);
and U17126 (N_17126,N_14056,N_12395);
nor U17127 (N_17127,N_14566,N_14541);
xor U17128 (N_17128,N_12210,N_12700);
nor U17129 (N_17129,N_12547,N_13237);
nand U17130 (N_17130,N_15252,N_12084);
nand U17131 (N_17131,N_15434,N_14950);
xor U17132 (N_17132,N_13054,N_14578);
nor U17133 (N_17133,N_13293,N_13215);
and U17134 (N_17134,N_13994,N_15708);
or U17135 (N_17135,N_12730,N_13350);
xor U17136 (N_17136,N_13795,N_13390);
nand U17137 (N_17137,N_15648,N_14800);
nand U17138 (N_17138,N_15214,N_15667);
and U17139 (N_17139,N_14667,N_13610);
nand U17140 (N_17140,N_13397,N_14077);
and U17141 (N_17141,N_12907,N_12803);
xnor U17142 (N_17142,N_13278,N_13979);
xor U17143 (N_17143,N_15656,N_13289);
nor U17144 (N_17144,N_12007,N_15835);
and U17145 (N_17145,N_14220,N_15522);
nor U17146 (N_17146,N_15443,N_15095);
nor U17147 (N_17147,N_14531,N_15478);
nor U17148 (N_17148,N_12376,N_15750);
and U17149 (N_17149,N_13681,N_14278);
xnor U17150 (N_17150,N_15919,N_14786);
and U17151 (N_17151,N_12456,N_15647);
nor U17152 (N_17152,N_14196,N_12061);
and U17153 (N_17153,N_13984,N_13904);
xor U17154 (N_17154,N_14200,N_14219);
and U17155 (N_17155,N_12879,N_14365);
nand U17156 (N_17156,N_14857,N_12819);
nand U17157 (N_17157,N_12687,N_13967);
xnor U17158 (N_17158,N_12478,N_15510);
nand U17159 (N_17159,N_12629,N_15065);
nor U17160 (N_17160,N_12552,N_13028);
nand U17161 (N_17161,N_14311,N_12787);
or U17162 (N_17162,N_14606,N_13969);
xnor U17163 (N_17163,N_14771,N_13059);
and U17164 (N_17164,N_14268,N_14553);
xor U17165 (N_17165,N_12352,N_13186);
and U17166 (N_17166,N_12189,N_15277);
and U17167 (N_17167,N_13026,N_13848);
and U17168 (N_17168,N_12221,N_15506);
nand U17169 (N_17169,N_14519,N_12080);
and U17170 (N_17170,N_13297,N_12132);
xor U17171 (N_17171,N_13842,N_13551);
xor U17172 (N_17172,N_12727,N_13342);
and U17173 (N_17173,N_13633,N_12341);
nand U17174 (N_17174,N_12980,N_13537);
xor U17175 (N_17175,N_14887,N_15121);
nand U17176 (N_17176,N_12241,N_12734);
or U17177 (N_17177,N_12838,N_14821);
and U17178 (N_17178,N_13057,N_12044);
and U17179 (N_17179,N_12282,N_15106);
and U17180 (N_17180,N_15160,N_14759);
nand U17181 (N_17181,N_15304,N_15046);
xnor U17182 (N_17182,N_12072,N_13243);
or U17183 (N_17183,N_14897,N_14809);
or U17184 (N_17184,N_12719,N_13508);
and U17185 (N_17185,N_13161,N_13929);
nand U17186 (N_17186,N_15795,N_13512);
and U17187 (N_17187,N_12449,N_15627);
or U17188 (N_17188,N_14079,N_15457);
or U17189 (N_17189,N_12860,N_12215);
xor U17190 (N_17190,N_12621,N_15894);
nor U17191 (N_17191,N_13694,N_14053);
nor U17192 (N_17192,N_12347,N_13094);
or U17193 (N_17193,N_14151,N_12301);
nor U17194 (N_17194,N_13087,N_15163);
xor U17195 (N_17195,N_13919,N_13349);
nand U17196 (N_17196,N_14319,N_13307);
nor U17197 (N_17197,N_12528,N_14713);
and U17198 (N_17198,N_15315,N_14698);
and U17199 (N_17199,N_12060,N_12588);
or U17200 (N_17200,N_13920,N_12863);
or U17201 (N_17201,N_13099,N_15666);
nand U17202 (N_17202,N_14842,N_15785);
or U17203 (N_17203,N_13082,N_15682);
nand U17204 (N_17204,N_13707,N_12622);
or U17205 (N_17205,N_13587,N_13262);
and U17206 (N_17206,N_13066,N_14970);
xor U17207 (N_17207,N_12138,N_13747);
or U17208 (N_17208,N_15467,N_14283);
nand U17209 (N_17209,N_13741,N_14846);
or U17210 (N_17210,N_12100,N_14034);
nor U17211 (N_17211,N_13619,N_12367);
nor U17212 (N_17212,N_13892,N_14475);
xor U17213 (N_17213,N_14712,N_14815);
and U17214 (N_17214,N_12557,N_15626);
nor U17215 (N_17215,N_13378,N_15807);
or U17216 (N_17216,N_14425,N_13220);
xnor U17217 (N_17217,N_13985,N_13414);
or U17218 (N_17218,N_12739,N_12078);
and U17219 (N_17219,N_14091,N_12693);
nor U17220 (N_17220,N_14247,N_12958);
xor U17221 (N_17221,N_15654,N_12165);
xnor U17222 (N_17222,N_12090,N_14120);
and U17223 (N_17223,N_12216,N_15751);
nand U17224 (N_17224,N_15705,N_14977);
and U17225 (N_17225,N_15241,N_13213);
or U17226 (N_17226,N_13854,N_12294);
or U17227 (N_17227,N_14215,N_13072);
nor U17228 (N_17228,N_14721,N_13236);
and U17229 (N_17229,N_12465,N_12397);
xor U17230 (N_17230,N_15465,N_12657);
nand U17231 (N_17231,N_14488,N_13926);
nand U17232 (N_17232,N_12668,N_15934);
and U17233 (N_17233,N_15436,N_15985);
or U17234 (N_17234,N_14417,N_13876);
and U17235 (N_17235,N_13632,N_15687);
or U17236 (N_17236,N_14740,N_12732);
or U17237 (N_17237,N_15941,N_15112);
or U17238 (N_17238,N_15310,N_15182);
xnor U17239 (N_17239,N_13417,N_13859);
xnor U17240 (N_17240,N_14850,N_14408);
nor U17241 (N_17241,N_14594,N_12428);
xor U17242 (N_17242,N_14395,N_12262);
and U17243 (N_17243,N_13708,N_14819);
or U17244 (N_17244,N_14749,N_12383);
xnor U17245 (N_17245,N_14356,N_13865);
or U17246 (N_17246,N_14181,N_15083);
nor U17247 (N_17247,N_14284,N_14683);
xor U17248 (N_17248,N_12276,N_12098);
and U17249 (N_17249,N_12207,N_14186);
xor U17250 (N_17250,N_14918,N_14195);
and U17251 (N_17251,N_14886,N_13834);
xor U17252 (N_17252,N_13015,N_13748);
nand U17253 (N_17253,N_15737,N_13083);
xor U17254 (N_17254,N_14128,N_14599);
nor U17255 (N_17255,N_15330,N_13479);
nor U17256 (N_17256,N_12810,N_15580);
xor U17257 (N_17257,N_15004,N_12443);
nand U17258 (N_17258,N_14132,N_15118);
or U17259 (N_17259,N_12147,N_13175);
nor U17260 (N_17260,N_14826,N_14577);
nor U17261 (N_17261,N_15615,N_14248);
nor U17262 (N_17262,N_15590,N_15037);
xor U17263 (N_17263,N_13888,N_12469);
nand U17264 (N_17264,N_12126,N_14472);
and U17265 (N_17265,N_14585,N_12299);
nor U17266 (N_17266,N_14936,N_13853);
nor U17267 (N_17267,N_13006,N_13561);
nand U17268 (N_17268,N_12447,N_13701);
and U17269 (N_17269,N_15374,N_14879);
or U17270 (N_17270,N_14177,N_15442);
and U17271 (N_17271,N_15614,N_15235);
nor U17272 (N_17272,N_14536,N_13594);
nand U17273 (N_17273,N_12120,N_12676);
nor U17274 (N_17274,N_12441,N_15805);
nand U17275 (N_17275,N_14035,N_12912);
nand U17276 (N_17276,N_15855,N_12985);
nand U17277 (N_17277,N_13010,N_13886);
nor U17278 (N_17278,N_15553,N_12917);
or U17279 (N_17279,N_15618,N_12245);
nand U17280 (N_17280,N_12632,N_14853);
or U17281 (N_17281,N_14663,N_12115);
and U17282 (N_17282,N_12521,N_14491);
and U17283 (N_17283,N_12812,N_13351);
nor U17284 (N_17284,N_13597,N_15402);
nor U17285 (N_17285,N_14404,N_15299);
nor U17286 (N_17286,N_14279,N_12411);
nand U17287 (N_17287,N_13114,N_15482);
or U17288 (N_17288,N_14046,N_14617);
nand U17289 (N_17289,N_14817,N_12293);
and U17290 (N_17290,N_14099,N_12998);
xor U17291 (N_17291,N_13673,N_14213);
nand U17292 (N_17292,N_14881,N_13019);
or U17293 (N_17293,N_14877,N_13067);
nand U17294 (N_17294,N_12171,N_13035);
nor U17295 (N_17295,N_13682,N_14263);
xor U17296 (N_17296,N_13073,N_15637);
and U17297 (N_17297,N_14549,N_12608);
or U17298 (N_17298,N_13056,N_14653);
xnor U17299 (N_17299,N_12471,N_15526);
nor U17300 (N_17300,N_12862,N_15342);
and U17301 (N_17301,N_13577,N_14336);
or U17302 (N_17302,N_14490,N_13216);
nor U17303 (N_17303,N_13327,N_12843);
or U17304 (N_17304,N_14237,N_15451);
and U17305 (N_17305,N_12875,N_14999);
nand U17306 (N_17306,N_13288,N_12756);
xnor U17307 (N_17307,N_15427,N_15289);
nand U17308 (N_17308,N_15842,N_13191);
or U17309 (N_17309,N_13720,N_14342);
or U17310 (N_17310,N_12774,N_14463);
nor U17311 (N_17311,N_12459,N_15970);
nand U17312 (N_17312,N_14801,N_15549);
nand U17313 (N_17313,N_13196,N_12337);
and U17314 (N_17314,N_14480,N_15068);
and U17315 (N_17315,N_12920,N_15584);
and U17316 (N_17316,N_14477,N_12890);
nor U17317 (N_17317,N_12074,N_15849);
nor U17318 (N_17318,N_15429,N_15527);
and U17319 (N_17319,N_15147,N_12067);
nand U17320 (N_17320,N_13398,N_13454);
nor U17321 (N_17321,N_12768,N_13906);
and U17322 (N_17322,N_12343,N_14203);
xor U17323 (N_17323,N_14755,N_12715);
or U17324 (N_17324,N_12791,N_12008);
nand U17325 (N_17325,N_12480,N_14442);
nor U17326 (N_17326,N_15044,N_12963);
nor U17327 (N_17327,N_13964,N_15520);
xnor U17328 (N_17328,N_13968,N_14338);
nand U17329 (N_17329,N_12506,N_13118);
and U17330 (N_17330,N_14548,N_12716);
xor U17331 (N_17331,N_15126,N_15607);
or U17332 (N_17332,N_13963,N_12283);
and U17333 (N_17333,N_12758,N_12420);
and U17334 (N_17334,N_13908,N_14435);
and U17335 (N_17335,N_15193,N_13227);
xor U17336 (N_17336,N_13757,N_13358);
or U17337 (N_17337,N_12515,N_14845);
nor U17338 (N_17338,N_13735,N_15301);
xor U17339 (N_17339,N_12103,N_13601);
or U17340 (N_17340,N_15850,N_15779);
xnor U17341 (N_17341,N_14736,N_15093);
or U17342 (N_17342,N_15468,N_14864);
xnor U17343 (N_17343,N_15331,N_13232);
nand U17344 (N_17344,N_12949,N_14131);
nor U17345 (N_17345,N_14741,N_13172);
nor U17346 (N_17346,N_12680,N_12519);
or U17347 (N_17347,N_13855,N_12251);
nor U17348 (N_17348,N_13533,N_14199);
or U17349 (N_17349,N_15048,N_15951);
and U17350 (N_17350,N_15077,N_14346);
or U17351 (N_17351,N_12372,N_14052);
and U17352 (N_17352,N_15856,N_12771);
and U17353 (N_17353,N_14812,N_14264);
xnor U17354 (N_17354,N_13877,N_15940);
xor U17355 (N_17355,N_12684,N_13256);
and U17356 (N_17356,N_15923,N_13563);
nor U17357 (N_17357,N_13560,N_15489);
nand U17358 (N_17358,N_12984,N_15435);
xor U17359 (N_17359,N_15268,N_12091);
nor U17360 (N_17360,N_14115,N_15053);
nand U17361 (N_17361,N_12806,N_14087);
or U17362 (N_17362,N_13447,N_13178);
or U17363 (N_17363,N_14882,N_13075);
and U17364 (N_17364,N_13335,N_15684);
nand U17365 (N_17365,N_12170,N_12747);
xor U17366 (N_17366,N_12409,N_15464);
or U17367 (N_17367,N_12876,N_13598);
and U17368 (N_17368,N_14986,N_13319);
or U17369 (N_17369,N_13445,N_14717);
xnor U17370 (N_17370,N_12695,N_12187);
nor U17371 (N_17371,N_14457,N_13600);
xnor U17372 (N_17372,N_15533,N_15778);
or U17373 (N_17373,N_12016,N_14560);
nand U17374 (N_17374,N_14656,N_14103);
nor U17375 (N_17375,N_13550,N_15363);
nand U17376 (N_17376,N_13254,N_13778);
xor U17377 (N_17377,N_12918,N_12317);
nand U17378 (N_17378,N_14054,N_14426);
nand U17379 (N_17379,N_14911,N_15582);
nand U17380 (N_17380,N_15777,N_14929);
nor U17381 (N_17381,N_15120,N_14693);
nand U17382 (N_17382,N_14217,N_13543);
nand U17383 (N_17383,N_13531,N_12413);
or U17384 (N_17384,N_12109,N_15480);
nor U17385 (N_17385,N_12686,N_14290);
xnor U17386 (N_17386,N_13153,N_12837);
or U17387 (N_17387,N_14469,N_12867);
or U17388 (N_17388,N_15721,N_12807);
nand U17389 (N_17389,N_15736,N_12973);
nand U17390 (N_17390,N_14332,N_15901);
nor U17391 (N_17391,N_13146,N_15963);
nand U17392 (N_17392,N_12188,N_12155);
or U17393 (N_17393,N_14192,N_15084);
xnor U17394 (N_17394,N_15343,N_12232);
and U17395 (N_17395,N_13159,N_12790);
and U17396 (N_17396,N_12133,N_14474);
xnor U17397 (N_17397,N_12853,N_15153);
or U17398 (N_17398,N_14592,N_14917);
and U17399 (N_17399,N_14942,N_15713);
or U17400 (N_17400,N_12800,N_13640);
nand U17401 (N_17401,N_13337,N_13294);
nor U17402 (N_17402,N_13023,N_14651);
xnor U17403 (N_17403,N_13675,N_13881);
nor U17404 (N_17404,N_12124,N_12190);
or U17405 (N_17405,N_13117,N_15225);
and U17406 (N_17406,N_14269,N_12298);
and U17407 (N_17407,N_12445,N_12533);
xor U17408 (N_17408,N_14144,N_12544);
nor U17409 (N_17409,N_12290,N_12569);
and U17410 (N_17410,N_13553,N_15305);
nand U17411 (N_17411,N_12796,N_15447);
or U17412 (N_17412,N_12966,N_13591);
xor U17413 (N_17413,N_13768,N_12033);
xnor U17414 (N_17414,N_12707,N_14558);
and U17415 (N_17415,N_13989,N_12313);
and U17416 (N_17416,N_15851,N_15258);
or U17417 (N_17417,N_14019,N_14101);
nor U17418 (N_17418,N_13192,N_13183);
xnor U17419 (N_17419,N_15107,N_12363);
nand U17420 (N_17420,N_13229,N_13538);
nor U17421 (N_17421,N_12613,N_12857);
or U17422 (N_17422,N_14650,N_12311);
xnor U17423 (N_17423,N_15773,N_15463);
xnor U17424 (N_17424,N_12149,N_12524);
and U17425 (N_17425,N_12541,N_12306);
and U17426 (N_17426,N_12472,N_13462);
xor U17427 (N_17427,N_13008,N_12931);
xnor U17428 (N_17428,N_15731,N_14542);
nand U17429 (N_17429,N_14639,N_15968);
and U17430 (N_17430,N_13125,N_15880);
nor U17431 (N_17431,N_14487,N_12391);
and U17432 (N_17432,N_13611,N_14298);
xor U17433 (N_17433,N_14367,N_13612);
nand U17434 (N_17434,N_12357,N_14422);
nor U17435 (N_17435,N_13556,N_13081);
xor U17436 (N_17436,N_13100,N_13394);
nand U17437 (N_17437,N_15296,N_14497);
or U17438 (N_17438,N_12669,N_15334);
xnor U17439 (N_17439,N_15233,N_15375);
xor U17440 (N_17440,N_15559,N_13634);
nand U17441 (N_17441,N_14730,N_14787);
and U17442 (N_17442,N_12256,N_13503);
nand U17443 (N_17443,N_13436,N_15767);
xor U17444 (N_17444,N_14102,N_15132);
xnor U17445 (N_17445,N_15816,N_15184);
and U17446 (N_17446,N_12333,N_15242);
xnor U17447 (N_17447,N_12509,N_15783);
nor U17448 (N_17448,N_12708,N_14563);
and U17449 (N_17449,N_13638,N_12136);
and U17450 (N_17450,N_14227,N_12027);
xnor U17451 (N_17451,N_12706,N_14750);
and U17452 (N_17452,N_13282,N_15453);
xnor U17453 (N_17453,N_12789,N_12035);
nand U17454 (N_17454,N_15131,N_12477);
nand U17455 (N_17455,N_15219,N_13736);
and U17456 (N_17456,N_13978,N_14516);
and U17457 (N_17457,N_14036,N_15746);
and U17458 (N_17458,N_12818,N_15954);
and U17459 (N_17459,N_14382,N_13620);
nand U17460 (N_17460,N_13422,N_15575);
and U17461 (N_17461,N_12236,N_12069);
xor U17462 (N_17462,N_13817,N_14596);
nor U17463 (N_17463,N_15718,N_15516);
nand U17464 (N_17464,N_13605,N_15168);
and U17465 (N_17465,N_15231,N_15677);
nor U17466 (N_17466,N_12950,N_12729);
nor U17467 (N_17467,N_14140,N_13206);
nor U17468 (N_17468,N_15324,N_14836);
and U17469 (N_17469,N_12900,N_15837);
xnor U17470 (N_17470,N_13725,N_12401);
xor U17471 (N_17471,N_15530,N_13025);
or U17472 (N_17472,N_12736,N_13123);
xnor U17473 (N_17473,N_14149,N_13824);
and U17474 (N_17474,N_14722,N_12405);
or U17475 (N_17475,N_13464,N_15201);
and U17476 (N_17476,N_15384,N_14657);
or U17477 (N_17477,N_15505,N_12577);
and U17478 (N_17478,N_14310,N_15812);
nand U17479 (N_17479,N_12871,N_14574);
or U17480 (N_17480,N_15603,N_12059);
xor U17481 (N_17481,N_12887,N_14837);
nor U17482 (N_17482,N_14116,N_13686);
and U17483 (N_17483,N_13700,N_12435);
xnor U17484 (N_17484,N_14704,N_15906);
nand U17485 (N_17485,N_14631,N_15944);
or U17486 (N_17486,N_13755,N_15349);
nor U17487 (N_17487,N_15801,N_12765);
nand U17488 (N_17488,N_15265,N_14757);
or U17489 (N_17489,N_12655,N_14261);
and U17490 (N_17490,N_12598,N_13265);
nor U17491 (N_17491,N_12286,N_14723);
nor U17492 (N_17492,N_13379,N_12891);
xor U17493 (N_17493,N_14072,N_12418);
or U17494 (N_17494,N_14998,N_15758);
nand U17495 (N_17495,N_15965,N_12199);
and U17496 (N_17496,N_12804,N_15966);
nand U17497 (N_17497,N_13609,N_15764);
nand U17498 (N_17498,N_13354,N_13878);
or U17499 (N_17499,N_15860,N_15391);
and U17500 (N_17500,N_14669,N_12307);
nand U17501 (N_17501,N_13134,N_15799);
and U17502 (N_17502,N_12981,N_15957);
nand U17503 (N_17503,N_12451,N_12612);
nand U17504 (N_17504,N_15723,N_14238);
or U17505 (N_17505,N_13334,N_12458);
nand U17506 (N_17506,N_15141,N_15545);
and U17507 (N_17507,N_13109,N_15058);
or U17508 (N_17508,N_13304,N_13995);
and U17509 (N_17509,N_12661,N_12760);
nand U17510 (N_17510,N_13096,N_12403);
nor U17511 (N_17511,N_13502,N_12664);
or U17512 (N_17512,N_14946,N_14027);
xor U17513 (N_17513,N_13189,N_14239);
and U17514 (N_17514,N_12054,N_13546);
or U17515 (N_17515,N_13525,N_15925);
and U17516 (N_17516,N_13104,N_13144);
xor U17517 (N_17517,N_15136,N_13729);
and U17518 (N_17518,N_13706,N_12163);
or U17519 (N_17519,N_12252,N_13396);
or U17520 (N_17520,N_13530,N_15042);
or U17521 (N_17521,N_13721,N_14416);
nand U17522 (N_17522,N_14473,N_12025);
and U17523 (N_17523,N_15123,N_12942);
or U17524 (N_17524,N_15699,N_13300);
and U17525 (N_17525,N_13951,N_12031);
or U17526 (N_17526,N_12110,N_12179);
nand U17527 (N_17527,N_13418,N_12527);
or U17528 (N_17528,N_14708,N_13009);
nand U17529 (N_17529,N_14754,N_12130);
and U17530 (N_17530,N_13890,N_13239);
and U17531 (N_17531,N_14232,N_12102);
nor U17532 (N_17532,N_14230,N_14100);
and U17533 (N_17533,N_15208,N_13051);
and U17534 (N_17534,N_15417,N_12322);
and U17535 (N_17535,N_13787,N_14892);
and U17536 (N_17536,N_12881,N_15177);
and U17537 (N_17537,N_14366,N_13583);
xnor U17538 (N_17538,N_14190,N_13260);
xor U17539 (N_17539,N_12360,N_15598);
and U17540 (N_17540,N_12957,N_14302);
and U17541 (N_17541,N_15561,N_12448);
nor U17542 (N_17542,N_13302,N_12437);
and U17543 (N_17543,N_12264,N_13991);
nand U17544 (N_17544,N_13582,N_14692);
xor U17545 (N_17545,N_12750,N_15495);
and U17546 (N_17546,N_15070,N_15501);
or U17547 (N_17547,N_14344,N_15909);
and U17548 (N_17548,N_15204,N_14711);
or U17549 (N_17549,N_14873,N_15563);
nand U17550 (N_17550,N_13517,N_15337);
nor U17551 (N_17551,N_14139,N_15975);
nor U17552 (N_17552,N_13003,N_13214);
nor U17553 (N_17553,N_13217,N_15988);
nand U17554 (N_17554,N_12644,N_14334);
xor U17555 (N_17555,N_13450,N_15620);
nor U17556 (N_17556,N_13158,N_15748);
nor U17557 (N_17557,N_14673,N_14393);
xnor U17558 (N_17558,N_14508,N_14325);
xor U17559 (N_17559,N_13895,N_15761);
xnor U17560 (N_17560,N_12350,N_15316);
and U17561 (N_17561,N_12370,N_13945);
xor U17562 (N_17562,N_13401,N_12600);
nor U17563 (N_17563,N_12531,N_13910);
or U17564 (N_17564,N_15809,N_14292);
xnor U17565 (N_17565,N_12712,N_15082);
xnor U17566 (N_17566,N_15806,N_14779);
xor U17567 (N_17567,N_13126,N_13529);
nand U17568 (N_17568,N_12643,N_15393);
xnor U17569 (N_17569,N_14436,N_15414);
or U17570 (N_17570,N_13038,N_14945);
nor U17571 (N_17571,N_15142,N_14832);
nand U17572 (N_17572,N_14804,N_13407);
nor U17573 (N_17573,N_15275,N_13435);
and U17574 (N_17574,N_12633,N_15524);
and U17575 (N_17575,N_15759,N_12573);
and U17576 (N_17576,N_12088,N_15345);
and U17577 (N_17577,N_14971,N_13338);
nand U17578 (N_17578,N_14224,N_14350);
and U17579 (N_17579,N_15062,N_12137);
and U17580 (N_17580,N_12504,N_12064);
nor U17581 (N_17581,N_12377,N_14896);
nor U17582 (N_17582,N_13219,N_12145);
nand U17583 (N_17583,N_15440,N_13363);
nand U17584 (N_17584,N_13759,N_15634);
nor U17585 (N_17585,N_13392,N_14952);
xor U17586 (N_17586,N_13860,N_12637);
nand U17587 (N_17587,N_14778,N_14059);
xnor U17588 (N_17588,N_12235,N_12673);
xor U17589 (N_17589,N_14872,N_12012);
nor U17590 (N_17590,N_14798,N_13833);
or U17591 (N_17591,N_14107,N_14075);
nand U17592 (N_17592,N_12763,N_14098);
nand U17593 (N_17593,N_12665,N_13372);
nor U17594 (N_17594,N_12499,N_14005);
nand U17595 (N_17595,N_12662,N_12783);
xnor U17596 (N_17596,N_14956,N_13996);
or U17597 (N_17597,N_14777,N_12414);
or U17598 (N_17598,N_15662,N_13915);
xor U17599 (N_17599,N_13279,N_15205);
nand U17600 (N_17600,N_15693,N_14630);
nor U17601 (N_17601,N_14584,N_14955);
nor U17602 (N_17602,N_14972,N_12144);
xor U17603 (N_17603,N_15858,N_14008);
and U17604 (N_17604,N_12400,N_14557);
and U17605 (N_17605,N_15134,N_14799);
xor U17606 (N_17606,N_15567,N_12104);
nand U17607 (N_17607,N_14424,N_15672);
nor U17608 (N_17608,N_15306,N_15355);
nor U17609 (N_17609,N_15755,N_15854);
xnor U17610 (N_17610,N_14210,N_14983);
nor U17611 (N_17611,N_13810,N_15430);
nand U17612 (N_17612,N_12991,N_15528);
nand U17613 (N_17613,N_13077,N_13884);
nor U17614 (N_17614,N_15251,N_12623);
nor U17615 (N_17615,N_15285,N_12951);
xor U17616 (N_17616,N_14370,N_14392);
and U17617 (N_17617,N_13958,N_14216);
nand U17618 (N_17618,N_14518,N_15884);
nor U17619 (N_17619,N_12438,N_13247);
and U17620 (N_17620,N_12582,N_15596);
or U17621 (N_17621,N_12492,N_13693);
xnor U17622 (N_17622,N_13204,N_14159);
or U17623 (N_17623,N_15556,N_13323);
or U17624 (N_17624,N_14271,N_15240);
and U17625 (N_17625,N_14010,N_12551);
or U17626 (N_17626,N_13137,N_15914);
and U17627 (N_17627,N_13949,N_14208);
nand U17628 (N_17628,N_13616,N_12292);
nor U17629 (N_17629,N_15025,N_15564);
nor U17630 (N_17630,N_15630,N_12779);
nand U17631 (N_17631,N_12300,N_14496);
nand U17632 (N_17632,N_12929,N_13269);
nor U17633 (N_17633,N_13726,N_12579);
or U17634 (N_17634,N_13695,N_12237);
or U17635 (N_17635,N_15228,N_14396);
and U17636 (N_17636,N_13858,N_13347);
or U17637 (N_17637,N_12231,N_15050);
nand U17638 (N_17638,N_13613,N_14695);
nor U17639 (N_17639,N_12101,N_12315);
xor U17640 (N_17640,N_14051,N_13516);
xor U17641 (N_17641,N_15943,N_12382);
or U17642 (N_17642,N_14499,N_15057);
nand U17643 (N_17643,N_12037,N_15938);
nor U17644 (N_17644,N_15129,N_14225);
xnor U17645 (N_17645,N_12822,N_12799);
nand U17646 (N_17646,N_15749,N_13750);
nor U17647 (N_17647,N_13440,N_14959);
xor U17648 (N_17648,N_12169,N_15895);
or U17649 (N_17649,N_14198,N_14766);
nor U17650 (N_17650,N_14400,N_13635);
xnor U17651 (N_17651,N_15433,N_15689);
nor U17652 (N_17652,N_12051,N_12416);
xor U17653 (N_17653,N_12811,N_12605);
and U17654 (N_17654,N_15452,N_14776);
or U17655 (N_17655,N_12518,N_14796);
xor U17656 (N_17656,N_15466,N_12995);
nand U17657 (N_17657,N_15054,N_14512);
nor U17658 (N_17658,N_15993,N_14871);
nor U17659 (N_17659,N_15977,N_15683);
or U17660 (N_17660,N_14922,N_12956);
and U17661 (N_17661,N_13775,N_14889);
or U17662 (N_17662,N_15336,N_12710);
xor U17663 (N_17663,N_14733,N_12393);
nor U17664 (N_17664,N_13570,N_14172);
nand U17665 (N_17665,N_12209,N_12762);
xnor U17666 (N_17666,N_12628,N_12585);
nand U17667 (N_17667,N_14938,N_15300);
or U17668 (N_17668,N_14272,N_15669);
or U17669 (N_17669,N_15508,N_15534);
and U17670 (N_17670,N_12134,N_13522);
nand U17671 (N_17671,N_13111,N_13305);
nand U17672 (N_17672,N_14676,N_15444);
xor U17673 (N_17673,N_15309,N_13903);
nor U17674 (N_17674,N_15665,N_12939);
or U17675 (N_17675,N_13131,N_13376);
xnor U17676 (N_17676,N_12898,N_14554);
and U17677 (N_17677,N_14629,N_12592);
nand U17678 (N_17678,N_14240,N_14040);
and U17679 (N_17679,N_12955,N_12203);
nor U17680 (N_17680,N_13331,N_14254);
nand U17681 (N_17681,N_13368,N_13389);
nor U17682 (N_17682,N_15917,N_14544);
nor U17683 (N_17683,N_12735,N_14539);
or U17684 (N_17684,N_12488,N_15088);
nand U17685 (N_17685,N_14647,N_15635);
or U17686 (N_17686,N_14025,N_13765);
xnor U17687 (N_17687,N_13724,N_13332);
and U17688 (N_17688,N_15964,N_15833);
nor U17689 (N_17689,N_15845,N_14405);
xor U17690 (N_17690,N_15644,N_13296);
nand U17691 (N_17691,N_13584,N_15642);
xor U17692 (N_17692,N_13714,N_12817);
xnor U17693 (N_17693,N_15585,N_13843);
and U17694 (N_17694,N_15359,N_13088);
xnor U17695 (N_17695,N_13900,N_15030);
xor U17696 (N_17696,N_15226,N_13839);
and U17697 (N_17697,N_15811,N_15344);
nor U17698 (N_17698,N_13188,N_13727);
xnor U17699 (N_17699,N_13667,N_12645);
or U17700 (N_17700,N_15385,N_12387);
or U17701 (N_17701,N_12461,N_13836);
or U17702 (N_17702,N_13875,N_15399);
nor U17703 (N_17703,N_12185,N_15624);
xor U17704 (N_17704,N_13329,N_12678);
nand U17705 (N_17705,N_15403,N_15903);
xnor U17706 (N_17706,N_13044,N_13791);
and U17707 (N_17707,N_14794,N_12108);
nand U17708 (N_17708,N_12172,N_15913);
nand U17709 (N_17709,N_12160,N_13492);
or U17710 (N_17710,N_12429,N_12249);
nor U17711 (N_17711,N_13497,N_12079);
nor U17712 (N_17712,N_13831,N_15479);
xor U17713 (N_17713,N_12297,N_15255);
xor U17714 (N_17714,N_15157,N_15595);
nand U17715 (N_17715,N_13359,N_12275);
xor U17716 (N_17716,N_13340,N_13142);
nand U17717 (N_17717,N_14304,N_14438);
nor U17718 (N_17718,N_13607,N_12670);
xor U17719 (N_17719,N_12168,N_13052);
nand U17720 (N_17720,N_13637,N_14511);
xor U17721 (N_17721,N_12965,N_12908);
nor U17722 (N_17722,N_15143,N_12601);
nand U17723 (N_17723,N_13649,N_15942);
nor U17724 (N_17724,N_14162,N_13737);
xor U17725 (N_17725,N_15485,N_13863);
or U17726 (N_17726,N_14039,N_15473);
or U17727 (N_17727,N_12845,N_14369);
xnor U17728 (N_17728,N_13071,N_15358);
and U17729 (N_17729,N_13093,N_15981);
nor U17730 (N_17730,N_13861,N_15317);
or U17731 (N_17731,N_12571,N_12258);
or U17732 (N_17732,N_12501,N_14957);
xnor U17733 (N_17733,N_14386,N_12638);
or U17734 (N_17734,N_15872,N_15972);
nand U17735 (N_17735,N_14064,N_12692);
nor U17736 (N_17736,N_14032,N_13129);
or U17737 (N_17737,N_14166,N_12757);
or U17738 (N_17738,N_15771,N_13829);
xnor U17739 (N_17739,N_14085,N_15594);
or U17740 (N_17740,N_13799,N_14904);
xor U17741 (N_17741,N_12575,N_12049);
xnor U17742 (N_17742,N_15657,N_14275);
nand U17743 (N_17743,N_15288,N_14861);
nand U17744 (N_17744,N_12896,N_12162);
nand U17745 (N_17745,N_14486,N_15073);
or U17746 (N_17746,N_15055,N_13972);
nand U17747 (N_17747,N_12967,N_12398);
nand U17748 (N_17748,N_13937,N_15589);
nor U17749 (N_17749,N_15704,N_13940);
and U17750 (N_17750,N_13617,N_13845);
and U17751 (N_17751,N_12722,N_12026);
xor U17752 (N_17752,N_13930,N_14680);
nand U17753 (N_17753,N_15571,N_14525);
nor U17754 (N_17754,N_12466,N_15303);
and U17755 (N_17755,N_15818,N_12482);
and U17756 (N_17756,N_15392,N_14586);
or U17757 (N_17757,N_12928,N_12549);
or U17758 (N_17758,N_14427,N_14802);
and U17759 (N_17759,N_15102,N_13788);
and U17760 (N_17760,N_12303,N_15861);
nor U17761 (N_17761,N_14537,N_12214);
or U17762 (N_17762,N_14849,N_12848);
nand U17763 (N_17763,N_15313,N_15069);
nor U17764 (N_17764,N_13571,N_13549);
or U17765 (N_17765,N_12897,N_15974);
or U17766 (N_17766,N_12446,N_15608);
and U17767 (N_17767,N_12151,N_14775);
nand U17768 (N_17768,N_13518,N_12491);
or U17769 (N_17769,N_15340,N_13135);
and U17770 (N_17770,N_15696,N_12660);
and U17771 (N_17771,N_15411,N_14452);
and U17772 (N_17772,N_15808,N_13203);
xor U17773 (N_17773,N_13352,N_12279);
nand U17774 (N_17774,N_15171,N_13428);
nor U17775 (N_17775,N_15273,N_13156);
nor U17776 (N_17776,N_13558,N_13974);
or U17777 (N_17777,N_13312,N_14964);
or U17778 (N_17778,N_12924,N_12836);
nor U17779 (N_17779,N_13383,N_12039);
or U17780 (N_17780,N_14921,N_14029);
nand U17781 (N_17781,N_13240,N_12166);
nor U17782 (N_17782,N_12513,N_14440);
and U17783 (N_17783,N_14296,N_15370);
nor U17784 (N_17784,N_12808,N_13264);
and U17785 (N_17785,N_14981,N_12093);
or U17786 (N_17786,N_14906,N_12048);
and U17787 (N_17787,N_15019,N_12043);
and U17788 (N_17788,N_15967,N_12542);
or U17789 (N_17789,N_14080,N_12248);
xnor U17790 (N_17790,N_12927,N_14561);
or U17791 (N_17791,N_12522,N_12619);
xor U17792 (N_17792,N_13460,N_14288);
and U17793 (N_17793,N_15655,N_13336);
or U17794 (N_17794,N_12688,N_12679);
xor U17795 (N_17795,N_15338,N_12916);
or U17796 (N_17796,N_15291,N_14468);
or U17797 (N_17797,N_12486,N_12852);
nor U17798 (N_17798,N_14773,N_14380);
and U17799 (N_17799,N_13651,N_12011);
nor U17800 (N_17800,N_14241,N_12006);
nor U17801 (N_17801,N_13080,N_14421);
xor U17802 (N_17802,N_13384,N_15697);
nand U17803 (N_17803,N_15832,N_14033);
nor U17804 (N_17804,N_14389,N_12563);
and U17805 (N_17805,N_14978,N_12058);
nor U17806 (N_17806,N_14277,N_13124);
nand U17807 (N_17807,N_12244,N_14529);
nand U17808 (N_17808,N_13656,N_14954);
nand U17809 (N_17809,N_13523,N_13303);
nor U17810 (N_17810,N_13973,N_14568);
and U17811 (N_17811,N_14862,N_15739);
or U17812 (N_17812,N_15260,N_15381);
nor U17813 (N_17813,N_15139,N_13856);
xor U17814 (N_17814,N_13841,N_14666);
xor U17815 (N_17815,N_15959,N_12296);
and U17816 (N_17816,N_14322,N_14844);
and U17817 (N_17817,N_12590,N_15793);
xnor U17818 (N_17818,N_13476,N_12052);
xor U17819 (N_17819,N_13955,N_14359);
or U17820 (N_17820,N_13740,N_15550);
nand U17821 (N_17821,N_14109,N_13652);
xor U17822 (N_17822,N_14347,N_13891);
nand U17823 (N_17823,N_14932,N_14854);
nand U17824 (N_17824,N_14206,N_15924);
nor U17825 (N_17825,N_14893,N_13672);
nand U17826 (N_17826,N_15284,N_15144);
nor U17827 (N_17827,N_13416,N_12609);
nor U17828 (N_17828,N_15552,N_14985);
or U17829 (N_17829,N_13494,N_15249);
nand U17830 (N_17830,N_15060,N_12529);
xnor U17831 (N_17831,N_14094,N_12348);
or U17832 (N_17832,N_12566,N_13639);
xor U17833 (N_17833,N_14018,N_15312);
xnor U17834 (N_17834,N_15823,N_14119);
xnor U17835 (N_17835,N_13474,N_15247);
nor U17836 (N_17836,N_12023,N_15623);
and U17837 (N_17837,N_14048,N_13174);
or U17838 (N_17838,N_13663,N_13524);
nor U17839 (N_17839,N_12699,N_15605);
nand U17840 (N_17840,N_15840,N_15658);
nor U17841 (N_17841,N_13559,N_14935);
xor U17842 (N_17842,N_14965,N_12032);
xnor U17843 (N_17843,N_14620,N_13999);
or U17844 (N_17844,N_12714,N_13956);
and U17845 (N_17845,N_12626,N_12197);
xnor U17846 (N_17846,N_13321,N_12474);
xor U17847 (N_17847,N_15784,N_13743);
nand U17848 (N_17848,N_14498,N_12200);
nor U17849 (N_17849,N_12243,N_12211);
xnor U17850 (N_17850,N_14340,N_15248);
nand U17851 (N_17851,N_15080,N_14875);
nand U17852 (N_17852,N_14433,N_13771);
xor U17853 (N_17853,N_15986,N_14943);
nand U17854 (N_17854,N_13070,N_12233);
nor U17855 (N_17855,N_13739,N_13804);
or U17856 (N_17856,N_14391,N_13593);
and U17857 (N_17857,N_13709,N_14987);
or U17858 (N_17858,N_15882,N_13762);
nand U17859 (N_17859,N_12068,N_15537);
and U17860 (N_17860,N_15546,N_14447);
or U17861 (N_17861,N_13670,N_12053);
nand U17862 (N_17862,N_14732,N_15640);
nand U17863 (N_17863,N_12893,N_15455);
nand U17864 (N_17864,N_14874,N_13370);
nand U17865 (N_17865,N_12234,N_13039);
or U17866 (N_17866,N_12576,N_15604);
xnor U17867 (N_17867,N_14674,N_14095);
and U17868 (N_17868,N_15000,N_12558);
and U17869 (N_17869,N_14255,N_12021);
xnor U17870 (N_17870,N_14170,N_14903);
nand U17871 (N_17871,N_13770,N_12066);
and U17872 (N_17872,N_12344,N_13024);
xor U17873 (N_17873,N_12431,N_15199);
xor U17874 (N_17874,N_12532,N_14246);
nor U17875 (N_17875,N_14164,N_12479);
and U17876 (N_17876,N_15405,N_12535);
or U17877 (N_17877,N_12559,N_14607);
xor U17878 (N_17878,N_13683,N_15675);
or U17879 (N_17879,N_13641,N_15283);
or U17880 (N_17880,N_15727,N_13595);
or U17881 (N_17881,N_14839,N_13809);
and U17882 (N_17882,N_15927,N_12798);
nand U17883 (N_17883,N_12894,N_13661);
nand U17884 (N_17884,N_15159,N_12520);
nand U17885 (N_17885,N_15502,N_13927);
and U17886 (N_17886,N_13588,N_14960);
nand U17887 (N_17887,N_12953,N_15999);
and U17888 (N_17888,N_15591,N_15211);
xnor U17889 (N_17889,N_13212,N_15539);
xnor U17890 (N_17890,N_13488,N_13542);
nor U17891 (N_17891,N_13515,N_12444);
nand U17892 (N_17892,N_13453,N_15412);
xnor U17893 (N_17893,N_14614,N_15203);
and U17894 (N_17894,N_15762,N_12323);
xnor U17895 (N_17895,N_15404,N_14013);
and U17896 (N_17896,N_13490,N_14910);
nand U17897 (N_17897,N_15741,N_14919);
nor U17898 (N_17898,N_13377,N_12034);
xnor U17899 (N_17899,N_12996,N_12940);
xnor U17900 (N_17900,N_12174,N_12273);
or U17901 (N_17901,N_13438,N_14337);
nor U17902 (N_17902,N_13116,N_12511);
and U17903 (N_17903,N_12092,N_13511);
or U17904 (N_17904,N_12331,N_13484);
or U17905 (N_17905,N_14748,N_14001);
nand U17906 (N_17906,N_15574,N_15494);
or U17907 (N_17907,N_12517,N_13224);
nor U17908 (N_17908,N_12923,N_15333);
nand U17909 (N_17909,N_15789,N_14818);
xnor U17910 (N_17910,N_14534,N_15844);
nor U17911 (N_17911,N_13948,N_13867);
and U17912 (N_17912,N_13796,N_12930);
nand U17913 (N_17913,N_14411,N_13119);
and U17914 (N_17914,N_12454,N_12268);
nor U17915 (N_17915,N_15814,N_14074);
or U17916 (N_17916,N_12153,N_14335);
xor U17917 (N_17917,N_14155,N_15210);
or U17918 (N_17918,N_15357,N_14726);
or U17919 (N_17919,N_15262,N_14564);
or U17920 (N_17920,N_15535,N_12572);
and U17921 (N_17921,N_15222,N_14245);
xnor U17922 (N_17922,N_12539,N_14378);
nand U17923 (N_17923,N_14744,N_12498);
nor U17924 (N_17924,N_15886,N_13385);
xnor U17925 (N_17925,N_15431,N_12213);
nor U17926 (N_17926,N_15332,N_14830);
nand U17927 (N_17927,N_12468,N_13179);
or U17928 (N_17928,N_12960,N_15051);
nand U17929 (N_17929,N_15323,N_12977);
or U17930 (N_17930,N_12152,N_13939);
xnor U17931 (N_17931,N_15562,N_15196);
nor U17932 (N_17932,N_15076,N_15398);
nor U17933 (N_17933,N_15588,N_15949);
nand U17934 (N_17934,N_12205,N_12127);
nand U17935 (N_17935,N_14089,N_13230);
nor U17936 (N_17936,N_15960,N_15821);
nand U17937 (N_17937,N_12685,N_12711);
nor U17938 (N_17938,N_15979,N_13140);
or U17939 (N_17939,N_12962,N_14505);
or U17940 (N_17940,N_15091,N_12014);
nand U17941 (N_17941,N_13231,N_15364);
and U17942 (N_17942,N_15039,N_13751);
nand U17943 (N_17943,N_14314,N_12555);
nand U17944 (N_17944,N_14274,N_13493);
xor U17945 (N_17945,N_12334,N_14176);
or U17946 (N_17946,N_15119,N_15663);
nor U17947 (N_17947,N_15593,N_14055);
or U17948 (N_17948,N_14974,N_15380);
xnor U17949 (N_17949,N_14925,N_14622);
and U17950 (N_17950,N_13311,N_15868);
or U17951 (N_17951,N_13873,N_15191);
and U17952 (N_17952,N_15953,N_14141);
nor U17953 (N_17953,N_12483,N_15362);
and U17954 (N_17954,N_15907,N_15239);
and U17955 (N_17955,N_12591,N_14379);
xor U17956 (N_17956,N_13195,N_14207);
nor U17957 (N_17957,N_12056,N_13457);
and U17958 (N_17958,N_15889,N_12111);
or U17959 (N_17959,N_14067,N_13235);
nor U17960 (N_17960,N_13328,N_13068);
nand U17961 (N_17961,N_13521,N_13959);
or U17962 (N_17962,N_12911,N_13045);
and U17963 (N_17963,N_13205,N_13932);
and U17964 (N_17964,N_13141,N_15800);
nor U17965 (N_17965,N_12709,N_12345);
nor U17966 (N_17966,N_15890,N_13690);
and U17967 (N_17967,N_12119,N_15698);
nor U17968 (N_17968,N_13167,N_12230);
or U17969 (N_17969,N_14437,N_12648);
nand U17970 (N_17970,N_12764,N_12550);
and U17971 (N_17971,N_14315,N_12567);
nand U17972 (N_17972,N_15606,N_14402);
xnor U17973 (N_17973,N_12476,N_14545);
nand U17974 (N_17974,N_15702,N_14948);
or U17975 (N_17975,N_14517,N_13468);
nor U17976 (N_17976,N_14221,N_15551);
nand U17977 (N_17977,N_12071,N_12726);
xnor U17978 (N_17978,N_14262,N_12880);
nor U17979 (N_17979,N_13816,N_12858);
nand U17980 (N_17980,N_15149,N_14572);
and U17981 (N_17981,N_15641,N_13781);
nor U17982 (N_17982,N_15394,N_15645);
nor U17983 (N_17983,N_12792,N_13463);
nor U17984 (N_17984,N_13564,N_15221);
nand U17985 (N_17985,N_12507,N_13982);
nor U17986 (N_17986,N_15010,N_15707);
nor U17987 (N_17987,N_13723,N_12250);
nor U17988 (N_17988,N_13596,N_12746);
nand U17989 (N_17989,N_15878,N_12886);
nand U17990 (N_17990,N_12869,N_14165);
or U17991 (N_17991,N_15726,N_12425);
nand U17992 (N_17992,N_15792,N_13047);
xnor U17993 (N_17993,N_15543,N_15224);
nand U17994 (N_17994,N_13263,N_15067);
nor U17995 (N_17995,N_14643,N_14961);
or U17996 (N_17996,N_14753,N_13181);
nor U17997 (N_17997,N_14678,N_13000);
or U17998 (N_17998,N_12947,N_15035);
nand U17999 (N_17999,N_14071,N_15518);
or U18000 (N_18000,N_14994,N_13195);
and U18001 (N_18001,N_13835,N_13739);
and U18002 (N_18002,N_12275,N_14176);
xor U18003 (N_18003,N_12739,N_14192);
nor U18004 (N_18004,N_15617,N_12832);
xnor U18005 (N_18005,N_15742,N_15031);
or U18006 (N_18006,N_13799,N_14605);
or U18007 (N_18007,N_12385,N_14779);
nand U18008 (N_18008,N_14219,N_12403);
nand U18009 (N_18009,N_12498,N_15693);
nor U18010 (N_18010,N_12521,N_12549);
or U18011 (N_18011,N_12506,N_15135);
nand U18012 (N_18012,N_12376,N_15463);
or U18013 (N_18013,N_14048,N_13056);
nor U18014 (N_18014,N_15230,N_14171);
nand U18015 (N_18015,N_14602,N_15946);
or U18016 (N_18016,N_13335,N_15120);
xnor U18017 (N_18017,N_14648,N_15622);
and U18018 (N_18018,N_13497,N_13847);
nor U18019 (N_18019,N_12981,N_15370);
nand U18020 (N_18020,N_12320,N_15431);
xnor U18021 (N_18021,N_15715,N_13812);
xor U18022 (N_18022,N_15266,N_12139);
nor U18023 (N_18023,N_13237,N_12296);
or U18024 (N_18024,N_13505,N_14973);
or U18025 (N_18025,N_12796,N_15114);
and U18026 (N_18026,N_14902,N_12972);
or U18027 (N_18027,N_15131,N_15513);
nor U18028 (N_18028,N_14549,N_14733);
nor U18029 (N_18029,N_14383,N_12548);
nor U18030 (N_18030,N_13808,N_12584);
and U18031 (N_18031,N_15076,N_13021);
nand U18032 (N_18032,N_13333,N_15768);
nor U18033 (N_18033,N_14461,N_13280);
nor U18034 (N_18034,N_14724,N_14160);
and U18035 (N_18035,N_14736,N_15787);
and U18036 (N_18036,N_14795,N_14749);
and U18037 (N_18037,N_12172,N_12913);
nor U18038 (N_18038,N_13422,N_12445);
nand U18039 (N_18039,N_14513,N_13019);
and U18040 (N_18040,N_12984,N_12410);
or U18041 (N_18041,N_14589,N_12335);
xnor U18042 (N_18042,N_14313,N_15247);
nor U18043 (N_18043,N_14162,N_15663);
xor U18044 (N_18044,N_12950,N_15702);
or U18045 (N_18045,N_14119,N_12244);
nand U18046 (N_18046,N_12049,N_15209);
nand U18047 (N_18047,N_15273,N_12401);
and U18048 (N_18048,N_15664,N_13868);
or U18049 (N_18049,N_15105,N_12826);
xnor U18050 (N_18050,N_13174,N_15511);
nand U18051 (N_18051,N_14101,N_15221);
xor U18052 (N_18052,N_15407,N_13621);
and U18053 (N_18053,N_13259,N_13621);
or U18054 (N_18054,N_13767,N_14227);
and U18055 (N_18055,N_14718,N_12590);
nor U18056 (N_18056,N_13764,N_15556);
or U18057 (N_18057,N_15501,N_14510);
and U18058 (N_18058,N_15369,N_15775);
and U18059 (N_18059,N_12945,N_15008);
nor U18060 (N_18060,N_14318,N_15300);
nand U18061 (N_18061,N_13023,N_12893);
and U18062 (N_18062,N_12451,N_12591);
xnor U18063 (N_18063,N_12804,N_12807);
nor U18064 (N_18064,N_12211,N_13277);
or U18065 (N_18065,N_14890,N_15363);
nand U18066 (N_18066,N_15395,N_13126);
nand U18067 (N_18067,N_14176,N_14665);
nor U18068 (N_18068,N_15649,N_14730);
or U18069 (N_18069,N_14564,N_13719);
nor U18070 (N_18070,N_13020,N_14793);
or U18071 (N_18071,N_15859,N_13950);
nor U18072 (N_18072,N_13040,N_14578);
and U18073 (N_18073,N_13563,N_15045);
or U18074 (N_18074,N_12686,N_12234);
nor U18075 (N_18075,N_13242,N_13737);
and U18076 (N_18076,N_13349,N_12538);
nor U18077 (N_18077,N_13295,N_12008);
xnor U18078 (N_18078,N_15488,N_14953);
nand U18079 (N_18079,N_14069,N_14779);
nand U18080 (N_18080,N_14216,N_13899);
xnor U18081 (N_18081,N_14757,N_14587);
nand U18082 (N_18082,N_14997,N_15298);
xor U18083 (N_18083,N_12046,N_15677);
xnor U18084 (N_18084,N_13620,N_12386);
or U18085 (N_18085,N_13083,N_14272);
nor U18086 (N_18086,N_14900,N_15550);
xor U18087 (N_18087,N_15734,N_12586);
xor U18088 (N_18088,N_14251,N_15881);
xnor U18089 (N_18089,N_12900,N_15958);
xor U18090 (N_18090,N_14154,N_13419);
or U18091 (N_18091,N_13560,N_15313);
or U18092 (N_18092,N_12847,N_13115);
nand U18093 (N_18093,N_12478,N_14482);
or U18094 (N_18094,N_12570,N_12028);
and U18095 (N_18095,N_14369,N_14301);
nand U18096 (N_18096,N_14180,N_12388);
or U18097 (N_18097,N_12334,N_15759);
xor U18098 (N_18098,N_12975,N_14267);
or U18099 (N_18099,N_14030,N_13744);
nor U18100 (N_18100,N_13593,N_14338);
nor U18101 (N_18101,N_15760,N_12166);
nand U18102 (N_18102,N_13276,N_14465);
nor U18103 (N_18103,N_13849,N_12907);
and U18104 (N_18104,N_14371,N_12653);
nor U18105 (N_18105,N_14930,N_14688);
or U18106 (N_18106,N_14563,N_13022);
nor U18107 (N_18107,N_12820,N_13047);
or U18108 (N_18108,N_13048,N_12472);
nand U18109 (N_18109,N_14930,N_12513);
nand U18110 (N_18110,N_14625,N_12906);
nand U18111 (N_18111,N_12660,N_12094);
and U18112 (N_18112,N_15545,N_15927);
or U18113 (N_18113,N_15683,N_15754);
and U18114 (N_18114,N_13994,N_14086);
xor U18115 (N_18115,N_14349,N_13361);
xnor U18116 (N_18116,N_14521,N_12735);
nor U18117 (N_18117,N_12003,N_13856);
xnor U18118 (N_18118,N_14422,N_15857);
nand U18119 (N_18119,N_15955,N_13827);
nor U18120 (N_18120,N_12336,N_14701);
nor U18121 (N_18121,N_14821,N_13150);
or U18122 (N_18122,N_15738,N_14569);
xnor U18123 (N_18123,N_12155,N_15735);
nand U18124 (N_18124,N_14322,N_14856);
xnor U18125 (N_18125,N_14679,N_13973);
xor U18126 (N_18126,N_15036,N_14627);
or U18127 (N_18127,N_12086,N_13626);
or U18128 (N_18128,N_13013,N_14373);
or U18129 (N_18129,N_15332,N_12283);
nand U18130 (N_18130,N_14702,N_14981);
nor U18131 (N_18131,N_14847,N_14737);
or U18132 (N_18132,N_15985,N_12816);
nand U18133 (N_18133,N_13886,N_12468);
nand U18134 (N_18134,N_15582,N_14068);
nand U18135 (N_18135,N_13171,N_12609);
or U18136 (N_18136,N_15819,N_13975);
or U18137 (N_18137,N_12363,N_12025);
nor U18138 (N_18138,N_13700,N_14686);
xnor U18139 (N_18139,N_14094,N_15263);
or U18140 (N_18140,N_14954,N_13618);
or U18141 (N_18141,N_14650,N_12828);
nand U18142 (N_18142,N_14146,N_15404);
xnor U18143 (N_18143,N_14570,N_13095);
and U18144 (N_18144,N_15588,N_14057);
and U18145 (N_18145,N_14180,N_14153);
nand U18146 (N_18146,N_12052,N_14576);
or U18147 (N_18147,N_14756,N_15792);
nand U18148 (N_18148,N_15278,N_15877);
and U18149 (N_18149,N_15236,N_13858);
nor U18150 (N_18150,N_12130,N_14334);
nand U18151 (N_18151,N_12034,N_14791);
nand U18152 (N_18152,N_12966,N_15812);
nor U18153 (N_18153,N_12741,N_13947);
nor U18154 (N_18154,N_15242,N_13550);
nand U18155 (N_18155,N_15878,N_13691);
nor U18156 (N_18156,N_14744,N_14684);
nand U18157 (N_18157,N_12942,N_12142);
nor U18158 (N_18158,N_14533,N_14855);
or U18159 (N_18159,N_12439,N_14216);
or U18160 (N_18160,N_15598,N_15461);
or U18161 (N_18161,N_13443,N_14811);
nor U18162 (N_18162,N_15295,N_14004);
or U18163 (N_18163,N_13390,N_13538);
nor U18164 (N_18164,N_15956,N_12553);
and U18165 (N_18165,N_12254,N_12218);
and U18166 (N_18166,N_12891,N_15231);
and U18167 (N_18167,N_15797,N_14407);
nand U18168 (N_18168,N_14567,N_14019);
nor U18169 (N_18169,N_15951,N_15019);
nand U18170 (N_18170,N_14040,N_15935);
nor U18171 (N_18171,N_15206,N_14774);
nand U18172 (N_18172,N_14655,N_14640);
xnor U18173 (N_18173,N_15446,N_12402);
nand U18174 (N_18174,N_12120,N_13429);
nand U18175 (N_18175,N_14698,N_12420);
and U18176 (N_18176,N_14350,N_12154);
and U18177 (N_18177,N_14583,N_12176);
or U18178 (N_18178,N_13536,N_12152);
nand U18179 (N_18179,N_13315,N_15654);
nor U18180 (N_18180,N_14247,N_12385);
or U18181 (N_18181,N_13275,N_14936);
xor U18182 (N_18182,N_12123,N_14102);
or U18183 (N_18183,N_14615,N_12533);
xnor U18184 (N_18184,N_15336,N_15164);
xor U18185 (N_18185,N_15676,N_14605);
nor U18186 (N_18186,N_13571,N_14677);
nand U18187 (N_18187,N_14954,N_14178);
and U18188 (N_18188,N_13261,N_12007);
xor U18189 (N_18189,N_13765,N_15908);
or U18190 (N_18190,N_13139,N_15181);
nand U18191 (N_18191,N_14076,N_12857);
nor U18192 (N_18192,N_12389,N_14735);
nor U18193 (N_18193,N_14081,N_13665);
xnor U18194 (N_18194,N_13053,N_15567);
nor U18195 (N_18195,N_13222,N_13429);
xor U18196 (N_18196,N_13794,N_13486);
xor U18197 (N_18197,N_15666,N_12676);
nor U18198 (N_18198,N_14369,N_15076);
nand U18199 (N_18199,N_14993,N_14318);
xor U18200 (N_18200,N_15949,N_12706);
nor U18201 (N_18201,N_15320,N_12203);
and U18202 (N_18202,N_12534,N_15622);
and U18203 (N_18203,N_12329,N_13398);
and U18204 (N_18204,N_15669,N_15962);
xor U18205 (N_18205,N_14582,N_15276);
nand U18206 (N_18206,N_15379,N_15835);
xor U18207 (N_18207,N_12314,N_12855);
xnor U18208 (N_18208,N_13636,N_15154);
nor U18209 (N_18209,N_15406,N_12956);
nand U18210 (N_18210,N_12058,N_14808);
xnor U18211 (N_18211,N_14877,N_12277);
nand U18212 (N_18212,N_12910,N_14586);
nor U18213 (N_18213,N_14531,N_13017);
nor U18214 (N_18214,N_14216,N_14740);
and U18215 (N_18215,N_12427,N_12134);
or U18216 (N_18216,N_12231,N_14394);
nor U18217 (N_18217,N_15094,N_13127);
or U18218 (N_18218,N_13797,N_13067);
and U18219 (N_18219,N_14822,N_14863);
nand U18220 (N_18220,N_15188,N_13057);
and U18221 (N_18221,N_13768,N_14937);
nand U18222 (N_18222,N_13955,N_15425);
xnor U18223 (N_18223,N_12659,N_14906);
or U18224 (N_18224,N_13506,N_14530);
nand U18225 (N_18225,N_12932,N_13168);
or U18226 (N_18226,N_13843,N_14272);
or U18227 (N_18227,N_12841,N_14361);
nand U18228 (N_18228,N_15613,N_13919);
and U18229 (N_18229,N_13210,N_15328);
or U18230 (N_18230,N_14641,N_14386);
xor U18231 (N_18231,N_15204,N_12264);
and U18232 (N_18232,N_15213,N_12565);
xor U18233 (N_18233,N_13718,N_13932);
nand U18234 (N_18234,N_13607,N_13527);
nor U18235 (N_18235,N_14584,N_14240);
nand U18236 (N_18236,N_13438,N_12034);
nand U18237 (N_18237,N_15761,N_13763);
or U18238 (N_18238,N_13772,N_14766);
or U18239 (N_18239,N_12854,N_13008);
xor U18240 (N_18240,N_13000,N_15694);
and U18241 (N_18241,N_15759,N_12184);
nand U18242 (N_18242,N_15467,N_13627);
nand U18243 (N_18243,N_14368,N_12570);
xor U18244 (N_18244,N_13706,N_15305);
and U18245 (N_18245,N_14712,N_12850);
and U18246 (N_18246,N_14334,N_13064);
or U18247 (N_18247,N_15765,N_14913);
and U18248 (N_18248,N_12903,N_14284);
and U18249 (N_18249,N_14745,N_15367);
nor U18250 (N_18250,N_14543,N_13486);
xnor U18251 (N_18251,N_12476,N_14348);
nor U18252 (N_18252,N_15749,N_14184);
xnor U18253 (N_18253,N_15190,N_14700);
nand U18254 (N_18254,N_13062,N_13596);
xor U18255 (N_18255,N_15755,N_14255);
nor U18256 (N_18256,N_12060,N_15455);
or U18257 (N_18257,N_15669,N_13103);
nand U18258 (N_18258,N_14208,N_14157);
nor U18259 (N_18259,N_15843,N_15994);
and U18260 (N_18260,N_14455,N_12038);
nand U18261 (N_18261,N_14997,N_14096);
nand U18262 (N_18262,N_15151,N_13445);
nand U18263 (N_18263,N_12030,N_14995);
or U18264 (N_18264,N_12824,N_14140);
nand U18265 (N_18265,N_12329,N_13361);
and U18266 (N_18266,N_14188,N_13031);
and U18267 (N_18267,N_15039,N_15541);
nand U18268 (N_18268,N_15390,N_15395);
nand U18269 (N_18269,N_12230,N_12131);
xnor U18270 (N_18270,N_15768,N_15685);
and U18271 (N_18271,N_13396,N_15377);
and U18272 (N_18272,N_15708,N_14243);
or U18273 (N_18273,N_12322,N_12837);
or U18274 (N_18274,N_12969,N_14617);
xnor U18275 (N_18275,N_14990,N_13034);
nand U18276 (N_18276,N_13165,N_12549);
nand U18277 (N_18277,N_13688,N_15727);
nor U18278 (N_18278,N_14738,N_12903);
xor U18279 (N_18279,N_14886,N_15978);
or U18280 (N_18280,N_13036,N_15830);
or U18281 (N_18281,N_14286,N_12593);
and U18282 (N_18282,N_13832,N_15434);
and U18283 (N_18283,N_12823,N_12363);
nor U18284 (N_18284,N_15789,N_13102);
or U18285 (N_18285,N_15602,N_14582);
nand U18286 (N_18286,N_15336,N_13608);
xor U18287 (N_18287,N_15163,N_14083);
or U18288 (N_18288,N_12882,N_14566);
xnor U18289 (N_18289,N_13680,N_14935);
and U18290 (N_18290,N_13207,N_14575);
or U18291 (N_18291,N_14753,N_13571);
nor U18292 (N_18292,N_15173,N_14917);
and U18293 (N_18293,N_14705,N_12491);
and U18294 (N_18294,N_14549,N_13869);
or U18295 (N_18295,N_13291,N_13350);
nor U18296 (N_18296,N_15360,N_14488);
nor U18297 (N_18297,N_15906,N_12874);
and U18298 (N_18298,N_13474,N_13743);
nand U18299 (N_18299,N_13001,N_14678);
or U18300 (N_18300,N_15900,N_12924);
or U18301 (N_18301,N_13552,N_12208);
nor U18302 (N_18302,N_14787,N_13952);
nand U18303 (N_18303,N_15544,N_15441);
xnor U18304 (N_18304,N_12924,N_13219);
and U18305 (N_18305,N_12933,N_13602);
or U18306 (N_18306,N_14334,N_13454);
nand U18307 (N_18307,N_14033,N_12708);
xor U18308 (N_18308,N_13179,N_14149);
nor U18309 (N_18309,N_12743,N_15560);
and U18310 (N_18310,N_14604,N_15316);
and U18311 (N_18311,N_13702,N_14542);
nor U18312 (N_18312,N_13106,N_12554);
nand U18313 (N_18313,N_12223,N_14399);
nor U18314 (N_18314,N_15958,N_12839);
or U18315 (N_18315,N_13624,N_12952);
nor U18316 (N_18316,N_13834,N_15729);
xor U18317 (N_18317,N_13419,N_12967);
xnor U18318 (N_18318,N_14857,N_12704);
nand U18319 (N_18319,N_13610,N_12261);
or U18320 (N_18320,N_13823,N_15658);
xor U18321 (N_18321,N_14816,N_12040);
or U18322 (N_18322,N_15684,N_13492);
nand U18323 (N_18323,N_12741,N_12317);
nor U18324 (N_18324,N_15979,N_14058);
and U18325 (N_18325,N_14876,N_14174);
xor U18326 (N_18326,N_15752,N_15738);
nor U18327 (N_18327,N_15891,N_13236);
xor U18328 (N_18328,N_14342,N_12062);
and U18329 (N_18329,N_15052,N_14074);
or U18330 (N_18330,N_13751,N_13906);
xor U18331 (N_18331,N_15583,N_12227);
nor U18332 (N_18332,N_15995,N_15338);
or U18333 (N_18333,N_12422,N_12043);
xnor U18334 (N_18334,N_13404,N_15474);
or U18335 (N_18335,N_13385,N_12113);
or U18336 (N_18336,N_14452,N_14338);
and U18337 (N_18337,N_15674,N_13709);
nor U18338 (N_18338,N_12326,N_13676);
nand U18339 (N_18339,N_15502,N_15794);
nor U18340 (N_18340,N_14212,N_13501);
xnor U18341 (N_18341,N_13189,N_14606);
nand U18342 (N_18342,N_12479,N_12754);
nor U18343 (N_18343,N_15155,N_14162);
nand U18344 (N_18344,N_12590,N_13551);
xor U18345 (N_18345,N_13995,N_14252);
xnor U18346 (N_18346,N_12347,N_15831);
and U18347 (N_18347,N_13043,N_12325);
and U18348 (N_18348,N_12236,N_14105);
xor U18349 (N_18349,N_15365,N_12576);
and U18350 (N_18350,N_13794,N_15965);
nand U18351 (N_18351,N_14148,N_12830);
nand U18352 (N_18352,N_13384,N_14178);
nor U18353 (N_18353,N_14070,N_14811);
or U18354 (N_18354,N_15743,N_13612);
or U18355 (N_18355,N_13485,N_15297);
xor U18356 (N_18356,N_15464,N_15166);
or U18357 (N_18357,N_13126,N_15919);
and U18358 (N_18358,N_13754,N_13146);
nor U18359 (N_18359,N_15356,N_14975);
xor U18360 (N_18360,N_12309,N_14061);
xnor U18361 (N_18361,N_13377,N_15374);
xnor U18362 (N_18362,N_14057,N_14013);
and U18363 (N_18363,N_14902,N_14890);
or U18364 (N_18364,N_13032,N_15960);
nor U18365 (N_18365,N_12816,N_15494);
xnor U18366 (N_18366,N_13780,N_15205);
and U18367 (N_18367,N_12142,N_14447);
or U18368 (N_18368,N_15083,N_15470);
or U18369 (N_18369,N_15239,N_15895);
and U18370 (N_18370,N_15029,N_12598);
nor U18371 (N_18371,N_13279,N_13603);
or U18372 (N_18372,N_15537,N_13650);
nand U18373 (N_18373,N_14665,N_12958);
or U18374 (N_18374,N_12059,N_12908);
or U18375 (N_18375,N_13290,N_14550);
and U18376 (N_18376,N_15678,N_13844);
or U18377 (N_18377,N_14277,N_14860);
nand U18378 (N_18378,N_14549,N_15004);
nor U18379 (N_18379,N_14227,N_13367);
xnor U18380 (N_18380,N_13392,N_13720);
nor U18381 (N_18381,N_13948,N_15802);
xnor U18382 (N_18382,N_15062,N_14893);
nand U18383 (N_18383,N_13913,N_12579);
xnor U18384 (N_18384,N_14102,N_12696);
xor U18385 (N_18385,N_15599,N_12989);
nor U18386 (N_18386,N_14795,N_13615);
xnor U18387 (N_18387,N_15323,N_15067);
xor U18388 (N_18388,N_12718,N_14730);
xor U18389 (N_18389,N_13789,N_15188);
nor U18390 (N_18390,N_12148,N_13102);
nor U18391 (N_18391,N_13028,N_15764);
xor U18392 (N_18392,N_12133,N_14149);
xor U18393 (N_18393,N_13942,N_14384);
nand U18394 (N_18394,N_15342,N_15833);
nor U18395 (N_18395,N_15441,N_15112);
xor U18396 (N_18396,N_15227,N_12767);
nor U18397 (N_18397,N_14589,N_13908);
nor U18398 (N_18398,N_13213,N_12307);
or U18399 (N_18399,N_13232,N_13086);
nor U18400 (N_18400,N_13819,N_12937);
xor U18401 (N_18401,N_12039,N_14061);
and U18402 (N_18402,N_14689,N_15739);
nand U18403 (N_18403,N_15554,N_15565);
nor U18404 (N_18404,N_12410,N_14057);
nand U18405 (N_18405,N_15785,N_15705);
or U18406 (N_18406,N_13318,N_13761);
xnor U18407 (N_18407,N_14766,N_15592);
nor U18408 (N_18408,N_13198,N_14254);
or U18409 (N_18409,N_12814,N_14569);
or U18410 (N_18410,N_15171,N_15296);
or U18411 (N_18411,N_12035,N_15106);
and U18412 (N_18412,N_15541,N_14844);
xor U18413 (N_18413,N_15881,N_15409);
or U18414 (N_18414,N_14048,N_12212);
xnor U18415 (N_18415,N_15569,N_13741);
xor U18416 (N_18416,N_12428,N_14602);
and U18417 (N_18417,N_12860,N_14194);
xor U18418 (N_18418,N_14148,N_13234);
nand U18419 (N_18419,N_15953,N_13659);
and U18420 (N_18420,N_13489,N_13364);
and U18421 (N_18421,N_15660,N_12546);
or U18422 (N_18422,N_14757,N_14841);
nand U18423 (N_18423,N_12713,N_12671);
xnor U18424 (N_18424,N_12610,N_12278);
and U18425 (N_18425,N_14710,N_12145);
or U18426 (N_18426,N_13079,N_12146);
nand U18427 (N_18427,N_12302,N_14908);
xor U18428 (N_18428,N_15342,N_15112);
nand U18429 (N_18429,N_14831,N_14031);
and U18430 (N_18430,N_12656,N_13575);
nor U18431 (N_18431,N_12840,N_14761);
nand U18432 (N_18432,N_13414,N_13280);
or U18433 (N_18433,N_14223,N_15770);
or U18434 (N_18434,N_15291,N_12780);
xnor U18435 (N_18435,N_13653,N_13487);
nand U18436 (N_18436,N_13025,N_15554);
xor U18437 (N_18437,N_14893,N_15891);
or U18438 (N_18438,N_14708,N_12911);
or U18439 (N_18439,N_13086,N_15484);
nand U18440 (N_18440,N_14438,N_13715);
or U18441 (N_18441,N_15948,N_14190);
xnor U18442 (N_18442,N_12811,N_13260);
nand U18443 (N_18443,N_14875,N_15628);
or U18444 (N_18444,N_12845,N_14080);
xnor U18445 (N_18445,N_13606,N_14110);
or U18446 (N_18446,N_13696,N_12694);
and U18447 (N_18447,N_12979,N_14917);
or U18448 (N_18448,N_14232,N_15071);
xnor U18449 (N_18449,N_14818,N_12887);
or U18450 (N_18450,N_15453,N_14150);
nand U18451 (N_18451,N_14005,N_15764);
nor U18452 (N_18452,N_15021,N_12490);
nor U18453 (N_18453,N_14324,N_12070);
and U18454 (N_18454,N_14399,N_13695);
or U18455 (N_18455,N_13695,N_14212);
or U18456 (N_18456,N_12966,N_15230);
xor U18457 (N_18457,N_15968,N_14346);
or U18458 (N_18458,N_14899,N_15581);
nor U18459 (N_18459,N_14395,N_13362);
nand U18460 (N_18460,N_13522,N_13392);
xnor U18461 (N_18461,N_13194,N_13111);
xnor U18462 (N_18462,N_13469,N_12136);
nor U18463 (N_18463,N_12356,N_14969);
or U18464 (N_18464,N_13332,N_13269);
xor U18465 (N_18465,N_15464,N_15543);
nand U18466 (N_18466,N_13637,N_13292);
nand U18467 (N_18467,N_14420,N_14259);
nor U18468 (N_18468,N_15008,N_15767);
or U18469 (N_18469,N_15598,N_14599);
xnor U18470 (N_18470,N_12665,N_14049);
or U18471 (N_18471,N_14356,N_14443);
or U18472 (N_18472,N_15257,N_14899);
xor U18473 (N_18473,N_14363,N_12667);
nand U18474 (N_18474,N_13752,N_13608);
nor U18475 (N_18475,N_12227,N_12122);
nor U18476 (N_18476,N_13599,N_15272);
and U18477 (N_18477,N_14968,N_13818);
and U18478 (N_18478,N_12481,N_12722);
and U18479 (N_18479,N_14569,N_15072);
and U18480 (N_18480,N_14581,N_12473);
nor U18481 (N_18481,N_15812,N_12881);
xnor U18482 (N_18482,N_13786,N_14078);
and U18483 (N_18483,N_13172,N_15889);
nor U18484 (N_18484,N_13547,N_12502);
xnor U18485 (N_18485,N_15056,N_14268);
and U18486 (N_18486,N_14552,N_14478);
nor U18487 (N_18487,N_12253,N_13144);
or U18488 (N_18488,N_12672,N_12190);
and U18489 (N_18489,N_14755,N_15409);
nor U18490 (N_18490,N_14995,N_12238);
nand U18491 (N_18491,N_12325,N_13330);
and U18492 (N_18492,N_12427,N_13877);
nor U18493 (N_18493,N_12773,N_12849);
nand U18494 (N_18494,N_12856,N_12962);
nor U18495 (N_18495,N_12825,N_13952);
xor U18496 (N_18496,N_15532,N_15866);
or U18497 (N_18497,N_15956,N_14770);
xor U18498 (N_18498,N_12022,N_13080);
nor U18499 (N_18499,N_12438,N_13766);
xnor U18500 (N_18500,N_14206,N_15477);
xor U18501 (N_18501,N_15348,N_13521);
xor U18502 (N_18502,N_13893,N_13378);
xnor U18503 (N_18503,N_12703,N_14744);
and U18504 (N_18504,N_13222,N_12912);
and U18505 (N_18505,N_15833,N_14335);
nor U18506 (N_18506,N_12886,N_15712);
nand U18507 (N_18507,N_12987,N_12420);
nor U18508 (N_18508,N_14762,N_15442);
nor U18509 (N_18509,N_15200,N_12085);
xnor U18510 (N_18510,N_15850,N_14569);
nand U18511 (N_18511,N_14275,N_13999);
or U18512 (N_18512,N_12068,N_12374);
or U18513 (N_18513,N_13807,N_14817);
and U18514 (N_18514,N_15923,N_15772);
and U18515 (N_18515,N_13028,N_14887);
xnor U18516 (N_18516,N_13494,N_12460);
xor U18517 (N_18517,N_15592,N_13737);
nand U18518 (N_18518,N_15381,N_14746);
and U18519 (N_18519,N_12723,N_13276);
nand U18520 (N_18520,N_12713,N_15358);
nor U18521 (N_18521,N_13477,N_13452);
nand U18522 (N_18522,N_13120,N_15480);
or U18523 (N_18523,N_13540,N_12317);
or U18524 (N_18524,N_14309,N_15241);
nand U18525 (N_18525,N_12975,N_14803);
nand U18526 (N_18526,N_12599,N_14189);
nor U18527 (N_18527,N_15101,N_12453);
nand U18528 (N_18528,N_12413,N_13172);
nor U18529 (N_18529,N_15057,N_13053);
nand U18530 (N_18530,N_15799,N_14596);
or U18531 (N_18531,N_12883,N_14802);
and U18532 (N_18532,N_14784,N_12076);
xor U18533 (N_18533,N_13158,N_14278);
or U18534 (N_18534,N_14322,N_15879);
nor U18535 (N_18535,N_14749,N_12266);
xnor U18536 (N_18536,N_12655,N_13312);
nor U18537 (N_18537,N_12712,N_14565);
nand U18538 (N_18538,N_15662,N_15375);
xnor U18539 (N_18539,N_14592,N_13519);
nand U18540 (N_18540,N_14968,N_14084);
nand U18541 (N_18541,N_12872,N_12348);
or U18542 (N_18542,N_15238,N_15441);
nor U18543 (N_18543,N_15760,N_13463);
or U18544 (N_18544,N_13564,N_15426);
or U18545 (N_18545,N_13808,N_12936);
xor U18546 (N_18546,N_13661,N_15669);
and U18547 (N_18547,N_12919,N_15899);
or U18548 (N_18548,N_15717,N_12662);
or U18549 (N_18549,N_15482,N_14395);
nor U18550 (N_18550,N_14464,N_12262);
nand U18551 (N_18551,N_14003,N_15826);
or U18552 (N_18552,N_15355,N_12186);
or U18553 (N_18553,N_13120,N_12007);
xor U18554 (N_18554,N_12608,N_15970);
nand U18555 (N_18555,N_14308,N_12633);
xor U18556 (N_18556,N_13714,N_12305);
and U18557 (N_18557,N_14055,N_13640);
and U18558 (N_18558,N_13844,N_15211);
or U18559 (N_18559,N_15795,N_13182);
xnor U18560 (N_18560,N_13044,N_13677);
xor U18561 (N_18561,N_12537,N_14619);
or U18562 (N_18562,N_15604,N_13657);
xor U18563 (N_18563,N_15643,N_12012);
and U18564 (N_18564,N_15765,N_14699);
nand U18565 (N_18565,N_12926,N_13169);
nand U18566 (N_18566,N_15474,N_15693);
nand U18567 (N_18567,N_15082,N_12466);
and U18568 (N_18568,N_15466,N_14816);
or U18569 (N_18569,N_13943,N_12212);
or U18570 (N_18570,N_13176,N_15981);
or U18571 (N_18571,N_12796,N_12432);
nand U18572 (N_18572,N_15740,N_13632);
or U18573 (N_18573,N_12285,N_14654);
nor U18574 (N_18574,N_14598,N_14758);
and U18575 (N_18575,N_13674,N_14248);
or U18576 (N_18576,N_15084,N_14072);
nor U18577 (N_18577,N_12249,N_12969);
nor U18578 (N_18578,N_13023,N_15420);
nor U18579 (N_18579,N_13284,N_12235);
nand U18580 (N_18580,N_12114,N_13837);
and U18581 (N_18581,N_15583,N_14678);
xnor U18582 (N_18582,N_13885,N_13284);
xnor U18583 (N_18583,N_12062,N_14766);
and U18584 (N_18584,N_14196,N_13661);
nand U18585 (N_18585,N_13845,N_13495);
and U18586 (N_18586,N_13920,N_15763);
and U18587 (N_18587,N_13555,N_14437);
nor U18588 (N_18588,N_15355,N_15926);
nand U18589 (N_18589,N_13673,N_14514);
nand U18590 (N_18590,N_13164,N_15236);
nor U18591 (N_18591,N_13701,N_14369);
xnor U18592 (N_18592,N_13439,N_14408);
nand U18593 (N_18593,N_13263,N_15103);
nand U18594 (N_18594,N_15630,N_12849);
xor U18595 (N_18595,N_13209,N_15344);
and U18596 (N_18596,N_12731,N_13074);
nand U18597 (N_18597,N_13309,N_14184);
and U18598 (N_18598,N_12323,N_13562);
xor U18599 (N_18599,N_15478,N_12291);
or U18600 (N_18600,N_15793,N_12047);
and U18601 (N_18601,N_13965,N_13094);
or U18602 (N_18602,N_12645,N_14928);
or U18603 (N_18603,N_12097,N_13037);
nor U18604 (N_18604,N_15197,N_14334);
and U18605 (N_18605,N_14114,N_12929);
and U18606 (N_18606,N_15977,N_14759);
and U18607 (N_18607,N_13589,N_15848);
xnor U18608 (N_18608,N_12161,N_13452);
nand U18609 (N_18609,N_14527,N_13251);
nor U18610 (N_18610,N_13276,N_13632);
nand U18611 (N_18611,N_13969,N_14302);
xnor U18612 (N_18612,N_14634,N_14995);
or U18613 (N_18613,N_15214,N_13688);
xor U18614 (N_18614,N_12782,N_12005);
xnor U18615 (N_18615,N_15393,N_12980);
or U18616 (N_18616,N_15279,N_15737);
nand U18617 (N_18617,N_14285,N_14380);
or U18618 (N_18618,N_15593,N_14221);
or U18619 (N_18619,N_14202,N_13764);
nand U18620 (N_18620,N_14954,N_14609);
and U18621 (N_18621,N_13107,N_15278);
and U18622 (N_18622,N_15593,N_14713);
nor U18623 (N_18623,N_14838,N_13998);
nor U18624 (N_18624,N_12018,N_13270);
and U18625 (N_18625,N_13584,N_15146);
and U18626 (N_18626,N_12126,N_12410);
nand U18627 (N_18627,N_14596,N_13720);
xor U18628 (N_18628,N_14265,N_15543);
nor U18629 (N_18629,N_12972,N_13683);
or U18630 (N_18630,N_14517,N_13926);
or U18631 (N_18631,N_13053,N_15528);
and U18632 (N_18632,N_12060,N_14925);
or U18633 (N_18633,N_12892,N_13950);
nor U18634 (N_18634,N_13804,N_13287);
xor U18635 (N_18635,N_12913,N_13942);
nor U18636 (N_18636,N_15538,N_14275);
or U18637 (N_18637,N_15275,N_15644);
xor U18638 (N_18638,N_12665,N_15007);
nand U18639 (N_18639,N_14421,N_12505);
and U18640 (N_18640,N_15730,N_14338);
nand U18641 (N_18641,N_14108,N_12924);
xor U18642 (N_18642,N_15291,N_13368);
nor U18643 (N_18643,N_15636,N_13275);
nor U18644 (N_18644,N_15928,N_12542);
xnor U18645 (N_18645,N_13052,N_12385);
xor U18646 (N_18646,N_12905,N_14333);
or U18647 (N_18647,N_14656,N_15166);
nor U18648 (N_18648,N_13189,N_15414);
nand U18649 (N_18649,N_14622,N_15666);
and U18650 (N_18650,N_14501,N_14010);
nor U18651 (N_18651,N_12955,N_15060);
or U18652 (N_18652,N_12340,N_12545);
xnor U18653 (N_18653,N_14253,N_14298);
nand U18654 (N_18654,N_13908,N_15748);
or U18655 (N_18655,N_13997,N_15128);
nor U18656 (N_18656,N_13367,N_14961);
nor U18657 (N_18657,N_15404,N_15557);
or U18658 (N_18658,N_14989,N_14074);
nand U18659 (N_18659,N_13830,N_15224);
xor U18660 (N_18660,N_15559,N_14141);
nor U18661 (N_18661,N_12453,N_12612);
or U18662 (N_18662,N_15208,N_14034);
or U18663 (N_18663,N_14844,N_14885);
xnor U18664 (N_18664,N_15825,N_12389);
or U18665 (N_18665,N_14240,N_12983);
xnor U18666 (N_18666,N_12523,N_13600);
or U18667 (N_18667,N_14306,N_13822);
and U18668 (N_18668,N_15364,N_12488);
nor U18669 (N_18669,N_12614,N_15103);
and U18670 (N_18670,N_12351,N_15925);
and U18671 (N_18671,N_13935,N_14371);
nor U18672 (N_18672,N_15442,N_13840);
nor U18673 (N_18673,N_15146,N_13916);
nor U18674 (N_18674,N_12497,N_12356);
or U18675 (N_18675,N_13213,N_14587);
and U18676 (N_18676,N_12998,N_12814);
nor U18677 (N_18677,N_14386,N_14861);
or U18678 (N_18678,N_15001,N_12142);
or U18679 (N_18679,N_13101,N_14295);
or U18680 (N_18680,N_12918,N_15796);
or U18681 (N_18681,N_12082,N_12006);
and U18682 (N_18682,N_13757,N_15334);
and U18683 (N_18683,N_13691,N_13777);
and U18684 (N_18684,N_12437,N_12171);
nand U18685 (N_18685,N_13373,N_12492);
nand U18686 (N_18686,N_12365,N_15640);
xnor U18687 (N_18687,N_14953,N_15154);
or U18688 (N_18688,N_15872,N_12191);
nand U18689 (N_18689,N_12395,N_13261);
or U18690 (N_18690,N_15615,N_12547);
xor U18691 (N_18691,N_14632,N_12241);
nand U18692 (N_18692,N_14830,N_15691);
and U18693 (N_18693,N_15825,N_14147);
xor U18694 (N_18694,N_14499,N_15435);
nor U18695 (N_18695,N_14008,N_12585);
or U18696 (N_18696,N_14457,N_12448);
nand U18697 (N_18697,N_14212,N_13362);
and U18698 (N_18698,N_14361,N_12395);
or U18699 (N_18699,N_15171,N_14636);
xor U18700 (N_18700,N_12649,N_13013);
nand U18701 (N_18701,N_15857,N_12958);
nand U18702 (N_18702,N_12117,N_15986);
or U18703 (N_18703,N_12590,N_12188);
nand U18704 (N_18704,N_12461,N_14960);
or U18705 (N_18705,N_12413,N_13998);
xnor U18706 (N_18706,N_15076,N_12200);
xnor U18707 (N_18707,N_12716,N_12250);
nand U18708 (N_18708,N_14680,N_12923);
xor U18709 (N_18709,N_13142,N_13577);
and U18710 (N_18710,N_15049,N_15382);
nor U18711 (N_18711,N_14336,N_14539);
and U18712 (N_18712,N_14863,N_14105);
nand U18713 (N_18713,N_15960,N_15157);
xor U18714 (N_18714,N_12005,N_12640);
nor U18715 (N_18715,N_14109,N_15694);
nand U18716 (N_18716,N_13220,N_12514);
xnor U18717 (N_18717,N_14821,N_12724);
or U18718 (N_18718,N_12195,N_12935);
nor U18719 (N_18719,N_15427,N_13434);
and U18720 (N_18720,N_14880,N_12483);
nand U18721 (N_18721,N_13478,N_14173);
nand U18722 (N_18722,N_12976,N_12458);
or U18723 (N_18723,N_14248,N_14638);
nand U18724 (N_18724,N_12401,N_13191);
xor U18725 (N_18725,N_15601,N_12845);
nand U18726 (N_18726,N_14987,N_13577);
xnor U18727 (N_18727,N_12995,N_14074);
nor U18728 (N_18728,N_12513,N_12436);
xnor U18729 (N_18729,N_13308,N_13512);
and U18730 (N_18730,N_14088,N_12040);
or U18731 (N_18731,N_13534,N_15471);
and U18732 (N_18732,N_13924,N_13534);
nand U18733 (N_18733,N_14050,N_13852);
xor U18734 (N_18734,N_15404,N_15756);
nor U18735 (N_18735,N_14753,N_13618);
nand U18736 (N_18736,N_15230,N_14360);
or U18737 (N_18737,N_12476,N_14997);
or U18738 (N_18738,N_12377,N_15311);
xnor U18739 (N_18739,N_14161,N_13111);
nand U18740 (N_18740,N_14699,N_13263);
and U18741 (N_18741,N_14503,N_14878);
nand U18742 (N_18742,N_12784,N_14538);
nor U18743 (N_18743,N_15387,N_15094);
and U18744 (N_18744,N_12652,N_15304);
nand U18745 (N_18745,N_12531,N_13632);
or U18746 (N_18746,N_14984,N_13783);
or U18747 (N_18747,N_12830,N_13856);
or U18748 (N_18748,N_14515,N_13352);
xor U18749 (N_18749,N_12340,N_14102);
and U18750 (N_18750,N_14187,N_12852);
and U18751 (N_18751,N_14856,N_14880);
xor U18752 (N_18752,N_12584,N_14963);
or U18753 (N_18753,N_15709,N_15220);
nand U18754 (N_18754,N_13655,N_15015);
nor U18755 (N_18755,N_14745,N_13025);
xnor U18756 (N_18756,N_14930,N_15546);
nor U18757 (N_18757,N_13220,N_12815);
nor U18758 (N_18758,N_14383,N_12230);
or U18759 (N_18759,N_13258,N_12495);
or U18760 (N_18760,N_13253,N_15287);
nand U18761 (N_18761,N_13528,N_12633);
or U18762 (N_18762,N_13517,N_13077);
xnor U18763 (N_18763,N_13457,N_15551);
and U18764 (N_18764,N_14810,N_15532);
nor U18765 (N_18765,N_14624,N_15550);
or U18766 (N_18766,N_12892,N_13229);
xor U18767 (N_18767,N_14712,N_13028);
nand U18768 (N_18768,N_13701,N_15190);
or U18769 (N_18769,N_15380,N_14705);
xor U18770 (N_18770,N_13438,N_14656);
xor U18771 (N_18771,N_13285,N_15511);
and U18772 (N_18772,N_13527,N_12396);
and U18773 (N_18773,N_12419,N_12024);
nor U18774 (N_18774,N_14454,N_12632);
or U18775 (N_18775,N_14783,N_12925);
and U18776 (N_18776,N_12263,N_12842);
xnor U18777 (N_18777,N_15562,N_14216);
nand U18778 (N_18778,N_13536,N_15845);
nand U18779 (N_18779,N_14171,N_12494);
nor U18780 (N_18780,N_12737,N_13165);
xnor U18781 (N_18781,N_13292,N_13514);
nand U18782 (N_18782,N_15920,N_13785);
or U18783 (N_18783,N_14064,N_13618);
nor U18784 (N_18784,N_14320,N_15262);
and U18785 (N_18785,N_15757,N_14446);
or U18786 (N_18786,N_14195,N_13743);
nand U18787 (N_18787,N_14755,N_14616);
nor U18788 (N_18788,N_13727,N_13802);
and U18789 (N_18789,N_14970,N_14370);
or U18790 (N_18790,N_15598,N_15424);
and U18791 (N_18791,N_15892,N_13064);
nor U18792 (N_18792,N_13871,N_14410);
xnor U18793 (N_18793,N_13474,N_13140);
or U18794 (N_18794,N_13272,N_14014);
and U18795 (N_18795,N_15386,N_14601);
nor U18796 (N_18796,N_14026,N_15322);
xor U18797 (N_18797,N_12363,N_15536);
nor U18798 (N_18798,N_14984,N_15698);
nor U18799 (N_18799,N_14507,N_14598);
nand U18800 (N_18800,N_12781,N_14873);
and U18801 (N_18801,N_12116,N_14096);
and U18802 (N_18802,N_12932,N_15031);
xor U18803 (N_18803,N_12093,N_15047);
or U18804 (N_18804,N_14125,N_15274);
nand U18805 (N_18805,N_15213,N_14388);
or U18806 (N_18806,N_15114,N_14373);
and U18807 (N_18807,N_13188,N_13360);
and U18808 (N_18808,N_14796,N_13434);
nand U18809 (N_18809,N_13172,N_15022);
nor U18810 (N_18810,N_12050,N_14752);
and U18811 (N_18811,N_13250,N_13630);
or U18812 (N_18812,N_15588,N_14769);
nor U18813 (N_18813,N_15897,N_14902);
xnor U18814 (N_18814,N_14414,N_14030);
or U18815 (N_18815,N_14629,N_14722);
nand U18816 (N_18816,N_12081,N_14586);
and U18817 (N_18817,N_14593,N_13989);
nand U18818 (N_18818,N_12575,N_14814);
or U18819 (N_18819,N_12021,N_14564);
and U18820 (N_18820,N_15710,N_15464);
or U18821 (N_18821,N_14228,N_15419);
and U18822 (N_18822,N_15625,N_15763);
nor U18823 (N_18823,N_13434,N_14641);
or U18824 (N_18824,N_12334,N_14368);
or U18825 (N_18825,N_15924,N_15785);
or U18826 (N_18826,N_14764,N_12281);
and U18827 (N_18827,N_12767,N_15624);
nand U18828 (N_18828,N_14917,N_12751);
and U18829 (N_18829,N_14580,N_13045);
or U18830 (N_18830,N_15788,N_15987);
and U18831 (N_18831,N_12782,N_12080);
or U18832 (N_18832,N_15935,N_13371);
or U18833 (N_18833,N_15871,N_12774);
and U18834 (N_18834,N_14174,N_15447);
or U18835 (N_18835,N_14520,N_13322);
or U18836 (N_18836,N_15202,N_13225);
nor U18837 (N_18837,N_12600,N_13664);
nor U18838 (N_18838,N_14835,N_12926);
xnor U18839 (N_18839,N_13019,N_13369);
xor U18840 (N_18840,N_13492,N_14006);
or U18841 (N_18841,N_13105,N_15953);
or U18842 (N_18842,N_14230,N_12272);
nor U18843 (N_18843,N_15282,N_14507);
nor U18844 (N_18844,N_12998,N_12536);
nand U18845 (N_18845,N_14857,N_15712);
or U18846 (N_18846,N_14674,N_15783);
nand U18847 (N_18847,N_14951,N_13409);
xor U18848 (N_18848,N_15492,N_14749);
and U18849 (N_18849,N_14439,N_13896);
and U18850 (N_18850,N_14261,N_15055);
or U18851 (N_18851,N_12951,N_15995);
or U18852 (N_18852,N_15106,N_14414);
nand U18853 (N_18853,N_12816,N_15722);
and U18854 (N_18854,N_14507,N_15136);
nor U18855 (N_18855,N_15929,N_15489);
nor U18856 (N_18856,N_15875,N_12873);
or U18857 (N_18857,N_13561,N_13192);
or U18858 (N_18858,N_15606,N_13757);
and U18859 (N_18859,N_15503,N_12607);
and U18860 (N_18860,N_13905,N_14636);
and U18861 (N_18861,N_13700,N_15351);
xor U18862 (N_18862,N_12357,N_13920);
nor U18863 (N_18863,N_12451,N_13755);
nand U18864 (N_18864,N_12930,N_12851);
xor U18865 (N_18865,N_13528,N_15884);
nand U18866 (N_18866,N_12848,N_14728);
and U18867 (N_18867,N_13342,N_15395);
xor U18868 (N_18868,N_15502,N_15956);
nand U18869 (N_18869,N_14128,N_12566);
xor U18870 (N_18870,N_13738,N_15728);
xnor U18871 (N_18871,N_14773,N_14754);
xnor U18872 (N_18872,N_12602,N_12516);
or U18873 (N_18873,N_15740,N_12344);
nand U18874 (N_18874,N_14492,N_12868);
nand U18875 (N_18875,N_12965,N_15861);
nand U18876 (N_18876,N_14301,N_14507);
or U18877 (N_18877,N_14246,N_14681);
xor U18878 (N_18878,N_13019,N_14819);
xnor U18879 (N_18879,N_14667,N_15717);
xnor U18880 (N_18880,N_15107,N_15591);
and U18881 (N_18881,N_15392,N_13377);
nand U18882 (N_18882,N_13809,N_14172);
xor U18883 (N_18883,N_15492,N_12790);
nor U18884 (N_18884,N_14383,N_15657);
and U18885 (N_18885,N_13464,N_12056);
xnor U18886 (N_18886,N_12872,N_13658);
and U18887 (N_18887,N_14014,N_12632);
nor U18888 (N_18888,N_14874,N_14180);
nor U18889 (N_18889,N_14861,N_14757);
or U18890 (N_18890,N_15856,N_15658);
xnor U18891 (N_18891,N_12031,N_13679);
nor U18892 (N_18892,N_13506,N_13633);
nor U18893 (N_18893,N_14609,N_14936);
nand U18894 (N_18894,N_15969,N_12030);
and U18895 (N_18895,N_13801,N_13117);
xnor U18896 (N_18896,N_14984,N_14347);
and U18897 (N_18897,N_12706,N_12118);
and U18898 (N_18898,N_12301,N_14225);
or U18899 (N_18899,N_15902,N_13904);
or U18900 (N_18900,N_12902,N_13574);
nor U18901 (N_18901,N_14338,N_13688);
xor U18902 (N_18902,N_12344,N_15025);
nor U18903 (N_18903,N_12875,N_13492);
nor U18904 (N_18904,N_12693,N_14840);
xor U18905 (N_18905,N_12500,N_15103);
nand U18906 (N_18906,N_14163,N_13631);
nor U18907 (N_18907,N_14395,N_15809);
or U18908 (N_18908,N_14623,N_13001);
nand U18909 (N_18909,N_15924,N_14738);
or U18910 (N_18910,N_15499,N_12138);
nand U18911 (N_18911,N_14291,N_15317);
xnor U18912 (N_18912,N_15639,N_12289);
and U18913 (N_18913,N_14882,N_15084);
xnor U18914 (N_18914,N_14790,N_13597);
and U18915 (N_18915,N_14651,N_12696);
xor U18916 (N_18916,N_14369,N_13885);
nand U18917 (N_18917,N_13382,N_12173);
or U18918 (N_18918,N_15159,N_14308);
xnor U18919 (N_18919,N_15460,N_14807);
and U18920 (N_18920,N_13661,N_13015);
and U18921 (N_18921,N_14858,N_12707);
or U18922 (N_18922,N_13173,N_14223);
xnor U18923 (N_18923,N_13658,N_12227);
nand U18924 (N_18924,N_13796,N_13344);
and U18925 (N_18925,N_15330,N_14273);
nand U18926 (N_18926,N_15732,N_14170);
or U18927 (N_18927,N_13512,N_13707);
xnor U18928 (N_18928,N_12653,N_13978);
or U18929 (N_18929,N_15643,N_13696);
nor U18930 (N_18930,N_15514,N_15521);
and U18931 (N_18931,N_12007,N_13647);
xor U18932 (N_18932,N_15767,N_15333);
xor U18933 (N_18933,N_13101,N_14784);
nand U18934 (N_18934,N_15704,N_14405);
nand U18935 (N_18935,N_15621,N_15127);
nand U18936 (N_18936,N_15587,N_12159);
nand U18937 (N_18937,N_13192,N_15252);
nand U18938 (N_18938,N_15540,N_15903);
or U18939 (N_18939,N_12891,N_13400);
or U18940 (N_18940,N_13593,N_15021);
nor U18941 (N_18941,N_14057,N_15920);
nand U18942 (N_18942,N_12985,N_12547);
nor U18943 (N_18943,N_13691,N_14162);
xor U18944 (N_18944,N_13011,N_13321);
or U18945 (N_18945,N_12975,N_14020);
nor U18946 (N_18946,N_12743,N_14399);
nor U18947 (N_18947,N_13049,N_14352);
nand U18948 (N_18948,N_12148,N_12398);
xor U18949 (N_18949,N_13009,N_13650);
nor U18950 (N_18950,N_14586,N_12411);
and U18951 (N_18951,N_13831,N_15188);
and U18952 (N_18952,N_13434,N_13143);
nand U18953 (N_18953,N_12870,N_15133);
or U18954 (N_18954,N_15185,N_12737);
nand U18955 (N_18955,N_13864,N_14613);
or U18956 (N_18956,N_14869,N_13348);
and U18957 (N_18957,N_13036,N_13196);
xor U18958 (N_18958,N_13888,N_12388);
nand U18959 (N_18959,N_14896,N_15349);
xor U18960 (N_18960,N_13775,N_12447);
or U18961 (N_18961,N_12523,N_13220);
or U18962 (N_18962,N_15305,N_15504);
nor U18963 (N_18963,N_12303,N_15280);
and U18964 (N_18964,N_12157,N_12018);
or U18965 (N_18965,N_14287,N_12486);
xor U18966 (N_18966,N_13069,N_14635);
nand U18967 (N_18967,N_14727,N_13015);
nor U18968 (N_18968,N_13866,N_15552);
and U18969 (N_18969,N_15007,N_13867);
nor U18970 (N_18970,N_15068,N_12558);
and U18971 (N_18971,N_12318,N_14955);
and U18972 (N_18972,N_12361,N_15362);
or U18973 (N_18973,N_15939,N_14962);
and U18974 (N_18974,N_15531,N_14516);
and U18975 (N_18975,N_12256,N_12854);
xor U18976 (N_18976,N_12883,N_14875);
xnor U18977 (N_18977,N_14440,N_12417);
nand U18978 (N_18978,N_13115,N_15688);
and U18979 (N_18979,N_13420,N_15781);
or U18980 (N_18980,N_15766,N_12197);
nand U18981 (N_18981,N_15388,N_12908);
or U18982 (N_18982,N_15133,N_15325);
nor U18983 (N_18983,N_13303,N_15642);
nand U18984 (N_18984,N_15755,N_14800);
nor U18985 (N_18985,N_13180,N_14040);
and U18986 (N_18986,N_13189,N_12360);
or U18987 (N_18987,N_12032,N_13212);
xor U18988 (N_18988,N_15355,N_13432);
nor U18989 (N_18989,N_13966,N_12086);
and U18990 (N_18990,N_12476,N_15412);
xor U18991 (N_18991,N_15331,N_13982);
nand U18992 (N_18992,N_13775,N_12037);
xnor U18993 (N_18993,N_14375,N_13704);
nor U18994 (N_18994,N_14296,N_15335);
or U18995 (N_18995,N_13245,N_13575);
xnor U18996 (N_18996,N_13769,N_13966);
nor U18997 (N_18997,N_12779,N_13900);
nor U18998 (N_18998,N_15263,N_15943);
xor U18999 (N_18999,N_15238,N_15642);
xor U19000 (N_19000,N_13058,N_12011);
or U19001 (N_19001,N_15473,N_14139);
nand U19002 (N_19002,N_15717,N_14856);
xor U19003 (N_19003,N_15631,N_15769);
or U19004 (N_19004,N_12551,N_13899);
nand U19005 (N_19005,N_14226,N_12397);
xor U19006 (N_19006,N_13852,N_13153);
xnor U19007 (N_19007,N_12605,N_14931);
and U19008 (N_19008,N_12081,N_13134);
or U19009 (N_19009,N_13570,N_13829);
xor U19010 (N_19010,N_12561,N_14376);
nor U19011 (N_19011,N_12348,N_15674);
nand U19012 (N_19012,N_13640,N_13485);
xor U19013 (N_19013,N_12729,N_13514);
or U19014 (N_19014,N_14967,N_13133);
nand U19015 (N_19015,N_13261,N_14923);
and U19016 (N_19016,N_15995,N_15286);
xnor U19017 (N_19017,N_12196,N_14271);
or U19018 (N_19018,N_14106,N_15308);
or U19019 (N_19019,N_14517,N_14013);
nor U19020 (N_19020,N_12384,N_12747);
xnor U19021 (N_19021,N_14404,N_14993);
xnor U19022 (N_19022,N_12598,N_14024);
and U19023 (N_19023,N_14196,N_13366);
nor U19024 (N_19024,N_13586,N_13207);
or U19025 (N_19025,N_13096,N_15260);
xor U19026 (N_19026,N_15920,N_13675);
xor U19027 (N_19027,N_14332,N_14540);
nand U19028 (N_19028,N_15216,N_12887);
or U19029 (N_19029,N_12547,N_15226);
and U19030 (N_19030,N_13004,N_14142);
xor U19031 (N_19031,N_15972,N_15284);
nor U19032 (N_19032,N_15274,N_13145);
or U19033 (N_19033,N_15697,N_15658);
nor U19034 (N_19034,N_13612,N_14938);
and U19035 (N_19035,N_13062,N_13204);
and U19036 (N_19036,N_13890,N_13815);
xor U19037 (N_19037,N_14301,N_13541);
xor U19038 (N_19038,N_13219,N_12676);
xor U19039 (N_19039,N_15377,N_15595);
or U19040 (N_19040,N_12224,N_15763);
or U19041 (N_19041,N_13098,N_12754);
nor U19042 (N_19042,N_12534,N_12567);
nor U19043 (N_19043,N_12228,N_15176);
nor U19044 (N_19044,N_14545,N_13468);
or U19045 (N_19045,N_14792,N_13493);
or U19046 (N_19046,N_15623,N_12885);
nand U19047 (N_19047,N_15907,N_15837);
nand U19048 (N_19048,N_14273,N_13193);
xnor U19049 (N_19049,N_13178,N_14083);
or U19050 (N_19050,N_14652,N_14274);
xor U19051 (N_19051,N_13270,N_12529);
and U19052 (N_19052,N_14334,N_12277);
or U19053 (N_19053,N_15169,N_12330);
xnor U19054 (N_19054,N_12222,N_13060);
nand U19055 (N_19055,N_15532,N_14757);
or U19056 (N_19056,N_14489,N_15600);
nand U19057 (N_19057,N_13086,N_12448);
xor U19058 (N_19058,N_13685,N_13690);
or U19059 (N_19059,N_13772,N_14575);
nor U19060 (N_19060,N_14575,N_12270);
and U19061 (N_19061,N_13174,N_13798);
nand U19062 (N_19062,N_14418,N_15175);
or U19063 (N_19063,N_13201,N_14648);
and U19064 (N_19064,N_14896,N_12799);
and U19065 (N_19065,N_13651,N_12679);
or U19066 (N_19066,N_15339,N_15508);
nor U19067 (N_19067,N_12861,N_15168);
or U19068 (N_19068,N_13524,N_14310);
or U19069 (N_19069,N_15954,N_13459);
nand U19070 (N_19070,N_15204,N_12825);
nand U19071 (N_19071,N_13750,N_12914);
or U19072 (N_19072,N_15890,N_12004);
nor U19073 (N_19073,N_15468,N_13261);
nand U19074 (N_19074,N_15865,N_12895);
or U19075 (N_19075,N_13430,N_15984);
and U19076 (N_19076,N_13167,N_14712);
nand U19077 (N_19077,N_12506,N_15862);
and U19078 (N_19078,N_13469,N_12384);
or U19079 (N_19079,N_12431,N_12312);
nor U19080 (N_19080,N_14571,N_15231);
nor U19081 (N_19081,N_13412,N_14786);
nand U19082 (N_19082,N_14291,N_12625);
and U19083 (N_19083,N_14148,N_12831);
xor U19084 (N_19084,N_15790,N_13476);
xor U19085 (N_19085,N_12735,N_13579);
nand U19086 (N_19086,N_15078,N_13485);
or U19087 (N_19087,N_15801,N_15033);
or U19088 (N_19088,N_14508,N_14648);
nor U19089 (N_19089,N_15530,N_12948);
and U19090 (N_19090,N_15110,N_15527);
xor U19091 (N_19091,N_12396,N_15110);
nor U19092 (N_19092,N_15084,N_13187);
or U19093 (N_19093,N_12281,N_13867);
or U19094 (N_19094,N_15095,N_13174);
or U19095 (N_19095,N_13135,N_12875);
xnor U19096 (N_19096,N_15837,N_12887);
xor U19097 (N_19097,N_13561,N_12778);
nor U19098 (N_19098,N_12649,N_14724);
or U19099 (N_19099,N_12309,N_13447);
nand U19100 (N_19100,N_12328,N_13384);
and U19101 (N_19101,N_14600,N_15429);
nor U19102 (N_19102,N_14138,N_15643);
or U19103 (N_19103,N_13349,N_12398);
xor U19104 (N_19104,N_15955,N_13912);
or U19105 (N_19105,N_14773,N_12518);
nand U19106 (N_19106,N_13974,N_12873);
xor U19107 (N_19107,N_14029,N_15639);
and U19108 (N_19108,N_12658,N_14580);
or U19109 (N_19109,N_15952,N_13627);
nor U19110 (N_19110,N_12551,N_12452);
nand U19111 (N_19111,N_13509,N_14700);
and U19112 (N_19112,N_14486,N_15354);
xor U19113 (N_19113,N_12674,N_15531);
xnor U19114 (N_19114,N_13165,N_15533);
xnor U19115 (N_19115,N_12911,N_15331);
xnor U19116 (N_19116,N_13725,N_15593);
nor U19117 (N_19117,N_13877,N_15097);
nand U19118 (N_19118,N_14829,N_12331);
or U19119 (N_19119,N_15182,N_14308);
nand U19120 (N_19120,N_14125,N_14535);
and U19121 (N_19121,N_14366,N_13445);
nor U19122 (N_19122,N_15943,N_13044);
nand U19123 (N_19123,N_12296,N_13853);
nor U19124 (N_19124,N_15140,N_15358);
or U19125 (N_19125,N_13130,N_15150);
or U19126 (N_19126,N_14674,N_14821);
nand U19127 (N_19127,N_15632,N_12868);
and U19128 (N_19128,N_14738,N_15962);
nand U19129 (N_19129,N_15614,N_15366);
xnor U19130 (N_19130,N_15197,N_15130);
or U19131 (N_19131,N_13246,N_14374);
or U19132 (N_19132,N_15511,N_15979);
nor U19133 (N_19133,N_14298,N_13375);
nand U19134 (N_19134,N_12055,N_12338);
and U19135 (N_19135,N_15845,N_15399);
and U19136 (N_19136,N_14008,N_13858);
xor U19137 (N_19137,N_14873,N_15532);
or U19138 (N_19138,N_13820,N_14388);
nor U19139 (N_19139,N_13738,N_13795);
xor U19140 (N_19140,N_14482,N_15624);
or U19141 (N_19141,N_14959,N_12884);
or U19142 (N_19142,N_12447,N_14993);
nor U19143 (N_19143,N_12842,N_14089);
nand U19144 (N_19144,N_15033,N_12909);
xor U19145 (N_19145,N_14658,N_13555);
and U19146 (N_19146,N_15490,N_13964);
and U19147 (N_19147,N_12721,N_12780);
nor U19148 (N_19148,N_13988,N_12687);
or U19149 (N_19149,N_12542,N_14301);
nor U19150 (N_19150,N_13179,N_13226);
or U19151 (N_19151,N_15906,N_13697);
xnor U19152 (N_19152,N_14453,N_14709);
nand U19153 (N_19153,N_14192,N_14757);
xnor U19154 (N_19154,N_15269,N_12993);
nor U19155 (N_19155,N_14124,N_14613);
nand U19156 (N_19156,N_15215,N_15217);
nand U19157 (N_19157,N_13264,N_13996);
nand U19158 (N_19158,N_13694,N_13022);
or U19159 (N_19159,N_15748,N_13615);
or U19160 (N_19160,N_12174,N_14274);
xnor U19161 (N_19161,N_14626,N_13693);
nor U19162 (N_19162,N_13444,N_14748);
xnor U19163 (N_19163,N_14613,N_14777);
or U19164 (N_19164,N_15525,N_15480);
nor U19165 (N_19165,N_15978,N_15431);
nand U19166 (N_19166,N_12468,N_12674);
nor U19167 (N_19167,N_13976,N_12933);
and U19168 (N_19168,N_15162,N_15668);
or U19169 (N_19169,N_12920,N_12802);
and U19170 (N_19170,N_15383,N_14133);
and U19171 (N_19171,N_13715,N_13386);
or U19172 (N_19172,N_15587,N_14832);
nand U19173 (N_19173,N_15790,N_14548);
nor U19174 (N_19174,N_15234,N_15386);
and U19175 (N_19175,N_13039,N_12167);
nor U19176 (N_19176,N_14940,N_13949);
xor U19177 (N_19177,N_14058,N_13489);
or U19178 (N_19178,N_12129,N_12305);
nor U19179 (N_19179,N_12086,N_12272);
xnor U19180 (N_19180,N_13090,N_13937);
xor U19181 (N_19181,N_12514,N_12129);
or U19182 (N_19182,N_13784,N_14992);
nor U19183 (N_19183,N_12584,N_12395);
nand U19184 (N_19184,N_14472,N_15885);
and U19185 (N_19185,N_13420,N_13649);
and U19186 (N_19186,N_15003,N_12529);
nand U19187 (N_19187,N_15686,N_12335);
nor U19188 (N_19188,N_12579,N_13943);
and U19189 (N_19189,N_15987,N_12675);
or U19190 (N_19190,N_12649,N_13826);
nand U19191 (N_19191,N_13022,N_14364);
or U19192 (N_19192,N_14045,N_13651);
and U19193 (N_19193,N_12525,N_15495);
and U19194 (N_19194,N_12329,N_12216);
and U19195 (N_19195,N_14454,N_12174);
nor U19196 (N_19196,N_12059,N_12404);
nor U19197 (N_19197,N_12908,N_13426);
and U19198 (N_19198,N_14536,N_15682);
and U19199 (N_19199,N_15531,N_13030);
nand U19200 (N_19200,N_12974,N_12088);
xnor U19201 (N_19201,N_14503,N_12358);
and U19202 (N_19202,N_12355,N_13844);
xor U19203 (N_19203,N_13491,N_13885);
xnor U19204 (N_19204,N_12246,N_14540);
nor U19205 (N_19205,N_13508,N_15505);
nand U19206 (N_19206,N_12099,N_13537);
and U19207 (N_19207,N_13460,N_13925);
and U19208 (N_19208,N_13184,N_14669);
and U19209 (N_19209,N_14238,N_14897);
or U19210 (N_19210,N_12486,N_14919);
nand U19211 (N_19211,N_12710,N_14306);
xnor U19212 (N_19212,N_15706,N_14258);
and U19213 (N_19213,N_15829,N_14190);
nand U19214 (N_19214,N_12190,N_14806);
nand U19215 (N_19215,N_12016,N_13352);
nand U19216 (N_19216,N_14523,N_13276);
and U19217 (N_19217,N_13139,N_12579);
nand U19218 (N_19218,N_15177,N_13437);
and U19219 (N_19219,N_13274,N_12746);
or U19220 (N_19220,N_12234,N_15799);
and U19221 (N_19221,N_15287,N_15284);
or U19222 (N_19222,N_12320,N_15376);
and U19223 (N_19223,N_13204,N_12435);
nor U19224 (N_19224,N_15054,N_13555);
and U19225 (N_19225,N_12157,N_12961);
nand U19226 (N_19226,N_13182,N_15908);
and U19227 (N_19227,N_15986,N_12035);
nand U19228 (N_19228,N_12333,N_15220);
nor U19229 (N_19229,N_12889,N_14472);
or U19230 (N_19230,N_15508,N_13514);
and U19231 (N_19231,N_13839,N_14635);
xor U19232 (N_19232,N_12143,N_13110);
or U19233 (N_19233,N_15211,N_15366);
and U19234 (N_19234,N_13750,N_14748);
nand U19235 (N_19235,N_14286,N_12382);
and U19236 (N_19236,N_12358,N_14929);
nand U19237 (N_19237,N_13951,N_15388);
nor U19238 (N_19238,N_14755,N_13143);
or U19239 (N_19239,N_12200,N_13834);
and U19240 (N_19240,N_13864,N_13595);
xor U19241 (N_19241,N_14950,N_12517);
xnor U19242 (N_19242,N_13946,N_15469);
nor U19243 (N_19243,N_13110,N_12507);
or U19244 (N_19244,N_13804,N_13388);
nor U19245 (N_19245,N_13195,N_14761);
nor U19246 (N_19246,N_12331,N_12301);
nand U19247 (N_19247,N_13120,N_14059);
xor U19248 (N_19248,N_14442,N_12986);
or U19249 (N_19249,N_12957,N_15963);
and U19250 (N_19250,N_12665,N_15416);
and U19251 (N_19251,N_12193,N_14340);
nor U19252 (N_19252,N_13358,N_13660);
nand U19253 (N_19253,N_13457,N_13569);
nand U19254 (N_19254,N_13584,N_13194);
and U19255 (N_19255,N_14159,N_14681);
nand U19256 (N_19256,N_12550,N_14492);
nand U19257 (N_19257,N_15823,N_13159);
xor U19258 (N_19258,N_14761,N_13982);
xnor U19259 (N_19259,N_13925,N_15673);
or U19260 (N_19260,N_15312,N_13356);
nand U19261 (N_19261,N_14104,N_14068);
or U19262 (N_19262,N_15651,N_13104);
nand U19263 (N_19263,N_12460,N_15115);
and U19264 (N_19264,N_15192,N_14836);
or U19265 (N_19265,N_12829,N_13715);
nand U19266 (N_19266,N_12137,N_15298);
nor U19267 (N_19267,N_14460,N_14052);
and U19268 (N_19268,N_12917,N_13314);
and U19269 (N_19269,N_12783,N_13869);
nor U19270 (N_19270,N_15300,N_13093);
or U19271 (N_19271,N_14286,N_15370);
xor U19272 (N_19272,N_14574,N_13199);
nand U19273 (N_19273,N_14752,N_14475);
nor U19274 (N_19274,N_14977,N_15741);
nand U19275 (N_19275,N_12554,N_12381);
or U19276 (N_19276,N_15822,N_13626);
xnor U19277 (N_19277,N_14037,N_14031);
and U19278 (N_19278,N_12182,N_15483);
and U19279 (N_19279,N_15716,N_14457);
xor U19280 (N_19280,N_15229,N_15665);
nor U19281 (N_19281,N_12665,N_14180);
or U19282 (N_19282,N_15481,N_14909);
and U19283 (N_19283,N_15458,N_15596);
and U19284 (N_19284,N_12011,N_15249);
xor U19285 (N_19285,N_14566,N_14543);
nor U19286 (N_19286,N_13596,N_15239);
xnor U19287 (N_19287,N_14431,N_15522);
nor U19288 (N_19288,N_15311,N_12639);
or U19289 (N_19289,N_14605,N_13036);
nand U19290 (N_19290,N_15758,N_15749);
or U19291 (N_19291,N_14275,N_14560);
nand U19292 (N_19292,N_15116,N_14535);
and U19293 (N_19293,N_12616,N_13377);
xor U19294 (N_19294,N_12482,N_14156);
xor U19295 (N_19295,N_12683,N_13278);
nor U19296 (N_19296,N_12880,N_15853);
nor U19297 (N_19297,N_14031,N_15266);
nor U19298 (N_19298,N_15872,N_14744);
xnor U19299 (N_19299,N_12143,N_14518);
and U19300 (N_19300,N_15305,N_12048);
nor U19301 (N_19301,N_14198,N_14788);
nand U19302 (N_19302,N_14297,N_14505);
xor U19303 (N_19303,N_12461,N_15662);
xnor U19304 (N_19304,N_14135,N_14284);
nor U19305 (N_19305,N_14289,N_15348);
nand U19306 (N_19306,N_12701,N_14549);
or U19307 (N_19307,N_12721,N_13188);
xnor U19308 (N_19308,N_15211,N_13912);
or U19309 (N_19309,N_15610,N_15008);
nand U19310 (N_19310,N_14632,N_13377);
and U19311 (N_19311,N_14201,N_12257);
xor U19312 (N_19312,N_15809,N_14454);
xnor U19313 (N_19313,N_12383,N_15272);
nor U19314 (N_19314,N_15861,N_13552);
xor U19315 (N_19315,N_15475,N_15641);
nand U19316 (N_19316,N_13166,N_14005);
xor U19317 (N_19317,N_13062,N_15566);
nor U19318 (N_19318,N_15446,N_12659);
and U19319 (N_19319,N_14355,N_13990);
nor U19320 (N_19320,N_13938,N_14240);
nand U19321 (N_19321,N_13848,N_14930);
or U19322 (N_19322,N_13978,N_15537);
and U19323 (N_19323,N_14427,N_15283);
or U19324 (N_19324,N_14685,N_14457);
xor U19325 (N_19325,N_14391,N_15994);
nor U19326 (N_19326,N_13519,N_15091);
or U19327 (N_19327,N_12259,N_15319);
xnor U19328 (N_19328,N_14135,N_12031);
and U19329 (N_19329,N_14297,N_15453);
nand U19330 (N_19330,N_15761,N_14895);
nand U19331 (N_19331,N_14477,N_14828);
nor U19332 (N_19332,N_12663,N_13093);
nor U19333 (N_19333,N_13086,N_15436);
nor U19334 (N_19334,N_12276,N_13015);
and U19335 (N_19335,N_12264,N_14182);
and U19336 (N_19336,N_13883,N_13462);
or U19337 (N_19337,N_12913,N_14788);
or U19338 (N_19338,N_14532,N_15088);
or U19339 (N_19339,N_15185,N_13557);
and U19340 (N_19340,N_15456,N_14190);
and U19341 (N_19341,N_12736,N_13852);
and U19342 (N_19342,N_13859,N_14990);
and U19343 (N_19343,N_13689,N_12914);
xnor U19344 (N_19344,N_12357,N_15995);
xor U19345 (N_19345,N_12624,N_14770);
nor U19346 (N_19346,N_12873,N_14160);
xnor U19347 (N_19347,N_15202,N_14864);
nor U19348 (N_19348,N_15838,N_12342);
xnor U19349 (N_19349,N_13075,N_13713);
or U19350 (N_19350,N_13139,N_15448);
or U19351 (N_19351,N_14961,N_13046);
nor U19352 (N_19352,N_14783,N_14306);
xor U19353 (N_19353,N_15587,N_12875);
nand U19354 (N_19354,N_15361,N_14595);
xor U19355 (N_19355,N_14011,N_12624);
or U19356 (N_19356,N_13509,N_14790);
nand U19357 (N_19357,N_14270,N_15251);
and U19358 (N_19358,N_14461,N_12213);
nor U19359 (N_19359,N_13634,N_13253);
and U19360 (N_19360,N_15641,N_13044);
nor U19361 (N_19361,N_15706,N_12236);
and U19362 (N_19362,N_14530,N_13253);
and U19363 (N_19363,N_12975,N_12121);
nand U19364 (N_19364,N_12784,N_14851);
or U19365 (N_19365,N_15968,N_14371);
and U19366 (N_19366,N_12178,N_12349);
nor U19367 (N_19367,N_14054,N_13987);
xnor U19368 (N_19368,N_13053,N_14782);
xnor U19369 (N_19369,N_12899,N_15275);
xnor U19370 (N_19370,N_13318,N_12706);
or U19371 (N_19371,N_14574,N_14394);
or U19372 (N_19372,N_12128,N_13703);
nor U19373 (N_19373,N_14863,N_15762);
xor U19374 (N_19374,N_13418,N_12303);
nand U19375 (N_19375,N_13904,N_14974);
nand U19376 (N_19376,N_13757,N_12947);
and U19377 (N_19377,N_13429,N_14370);
or U19378 (N_19378,N_12098,N_12675);
xnor U19379 (N_19379,N_14150,N_14453);
or U19380 (N_19380,N_15721,N_14707);
nand U19381 (N_19381,N_14971,N_12167);
xnor U19382 (N_19382,N_12423,N_14442);
nor U19383 (N_19383,N_12608,N_12373);
nand U19384 (N_19384,N_12079,N_12129);
and U19385 (N_19385,N_13137,N_13140);
nor U19386 (N_19386,N_12840,N_14671);
and U19387 (N_19387,N_15750,N_13370);
xor U19388 (N_19388,N_14901,N_14196);
and U19389 (N_19389,N_14307,N_13197);
xor U19390 (N_19390,N_15021,N_12553);
or U19391 (N_19391,N_15737,N_15299);
or U19392 (N_19392,N_12058,N_13597);
nand U19393 (N_19393,N_15689,N_15681);
xnor U19394 (N_19394,N_12089,N_12413);
and U19395 (N_19395,N_12935,N_15216);
xnor U19396 (N_19396,N_12351,N_14205);
xor U19397 (N_19397,N_14365,N_12118);
and U19398 (N_19398,N_15340,N_13865);
or U19399 (N_19399,N_14739,N_13035);
nand U19400 (N_19400,N_13456,N_13695);
and U19401 (N_19401,N_13859,N_15604);
xor U19402 (N_19402,N_13686,N_13014);
nor U19403 (N_19403,N_13257,N_14764);
nor U19404 (N_19404,N_14204,N_15038);
or U19405 (N_19405,N_13193,N_14500);
nand U19406 (N_19406,N_15072,N_12125);
nor U19407 (N_19407,N_13667,N_15832);
nor U19408 (N_19408,N_13087,N_14703);
or U19409 (N_19409,N_12673,N_14470);
nor U19410 (N_19410,N_14472,N_12781);
and U19411 (N_19411,N_13485,N_12918);
nor U19412 (N_19412,N_12557,N_14122);
or U19413 (N_19413,N_14098,N_13014);
and U19414 (N_19414,N_14375,N_15389);
nand U19415 (N_19415,N_15943,N_15088);
and U19416 (N_19416,N_13081,N_12979);
or U19417 (N_19417,N_12007,N_15726);
and U19418 (N_19418,N_14750,N_15772);
xnor U19419 (N_19419,N_12290,N_13082);
or U19420 (N_19420,N_15468,N_14846);
and U19421 (N_19421,N_13168,N_14084);
xnor U19422 (N_19422,N_12696,N_14955);
xor U19423 (N_19423,N_12298,N_15365);
nand U19424 (N_19424,N_15451,N_12305);
and U19425 (N_19425,N_13914,N_14330);
and U19426 (N_19426,N_13219,N_13340);
nor U19427 (N_19427,N_13172,N_12357);
xor U19428 (N_19428,N_12412,N_12720);
xnor U19429 (N_19429,N_15145,N_12985);
xor U19430 (N_19430,N_15013,N_13030);
nor U19431 (N_19431,N_12353,N_15210);
nand U19432 (N_19432,N_15909,N_13134);
nand U19433 (N_19433,N_15130,N_15825);
or U19434 (N_19434,N_15986,N_12486);
nor U19435 (N_19435,N_12979,N_12927);
xnor U19436 (N_19436,N_12415,N_12031);
xor U19437 (N_19437,N_14450,N_14524);
or U19438 (N_19438,N_15051,N_15603);
and U19439 (N_19439,N_15227,N_14015);
nand U19440 (N_19440,N_12363,N_15596);
nor U19441 (N_19441,N_13364,N_12592);
or U19442 (N_19442,N_14142,N_15671);
or U19443 (N_19443,N_13455,N_12134);
and U19444 (N_19444,N_13624,N_13546);
nand U19445 (N_19445,N_15837,N_13987);
or U19446 (N_19446,N_14598,N_12701);
and U19447 (N_19447,N_12343,N_15552);
nand U19448 (N_19448,N_15703,N_15138);
xnor U19449 (N_19449,N_13980,N_15479);
xor U19450 (N_19450,N_15174,N_12043);
xnor U19451 (N_19451,N_13781,N_15521);
or U19452 (N_19452,N_14220,N_12261);
nor U19453 (N_19453,N_14885,N_15049);
xnor U19454 (N_19454,N_15416,N_15457);
nand U19455 (N_19455,N_14004,N_12495);
xnor U19456 (N_19456,N_15291,N_12757);
xor U19457 (N_19457,N_14422,N_13570);
and U19458 (N_19458,N_14792,N_13916);
nand U19459 (N_19459,N_12029,N_14491);
xnor U19460 (N_19460,N_13496,N_15039);
or U19461 (N_19461,N_12148,N_14752);
or U19462 (N_19462,N_15758,N_12674);
nand U19463 (N_19463,N_15382,N_13104);
nand U19464 (N_19464,N_15947,N_13838);
nor U19465 (N_19465,N_14350,N_13375);
xor U19466 (N_19466,N_13863,N_15177);
or U19467 (N_19467,N_13795,N_12300);
xor U19468 (N_19468,N_14375,N_15200);
and U19469 (N_19469,N_15046,N_14049);
nand U19470 (N_19470,N_12780,N_14728);
and U19471 (N_19471,N_13910,N_13551);
xor U19472 (N_19472,N_15264,N_14795);
nand U19473 (N_19473,N_14950,N_12721);
xnor U19474 (N_19474,N_13818,N_13314);
xnor U19475 (N_19475,N_14961,N_13904);
xor U19476 (N_19476,N_15117,N_12905);
nand U19477 (N_19477,N_14157,N_14323);
nand U19478 (N_19478,N_12213,N_15025);
nand U19479 (N_19479,N_12375,N_15951);
nand U19480 (N_19480,N_15114,N_14980);
nor U19481 (N_19481,N_15329,N_15870);
xor U19482 (N_19482,N_12720,N_14796);
xnor U19483 (N_19483,N_14474,N_15490);
or U19484 (N_19484,N_15122,N_14059);
nand U19485 (N_19485,N_13465,N_12648);
nand U19486 (N_19486,N_15413,N_13157);
xnor U19487 (N_19487,N_15061,N_12158);
or U19488 (N_19488,N_13824,N_13711);
xnor U19489 (N_19489,N_14713,N_14274);
nand U19490 (N_19490,N_15834,N_12104);
or U19491 (N_19491,N_15404,N_14704);
nand U19492 (N_19492,N_12063,N_13212);
and U19493 (N_19493,N_13962,N_13007);
or U19494 (N_19494,N_12086,N_12762);
xor U19495 (N_19495,N_12411,N_13624);
or U19496 (N_19496,N_12726,N_13146);
or U19497 (N_19497,N_15285,N_15058);
nor U19498 (N_19498,N_13562,N_14201);
nand U19499 (N_19499,N_13068,N_12527);
nand U19500 (N_19500,N_14004,N_13993);
and U19501 (N_19501,N_13472,N_14495);
and U19502 (N_19502,N_14215,N_12254);
nand U19503 (N_19503,N_12510,N_14605);
and U19504 (N_19504,N_15022,N_13497);
or U19505 (N_19505,N_13005,N_13159);
nand U19506 (N_19506,N_13390,N_14839);
nand U19507 (N_19507,N_12130,N_14248);
and U19508 (N_19508,N_12115,N_13582);
nand U19509 (N_19509,N_13016,N_14735);
xor U19510 (N_19510,N_13314,N_15438);
xor U19511 (N_19511,N_13148,N_15412);
nor U19512 (N_19512,N_15204,N_13145);
and U19513 (N_19513,N_13958,N_14184);
nor U19514 (N_19514,N_13450,N_13544);
nand U19515 (N_19515,N_15904,N_15506);
nor U19516 (N_19516,N_13003,N_12451);
and U19517 (N_19517,N_14277,N_12081);
xor U19518 (N_19518,N_13105,N_13888);
nor U19519 (N_19519,N_14365,N_12092);
nand U19520 (N_19520,N_15705,N_15787);
xnor U19521 (N_19521,N_15258,N_12634);
and U19522 (N_19522,N_14110,N_12045);
and U19523 (N_19523,N_15688,N_14069);
or U19524 (N_19524,N_12358,N_15641);
nor U19525 (N_19525,N_15728,N_15490);
nand U19526 (N_19526,N_12608,N_12001);
xnor U19527 (N_19527,N_15605,N_15981);
nor U19528 (N_19528,N_15851,N_13707);
nor U19529 (N_19529,N_15964,N_14198);
or U19530 (N_19530,N_12276,N_12476);
and U19531 (N_19531,N_12042,N_14839);
and U19532 (N_19532,N_14073,N_14923);
or U19533 (N_19533,N_13911,N_14219);
xnor U19534 (N_19534,N_14450,N_15491);
nand U19535 (N_19535,N_14231,N_15233);
and U19536 (N_19536,N_14473,N_13571);
or U19537 (N_19537,N_14667,N_13967);
or U19538 (N_19538,N_15414,N_13707);
xnor U19539 (N_19539,N_12944,N_14758);
nand U19540 (N_19540,N_12353,N_14356);
or U19541 (N_19541,N_12245,N_14578);
or U19542 (N_19542,N_13410,N_14324);
nand U19543 (N_19543,N_12133,N_13785);
xor U19544 (N_19544,N_13418,N_15786);
or U19545 (N_19545,N_13073,N_12152);
xnor U19546 (N_19546,N_12288,N_12875);
nor U19547 (N_19547,N_15717,N_15535);
or U19548 (N_19548,N_12549,N_14384);
xnor U19549 (N_19549,N_12504,N_13400);
nand U19550 (N_19550,N_15636,N_12127);
or U19551 (N_19551,N_14181,N_15151);
nor U19552 (N_19552,N_14605,N_12370);
and U19553 (N_19553,N_13694,N_14395);
nor U19554 (N_19554,N_14305,N_13805);
or U19555 (N_19555,N_13772,N_13055);
xor U19556 (N_19556,N_13635,N_15794);
xnor U19557 (N_19557,N_15422,N_15131);
or U19558 (N_19558,N_13190,N_15617);
xnor U19559 (N_19559,N_12655,N_14644);
or U19560 (N_19560,N_13489,N_13466);
nor U19561 (N_19561,N_13552,N_13676);
nor U19562 (N_19562,N_14131,N_14813);
xor U19563 (N_19563,N_14008,N_12519);
xor U19564 (N_19564,N_15476,N_12093);
or U19565 (N_19565,N_15264,N_14351);
nor U19566 (N_19566,N_15203,N_13192);
or U19567 (N_19567,N_13591,N_12076);
and U19568 (N_19568,N_12986,N_12241);
nor U19569 (N_19569,N_14528,N_15328);
nor U19570 (N_19570,N_13814,N_13790);
nand U19571 (N_19571,N_13547,N_14571);
nor U19572 (N_19572,N_14422,N_15851);
and U19573 (N_19573,N_13655,N_13153);
or U19574 (N_19574,N_14092,N_15638);
nor U19575 (N_19575,N_12299,N_12392);
nand U19576 (N_19576,N_12076,N_12387);
xor U19577 (N_19577,N_14030,N_14659);
and U19578 (N_19578,N_13303,N_12148);
or U19579 (N_19579,N_13313,N_12432);
xnor U19580 (N_19580,N_13241,N_14913);
nor U19581 (N_19581,N_13178,N_14185);
and U19582 (N_19582,N_13334,N_14409);
or U19583 (N_19583,N_15326,N_12127);
and U19584 (N_19584,N_14143,N_14204);
or U19585 (N_19585,N_14624,N_13191);
xnor U19586 (N_19586,N_15236,N_12390);
xor U19587 (N_19587,N_13363,N_14563);
nor U19588 (N_19588,N_12525,N_13927);
nand U19589 (N_19589,N_14368,N_15742);
xnor U19590 (N_19590,N_13507,N_12774);
nand U19591 (N_19591,N_12082,N_15671);
nor U19592 (N_19592,N_14705,N_13494);
xor U19593 (N_19593,N_14178,N_12288);
xor U19594 (N_19594,N_14865,N_12508);
nand U19595 (N_19595,N_12124,N_13921);
nor U19596 (N_19596,N_13136,N_12775);
nand U19597 (N_19597,N_15850,N_13327);
nor U19598 (N_19598,N_12498,N_15225);
xor U19599 (N_19599,N_15491,N_15513);
and U19600 (N_19600,N_13594,N_15196);
and U19601 (N_19601,N_12500,N_15503);
nand U19602 (N_19602,N_12997,N_15265);
and U19603 (N_19603,N_15606,N_14638);
xnor U19604 (N_19604,N_13016,N_14453);
and U19605 (N_19605,N_12311,N_12733);
xor U19606 (N_19606,N_12275,N_13081);
nor U19607 (N_19607,N_15149,N_14063);
and U19608 (N_19608,N_14471,N_12105);
xor U19609 (N_19609,N_15142,N_13625);
nor U19610 (N_19610,N_14650,N_15878);
and U19611 (N_19611,N_14593,N_12191);
or U19612 (N_19612,N_14380,N_12325);
or U19613 (N_19613,N_14458,N_13448);
and U19614 (N_19614,N_14251,N_12862);
nor U19615 (N_19615,N_12582,N_13003);
or U19616 (N_19616,N_15030,N_14877);
nor U19617 (N_19617,N_15155,N_14354);
or U19618 (N_19618,N_12893,N_15881);
xor U19619 (N_19619,N_13465,N_15792);
nand U19620 (N_19620,N_14755,N_13219);
xnor U19621 (N_19621,N_13215,N_12161);
nand U19622 (N_19622,N_14481,N_14971);
xnor U19623 (N_19623,N_13581,N_15883);
nand U19624 (N_19624,N_13516,N_13501);
nor U19625 (N_19625,N_15582,N_12708);
nor U19626 (N_19626,N_12350,N_13619);
nor U19627 (N_19627,N_14703,N_12680);
nand U19628 (N_19628,N_14055,N_14519);
or U19629 (N_19629,N_13182,N_13232);
xor U19630 (N_19630,N_12870,N_14670);
nand U19631 (N_19631,N_12286,N_14070);
or U19632 (N_19632,N_14629,N_12771);
or U19633 (N_19633,N_13779,N_15241);
nand U19634 (N_19634,N_13511,N_15482);
nand U19635 (N_19635,N_12531,N_13847);
and U19636 (N_19636,N_14625,N_12910);
xor U19637 (N_19637,N_15887,N_15826);
or U19638 (N_19638,N_14875,N_15456);
xnor U19639 (N_19639,N_14087,N_15582);
xor U19640 (N_19640,N_13995,N_15755);
xnor U19641 (N_19641,N_13927,N_12484);
xnor U19642 (N_19642,N_12803,N_13114);
xnor U19643 (N_19643,N_14366,N_13967);
nor U19644 (N_19644,N_13938,N_13416);
or U19645 (N_19645,N_12687,N_14071);
xnor U19646 (N_19646,N_13580,N_12736);
nand U19647 (N_19647,N_12034,N_13736);
or U19648 (N_19648,N_13134,N_14774);
or U19649 (N_19649,N_15287,N_12963);
xor U19650 (N_19650,N_13646,N_12496);
xnor U19651 (N_19651,N_15888,N_12006);
xor U19652 (N_19652,N_12157,N_14803);
nor U19653 (N_19653,N_12042,N_15756);
or U19654 (N_19654,N_14016,N_14312);
xor U19655 (N_19655,N_15244,N_13367);
xor U19656 (N_19656,N_13628,N_12161);
or U19657 (N_19657,N_12057,N_14381);
xor U19658 (N_19658,N_13505,N_15431);
or U19659 (N_19659,N_12236,N_13908);
and U19660 (N_19660,N_12832,N_13051);
nor U19661 (N_19661,N_12126,N_12030);
xnor U19662 (N_19662,N_13832,N_15715);
or U19663 (N_19663,N_12266,N_15635);
xor U19664 (N_19664,N_12778,N_13664);
nand U19665 (N_19665,N_12131,N_14278);
nand U19666 (N_19666,N_15907,N_13571);
or U19667 (N_19667,N_13049,N_13330);
nand U19668 (N_19668,N_14604,N_13928);
or U19669 (N_19669,N_15445,N_15476);
xor U19670 (N_19670,N_12982,N_13529);
or U19671 (N_19671,N_12021,N_12816);
nor U19672 (N_19672,N_15827,N_15028);
or U19673 (N_19673,N_12312,N_12971);
xor U19674 (N_19674,N_12119,N_13595);
nor U19675 (N_19675,N_12552,N_15783);
nor U19676 (N_19676,N_15119,N_15573);
xor U19677 (N_19677,N_15157,N_13907);
xor U19678 (N_19678,N_14929,N_14549);
xnor U19679 (N_19679,N_12572,N_15679);
nand U19680 (N_19680,N_14560,N_15335);
xnor U19681 (N_19681,N_13333,N_15511);
nor U19682 (N_19682,N_12142,N_15730);
or U19683 (N_19683,N_13864,N_12323);
and U19684 (N_19684,N_15088,N_15129);
nor U19685 (N_19685,N_12337,N_15694);
or U19686 (N_19686,N_15417,N_13319);
nand U19687 (N_19687,N_13545,N_14906);
nand U19688 (N_19688,N_15575,N_13533);
nor U19689 (N_19689,N_14730,N_13547);
or U19690 (N_19690,N_12907,N_13224);
or U19691 (N_19691,N_13257,N_14845);
or U19692 (N_19692,N_15387,N_14523);
or U19693 (N_19693,N_14267,N_15549);
nand U19694 (N_19694,N_14578,N_13488);
nor U19695 (N_19695,N_13398,N_14763);
and U19696 (N_19696,N_12367,N_12290);
xnor U19697 (N_19697,N_12440,N_12152);
nand U19698 (N_19698,N_13516,N_12161);
nor U19699 (N_19699,N_13790,N_13281);
nor U19700 (N_19700,N_15345,N_14028);
nor U19701 (N_19701,N_12910,N_14015);
xor U19702 (N_19702,N_14197,N_13894);
nand U19703 (N_19703,N_15373,N_15999);
or U19704 (N_19704,N_15110,N_12743);
and U19705 (N_19705,N_12324,N_15113);
or U19706 (N_19706,N_12248,N_12699);
or U19707 (N_19707,N_15292,N_14346);
xnor U19708 (N_19708,N_13451,N_12951);
xor U19709 (N_19709,N_14859,N_13013);
and U19710 (N_19710,N_15220,N_15799);
xor U19711 (N_19711,N_12884,N_13411);
xnor U19712 (N_19712,N_15313,N_12260);
nand U19713 (N_19713,N_14229,N_13192);
xor U19714 (N_19714,N_12877,N_14462);
nand U19715 (N_19715,N_15185,N_14373);
nand U19716 (N_19716,N_15049,N_14926);
nand U19717 (N_19717,N_13525,N_12839);
nor U19718 (N_19718,N_13287,N_12815);
and U19719 (N_19719,N_14765,N_15341);
nor U19720 (N_19720,N_12270,N_14821);
and U19721 (N_19721,N_15912,N_15970);
and U19722 (N_19722,N_15045,N_15457);
xor U19723 (N_19723,N_13662,N_14936);
and U19724 (N_19724,N_14187,N_12927);
nor U19725 (N_19725,N_15814,N_14648);
nor U19726 (N_19726,N_12229,N_13010);
nand U19727 (N_19727,N_13354,N_15278);
xnor U19728 (N_19728,N_12023,N_13189);
nand U19729 (N_19729,N_14944,N_12320);
nor U19730 (N_19730,N_15704,N_14554);
nor U19731 (N_19731,N_14079,N_13480);
and U19732 (N_19732,N_13790,N_14859);
or U19733 (N_19733,N_14148,N_13168);
or U19734 (N_19734,N_13430,N_13384);
or U19735 (N_19735,N_13752,N_15546);
nor U19736 (N_19736,N_14517,N_14856);
nand U19737 (N_19737,N_15374,N_14406);
nor U19738 (N_19738,N_12848,N_13456);
nand U19739 (N_19739,N_15781,N_13986);
and U19740 (N_19740,N_14734,N_15895);
nand U19741 (N_19741,N_12043,N_15140);
xor U19742 (N_19742,N_15963,N_15974);
nand U19743 (N_19743,N_13303,N_14734);
nand U19744 (N_19744,N_12067,N_15736);
xnor U19745 (N_19745,N_14405,N_12380);
xnor U19746 (N_19746,N_13456,N_12081);
nand U19747 (N_19747,N_12598,N_15992);
nor U19748 (N_19748,N_12029,N_13748);
xnor U19749 (N_19749,N_13167,N_14731);
nand U19750 (N_19750,N_14070,N_12449);
xor U19751 (N_19751,N_15053,N_14479);
nor U19752 (N_19752,N_14717,N_13751);
and U19753 (N_19753,N_15600,N_14883);
xnor U19754 (N_19754,N_12052,N_14866);
or U19755 (N_19755,N_13025,N_12240);
nor U19756 (N_19756,N_12737,N_13802);
or U19757 (N_19757,N_13696,N_15649);
or U19758 (N_19758,N_13014,N_13911);
or U19759 (N_19759,N_15222,N_14939);
and U19760 (N_19760,N_13255,N_13928);
or U19761 (N_19761,N_13079,N_15550);
xor U19762 (N_19762,N_13402,N_13951);
and U19763 (N_19763,N_15032,N_15290);
xor U19764 (N_19764,N_14765,N_14213);
nand U19765 (N_19765,N_12293,N_12467);
nor U19766 (N_19766,N_13904,N_12139);
nor U19767 (N_19767,N_14358,N_14918);
or U19768 (N_19768,N_13926,N_14766);
nor U19769 (N_19769,N_14994,N_15594);
and U19770 (N_19770,N_12920,N_15260);
or U19771 (N_19771,N_15572,N_15119);
and U19772 (N_19772,N_14915,N_12172);
nor U19773 (N_19773,N_14600,N_13741);
nor U19774 (N_19774,N_13570,N_13254);
xor U19775 (N_19775,N_14831,N_12467);
nand U19776 (N_19776,N_14378,N_14165);
xor U19777 (N_19777,N_12796,N_13381);
xor U19778 (N_19778,N_14774,N_15855);
or U19779 (N_19779,N_14008,N_12245);
and U19780 (N_19780,N_12851,N_14764);
nand U19781 (N_19781,N_14059,N_14040);
xor U19782 (N_19782,N_14242,N_14362);
and U19783 (N_19783,N_14618,N_12573);
xor U19784 (N_19784,N_12719,N_12465);
and U19785 (N_19785,N_14718,N_13932);
and U19786 (N_19786,N_15383,N_14299);
nand U19787 (N_19787,N_12571,N_13130);
nand U19788 (N_19788,N_13886,N_13366);
or U19789 (N_19789,N_14355,N_13620);
xor U19790 (N_19790,N_13548,N_14218);
or U19791 (N_19791,N_12599,N_15737);
nand U19792 (N_19792,N_14765,N_14907);
nor U19793 (N_19793,N_12104,N_13536);
xor U19794 (N_19794,N_13720,N_12959);
nor U19795 (N_19795,N_15323,N_15745);
or U19796 (N_19796,N_12413,N_12053);
nor U19797 (N_19797,N_12911,N_14824);
xor U19798 (N_19798,N_15387,N_13903);
and U19799 (N_19799,N_12566,N_14048);
and U19800 (N_19800,N_15818,N_12897);
or U19801 (N_19801,N_15784,N_15529);
nand U19802 (N_19802,N_14235,N_13192);
and U19803 (N_19803,N_14141,N_12194);
nand U19804 (N_19804,N_12234,N_14957);
nor U19805 (N_19805,N_12503,N_13146);
nand U19806 (N_19806,N_14886,N_13568);
nor U19807 (N_19807,N_12429,N_13385);
and U19808 (N_19808,N_13992,N_13795);
xnor U19809 (N_19809,N_15582,N_15122);
nor U19810 (N_19810,N_14892,N_15317);
or U19811 (N_19811,N_14969,N_13206);
nand U19812 (N_19812,N_14926,N_14017);
or U19813 (N_19813,N_12913,N_12723);
nand U19814 (N_19814,N_15254,N_12941);
or U19815 (N_19815,N_14659,N_15850);
or U19816 (N_19816,N_13445,N_13151);
or U19817 (N_19817,N_12330,N_12778);
xor U19818 (N_19818,N_14457,N_12543);
xor U19819 (N_19819,N_12582,N_13893);
or U19820 (N_19820,N_14808,N_14497);
nand U19821 (N_19821,N_14861,N_13174);
or U19822 (N_19822,N_13394,N_15929);
nand U19823 (N_19823,N_13156,N_15399);
xnor U19824 (N_19824,N_15496,N_14011);
xor U19825 (N_19825,N_14823,N_13689);
nor U19826 (N_19826,N_13483,N_15663);
nand U19827 (N_19827,N_13819,N_15965);
xnor U19828 (N_19828,N_12261,N_15775);
and U19829 (N_19829,N_12590,N_13231);
nor U19830 (N_19830,N_13051,N_15672);
nor U19831 (N_19831,N_12604,N_12037);
nor U19832 (N_19832,N_12677,N_12089);
nor U19833 (N_19833,N_15082,N_12164);
and U19834 (N_19834,N_15589,N_14004);
nand U19835 (N_19835,N_13531,N_14669);
or U19836 (N_19836,N_14230,N_13642);
nor U19837 (N_19837,N_15074,N_14538);
nor U19838 (N_19838,N_14308,N_14865);
nand U19839 (N_19839,N_12253,N_13781);
xnor U19840 (N_19840,N_13792,N_15400);
and U19841 (N_19841,N_13389,N_14632);
or U19842 (N_19842,N_12137,N_12412);
or U19843 (N_19843,N_15719,N_14994);
xor U19844 (N_19844,N_12738,N_15738);
nor U19845 (N_19845,N_14525,N_15391);
nand U19846 (N_19846,N_15204,N_14121);
or U19847 (N_19847,N_15926,N_14773);
and U19848 (N_19848,N_14549,N_12227);
and U19849 (N_19849,N_12060,N_15850);
nor U19850 (N_19850,N_12738,N_14306);
nor U19851 (N_19851,N_13669,N_14272);
nor U19852 (N_19852,N_13340,N_15605);
nand U19853 (N_19853,N_13778,N_12227);
nand U19854 (N_19854,N_12365,N_14289);
xor U19855 (N_19855,N_15785,N_15307);
and U19856 (N_19856,N_14748,N_13587);
or U19857 (N_19857,N_14549,N_14478);
xor U19858 (N_19858,N_14383,N_13294);
nor U19859 (N_19859,N_15178,N_12359);
and U19860 (N_19860,N_15066,N_14410);
xor U19861 (N_19861,N_13408,N_13540);
nand U19862 (N_19862,N_13540,N_13598);
nor U19863 (N_19863,N_12151,N_12888);
or U19864 (N_19864,N_13181,N_13646);
nor U19865 (N_19865,N_15790,N_13089);
nor U19866 (N_19866,N_12394,N_12078);
or U19867 (N_19867,N_12530,N_14018);
nor U19868 (N_19868,N_13090,N_15660);
xor U19869 (N_19869,N_15004,N_13816);
nand U19870 (N_19870,N_15570,N_13026);
nand U19871 (N_19871,N_14428,N_12348);
nand U19872 (N_19872,N_15283,N_15035);
nand U19873 (N_19873,N_12096,N_13644);
nor U19874 (N_19874,N_12529,N_14916);
nor U19875 (N_19875,N_14536,N_15330);
xor U19876 (N_19876,N_14007,N_12771);
xor U19877 (N_19877,N_14244,N_13069);
or U19878 (N_19878,N_14759,N_13022);
nand U19879 (N_19879,N_12522,N_15696);
nor U19880 (N_19880,N_12559,N_12226);
nand U19881 (N_19881,N_14494,N_14109);
nand U19882 (N_19882,N_15431,N_12962);
nand U19883 (N_19883,N_13436,N_14627);
nand U19884 (N_19884,N_12056,N_13163);
xnor U19885 (N_19885,N_14499,N_14111);
nand U19886 (N_19886,N_13742,N_15958);
and U19887 (N_19887,N_13172,N_14174);
nor U19888 (N_19888,N_15696,N_14023);
nor U19889 (N_19889,N_15024,N_12326);
nor U19890 (N_19890,N_13208,N_15948);
and U19891 (N_19891,N_15877,N_13714);
xor U19892 (N_19892,N_15812,N_14718);
or U19893 (N_19893,N_12322,N_15271);
or U19894 (N_19894,N_13832,N_13995);
and U19895 (N_19895,N_13223,N_13690);
and U19896 (N_19896,N_13594,N_14390);
nor U19897 (N_19897,N_13875,N_15975);
nand U19898 (N_19898,N_15114,N_13935);
or U19899 (N_19899,N_13914,N_15502);
xor U19900 (N_19900,N_13666,N_15310);
and U19901 (N_19901,N_13325,N_15728);
nor U19902 (N_19902,N_14332,N_14065);
and U19903 (N_19903,N_13003,N_15387);
nor U19904 (N_19904,N_13990,N_14395);
nor U19905 (N_19905,N_14463,N_12808);
nor U19906 (N_19906,N_14856,N_13044);
nor U19907 (N_19907,N_12621,N_12078);
and U19908 (N_19908,N_13919,N_15609);
nor U19909 (N_19909,N_12196,N_13239);
nand U19910 (N_19910,N_13138,N_12041);
xnor U19911 (N_19911,N_15216,N_13681);
nor U19912 (N_19912,N_13682,N_14627);
and U19913 (N_19913,N_14785,N_14416);
and U19914 (N_19914,N_15226,N_12263);
xnor U19915 (N_19915,N_14327,N_14188);
nor U19916 (N_19916,N_12417,N_12604);
nor U19917 (N_19917,N_14654,N_13694);
nor U19918 (N_19918,N_13152,N_15366);
xor U19919 (N_19919,N_15483,N_15336);
xor U19920 (N_19920,N_13059,N_14689);
or U19921 (N_19921,N_13270,N_13055);
and U19922 (N_19922,N_12004,N_13620);
nor U19923 (N_19923,N_15927,N_14511);
or U19924 (N_19924,N_12826,N_13563);
xor U19925 (N_19925,N_15084,N_14884);
xnor U19926 (N_19926,N_14671,N_12449);
and U19927 (N_19927,N_12627,N_13142);
nand U19928 (N_19928,N_15644,N_13659);
nand U19929 (N_19929,N_12114,N_12874);
xnor U19930 (N_19930,N_12125,N_14008);
or U19931 (N_19931,N_14873,N_13611);
nor U19932 (N_19932,N_15097,N_14165);
or U19933 (N_19933,N_14009,N_15626);
nor U19934 (N_19934,N_13016,N_13696);
and U19935 (N_19935,N_15783,N_13212);
and U19936 (N_19936,N_14168,N_15281);
xnor U19937 (N_19937,N_12707,N_12126);
and U19938 (N_19938,N_14749,N_15891);
xor U19939 (N_19939,N_15636,N_15237);
nand U19940 (N_19940,N_12581,N_13924);
nand U19941 (N_19941,N_15112,N_13872);
xor U19942 (N_19942,N_15341,N_12171);
or U19943 (N_19943,N_13891,N_13551);
nand U19944 (N_19944,N_14747,N_14929);
nand U19945 (N_19945,N_15668,N_12641);
and U19946 (N_19946,N_13146,N_15287);
nand U19947 (N_19947,N_14189,N_13012);
nand U19948 (N_19948,N_13522,N_14304);
nand U19949 (N_19949,N_15627,N_14144);
nand U19950 (N_19950,N_13025,N_14952);
nand U19951 (N_19951,N_15867,N_15207);
and U19952 (N_19952,N_14908,N_12453);
nand U19953 (N_19953,N_15069,N_15750);
nand U19954 (N_19954,N_12357,N_14166);
xor U19955 (N_19955,N_12167,N_15598);
xnor U19956 (N_19956,N_12551,N_13720);
or U19957 (N_19957,N_13669,N_14496);
nand U19958 (N_19958,N_15288,N_14406);
xor U19959 (N_19959,N_15435,N_15309);
and U19960 (N_19960,N_14869,N_15895);
xnor U19961 (N_19961,N_14638,N_13432);
and U19962 (N_19962,N_15385,N_13443);
xnor U19963 (N_19963,N_13498,N_14978);
nor U19964 (N_19964,N_12883,N_15590);
nor U19965 (N_19965,N_15328,N_15344);
nand U19966 (N_19966,N_12734,N_14425);
or U19967 (N_19967,N_15024,N_14386);
or U19968 (N_19968,N_15184,N_15442);
and U19969 (N_19969,N_12362,N_15781);
or U19970 (N_19970,N_14329,N_13509);
xor U19971 (N_19971,N_13860,N_14041);
xnor U19972 (N_19972,N_15646,N_12796);
nand U19973 (N_19973,N_12532,N_13161);
and U19974 (N_19974,N_15143,N_13319);
and U19975 (N_19975,N_15194,N_14812);
and U19976 (N_19976,N_14149,N_14399);
and U19977 (N_19977,N_12100,N_12547);
xor U19978 (N_19978,N_14485,N_13146);
and U19979 (N_19979,N_12248,N_15959);
and U19980 (N_19980,N_12501,N_13409);
xnor U19981 (N_19981,N_13574,N_12704);
xnor U19982 (N_19982,N_12347,N_12070);
or U19983 (N_19983,N_15705,N_15347);
xor U19984 (N_19984,N_13745,N_12815);
and U19985 (N_19985,N_15255,N_13596);
nand U19986 (N_19986,N_12698,N_13709);
or U19987 (N_19987,N_15537,N_13758);
nor U19988 (N_19988,N_15758,N_14915);
and U19989 (N_19989,N_14189,N_15010);
and U19990 (N_19990,N_15888,N_12283);
nor U19991 (N_19991,N_13444,N_13155);
xor U19992 (N_19992,N_15823,N_12904);
xnor U19993 (N_19993,N_13180,N_12377);
or U19994 (N_19994,N_15075,N_12032);
or U19995 (N_19995,N_12568,N_13586);
or U19996 (N_19996,N_15128,N_14753);
or U19997 (N_19997,N_15557,N_13459);
nand U19998 (N_19998,N_15497,N_15612);
and U19999 (N_19999,N_15093,N_15451);
xor UO_0 (O_0,N_16522,N_17210);
nor UO_1 (O_1,N_17997,N_16863);
nand UO_2 (O_2,N_16166,N_16798);
nand UO_3 (O_3,N_17299,N_18348);
xor UO_4 (O_4,N_19005,N_18038);
nand UO_5 (O_5,N_19469,N_18634);
or UO_6 (O_6,N_16406,N_18980);
nand UO_7 (O_7,N_18702,N_19416);
nand UO_8 (O_8,N_16799,N_18711);
nand UO_9 (O_9,N_17659,N_18575);
or UO_10 (O_10,N_16768,N_16700);
xnor UO_11 (O_11,N_18805,N_16088);
or UO_12 (O_12,N_17360,N_17294);
nor UO_13 (O_13,N_19243,N_18190);
or UO_14 (O_14,N_19531,N_17045);
and UO_15 (O_15,N_18914,N_17792);
nand UO_16 (O_16,N_17197,N_16380);
xor UO_17 (O_17,N_18731,N_17035);
or UO_18 (O_18,N_19484,N_18395);
or UO_19 (O_19,N_18464,N_17160);
and UO_20 (O_20,N_16311,N_19767);
xnor UO_21 (O_21,N_18768,N_18096);
xnor UO_22 (O_22,N_18376,N_18859);
and UO_23 (O_23,N_17368,N_19714);
and UO_24 (O_24,N_17874,N_17136);
and UO_25 (O_25,N_17679,N_19613);
xnor UO_26 (O_26,N_19411,N_19683);
nor UO_27 (O_27,N_18403,N_19997);
nor UO_28 (O_28,N_16655,N_16355);
and UO_29 (O_29,N_16167,N_18443);
nand UO_30 (O_30,N_19021,N_18669);
and UO_31 (O_31,N_16714,N_18465);
and UO_32 (O_32,N_18362,N_18215);
or UO_33 (O_33,N_17575,N_16640);
or UO_34 (O_34,N_19582,N_18142);
nor UO_35 (O_35,N_16667,N_18367);
or UO_36 (O_36,N_19522,N_16690);
and UO_37 (O_37,N_16297,N_18624);
nand UO_38 (O_38,N_17004,N_16412);
nand UO_39 (O_39,N_19998,N_16010);
nor UO_40 (O_40,N_16984,N_17795);
nand UO_41 (O_41,N_16260,N_16299);
and UO_42 (O_42,N_16516,N_17156);
or UO_43 (O_43,N_18984,N_16344);
or UO_44 (O_44,N_17242,N_19149);
nand UO_45 (O_45,N_19177,N_18268);
nor UO_46 (O_46,N_17821,N_18637);
nor UO_47 (O_47,N_16615,N_16679);
or UO_48 (O_48,N_19832,N_19989);
xor UO_49 (O_49,N_19318,N_19829);
and UO_50 (O_50,N_19758,N_16880);
xor UO_51 (O_51,N_18246,N_17396);
xor UO_52 (O_52,N_16231,N_17304);
xor UO_53 (O_53,N_18595,N_16122);
xor UO_54 (O_54,N_17765,N_16481);
and UO_55 (O_55,N_17616,N_16764);
or UO_56 (O_56,N_16000,N_19385);
nor UO_57 (O_57,N_18265,N_19082);
and UO_58 (O_58,N_18930,N_18204);
and UO_59 (O_59,N_18791,N_19399);
or UO_60 (O_60,N_16830,N_17651);
or UO_61 (O_61,N_19198,N_16549);
xor UO_62 (O_62,N_18423,N_19509);
or UO_63 (O_63,N_18559,N_17001);
xor UO_64 (O_64,N_17929,N_16317);
xor UO_65 (O_65,N_16857,N_18703);
or UO_66 (O_66,N_17329,N_18679);
or UO_67 (O_67,N_16797,N_16011);
nor UO_68 (O_68,N_19612,N_16755);
xor UO_69 (O_69,N_17643,N_16420);
xor UO_70 (O_70,N_17948,N_17243);
and UO_71 (O_71,N_17164,N_16821);
and UO_72 (O_72,N_16532,N_19270);
and UO_73 (O_73,N_18767,N_17232);
nand UO_74 (O_74,N_19206,N_18554);
and UO_75 (O_75,N_19859,N_19419);
and UO_76 (O_76,N_19757,N_18912);
nand UO_77 (O_77,N_17280,N_17859);
or UO_78 (O_78,N_19902,N_17278);
xnor UO_79 (O_79,N_17646,N_17829);
nand UO_80 (O_80,N_18809,N_18946);
nand UO_81 (O_81,N_18460,N_17302);
nand UO_82 (O_82,N_17502,N_19554);
nor UO_83 (O_83,N_16001,N_18401);
and UO_84 (O_84,N_16988,N_16177);
nor UO_85 (O_85,N_18184,N_16064);
and UO_86 (O_86,N_16841,N_18343);
or UO_87 (O_87,N_16007,N_17257);
or UO_88 (O_88,N_18999,N_18089);
nor UO_89 (O_89,N_16720,N_16120);
nor UO_90 (O_90,N_18968,N_18596);
nand UO_91 (O_91,N_19065,N_18514);
and UO_92 (O_92,N_19527,N_17328);
and UO_93 (O_93,N_18099,N_17816);
xor UO_94 (O_94,N_17837,N_18932);
and UO_95 (O_95,N_19638,N_17872);
xnor UO_96 (O_96,N_19211,N_16588);
or UO_97 (O_97,N_17227,N_18032);
xor UO_98 (O_98,N_18762,N_16660);
nor UO_99 (O_99,N_17135,N_16336);
nand UO_100 (O_100,N_16652,N_17336);
nor UO_101 (O_101,N_19293,N_19749);
xnor UO_102 (O_102,N_18926,N_19954);
and UO_103 (O_103,N_19508,N_17363);
or UO_104 (O_104,N_17926,N_19456);
nand UO_105 (O_105,N_17256,N_18827);
nor UO_106 (O_106,N_18441,N_18123);
xnor UO_107 (O_107,N_16195,N_17132);
nand UO_108 (O_108,N_16215,N_18847);
xnor UO_109 (O_109,N_16550,N_18192);
xnor UO_110 (O_110,N_19498,N_19855);
and UO_111 (O_111,N_19686,N_18951);
and UO_112 (O_112,N_16298,N_18477);
or UO_113 (O_113,N_16974,N_19425);
nor UO_114 (O_114,N_19312,N_18720);
nor UO_115 (O_115,N_19471,N_19112);
nand UO_116 (O_116,N_18272,N_16090);
nand UO_117 (O_117,N_18836,N_19172);
and UO_118 (O_118,N_19279,N_19427);
nor UO_119 (O_119,N_18838,N_19487);
nand UO_120 (O_120,N_18752,N_16952);
nor UO_121 (O_121,N_19217,N_18700);
and UO_122 (O_122,N_19486,N_17901);
nor UO_123 (O_123,N_16711,N_16484);
nand UO_124 (O_124,N_18977,N_16753);
or UO_125 (O_125,N_18681,N_18668);
nor UO_126 (O_126,N_18356,N_17216);
xor UO_127 (O_127,N_18100,N_16480);
nor UO_128 (O_128,N_18137,N_16659);
xor UO_129 (O_129,N_17514,N_16409);
or UO_130 (O_130,N_17885,N_18843);
xnor UO_131 (O_131,N_18738,N_16770);
xor UO_132 (O_132,N_17196,N_17784);
or UO_133 (O_133,N_18378,N_19822);
or UO_134 (O_134,N_19164,N_18739);
nor UO_135 (O_135,N_18128,N_18852);
nand UO_136 (O_136,N_19039,N_19587);
and UO_137 (O_137,N_17460,N_18650);
nor UO_138 (O_138,N_19881,N_16047);
and UO_139 (O_139,N_18025,N_16892);
nand UO_140 (O_140,N_18018,N_18665);
or UO_141 (O_141,N_19374,N_18026);
nand UO_142 (O_142,N_19864,N_18744);
xor UO_143 (O_143,N_17780,N_17137);
nor UO_144 (O_144,N_18664,N_18566);
or UO_145 (O_145,N_17843,N_16566);
or UO_146 (O_146,N_16022,N_18396);
xor UO_147 (O_147,N_16489,N_19212);
nand UO_148 (O_148,N_17042,N_18715);
nor UO_149 (O_149,N_19200,N_17595);
xnor UO_150 (O_150,N_17127,N_16440);
and UO_151 (O_151,N_16191,N_17857);
or UO_152 (O_152,N_18214,N_18522);
xor UO_153 (O_153,N_19185,N_17725);
or UO_154 (O_154,N_17211,N_19047);
nand UO_155 (O_155,N_19146,N_17582);
nor UO_156 (O_156,N_16668,N_18411);
nor UO_157 (O_157,N_18437,N_17676);
or UO_158 (O_158,N_19052,N_16779);
and UO_159 (O_159,N_16185,N_19151);
xnor UO_160 (O_160,N_16091,N_18986);
or UO_161 (O_161,N_17672,N_18918);
or UO_162 (O_162,N_17204,N_16671);
xnor UO_163 (O_163,N_19091,N_18920);
nand UO_164 (O_164,N_18122,N_16767);
nand UO_165 (O_165,N_19978,N_18855);
nor UO_166 (O_166,N_16742,N_19721);
xnor UO_167 (O_167,N_18510,N_18492);
or UO_168 (O_168,N_19593,N_18931);
or UO_169 (O_169,N_16067,N_19872);
and UO_170 (O_170,N_19084,N_19866);
nor UO_171 (O_171,N_19193,N_17645);
nand UO_172 (O_172,N_18888,N_18036);
or UO_173 (O_173,N_17070,N_16369);
or UO_174 (O_174,N_16851,N_18628);
xnor UO_175 (O_175,N_16994,N_19547);
xnor UO_176 (O_176,N_19067,N_17762);
and UO_177 (O_177,N_19976,N_16171);
nor UO_178 (O_178,N_16696,N_16207);
nand UO_179 (O_179,N_16479,N_17075);
nor UO_180 (O_180,N_18062,N_16424);
or UO_181 (O_181,N_18483,N_19496);
and UO_182 (O_182,N_19643,N_18307);
nor UO_183 (O_183,N_16026,N_18282);
nand UO_184 (O_184,N_16145,N_17823);
nor UO_185 (O_185,N_17714,N_18033);
or UO_186 (O_186,N_17629,N_19993);
and UO_187 (O_187,N_17067,N_18217);
or UO_188 (O_188,N_17634,N_16390);
or UO_189 (O_189,N_19734,N_19801);
or UO_190 (O_190,N_18779,N_19489);
nor UO_191 (O_191,N_18910,N_17908);
or UO_192 (O_192,N_16657,N_17772);
and UO_193 (O_193,N_19969,N_19950);
nand UO_194 (O_194,N_17979,N_18004);
xnor UO_195 (O_195,N_17150,N_16492);
and UO_196 (O_196,N_19062,N_17801);
xnor UO_197 (O_197,N_16748,N_17025);
or UO_198 (O_198,N_16300,N_16036);
xor UO_199 (O_199,N_19504,N_19083);
and UO_200 (O_200,N_16396,N_17056);
xnor UO_201 (O_201,N_18675,N_17126);
nand UO_202 (O_202,N_17661,N_19803);
xor UO_203 (O_203,N_16105,N_17357);
xor UO_204 (O_204,N_17812,N_17149);
nor UO_205 (O_205,N_17415,N_17238);
nor UO_206 (O_206,N_17726,N_16025);
nor UO_207 (O_207,N_16334,N_17544);
nand UO_208 (O_208,N_17555,N_19979);
nor UO_209 (O_209,N_17303,N_19136);
xnor UO_210 (O_210,N_16383,N_16999);
and UO_211 (O_211,N_18651,N_19566);
and UO_212 (O_212,N_18722,N_19123);
and UO_213 (O_213,N_16648,N_16848);
nand UO_214 (O_214,N_19704,N_19611);
nor UO_215 (O_215,N_16243,N_17254);
nand UO_216 (O_216,N_16482,N_17028);
and UO_217 (O_217,N_16109,N_16159);
and UO_218 (O_218,N_18727,N_16624);
nor UO_219 (O_219,N_18901,N_18372);
nor UO_220 (O_220,N_19434,N_17339);
or UO_221 (O_221,N_17319,N_17259);
nor UO_222 (O_222,N_18922,N_19706);
xor UO_223 (O_223,N_18763,N_17621);
and UO_224 (O_224,N_18289,N_17247);
or UO_225 (O_225,N_18242,N_18470);
or UO_226 (O_226,N_19322,N_16259);
xor UO_227 (O_227,N_16018,N_19807);
nor UO_228 (O_228,N_17826,N_19996);
and UO_229 (O_229,N_16541,N_17050);
and UO_230 (O_230,N_18229,N_18793);
nor UO_231 (O_231,N_16600,N_19712);
and UO_232 (O_232,N_18328,N_19906);
and UO_233 (O_233,N_18663,N_16783);
and UO_234 (O_234,N_16180,N_19988);
nor UO_235 (O_235,N_18380,N_16864);
xor UO_236 (O_236,N_16617,N_17226);
or UO_237 (O_237,N_19971,N_19835);
nand UO_238 (O_238,N_19924,N_16096);
or UO_239 (O_239,N_19275,N_17938);
nand UO_240 (O_240,N_17928,N_18237);
xor UO_241 (O_241,N_16603,N_17377);
and UO_242 (O_242,N_17763,N_16237);
and UO_243 (O_243,N_19607,N_17738);
nor UO_244 (O_244,N_19584,N_16578);
xor UO_245 (O_245,N_19184,N_16203);
nand UO_246 (O_246,N_18875,N_17855);
and UO_247 (O_247,N_18754,N_16097);
nand UO_248 (O_248,N_17061,N_18556);
and UO_249 (O_249,N_18241,N_19301);
nand UO_250 (O_250,N_17891,N_17802);
and UO_251 (O_251,N_16840,N_17691);
or UO_252 (O_252,N_16200,N_17919);
nor UO_253 (O_253,N_19980,N_18654);
and UO_254 (O_254,N_19328,N_19131);
xnor UO_255 (O_255,N_18864,N_17214);
nor UO_256 (O_256,N_17486,N_16012);
nand UO_257 (O_257,N_18132,N_16020);
xnor UO_258 (O_258,N_16608,N_16687);
or UO_259 (O_259,N_16750,N_16471);
nand UO_260 (O_260,N_19763,N_17131);
nand UO_261 (O_261,N_18604,N_19379);
and UO_262 (O_262,N_18106,N_18306);
xor UO_263 (O_263,N_16876,N_19348);
or UO_264 (O_264,N_16388,N_17833);
xnor UO_265 (O_265,N_17584,N_18295);
nor UO_266 (O_266,N_16136,N_16784);
nor UO_267 (O_267,N_18549,N_16956);
and UO_268 (O_268,N_17323,N_18680);
nand UO_269 (O_269,N_18737,N_16151);
and UO_270 (O_270,N_19233,N_16322);
xnor UO_271 (O_271,N_19899,N_19404);
nor UO_272 (O_272,N_19608,N_18301);
and UO_273 (O_273,N_18954,N_18899);
xor UO_274 (O_274,N_17391,N_18098);
xor UO_275 (O_275,N_19926,N_18167);
or UO_276 (O_276,N_19170,N_18339);
xor UO_277 (O_277,N_17369,N_17783);
xor UO_278 (O_278,N_17036,N_17804);
xor UO_279 (O_279,N_17677,N_16654);
nor UO_280 (O_280,N_16294,N_19179);
nand UO_281 (O_281,N_19147,N_19839);
and UO_282 (O_282,N_17417,N_16288);
nor UO_283 (O_283,N_19828,N_19232);
nand UO_284 (O_284,N_17069,N_17382);
nor UO_285 (O_285,N_19506,N_18746);
xor UO_286 (O_286,N_18733,N_18959);
nand UO_287 (O_287,N_18338,N_19664);
nor UO_288 (O_288,N_17237,N_16610);
or UO_289 (O_289,N_18068,N_19141);
nor UO_290 (O_290,N_18294,N_19020);
or UO_291 (O_291,N_18742,N_19648);
nor UO_292 (O_292,N_18133,N_17295);
nand UO_293 (O_293,N_16147,N_17317);
nand UO_294 (O_294,N_16179,N_19947);
xor UO_295 (O_295,N_16692,N_17552);
and UO_296 (O_296,N_16803,N_17916);
nor UO_297 (O_297,N_19851,N_19285);
or UO_298 (O_298,N_17894,N_19795);
xor UO_299 (O_299,N_19175,N_17176);
xor UO_300 (O_300,N_18005,N_16553);
nand UO_301 (O_301,N_19304,N_19462);
xnor UO_302 (O_302,N_17161,N_19367);
and UO_303 (O_303,N_18428,N_18063);
xor UO_304 (O_304,N_18511,N_19676);
or UO_305 (O_305,N_16724,N_18885);
or UO_306 (O_306,N_17038,N_16134);
or UO_307 (O_307,N_17572,N_16221);
nand UO_308 (O_308,N_17615,N_17824);
and UO_309 (O_309,N_17927,N_16596);
or UO_310 (O_310,N_19781,N_17682);
or UO_311 (O_311,N_19138,N_17694);
or UO_312 (O_312,N_19287,N_17605);
or UO_313 (O_313,N_16626,N_17776);
nand UO_314 (O_314,N_18906,N_16635);
nand UO_315 (O_315,N_16514,N_19655);
or UO_316 (O_316,N_19236,N_17098);
nand UO_317 (O_317,N_19754,N_18269);
xor UO_318 (O_318,N_18054,N_19891);
nor UO_319 (O_319,N_17383,N_16506);
and UO_320 (O_320,N_18420,N_18748);
or UO_321 (O_321,N_16865,N_18187);
or UO_322 (O_322,N_17110,N_16158);
and UO_323 (O_323,N_19122,N_16107);
and UO_324 (O_324,N_19837,N_16157);
nor UO_325 (O_325,N_19327,N_19838);
nand UO_326 (O_326,N_17794,N_17096);
xnor UO_327 (O_327,N_19480,N_19896);
and UO_328 (O_328,N_18495,N_18568);
nand UO_329 (O_329,N_18124,N_17593);
nor UO_330 (O_330,N_18115,N_16859);
nand UO_331 (O_331,N_16616,N_19197);
xor UO_332 (O_332,N_17771,N_16080);
and UO_333 (O_333,N_17587,N_17969);
and UO_334 (O_334,N_19684,N_18799);
or UO_335 (O_335,N_19408,N_18983);
xnor UO_336 (O_336,N_16428,N_16936);
xor UO_337 (O_337,N_18548,N_17981);
and UO_338 (O_338,N_17100,N_17297);
nand UO_339 (O_339,N_16649,N_16366);
nand UO_340 (O_340,N_18486,N_19037);
nor UO_341 (O_341,N_18882,N_18239);
nor UO_342 (O_342,N_19741,N_18760);
xor UO_343 (O_343,N_16272,N_18958);
nand UO_344 (O_344,N_18829,N_18755);
or UO_345 (O_345,N_18974,N_16987);
nor UO_346 (O_346,N_19247,N_16607);
nand UO_347 (O_347,N_16308,N_18172);
nand UO_348 (O_348,N_17500,N_16446);
and UO_349 (O_349,N_17086,N_16003);
nand UO_350 (O_350,N_18415,N_19873);
or UO_351 (O_351,N_17890,N_17082);
xor UO_352 (O_352,N_17856,N_16345);
nor UO_353 (O_353,N_19239,N_17750);
and UO_354 (O_354,N_16321,N_19423);
nand UO_355 (O_355,N_18145,N_19695);
nor UO_356 (O_356,N_16385,N_16703);
or UO_357 (O_357,N_19451,N_16443);
nand UO_358 (O_358,N_17732,N_17849);
nor UO_359 (O_359,N_18081,N_16431);
xnor UO_360 (O_360,N_17546,N_17314);
xor UO_361 (O_361,N_17130,N_18712);
or UO_362 (O_362,N_18693,N_18751);
or UO_363 (O_363,N_19078,N_18523);
and UO_364 (O_364,N_16873,N_16877);
nand UO_365 (O_365,N_19373,N_16732);
and UO_366 (O_366,N_19844,N_18402);
nor UO_367 (O_367,N_19011,N_17171);
or UO_368 (O_368,N_19799,N_18070);
xor UO_369 (O_369,N_18206,N_19101);
nand UO_370 (O_370,N_17747,N_16213);
xnor UO_371 (O_371,N_16813,N_18171);
nand UO_372 (O_372,N_18456,N_16869);
or UO_373 (O_373,N_17422,N_19266);
and UO_374 (O_374,N_18302,N_18661);
and UO_375 (O_375,N_17400,N_16350);
xor UO_376 (O_376,N_16309,N_17509);
or UO_377 (O_377,N_18388,N_16972);
nor UO_378 (O_378,N_19392,N_19004);
nor UO_379 (O_379,N_19772,N_17505);
nor UO_380 (O_380,N_16005,N_18230);
nand UO_381 (O_381,N_16124,N_18413);
or UO_382 (O_382,N_16371,N_19669);
nand UO_383 (O_383,N_19645,N_18406);
or UO_384 (O_384,N_18009,N_16547);
and UO_385 (O_385,N_19228,N_17285);
or UO_386 (O_386,N_18478,N_18150);
or UO_387 (O_387,N_19700,N_16353);
xor UO_388 (O_388,N_19879,N_18039);
xnor UO_389 (O_389,N_17439,N_18987);
and UO_390 (O_390,N_18463,N_19794);
nand UO_391 (O_391,N_17695,N_19771);
or UO_392 (O_392,N_19230,N_18476);
xnor UO_393 (O_393,N_16573,N_18012);
or UO_394 (O_394,N_16181,N_18813);
and UO_395 (O_395,N_16236,N_19364);
nand UO_396 (O_396,N_19647,N_17031);
or UO_397 (O_397,N_16745,N_18662);
nor UO_398 (O_398,N_18078,N_19719);
nor UO_399 (O_399,N_19768,N_18034);
nand UO_400 (O_400,N_16264,N_17915);
nand UO_401 (O_401,N_16086,N_16918);
or UO_402 (O_402,N_19511,N_16472);
or UO_403 (O_403,N_18092,N_17245);
xor UO_404 (O_404,N_19255,N_17565);
or UO_405 (O_405,N_19736,N_16331);
nor UO_406 (O_406,N_17266,N_18682);
nor UO_407 (O_407,N_17865,N_16699);
and UO_408 (O_408,N_18504,N_16401);
nand UO_409 (O_409,N_17088,N_18505);
and UO_410 (O_410,N_19623,N_17551);
or UO_411 (O_411,N_19882,N_19620);
and UO_412 (O_412,N_19139,N_19460);
and UO_413 (O_413,N_17425,N_16224);
and UO_414 (O_414,N_19386,N_16028);
or UO_415 (O_415,N_17491,N_18804);
or UO_416 (O_416,N_16330,N_16302);
or UO_417 (O_417,N_19278,N_17332);
or UO_418 (O_418,N_16512,N_19010);
xor UO_419 (O_419,N_17355,N_17206);
nand UO_420 (O_420,N_17701,N_17513);
nand UO_421 (O_421,N_16964,N_17289);
and UO_422 (O_422,N_18258,N_17047);
xnor UO_423 (O_423,N_16265,N_16169);
nand UO_424 (O_424,N_16656,N_16631);
or UO_425 (O_425,N_19148,N_17309);
and UO_426 (O_426,N_18203,N_17352);
xor UO_427 (O_427,N_18417,N_16536);
nor UO_428 (O_428,N_16470,N_19939);
or UO_429 (O_429,N_16910,N_18213);
nor UO_430 (O_430,N_19850,N_19674);
and UO_431 (O_431,N_19665,N_18871);
or UO_432 (O_432,N_19048,N_17198);
nand UO_433 (O_433,N_17600,N_16976);
nor UO_434 (O_434,N_18366,N_19809);
xor UO_435 (O_435,N_16202,N_16033);
and UO_436 (O_436,N_16780,N_18839);
and UO_437 (O_437,N_19267,N_16658);
and UO_438 (O_438,N_16115,N_16718);
xor UO_439 (O_439,N_18814,N_17434);
xnor UO_440 (O_440,N_19436,N_18543);
xnor UO_441 (O_441,N_19249,N_17464);
or UO_442 (O_442,N_17921,N_17869);
nand UO_443 (O_443,N_16360,N_16681);
nand UO_444 (O_444,N_18351,N_17854);
nor UO_445 (O_445,N_17971,N_17527);
nand UO_446 (O_446,N_17523,N_17719);
nand UO_447 (O_447,N_18317,N_17773);
nand UO_448 (O_448,N_18745,N_17624);
and UO_449 (O_449,N_18580,N_18175);
nor UO_450 (O_450,N_18455,N_16044);
nand UO_451 (O_451,N_19492,N_18074);
or UO_452 (O_452,N_16737,N_18238);
nor UO_453 (O_453,N_17330,N_19792);
nand UO_454 (O_454,N_16849,N_16439);
nor UO_455 (O_455,N_17566,N_17395);
and UO_456 (O_456,N_18724,N_16828);
xnor UO_457 (O_457,N_18393,N_19709);
and UO_458 (O_458,N_18718,N_19295);
or UO_459 (O_459,N_19113,N_17602);
nor UO_460 (O_460,N_18143,N_17723);
and UO_461 (O_461,N_17483,N_19717);
nand UO_462 (O_462,N_19009,N_19619);
or UO_463 (O_463,N_17592,N_17904);
xnor UO_464 (O_464,N_17215,N_18164);
nand UO_465 (O_465,N_19773,N_18971);
nor UO_466 (O_466,N_16072,N_16327);
and UO_467 (O_467,N_19129,N_16214);
and UO_468 (O_468,N_18196,N_19111);
and UO_469 (O_469,N_16199,N_18458);
or UO_470 (O_470,N_16807,N_19412);
nor UO_471 (O_471,N_17984,N_18646);
nor UO_472 (O_472,N_16103,N_16139);
nand UO_473 (O_473,N_17481,N_17957);
nor UO_474 (O_474,N_19488,N_19237);
nor UO_475 (O_475,N_16664,N_18061);
or UO_476 (O_476,N_19907,N_16442);
nor UO_477 (O_477,N_19263,N_16283);
nor UO_478 (O_478,N_17416,N_19535);
xnor UO_479 (O_479,N_18273,N_19325);
or UO_480 (O_480,N_16762,N_17716);
xor UO_481 (O_481,N_18766,N_18826);
and UO_482 (O_482,N_19225,N_19894);
and UO_483 (O_483,N_18473,N_16619);
or UO_484 (O_484,N_18221,N_19682);
or UO_485 (O_485,N_16146,N_18116);
nor UO_486 (O_486,N_19689,N_18015);
and UO_487 (O_487,N_16827,N_18508);
or UO_488 (O_488,N_19743,N_18365);
and UO_489 (O_489,N_17106,N_19595);
xnor UO_490 (O_490,N_18064,N_18607);
or UO_491 (O_491,N_18430,N_17667);
and UO_492 (O_492,N_17737,N_16786);
nor UO_493 (O_493,N_19105,N_18071);
and UO_494 (O_494,N_17021,N_19168);
xor UO_495 (O_495,N_16609,N_16451);
nor UO_496 (O_496,N_19368,N_19942);
xor UO_497 (O_497,N_16676,N_19452);
or UO_498 (O_498,N_18743,N_17006);
xnor UO_499 (O_499,N_16824,N_18364);
or UO_500 (O_500,N_19025,N_18429);
and UO_501 (O_501,N_17046,N_18632);
and UO_502 (O_502,N_19118,N_16815);
or UO_503 (O_503,N_18848,N_17548);
xnor UO_504 (O_504,N_17079,N_17458);
nor UO_505 (O_505,N_17966,N_17044);
xor UO_506 (O_506,N_18978,N_16423);
and UO_507 (O_507,N_17530,N_18412);
nand UO_508 (O_508,N_16421,N_17992);
or UO_509 (O_509,N_19366,N_18583);
xnor UO_510 (O_510,N_19533,N_19530);
and UO_511 (O_511,N_16576,N_16053);
xor UO_512 (O_512,N_18788,N_19213);
xor UO_513 (O_513,N_16287,N_18570);
xor UO_514 (O_514,N_19725,N_18835);
nor UO_515 (O_515,N_19218,N_16293);
and UO_516 (O_516,N_19789,N_17576);
and UO_517 (O_517,N_16381,N_18994);
or UO_518 (O_518,N_19095,N_17385);
nand UO_519 (O_519,N_19812,N_18617);
and UO_520 (O_520,N_18292,N_16574);
and UO_521 (O_521,N_19072,N_19094);
xnor UO_522 (O_522,N_17522,N_18474);
and UO_523 (O_523,N_18442,N_17490);
nor UO_524 (O_524,N_18537,N_17354);
nand UO_525 (O_525,N_18083,N_17879);
or UO_526 (O_526,N_19042,N_18943);
nor UO_527 (O_527,N_19341,N_16906);
xor UO_528 (O_528,N_19294,N_17935);
and UO_529 (O_529,N_17074,N_18687);
and UO_530 (O_530,N_19999,N_19432);
xnor UO_531 (O_531,N_18710,N_17340);
nand UO_532 (O_532,N_16789,N_19690);
nand UO_533 (O_533,N_18658,N_16695);
or UO_534 (O_534,N_18201,N_19277);
and UO_535 (O_535,N_19409,N_18136);
xnor UO_536 (O_536,N_17426,N_19868);
and UO_537 (O_537,N_17724,N_18872);
and UO_538 (O_538,N_19598,N_19207);
nand UO_539 (O_539,N_18384,N_16647);
nor UO_540 (O_540,N_17610,N_16919);
or UO_541 (O_541,N_16437,N_16763);
or UO_542 (O_542,N_18284,N_19808);
nor UO_543 (O_543,N_17022,N_17186);
nor UO_544 (O_544,N_19858,N_19816);
xor UO_545 (O_545,N_19150,N_18884);
xnor UO_546 (O_546,N_18961,N_17389);
xor UO_547 (O_547,N_18660,N_16728);
nor UO_548 (O_548,N_16054,N_16751);
xor UO_549 (O_549,N_19628,N_18014);
xnor UO_550 (O_550,N_17147,N_17573);
and UO_551 (O_551,N_18587,N_17950);
nand UO_552 (O_552,N_17279,N_16605);
nand UO_553 (O_553,N_19444,N_16176);
nor UO_554 (O_554,N_18157,N_19845);
nand UO_555 (O_555,N_19961,N_17805);
xnor UO_556 (O_556,N_19574,N_16822);
nor UO_557 (O_557,N_16975,N_17713);
nor UO_558 (O_558,N_17476,N_17990);
or UO_559 (O_559,N_18330,N_18605);
nor UO_560 (O_560,N_16349,N_18358);
xor UO_561 (O_561,N_18801,N_18941);
xor UO_562 (O_562,N_19058,N_16277);
nand UO_563 (O_563,N_17851,N_19982);
xor UO_564 (O_564,N_17097,N_18467);
xor UO_565 (O_565,N_18013,N_17471);
and UO_566 (O_566,N_19804,N_16979);
nor UO_567 (O_567,N_19813,N_18152);
xor UO_568 (O_568,N_18708,N_18528);
nor UO_569 (O_569,N_19120,N_16337);
or UO_570 (O_570,N_16240,N_18638);
and UO_571 (O_571,N_16582,N_19745);
nor UO_572 (O_572,N_17721,N_16968);
or UO_573 (O_573,N_19892,N_17268);
or UO_574 (O_574,N_19519,N_17993);
xnor UO_575 (O_575,N_19049,N_16613);
and UO_576 (O_576,N_18266,N_18985);
and UO_577 (O_577,N_17123,N_17349);
xor UO_578 (O_578,N_19463,N_19383);
nor UO_579 (O_579,N_16049,N_18991);
or UO_580 (O_580,N_16089,N_18798);
nor UO_581 (O_581,N_16211,N_19337);
nand UO_582 (O_582,N_18193,N_18892);
nor UO_583 (O_583,N_17468,N_19874);
nand UO_584 (O_584,N_19395,N_18896);
or UO_585 (O_585,N_16485,N_16969);
or UO_586 (O_586,N_16960,N_18027);
and UO_587 (O_587,N_18671,N_16121);
nor UO_588 (O_588,N_18427,N_17868);
xnor UO_589 (O_589,N_16425,N_16878);
nand UO_590 (O_590,N_17093,N_16820);
nand UO_591 (O_591,N_17543,N_19820);
xnor UO_592 (O_592,N_18432,N_17554);
nor UO_593 (O_593,N_18551,N_18182);
xor UO_594 (O_594,N_17455,N_16093);
or UO_595 (O_595,N_18323,N_16896);
xor UO_596 (O_596,N_16705,N_17213);
nor UO_597 (O_597,N_16268,N_17091);
nand UO_598 (O_598,N_19475,N_16543);
and UO_599 (O_599,N_17813,N_19718);
nand UO_600 (O_600,N_18525,N_17963);
or UO_601 (O_601,N_17911,N_19630);
nand UO_602 (O_602,N_19916,N_19448);
nand UO_603 (O_603,N_16465,N_16364);
and UO_604 (O_604,N_19770,N_19018);
and UO_605 (O_605,N_16315,N_16511);
or UO_606 (O_606,N_18863,N_16835);
nand UO_607 (O_607,N_19726,N_17655);
and UO_608 (O_608,N_18017,N_18726);
xor UO_609 (O_609,N_17607,N_16318);
and UO_610 (O_610,N_16312,N_19445);
xnor UO_611 (O_611,N_16746,N_17059);
nand UO_612 (O_612,N_17956,N_19545);
nor UO_613 (O_613,N_17944,N_16368);
or UO_614 (O_614,N_17051,N_16802);
and UO_615 (O_615,N_19660,N_17408);
xor UO_616 (O_616,N_17626,N_17586);
xnor UO_617 (O_617,N_18540,N_16189);
nand UO_618 (O_618,N_17270,N_16085);
nor UO_619 (O_619,N_18861,N_18363);
or UO_620 (O_620,N_16875,N_17899);
nor UO_621 (O_621,N_18904,N_17095);
nand UO_622 (O_622,N_16263,N_18927);
nor UO_623 (O_623,N_16119,N_19201);
nand UO_624 (O_624,N_16686,N_17913);
and UO_625 (O_625,N_18337,N_17508);
nand UO_626 (O_626,N_19585,N_19922);
nand UO_627 (O_627,N_19521,N_17078);
or UO_628 (O_628,N_18667,N_17658);
or UO_629 (O_629,N_18948,N_18207);
nand UO_630 (O_630,N_18616,N_16296);
and UO_631 (O_631,N_17775,N_19621);
and UO_632 (O_632,N_19787,N_18840);
or UO_633 (O_633,N_16707,N_18031);
nor UO_634 (O_634,N_18623,N_16427);
xor UO_635 (O_635,N_17947,N_18786);
or UO_636 (O_636,N_18553,N_16805);
or UO_637 (O_637,N_18701,N_19036);
and UO_638 (O_638,N_19715,N_18819);
nor UO_639 (O_639,N_19537,N_18685);
xnor UO_640 (O_640,N_16210,N_17414);
and UO_641 (O_641,N_17258,N_16501);
nor UO_642 (O_642,N_18841,N_18516);
or UO_643 (O_643,N_19663,N_19167);
or UO_644 (O_644,N_17077,N_19705);
nand UO_645 (O_645,N_18210,N_17440);
xor UO_646 (O_646,N_16565,N_16418);
xnor UO_647 (O_647,N_19626,N_17568);
nand UO_648 (O_648,N_19666,N_19699);
or UO_649 (O_649,N_18891,N_19202);
or UO_650 (O_650,N_18902,N_19483);
nor UO_651 (O_651,N_18228,N_17341);
xor UO_652 (O_652,N_19510,N_16374);
or UO_653 (O_653,N_18274,N_17477);
or UO_654 (O_654,N_16944,N_17815);
xor UO_655 (O_655,N_18598,N_18060);
or UO_656 (O_656,N_16379,N_18789);
and UO_657 (O_657,N_16946,N_17799);
or UO_658 (O_658,N_19331,N_17688);
nor UO_659 (O_659,N_16529,N_16794);
xor UO_660 (O_660,N_16127,N_17361);
nand UO_661 (O_661,N_17652,N_19075);
xor UO_662 (O_662,N_17221,N_17517);
nor UO_663 (O_663,N_19994,N_18732);
nor UO_664 (O_664,N_16554,N_18905);
nand UO_665 (O_665,N_17895,N_19254);
or UO_666 (O_666,N_16953,N_16208);
nor UO_667 (O_667,N_18202,N_17564);
nand UO_668 (O_668,N_17166,N_18399);
or UO_669 (O_669,N_18409,N_17461);
nand UO_670 (O_670,N_16674,N_16370);
or UO_671 (O_671,N_18593,N_19221);
or UO_672 (O_672,N_17301,N_19934);
nand UO_673 (O_673,N_19629,N_19241);
or UO_674 (O_674,N_16810,N_16435);
nor UO_675 (O_675,N_18759,N_18979);
or UO_676 (O_676,N_19897,N_18996);
nand UO_677 (O_677,N_18833,N_18967);
or UO_678 (O_678,N_18609,N_18590);
or UO_679 (O_679,N_17871,N_16027);
and UO_680 (O_680,N_16419,N_16252);
xor UO_681 (O_681,N_19400,N_17203);
nor UO_682 (O_682,N_17387,N_17298);
nor UO_683 (O_683,N_17411,N_16954);
nor UO_684 (O_684,N_18889,N_19477);
and UO_685 (O_685,N_16411,N_17683);
nand UO_686 (O_686,N_17620,N_16123);
or UO_687 (O_687,N_16540,N_18962);
nand UO_688 (O_688,N_16862,N_18454);
and UO_689 (O_689,N_17660,N_16866);
nand UO_690 (O_690,N_17068,N_18250);
and UO_691 (O_691,N_18810,N_19443);
nor UO_692 (O_692,N_19406,N_19798);
nand UO_693 (O_693,N_16967,N_17489);
or UO_694 (O_694,N_16843,N_17518);
xor UO_695 (O_695,N_17898,N_16685);
xor UO_696 (O_696,N_17757,N_19397);
nor UO_697 (O_697,N_19544,N_18262);
xor UO_698 (O_698,N_16634,N_16888);
and UO_699 (O_699,N_17735,N_19426);
xor UO_700 (O_700,N_18006,N_17284);
and UO_701 (O_701,N_18446,N_18673);
and UO_702 (O_702,N_16301,N_19854);
and UO_703 (O_703,N_16893,N_17162);
nor UO_704 (O_704,N_17764,N_18536);
nor UO_705 (O_705,N_17407,N_17870);
or UO_706 (O_706,N_19546,N_18311);
nand UO_707 (O_707,N_16040,N_16867);
xor UO_708 (O_708,N_16868,N_17165);
nand UO_709 (O_709,N_19022,N_17766);
nand UO_710 (O_710,N_17560,N_17463);
xnor UO_711 (O_711,N_18189,N_18496);
nor UO_712 (O_712,N_17250,N_17529);
and UO_713 (O_713,N_17085,N_19424);
nand UO_714 (O_714,N_17485,N_16623);
nand UO_715 (O_715,N_18966,N_17212);
and UO_716 (O_716,N_16845,N_17080);
nor UO_717 (O_717,N_16478,N_18357);
or UO_718 (O_718,N_16666,N_17803);
nand UO_719 (O_719,N_19815,N_19834);
and UO_720 (O_720,N_19377,N_19501);
nor UO_721 (O_721,N_16187,N_18488);
and UO_722 (O_722,N_17055,N_17983);
xnor UO_723 (O_723,N_19948,N_16463);
xnor UO_724 (O_724,N_16955,N_16197);
xor UO_725 (O_725,N_18585,N_16487);
nor UO_726 (O_726,N_18000,N_18394);
nor UO_727 (O_727,N_17333,N_17722);
or UO_728 (O_728,N_19991,N_19482);
or UO_729 (O_729,N_17867,N_19143);
or UO_730 (O_730,N_16032,N_19673);
or UO_731 (O_731,N_17375,N_17578);
and UO_732 (O_732,N_17810,N_16998);
and UO_733 (O_733,N_17603,N_17350);
or UO_734 (O_734,N_16898,N_18459);
nor UO_735 (O_735,N_19029,N_16899);
or UO_736 (O_736,N_18329,N_19677);
nor UO_737 (O_737,N_18812,N_16148);
and UO_738 (O_738,N_19465,N_19453);
xnor UO_739 (O_739,N_19104,N_19313);
and UO_740 (O_740,N_18655,N_17630);
nand UO_741 (O_741,N_18386,N_19097);
and UO_742 (O_742,N_17536,N_16467);
nand UO_743 (O_743,N_18240,N_19108);
and UO_744 (O_744,N_17943,N_19740);
nand UO_745 (O_745,N_19871,N_17519);
nor UO_746 (O_746,N_17190,N_17907);
nor UO_747 (O_747,N_17241,N_16962);
xnor UO_748 (O_748,N_17153,N_17374);
xnor UO_749 (O_749,N_17052,N_19459);
nand UO_750 (O_750,N_19073,N_18360);
or UO_751 (O_751,N_17553,N_19780);
and UO_752 (O_752,N_18090,N_19188);
xor UO_753 (O_753,N_19568,N_18044);
nand UO_754 (O_754,N_16460,N_18041);
nand UO_755 (O_755,N_17700,N_19245);
xor UO_756 (O_756,N_17539,N_18714);
and UO_757 (O_757,N_16909,N_16505);
nor UO_758 (O_758,N_17952,N_16930);
xnor UO_759 (O_759,N_19421,N_17888);
nor UO_760 (O_760,N_18468,N_17459);
nand UO_761 (O_761,N_17469,N_17731);
and UO_762 (O_762,N_19756,N_17117);
nor UO_763 (O_763,N_17020,N_17989);
nand UO_764 (O_764,N_16056,N_18784);
or UO_765 (O_765,N_18140,N_19155);
or UO_766 (O_766,N_16048,N_19045);
or UO_767 (O_767,N_16650,N_19309);
nor UO_768 (O_768,N_16860,N_19923);
or UO_769 (O_769,N_17346,N_16447);
xor UO_770 (O_770,N_17138,N_18101);
xor UO_771 (O_771,N_17756,N_17386);
xor UO_772 (O_772,N_19089,N_18208);
nand UO_773 (O_773,N_18346,N_17424);
or UO_774 (O_774,N_19548,N_16934);
xnor UO_775 (O_775,N_18002,N_19286);
or UO_776 (O_776,N_16462,N_16620);
xor UO_777 (O_777,N_16094,N_16261);
nand UO_778 (O_778,N_18019,N_18043);
and UO_779 (O_779,N_18934,N_17625);
nand UO_780 (O_780,N_19657,N_17846);
and UO_781 (O_781,N_17743,N_17759);
xor UO_782 (O_782,N_16537,N_16035);
xor UO_783 (O_783,N_17831,N_18656);
xnor UO_784 (O_784,N_16004,N_17393);
nand UO_785 (O_785,N_18310,N_16564);
xor UO_786 (O_786,N_18612,N_18533);
xor UO_787 (O_787,N_19403,N_17670);
nand UO_788 (O_788,N_19464,N_16889);
and UO_789 (O_789,N_19054,N_16061);
or UO_790 (O_790,N_19538,N_17834);
xor UO_791 (O_791,N_16351,N_16725);
or UO_792 (O_792,N_18606,N_17549);
nand UO_793 (O_793,N_17023,N_16709);
and UO_794 (O_794,N_16682,N_16024);
nor UO_795 (O_795,N_19438,N_16526);
and UO_796 (O_796,N_16254,N_17184);
nor UO_797 (O_797,N_17099,N_16844);
nand UO_798 (O_798,N_16128,N_17436);
nand UO_799 (O_799,N_19883,N_19479);
nand UO_800 (O_800,N_19393,N_16765);
and UO_801 (O_801,N_16793,N_19499);
nor UO_802 (O_802,N_17418,N_19137);
and UO_803 (O_803,N_16324,N_18695);
nor UO_804 (O_804,N_16510,N_17431);
xnor UO_805 (O_805,N_19616,N_18449);
nand UO_806 (O_806,N_18391,N_17863);
and UO_807 (O_807,N_16356,N_18138);
nor UO_808 (O_808,N_18355,N_18254);
nand UO_809 (O_809,N_17591,N_18147);
nand UO_810 (O_810,N_17348,N_17703);
nand UO_811 (O_811,N_16598,N_17962);
nand UO_812 (O_812,N_16963,N_17945);
or UO_813 (O_813,N_17252,N_17599);
xor UO_814 (O_814,N_18315,N_18091);
nor UO_815 (O_815,N_17478,N_18717);
and UO_816 (O_816,N_17842,N_19502);
or UO_817 (O_817,N_19378,N_17207);
or UO_818 (O_818,N_19356,N_17199);
xor UO_819 (O_819,N_17588,N_18095);
and UO_820 (O_820,N_18344,N_17413);
nor UO_821 (O_821,N_19955,N_19116);
or UO_822 (O_822,N_19028,N_17848);
nand UO_823 (O_823,N_19678,N_19884);
nand UO_824 (O_824,N_17310,N_17745);
and UO_825 (O_825,N_17648,N_19334);
nand UO_826 (O_826,N_16068,N_18886);
and UO_827 (O_827,N_18610,N_19130);
nand UO_828 (O_828,N_18153,N_16289);
nor UO_829 (O_829,N_19634,N_17065);
xor UO_830 (O_830,N_18757,N_17937);
xor UO_831 (O_831,N_17976,N_18480);
and UO_832 (O_832,N_17427,N_16354);
and UO_833 (O_833,N_17475,N_18161);
and UO_834 (O_834,N_16429,N_19900);
nand UO_835 (O_835,N_17401,N_16209);
xor UO_836 (O_836,N_16149,N_18770);
xnor UO_837 (O_837,N_17109,N_16662);
nand UO_838 (O_838,N_16069,N_18199);
nor UO_839 (O_839,N_18802,N_17370);
nor UO_840 (O_840,N_18371,N_19959);
nor UO_841 (O_841,N_16445,N_17687);
and UO_842 (O_842,N_17373,N_16082);
and UO_843 (O_843,N_17029,N_17836);
or UO_844 (O_844,N_19875,N_18050);
or UO_845 (O_845,N_19945,N_19032);
nand UO_846 (O_846,N_16903,N_19825);
xnor UO_847 (O_847,N_18823,N_16365);
nand UO_848 (O_848,N_18322,N_19570);
nand UO_849 (O_849,N_18320,N_17883);
and UO_850 (O_850,N_17657,N_16897);
and UO_851 (O_851,N_19079,N_16394);
nor UO_852 (O_852,N_17598,N_19355);
nor UO_853 (O_853,N_17265,N_16144);
or UO_854 (O_854,N_18285,N_17767);
and UO_855 (O_855,N_17924,N_18341);
or UO_856 (O_856,N_19474,N_19314);
nand UO_857 (O_857,N_18016,N_18127);
or UO_858 (O_858,N_18318,N_16782);
nor UO_859 (O_859,N_17026,N_19310);
and UO_860 (O_860,N_18519,N_19338);
and UO_861 (O_861,N_18895,N_19555);
xor UO_862 (O_862,N_17343,N_19653);
or UO_863 (O_863,N_16407,N_19928);
and UO_864 (O_864,N_17209,N_17727);
or UO_865 (O_865,N_18691,N_17965);
xor UO_866 (O_866,N_16404,N_19389);
nor UO_867 (O_867,N_17752,N_19442);
nor UO_868 (O_868,N_18502,N_17403);
or UO_869 (O_869,N_18876,N_18603);
or UO_870 (O_870,N_18666,N_19577);
nor UO_871 (O_871,N_19128,N_16415);
xor UO_872 (O_872,N_16310,N_16766);
nand UO_873 (O_873,N_19273,N_17040);
xor UO_874 (O_874,N_17542,N_19208);
nor UO_875 (O_875,N_16313,N_19602);
nor UO_876 (O_876,N_19281,N_19774);
and UO_877 (O_877,N_19369,N_19877);
and UO_878 (O_878,N_16392,N_19087);
nand UO_879 (O_879,N_17073,N_17681);
and UO_880 (O_880,N_16160,N_18572);
xnor UO_881 (O_881,N_19380,N_16567);
and UO_882 (O_882,N_19696,N_18592);
xnor UO_883 (O_883,N_19210,N_18982);
nor UO_884 (O_884,N_16132,N_18574);
nor UO_885 (O_885,N_19956,N_16373);
xnor UO_886 (O_886,N_19023,N_19797);
nor UO_887 (O_887,N_17380,N_16077);
or UO_888 (O_888,N_18547,N_19583);
and UO_889 (O_889,N_17102,N_16642);
and UO_890 (O_890,N_16138,N_16778);
nand UO_891 (O_891,N_19160,N_17973);
nor UO_892 (O_892,N_17187,N_17754);
nor UO_893 (O_893,N_19166,N_16083);
nand UO_894 (O_894,N_18741,N_18728);
nor UO_895 (O_895,N_19439,N_19724);
nor UO_896 (O_896,N_19169,N_19728);
and UO_897 (O_897,N_16062,N_16806);
or UO_898 (O_898,N_18613,N_16059);
nand UO_899 (O_899,N_18227,N_17644);
xnor UO_900 (O_900,N_16850,N_16192);
and UO_901 (O_901,N_19405,N_16638);
nor UO_902 (O_902,N_17507,N_19910);
xnor UO_903 (O_903,N_19777,N_18621);
nor UO_904 (O_904,N_16432,N_18345);
and UO_905 (O_905,N_19242,N_19842);
nor UO_906 (O_906,N_17623,N_18052);
and UO_907 (O_907,N_19349,N_16100);
or UO_908 (O_908,N_17498,N_19823);
nand UO_909 (O_909,N_16218,N_19490);
xnor UO_910 (O_910,N_16890,N_17557);
and UO_911 (O_911,N_17967,N_19867);
xor UO_912 (O_912,N_19654,N_17707);
nand UO_913 (O_913,N_16579,N_16990);
and UO_914 (O_914,N_18925,N_18707);
or UO_915 (O_915,N_19800,N_18327);
nand UO_916 (O_916,N_18600,N_18542);
or UO_917 (O_917,N_16389,N_18988);
nand UO_918 (O_918,N_16174,N_17291);
and UO_919 (O_919,N_19158,N_18530);
and UO_920 (O_920,N_18200,N_17991);
nor UO_921 (O_921,N_17115,N_19680);
nand UO_922 (O_922,N_19125,N_16226);
and UO_923 (O_923,N_17202,N_18249);
and UO_924 (O_924,N_18424,N_18781);
or UO_925 (O_925,N_18776,N_17673);
nor UO_926 (O_926,N_18837,N_18818);
nor UO_927 (O_927,N_16531,N_19227);
xor UO_928 (O_928,N_17140,N_18162);
nand UO_929 (O_929,N_16397,N_17817);
and UO_930 (O_930,N_17039,N_17367);
nor UO_931 (O_931,N_18834,N_17010);
nand UO_932 (O_932,N_18264,N_17873);
nand UO_933 (O_933,N_16738,N_18563);
nand UO_934 (O_934,N_18842,N_17665);
nand UO_935 (O_935,N_19250,N_17092);
xnor UO_936 (O_936,N_18287,N_19468);
nor UO_937 (O_937,N_16761,N_18188);
nor UO_938 (O_938,N_18383,N_17933);
nand UO_939 (O_939,N_19836,N_16597);
nand UO_940 (O_940,N_19248,N_17547);
nand UO_941 (O_941,N_16483,N_19413);
or UO_942 (O_942,N_18491,N_18298);
nor UO_943 (O_943,N_16534,N_19110);
nor UO_944 (O_944,N_18280,N_19365);
nor UO_945 (O_945,N_19319,N_18047);
and UO_946 (O_946,N_16241,N_19203);
xnor UO_947 (O_947,N_16450,N_16279);
nand UO_948 (O_948,N_17451,N_19856);
nand UO_949 (O_949,N_16276,N_18382);
or UO_950 (O_950,N_16950,N_16271);
nor UO_951 (O_951,N_18163,N_16066);
xnor UO_952 (O_952,N_18001,N_19068);
or UO_953 (O_953,N_19472,N_17635);
and UO_954 (O_954,N_18170,N_19732);
or UO_955 (O_955,N_19738,N_18211);
or UO_956 (O_956,N_16332,N_16717);
and UO_957 (O_957,N_19592,N_17347);
or UO_958 (O_958,N_17639,N_18964);
nor UO_959 (O_959,N_19026,N_18868);
and UO_960 (O_960,N_18811,N_17613);
xor UO_961 (O_961,N_16057,N_16466);
xnor UO_962 (O_962,N_19846,N_18903);
nor UO_963 (O_963,N_19633,N_16143);
and UO_964 (O_964,N_17860,N_17583);
nor UO_965 (O_965,N_19050,N_18121);
xor UO_966 (O_966,N_17906,N_17540);
nor UO_967 (O_967,N_16595,N_16129);
or UO_968 (O_968,N_17084,N_16913);
xor UO_969 (O_969,N_17760,N_17852);
or UO_970 (O_970,N_16520,N_16804);
xnor UO_971 (O_971,N_19753,N_16575);
or UO_972 (O_972,N_16305,N_18771);
or UO_973 (O_973,N_17736,N_17229);
and UO_974 (O_974,N_19830,N_16230);
nor UO_975 (O_975,N_19288,N_19525);
or UO_976 (O_976,N_19119,N_19729);
and UO_977 (O_977,N_19190,N_18416);
and UO_978 (O_978,N_17143,N_19559);
nand UO_979 (O_979,N_16966,N_19505);
nand UO_980 (O_980,N_18448,N_18506);
nor UO_981 (O_981,N_17637,N_19814);
xor UO_982 (O_982,N_19157,N_18392);
and UO_983 (O_983,N_19066,N_16571);
or UO_984 (O_984,N_16677,N_16494);
and UO_985 (O_985,N_16733,N_18952);
xor UO_986 (O_986,N_17686,N_17178);
or UO_987 (O_987,N_16646,N_18144);
and UO_988 (O_988,N_17970,N_17520);
nor UO_989 (O_989,N_18867,N_18247);
nor UO_990 (O_990,N_16842,N_17054);
and UO_991 (O_991,N_17435,N_18643);
and UO_992 (O_992,N_19550,N_18023);
xor UO_993 (O_993,N_18020,N_16417);
or UO_994 (O_994,N_16140,N_19513);
and UO_995 (O_995,N_16535,N_18130);
or UO_996 (O_996,N_18191,N_18866);
or UO_997 (O_997,N_16989,N_19707);
nand UO_998 (O_998,N_16060,N_19599);
nor UO_999 (O_999,N_18844,N_18550);
and UO_1000 (O_1000,N_17881,N_19852);
xnor UO_1001 (O_1001,N_19428,N_19420);
and UO_1002 (O_1002,N_19627,N_18591);
xor UO_1003 (O_1003,N_16978,N_17875);
and UO_1004 (O_1004,N_17589,N_16031);
or UO_1005 (O_1005,N_16614,N_17985);
and UO_1006 (O_1006,N_16716,N_17934);
xor UO_1007 (O_1007,N_19384,N_18713);
nor UO_1008 (O_1008,N_17741,N_19019);
nor UO_1009 (O_1009,N_16731,N_19543);
and UO_1010 (O_1010,N_19640,N_18046);
nor UO_1011 (O_1011,N_19636,N_17225);
nor UO_1012 (O_1012,N_18303,N_19046);
or UO_1013 (O_1013,N_16773,N_16560);
or UO_1014 (O_1014,N_18716,N_19422);
and UO_1015 (O_1015,N_18792,N_19391);
nand UO_1016 (O_1016,N_16861,N_16347);
or UO_1017 (O_1017,N_19495,N_17531);
and UO_1018 (O_1018,N_16348,N_16178);
and UO_1019 (O_1019,N_19071,N_16882);
nand UO_1020 (O_1020,N_16253,N_18897);
and UO_1021 (O_1021,N_16781,N_16922);
nor UO_1022 (O_1022,N_16580,N_19597);
nand UO_1023 (O_1023,N_16643,N_18253);
or UO_1024 (O_1024,N_16759,N_18434);
xor UO_1025 (O_1025,N_16900,N_16528);
nand UO_1026 (O_1026,N_17570,N_17316);
or UO_1027 (O_1027,N_18316,N_19401);
nand UO_1028 (O_1028,N_17830,N_18342);
nand UO_1029 (O_1029,N_18135,N_16747);
or UO_1030 (O_1030,N_18040,N_16644);
xor UO_1031 (O_1031,N_18531,N_17002);
and UO_1032 (O_1032,N_18824,N_19390);
nor UO_1033 (O_1033,N_17371,N_18461);
nand UO_1034 (O_1034,N_17835,N_17181);
nand UO_1035 (O_1035,N_19681,N_19644);
nand UO_1036 (O_1036,N_17248,N_18319);
nand UO_1037 (O_1037,N_17900,N_17951);
nand UO_1038 (O_1038,N_16198,N_19231);
and UO_1039 (O_1039,N_17861,N_19869);
nand UO_1040 (O_1040,N_17887,N_17653);
nor UO_1041 (O_1041,N_17685,N_19060);
xnor UO_1042 (O_1042,N_17923,N_17958);
nor UO_1043 (O_1043,N_19353,N_17496);
xor UO_1044 (O_1044,N_19027,N_17545);
or UO_1045 (O_1045,N_19723,N_18452);
nor UO_1046 (O_1046,N_16920,N_16041);
or UO_1047 (O_1047,N_18619,N_19276);
or UO_1048 (O_1048,N_19031,N_16833);
xor UO_1049 (O_1049,N_19102,N_19658);
and UO_1050 (O_1050,N_19316,N_19336);
xor UO_1051 (O_1051,N_16907,N_18220);
or UO_1052 (O_1052,N_16242,N_16713);
nand UO_1053 (O_1053,N_18794,N_18524);
nand UO_1054 (O_1054,N_18936,N_19388);
or UO_1055 (O_1055,N_16524,N_16923);
xnor UO_1056 (O_1056,N_19142,N_19981);
nor UO_1057 (O_1057,N_19099,N_17219);
nand UO_1058 (O_1058,N_16939,N_16116);
or UO_1059 (O_1059,N_16499,N_18065);
nor UO_1060 (O_1060,N_18324,N_16014);
and UO_1061 (O_1061,N_16172,N_16410);
and UO_1062 (O_1062,N_17574,N_16170);
nand UO_1063 (O_1063,N_19558,N_19359);
nand UO_1064 (O_1064,N_19549,N_19581);
or UO_1065 (O_1065,N_17884,N_16125);
xnor UO_1066 (O_1066,N_19251,N_18313);
and UO_1067 (O_1067,N_17689,N_17188);
nor UO_1068 (O_1068,N_18134,N_17482);
nand UO_1069 (O_1069,N_18212,N_18594);
and UO_1070 (O_1070,N_17882,N_16382);
nor UO_1071 (O_1071,N_17739,N_18816);
nand UO_1072 (O_1072,N_19077,N_19765);
nand UO_1073 (O_1073,N_19688,N_16983);
or UO_1074 (O_1074,N_17786,N_18244);
xnor UO_1075 (O_1075,N_17246,N_19716);
or UO_1076 (O_1076,N_17501,N_18077);
nor UO_1077 (O_1077,N_16101,N_16785);
and UO_1078 (O_1078,N_16719,N_19372);
or UO_1079 (O_1079,N_16384,N_17939);
xor UO_1080 (O_1080,N_17942,N_18251);
nor UO_1081 (O_1081,N_18333,N_19057);
or UO_1082 (O_1082,N_18998,N_17638);
nand UO_1083 (O_1083,N_16205,N_17806);
and UO_1084 (O_1084,N_17779,N_18479);
nor UO_1085 (O_1085,N_19805,N_18234);
or UO_1086 (O_1086,N_18775,N_18569);
and UO_1087 (O_1087,N_19904,N_17320);
and UO_1088 (O_1088,N_19024,N_19983);
xnor UO_1089 (O_1089,N_17541,N_18652);
and UO_1090 (O_1090,N_16901,N_17715);
xor UO_1091 (O_1091,N_17076,N_16092);
xnor UO_1092 (O_1092,N_19951,N_18796);
nor UO_1093 (O_1093,N_18037,N_19298);
nor UO_1094 (O_1094,N_16245,N_17263);
and UO_1095 (O_1095,N_19742,N_17112);
or UO_1096 (O_1096,N_16915,N_17293);
xor UO_1097 (O_1097,N_19282,N_19746);
and UO_1098 (O_1098,N_16561,N_16894);
xor UO_1099 (O_1099,N_18780,N_16569);
and UO_1100 (O_1100,N_17274,N_19600);
xor UO_1101 (O_1101,N_19455,N_18066);
and UO_1102 (O_1102,N_18304,N_19258);
xor UO_1103 (O_1103,N_19526,N_18670);
and UO_1104 (O_1104,N_17561,N_17013);
and UO_1105 (O_1105,N_16816,N_17753);
nor UO_1106 (O_1106,N_19466,N_18534);
nor UO_1107 (O_1107,N_17619,N_17902);
xor UO_1108 (O_1108,N_18586,N_18845);
xor UO_1109 (O_1109,N_19515,N_16949);
xor UO_1110 (O_1110,N_17335,N_19733);
nand UO_1111 (O_1111,N_18475,N_19730);
or UO_1112 (O_1112,N_18271,N_16217);
xnor UO_1113 (O_1113,N_18627,N_19624);
nand UO_1114 (O_1114,N_19284,N_19672);
nor UO_1115 (O_1115,N_19788,N_17452);
xnor UO_1116 (O_1116,N_16823,N_18618);
and UO_1117 (O_1117,N_18245,N_17271);
and UO_1118 (O_1118,N_17419,N_16475);
nand UO_1119 (O_1119,N_19778,N_19890);
nand UO_1120 (O_1120,N_18807,N_16611);
nor UO_1121 (O_1121,N_19297,N_16669);
xor UO_1122 (O_1122,N_16314,N_19635);
and UO_1123 (O_1123,N_18963,N_19051);
or UO_1124 (O_1124,N_16587,N_16323);
or UO_1125 (O_1125,N_19107,N_17844);
nor UO_1126 (O_1126,N_16285,N_17322);
xor UO_1127 (O_1127,N_19514,N_19339);
nor UO_1128 (O_1128,N_18900,N_16933);
xor UO_1129 (O_1129,N_18368,N_19958);
or UO_1130 (O_1130,N_17048,N_16945);
or UO_1131 (O_1131,N_18008,N_18815);
or UO_1132 (O_1132,N_17480,N_16675);
nor UO_1133 (O_1133,N_18777,N_17941);
xnor UO_1134 (O_1134,N_16251,N_19565);
and UO_1135 (O_1135,N_16491,N_16645);
xnor UO_1136 (O_1136,N_19843,N_17968);
or UO_1137 (O_1137,N_17466,N_16227);
nand UO_1138 (O_1138,N_17820,N_17594);
nand UO_1139 (O_1139,N_18949,N_16555);
nand UO_1140 (O_1140,N_17998,N_19790);
xor UO_1141 (O_1141,N_19006,N_16518);
and UO_1142 (O_1142,N_17974,N_18915);
nand UO_1143 (O_1143,N_16548,N_19936);
xor UO_1144 (O_1144,N_16325,N_17233);
xor UO_1145 (O_1145,N_16071,N_18797);
and UO_1146 (O_1146,N_16398,N_17729);
nor UO_1147 (O_1147,N_18644,N_19517);
or UO_1148 (O_1148,N_18749,N_19541);
nand UO_1149 (O_1149,N_17292,N_16438);
and UO_1150 (O_1150,N_16246,N_16058);
or UO_1151 (O_1151,N_16592,N_16995);
nand UO_1152 (O_1152,N_17744,N_16694);
or UO_1153 (O_1153,N_18851,N_19315);
nand UO_1154 (O_1154,N_18641,N_19694);
and UO_1155 (O_1155,N_17185,N_16530);
nor UO_1156 (O_1156,N_19195,N_17193);
and UO_1157 (O_1157,N_19470,N_16405);
and UO_1158 (O_1158,N_17428,N_16131);
and UO_1159 (O_1159,N_17005,N_17808);
and UO_1160 (O_1160,N_18546,N_16212);
xnor UO_1161 (O_1161,N_18057,N_17111);
or UO_1162 (O_1162,N_17057,N_18410);
nor UO_1163 (O_1163,N_18148,N_19943);
nand UO_1164 (O_1164,N_19154,N_18275);
nand UO_1165 (O_1165,N_17853,N_18808);
nand UO_1166 (O_1166,N_19069,N_19786);
or UO_1167 (O_1167,N_17495,N_16736);
xor UO_1168 (O_1168,N_18088,N_16734);
and UO_1169 (O_1169,N_17177,N_19752);
nor UO_1170 (O_1170,N_19407,N_16991);
nor UO_1171 (O_1171,N_16683,N_19199);
and UO_1172 (O_1172,N_17889,N_19571);
and UO_1173 (O_1173,N_19915,N_19833);
or UO_1174 (O_1174,N_18512,N_18385);
or UO_1175 (O_1175,N_19402,N_17313);
nand UO_1176 (O_1176,N_17453,N_18879);
and UO_1177 (O_1177,N_17089,N_18058);
nand UO_1178 (O_1178,N_19269,N_17579);
xor UO_1179 (O_1179,N_19625,N_16590);
or UO_1180 (O_1180,N_16038,N_18846);
xor UO_1181 (O_1181,N_19092,N_17769);
xor UO_1182 (O_1182,N_16286,N_18787);
or UO_1183 (O_1183,N_19831,N_18697);
and UO_1184 (O_1184,N_18919,N_18185);
or UO_1185 (O_1185,N_16155,N_19957);
xnor UO_1186 (O_1186,N_17562,N_18862);
nand UO_1187 (O_1187,N_18314,N_18139);
and UO_1188 (O_1188,N_18917,N_18296);
nand UO_1189 (O_1189,N_19234,N_18444);
nor UO_1190 (O_1190,N_16508,N_16023);
and UO_1191 (O_1191,N_16267,N_19667);
and UO_1192 (O_1192,N_18118,N_17785);
or UO_1193 (O_1193,N_18790,N_16257);
nand UO_1194 (O_1194,N_16362,N_19173);
and UO_1195 (O_1195,N_18117,N_18325);
and UO_1196 (O_1196,N_17276,N_17062);
xnor UO_1197 (O_1197,N_19115,N_18279);
xnor UO_1198 (O_1198,N_18390,N_19766);
nand UO_1199 (O_1199,N_17420,N_16079);
nand UO_1200 (O_1200,N_17484,N_19458);
xor UO_1201 (O_1201,N_18773,N_16817);
and UO_1202 (O_1202,N_16938,N_16223);
xnor UO_1203 (O_1203,N_16729,N_19174);
and UO_1204 (O_1204,N_17521,N_18806);
and UO_1205 (O_1205,N_19345,N_17182);
or UO_1206 (O_1206,N_17311,N_19012);
xor UO_1207 (O_1207,N_18290,N_18729);
nand UO_1208 (O_1208,N_17647,N_16837);
xnor UO_1209 (O_1209,N_16009,N_19963);
nor UO_1210 (O_1210,N_18683,N_19311);
nor UO_1211 (O_1211,N_17433,N_16303);
or UO_1212 (O_1212,N_16826,N_18466);
nand UO_1213 (O_1213,N_19649,N_17733);
or UO_1214 (O_1214,N_19933,N_19944);
nor UO_1215 (O_1215,N_16074,N_18226);
nor UO_1216 (O_1216,N_18235,N_18482);
or UO_1217 (O_1217,N_19806,N_17533);
and UO_1218 (O_1218,N_16739,N_17809);
and UO_1219 (O_1219,N_16924,N_18990);
xor UO_1220 (O_1220,N_19491,N_16391);
nand UO_1221 (O_1221,N_17601,N_16052);
or UO_1222 (O_1222,N_17472,N_16986);
nor UO_1223 (O_1223,N_18558,N_16408);
and UO_1224 (O_1224,N_17018,N_17720);
nor UO_1225 (O_1225,N_17249,N_18830);
nor UO_1226 (O_1226,N_17488,N_19109);
nor UO_1227 (O_1227,N_17571,N_16436);
and UO_1228 (O_1228,N_19257,N_17479);
or UO_1229 (O_1229,N_16839,N_17158);
or UO_1230 (O_1230,N_19346,N_17366);
xnor UO_1231 (O_1231,N_17327,N_18232);
nand UO_1232 (O_1232,N_18630,N_19361);
or UO_1233 (O_1233,N_18898,N_18944);
or UO_1234 (O_1234,N_17308,N_18857);
nor UO_1235 (O_1235,N_16075,N_18435);
nand UO_1236 (O_1236,N_16633,N_19056);
and UO_1237 (O_1237,N_17822,N_19711);
nor UO_1238 (O_1238,N_16800,N_18107);
or UO_1239 (O_1239,N_17230,N_16519);
xor UO_1240 (O_1240,N_16500,N_16872);
or UO_1241 (O_1241,N_17800,N_16338);
xnor UO_1242 (O_1242,N_18853,N_17262);
xor UO_1243 (O_1243,N_19398,N_16459);
nor UO_1244 (O_1244,N_19710,N_17774);
and UO_1245 (O_1245,N_18431,N_17559);
xnor UO_1246 (O_1246,N_16441,N_19927);
nor UO_1247 (O_1247,N_17631,N_18942);
or UO_1248 (O_1248,N_18126,N_16228);
nor UO_1249 (O_1249,N_18734,N_17789);
xor UO_1250 (O_1250,N_17359,N_18028);
nor UO_1251 (O_1251,N_17680,N_19307);
or UO_1252 (O_1252,N_19290,N_18581);
or UO_1253 (O_1253,N_18457,N_18576);
xnor UO_1254 (O_1254,N_16618,N_17342);
nand UO_1255 (O_1255,N_17876,N_16050);
or UO_1256 (O_1256,N_19291,N_17528);
and UO_1257 (O_1257,N_17811,N_18501);
xnor UO_1258 (O_1258,N_16444,N_18160);
xor UO_1259 (O_1259,N_19274,N_16776);
xnor UO_1260 (O_1260,N_18389,N_17307);
nor UO_1261 (O_1261,N_19450,N_16722);
or UO_1262 (O_1262,N_18560,N_17378);
nand UO_1263 (O_1263,N_17850,N_18049);
nor UO_1264 (O_1264,N_18353,N_19080);
nor UO_1265 (O_1265,N_16498,N_16760);
or UO_1266 (O_1266,N_16819,N_16175);
nand UO_1267 (O_1267,N_16940,N_18067);
nand UO_1268 (O_1268,N_16448,N_17345);
nor UO_1269 (O_1269,N_16743,N_16497);
nor UO_1270 (O_1270,N_19764,N_17510);
or UO_1271 (O_1271,N_16503,N_18517);
or UO_1272 (O_1272,N_16559,N_16916);
and UO_1273 (O_1273,N_18599,N_17094);
xnor UO_1274 (O_1274,N_17033,N_19132);
nand UO_1275 (O_1275,N_17228,N_17525);
xor UO_1276 (O_1276,N_16525,N_17917);
or UO_1277 (O_1277,N_16545,N_16651);
nand UO_1278 (O_1278,N_17512,N_19070);
xor UO_1279 (O_1279,N_17334,N_16911);
nand UO_1280 (O_1280,N_17273,N_17705);
xor UO_1281 (O_1281,N_16941,N_19968);
and UO_1282 (O_1282,N_17409,N_19903);
and UO_1283 (O_1283,N_18024,N_16591);
nor UO_1284 (O_1284,N_17172,N_18588);
and UO_1285 (O_1285,N_19779,N_19631);
and UO_1286 (O_1286,N_17041,N_16126);
and UO_1287 (O_1287,N_17454,N_19727);
xnor UO_1288 (O_1288,N_17959,N_16030);
xnor UO_1289 (O_1289,N_19153,N_17467);
or UO_1290 (O_1290,N_16190,N_18602);
nand UO_1291 (O_1291,N_18256,N_18109);
xor UO_1292 (O_1292,N_16630,N_17712);
or UO_1293 (O_1293,N_19235,N_19783);
nand UO_1294 (O_1294,N_18597,N_16925);
or UO_1295 (O_1295,N_18112,N_16792);
xnor UO_1296 (O_1296,N_17142,N_16250);
xor UO_1297 (O_1297,N_16672,N_17674);
and UO_1298 (O_1298,N_16163,N_16993);
xor UO_1299 (O_1299,N_16229,N_18557);
xor UO_1300 (O_1300,N_18887,N_17189);
nand UO_1301 (O_1301,N_18894,N_16295);
or UO_1302 (O_1302,N_19905,N_16948);
nand UO_1303 (O_1303,N_19222,N_19703);
xor UO_1304 (O_1304,N_19512,N_16606);
nand UO_1305 (O_1305,N_16403,N_19967);
xnor UO_1306 (O_1306,N_16266,N_18129);
or UO_1307 (O_1307,N_17175,N_18820);
nand UO_1308 (O_1308,N_19001,N_19848);
nand UO_1309 (O_1309,N_16852,N_18648);
nor UO_1310 (O_1310,N_19975,N_16568);
nand UO_1311 (O_1311,N_18183,N_18577);
xnor UO_1312 (O_1312,N_16275,N_17053);
nand UO_1313 (O_1313,N_19893,N_17103);
xnor UO_1314 (O_1314,N_16118,N_18114);
nand UO_1315 (O_1315,N_18222,N_18938);
and UO_1316 (O_1316,N_18270,N_17781);
nor UO_1317 (O_1317,N_16141,N_17141);
or UO_1318 (O_1318,N_19748,N_18433);
nand UO_1319 (O_1319,N_17678,N_16723);
and UO_1320 (O_1320,N_16957,N_16455);
nand UO_1321 (O_1321,N_17892,N_16749);
xor UO_1322 (O_1322,N_17146,N_17912);
nand UO_1323 (O_1323,N_19081,N_19911);
nand UO_1324 (O_1324,N_17120,N_18102);
or UO_1325 (O_1325,N_17717,N_19941);
xor UO_1326 (O_1326,N_17930,N_19751);
nand UO_1327 (O_1327,N_19209,N_17083);
nor UO_1328 (O_1328,N_18086,N_17932);
xnor UO_1329 (O_1329,N_19382,N_18870);
nor UO_1330 (O_1330,N_18589,N_18179);
xor UO_1331 (O_1331,N_16795,N_18174);
and UO_1332 (O_1332,N_19265,N_16496);
or UO_1333 (O_1333,N_16791,N_17220);
xor UO_1334 (O_1334,N_17642,N_16693);
and UO_1335 (O_1335,N_16152,N_17337);
or UO_1336 (O_1336,N_17406,N_16958);
or UO_1337 (O_1337,N_16244,N_17832);
or UO_1338 (O_1338,N_16527,N_17260);
nand UO_1339 (O_1339,N_18694,N_19396);
nand UO_1340 (O_1340,N_17914,N_18218);
xnor UO_1341 (O_1341,N_18611,N_19159);
xor UO_1342 (O_1342,N_17444,N_16154);
nand UO_1343 (O_1343,N_19990,N_16393);
xor UO_1344 (O_1344,N_17384,N_19417);
nand UO_1345 (O_1345,N_16542,N_16583);
xor UO_1346 (O_1346,N_19580,N_16002);
nand UO_1347 (O_1347,N_19796,N_17936);
and UO_1348 (O_1348,N_19076,N_17122);
and UO_1349 (O_1349,N_19524,N_18730);
or UO_1350 (O_1350,N_19457,N_19930);
or UO_1351 (O_1351,N_18030,N_16521);
xor UO_1352 (O_1352,N_18119,N_19579);
nor UO_1353 (O_1353,N_19610,N_17953);
xnor UO_1354 (O_1354,N_19441,N_16130);
xnor UO_1355 (O_1355,N_16831,N_18684);
nand UO_1356 (O_1356,N_18350,N_18929);
or UO_1357 (O_1357,N_19588,N_19055);
xnor UO_1358 (O_1358,N_16854,N_17922);
nand UO_1359 (O_1359,N_18677,N_16377);
or UO_1360 (O_1360,N_19433,N_18935);
nor UO_1361 (O_1361,N_19811,N_16255);
nand UO_1362 (O_1362,N_19215,N_17462);
and UO_1363 (O_1363,N_17287,N_19358);
nand UO_1364 (O_1364,N_17596,N_16114);
nor UO_1365 (O_1365,N_17825,N_17709);
xor UO_1366 (O_1366,N_17711,N_17697);
and UO_1367 (O_1367,N_17398,N_17064);
or UO_1368 (O_1368,N_18498,N_19847);
nor UO_1369 (O_1369,N_16434,N_18753);
and UO_1370 (O_1370,N_16787,N_19642);
and UO_1371 (O_1371,N_18676,N_19256);
and UO_1372 (O_1372,N_19617,N_17283);
or UO_1373 (O_1373,N_18535,N_19722);
xnor UO_1374 (O_1374,N_19375,N_16884);
nor UO_1375 (O_1375,N_17493,N_16504);
nor UO_1376 (O_1376,N_17105,N_19937);
xnor UO_1377 (O_1377,N_18883,N_18397);
or UO_1378 (O_1378,N_18782,N_16965);
or UO_1379 (O_1379,N_17124,N_16065);
or UO_1380 (O_1380,N_19096,N_17692);
xor UO_1381 (O_1381,N_19901,N_16248);
xor UO_1382 (O_1382,N_18657,N_17798);
or UO_1383 (O_1383,N_16037,N_19972);
nand UO_1384 (O_1384,N_17392,N_16307);
and UO_1385 (O_1385,N_17277,N_17125);
or UO_1386 (O_1386,N_16891,N_18053);
nor UO_1387 (O_1387,N_18783,N_18297);
or UO_1388 (O_1388,N_19100,N_19103);
nor UO_1389 (O_1389,N_18890,N_17244);
and UO_1390 (O_1390,N_19775,N_16340);
nor UO_1391 (O_1391,N_16102,N_18105);
xor UO_1392 (O_1392,N_18178,N_16829);
nor UO_1393 (O_1393,N_17866,N_19140);
nor UO_1394 (O_1394,N_17296,N_16333);
and UO_1395 (O_1395,N_16335,N_19919);
and UO_1396 (O_1396,N_19308,N_17961);
nand UO_1397 (O_1397,N_16926,N_18865);
or UO_1398 (O_1398,N_18349,N_17538);
xnor UO_1399 (O_1399,N_17365,N_18764);
nand UO_1400 (O_1400,N_19708,N_18526);
xnor UO_1401 (O_1401,N_16585,N_17581);
nor UO_1402 (O_1402,N_17465,N_16233);
nor UO_1403 (O_1403,N_19418,N_18678);
nor UO_1404 (O_1404,N_16937,N_17994);
xor UO_1405 (O_1405,N_17027,N_17058);
and UO_1406 (O_1406,N_17169,N_16474);
xnor UO_1407 (O_1407,N_18800,N_19163);
nor UO_1408 (O_1408,N_18515,N_17015);
xor UO_1409 (O_1409,N_19921,N_16678);
nand UO_1410 (O_1410,N_19962,N_17200);
xnor UO_1411 (O_1411,N_19351,N_18293);
and UO_1412 (O_1412,N_16372,N_18151);
xnor UO_1413 (O_1413,N_16809,N_19152);
nor UO_1414 (O_1414,N_18387,N_16486);
nand UO_1415 (O_1415,N_18255,N_19238);
nor UO_1416 (O_1416,N_16416,N_17524);
and UO_1417 (O_1417,N_19134,N_16517);
or UO_1418 (O_1418,N_17999,N_16980);
nor UO_1419 (O_1419,N_16701,N_18908);
or UO_1420 (O_1420,N_17954,N_18849);
or UO_1421 (O_1421,N_17749,N_18947);
nor UO_1422 (O_1422,N_16357,N_16280);
or UO_1423 (O_1423,N_19264,N_18048);
nand UO_1424 (O_1424,N_17261,N_16558);
nand UO_1425 (O_1425,N_18976,N_17201);
xnor UO_1426 (O_1426,N_18073,N_18029);
nor UO_1427 (O_1427,N_19220,N_18450);
nand UO_1428 (O_1428,N_17787,N_16985);
and UO_1429 (O_1429,N_16270,N_18620);
and UO_1430 (O_1430,N_18565,N_17445);
nand UO_1431 (O_1431,N_17980,N_17331);
nand UO_1432 (O_1432,N_19191,N_16258);
xor UO_1433 (O_1433,N_16422,N_16426);
or UO_1434 (O_1434,N_18419,N_19219);
nand UO_1435 (O_1435,N_19354,N_17344);
or UO_1436 (O_1436,N_17684,N_16706);
nand UO_1437 (O_1437,N_16262,N_18803);
xor UO_1438 (O_1438,N_17497,N_17706);
or UO_1439 (O_1439,N_17421,N_19000);
xor UO_1440 (O_1440,N_17827,N_19737);
nand UO_1441 (O_1441,N_18097,N_17663);
or UO_1442 (O_1442,N_16367,N_16164);
or UO_1443 (O_1443,N_16112,N_17145);
nor UO_1444 (O_1444,N_18913,N_19033);
xor UO_1445 (O_1445,N_19414,N_16513);
xor UO_1446 (O_1446,N_19562,N_18497);
nand UO_1447 (O_1447,N_19876,N_19671);
nor UO_1448 (O_1448,N_17179,N_18042);
nand UO_1449 (O_1449,N_17217,N_16702);
nand UO_1450 (O_1450,N_16612,N_16358);
nand UO_1451 (O_1451,N_16453,N_19156);
xnor UO_1452 (O_1452,N_16087,N_17032);
nor UO_1453 (O_1453,N_19739,N_18146);
xnor UO_1454 (O_1454,N_17492,N_19920);
nor UO_1455 (O_1455,N_17777,N_19214);
xor UO_1456 (O_1456,N_19735,N_17791);
nand UO_1457 (O_1457,N_18487,N_16730);
or UO_1458 (O_1458,N_17949,N_18937);
and UO_1459 (O_1459,N_18981,N_17376);
or UO_1460 (O_1460,N_17159,N_17778);
and UO_1461 (O_1461,N_16193,N_17412);
xnor UO_1462 (O_1462,N_17119,N_16593);
nand UO_1463 (O_1463,N_18699,N_19030);
or UO_1464 (O_1464,N_19180,N_16430);
xor UO_1465 (O_1465,N_18921,N_17234);
xnor UO_1466 (O_1466,N_17007,N_17107);
nand UO_1467 (O_1467,N_18686,N_16599);
nand UO_1468 (O_1468,N_18973,N_19687);
xnor UO_1469 (O_1469,N_18300,N_16281);
xnor UO_1470 (O_1470,N_19335,N_18209);
nand UO_1471 (O_1471,N_17104,N_19973);
nor UO_1472 (O_1472,N_18584,N_17195);
xnor UO_1473 (O_1473,N_18761,N_17397);
xor UO_1474 (O_1474,N_18422,N_17864);
nand UO_1475 (O_1475,N_16932,N_19670);
nand UO_1476 (O_1476,N_19272,N_19865);
or UO_1477 (O_1477,N_19321,N_18689);
nand UO_1478 (O_1478,N_18878,N_18955);
xor UO_1479 (O_1479,N_18705,N_19176);
xnor UO_1480 (O_1480,N_17063,N_16400);
nor UO_1481 (O_1481,N_16161,N_17116);
nand UO_1482 (O_1482,N_19507,N_16970);
nand UO_1483 (O_1483,N_16165,N_17704);
xor UO_1484 (O_1484,N_18110,N_17356);
nand UO_1485 (O_1485,N_16454,N_17537);
xor UO_1486 (O_1486,N_16581,N_16942);
nand UO_1487 (O_1487,N_18509,N_18075);
or UO_1488 (O_1488,N_19826,N_18299);
nand UO_1489 (O_1489,N_16774,N_17675);
and UO_1490 (O_1490,N_17312,N_16495);
xnor UO_1491 (O_1491,N_16811,N_18772);
nand UO_1492 (O_1492,N_17017,N_17024);
nor UO_1493 (O_1493,N_18975,N_18155);
or UO_1494 (O_1494,N_17305,N_18645);
xnor UO_1495 (O_1495,N_17782,N_17818);
nor UO_1496 (O_1496,N_16943,N_18909);
and UO_1497 (O_1497,N_18197,N_19161);
or UO_1498 (O_1498,N_19476,N_19960);
and UO_1499 (O_1499,N_18045,N_19229);
nor UO_1500 (O_1500,N_17690,N_19693);
xnor UO_1501 (O_1501,N_16584,N_17986);
and UO_1502 (O_1502,N_17081,N_17845);
nor UO_1503 (O_1503,N_16902,N_16343);
and UO_1504 (O_1504,N_17515,N_18243);
and UO_1505 (O_1505,N_16552,N_16413);
or UO_1506 (O_1506,N_19289,N_19720);
and UO_1507 (O_1507,N_18011,N_18231);
nand UO_1508 (O_1508,N_17224,N_16319);
or UO_1509 (O_1509,N_18747,N_19306);
xor UO_1510 (O_1510,N_17503,N_17060);
xnor UO_1511 (O_1511,N_18924,N_17590);
nand UO_1512 (O_1512,N_19802,N_16895);
or UO_1513 (O_1513,N_17012,N_19885);
and UO_1514 (O_1514,N_16188,N_17858);
or UO_1515 (O_1515,N_16622,N_17473);
nor UO_1516 (O_1516,N_19041,N_17728);
nor UO_1517 (O_1517,N_19949,N_19090);
and UO_1518 (O_1518,N_18579,N_16292);
and UO_1519 (O_1519,N_18158,N_17152);
nand UO_1520 (O_1520,N_19880,N_16219);
and UO_1521 (O_1521,N_17669,N_16222);
and UO_1522 (O_1522,N_18080,N_18490);
nand UO_1523 (O_1523,N_17390,N_18825);
or UO_1524 (O_1524,N_19556,N_17016);
xnor UO_1525 (O_1525,N_19299,N_19898);
nand UO_1526 (O_1526,N_16726,N_18642);
xnor UO_1527 (O_1527,N_18177,N_18331);
and UO_1528 (O_1528,N_18414,N_18571);
xnor UO_1529 (O_1529,N_16740,N_16099);
nand UO_1530 (O_1530,N_17819,N_16961);
nand UO_1531 (O_1531,N_17880,N_16639);
or UO_1532 (O_1532,N_19935,N_16457);
or UO_1533 (O_1533,N_16150,N_16182);
nor UO_1534 (O_1534,N_19162,N_17066);
nor UO_1535 (O_1535,N_17442,N_16691);
or UO_1536 (O_1536,N_19601,N_16282);
nor UO_1537 (O_1537,N_19849,N_19121);
and UO_1538 (O_1538,N_16284,N_19840);
xor UO_1539 (O_1539,N_16836,N_18555);
and UO_1540 (O_1540,N_18723,N_16712);
nand UO_1541 (O_1541,N_17920,N_16914);
nand UO_1542 (O_1542,N_17168,N_17535);
and UO_1543 (O_1543,N_19965,N_17351);
nand UO_1544 (O_1544,N_19106,N_18672);
nor UO_1545 (O_1545,N_17223,N_16386);
or UO_1546 (O_1546,N_19661,N_17155);
xor UO_1547 (O_1547,N_17577,N_18484);
or UO_1548 (O_1548,N_19702,N_19035);
and UO_1549 (O_1549,N_16572,N_18400);
xnor UO_1550 (O_1550,N_18494,N_18756);
nor UO_1551 (O_1551,N_19449,N_18500);
nand UO_1552 (O_1552,N_17995,N_18709);
or UO_1553 (O_1553,N_18629,N_19300);
and UO_1554 (O_1554,N_18873,N_16168);
and UO_1555 (O_1555,N_16395,N_16290);
and UO_1556 (O_1556,N_19618,N_18960);
or UO_1557 (O_1557,N_16352,N_19697);
xnor UO_1558 (O_1558,N_16320,N_16808);
xnor UO_1559 (O_1559,N_18725,N_16621);
and UO_1560 (O_1560,N_16921,N_19810);
or UO_1561 (O_1561,N_18335,N_18369);
nor UO_1562 (O_1562,N_18874,N_18165);
nor UO_1563 (O_1563,N_19303,N_18010);
or UO_1564 (O_1564,N_18374,N_18916);
xor UO_1565 (O_1565,N_19494,N_19340);
and UO_1566 (O_1566,N_18945,N_18056);
or UO_1567 (O_1567,N_17448,N_17617);
nor UO_1568 (O_1568,N_19189,N_16538);
and UO_1569 (O_1569,N_17622,N_19145);
xnor UO_1570 (O_1570,N_18149,N_16887);
nor UO_1571 (O_1571,N_16095,N_17014);
nand UO_1572 (O_1572,N_16247,N_16752);
and UO_1573 (O_1573,N_19252,N_16186);
nor UO_1574 (O_1574,N_19536,N_19292);
nor UO_1575 (O_1575,N_19863,N_16204);
nor UO_1576 (O_1576,N_16947,N_18928);
xor UO_1577 (O_1577,N_19769,N_16399);
xor UO_1578 (O_1578,N_16111,N_18485);
and UO_1579 (O_1579,N_16757,N_17208);
or UO_1580 (O_1580,N_18719,N_18021);
nor UO_1581 (O_1581,N_16274,N_19590);
nand UO_1582 (O_1582,N_19357,N_17139);
nand UO_1583 (O_1583,N_16216,N_16971);
nor UO_1584 (O_1584,N_19540,N_17151);
or UO_1585 (O_1585,N_16982,N_19594);
and UO_1586 (O_1586,N_19542,N_19821);
nand UO_1587 (O_1587,N_18740,N_16886);
nand UO_1588 (O_1588,N_19908,N_16076);
xor UO_1589 (O_1589,N_18236,N_19329);
and UO_1590 (O_1590,N_18503,N_17388);
xor UO_1591 (O_1591,N_16515,N_19639);
and UO_1592 (O_1592,N_17487,N_18659);
or UO_1593 (O_1593,N_19701,N_17627);
nor UO_1594 (O_1594,N_17318,N_18263);
and UO_1595 (O_1595,N_16959,N_18259);
and UO_1596 (O_1596,N_18831,N_17662);
xnor UO_1597 (O_1597,N_17664,N_19952);
nor UO_1598 (O_1598,N_16912,N_19569);
or UO_1599 (O_1599,N_16414,N_19887);
nand UO_1600 (O_1600,N_16098,N_18407);
xor UO_1601 (O_1601,N_16885,N_18706);
or UO_1602 (O_1602,N_19886,N_16449);
nand UO_1603 (O_1603,N_16551,N_19324);
and UO_1604 (O_1604,N_16220,N_16081);
xnor UO_1605 (O_1605,N_16670,N_17381);
nand UO_1606 (O_1606,N_16727,N_19782);
nand UO_1607 (O_1607,N_16602,N_16073);
xor UO_1608 (O_1608,N_17325,N_19691);
nand UO_1609 (O_1609,N_17702,N_19302);
nand UO_1610 (O_1610,N_18850,N_18405);
nand UO_1611 (O_1611,N_16238,N_17443);
nand UO_1612 (O_1612,N_16456,N_19614);
nand UO_1613 (O_1613,N_19467,N_19493);
and UO_1614 (O_1614,N_18626,N_18778);
nor UO_1615 (O_1615,N_19572,N_16796);
xnor UO_1616 (O_1616,N_17698,N_17896);
nand UO_1617 (O_1617,N_17410,N_18880);
nor UO_1618 (O_1618,N_19196,N_18992);
nor UO_1619 (O_1619,N_18111,N_17170);
nor UO_1620 (O_1620,N_17790,N_17516);
xnor UO_1621 (O_1621,N_17019,N_18267);
or UO_1622 (O_1622,N_18636,N_16063);
and UO_1623 (O_1623,N_17192,N_18911);
nor UO_1624 (O_1624,N_19187,N_18965);
or UO_1625 (O_1625,N_18309,N_16589);
or UO_1626 (O_1626,N_19053,N_18893);
nand UO_1627 (O_1627,N_17640,N_16034);
or UO_1628 (O_1628,N_18828,N_18205);
or UO_1629 (O_1629,N_16847,N_19539);
and UO_1630 (O_1630,N_17946,N_16928);
and UO_1631 (O_1631,N_17668,N_17290);
and UO_1632 (O_1632,N_18168,N_16201);
or UO_1633 (O_1633,N_16744,N_16104);
nand UO_1634 (O_1634,N_19692,N_17925);
nand UO_1635 (O_1635,N_18224,N_18169);
xor UO_1636 (O_1636,N_18332,N_16156);
or UO_1637 (O_1637,N_17157,N_19497);
and UO_1638 (O_1638,N_19561,N_17180);
nor UO_1639 (O_1639,N_17504,N_17940);
nor UO_1640 (O_1640,N_17072,N_19987);
nand UO_1641 (O_1641,N_16825,N_19226);
nand UO_1642 (O_1642,N_19114,N_19841);
xor UO_1643 (O_1643,N_17788,N_18336);
or UO_1644 (O_1644,N_18408,N_19127);
nand UO_1645 (O_1645,N_16473,N_19205);
nand UO_1646 (O_1646,N_17338,N_18462);
xnor UO_1647 (O_1647,N_19088,N_18195);
nor UO_1648 (O_1648,N_16697,N_19016);
or UO_1649 (O_1649,N_16981,N_16013);
or UO_1650 (O_1650,N_19454,N_16641);
nor UO_1651 (O_1651,N_19888,N_16021);
xnor UO_1652 (O_1652,N_16790,N_16234);
nand UO_1653 (O_1653,N_17532,N_18972);
xnor UO_1654 (O_1654,N_17043,N_18856);
and UO_1655 (O_1655,N_17730,N_19656);
nand UO_1656 (O_1656,N_17931,N_16509);
xnor UO_1657 (O_1657,N_16855,N_19271);
or UO_1658 (O_1658,N_19063,N_17205);
nand UO_1659 (O_1659,N_19178,N_17000);
nand UO_1660 (O_1660,N_19586,N_17306);
xnor UO_1661 (O_1661,N_18631,N_18219);
xnor UO_1662 (O_1662,N_17955,N_18176);
nor UO_1663 (O_1663,N_18795,N_18418);
or UO_1664 (O_1664,N_17235,N_18084);
nand UO_1665 (O_1665,N_17740,N_19529);
and UO_1666 (O_1666,N_17768,N_19551);
and UO_1667 (O_1667,N_16684,N_17364);
xnor UO_1668 (O_1668,N_19563,N_18698);
or UO_1669 (O_1669,N_17321,N_17470);
or UO_1670 (O_1670,N_19791,N_16008);
nand UO_1671 (O_1671,N_17612,N_19747);
nor UO_1672 (O_1672,N_17114,N_17758);
xnor UO_1673 (O_1673,N_18377,N_19870);
xnor UO_1674 (O_1674,N_17008,N_17264);
nor UO_1675 (O_1675,N_16858,N_17708);
and UO_1676 (O_1676,N_19015,N_16604);
or UO_1677 (O_1677,N_19223,N_19194);
nor UO_1678 (O_1678,N_19557,N_19862);
nor UO_1679 (O_1679,N_18564,N_19762);
or UO_1680 (O_1680,N_19305,N_16661);
or UO_1681 (O_1681,N_16469,N_18347);
and UO_1682 (O_1682,N_19925,N_17633);
nor UO_1683 (O_1683,N_19244,N_19043);
or UO_1684 (O_1684,N_18674,N_16556);
and UO_1685 (O_1685,N_19609,N_18544);
and UO_1686 (O_1686,N_19038,N_19461);
and UO_1687 (O_1687,N_19992,N_17402);
nor UO_1688 (O_1688,N_18104,N_16458);
xnor UO_1689 (O_1689,N_19552,N_16586);
and UO_1690 (O_1690,N_16108,N_17441);
and UO_1691 (O_1691,N_16775,N_17807);
nand UO_1692 (O_1692,N_18248,N_18223);
or UO_1693 (O_1693,N_18639,N_18278);
and UO_1694 (O_1694,N_19520,N_17457);
nor UO_1695 (O_1695,N_16771,N_19573);
nor UO_1696 (O_1696,N_19017,N_19165);
or UO_1697 (O_1697,N_18198,N_16562);
or UO_1698 (O_1698,N_18354,N_18361);
nor UO_1699 (O_1699,N_19144,N_19641);
and UO_1700 (O_1700,N_16754,N_16452);
xor UO_1701 (O_1701,N_16476,N_19014);
and UO_1702 (O_1702,N_16997,N_16846);
nand UO_1703 (O_1703,N_16929,N_17847);
and UO_1704 (O_1704,N_18370,N_16043);
or UO_1705 (O_1705,N_16184,N_17511);
nand UO_1706 (O_1706,N_19360,N_17650);
or UO_1707 (O_1707,N_16905,N_19261);
or UO_1708 (O_1708,N_19253,N_18072);
nor UO_1709 (O_1709,N_16715,N_18436);
nor UO_1710 (O_1710,N_18881,N_16173);
nand UO_1711 (O_1711,N_19350,N_17144);
or UO_1712 (O_1712,N_19437,N_17034);
nand UO_1713 (O_1713,N_18832,N_18539);
or UO_1714 (O_1714,N_19415,N_18398);
xor UO_1715 (O_1715,N_18421,N_16557);
or UO_1716 (O_1716,N_17437,N_19853);
xor UO_1717 (O_1717,N_16502,N_19940);
or UO_1718 (O_1718,N_18541,N_16046);
nor UO_1719 (O_1719,N_17797,N_18529);
or UO_1720 (O_1720,N_16533,N_19326);
and UO_1721 (O_1721,N_16832,N_18601);
xor UO_1722 (O_1722,N_19977,N_16339);
nor UO_1723 (O_1723,N_16329,N_18381);
nand UO_1724 (O_1724,N_18785,N_18822);
or UO_1725 (O_1725,N_17315,N_17154);
and UO_1726 (O_1726,N_16306,N_17049);
nor UO_1727 (O_1727,N_17118,N_18194);
xnor UO_1728 (O_1728,N_18438,N_18521);
and UO_1729 (O_1729,N_17609,N_17071);
nand UO_1730 (O_1730,N_19370,N_16017);
or UO_1731 (O_1731,N_18614,N_16756);
and UO_1732 (O_1732,N_17194,N_18453);
or UO_1733 (O_1733,N_16070,N_17282);
and UO_1734 (O_1734,N_19518,N_18950);
nor UO_1735 (O_1735,N_17251,N_18022);
or UO_1736 (O_1736,N_16879,N_19931);
and UO_1737 (O_1737,N_16135,N_18562);
nand UO_1738 (O_1738,N_19564,N_17710);
nand UO_1739 (O_1739,N_16698,N_18035);
and UO_1740 (O_1740,N_16777,N_19909);
xor UO_1741 (O_1741,N_18120,N_16856);
nor UO_1742 (O_1742,N_16256,N_16239);
nor UO_1743 (O_1743,N_16235,N_17506);
and UO_1744 (O_1744,N_19985,N_18003);
or UO_1745 (O_1745,N_19085,N_17654);
nor UO_1746 (O_1746,N_18750,N_19317);
xor UO_1747 (O_1747,N_16291,N_18608);
nor UO_1748 (O_1748,N_16019,N_17656);
or UO_1749 (O_1749,N_17699,N_16688);
nand UO_1750 (O_1750,N_19333,N_17101);
nor UO_1751 (O_1751,N_19447,N_16625);
or UO_1752 (O_1752,N_17526,N_18649);
nand UO_1753 (O_1753,N_16637,N_16704);
and UO_1754 (O_1754,N_19013,N_17580);
xnor UO_1755 (O_1755,N_17693,N_16488);
or UO_1756 (O_1756,N_16628,N_16342);
xor UO_1757 (O_1757,N_18334,N_19371);
nand UO_1758 (O_1758,N_18721,N_16055);
or UO_1759 (O_1759,N_19429,N_19659);
or UO_1760 (O_1760,N_16206,N_17430);
nor UO_1761 (O_1761,N_17569,N_18472);
nor UO_1762 (O_1762,N_19785,N_16577);
nand UO_1763 (O_1763,N_19362,N_19755);
xor UO_1764 (O_1764,N_16273,N_16269);
nor UO_1765 (O_1765,N_18869,N_19347);
nor UO_1766 (O_1766,N_17494,N_16477);
nor UO_1767 (O_1767,N_18261,N_16363);
xnor UO_1768 (O_1768,N_19186,N_18055);
nor UO_1769 (O_1769,N_19606,N_19332);
nand UO_1770 (O_1770,N_18085,N_17326);
and UO_1771 (O_1771,N_16629,N_19280);
and UO_1772 (O_1772,N_16051,N_17838);
and UO_1773 (O_1773,N_19064,N_19591);
xor UO_1774 (O_1774,N_17604,N_18997);
and UO_1775 (O_1775,N_16249,N_17218);
nor UO_1776 (O_1776,N_19895,N_18312);
nand UO_1777 (O_1777,N_16133,N_19002);
xor UO_1778 (O_1778,N_19135,N_16341);
or UO_1779 (O_1779,N_16814,N_17174);
nand UO_1780 (O_1780,N_19986,N_18225);
or UO_1781 (O_1781,N_18340,N_19344);
nand UO_1782 (O_1782,N_19603,N_18858);
nand UO_1783 (O_1783,N_16402,N_19394);
nand UO_1784 (O_1784,N_17903,N_18426);
nand UO_1785 (O_1785,N_16632,N_17618);
xnor UO_1786 (O_1786,N_16162,N_16461);
nor UO_1787 (O_1787,N_18093,N_17113);
or UO_1788 (O_1788,N_16741,N_19363);
or UO_1789 (O_1789,N_18647,N_18567);
and UO_1790 (O_1790,N_17840,N_19516);
nor UO_1791 (O_1791,N_17761,N_16908);
or UO_1792 (O_1792,N_19668,N_19320);
or UO_1793 (O_1793,N_19008,N_17909);
xnor UO_1794 (O_1794,N_16563,N_16931);
and UO_1795 (O_1795,N_17353,N_18765);
nand UO_1796 (O_1796,N_16110,N_19622);
and UO_1797 (O_1797,N_17793,N_17977);
and UO_1798 (O_1798,N_17404,N_16232);
xor UO_1799 (O_1799,N_19889,N_16464);
and UO_1800 (O_1800,N_18578,N_19731);
and UO_1801 (O_1801,N_16278,N_19652);
or UO_1802 (O_1802,N_17960,N_16996);
nor UO_1803 (O_1803,N_16801,N_18615);
nor UO_1804 (O_1804,N_17108,N_16078);
nor UO_1805 (O_1805,N_19007,N_16758);
and UO_1806 (O_1806,N_18513,N_19061);
nand UO_1807 (O_1807,N_17030,N_16594);
or UO_1808 (O_1808,N_17814,N_19575);
and UO_1809 (O_1809,N_19481,N_18956);
nand UO_1810 (O_1810,N_17438,N_19576);
nand UO_1811 (O_1811,N_18326,N_17267);
xnor UO_1812 (O_1812,N_16015,N_17456);
or UO_1813 (O_1813,N_18007,N_17253);
and UO_1814 (O_1814,N_18087,N_18640);
and UO_1815 (O_1815,N_16029,N_17090);
xor UO_1816 (O_1816,N_18404,N_17281);
nand UO_1817 (O_1817,N_16194,N_19938);
nor UO_1818 (O_1818,N_17003,N_18260);
xnor UO_1819 (O_1819,N_18923,N_19262);
xor UO_1820 (O_1820,N_18166,N_19192);
xor UO_1821 (O_1821,N_19966,N_16045);
xor UO_1822 (O_1822,N_19532,N_16084);
nor UO_1823 (O_1823,N_19040,N_17628);
xor UO_1824 (O_1824,N_19824,N_16812);
or UO_1825 (O_1825,N_17183,N_16838);
xnor UO_1826 (O_1826,N_16881,N_18696);
or UO_1827 (O_1827,N_16304,N_17405);
and UO_1828 (O_1828,N_17429,N_18082);
or UO_1829 (O_1829,N_19204,N_19953);
nand UO_1830 (O_1830,N_16225,N_18545);
and UO_1831 (O_1831,N_17236,N_18532);
nor UO_1832 (O_1832,N_19343,N_19589);
nor UO_1833 (O_1833,N_16992,N_19784);
nor UO_1834 (O_1834,N_19651,N_18094);
or UO_1835 (O_1835,N_18582,N_18113);
and UO_1836 (O_1836,N_16039,N_18758);
xor UO_1837 (O_1837,N_19713,N_17839);
and UO_1838 (O_1838,N_18375,N_18059);
xor UO_1839 (O_1839,N_19560,N_18933);
or UO_1840 (O_1840,N_17878,N_17394);
nor UO_1841 (O_1841,N_18507,N_17886);
nand UO_1842 (O_1842,N_18305,N_19932);
and UO_1843 (O_1843,N_17534,N_19224);
xnor UO_1844 (O_1844,N_19861,N_19381);
nor UO_1845 (O_1845,N_16359,N_18993);
or UO_1846 (O_1846,N_18233,N_16665);
nor UO_1847 (O_1847,N_17718,N_19528);
nor UO_1848 (O_1848,N_17585,N_17191);
xnor UO_1849 (O_1849,N_16627,N_16673);
nand UO_1850 (O_1850,N_18493,N_17447);
or UO_1851 (O_1851,N_17978,N_19074);
or UO_1852 (O_1852,N_17300,N_16326);
or UO_1853 (O_1853,N_17987,N_18704);
and UO_1854 (O_1854,N_18989,N_19605);
xnor UO_1855 (O_1855,N_17222,N_17358);
and UO_1856 (O_1856,N_18108,N_17499);
xor UO_1857 (O_1857,N_19296,N_17910);
or UO_1858 (O_1858,N_16523,N_19182);
nand UO_1859 (O_1859,N_16117,N_19431);
xnor UO_1860 (O_1860,N_17269,N_17841);
nor UO_1861 (O_1861,N_18076,N_18735);
nand UO_1862 (O_1862,N_19183,N_19342);
nand UO_1863 (O_1863,N_19216,N_16772);
xnor UO_1864 (O_1864,N_17597,N_17167);
nor UO_1865 (O_1865,N_18995,N_16689);
xnor UO_1866 (O_1866,N_19860,N_16735);
or UO_1867 (O_1867,N_17563,N_18286);
nor UO_1868 (O_1868,N_16378,N_19478);
nand UO_1869 (O_1869,N_16153,N_18970);
nor UO_1870 (O_1870,N_19446,N_16708);
nor UO_1871 (O_1871,N_19750,N_16951);
and UO_1872 (O_1872,N_18622,N_19970);
xor UO_1873 (O_1873,N_18573,N_18471);
xnor UO_1874 (O_1874,N_17556,N_18425);
nand UO_1875 (O_1875,N_18860,N_16680);
nand UO_1876 (O_1876,N_18276,N_17641);
or UO_1877 (O_1877,N_17474,N_18257);
nand UO_1878 (O_1878,N_19760,N_17423);
and UO_1879 (O_1879,N_18186,N_18817);
and UO_1880 (O_1880,N_17148,N_19126);
xnor UO_1881 (O_1881,N_19857,N_17649);
and UO_1882 (O_1882,N_19133,N_18489);
or UO_1883 (O_1883,N_18774,N_17905);
or UO_1884 (O_1884,N_17988,N_17748);
xor UO_1885 (O_1885,N_16493,N_19698);
or UO_1886 (O_1886,N_19503,N_19430);
or UO_1887 (O_1887,N_17133,N_19964);
nand UO_1888 (O_1888,N_19500,N_17449);
or UO_1889 (O_1889,N_18969,N_18373);
and UO_1890 (O_1890,N_16183,N_17862);
and UO_1891 (O_1891,N_17742,N_16834);
and UO_1892 (O_1892,N_17982,N_19171);
and UO_1893 (O_1893,N_16853,N_16874);
and UO_1894 (O_1894,N_16769,N_17446);
nor UO_1895 (O_1895,N_18538,N_19059);
xor UO_1896 (O_1896,N_19604,N_16973);
xor UO_1897 (O_1897,N_19819,N_18469);
and UO_1898 (O_1898,N_18561,N_16788);
nor UO_1899 (O_1899,N_19034,N_18321);
and UO_1900 (O_1900,N_18518,N_17608);
nor UO_1901 (O_1901,N_17964,N_18940);
xor UO_1902 (O_1902,N_17567,N_17450);
nand UO_1903 (O_1903,N_19759,N_16721);
nand UO_1904 (O_1904,N_19615,N_16636);
xor UO_1905 (O_1905,N_19679,N_19323);
nand UO_1906 (O_1906,N_18125,N_19534);
or UO_1907 (O_1907,N_19646,N_18359);
and UO_1908 (O_1908,N_16375,N_18451);
or UO_1909 (O_1909,N_18079,N_19117);
nor UO_1910 (O_1910,N_18953,N_19093);
xor UO_1911 (O_1911,N_19473,N_17324);
nor UO_1912 (O_1912,N_17893,N_16871);
or UO_1913 (O_1913,N_18692,N_16904);
xor UO_1914 (O_1914,N_17996,N_17972);
xor UO_1915 (O_1915,N_16546,N_18552);
or UO_1916 (O_1916,N_16042,N_19044);
xor UO_1917 (O_1917,N_18283,N_18445);
or UO_1918 (O_1918,N_19440,N_19827);
or UO_1919 (O_1919,N_17129,N_16106);
nor UO_1920 (O_1920,N_19685,N_16196);
nor UO_1921 (O_1921,N_17770,N_19917);
and UO_1922 (O_1922,N_18141,N_18821);
or UO_1923 (O_1923,N_17399,N_18352);
or UO_1924 (O_1924,N_19246,N_18154);
nand UO_1925 (O_1925,N_17379,N_17011);
nor UO_1926 (O_1926,N_19650,N_18499);
and UO_1927 (O_1927,N_16818,N_16539);
xnor UO_1928 (O_1928,N_19352,N_19776);
and UO_1929 (O_1929,N_18252,N_19912);
nor UO_1930 (O_1930,N_19578,N_17240);
and UO_1931 (O_1931,N_16935,N_18131);
nor UO_1932 (O_1932,N_17009,N_18439);
nor UO_1933 (O_1933,N_18291,N_18180);
nand UO_1934 (O_1934,N_18069,N_18653);
nand UO_1935 (O_1935,N_17751,N_17696);
nand UO_1936 (O_1936,N_19946,N_19913);
nor UO_1937 (O_1937,N_18447,N_16346);
or UO_1938 (O_1938,N_16361,N_19124);
or UO_1939 (O_1939,N_18854,N_19637);
and UO_1940 (O_1940,N_17163,N_18625);
or UO_1941 (O_1941,N_18159,N_18288);
nor UO_1942 (O_1942,N_19410,N_17636);
nor UO_1943 (O_1943,N_18156,N_18688);
nor UO_1944 (O_1944,N_19974,N_19662);
xor UO_1945 (O_1945,N_18308,N_18939);
and UO_1946 (O_1946,N_17550,N_19268);
nand UO_1947 (O_1947,N_18527,N_16883);
and UO_1948 (O_1948,N_16544,N_16663);
and UO_1949 (O_1949,N_17239,N_19995);
nand UO_1950 (O_1950,N_16468,N_18769);
nand UO_1951 (O_1951,N_16376,N_19761);
and UO_1952 (O_1952,N_17611,N_17918);
xor UO_1953 (O_1953,N_18690,N_19435);
xnor UO_1954 (O_1954,N_16328,N_17877);
nor UO_1955 (O_1955,N_16490,N_17796);
nand UO_1956 (O_1956,N_19553,N_18957);
and UO_1957 (O_1957,N_18481,N_17087);
nand UO_1958 (O_1958,N_18520,N_17372);
or UO_1959 (O_1959,N_18103,N_18379);
and UO_1960 (O_1960,N_17614,N_19523);
and UO_1961 (O_1961,N_19818,N_19098);
nand UO_1962 (O_1962,N_17606,N_19387);
nor UO_1963 (O_1963,N_19260,N_17746);
nand UO_1964 (O_1964,N_19259,N_19181);
and UO_1965 (O_1965,N_17755,N_17286);
nand UO_1966 (O_1966,N_18736,N_19567);
or UO_1967 (O_1967,N_19878,N_18051);
nand UO_1968 (O_1968,N_16016,N_19914);
and UO_1969 (O_1969,N_19330,N_16137);
or UO_1970 (O_1970,N_16316,N_16113);
xor UO_1971 (O_1971,N_17121,N_16006);
xor UO_1972 (O_1972,N_17173,N_17275);
xor UO_1973 (O_1973,N_17671,N_16710);
nand UO_1974 (O_1974,N_18181,N_18633);
nor UO_1975 (O_1975,N_19376,N_18281);
nor UO_1976 (O_1976,N_19744,N_18877);
nor UO_1977 (O_1977,N_16870,N_16507);
xnor UO_1978 (O_1978,N_16142,N_18216);
and UO_1979 (O_1979,N_17037,N_18440);
xnor UO_1980 (O_1980,N_16917,N_17288);
and UO_1981 (O_1981,N_18277,N_17734);
or UO_1982 (O_1982,N_19632,N_19003);
nor UO_1983 (O_1983,N_17362,N_19086);
nor UO_1984 (O_1984,N_19240,N_17897);
nor UO_1985 (O_1985,N_17828,N_16927);
nor UO_1986 (O_1986,N_16433,N_18173);
nand UO_1987 (O_1987,N_19596,N_17272);
xnor UO_1988 (O_1988,N_16387,N_17255);
or UO_1989 (O_1989,N_19817,N_16653);
xnor UO_1990 (O_1990,N_16570,N_16601);
nand UO_1991 (O_1991,N_17558,N_19929);
xor UO_1992 (O_1992,N_19984,N_16977);
nor UO_1993 (O_1993,N_19793,N_17975);
nand UO_1994 (O_1994,N_18635,N_17432);
and UO_1995 (O_1995,N_17128,N_17134);
nor UO_1996 (O_1996,N_17666,N_19675);
nand UO_1997 (O_1997,N_17231,N_18907);
xor UO_1998 (O_1998,N_17632,N_19283);
nand UO_1999 (O_1999,N_19918,N_19485);
xor UO_2000 (O_2000,N_18881,N_19922);
xnor UO_2001 (O_2001,N_19221,N_17870);
xor UO_2002 (O_2002,N_18038,N_16029);
xnor UO_2003 (O_2003,N_18082,N_16330);
and UO_2004 (O_2004,N_17489,N_19260);
or UO_2005 (O_2005,N_18328,N_18911);
nand UO_2006 (O_2006,N_17777,N_19334);
xnor UO_2007 (O_2007,N_17772,N_19289);
and UO_2008 (O_2008,N_16720,N_19064);
nand UO_2009 (O_2009,N_18125,N_17652);
nand UO_2010 (O_2010,N_18528,N_17679);
xnor UO_2011 (O_2011,N_18046,N_18729);
xor UO_2012 (O_2012,N_16382,N_19875);
nor UO_2013 (O_2013,N_16603,N_17972);
or UO_2014 (O_2014,N_17237,N_19898);
and UO_2015 (O_2015,N_19442,N_19740);
nand UO_2016 (O_2016,N_18638,N_18965);
and UO_2017 (O_2017,N_17031,N_17839);
nor UO_2018 (O_2018,N_16435,N_17835);
or UO_2019 (O_2019,N_16757,N_17108);
and UO_2020 (O_2020,N_17717,N_16275);
nand UO_2021 (O_2021,N_18491,N_19946);
nor UO_2022 (O_2022,N_17685,N_16720);
nor UO_2023 (O_2023,N_19243,N_17032);
xor UO_2024 (O_2024,N_19832,N_16554);
nand UO_2025 (O_2025,N_18236,N_17269);
and UO_2026 (O_2026,N_16452,N_19580);
nand UO_2027 (O_2027,N_18030,N_19445);
nand UO_2028 (O_2028,N_17064,N_17351);
nand UO_2029 (O_2029,N_18597,N_17645);
xor UO_2030 (O_2030,N_19737,N_19646);
xnor UO_2031 (O_2031,N_16398,N_19700);
and UO_2032 (O_2032,N_18903,N_17933);
xor UO_2033 (O_2033,N_16411,N_18261);
and UO_2034 (O_2034,N_17262,N_17163);
and UO_2035 (O_2035,N_17511,N_17514);
or UO_2036 (O_2036,N_16931,N_17902);
xnor UO_2037 (O_2037,N_17919,N_18707);
xnor UO_2038 (O_2038,N_18898,N_16427);
and UO_2039 (O_2039,N_19817,N_18494);
or UO_2040 (O_2040,N_16000,N_16352);
or UO_2041 (O_2041,N_18391,N_17789);
or UO_2042 (O_2042,N_16665,N_18620);
nor UO_2043 (O_2043,N_17185,N_17549);
and UO_2044 (O_2044,N_19380,N_18223);
xnor UO_2045 (O_2045,N_16397,N_18710);
xnor UO_2046 (O_2046,N_19952,N_19111);
xnor UO_2047 (O_2047,N_19466,N_17654);
or UO_2048 (O_2048,N_19051,N_19087);
and UO_2049 (O_2049,N_16328,N_16893);
and UO_2050 (O_2050,N_17136,N_18976);
xor UO_2051 (O_2051,N_19456,N_18438);
nor UO_2052 (O_2052,N_18258,N_16601);
and UO_2053 (O_2053,N_16462,N_16021);
nor UO_2054 (O_2054,N_18515,N_16345);
or UO_2055 (O_2055,N_16985,N_17557);
and UO_2056 (O_2056,N_17505,N_18043);
xor UO_2057 (O_2057,N_16477,N_19433);
or UO_2058 (O_2058,N_19551,N_18795);
xnor UO_2059 (O_2059,N_18578,N_18748);
or UO_2060 (O_2060,N_18257,N_17675);
and UO_2061 (O_2061,N_18954,N_18114);
or UO_2062 (O_2062,N_17663,N_16498);
xor UO_2063 (O_2063,N_17806,N_18726);
and UO_2064 (O_2064,N_19251,N_18922);
nor UO_2065 (O_2065,N_17040,N_17992);
xor UO_2066 (O_2066,N_16670,N_16676);
or UO_2067 (O_2067,N_18459,N_18805);
nor UO_2068 (O_2068,N_17255,N_18927);
and UO_2069 (O_2069,N_19234,N_18155);
xnor UO_2070 (O_2070,N_17172,N_18125);
or UO_2071 (O_2071,N_17896,N_17891);
nand UO_2072 (O_2072,N_16312,N_16130);
nor UO_2073 (O_2073,N_17015,N_18342);
nand UO_2074 (O_2074,N_18251,N_19895);
and UO_2075 (O_2075,N_17433,N_18446);
xor UO_2076 (O_2076,N_19255,N_19192);
nand UO_2077 (O_2077,N_18998,N_18552);
and UO_2078 (O_2078,N_19817,N_19487);
nand UO_2079 (O_2079,N_19497,N_19272);
or UO_2080 (O_2080,N_16807,N_18543);
xnor UO_2081 (O_2081,N_19872,N_18950);
nor UO_2082 (O_2082,N_19604,N_19605);
nand UO_2083 (O_2083,N_17966,N_17627);
xor UO_2084 (O_2084,N_16714,N_17354);
and UO_2085 (O_2085,N_16798,N_17652);
or UO_2086 (O_2086,N_16108,N_16048);
or UO_2087 (O_2087,N_17097,N_17691);
xnor UO_2088 (O_2088,N_18282,N_17129);
nand UO_2089 (O_2089,N_18942,N_18238);
or UO_2090 (O_2090,N_17313,N_18692);
or UO_2091 (O_2091,N_18828,N_19437);
nor UO_2092 (O_2092,N_17349,N_19630);
nand UO_2093 (O_2093,N_16841,N_19569);
nand UO_2094 (O_2094,N_16082,N_19523);
and UO_2095 (O_2095,N_16309,N_16107);
nor UO_2096 (O_2096,N_17801,N_16810);
nor UO_2097 (O_2097,N_16303,N_19898);
nand UO_2098 (O_2098,N_16998,N_18935);
or UO_2099 (O_2099,N_19968,N_19762);
and UO_2100 (O_2100,N_16079,N_16138);
or UO_2101 (O_2101,N_18812,N_18036);
nor UO_2102 (O_2102,N_16500,N_18379);
nand UO_2103 (O_2103,N_16613,N_17921);
xnor UO_2104 (O_2104,N_18107,N_17834);
or UO_2105 (O_2105,N_18127,N_19650);
or UO_2106 (O_2106,N_19306,N_19884);
xnor UO_2107 (O_2107,N_17350,N_17756);
and UO_2108 (O_2108,N_19800,N_18888);
and UO_2109 (O_2109,N_17651,N_17709);
xor UO_2110 (O_2110,N_18134,N_16230);
or UO_2111 (O_2111,N_18895,N_19997);
nand UO_2112 (O_2112,N_17862,N_16188);
nand UO_2113 (O_2113,N_17657,N_16320);
xnor UO_2114 (O_2114,N_16740,N_17664);
nor UO_2115 (O_2115,N_17509,N_19843);
or UO_2116 (O_2116,N_19250,N_16905);
or UO_2117 (O_2117,N_16221,N_17172);
or UO_2118 (O_2118,N_19114,N_18736);
nor UO_2119 (O_2119,N_19784,N_19904);
or UO_2120 (O_2120,N_19461,N_16130);
xor UO_2121 (O_2121,N_17333,N_19411);
or UO_2122 (O_2122,N_17956,N_16678);
and UO_2123 (O_2123,N_16679,N_19413);
nor UO_2124 (O_2124,N_18774,N_16189);
and UO_2125 (O_2125,N_16379,N_16700);
and UO_2126 (O_2126,N_16649,N_17674);
nand UO_2127 (O_2127,N_16573,N_17850);
xnor UO_2128 (O_2128,N_19096,N_16587);
xor UO_2129 (O_2129,N_19260,N_19222);
nor UO_2130 (O_2130,N_17996,N_18718);
nor UO_2131 (O_2131,N_19749,N_19967);
or UO_2132 (O_2132,N_18696,N_19915);
nand UO_2133 (O_2133,N_16193,N_17156);
nor UO_2134 (O_2134,N_16027,N_16225);
and UO_2135 (O_2135,N_17032,N_19865);
or UO_2136 (O_2136,N_19232,N_16757);
nand UO_2137 (O_2137,N_19312,N_16003);
or UO_2138 (O_2138,N_18623,N_18953);
and UO_2139 (O_2139,N_19098,N_16738);
nor UO_2140 (O_2140,N_17540,N_18380);
or UO_2141 (O_2141,N_19187,N_16473);
nand UO_2142 (O_2142,N_17471,N_19257);
and UO_2143 (O_2143,N_19846,N_18726);
nand UO_2144 (O_2144,N_17554,N_17791);
or UO_2145 (O_2145,N_16575,N_17099);
nand UO_2146 (O_2146,N_16728,N_17140);
nand UO_2147 (O_2147,N_19320,N_17819);
nand UO_2148 (O_2148,N_16353,N_16841);
xor UO_2149 (O_2149,N_17543,N_18414);
or UO_2150 (O_2150,N_17197,N_18036);
or UO_2151 (O_2151,N_19819,N_16143);
nand UO_2152 (O_2152,N_19637,N_18383);
xnor UO_2153 (O_2153,N_16249,N_16798);
nand UO_2154 (O_2154,N_17999,N_17109);
nand UO_2155 (O_2155,N_17231,N_17097);
and UO_2156 (O_2156,N_17131,N_17963);
and UO_2157 (O_2157,N_18357,N_17926);
nor UO_2158 (O_2158,N_17912,N_16052);
nor UO_2159 (O_2159,N_19077,N_19732);
or UO_2160 (O_2160,N_19021,N_18133);
xnor UO_2161 (O_2161,N_18902,N_19564);
nand UO_2162 (O_2162,N_19203,N_19428);
nor UO_2163 (O_2163,N_19363,N_16403);
and UO_2164 (O_2164,N_19417,N_16628);
or UO_2165 (O_2165,N_18162,N_18671);
xor UO_2166 (O_2166,N_16428,N_18971);
nor UO_2167 (O_2167,N_18188,N_17450);
and UO_2168 (O_2168,N_16006,N_16282);
xor UO_2169 (O_2169,N_16592,N_19914);
nor UO_2170 (O_2170,N_18990,N_16063);
and UO_2171 (O_2171,N_16848,N_17477);
nor UO_2172 (O_2172,N_17823,N_17087);
nor UO_2173 (O_2173,N_16335,N_18002);
or UO_2174 (O_2174,N_16907,N_19018);
nand UO_2175 (O_2175,N_18122,N_17239);
nand UO_2176 (O_2176,N_19288,N_16746);
or UO_2177 (O_2177,N_16741,N_17083);
and UO_2178 (O_2178,N_16656,N_19107);
nand UO_2179 (O_2179,N_18301,N_19939);
and UO_2180 (O_2180,N_17778,N_17684);
or UO_2181 (O_2181,N_17965,N_19861);
nand UO_2182 (O_2182,N_17933,N_19514);
nor UO_2183 (O_2183,N_18555,N_16396);
nand UO_2184 (O_2184,N_18554,N_16528);
nor UO_2185 (O_2185,N_18183,N_18698);
and UO_2186 (O_2186,N_18574,N_18658);
and UO_2187 (O_2187,N_18158,N_19436);
or UO_2188 (O_2188,N_18013,N_17885);
xnor UO_2189 (O_2189,N_18469,N_16117);
nand UO_2190 (O_2190,N_19872,N_17103);
or UO_2191 (O_2191,N_16035,N_17794);
xor UO_2192 (O_2192,N_18726,N_19133);
nor UO_2193 (O_2193,N_16902,N_17264);
or UO_2194 (O_2194,N_16103,N_17502);
xor UO_2195 (O_2195,N_18789,N_17162);
nand UO_2196 (O_2196,N_18296,N_19356);
and UO_2197 (O_2197,N_16507,N_17701);
nor UO_2198 (O_2198,N_16956,N_17659);
xnor UO_2199 (O_2199,N_17922,N_17833);
and UO_2200 (O_2200,N_17268,N_19010);
nand UO_2201 (O_2201,N_17331,N_16433);
and UO_2202 (O_2202,N_18226,N_18783);
xor UO_2203 (O_2203,N_19537,N_17646);
xor UO_2204 (O_2204,N_17096,N_16447);
or UO_2205 (O_2205,N_17540,N_18959);
nand UO_2206 (O_2206,N_19626,N_17357);
nor UO_2207 (O_2207,N_19435,N_18408);
nand UO_2208 (O_2208,N_17092,N_17938);
nor UO_2209 (O_2209,N_19235,N_17047);
and UO_2210 (O_2210,N_17808,N_17855);
or UO_2211 (O_2211,N_19334,N_17223);
nor UO_2212 (O_2212,N_17578,N_17065);
nor UO_2213 (O_2213,N_19733,N_17677);
nand UO_2214 (O_2214,N_17662,N_18042);
xor UO_2215 (O_2215,N_18110,N_18900);
and UO_2216 (O_2216,N_19344,N_17157);
or UO_2217 (O_2217,N_18620,N_17582);
xnor UO_2218 (O_2218,N_16909,N_16458);
nor UO_2219 (O_2219,N_19146,N_17207);
nand UO_2220 (O_2220,N_18457,N_16610);
nand UO_2221 (O_2221,N_19276,N_16405);
or UO_2222 (O_2222,N_17698,N_18936);
xnor UO_2223 (O_2223,N_18792,N_19262);
and UO_2224 (O_2224,N_17659,N_17496);
or UO_2225 (O_2225,N_19989,N_19163);
or UO_2226 (O_2226,N_16591,N_18180);
or UO_2227 (O_2227,N_16038,N_17881);
nor UO_2228 (O_2228,N_19099,N_18546);
or UO_2229 (O_2229,N_17443,N_19787);
or UO_2230 (O_2230,N_18819,N_17337);
and UO_2231 (O_2231,N_18097,N_18470);
nor UO_2232 (O_2232,N_17778,N_17276);
xnor UO_2233 (O_2233,N_19371,N_17549);
and UO_2234 (O_2234,N_16013,N_18018);
nand UO_2235 (O_2235,N_16121,N_16302);
or UO_2236 (O_2236,N_16316,N_17841);
nor UO_2237 (O_2237,N_19086,N_16965);
or UO_2238 (O_2238,N_17027,N_19647);
xor UO_2239 (O_2239,N_17344,N_17390);
or UO_2240 (O_2240,N_16080,N_17597);
or UO_2241 (O_2241,N_19518,N_16472);
xor UO_2242 (O_2242,N_17968,N_18927);
nor UO_2243 (O_2243,N_18788,N_19498);
and UO_2244 (O_2244,N_16458,N_18512);
xnor UO_2245 (O_2245,N_17467,N_16883);
nand UO_2246 (O_2246,N_18964,N_16311);
or UO_2247 (O_2247,N_16862,N_19025);
xnor UO_2248 (O_2248,N_17224,N_17374);
and UO_2249 (O_2249,N_16692,N_16761);
nor UO_2250 (O_2250,N_18537,N_19616);
nor UO_2251 (O_2251,N_17538,N_18870);
nor UO_2252 (O_2252,N_17856,N_16545);
xnor UO_2253 (O_2253,N_16460,N_18589);
and UO_2254 (O_2254,N_18908,N_17763);
nor UO_2255 (O_2255,N_19763,N_18292);
xor UO_2256 (O_2256,N_19795,N_17547);
or UO_2257 (O_2257,N_18525,N_17971);
or UO_2258 (O_2258,N_18100,N_19915);
nand UO_2259 (O_2259,N_17528,N_16566);
nor UO_2260 (O_2260,N_19632,N_17847);
nand UO_2261 (O_2261,N_18756,N_17380);
nor UO_2262 (O_2262,N_17169,N_19020);
xnor UO_2263 (O_2263,N_19826,N_19240);
or UO_2264 (O_2264,N_19607,N_17330);
nor UO_2265 (O_2265,N_18566,N_16817);
and UO_2266 (O_2266,N_16319,N_19223);
nor UO_2267 (O_2267,N_18860,N_17321);
and UO_2268 (O_2268,N_19586,N_16231);
and UO_2269 (O_2269,N_19059,N_18488);
nor UO_2270 (O_2270,N_19980,N_19249);
or UO_2271 (O_2271,N_18270,N_19819);
or UO_2272 (O_2272,N_18893,N_17998);
nand UO_2273 (O_2273,N_19477,N_18659);
or UO_2274 (O_2274,N_16253,N_19364);
xor UO_2275 (O_2275,N_16878,N_19921);
and UO_2276 (O_2276,N_18885,N_17306);
xnor UO_2277 (O_2277,N_16486,N_19016);
xor UO_2278 (O_2278,N_17404,N_18917);
xor UO_2279 (O_2279,N_19663,N_19176);
nor UO_2280 (O_2280,N_19253,N_16530);
and UO_2281 (O_2281,N_19519,N_19879);
and UO_2282 (O_2282,N_16888,N_19742);
nor UO_2283 (O_2283,N_18980,N_17742);
and UO_2284 (O_2284,N_19473,N_18102);
or UO_2285 (O_2285,N_19769,N_16812);
or UO_2286 (O_2286,N_17309,N_16906);
xnor UO_2287 (O_2287,N_18190,N_16062);
xor UO_2288 (O_2288,N_19413,N_19861);
xor UO_2289 (O_2289,N_16466,N_17743);
xnor UO_2290 (O_2290,N_17905,N_18069);
nor UO_2291 (O_2291,N_18810,N_19465);
nor UO_2292 (O_2292,N_18697,N_19162);
and UO_2293 (O_2293,N_16979,N_17512);
or UO_2294 (O_2294,N_18955,N_18719);
nor UO_2295 (O_2295,N_16656,N_18307);
or UO_2296 (O_2296,N_18129,N_18703);
and UO_2297 (O_2297,N_19226,N_18278);
nor UO_2298 (O_2298,N_19348,N_17384);
or UO_2299 (O_2299,N_16324,N_17821);
nand UO_2300 (O_2300,N_17503,N_16520);
nand UO_2301 (O_2301,N_16894,N_18259);
nor UO_2302 (O_2302,N_17883,N_19736);
and UO_2303 (O_2303,N_18216,N_17269);
nor UO_2304 (O_2304,N_17928,N_17779);
nand UO_2305 (O_2305,N_18266,N_18338);
and UO_2306 (O_2306,N_19753,N_17965);
and UO_2307 (O_2307,N_17139,N_18623);
and UO_2308 (O_2308,N_18311,N_17678);
nor UO_2309 (O_2309,N_17370,N_19648);
or UO_2310 (O_2310,N_19409,N_16273);
nand UO_2311 (O_2311,N_17266,N_18550);
and UO_2312 (O_2312,N_17438,N_18799);
and UO_2313 (O_2313,N_17619,N_19218);
or UO_2314 (O_2314,N_16049,N_16589);
nor UO_2315 (O_2315,N_16863,N_16845);
or UO_2316 (O_2316,N_19957,N_16477);
nor UO_2317 (O_2317,N_16022,N_17131);
nor UO_2318 (O_2318,N_18221,N_18932);
nand UO_2319 (O_2319,N_19978,N_18625);
nand UO_2320 (O_2320,N_19795,N_18716);
and UO_2321 (O_2321,N_16477,N_17656);
nor UO_2322 (O_2322,N_16166,N_16391);
nand UO_2323 (O_2323,N_17559,N_17107);
xor UO_2324 (O_2324,N_18251,N_18069);
or UO_2325 (O_2325,N_17020,N_18324);
nor UO_2326 (O_2326,N_16153,N_17467);
and UO_2327 (O_2327,N_18814,N_19919);
xor UO_2328 (O_2328,N_16430,N_18320);
nor UO_2329 (O_2329,N_19117,N_19092);
and UO_2330 (O_2330,N_19847,N_18072);
or UO_2331 (O_2331,N_18069,N_19283);
nand UO_2332 (O_2332,N_16750,N_19383);
xor UO_2333 (O_2333,N_19153,N_16679);
nand UO_2334 (O_2334,N_17757,N_17143);
xnor UO_2335 (O_2335,N_19415,N_17306);
or UO_2336 (O_2336,N_19001,N_18887);
nand UO_2337 (O_2337,N_17531,N_17661);
xor UO_2338 (O_2338,N_17735,N_16856);
or UO_2339 (O_2339,N_18147,N_18021);
and UO_2340 (O_2340,N_19580,N_16553);
and UO_2341 (O_2341,N_17850,N_16748);
or UO_2342 (O_2342,N_19100,N_16782);
or UO_2343 (O_2343,N_16474,N_19229);
xnor UO_2344 (O_2344,N_17675,N_17930);
or UO_2345 (O_2345,N_16360,N_16612);
xnor UO_2346 (O_2346,N_16116,N_17837);
nor UO_2347 (O_2347,N_19184,N_19186);
xor UO_2348 (O_2348,N_17224,N_16105);
nor UO_2349 (O_2349,N_18905,N_17809);
nand UO_2350 (O_2350,N_17015,N_16146);
nor UO_2351 (O_2351,N_18939,N_17386);
nand UO_2352 (O_2352,N_17929,N_17247);
or UO_2353 (O_2353,N_17412,N_18178);
nor UO_2354 (O_2354,N_18214,N_17696);
and UO_2355 (O_2355,N_17694,N_16549);
nor UO_2356 (O_2356,N_19187,N_16289);
or UO_2357 (O_2357,N_19848,N_17779);
and UO_2358 (O_2358,N_17205,N_18202);
nor UO_2359 (O_2359,N_16378,N_18061);
and UO_2360 (O_2360,N_18551,N_18978);
or UO_2361 (O_2361,N_19607,N_16198);
nand UO_2362 (O_2362,N_18553,N_19563);
or UO_2363 (O_2363,N_16086,N_17502);
and UO_2364 (O_2364,N_18214,N_17381);
or UO_2365 (O_2365,N_18939,N_16530);
and UO_2366 (O_2366,N_16014,N_18280);
or UO_2367 (O_2367,N_18552,N_17584);
nand UO_2368 (O_2368,N_18104,N_18221);
or UO_2369 (O_2369,N_18066,N_16860);
xor UO_2370 (O_2370,N_16353,N_18784);
nand UO_2371 (O_2371,N_17074,N_19858);
nand UO_2372 (O_2372,N_19666,N_18806);
nand UO_2373 (O_2373,N_17444,N_19176);
xnor UO_2374 (O_2374,N_16215,N_18803);
and UO_2375 (O_2375,N_18608,N_18643);
nand UO_2376 (O_2376,N_16975,N_18967);
and UO_2377 (O_2377,N_16147,N_16691);
and UO_2378 (O_2378,N_16418,N_19588);
or UO_2379 (O_2379,N_19111,N_18068);
nor UO_2380 (O_2380,N_18347,N_18554);
nand UO_2381 (O_2381,N_17535,N_19458);
and UO_2382 (O_2382,N_18397,N_19600);
and UO_2383 (O_2383,N_17180,N_17819);
and UO_2384 (O_2384,N_18560,N_19323);
and UO_2385 (O_2385,N_17827,N_18432);
nor UO_2386 (O_2386,N_16510,N_17170);
nand UO_2387 (O_2387,N_16252,N_18853);
xor UO_2388 (O_2388,N_18311,N_19891);
xor UO_2389 (O_2389,N_17546,N_18958);
nand UO_2390 (O_2390,N_18060,N_17372);
and UO_2391 (O_2391,N_19932,N_16468);
or UO_2392 (O_2392,N_18192,N_16251);
xnor UO_2393 (O_2393,N_17735,N_19886);
nor UO_2394 (O_2394,N_19807,N_18973);
xor UO_2395 (O_2395,N_17161,N_19804);
xnor UO_2396 (O_2396,N_16358,N_16478);
or UO_2397 (O_2397,N_16586,N_17892);
and UO_2398 (O_2398,N_16654,N_16665);
nand UO_2399 (O_2399,N_17924,N_19042);
or UO_2400 (O_2400,N_17245,N_17100);
nand UO_2401 (O_2401,N_16489,N_19840);
nand UO_2402 (O_2402,N_19806,N_16670);
or UO_2403 (O_2403,N_18853,N_17734);
nand UO_2404 (O_2404,N_19110,N_18758);
nor UO_2405 (O_2405,N_18276,N_16048);
nand UO_2406 (O_2406,N_16944,N_16228);
or UO_2407 (O_2407,N_16297,N_16737);
or UO_2408 (O_2408,N_16812,N_16926);
nor UO_2409 (O_2409,N_16824,N_17658);
xor UO_2410 (O_2410,N_17252,N_18199);
and UO_2411 (O_2411,N_16423,N_19318);
nor UO_2412 (O_2412,N_18252,N_17874);
xor UO_2413 (O_2413,N_18529,N_19033);
nand UO_2414 (O_2414,N_18290,N_19747);
and UO_2415 (O_2415,N_18023,N_19171);
nand UO_2416 (O_2416,N_18108,N_19143);
nand UO_2417 (O_2417,N_17290,N_19287);
and UO_2418 (O_2418,N_18073,N_16102);
and UO_2419 (O_2419,N_16395,N_18823);
and UO_2420 (O_2420,N_19464,N_17574);
or UO_2421 (O_2421,N_17559,N_19393);
or UO_2422 (O_2422,N_18396,N_17684);
and UO_2423 (O_2423,N_18582,N_19834);
and UO_2424 (O_2424,N_17368,N_18261);
and UO_2425 (O_2425,N_17153,N_19488);
xor UO_2426 (O_2426,N_19177,N_17336);
xor UO_2427 (O_2427,N_18869,N_18142);
nor UO_2428 (O_2428,N_19722,N_18536);
or UO_2429 (O_2429,N_19953,N_19705);
xnor UO_2430 (O_2430,N_19442,N_17581);
and UO_2431 (O_2431,N_16873,N_17193);
nor UO_2432 (O_2432,N_17095,N_19627);
nand UO_2433 (O_2433,N_16162,N_18622);
nand UO_2434 (O_2434,N_16503,N_16803);
xor UO_2435 (O_2435,N_19955,N_18351);
nor UO_2436 (O_2436,N_19271,N_17080);
and UO_2437 (O_2437,N_17396,N_17741);
and UO_2438 (O_2438,N_18101,N_18426);
xor UO_2439 (O_2439,N_18470,N_16031);
xnor UO_2440 (O_2440,N_18754,N_18075);
xnor UO_2441 (O_2441,N_18496,N_19457);
nand UO_2442 (O_2442,N_19820,N_19670);
and UO_2443 (O_2443,N_18472,N_16107);
nand UO_2444 (O_2444,N_17569,N_18078);
nand UO_2445 (O_2445,N_16757,N_17352);
nand UO_2446 (O_2446,N_18968,N_18984);
xor UO_2447 (O_2447,N_17817,N_18869);
or UO_2448 (O_2448,N_16479,N_17280);
nand UO_2449 (O_2449,N_19457,N_16591);
nor UO_2450 (O_2450,N_16759,N_19710);
nor UO_2451 (O_2451,N_19365,N_18275);
xor UO_2452 (O_2452,N_19635,N_18479);
and UO_2453 (O_2453,N_17463,N_17453);
or UO_2454 (O_2454,N_19499,N_16874);
or UO_2455 (O_2455,N_17749,N_16924);
xnor UO_2456 (O_2456,N_19725,N_18705);
nor UO_2457 (O_2457,N_19914,N_19986);
xnor UO_2458 (O_2458,N_19025,N_19070);
nor UO_2459 (O_2459,N_19041,N_19260);
nand UO_2460 (O_2460,N_19518,N_19559);
nor UO_2461 (O_2461,N_18593,N_19951);
and UO_2462 (O_2462,N_18972,N_17200);
and UO_2463 (O_2463,N_19631,N_18267);
nor UO_2464 (O_2464,N_16273,N_18445);
nor UO_2465 (O_2465,N_17873,N_19767);
and UO_2466 (O_2466,N_17182,N_16789);
nor UO_2467 (O_2467,N_17795,N_19660);
or UO_2468 (O_2468,N_18205,N_17536);
or UO_2469 (O_2469,N_17437,N_19533);
nand UO_2470 (O_2470,N_18346,N_17347);
and UO_2471 (O_2471,N_17398,N_17995);
or UO_2472 (O_2472,N_18932,N_17854);
nor UO_2473 (O_2473,N_18783,N_18604);
and UO_2474 (O_2474,N_17577,N_19394);
nand UO_2475 (O_2475,N_16643,N_18876);
xnor UO_2476 (O_2476,N_16428,N_18630);
or UO_2477 (O_2477,N_16560,N_16160);
nor UO_2478 (O_2478,N_19737,N_19011);
and UO_2479 (O_2479,N_18978,N_19191);
and UO_2480 (O_2480,N_18438,N_19634);
xnor UO_2481 (O_2481,N_18452,N_19368);
and UO_2482 (O_2482,N_19422,N_19492);
xnor UO_2483 (O_2483,N_19001,N_18619);
xor UO_2484 (O_2484,N_16761,N_18352);
or UO_2485 (O_2485,N_18628,N_18196);
or UO_2486 (O_2486,N_16980,N_18215);
or UO_2487 (O_2487,N_16297,N_17621);
nor UO_2488 (O_2488,N_18468,N_17788);
xnor UO_2489 (O_2489,N_18745,N_19470);
nor UO_2490 (O_2490,N_17640,N_16997);
and UO_2491 (O_2491,N_16374,N_17675);
nor UO_2492 (O_2492,N_16078,N_17636);
or UO_2493 (O_2493,N_17241,N_17831);
nand UO_2494 (O_2494,N_16932,N_18561);
xnor UO_2495 (O_2495,N_19464,N_19281);
nand UO_2496 (O_2496,N_17941,N_17186);
nand UO_2497 (O_2497,N_16500,N_18507);
and UO_2498 (O_2498,N_17751,N_19425);
and UO_2499 (O_2499,N_17421,N_18696);
endmodule