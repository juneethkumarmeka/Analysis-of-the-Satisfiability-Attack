module basic_500_3000_500_15_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_479,In_307);
nand U1 (N_1,In_362,In_84);
nand U2 (N_2,In_211,In_258);
and U3 (N_3,In_234,In_92);
nor U4 (N_4,In_207,In_315);
nand U5 (N_5,In_169,In_311);
nand U6 (N_6,In_320,In_344);
nor U7 (N_7,In_420,In_67);
or U8 (N_8,In_0,In_284);
xor U9 (N_9,In_221,In_236);
nor U10 (N_10,In_225,In_329);
or U11 (N_11,In_488,In_109);
nor U12 (N_12,In_251,In_465);
and U13 (N_13,In_399,In_499);
or U14 (N_14,In_494,In_228);
xor U15 (N_15,In_66,In_418);
nand U16 (N_16,In_456,In_272);
xnor U17 (N_17,In_222,In_128);
or U18 (N_18,In_203,In_87);
nor U19 (N_19,In_191,In_4);
and U20 (N_20,In_215,In_496);
xor U21 (N_21,In_247,In_47);
nor U22 (N_22,In_59,In_483);
and U23 (N_23,In_235,In_202);
and U24 (N_24,In_130,In_46);
and U25 (N_25,In_93,In_440);
nor U26 (N_26,In_490,In_40);
nor U27 (N_27,In_83,In_41);
or U28 (N_28,In_184,In_357);
or U29 (N_29,In_413,In_133);
nor U30 (N_30,In_443,In_398);
xnor U31 (N_31,In_308,In_190);
xor U32 (N_32,In_462,In_101);
xnor U33 (N_33,In_178,In_147);
and U34 (N_34,In_121,In_444);
or U35 (N_35,In_277,In_297);
nor U36 (N_36,In_115,In_13);
nand U37 (N_37,In_259,In_437);
or U38 (N_38,In_82,In_487);
nor U39 (N_39,In_339,In_233);
and U40 (N_40,In_127,In_60);
or U41 (N_41,In_267,In_38);
and U42 (N_42,In_52,In_466);
nor U43 (N_43,In_55,In_154);
nor U44 (N_44,In_396,In_112);
xor U45 (N_45,In_194,In_209);
and U46 (N_46,In_15,In_469);
nor U47 (N_47,In_114,In_160);
and U48 (N_48,In_438,In_69);
and U49 (N_49,In_368,In_238);
nor U50 (N_50,In_250,In_102);
nand U51 (N_51,In_255,In_376);
nand U52 (N_52,In_150,In_419);
xor U53 (N_53,In_261,In_116);
xor U54 (N_54,In_390,In_324);
or U55 (N_55,In_491,In_343);
and U56 (N_56,In_355,In_54);
nand U57 (N_57,In_91,In_423);
and U58 (N_58,In_275,In_64);
nand U59 (N_59,In_493,In_135);
nand U60 (N_60,In_379,In_432);
xnor U61 (N_61,In_156,In_6);
nand U62 (N_62,In_361,In_472);
or U63 (N_63,In_192,In_338);
or U64 (N_64,In_220,In_463);
nand U65 (N_65,In_380,In_268);
and U66 (N_66,In_484,In_172);
nand U67 (N_67,In_45,In_245);
nand U68 (N_68,In_14,In_446);
nor U69 (N_69,In_336,In_134);
nor U70 (N_70,In_348,In_240);
nor U71 (N_71,In_241,In_212);
xnor U72 (N_72,In_205,In_57);
or U73 (N_73,In_18,In_447);
or U74 (N_74,In_283,In_181);
xor U75 (N_75,In_198,In_206);
nand U76 (N_76,In_435,In_36);
xnor U77 (N_77,In_170,In_177);
and U78 (N_78,In_131,In_327);
nand U79 (N_79,In_152,In_303);
nor U80 (N_80,In_249,In_86);
or U81 (N_81,In_281,In_313);
xor U82 (N_82,In_468,In_481);
nand U83 (N_83,In_351,In_22);
nor U84 (N_84,In_319,In_299);
nand U85 (N_85,In_180,In_157);
nand U86 (N_86,In_142,In_291);
nor U87 (N_87,In_95,In_372);
and U88 (N_88,In_79,In_185);
or U89 (N_89,In_53,In_23);
and U90 (N_90,In_371,In_388);
and U91 (N_91,In_226,In_270);
nor U92 (N_92,In_35,In_8);
nor U93 (N_93,In_495,In_337);
xor U94 (N_94,In_98,In_309);
and U95 (N_95,In_44,In_364);
and U96 (N_96,In_56,In_402);
and U97 (N_97,In_401,In_293);
or U98 (N_98,In_25,In_197);
xnor U99 (N_99,In_76,In_5);
and U100 (N_100,In_457,In_171);
nor U101 (N_101,In_410,In_394);
nor U102 (N_102,In_246,In_416);
nor U103 (N_103,In_100,In_471);
and U104 (N_104,In_143,In_391);
or U105 (N_105,In_331,In_218);
nand U106 (N_106,In_189,In_480);
nand U107 (N_107,In_411,In_70);
and U108 (N_108,In_378,In_237);
nor U109 (N_109,In_162,In_335);
xor U110 (N_110,In_2,In_365);
and U111 (N_111,In_49,In_153);
xor U112 (N_112,In_434,In_385);
and U113 (N_113,In_19,In_295);
nand U114 (N_114,In_395,In_405);
nor U115 (N_115,In_108,In_455);
nand U116 (N_116,In_296,In_386);
nand U117 (N_117,In_350,In_298);
and U118 (N_118,In_342,In_289);
nor U119 (N_119,In_467,In_408);
or U120 (N_120,In_294,In_120);
xor U121 (N_121,In_369,In_263);
nand U122 (N_122,In_353,In_43);
nor U123 (N_123,In_474,In_118);
and U124 (N_124,In_155,In_370);
or U125 (N_125,In_227,In_132);
nor U126 (N_126,In_454,In_477);
xnor U127 (N_127,In_124,In_166);
xor U128 (N_128,In_78,In_193);
xor U129 (N_129,In_11,In_269);
nor U130 (N_130,In_266,In_183);
nand U131 (N_131,In_244,In_424);
nor U132 (N_132,In_204,In_39);
and U133 (N_133,In_210,In_97);
and U134 (N_134,In_9,In_302);
xnor U135 (N_135,In_312,In_103);
and U136 (N_136,In_174,In_288);
nor U137 (N_137,In_326,In_145);
and U138 (N_138,In_290,In_99);
xor U139 (N_139,In_450,In_34);
nor U140 (N_140,In_224,In_200);
xor U141 (N_141,In_347,In_285);
and U142 (N_142,In_397,In_146);
xnor U143 (N_143,In_179,In_85);
nor U144 (N_144,In_393,In_163);
and U145 (N_145,In_88,In_51);
and U146 (N_146,In_129,In_201);
nand U147 (N_147,In_136,In_30);
or U148 (N_148,In_188,In_341);
or U149 (N_149,In_485,In_107);
xor U150 (N_150,In_445,In_28);
nor U151 (N_151,In_415,In_317);
and U152 (N_152,In_328,In_3);
and U153 (N_153,In_77,In_453);
or U154 (N_154,In_300,In_256);
xnor U155 (N_155,In_243,In_216);
or U156 (N_156,In_126,In_306);
nand U157 (N_157,In_187,In_213);
or U158 (N_158,In_72,In_33);
nor U159 (N_159,In_223,In_219);
and U160 (N_160,In_400,In_158);
nor U161 (N_161,In_403,In_404);
nor U162 (N_162,In_117,In_63);
xor U163 (N_163,In_433,In_470);
xor U164 (N_164,In_122,In_42);
and U165 (N_165,In_325,In_492);
nand U166 (N_166,In_274,In_473);
nand U167 (N_167,In_17,In_497);
nand U168 (N_168,In_374,In_20);
nor U169 (N_169,In_359,In_429);
and U170 (N_170,In_32,In_367);
or U171 (N_171,In_358,In_29);
or U172 (N_172,In_125,In_31);
nor U173 (N_173,In_217,In_425);
or U174 (N_174,In_140,In_486);
nor U175 (N_175,In_75,In_356);
or U176 (N_176,In_37,In_330);
nor U177 (N_177,In_231,In_141);
or U178 (N_178,In_175,In_90);
and U179 (N_179,In_301,In_196);
xor U180 (N_180,In_304,In_248);
or U181 (N_181,In_366,In_242);
and U182 (N_182,In_292,In_26);
xor U183 (N_183,In_164,In_61);
or U184 (N_184,In_278,In_199);
nand U185 (N_185,In_360,In_73);
nor U186 (N_186,In_373,In_286);
xnor U187 (N_187,In_229,In_239);
nor U188 (N_188,In_186,In_254);
and U189 (N_189,In_449,In_68);
nand U190 (N_190,In_159,In_214);
xor U191 (N_191,In_138,In_458);
xnor U192 (N_192,In_305,In_441);
xnor U193 (N_193,In_161,In_406);
nand U194 (N_194,In_273,In_173);
or U195 (N_195,In_321,In_382);
xnor U196 (N_196,In_111,In_460);
and U197 (N_197,In_113,In_276);
nor U198 (N_198,In_230,In_94);
xnor U199 (N_199,In_260,In_81);
nor U200 (N_200,N_149,N_47);
and U201 (N_201,N_187,N_84);
or U202 (N_202,N_116,N_49);
or U203 (N_203,N_120,N_184);
nand U204 (N_204,In_148,N_72);
and U205 (N_205,N_97,In_80);
or U206 (N_206,N_109,In_182);
nor U207 (N_207,In_282,In_176);
and U208 (N_208,In_318,N_167);
and U209 (N_209,N_15,N_8);
xnor U210 (N_210,N_65,N_115);
and U211 (N_211,N_4,N_28);
nor U212 (N_212,N_144,N_190);
and U213 (N_213,In_123,In_208);
nor U214 (N_214,N_95,N_148);
nor U215 (N_215,In_414,N_102);
nand U216 (N_216,N_106,N_127);
and U217 (N_217,N_36,N_16);
nor U218 (N_218,N_44,N_98);
nor U219 (N_219,In_144,N_87);
xor U220 (N_220,N_3,In_459);
nand U221 (N_221,In_1,N_21);
or U222 (N_222,N_59,N_179);
and U223 (N_223,In_489,In_62);
or U224 (N_224,N_132,N_197);
or U225 (N_225,N_56,N_43);
nor U226 (N_226,N_156,In_427);
nor U227 (N_227,N_171,In_349);
and U228 (N_228,N_76,N_101);
or U229 (N_229,In_314,In_451);
nand U230 (N_230,In_334,N_118);
xnor U231 (N_231,N_129,N_93);
xnor U232 (N_232,In_431,N_29);
nand U233 (N_233,N_54,N_74);
xnor U234 (N_234,N_42,In_12);
nand U235 (N_235,N_182,N_178);
nand U236 (N_236,N_73,In_279);
xnor U237 (N_237,N_165,N_153);
and U238 (N_238,N_113,In_352);
nor U239 (N_239,In_10,In_271);
nor U240 (N_240,N_166,N_62);
nand U241 (N_241,N_2,In_232);
nor U242 (N_242,N_196,In_105);
xnor U243 (N_243,N_75,In_74);
nor U244 (N_244,N_5,N_80);
nand U245 (N_245,N_157,N_22);
nand U246 (N_246,N_195,N_199);
or U247 (N_247,In_167,In_428);
xnor U248 (N_248,N_40,In_333);
nor U249 (N_249,N_27,In_165);
nand U250 (N_250,N_60,N_161);
nand U251 (N_251,In_71,N_136);
xor U252 (N_252,N_31,N_53);
nand U253 (N_253,N_20,In_422);
nand U254 (N_254,N_33,N_0);
and U255 (N_255,N_188,N_96);
xnor U256 (N_256,N_143,N_107);
or U257 (N_257,N_14,N_38);
and U258 (N_258,N_13,N_145);
and U259 (N_259,N_126,N_58);
nand U260 (N_260,In_475,N_192);
and U261 (N_261,In_354,In_65);
or U262 (N_262,N_173,N_68);
and U263 (N_263,In_323,In_16);
nand U264 (N_264,N_34,N_194);
and U265 (N_265,N_82,In_384);
nand U266 (N_266,N_185,N_19);
and U267 (N_267,In_498,In_332);
nor U268 (N_268,In_106,N_152);
or U269 (N_269,N_94,In_452);
nand U270 (N_270,N_128,N_183);
and U271 (N_271,N_12,N_81);
nor U272 (N_272,In_119,N_25);
nor U273 (N_273,N_154,N_110);
nand U274 (N_274,In_137,N_150);
nor U275 (N_275,N_146,N_92);
or U276 (N_276,In_149,N_122);
and U277 (N_277,In_407,N_158);
nand U278 (N_278,N_6,N_191);
xor U279 (N_279,In_389,N_64);
nand U280 (N_280,N_46,In_340);
xnor U281 (N_281,N_155,N_162);
xor U282 (N_282,In_287,N_99);
or U283 (N_283,N_169,N_181);
or U284 (N_284,N_57,N_90);
nand U285 (N_285,N_121,N_163);
nor U286 (N_286,N_134,N_51);
and U287 (N_287,N_7,In_322);
nor U288 (N_288,N_105,In_387);
and U289 (N_289,In_104,N_91);
xnor U290 (N_290,N_138,In_265);
xor U291 (N_291,N_160,N_170);
xnor U292 (N_292,In_24,In_482);
or U293 (N_293,In_409,N_103);
nand U294 (N_294,N_141,In_21);
or U295 (N_295,N_135,In_168);
nor U296 (N_296,N_172,N_52);
xor U297 (N_297,N_131,In_375);
nor U298 (N_298,In_310,N_186);
nor U299 (N_299,N_140,In_436);
nand U300 (N_300,N_124,In_257);
nor U301 (N_301,N_48,N_37);
nor U302 (N_302,In_252,N_79);
xnor U303 (N_303,In_430,N_198);
and U304 (N_304,In_363,In_195);
or U305 (N_305,N_176,In_345);
or U306 (N_306,In_48,In_264);
and U307 (N_307,N_177,In_442);
nor U308 (N_308,N_117,N_77);
nand U309 (N_309,N_69,In_58);
and U310 (N_310,N_108,N_193);
and U311 (N_311,N_63,N_32);
nor U312 (N_312,In_392,N_50);
nor U313 (N_313,In_426,In_280);
nand U314 (N_314,In_381,N_55);
or U315 (N_315,N_130,N_180);
and U316 (N_316,N_86,In_89);
nand U317 (N_317,N_174,In_383);
or U318 (N_318,In_439,N_112);
and U319 (N_319,N_35,In_253);
and U320 (N_320,N_151,N_175);
nor U321 (N_321,In_417,In_262);
xnor U322 (N_322,N_88,N_71);
or U323 (N_323,N_137,N_30);
nand U324 (N_324,N_41,N_168);
nand U325 (N_325,N_147,In_27);
or U326 (N_326,N_119,N_61);
or U327 (N_327,N_123,N_139);
nand U328 (N_328,N_85,N_142);
or U329 (N_329,N_189,In_448);
or U330 (N_330,In_461,In_316);
xnor U331 (N_331,N_66,N_39);
xor U332 (N_332,In_7,N_9);
nand U333 (N_333,N_18,In_151);
xor U334 (N_334,In_478,N_78);
and U335 (N_335,N_159,N_83);
or U336 (N_336,N_10,N_17);
and U337 (N_337,N_125,N_111);
xnor U338 (N_338,In_464,In_96);
and U339 (N_339,In_50,N_67);
and U340 (N_340,N_11,In_476);
or U341 (N_341,N_70,N_23);
and U342 (N_342,N_45,In_377);
nor U343 (N_343,N_114,N_133);
nand U344 (N_344,N_89,N_24);
and U345 (N_345,N_100,In_110);
nor U346 (N_346,In_421,In_346);
and U347 (N_347,In_412,N_1);
nor U348 (N_348,In_139,N_164);
and U349 (N_349,N_26,N_104);
or U350 (N_350,N_124,N_77);
nand U351 (N_351,In_176,In_265);
nor U352 (N_352,N_93,N_94);
and U353 (N_353,N_73,N_189);
xor U354 (N_354,N_162,N_64);
and U355 (N_355,N_39,In_265);
xor U356 (N_356,In_383,N_137);
nand U357 (N_357,N_109,In_165);
xor U358 (N_358,N_168,In_264);
nand U359 (N_359,In_334,N_109);
and U360 (N_360,N_118,In_352);
or U361 (N_361,In_253,N_189);
nand U362 (N_362,N_164,In_280);
xor U363 (N_363,N_161,N_80);
and U364 (N_364,In_448,N_19);
or U365 (N_365,In_62,N_113);
or U366 (N_366,N_53,N_35);
nor U367 (N_367,N_39,N_23);
nand U368 (N_368,In_257,In_139);
or U369 (N_369,N_56,N_48);
or U370 (N_370,N_133,N_8);
xor U371 (N_371,N_125,In_478);
nand U372 (N_372,In_426,In_428);
and U373 (N_373,N_34,In_316);
xnor U374 (N_374,N_74,N_70);
nor U375 (N_375,N_105,N_123);
nor U376 (N_376,N_61,N_153);
and U377 (N_377,N_154,N_32);
xor U378 (N_378,N_0,In_340);
xnor U379 (N_379,N_104,In_489);
or U380 (N_380,N_6,N_165);
or U381 (N_381,In_442,N_161);
xnor U382 (N_382,N_175,In_10);
or U383 (N_383,N_68,In_50);
xnor U384 (N_384,N_119,In_119);
nor U385 (N_385,N_152,N_78);
nand U386 (N_386,In_168,N_40);
xnor U387 (N_387,In_349,N_10);
or U388 (N_388,N_125,N_35);
xnor U389 (N_389,N_65,In_340);
and U390 (N_390,In_105,In_62);
xor U391 (N_391,N_143,N_188);
xor U392 (N_392,In_422,In_381);
and U393 (N_393,N_8,In_208);
or U394 (N_394,In_271,N_187);
or U395 (N_395,In_12,N_166);
xnor U396 (N_396,In_340,N_94);
or U397 (N_397,In_139,In_448);
or U398 (N_398,N_142,In_10);
nand U399 (N_399,In_322,N_48);
xnor U400 (N_400,N_265,N_232);
nand U401 (N_401,N_294,N_276);
nand U402 (N_402,N_318,N_213);
nand U403 (N_403,N_204,N_254);
or U404 (N_404,N_336,N_343);
nand U405 (N_405,N_351,N_302);
xor U406 (N_406,N_348,N_396);
or U407 (N_407,N_297,N_205);
or U408 (N_408,N_378,N_328);
xnor U409 (N_409,N_299,N_372);
and U410 (N_410,N_275,N_218);
xnor U411 (N_411,N_390,N_251);
or U412 (N_412,N_235,N_236);
and U413 (N_413,N_356,N_341);
xnor U414 (N_414,N_360,N_370);
nor U415 (N_415,N_287,N_367);
nand U416 (N_416,N_329,N_395);
nor U417 (N_417,N_292,N_286);
and U418 (N_418,N_371,N_266);
or U419 (N_419,N_353,N_337);
nor U420 (N_420,N_375,N_221);
nand U421 (N_421,N_262,N_386);
and U422 (N_422,N_344,N_206);
xor U423 (N_423,N_284,N_285);
nor U424 (N_424,N_305,N_354);
xor U425 (N_425,N_338,N_200);
nand U426 (N_426,N_248,N_303);
xnor U427 (N_427,N_228,N_282);
and U428 (N_428,N_330,N_322);
or U429 (N_429,N_224,N_227);
nor U430 (N_430,N_393,N_258);
nor U431 (N_431,N_345,N_212);
or U432 (N_432,N_243,N_387);
xor U433 (N_433,N_270,N_382);
nand U434 (N_434,N_374,N_398);
and U435 (N_435,N_268,N_263);
nor U436 (N_436,N_277,N_225);
nand U437 (N_437,N_256,N_376);
and U438 (N_438,N_342,N_321);
and U439 (N_439,N_239,N_310);
nor U440 (N_440,N_267,N_269);
or U441 (N_441,N_392,N_234);
nand U442 (N_442,N_365,N_332);
xnor U443 (N_443,N_340,N_257);
or U444 (N_444,N_230,N_250);
xnor U445 (N_445,N_229,N_333);
nand U446 (N_446,N_201,N_331);
or U447 (N_447,N_242,N_352);
or U448 (N_448,N_355,N_347);
nand U449 (N_449,N_309,N_226);
and U450 (N_450,N_291,N_249);
xnor U451 (N_451,N_272,N_209);
nor U452 (N_452,N_397,N_279);
xor U453 (N_453,N_308,N_237);
nand U454 (N_454,N_389,N_203);
or U455 (N_455,N_307,N_346);
xnor U456 (N_456,N_274,N_383);
nand U457 (N_457,N_281,N_364);
nor U458 (N_458,N_246,N_244);
or U459 (N_459,N_293,N_306);
and U460 (N_460,N_369,N_253);
xnor U461 (N_461,N_207,N_252);
nand U462 (N_462,N_300,N_315);
and U463 (N_463,N_381,N_339);
nor U464 (N_464,N_289,N_264);
nor U465 (N_465,N_358,N_399);
or U466 (N_466,N_314,N_368);
nand U467 (N_467,N_311,N_359);
nor U468 (N_468,N_349,N_241);
nand U469 (N_469,N_202,N_335);
and U470 (N_470,N_220,N_324);
nor U471 (N_471,N_255,N_301);
and U472 (N_472,N_211,N_384);
nor U473 (N_473,N_216,N_350);
and U474 (N_474,N_357,N_316);
xnor U475 (N_475,N_394,N_327);
xnor U476 (N_476,N_231,N_326);
or U477 (N_477,N_377,N_288);
and U478 (N_478,N_215,N_325);
xor U479 (N_479,N_223,N_313);
and U480 (N_480,N_245,N_283);
and U481 (N_481,N_363,N_260);
nand U482 (N_482,N_319,N_240);
and U483 (N_483,N_222,N_388);
nor U484 (N_484,N_361,N_312);
nand U485 (N_485,N_296,N_233);
xor U486 (N_486,N_217,N_208);
or U487 (N_487,N_366,N_334);
or U488 (N_488,N_380,N_247);
or U489 (N_489,N_373,N_271);
nand U490 (N_490,N_295,N_290);
xor U491 (N_491,N_280,N_362);
nand U492 (N_492,N_259,N_214);
nand U493 (N_493,N_317,N_210);
nand U494 (N_494,N_298,N_323);
or U495 (N_495,N_379,N_219);
or U496 (N_496,N_238,N_278);
xnor U497 (N_497,N_391,N_320);
or U498 (N_498,N_304,N_273);
nor U499 (N_499,N_261,N_385);
or U500 (N_500,N_360,N_236);
xnor U501 (N_501,N_395,N_322);
nor U502 (N_502,N_337,N_247);
nor U503 (N_503,N_289,N_267);
or U504 (N_504,N_285,N_361);
and U505 (N_505,N_290,N_230);
nor U506 (N_506,N_301,N_398);
nor U507 (N_507,N_218,N_236);
nor U508 (N_508,N_251,N_283);
and U509 (N_509,N_266,N_259);
and U510 (N_510,N_317,N_339);
xnor U511 (N_511,N_217,N_290);
xnor U512 (N_512,N_295,N_345);
nor U513 (N_513,N_255,N_223);
nand U514 (N_514,N_219,N_359);
xnor U515 (N_515,N_335,N_204);
or U516 (N_516,N_320,N_229);
nor U517 (N_517,N_334,N_229);
or U518 (N_518,N_250,N_350);
nor U519 (N_519,N_210,N_376);
nand U520 (N_520,N_257,N_398);
nand U521 (N_521,N_278,N_300);
nor U522 (N_522,N_306,N_369);
and U523 (N_523,N_201,N_229);
and U524 (N_524,N_297,N_360);
xnor U525 (N_525,N_344,N_327);
xor U526 (N_526,N_259,N_324);
or U527 (N_527,N_282,N_379);
nand U528 (N_528,N_234,N_371);
nand U529 (N_529,N_339,N_233);
or U530 (N_530,N_300,N_294);
xor U531 (N_531,N_391,N_253);
xnor U532 (N_532,N_273,N_299);
or U533 (N_533,N_354,N_322);
or U534 (N_534,N_249,N_237);
or U535 (N_535,N_298,N_243);
nor U536 (N_536,N_206,N_360);
xor U537 (N_537,N_332,N_251);
xor U538 (N_538,N_287,N_372);
or U539 (N_539,N_382,N_367);
and U540 (N_540,N_291,N_386);
xor U541 (N_541,N_252,N_211);
or U542 (N_542,N_294,N_267);
or U543 (N_543,N_247,N_343);
xnor U544 (N_544,N_225,N_227);
or U545 (N_545,N_280,N_240);
or U546 (N_546,N_258,N_306);
or U547 (N_547,N_359,N_281);
and U548 (N_548,N_318,N_203);
or U549 (N_549,N_218,N_296);
and U550 (N_550,N_281,N_350);
nand U551 (N_551,N_200,N_258);
or U552 (N_552,N_357,N_265);
nor U553 (N_553,N_374,N_301);
nand U554 (N_554,N_369,N_360);
and U555 (N_555,N_216,N_295);
xnor U556 (N_556,N_363,N_223);
nand U557 (N_557,N_202,N_220);
xor U558 (N_558,N_202,N_262);
or U559 (N_559,N_202,N_320);
and U560 (N_560,N_259,N_346);
and U561 (N_561,N_223,N_210);
or U562 (N_562,N_384,N_212);
nand U563 (N_563,N_387,N_201);
and U564 (N_564,N_289,N_380);
nand U565 (N_565,N_282,N_384);
xor U566 (N_566,N_223,N_383);
or U567 (N_567,N_371,N_380);
or U568 (N_568,N_291,N_240);
xor U569 (N_569,N_275,N_297);
xnor U570 (N_570,N_370,N_357);
nand U571 (N_571,N_256,N_227);
nand U572 (N_572,N_227,N_239);
xor U573 (N_573,N_220,N_294);
nand U574 (N_574,N_374,N_273);
and U575 (N_575,N_309,N_297);
nor U576 (N_576,N_247,N_387);
xnor U577 (N_577,N_372,N_292);
xnor U578 (N_578,N_361,N_223);
or U579 (N_579,N_235,N_258);
xnor U580 (N_580,N_218,N_375);
and U581 (N_581,N_289,N_331);
nor U582 (N_582,N_246,N_306);
xor U583 (N_583,N_225,N_251);
nand U584 (N_584,N_264,N_384);
nor U585 (N_585,N_359,N_295);
or U586 (N_586,N_395,N_249);
or U587 (N_587,N_249,N_239);
and U588 (N_588,N_288,N_271);
nor U589 (N_589,N_243,N_257);
and U590 (N_590,N_372,N_274);
or U591 (N_591,N_259,N_307);
nand U592 (N_592,N_355,N_209);
nor U593 (N_593,N_245,N_354);
and U594 (N_594,N_240,N_290);
or U595 (N_595,N_379,N_373);
or U596 (N_596,N_215,N_295);
xnor U597 (N_597,N_216,N_247);
or U598 (N_598,N_351,N_210);
nand U599 (N_599,N_331,N_271);
xnor U600 (N_600,N_406,N_583);
nor U601 (N_601,N_504,N_509);
nor U602 (N_602,N_564,N_493);
nand U603 (N_603,N_586,N_405);
nor U604 (N_604,N_488,N_501);
xnor U605 (N_605,N_528,N_508);
or U606 (N_606,N_458,N_427);
or U607 (N_607,N_574,N_507);
and U608 (N_608,N_432,N_592);
nand U609 (N_609,N_527,N_510);
nand U610 (N_610,N_566,N_428);
xnor U611 (N_611,N_489,N_479);
or U612 (N_612,N_598,N_498);
and U613 (N_613,N_554,N_429);
nor U614 (N_614,N_518,N_536);
nor U615 (N_615,N_473,N_588);
xor U616 (N_616,N_469,N_494);
and U617 (N_617,N_578,N_459);
and U618 (N_618,N_419,N_539);
and U619 (N_619,N_475,N_482);
nand U620 (N_620,N_410,N_506);
or U621 (N_621,N_434,N_400);
xor U622 (N_622,N_495,N_579);
nor U623 (N_623,N_415,N_462);
or U624 (N_624,N_562,N_483);
nand U625 (N_625,N_572,N_446);
nor U626 (N_626,N_442,N_590);
or U627 (N_627,N_407,N_435);
nand U628 (N_628,N_521,N_550);
nor U629 (N_629,N_496,N_552);
nand U630 (N_630,N_546,N_532);
nor U631 (N_631,N_444,N_584);
nor U632 (N_632,N_457,N_481);
nand U633 (N_633,N_451,N_466);
xor U634 (N_634,N_557,N_471);
xor U635 (N_635,N_591,N_454);
and U636 (N_636,N_593,N_450);
xor U637 (N_637,N_412,N_478);
and U638 (N_638,N_447,N_487);
xor U639 (N_639,N_426,N_589);
and U640 (N_640,N_558,N_573);
xor U641 (N_641,N_570,N_548);
xnor U642 (N_642,N_575,N_505);
and U643 (N_643,N_499,N_549);
and U644 (N_644,N_438,N_533);
xnor U645 (N_645,N_571,N_529);
nand U646 (N_646,N_581,N_526);
and U647 (N_647,N_491,N_551);
nand U648 (N_648,N_561,N_514);
and U649 (N_649,N_404,N_472);
xor U650 (N_650,N_480,N_567);
and U651 (N_651,N_594,N_530);
xnor U652 (N_652,N_439,N_492);
or U653 (N_653,N_416,N_455);
nand U654 (N_654,N_534,N_547);
nand U655 (N_655,N_531,N_500);
xor U656 (N_656,N_461,N_467);
nand U657 (N_657,N_502,N_477);
nor U658 (N_658,N_585,N_409);
and U659 (N_659,N_420,N_587);
xnor U660 (N_660,N_470,N_555);
xnor U661 (N_661,N_453,N_443);
xor U662 (N_662,N_503,N_441);
nand U663 (N_663,N_541,N_417);
nor U664 (N_664,N_485,N_545);
or U665 (N_665,N_411,N_513);
xor U666 (N_666,N_595,N_456);
or U667 (N_667,N_452,N_497);
xnor U668 (N_668,N_544,N_413);
xor U669 (N_669,N_486,N_538);
and U670 (N_670,N_421,N_516);
xor U671 (N_671,N_474,N_484);
nor U672 (N_672,N_596,N_565);
xnor U673 (N_673,N_408,N_403);
or U674 (N_674,N_517,N_423);
nor U675 (N_675,N_568,N_464);
or U676 (N_676,N_597,N_511);
nand U677 (N_677,N_522,N_418);
or U678 (N_678,N_433,N_525);
or U679 (N_679,N_476,N_512);
and U680 (N_680,N_515,N_424);
or U681 (N_681,N_576,N_449);
and U682 (N_682,N_577,N_542);
or U683 (N_683,N_540,N_537);
nor U684 (N_684,N_580,N_520);
or U685 (N_685,N_448,N_556);
or U686 (N_686,N_582,N_440);
nor U687 (N_687,N_422,N_524);
nor U688 (N_688,N_543,N_425);
and U689 (N_689,N_563,N_569);
xnor U690 (N_690,N_401,N_465);
nor U691 (N_691,N_436,N_559);
nand U692 (N_692,N_519,N_523);
xor U693 (N_693,N_431,N_490);
nand U694 (N_694,N_460,N_414);
and U695 (N_695,N_402,N_463);
nor U696 (N_696,N_445,N_468);
nand U697 (N_697,N_553,N_535);
nand U698 (N_698,N_560,N_437);
or U699 (N_699,N_430,N_599);
nor U700 (N_700,N_460,N_405);
nand U701 (N_701,N_584,N_437);
and U702 (N_702,N_470,N_445);
or U703 (N_703,N_575,N_547);
or U704 (N_704,N_453,N_481);
xnor U705 (N_705,N_404,N_478);
or U706 (N_706,N_495,N_402);
nand U707 (N_707,N_485,N_585);
xor U708 (N_708,N_544,N_532);
and U709 (N_709,N_517,N_561);
or U710 (N_710,N_563,N_534);
nor U711 (N_711,N_426,N_560);
and U712 (N_712,N_509,N_517);
nor U713 (N_713,N_504,N_464);
or U714 (N_714,N_519,N_435);
and U715 (N_715,N_547,N_544);
and U716 (N_716,N_480,N_484);
nor U717 (N_717,N_470,N_506);
and U718 (N_718,N_562,N_593);
nand U719 (N_719,N_420,N_522);
nor U720 (N_720,N_434,N_513);
xnor U721 (N_721,N_463,N_492);
and U722 (N_722,N_577,N_498);
and U723 (N_723,N_594,N_591);
or U724 (N_724,N_520,N_446);
and U725 (N_725,N_557,N_523);
xor U726 (N_726,N_518,N_514);
or U727 (N_727,N_448,N_553);
and U728 (N_728,N_486,N_480);
nor U729 (N_729,N_425,N_539);
or U730 (N_730,N_501,N_549);
and U731 (N_731,N_421,N_402);
or U732 (N_732,N_483,N_484);
or U733 (N_733,N_540,N_556);
nand U734 (N_734,N_428,N_530);
nand U735 (N_735,N_571,N_568);
nor U736 (N_736,N_497,N_525);
and U737 (N_737,N_488,N_537);
and U738 (N_738,N_496,N_559);
or U739 (N_739,N_433,N_491);
and U740 (N_740,N_573,N_524);
and U741 (N_741,N_494,N_526);
xnor U742 (N_742,N_484,N_461);
nor U743 (N_743,N_578,N_473);
nand U744 (N_744,N_510,N_477);
nor U745 (N_745,N_498,N_516);
or U746 (N_746,N_439,N_532);
xor U747 (N_747,N_445,N_548);
nand U748 (N_748,N_545,N_458);
or U749 (N_749,N_490,N_552);
xnor U750 (N_750,N_496,N_551);
and U751 (N_751,N_536,N_559);
and U752 (N_752,N_409,N_559);
nor U753 (N_753,N_532,N_454);
nand U754 (N_754,N_548,N_550);
nand U755 (N_755,N_515,N_532);
xor U756 (N_756,N_488,N_466);
xor U757 (N_757,N_421,N_573);
and U758 (N_758,N_491,N_481);
nand U759 (N_759,N_435,N_438);
nor U760 (N_760,N_422,N_547);
nor U761 (N_761,N_554,N_538);
or U762 (N_762,N_437,N_578);
and U763 (N_763,N_544,N_519);
nor U764 (N_764,N_429,N_595);
nand U765 (N_765,N_543,N_404);
or U766 (N_766,N_592,N_452);
nor U767 (N_767,N_471,N_559);
nor U768 (N_768,N_474,N_460);
xnor U769 (N_769,N_481,N_436);
nand U770 (N_770,N_464,N_433);
and U771 (N_771,N_559,N_487);
nor U772 (N_772,N_506,N_468);
or U773 (N_773,N_582,N_519);
nor U774 (N_774,N_405,N_589);
nand U775 (N_775,N_503,N_567);
or U776 (N_776,N_517,N_593);
or U777 (N_777,N_520,N_425);
or U778 (N_778,N_531,N_476);
nand U779 (N_779,N_471,N_421);
or U780 (N_780,N_450,N_517);
xnor U781 (N_781,N_550,N_589);
nand U782 (N_782,N_584,N_428);
xor U783 (N_783,N_588,N_506);
or U784 (N_784,N_507,N_515);
nor U785 (N_785,N_490,N_520);
nand U786 (N_786,N_535,N_515);
xor U787 (N_787,N_429,N_523);
or U788 (N_788,N_453,N_527);
nand U789 (N_789,N_512,N_573);
nand U790 (N_790,N_517,N_476);
and U791 (N_791,N_471,N_508);
xnor U792 (N_792,N_503,N_564);
xnor U793 (N_793,N_447,N_417);
nand U794 (N_794,N_454,N_432);
or U795 (N_795,N_482,N_421);
and U796 (N_796,N_578,N_566);
or U797 (N_797,N_438,N_486);
xnor U798 (N_798,N_536,N_498);
and U799 (N_799,N_440,N_451);
nor U800 (N_800,N_608,N_775);
nor U801 (N_801,N_754,N_732);
and U802 (N_802,N_721,N_626);
xor U803 (N_803,N_793,N_679);
xnor U804 (N_804,N_644,N_717);
and U805 (N_805,N_785,N_733);
xnor U806 (N_806,N_718,N_791);
xnor U807 (N_807,N_629,N_604);
nor U808 (N_808,N_725,N_739);
and U809 (N_809,N_690,N_784);
nand U810 (N_810,N_705,N_702);
nor U811 (N_811,N_695,N_602);
xor U812 (N_812,N_688,N_756);
xor U813 (N_813,N_786,N_744);
and U814 (N_814,N_681,N_749);
xnor U815 (N_815,N_663,N_689);
nand U816 (N_816,N_704,N_646);
nand U817 (N_817,N_669,N_778);
or U818 (N_818,N_783,N_700);
xor U819 (N_819,N_710,N_694);
nor U820 (N_820,N_622,N_618);
nor U821 (N_821,N_649,N_781);
or U822 (N_822,N_790,N_737);
xor U823 (N_823,N_678,N_621);
nand U824 (N_824,N_730,N_788);
nand U825 (N_825,N_712,N_656);
xnor U826 (N_826,N_797,N_672);
or U827 (N_827,N_610,N_606);
or U828 (N_828,N_674,N_625);
nor U829 (N_829,N_600,N_643);
nor U830 (N_830,N_796,N_657);
or U831 (N_831,N_763,N_671);
nor U832 (N_832,N_627,N_652);
nor U833 (N_833,N_765,N_799);
nand U834 (N_834,N_740,N_697);
nor U835 (N_835,N_770,N_650);
nand U836 (N_836,N_738,N_758);
nand U837 (N_837,N_664,N_642);
and U838 (N_838,N_706,N_614);
nand U839 (N_839,N_611,N_624);
and U840 (N_840,N_773,N_637);
and U841 (N_841,N_728,N_794);
nor U842 (N_842,N_707,N_759);
nand U843 (N_843,N_751,N_632);
xnor U844 (N_844,N_641,N_683);
nor U845 (N_845,N_771,N_777);
xnor U846 (N_846,N_684,N_753);
nor U847 (N_847,N_722,N_693);
nor U848 (N_848,N_620,N_692);
nor U849 (N_849,N_743,N_605);
nand U850 (N_850,N_601,N_655);
and U851 (N_851,N_651,N_798);
nor U852 (N_852,N_701,N_768);
nand U853 (N_853,N_764,N_638);
xor U854 (N_854,N_731,N_667);
and U855 (N_855,N_660,N_619);
and U856 (N_856,N_760,N_680);
xor U857 (N_857,N_750,N_654);
nand U858 (N_858,N_696,N_699);
xnor U859 (N_859,N_726,N_691);
nand U860 (N_860,N_686,N_714);
xnor U861 (N_861,N_761,N_630);
nand U862 (N_862,N_742,N_616);
or U863 (N_863,N_787,N_780);
and U864 (N_864,N_716,N_727);
or U865 (N_865,N_746,N_673);
nor U866 (N_866,N_719,N_752);
or U867 (N_867,N_645,N_762);
or U868 (N_868,N_757,N_789);
nor U869 (N_869,N_617,N_748);
or U870 (N_870,N_635,N_665);
nor U871 (N_871,N_687,N_703);
or U872 (N_872,N_668,N_676);
nand U873 (N_873,N_747,N_607);
or U874 (N_874,N_698,N_767);
xor U875 (N_875,N_709,N_662);
nand U876 (N_876,N_772,N_711);
or U877 (N_877,N_774,N_659);
or U878 (N_878,N_658,N_735);
and U879 (N_879,N_782,N_685);
and U880 (N_880,N_708,N_628);
nor U881 (N_881,N_609,N_623);
or U882 (N_882,N_779,N_682);
and U883 (N_883,N_653,N_661);
or U884 (N_884,N_648,N_666);
nor U885 (N_885,N_729,N_639);
nand U886 (N_886,N_636,N_776);
or U887 (N_887,N_766,N_723);
nor U888 (N_888,N_633,N_640);
nor U889 (N_889,N_736,N_795);
or U890 (N_890,N_634,N_715);
nor U891 (N_891,N_745,N_631);
nor U892 (N_892,N_713,N_755);
xor U893 (N_893,N_615,N_612);
xor U894 (N_894,N_677,N_675);
nor U895 (N_895,N_724,N_670);
and U896 (N_896,N_603,N_769);
xnor U897 (N_897,N_613,N_720);
and U898 (N_898,N_647,N_734);
nand U899 (N_899,N_792,N_741);
or U900 (N_900,N_632,N_780);
or U901 (N_901,N_752,N_742);
nand U902 (N_902,N_681,N_777);
nor U903 (N_903,N_611,N_744);
nor U904 (N_904,N_654,N_670);
xnor U905 (N_905,N_636,N_718);
and U906 (N_906,N_668,N_784);
nand U907 (N_907,N_734,N_719);
or U908 (N_908,N_673,N_645);
or U909 (N_909,N_662,N_790);
nor U910 (N_910,N_678,N_697);
or U911 (N_911,N_732,N_658);
nor U912 (N_912,N_687,N_690);
nand U913 (N_913,N_613,N_787);
xor U914 (N_914,N_738,N_785);
and U915 (N_915,N_654,N_793);
xor U916 (N_916,N_714,N_705);
or U917 (N_917,N_789,N_675);
nor U918 (N_918,N_630,N_751);
xor U919 (N_919,N_623,N_676);
nor U920 (N_920,N_621,N_761);
or U921 (N_921,N_658,N_606);
or U922 (N_922,N_657,N_649);
or U923 (N_923,N_719,N_642);
or U924 (N_924,N_790,N_646);
or U925 (N_925,N_737,N_748);
nand U926 (N_926,N_753,N_794);
nor U927 (N_927,N_718,N_643);
nand U928 (N_928,N_674,N_744);
nand U929 (N_929,N_664,N_671);
and U930 (N_930,N_764,N_797);
xnor U931 (N_931,N_622,N_728);
nand U932 (N_932,N_654,N_743);
xor U933 (N_933,N_669,N_662);
nor U934 (N_934,N_615,N_711);
or U935 (N_935,N_742,N_710);
xor U936 (N_936,N_638,N_718);
nor U937 (N_937,N_710,N_724);
and U938 (N_938,N_619,N_736);
xnor U939 (N_939,N_635,N_626);
nand U940 (N_940,N_646,N_729);
or U941 (N_941,N_767,N_714);
or U942 (N_942,N_791,N_776);
or U943 (N_943,N_715,N_714);
nor U944 (N_944,N_764,N_706);
nand U945 (N_945,N_704,N_675);
nand U946 (N_946,N_603,N_621);
nor U947 (N_947,N_691,N_711);
nor U948 (N_948,N_695,N_643);
xor U949 (N_949,N_741,N_667);
nor U950 (N_950,N_738,N_765);
and U951 (N_951,N_790,N_601);
nor U952 (N_952,N_691,N_722);
xnor U953 (N_953,N_740,N_797);
xor U954 (N_954,N_604,N_683);
nand U955 (N_955,N_732,N_628);
xnor U956 (N_956,N_644,N_748);
nor U957 (N_957,N_641,N_677);
nand U958 (N_958,N_674,N_619);
nor U959 (N_959,N_720,N_770);
and U960 (N_960,N_761,N_794);
or U961 (N_961,N_794,N_747);
or U962 (N_962,N_730,N_611);
or U963 (N_963,N_787,N_639);
nand U964 (N_964,N_741,N_798);
nor U965 (N_965,N_617,N_649);
nand U966 (N_966,N_696,N_720);
and U967 (N_967,N_720,N_726);
nand U968 (N_968,N_644,N_690);
nor U969 (N_969,N_756,N_621);
nor U970 (N_970,N_659,N_604);
or U971 (N_971,N_716,N_776);
or U972 (N_972,N_725,N_642);
nand U973 (N_973,N_767,N_656);
nor U974 (N_974,N_676,N_775);
or U975 (N_975,N_764,N_782);
xnor U976 (N_976,N_734,N_690);
or U977 (N_977,N_692,N_608);
and U978 (N_978,N_664,N_726);
or U979 (N_979,N_756,N_691);
nor U980 (N_980,N_622,N_715);
nor U981 (N_981,N_668,N_769);
nand U982 (N_982,N_684,N_653);
nor U983 (N_983,N_774,N_710);
xnor U984 (N_984,N_635,N_780);
nor U985 (N_985,N_757,N_695);
xnor U986 (N_986,N_733,N_688);
nand U987 (N_987,N_789,N_659);
xnor U988 (N_988,N_704,N_709);
xor U989 (N_989,N_773,N_667);
xnor U990 (N_990,N_679,N_757);
xnor U991 (N_991,N_652,N_649);
and U992 (N_992,N_725,N_772);
xor U993 (N_993,N_784,N_666);
or U994 (N_994,N_636,N_694);
or U995 (N_995,N_793,N_708);
and U996 (N_996,N_683,N_650);
and U997 (N_997,N_746,N_694);
or U998 (N_998,N_734,N_602);
and U999 (N_999,N_741,N_745);
or U1000 (N_1000,N_801,N_966);
or U1001 (N_1001,N_811,N_907);
nor U1002 (N_1002,N_950,N_842);
and U1003 (N_1003,N_844,N_882);
xnor U1004 (N_1004,N_909,N_984);
or U1005 (N_1005,N_883,N_917);
or U1006 (N_1006,N_999,N_833);
nand U1007 (N_1007,N_873,N_805);
nor U1008 (N_1008,N_856,N_860);
xnor U1009 (N_1009,N_922,N_812);
or U1010 (N_1010,N_925,N_932);
nand U1011 (N_1011,N_910,N_979);
or U1012 (N_1012,N_946,N_924);
nand U1013 (N_1013,N_977,N_954);
nand U1014 (N_1014,N_978,N_821);
and U1015 (N_1015,N_852,N_838);
and U1016 (N_1016,N_847,N_969);
nor U1017 (N_1017,N_993,N_952);
nor U1018 (N_1018,N_964,N_988);
xor U1019 (N_1019,N_867,N_895);
or U1020 (N_1020,N_976,N_951);
nand U1021 (N_1021,N_850,N_937);
xnor U1022 (N_1022,N_918,N_904);
xor U1023 (N_1023,N_846,N_871);
nand U1024 (N_1024,N_959,N_906);
and U1025 (N_1025,N_935,N_949);
nand U1026 (N_1026,N_930,N_943);
nand U1027 (N_1027,N_898,N_824);
nor U1028 (N_1028,N_902,N_929);
xor U1029 (N_1029,N_896,N_859);
nor U1030 (N_1030,N_986,N_914);
xor U1031 (N_1031,N_862,N_828);
nand U1032 (N_1032,N_920,N_884);
nor U1033 (N_1033,N_853,N_928);
or U1034 (N_1034,N_939,N_972);
or U1035 (N_1035,N_848,N_897);
xnor U1036 (N_1036,N_879,N_892);
xor U1037 (N_1037,N_835,N_877);
and U1038 (N_1038,N_894,N_820);
nand U1039 (N_1039,N_815,N_938);
and U1040 (N_1040,N_825,N_818);
nor U1041 (N_1041,N_840,N_822);
nand U1042 (N_1042,N_921,N_890);
nand U1043 (N_1043,N_916,N_983);
nor U1044 (N_1044,N_970,N_900);
xnor U1045 (N_1045,N_808,N_899);
or U1046 (N_1046,N_913,N_989);
and U1047 (N_1047,N_807,N_885);
nor U1048 (N_1048,N_868,N_886);
nand U1049 (N_1049,N_874,N_936);
nand U1050 (N_1050,N_870,N_905);
and U1051 (N_1051,N_995,N_948);
or U1052 (N_1052,N_962,N_875);
xnor U1053 (N_1053,N_934,N_987);
and U1054 (N_1054,N_931,N_804);
xnor U1055 (N_1055,N_891,N_857);
nand U1056 (N_1056,N_827,N_958);
nand U1057 (N_1057,N_841,N_947);
nor U1058 (N_1058,N_854,N_830);
or U1059 (N_1059,N_865,N_861);
nand U1060 (N_1060,N_887,N_814);
and U1061 (N_1061,N_982,N_802);
and U1062 (N_1062,N_869,N_927);
or U1063 (N_1063,N_961,N_863);
xnor U1064 (N_1064,N_911,N_965);
nor U1065 (N_1065,N_858,N_919);
or U1066 (N_1066,N_888,N_994);
nand U1067 (N_1067,N_998,N_834);
and U1068 (N_1068,N_876,N_878);
or U1069 (N_1069,N_880,N_809);
xnor U1070 (N_1070,N_960,N_851);
nor U1071 (N_1071,N_893,N_800);
xor U1072 (N_1072,N_985,N_941);
nor U1073 (N_1073,N_992,N_832);
or U1074 (N_1074,N_971,N_849);
nor U1075 (N_1075,N_975,N_903);
or U1076 (N_1076,N_819,N_837);
nand U1077 (N_1077,N_945,N_956);
nand U1078 (N_1078,N_940,N_901);
nand U1079 (N_1079,N_967,N_803);
xor U1080 (N_1080,N_806,N_817);
xnor U1081 (N_1081,N_926,N_881);
or U1082 (N_1082,N_855,N_839);
nor U1083 (N_1083,N_963,N_912);
nand U1084 (N_1084,N_974,N_944);
or U1085 (N_1085,N_990,N_968);
nor U1086 (N_1086,N_831,N_889);
nand U1087 (N_1087,N_953,N_872);
nand U1088 (N_1088,N_973,N_816);
nor U1089 (N_1089,N_908,N_810);
or U1090 (N_1090,N_933,N_923);
xnor U1091 (N_1091,N_845,N_981);
nor U1092 (N_1092,N_826,N_997);
nor U1093 (N_1093,N_866,N_843);
and U1094 (N_1094,N_957,N_955);
or U1095 (N_1095,N_942,N_996);
nand U1096 (N_1096,N_813,N_864);
xnor U1097 (N_1097,N_991,N_915);
nor U1098 (N_1098,N_980,N_829);
xnor U1099 (N_1099,N_836,N_823);
and U1100 (N_1100,N_977,N_971);
and U1101 (N_1101,N_840,N_817);
nor U1102 (N_1102,N_855,N_853);
nor U1103 (N_1103,N_908,N_895);
nor U1104 (N_1104,N_877,N_812);
nand U1105 (N_1105,N_862,N_963);
or U1106 (N_1106,N_819,N_979);
and U1107 (N_1107,N_893,N_806);
xnor U1108 (N_1108,N_823,N_888);
nor U1109 (N_1109,N_830,N_958);
nor U1110 (N_1110,N_896,N_900);
and U1111 (N_1111,N_867,N_959);
or U1112 (N_1112,N_881,N_876);
or U1113 (N_1113,N_979,N_820);
nor U1114 (N_1114,N_911,N_950);
and U1115 (N_1115,N_913,N_822);
xnor U1116 (N_1116,N_938,N_963);
or U1117 (N_1117,N_821,N_924);
and U1118 (N_1118,N_934,N_817);
nor U1119 (N_1119,N_930,N_879);
xnor U1120 (N_1120,N_966,N_807);
nand U1121 (N_1121,N_985,N_997);
and U1122 (N_1122,N_982,N_852);
or U1123 (N_1123,N_924,N_819);
nand U1124 (N_1124,N_854,N_866);
and U1125 (N_1125,N_837,N_881);
xor U1126 (N_1126,N_906,N_953);
nand U1127 (N_1127,N_948,N_938);
and U1128 (N_1128,N_972,N_863);
nand U1129 (N_1129,N_838,N_937);
and U1130 (N_1130,N_890,N_869);
or U1131 (N_1131,N_852,N_843);
and U1132 (N_1132,N_977,N_985);
xnor U1133 (N_1133,N_873,N_966);
nor U1134 (N_1134,N_829,N_828);
nand U1135 (N_1135,N_851,N_874);
or U1136 (N_1136,N_895,N_869);
and U1137 (N_1137,N_968,N_889);
xnor U1138 (N_1138,N_906,N_875);
nand U1139 (N_1139,N_978,N_828);
and U1140 (N_1140,N_918,N_917);
nor U1141 (N_1141,N_821,N_919);
xor U1142 (N_1142,N_933,N_997);
or U1143 (N_1143,N_907,N_823);
and U1144 (N_1144,N_968,N_838);
nand U1145 (N_1145,N_881,N_842);
nor U1146 (N_1146,N_968,N_880);
or U1147 (N_1147,N_968,N_957);
nand U1148 (N_1148,N_898,N_935);
nor U1149 (N_1149,N_813,N_960);
and U1150 (N_1150,N_934,N_812);
nor U1151 (N_1151,N_853,N_877);
or U1152 (N_1152,N_929,N_999);
and U1153 (N_1153,N_865,N_883);
and U1154 (N_1154,N_949,N_840);
nand U1155 (N_1155,N_994,N_968);
or U1156 (N_1156,N_971,N_935);
nand U1157 (N_1157,N_918,N_833);
nor U1158 (N_1158,N_875,N_863);
and U1159 (N_1159,N_967,N_930);
xor U1160 (N_1160,N_964,N_926);
and U1161 (N_1161,N_823,N_806);
nor U1162 (N_1162,N_954,N_941);
and U1163 (N_1163,N_986,N_907);
nand U1164 (N_1164,N_810,N_873);
nand U1165 (N_1165,N_914,N_895);
nand U1166 (N_1166,N_849,N_870);
nor U1167 (N_1167,N_822,N_914);
xnor U1168 (N_1168,N_907,N_894);
xnor U1169 (N_1169,N_837,N_948);
nand U1170 (N_1170,N_943,N_993);
xnor U1171 (N_1171,N_958,N_889);
xor U1172 (N_1172,N_849,N_819);
xor U1173 (N_1173,N_842,N_990);
nand U1174 (N_1174,N_818,N_831);
nand U1175 (N_1175,N_877,N_982);
nor U1176 (N_1176,N_962,N_837);
nor U1177 (N_1177,N_890,N_889);
xor U1178 (N_1178,N_985,N_827);
nand U1179 (N_1179,N_936,N_900);
nor U1180 (N_1180,N_922,N_958);
nor U1181 (N_1181,N_829,N_905);
or U1182 (N_1182,N_860,N_886);
nand U1183 (N_1183,N_826,N_875);
nand U1184 (N_1184,N_811,N_968);
nor U1185 (N_1185,N_889,N_995);
or U1186 (N_1186,N_984,N_920);
and U1187 (N_1187,N_832,N_819);
or U1188 (N_1188,N_826,N_921);
and U1189 (N_1189,N_872,N_886);
nand U1190 (N_1190,N_905,N_917);
nor U1191 (N_1191,N_812,N_830);
and U1192 (N_1192,N_932,N_816);
nand U1193 (N_1193,N_800,N_880);
xor U1194 (N_1194,N_998,N_822);
nand U1195 (N_1195,N_889,N_988);
and U1196 (N_1196,N_888,N_835);
or U1197 (N_1197,N_846,N_832);
xor U1198 (N_1198,N_995,N_941);
nand U1199 (N_1199,N_976,N_903);
or U1200 (N_1200,N_1148,N_1016);
nor U1201 (N_1201,N_1163,N_1146);
and U1202 (N_1202,N_1137,N_1097);
nand U1203 (N_1203,N_1076,N_1136);
nor U1204 (N_1204,N_1021,N_1064);
and U1205 (N_1205,N_1145,N_1094);
or U1206 (N_1206,N_1167,N_1014);
xnor U1207 (N_1207,N_1179,N_1173);
xor U1208 (N_1208,N_1074,N_1026);
nand U1209 (N_1209,N_1098,N_1010);
and U1210 (N_1210,N_1170,N_1030);
nor U1211 (N_1211,N_1000,N_1187);
nand U1212 (N_1212,N_1154,N_1195);
or U1213 (N_1213,N_1180,N_1058);
or U1214 (N_1214,N_1156,N_1194);
or U1215 (N_1215,N_1018,N_1055);
nor U1216 (N_1216,N_1034,N_1035);
nand U1217 (N_1217,N_1158,N_1181);
nand U1218 (N_1218,N_1183,N_1114);
or U1219 (N_1219,N_1106,N_1117);
xor U1220 (N_1220,N_1066,N_1073);
nor U1221 (N_1221,N_1001,N_1025);
nand U1222 (N_1222,N_1006,N_1165);
nor U1223 (N_1223,N_1063,N_1152);
or U1224 (N_1224,N_1123,N_1115);
nor U1225 (N_1225,N_1157,N_1101);
nor U1226 (N_1226,N_1088,N_1028);
and U1227 (N_1227,N_1056,N_1083);
nand U1228 (N_1228,N_1011,N_1038);
nand U1229 (N_1229,N_1048,N_1050);
and U1230 (N_1230,N_1060,N_1081);
or U1231 (N_1231,N_1189,N_1052);
xor U1232 (N_1232,N_1119,N_1171);
nor U1233 (N_1233,N_1082,N_1109);
or U1234 (N_1234,N_1015,N_1140);
nor U1235 (N_1235,N_1144,N_1032);
nand U1236 (N_1236,N_1040,N_1182);
or U1237 (N_1237,N_1107,N_1031);
nand U1238 (N_1238,N_1022,N_1166);
or U1239 (N_1239,N_1044,N_1139);
nand U1240 (N_1240,N_1005,N_1065);
xnor U1241 (N_1241,N_1135,N_1104);
nor U1242 (N_1242,N_1150,N_1147);
and U1243 (N_1243,N_1077,N_1124);
xor U1244 (N_1244,N_1009,N_1125);
nor U1245 (N_1245,N_1199,N_1057);
or U1246 (N_1246,N_1142,N_1113);
or U1247 (N_1247,N_1196,N_1069);
nand U1248 (N_1248,N_1037,N_1129);
nor U1249 (N_1249,N_1062,N_1095);
and U1250 (N_1250,N_1185,N_1138);
and U1251 (N_1251,N_1086,N_1085);
nor U1252 (N_1252,N_1174,N_1169);
nor U1253 (N_1253,N_1079,N_1061);
and U1254 (N_1254,N_1177,N_1188);
xnor U1255 (N_1255,N_1121,N_1153);
nor U1256 (N_1256,N_1172,N_1127);
xor U1257 (N_1257,N_1023,N_1004);
and U1258 (N_1258,N_1143,N_1036);
and U1259 (N_1259,N_1007,N_1013);
or U1260 (N_1260,N_1161,N_1134);
and U1261 (N_1261,N_1111,N_1198);
nor U1262 (N_1262,N_1017,N_1133);
nor U1263 (N_1263,N_1116,N_1197);
nand U1264 (N_1264,N_1108,N_1002);
nor U1265 (N_1265,N_1175,N_1128);
or U1266 (N_1266,N_1184,N_1049);
nor U1267 (N_1267,N_1019,N_1042);
xor U1268 (N_1268,N_1100,N_1008);
nor U1269 (N_1269,N_1029,N_1103);
xnor U1270 (N_1270,N_1084,N_1132);
nor U1271 (N_1271,N_1054,N_1168);
nand U1272 (N_1272,N_1155,N_1162);
and U1273 (N_1273,N_1047,N_1039);
and U1274 (N_1274,N_1024,N_1122);
or U1275 (N_1275,N_1093,N_1012);
nor U1276 (N_1276,N_1091,N_1003);
xor U1277 (N_1277,N_1176,N_1130);
and U1278 (N_1278,N_1059,N_1164);
and U1279 (N_1279,N_1092,N_1099);
nor U1280 (N_1280,N_1033,N_1051);
or U1281 (N_1281,N_1105,N_1078);
nand U1282 (N_1282,N_1141,N_1112);
xor U1283 (N_1283,N_1193,N_1159);
nor U1284 (N_1284,N_1071,N_1149);
or U1285 (N_1285,N_1178,N_1053);
nor U1286 (N_1286,N_1043,N_1110);
nand U1287 (N_1287,N_1090,N_1120);
xnor U1288 (N_1288,N_1041,N_1131);
and U1289 (N_1289,N_1046,N_1045);
nand U1290 (N_1290,N_1072,N_1027);
and U1291 (N_1291,N_1186,N_1096);
or U1292 (N_1292,N_1089,N_1191);
nor U1293 (N_1293,N_1087,N_1080);
or U1294 (N_1294,N_1118,N_1192);
or U1295 (N_1295,N_1160,N_1190);
xor U1296 (N_1296,N_1151,N_1126);
nand U1297 (N_1297,N_1075,N_1102);
xnor U1298 (N_1298,N_1020,N_1068);
nor U1299 (N_1299,N_1070,N_1067);
xor U1300 (N_1300,N_1131,N_1120);
xnor U1301 (N_1301,N_1156,N_1176);
nand U1302 (N_1302,N_1115,N_1110);
or U1303 (N_1303,N_1018,N_1120);
or U1304 (N_1304,N_1160,N_1047);
nand U1305 (N_1305,N_1079,N_1008);
nand U1306 (N_1306,N_1195,N_1171);
nor U1307 (N_1307,N_1104,N_1136);
nand U1308 (N_1308,N_1010,N_1127);
xor U1309 (N_1309,N_1107,N_1032);
nor U1310 (N_1310,N_1012,N_1109);
nand U1311 (N_1311,N_1029,N_1133);
and U1312 (N_1312,N_1135,N_1074);
or U1313 (N_1313,N_1079,N_1125);
or U1314 (N_1314,N_1069,N_1067);
nor U1315 (N_1315,N_1003,N_1189);
or U1316 (N_1316,N_1119,N_1052);
and U1317 (N_1317,N_1023,N_1033);
nand U1318 (N_1318,N_1054,N_1104);
or U1319 (N_1319,N_1190,N_1076);
xnor U1320 (N_1320,N_1072,N_1116);
and U1321 (N_1321,N_1074,N_1165);
and U1322 (N_1322,N_1085,N_1018);
xor U1323 (N_1323,N_1084,N_1064);
and U1324 (N_1324,N_1170,N_1126);
nor U1325 (N_1325,N_1060,N_1003);
or U1326 (N_1326,N_1132,N_1163);
and U1327 (N_1327,N_1115,N_1192);
nand U1328 (N_1328,N_1196,N_1113);
nor U1329 (N_1329,N_1160,N_1040);
nand U1330 (N_1330,N_1156,N_1081);
xnor U1331 (N_1331,N_1099,N_1036);
or U1332 (N_1332,N_1119,N_1025);
nand U1333 (N_1333,N_1053,N_1079);
and U1334 (N_1334,N_1199,N_1110);
nor U1335 (N_1335,N_1048,N_1006);
nand U1336 (N_1336,N_1135,N_1152);
nand U1337 (N_1337,N_1103,N_1150);
or U1338 (N_1338,N_1098,N_1174);
xor U1339 (N_1339,N_1172,N_1085);
nand U1340 (N_1340,N_1043,N_1006);
xnor U1341 (N_1341,N_1059,N_1049);
xor U1342 (N_1342,N_1112,N_1065);
nor U1343 (N_1343,N_1146,N_1085);
nor U1344 (N_1344,N_1142,N_1080);
or U1345 (N_1345,N_1194,N_1033);
and U1346 (N_1346,N_1102,N_1171);
nand U1347 (N_1347,N_1057,N_1116);
nor U1348 (N_1348,N_1085,N_1108);
or U1349 (N_1349,N_1150,N_1163);
xor U1350 (N_1350,N_1151,N_1018);
xor U1351 (N_1351,N_1185,N_1122);
nand U1352 (N_1352,N_1032,N_1163);
nand U1353 (N_1353,N_1013,N_1138);
nor U1354 (N_1354,N_1130,N_1154);
xor U1355 (N_1355,N_1053,N_1133);
xor U1356 (N_1356,N_1191,N_1048);
or U1357 (N_1357,N_1035,N_1170);
xnor U1358 (N_1358,N_1040,N_1028);
xnor U1359 (N_1359,N_1105,N_1000);
xnor U1360 (N_1360,N_1138,N_1001);
xnor U1361 (N_1361,N_1063,N_1078);
or U1362 (N_1362,N_1117,N_1052);
nand U1363 (N_1363,N_1192,N_1013);
or U1364 (N_1364,N_1005,N_1019);
or U1365 (N_1365,N_1100,N_1054);
and U1366 (N_1366,N_1192,N_1189);
and U1367 (N_1367,N_1014,N_1059);
nor U1368 (N_1368,N_1078,N_1053);
nor U1369 (N_1369,N_1195,N_1081);
xnor U1370 (N_1370,N_1101,N_1021);
and U1371 (N_1371,N_1039,N_1050);
nor U1372 (N_1372,N_1092,N_1093);
or U1373 (N_1373,N_1056,N_1191);
xnor U1374 (N_1374,N_1146,N_1060);
xnor U1375 (N_1375,N_1058,N_1162);
or U1376 (N_1376,N_1067,N_1004);
or U1377 (N_1377,N_1082,N_1085);
and U1378 (N_1378,N_1182,N_1013);
or U1379 (N_1379,N_1023,N_1002);
or U1380 (N_1380,N_1110,N_1154);
xor U1381 (N_1381,N_1159,N_1047);
nand U1382 (N_1382,N_1178,N_1192);
nor U1383 (N_1383,N_1129,N_1036);
xor U1384 (N_1384,N_1137,N_1109);
or U1385 (N_1385,N_1193,N_1107);
or U1386 (N_1386,N_1044,N_1010);
and U1387 (N_1387,N_1143,N_1110);
and U1388 (N_1388,N_1103,N_1030);
xor U1389 (N_1389,N_1126,N_1005);
nor U1390 (N_1390,N_1040,N_1143);
nor U1391 (N_1391,N_1017,N_1009);
nor U1392 (N_1392,N_1035,N_1129);
nor U1393 (N_1393,N_1085,N_1196);
or U1394 (N_1394,N_1078,N_1114);
xor U1395 (N_1395,N_1037,N_1066);
nor U1396 (N_1396,N_1034,N_1183);
nor U1397 (N_1397,N_1001,N_1174);
or U1398 (N_1398,N_1054,N_1199);
nor U1399 (N_1399,N_1156,N_1187);
xnor U1400 (N_1400,N_1314,N_1301);
nand U1401 (N_1401,N_1380,N_1322);
and U1402 (N_1402,N_1254,N_1331);
xor U1403 (N_1403,N_1206,N_1205);
nor U1404 (N_1404,N_1283,N_1368);
or U1405 (N_1405,N_1366,N_1381);
or U1406 (N_1406,N_1327,N_1256);
and U1407 (N_1407,N_1321,N_1232);
nor U1408 (N_1408,N_1284,N_1318);
xnor U1409 (N_1409,N_1388,N_1377);
and U1410 (N_1410,N_1278,N_1299);
or U1411 (N_1411,N_1364,N_1297);
nor U1412 (N_1412,N_1204,N_1213);
or U1413 (N_1413,N_1371,N_1344);
and U1414 (N_1414,N_1326,N_1243);
nand U1415 (N_1415,N_1212,N_1316);
nor U1416 (N_1416,N_1233,N_1295);
nand U1417 (N_1417,N_1348,N_1202);
or U1418 (N_1418,N_1290,N_1208);
or U1419 (N_1419,N_1245,N_1216);
and U1420 (N_1420,N_1241,N_1360);
and U1421 (N_1421,N_1385,N_1308);
or U1422 (N_1422,N_1200,N_1319);
nand U1423 (N_1423,N_1342,N_1221);
and U1424 (N_1424,N_1207,N_1305);
nand U1425 (N_1425,N_1210,N_1333);
nor U1426 (N_1426,N_1337,N_1362);
and U1427 (N_1427,N_1332,N_1230);
nor U1428 (N_1428,N_1335,N_1397);
xor U1429 (N_1429,N_1357,N_1261);
or U1430 (N_1430,N_1272,N_1279);
nand U1431 (N_1431,N_1258,N_1323);
nand U1432 (N_1432,N_1235,N_1373);
or U1433 (N_1433,N_1352,N_1359);
xnor U1434 (N_1434,N_1236,N_1361);
nor U1435 (N_1435,N_1265,N_1351);
or U1436 (N_1436,N_1383,N_1292);
and U1437 (N_1437,N_1238,N_1313);
or U1438 (N_1438,N_1363,N_1345);
nor U1439 (N_1439,N_1274,N_1334);
xor U1440 (N_1440,N_1281,N_1309);
and U1441 (N_1441,N_1220,N_1294);
nor U1442 (N_1442,N_1240,N_1382);
or U1443 (N_1443,N_1250,N_1311);
or U1444 (N_1444,N_1237,N_1307);
and U1445 (N_1445,N_1354,N_1339);
nor U1446 (N_1446,N_1253,N_1346);
nor U1447 (N_1447,N_1289,N_1248);
nand U1448 (N_1448,N_1328,N_1214);
nor U1449 (N_1449,N_1217,N_1262);
nand U1450 (N_1450,N_1277,N_1276);
or U1451 (N_1451,N_1247,N_1387);
nand U1452 (N_1452,N_1201,N_1365);
or U1453 (N_1453,N_1280,N_1251);
nor U1454 (N_1454,N_1341,N_1264);
nand U1455 (N_1455,N_1392,N_1255);
nand U1456 (N_1456,N_1367,N_1347);
nand U1457 (N_1457,N_1288,N_1209);
and U1458 (N_1458,N_1399,N_1393);
or U1459 (N_1459,N_1229,N_1390);
or U1460 (N_1460,N_1325,N_1350);
nor U1461 (N_1461,N_1302,N_1372);
nor U1462 (N_1462,N_1394,N_1315);
or U1463 (N_1463,N_1374,N_1376);
nor U1464 (N_1464,N_1239,N_1343);
and U1465 (N_1465,N_1222,N_1267);
nor U1466 (N_1466,N_1203,N_1231);
nor U1467 (N_1467,N_1353,N_1268);
xor U1468 (N_1468,N_1398,N_1211);
or U1469 (N_1469,N_1270,N_1225);
xnor U1470 (N_1470,N_1396,N_1273);
nor U1471 (N_1471,N_1293,N_1330);
xnor U1472 (N_1472,N_1215,N_1375);
and U1473 (N_1473,N_1244,N_1349);
or U1474 (N_1474,N_1298,N_1338);
or U1475 (N_1475,N_1355,N_1304);
and U1476 (N_1476,N_1324,N_1356);
nor U1477 (N_1477,N_1291,N_1306);
and U1478 (N_1478,N_1246,N_1227);
nand U1479 (N_1479,N_1389,N_1219);
nand U1480 (N_1480,N_1358,N_1226);
and U1481 (N_1481,N_1310,N_1263);
nand U1482 (N_1482,N_1391,N_1257);
or U1483 (N_1483,N_1300,N_1218);
xor U1484 (N_1484,N_1296,N_1260);
xor U1485 (N_1485,N_1287,N_1259);
nand U1486 (N_1486,N_1303,N_1275);
or U1487 (N_1487,N_1285,N_1378);
or U1488 (N_1488,N_1320,N_1317);
or U1489 (N_1489,N_1340,N_1271);
xor U1490 (N_1490,N_1369,N_1269);
nand U1491 (N_1491,N_1223,N_1234);
nor U1492 (N_1492,N_1384,N_1329);
nand U1493 (N_1493,N_1312,N_1282);
xor U1494 (N_1494,N_1395,N_1242);
nand U1495 (N_1495,N_1224,N_1266);
or U1496 (N_1496,N_1379,N_1370);
or U1497 (N_1497,N_1252,N_1228);
and U1498 (N_1498,N_1386,N_1249);
or U1499 (N_1499,N_1336,N_1286);
nand U1500 (N_1500,N_1214,N_1230);
nor U1501 (N_1501,N_1232,N_1331);
or U1502 (N_1502,N_1288,N_1262);
xor U1503 (N_1503,N_1369,N_1324);
xor U1504 (N_1504,N_1374,N_1200);
nor U1505 (N_1505,N_1268,N_1229);
and U1506 (N_1506,N_1383,N_1244);
xnor U1507 (N_1507,N_1267,N_1250);
xnor U1508 (N_1508,N_1339,N_1220);
or U1509 (N_1509,N_1357,N_1291);
nand U1510 (N_1510,N_1343,N_1219);
and U1511 (N_1511,N_1341,N_1382);
and U1512 (N_1512,N_1388,N_1284);
xnor U1513 (N_1513,N_1281,N_1320);
or U1514 (N_1514,N_1271,N_1343);
and U1515 (N_1515,N_1200,N_1281);
nand U1516 (N_1516,N_1332,N_1327);
or U1517 (N_1517,N_1379,N_1286);
and U1518 (N_1518,N_1303,N_1377);
and U1519 (N_1519,N_1307,N_1346);
or U1520 (N_1520,N_1396,N_1287);
xor U1521 (N_1521,N_1208,N_1253);
nand U1522 (N_1522,N_1227,N_1244);
and U1523 (N_1523,N_1375,N_1316);
nor U1524 (N_1524,N_1310,N_1228);
or U1525 (N_1525,N_1247,N_1318);
and U1526 (N_1526,N_1313,N_1369);
nor U1527 (N_1527,N_1353,N_1256);
nand U1528 (N_1528,N_1210,N_1271);
xor U1529 (N_1529,N_1210,N_1285);
xor U1530 (N_1530,N_1317,N_1329);
or U1531 (N_1531,N_1339,N_1301);
xor U1532 (N_1532,N_1364,N_1368);
or U1533 (N_1533,N_1385,N_1378);
or U1534 (N_1534,N_1393,N_1210);
nand U1535 (N_1535,N_1204,N_1242);
or U1536 (N_1536,N_1290,N_1387);
or U1537 (N_1537,N_1350,N_1310);
nand U1538 (N_1538,N_1218,N_1319);
and U1539 (N_1539,N_1298,N_1345);
and U1540 (N_1540,N_1373,N_1362);
nand U1541 (N_1541,N_1385,N_1334);
nor U1542 (N_1542,N_1223,N_1388);
nand U1543 (N_1543,N_1234,N_1249);
nand U1544 (N_1544,N_1328,N_1226);
nand U1545 (N_1545,N_1273,N_1257);
nor U1546 (N_1546,N_1269,N_1394);
nor U1547 (N_1547,N_1376,N_1318);
xnor U1548 (N_1548,N_1255,N_1382);
nand U1549 (N_1549,N_1312,N_1324);
nor U1550 (N_1550,N_1317,N_1284);
xnor U1551 (N_1551,N_1239,N_1268);
xor U1552 (N_1552,N_1313,N_1305);
and U1553 (N_1553,N_1219,N_1393);
or U1554 (N_1554,N_1210,N_1361);
or U1555 (N_1555,N_1335,N_1398);
or U1556 (N_1556,N_1393,N_1267);
and U1557 (N_1557,N_1260,N_1338);
nor U1558 (N_1558,N_1324,N_1374);
xor U1559 (N_1559,N_1362,N_1385);
and U1560 (N_1560,N_1382,N_1228);
xnor U1561 (N_1561,N_1355,N_1261);
nand U1562 (N_1562,N_1338,N_1304);
xor U1563 (N_1563,N_1246,N_1357);
xor U1564 (N_1564,N_1326,N_1298);
and U1565 (N_1565,N_1257,N_1231);
or U1566 (N_1566,N_1234,N_1241);
and U1567 (N_1567,N_1290,N_1310);
nand U1568 (N_1568,N_1250,N_1392);
or U1569 (N_1569,N_1241,N_1320);
and U1570 (N_1570,N_1353,N_1392);
nand U1571 (N_1571,N_1264,N_1270);
and U1572 (N_1572,N_1300,N_1302);
nand U1573 (N_1573,N_1242,N_1309);
xor U1574 (N_1574,N_1365,N_1252);
or U1575 (N_1575,N_1306,N_1333);
xor U1576 (N_1576,N_1365,N_1373);
nand U1577 (N_1577,N_1256,N_1246);
xnor U1578 (N_1578,N_1399,N_1383);
xnor U1579 (N_1579,N_1247,N_1377);
nor U1580 (N_1580,N_1351,N_1287);
or U1581 (N_1581,N_1281,N_1262);
nor U1582 (N_1582,N_1340,N_1384);
nor U1583 (N_1583,N_1287,N_1352);
and U1584 (N_1584,N_1366,N_1279);
nor U1585 (N_1585,N_1364,N_1218);
xor U1586 (N_1586,N_1340,N_1233);
nand U1587 (N_1587,N_1347,N_1321);
and U1588 (N_1588,N_1292,N_1319);
nor U1589 (N_1589,N_1377,N_1385);
and U1590 (N_1590,N_1397,N_1228);
and U1591 (N_1591,N_1308,N_1351);
xor U1592 (N_1592,N_1302,N_1228);
xor U1593 (N_1593,N_1215,N_1354);
nor U1594 (N_1594,N_1356,N_1311);
xor U1595 (N_1595,N_1350,N_1233);
and U1596 (N_1596,N_1215,N_1369);
nor U1597 (N_1597,N_1201,N_1312);
xor U1598 (N_1598,N_1252,N_1216);
nand U1599 (N_1599,N_1397,N_1262);
and U1600 (N_1600,N_1547,N_1536);
nand U1601 (N_1601,N_1521,N_1434);
or U1602 (N_1602,N_1466,N_1431);
and U1603 (N_1603,N_1563,N_1472);
nor U1604 (N_1604,N_1576,N_1533);
nand U1605 (N_1605,N_1426,N_1528);
xnor U1606 (N_1606,N_1580,N_1441);
and U1607 (N_1607,N_1428,N_1541);
nand U1608 (N_1608,N_1475,N_1575);
nand U1609 (N_1609,N_1566,N_1438);
nor U1610 (N_1610,N_1482,N_1476);
nor U1611 (N_1611,N_1499,N_1460);
and U1612 (N_1612,N_1500,N_1411);
nand U1613 (N_1613,N_1561,N_1590);
xnor U1614 (N_1614,N_1595,N_1435);
nor U1615 (N_1615,N_1458,N_1470);
nor U1616 (N_1616,N_1490,N_1456);
and U1617 (N_1617,N_1447,N_1542);
nand U1618 (N_1618,N_1425,N_1504);
xor U1619 (N_1619,N_1584,N_1468);
xor U1620 (N_1620,N_1400,N_1488);
or U1621 (N_1621,N_1571,N_1556);
and U1622 (N_1622,N_1477,N_1577);
nand U1623 (N_1623,N_1471,N_1424);
nand U1624 (N_1624,N_1495,N_1529);
or U1625 (N_1625,N_1493,N_1506);
nand U1626 (N_1626,N_1420,N_1513);
and U1627 (N_1627,N_1519,N_1502);
or U1628 (N_1628,N_1412,N_1432);
or U1629 (N_1629,N_1419,N_1474);
or U1630 (N_1630,N_1473,N_1484);
nand U1631 (N_1631,N_1544,N_1408);
or U1632 (N_1632,N_1436,N_1594);
xnor U1633 (N_1633,N_1537,N_1463);
and U1634 (N_1634,N_1546,N_1581);
and U1635 (N_1635,N_1596,N_1453);
and U1636 (N_1636,N_1481,N_1559);
nand U1637 (N_1637,N_1413,N_1509);
nand U1638 (N_1638,N_1457,N_1443);
nor U1639 (N_1639,N_1440,N_1496);
nor U1640 (N_1640,N_1416,N_1538);
nor U1641 (N_1641,N_1406,N_1491);
or U1642 (N_1642,N_1409,N_1508);
and U1643 (N_1643,N_1564,N_1540);
or U1644 (N_1644,N_1497,N_1422);
and U1645 (N_1645,N_1524,N_1445);
xnor U1646 (N_1646,N_1573,N_1557);
nand U1647 (N_1647,N_1478,N_1514);
and U1648 (N_1648,N_1523,N_1585);
nor U1649 (N_1649,N_1515,N_1574);
nor U1650 (N_1650,N_1592,N_1427);
nor U1651 (N_1651,N_1492,N_1589);
or U1652 (N_1652,N_1461,N_1516);
or U1653 (N_1653,N_1505,N_1593);
nor U1654 (N_1654,N_1494,N_1568);
and U1655 (N_1655,N_1562,N_1455);
xnor U1656 (N_1656,N_1503,N_1415);
nor U1657 (N_1657,N_1549,N_1554);
and U1658 (N_1658,N_1565,N_1532);
nand U1659 (N_1659,N_1558,N_1483);
and U1660 (N_1660,N_1526,N_1437);
nor U1661 (N_1661,N_1464,N_1579);
xnor U1662 (N_1662,N_1433,N_1583);
and U1663 (N_1663,N_1429,N_1454);
and U1664 (N_1664,N_1548,N_1489);
nor U1665 (N_1665,N_1407,N_1530);
xor U1666 (N_1666,N_1553,N_1403);
xor U1667 (N_1667,N_1487,N_1405);
xor U1668 (N_1668,N_1479,N_1517);
and U1669 (N_1669,N_1418,N_1498);
or U1670 (N_1670,N_1401,N_1551);
nor U1671 (N_1671,N_1522,N_1512);
xnor U1672 (N_1672,N_1421,N_1423);
xor U1673 (N_1673,N_1598,N_1511);
nor U1674 (N_1674,N_1410,N_1480);
or U1675 (N_1675,N_1501,N_1507);
or U1676 (N_1676,N_1525,N_1459);
xor U1677 (N_1677,N_1402,N_1404);
nor U1678 (N_1678,N_1417,N_1467);
and U1679 (N_1679,N_1555,N_1451);
nand U1680 (N_1680,N_1527,N_1578);
and U1681 (N_1681,N_1465,N_1510);
and U1682 (N_1682,N_1582,N_1570);
xnor U1683 (N_1683,N_1442,N_1545);
nand U1684 (N_1684,N_1518,N_1539);
and U1685 (N_1685,N_1414,N_1452);
or U1686 (N_1686,N_1531,N_1586);
nor U1687 (N_1687,N_1588,N_1599);
or U1688 (N_1688,N_1450,N_1485);
nor U1689 (N_1689,N_1567,N_1520);
xor U1690 (N_1690,N_1591,N_1462);
nor U1691 (N_1691,N_1572,N_1597);
xnor U1692 (N_1692,N_1444,N_1560);
nand U1693 (N_1693,N_1439,N_1449);
nand U1694 (N_1694,N_1534,N_1587);
nor U1695 (N_1695,N_1550,N_1552);
nor U1696 (N_1696,N_1535,N_1486);
xor U1697 (N_1697,N_1448,N_1569);
nand U1698 (N_1698,N_1446,N_1543);
or U1699 (N_1699,N_1469,N_1430);
nand U1700 (N_1700,N_1497,N_1493);
xnor U1701 (N_1701,N_1448,N_1505);
and U1702 (N_1702,N_1429,N_1508);
and U1703 (N_1703,N_1548,N_1451);
and U1704 (N_1704,N_1450,N_1463);
or U1705 (N_1705,N_1529,N_1507);
or U1706 (N_1706,N_1583,N_1518);
nand U1707 (N_1707,N_1540,N_1551);
nor U1708 (N_1708,N_1545,N_1597);
nor U1709 (N_1709,N_1467,N_1520);
and U1710 (N_1710,N_1537,N_1566);
xor U1711 (N_1711,N_1463,N_1567);
and U1712 (N_1712,N_1556,N_1531);
xor U1713 (N_1713,N_1472,N_1530);
nor U1714 (N_1714,N_1444,N_1590);
nor U1715 (N_1715,N_1514,N_1554);
xor U1716 (N_1716,N_1451,N_1458);
and U1717 (N_1717,N_1558,N_1477);
or U1718 (N_1718,N_1527,N_1574);
or U1719 (N_1719,N_1411,N_1448);
xnor U1720 (N_1720,N_1515,N_1468);
and U1721 (N_1721,N_1404,N_1553);
nand U1722 (N_1722,N_1468,N_1583);
xor U1723 (N_1723,N_1444,N_1404);
nand U1724 (N_1724,N_1554,N_1486);
nor U1725 (N_1725,N_1592,N_1475);
xnor U1726 (N_1726,N_1567,N_1435);
and U1727 (N_1727,N_1478,N_1566);
and U1728 (N_1728,N_1497,N_1506);
or U1729 (N_1729,N_1551,N_1531);
xor U1730 (N_1730,N_1599,N_1552);
and U1731 (N_1731,N_1538,N_1474);
xor U1732 (N_1732,N_1592,N_1570);
or U1733 (N_1733,N_1535,N_1433);
and U1734 (N_1734,N_1405,N_1491);
and U1735 (N_1735,N_1552,N_1516);
nor U1736 (N_1736,N_1455,N_1502);
or U1737 (N_1737,N_1488,N_1557);
and U1738 (N_1738,N_1443,N_1434);
nor U1739 (N_1739,N_1518,N_1445);
or U1740 (N_1740,N_1436,N_1588);
and U1741 (N_1741,N_1540,N_1464);
nand U1742 (N_1742,N_1498,N_1593);
xor U1743 (N_1743,N_1478,N_1592);
nand U1744 (N_1744,N_1565,N_1595);
or U1745 (N_1745,N_1541,N_1568);
xnor U1746 (N_1746,N_1586,N_1482);
and U1747 (N_1747,N_1409,N_1580);
nor U1748 (N_1748,N_1551,N_1453);
xor U1749 (N_1749,N_1532,N_1494);
and U1750 (N_1750,N_1506,N_1598);
or U1751 (N_1751,N_1455,N_1532);
nor U1752 (N_1752,N_1548,N_1403);
or U1753 (N_1753,N_1438,N_1533);
xor U1754 (N_1754,N_1419,N_1504);
nand U1755 (N_1755,N_1555,N_1527);
nand U1756 (N_1756,N_1465,N_1546);
and U1757 (N_1757,N_1495,N_1559);
or U1758 (N_1758,N_1440,N_1478);
and U1759 (N_1759,N_1576,N_1487);
xnor U1760 (N_1760,N_1456,N_1492);
or U1761 (N_1761,N_1462,N_1513);
nor U1762 (N_1762,N_1573,N_1514);
xnor U1763 (N_1763,N_1566,N_1484);
nor U1764 (N_1764,N_1415,N_1418);
nor U1765 (N_1765,N_1546,N_1494);
xnor U1766 (N_1766,N_1469,N_1405);
nand U1767 (N_1767,N_1527,N_1425);
nand U1768 (N_1768,N_1531,N_1541);
nand U1769 (N_1769,N_1503,N_1465);
nor U1770 (N_1770,N_1462,N_1469);
nand U1771 (N_1771,N_1554,N_1533);
xor U1772 (N_1772,N_1591,N_1556);
xnor U1773 (N_1773,N_1497,N_1541);
or U1774 (N_1774,N_1559,N_1467);
or U1775 (N_1775,N_1441,N_1494);
nand U1776 (N_1776,N_1462,N_1514);
nor U1777 (N_1777,N_1565,N_1474);
or U1778 (N_1778,N_1530,N_1575);
nand U1779 (N_1779,N_1565,N_1404);
and U1780 (N_1780,N_1508,N_1537);
nor U1781 (N_1781,N_1441,N_1511);
nor U1782 (N_1782,N_1453,N_1553);
and U1783 (N_1783,N_1449,N_1442);
nand U1784 (N_1784,N_1537,N_1518);
nor U1785 (N_1785,N_1552,N_1593);
nand U1786 (N_1786,N_1590,N_1523);
or U1787 (N_1787,N_1512,N_1559);
nand U1788 (N_1788,N_1475,N_1439);
xnor U1789 (N_1789,N_1472,N_1525);
or U1790 (N_1790,N_1537,N_1492);
nand U1791 (N_1791,N_1549,N_1553);
and U1792 (N_1792,N_1551,N_1406);
and U1793 (N_1793,N_1404,N_1448);
nor U1794 (N_1794,N_1535,N_1436);
nand U1795 (N_1795,N_1463,N_1402);
nand U1796 (N_1796,N_1448,N_1421);
or U1797 (N_1797,N_1502,N_1595);
or U1798 (N_1798,N_1492,N_1522);
or U1799 (N_1799,N_1546,N_1503);
nand U1800 (N_1800,N_1670,N_1762);
xnor U1801 (N_1801,N_1633,N_1799);
nand U1802 (N_1802,N_1656,N_1749);
or U1803 (N_1803,N_1754,N_1730);
xnor U1804 (N_1804,N_1751,N_1657);
nor U1805 (N_1805,N_1667,N_1700);
or U1806 (N_1806,N_1697,N_1776);
nor U1807 (N_1807,N_1734,N_1778);
and U1808 (N_1808,N_1757,N_1611);
xnor U1809 (N_1809,N_1648,N_1647);
nand U1810 (N_1810,N_1626,N_1682);
nand U1811 (N_1811,N_1732,N_1796);
or U1812 (N_1812,N_1737,N_1678);
nand U1813 (N_1813,N_1606,N_1688);
and U1814 (N_1814,N_1654,N_1694);
nor U1815 (N_1815,N_1690,N_1660);
or U1816 (N_1816,N_1603,N_1781);
and U1817 (N_1817,N_1637,N_1679);
nor U1818 (N_1818,N_1729,N_1768);
or U1819 (N_1819,N_1634,N_1775);
nand U1820 (N_1820,N_1613,N_1790);
xnor U1821 (N_1821,N_1643,N_1738);
or U1822 (N_1822,N_1722,N_1696);
and U1823 (N_1823,N_1675,N_1793);
or U1824 (N_1824,N_1714,N_1771);
or U1825 (N_1825,N_1685,N_1630);
and U1826 (N_1826,N_1784,N_1689);
and U1827 (N_1827,N_1604,N_1713);
nor U1828 (N_1828,N_1641,N_1698);
and U1829 (N_1829,N_1745,N_1725);
nor U1830 (N_1830,N_1780,N_1774);
and U1831 (N_1831,N_1798,N_1644);
nand U1832 (N_1832,N_1652,N_1632);
nand U1833 (N_1833,N_1707,N_1674);
nor U1834 (N_1834,N_1773,N_1770);
or U1835 (N_1835,N_1686,N_1691);
nand U1836 (N_1836,N_1721,N_1761);
nor U1837 (N_1837,N_1727,N_1699);
nor U1838 (N_1838,N_1795,N_1638);
or U1839 (N_1839,N_1785,N_1742);
nor U1840 (N_1840,N_1653,N_1709);
and U1841 (N_1841,N_1607,N_1706);
and U1842 (N_1842,N_1642,N_1792);
and U1843 (N_1843,N_1731,N_1625);
nor U1844 (N_1844,N_1602,N_1759);
nor U1845 (N_1845,N_1623,N_1684);
and U1846 (N_1846,N_1600,N_1758);
or U1847 (N_1847,N_1646,N_1763);
xor U1848 (N_1848,N_1621,N_1708);
or U1849 (N_1849,N_1736,N_1635);
xnor U1850 (N_1850,N_1767,N_1787);
or U1851 (N_1851,N_1664,N_1692);
xnor U1852 (N_1852,N_1662,N_1609);
nor U1853 (N_1853,N_1733,N_1628);
nand U1854 (N_1854,N_1605,N_1739);
or U1855 (N_1855,N_1741,N_1726);
xnor U1856 (N_1856,N_1693,N_1743);
xor U1857 (N_1857,N_1677,N_1710);
nor U1858 (N_1858,N_1665,N_1619);
nand U1859 (N_1859,N_1723,N_1614);
nor U1860 (N_1860,N_1748,N_1612);
and U1861 (N_1861,N_1711,N_1719);
xor U1862 (N_1862,N_1636,N_1772);
nor U1863 (N_1863,N_1673,N_1764);
or U1864 (N_1864,N_1794,N_1712);
or U1865 (N_1865,N_1720,N_1655);
or U1866 (N_1866,N_1610,N_1788);
and U1867 (N_1867,N_1649,N_1695);
nand U1868 (N_1868,N_1620,N_1615);
or U1869 (N_1869,N_1631,N_1783);
nand U1870 (N_1870,N_1617,N_1661);
nor U1871 (N_1871,N_1629,N_1683);
or U1872 (N_1872,N_1608,N_1715);
or U1873 (N_1873,N_1658,N_1766);
or U1874 (N_1874,N_1671,N_1797);
nand U1875 (N_1875,N_1645,N_1760);
xor U1876 (N_1876,N_1716,N_1755);
xnor U1877 (N_1877,N_1701,N_1650);
nor U1878 (N_1878,N_1747,N_1791);
or U1879 (N_1879,N_1601,N_1668);
nand U1880 (N_1880,N_1718,N_1779);
xor U1881 (N_1881,N_1676,N_1681);
nand U1882 (N_1882,N_1666,N_1752);
and U1883 (N_1883,N_1672,N_1717);
or U1884 (N_1884,N_1624,N_1687);
nor U1885 (N_1885,N_1703,N_1616);
nor U1886 (N_1886,N_1744,N_1680);
xnor U1887 (N_1887,N_1782,N_1663);
nor U1888 (N_1888,N_1705,N_1753);
nand U1889 (N_1889,N_1728,N_1740);
nand U1890 (N_1890,N_1765,N_1659);
nor U1891 (N_1891,N_1746,N_1618);
nor U1892 (N_1892,N_1639,N_1622);
or U1893 (N_1893,N_1789,N_1769);
and U1894 (N_1894,N_1704,N_1640);
xor U1895 (N_1895,N_1756,N_1627);
nor U1896 (N_1896,N_1702,N_1724);
nor U1897 (N_1897,N_1750,N_1735);
or U1898 (N_1898,N_1786,N_1777);
xor U1899 (N_1899,N_1651,N_1669);
nor U1900 (N_1900,N_1744,N_1612);
or U1901 (N_1901,N_1733,N_1711);
and U1902 (N_1902,N_1782,N_1797);
nand U1903 (N_1903,N_1791,N_1787);
nor U1904 (N_1904,N_1794,N_1739);
nand U1905 (N_1905,N_1735,N_1765);
or U1906 (N_1906,N_1797,N_1683);
nor U1907 (N_1907,N_1746,N_1608);
nor U1908 (N_1908,N_1703,N_1740);
and U1909 (N_1909,N_1792,N_1650);
or U1910 (N_1910,N_1696,N_1613);
nand U1911 (N_1911,N_1676,N_1680);
and U1912 (N_1912,N_1712,N_1633);
nor U1913 (N_1913,N_1646,N_1781);
nand U1914 (N_1914,N_1619,N_1601);
nand U1915 (N_1915,N_1674,N_1746);
nand U1916 (N_1916,N_1673,N_1793);
nand U1917 (N_1917,N_1720,N_1679);
and U1918 (N_1918,N_1717,N_1652);
xnor U1919 (N_1919,N_1688,N_1610);
and U1920 (N_1920,N_1678,N_1791);
and U1921 (N_1921,N_1788,N_1757);
or U1922 (N_1922,N_1664,N_1739);
xnor U1923 (N_1923,N_1743,N_1779);
or U1924 (N_1924,N_1672,N_1654);
and U1925 (N_1925,N_1619,N_1789);
or U1926 (N_1926,N_1672,N_1788);
nor U1927 (N_1927,N_1640,N_1733);
nand U1928 (N_1928,N_1626,N_1625);
or U1929 (N_1929,N_1611,N_1608);
nor U1930 (N_1930,N_1695,N_1799);
xor U1931 (N_1931,N_1612,N_1662);
nand U1932 (N_1932,N_1769,N_1757);
and U1933 (N_1933,N_1682,N_1709);
nand U1934 (N_1934,N_1666,N_1603);
or U1935 (N_1935,N_1729,N_1620);
nor U1936 (N_1936,N_1606,N_1785);
xor U1937 (N_1937,N_1721,N_1769);
nor U1938 (N_1938,N_1715,N_1782);
nand U1939 (N_1939,N_1751,N_1760);
and U1940 (N_1940,N_1608,N_1733);
xor U1941 (N_1941,N_1757,N_1741);
xor U1942 (N_1942,N_1682,N_1672);
xnor U1943 (N_1943,N_1792,N_1726);
xnor U1944 (N_1944,N_1797,N_1743);
and U1945 (N_1945,N_1762,N_1744);
nor U1946 (N_1946,N_1677,N_1640);
and U1947 (N_1947,N_1607,N_1636);
xnor U1948 (N_1948,N_1690,N_1684);
or U1949 (N_1949,N_1750,N_1619);
and U1950 (N_1950,N_1621,N_1796);
or U1951 (N_1951,N_1792,N_1699);
or U1952 (N_1952,N_1633,N_1642);
xnor U1953 (N_1953,N_1669,N_1636);
nor U1954 (N_1954,N_1692,N_1673);
xor U1955 (N_1955,N_1642,N_1605);
nor U1956 (N_1956,N_1732,N_1645);
and U1957 (N_1957,N_1753,N_1624);
nor U1958 (N_1958,N_1633,N_1779);
nor U1959 (N_1959,N_1727,N_1730);
or U1960 (N_1960,N_1744,N_1778);
nor U1961 (N_1961,N_1700,N_1615);
or U1962 (N_1962,N_1705,N_1703);
or U1963 (N_1963,N_1672,N_1651);
nand U1964 (N_1964,N_1618,N_1716);
or U1965 (N_1965,N_1657,N_1766);
xnor U1966 (N_1966,N_1785,N_1692);
or U1967 (N_1967,N_1792,N_1772);
and U1968 (N_1968,N_1787,N_1674);
nor U1969 (N_1969,N_1628,N_1638);
and U1970 (N_1970,N_1698,N_1622);
nand U1971 (N_1971,N_1638,N_1671);
xor U1972 (N_1972,N_1785,N_1780);
xor U1973 (N_1973,N_1745,N_1605);
nor U1974 (N_1974,N_1715,N_1653);
or U1975 (N_1975,N_1697,N_1653);
nor U1976 (N_1976,N_1697,N_1758);
nand U1977 (N_1977,N_1746,N_1743);
nand U1978 (N_1978,N_1665,N_1734);
nor U1979 (N_1979,N_1600,N_1610);
nand U1980 (N_1980,N_1699,N_1653);
nor U1981 (N_1981,N_1783,N_1738);
nor U1982 (N_1982,N_1708,N_1651);
and U1983 (N_1983,N_1731,N_1705);
nor U1984 (N_1984,N_1767,N_1743);
nor U1985 (N_1985,N_1797,N_1756);
xnor U1986 (N_1986,N_1617,N_1695);
or U1987 (N_1987,N_1618,N_1632);
nand U1988 (N_1988,N_1794,N_1697);
nor U1989 (N_1989,N_1740,N_1794);
or U1990 (N_1990,N_1722,N_1644);
nor U1991 (N_1991,N_1639,N_1756);
and U1992 (N_1992,N_1684,N_1721);
nand U1993 (N_1993,N_1701,N_1642);
and U1994 (N_1994,N_1773,N_1782);
nor U1995 (N_1995,N_1747,N_1761);
and U1996 (N_1996,N_1746,N_1752);
xnor U1997 (N_1997,N_1604,N_1605);
xnor U1998 (N_1998,N_1793,N_1602);
nor U1999 (N_1999,N_1677,N_1713);
nand U2000 (N_2000,N_1895,N_1920);
or U2001 (N_2001,N_1987,N_1910);
xor U2002 (N_2002,N_1878,N_1867);
and U2003 (N_2003,N_1966,N_1834);
nor U2004 (N_2004,N_1958,N_1884);
nor U2005 (N_2005,N_1997,N_1840);
and U2006 (N_2006,N_1870,N_1925);
xnor U2007 (N_2007,N_1847,N_1805);
and U2008 (N_2008,N_1818,N_1892);
xnor U2009 (N_2009,N_1860,N_1983);
nor U2010 (N_2010,N_1957,N_1822);
nor U2011 (N_2011,N_1941,N_1896);
xor U2012 (N_2012,N_1981,N_1861);
and U2013 (N_2013,N_1857,N_1801);
and U2014 (N_2014,N_1943,N_1890);
nor U2015 (N_2015,N_1819,N_1820);
or U2016 (N_2016,N_1841,N_1998);
nand U2017 (N_2017,N_1931,N_1869);
and U2018 (N_2018,N_1855,N_1944);
nand U2019 (N_2019,N_1969,N_1811);
nor U2020 (N_2020,N_1833,N_1810);
nor U2021 (N_2021,N_1883,N_1832);
nand U2022 (N_2022,N_1826,N_1946);
and U2023 (N_2023,N_1924,N_1823);
xor U2024 (N_2024,N_1898,N_1971);
and U2025 (N_2025,N_1846,N_1942);
xnor U2026 (N_2026,N_1972,N_1836);
or U2027 (N_2027,N_1843,N_1901);
nor U2028 (N_2028,N_1885,N_1916);
nor U2029 (N_2029,N_1992,N_1927);
and U2030 (N_2030,N_1813,N_1935);
or U2031 (N_2031,N_1874,N_1933);
nand U2032 (N_2032,N_1871,N_1975);
nor U2033 (N_2033,N_1950,N_1868);
and U2034 (N_2034,N_1854,N_1959);
and U2035 (N_2035,N_1940,N_1937);
nor U2036 (N_2036,N_1915,N_1963);
xor U2037 (N_2037,N_1881,N_1835);
nor U2038 (N_2038,N_1995,N_1979);
nor U2039 (N_2039,N_1852,N_1825);
nor U2040 (N_2040,N_1990,N_1906);
xor U2041 (N_2041,N_1956,N_1803);
nor U2042 (N_2042,N_1917,N_1918);
nor U2043 (N_2043,N_1888,N_1951);
or U2044 (N_2044,N_1817,N_1945);
or U2045 (N_2045,N_1954,N_1856);
nor U2046 (N_2046,N_1902,N_1879);
and U2047 (N_2047,N_1932,N_1842);
xnor U2048 (N_2048,N_1815,N_1947);
or U2049 (N_2049,N_1982,N_1988);
xor U2050 (N_2050,N_1991,N_1904);
or U2051 (N_2051,N_1934,N_1827);
nand U2052 (N_2052,N_1919,N_1965);
or U2053 (N_2053,N_1865,N_1891);
nor U2054 (N_2054,N_1968,N_1866);
nand U2055 (N_2055,N_1912,N_1911);
xnor U2056 (N_2056,N_1922,N_1845);
and U2057 (N_2057,N_1844,N_1980);
or U2058 (N_2058,N_1887,N_1814);
xnor U2059 (N_2059,N_1936,N_1962);
and U2060 (N_2060,N_1996,N_1985);
and U2061 (N_2061,N_1889,N_1930);
xor U2062 (N_2062,N_1921,N_1804);
and U2063 (N_2063,N_1913,N_1830);
and U2064 (N_2064,N_1948,N_1923);
nand U2065 (N_2065,N_1955,N_1806);
nor U2066 (N_2066,N_1876,N_1964);
and U2067 (N_2067,N_1807,N_1899);
xor U2068 (N_2068,N_1863,N_1999);
xor U2069 (N_2069,N_1849,N_1821);
nor U2070 (N_2070,N_1812,N_1909);
nand U2071 (N_2071,N_1974,N_1929);
and U2072 (N_2072,N_1953,N_1926);
and U2073 (N_2073,N_1967,N_1952);
and U2074 (N_2074,N_1984,N_1838);
and U2075 (N_2075,N_1986,N_1993);
and U2076 (N_2076,N_1851,N_1976);
nand U2077 (N_2077,N_1872,N_1824);
nand U2078 (N_2078,N_1882,N_1831);
or U2079 (N_2079,N_1839,N_1864);
xor U2080 (N_2080,N_1949,N_1816);
or U2081 (N_2081,N_1928,N_1853);
and U2082 (N_2082,N_1873,N_1875);
and U2083 (N_2083,N_1905,N_1850);
or U2084 (N_2084,N_1828,N_1894);
or U2085 (N_2085,N_1938,N_1877);
or U2086 (N_2086,N_1994,N_1960);
xor U2087 (N_2087,N_1802,N_1907);
xnor U2088 (N_2088,N_1809,N_1908);
xor U2089 (N_2089,N_1903,N_1862);
xor U2090 (N_2090,N_1961,N_1848);
and U2091 (N_2091,N_1886,N_1939);
or U2092 (N_2092,N_1829,N_1897);
nand U2093 (N_2093,N_1808,N_1893);
xor U2094 (N_2094,N_1970,N_1800);
nor U2095 (N_2095,N_1978,N_1977);
nor U2096 (N_2096,N_1914,N_1837);
nand U2097 (N_2097,N_1973,N_1900);
or U2098 (N_2098,N_1858,N_1989);
or U2099 (N_2099,N_1859,N_1880);
or U2100 (N_2100,N_1862,N_1848);
nor U2101 (N_2101,N_1861,N_1850);
xnor U2102 (N_2102,N_1858,N_1874);
nand U2103 (N_2103,N_1841,N_1946);
xnor U2104 (N_2104,N_1917,N_1982);
or U2105 (N_2105,N_1931,N_1866);
and U2106 (N_2106,N_1886,N_1889);
or U2107 (N_2107,N_1834,N_1844);
or U2108 (N_2108,N_1807,N_1863);
nor U2109 (N_2109,N_1828,N_1984);
nor U2110 (N_2110,N_1959,N_1852);
nor U2111 (N_2111,N_1938,N_1817);
and U2112 (N_2112,N_1822,N_1947);
and U2113 (N_2113,N_1851,N_1906);
nand U2114 (N_2114,N_1972,N_1827);
nand U2115 (N_2115,N_1905,N_1887);
and U2116 (N_2116,N_1960,N_1894);
or U2117 (N_2117,N_1934,N_1824);
xnor U2118 (N_2118,N_1808,N_1895);
nand U2119 (N_2119,N_1974,N_1933);
and U2120 (N_2120,N_1924,N_1947);
and U2121 (N_2121,N_1948,N_1900);
nor U2122 (N_2122,N_1979,N_1878);
nor U2123 (N_2123,N_1951,N_1933);
or U2124 (N_2124,N_1831,N_1843);
xnor U2125 (N_2125,N_1935,N_1920);
and U2126 (N_2126,N_1832,N_1950);
nor U2127 (N_2127,N_1994,N_1881);
and U2128 (N_2128,N_1885,N_1874);
nor U2129 (N_2129,N_1893,N_1890);
xor U2130 (N_2130,N_1806,N_1873);
xor U2131 (N_2131,N_1931,N_1836);
nand U2132 (N_2132,N_1850,N_1896);
xnor U2133 (N_2133,N_1845,N_1809);
xor U2134 (N_2134,N_1921,N_1978);
nor U2135 (N_2135,N_1864,N_1962);
xnor U2136 (N_2136,N_1871,N_1939);
and U2137 (N_2137,N_1909,N_1992);
xnor U2138 (N_2138,N_1978,N_1909);
xnor U2139 (N_2139,N_1964,N_1983);
and U2140 (N_2140,N_1922,N_1909);
xor U2141 (N_2141,N_1815,N_1847);
and U2142 (N_2142,N_1855,N_1928);
and U2143 (N_2143,N_1804,N_1867);
or U2144 (N_2144,N_1861,N_1837);
xor U2145 (N_2145,N_1950,N_1992);
xor U2146 (N_2146,N_1902,N_1960);
nor U2147 (N_2147,N_1924,N_1993);
and U2148 (N_2148,N_1870,N_1859);
xnor U2149 (N_2149,N_1999,N_1932);
or U2150 (N_2150,N_1938,N_1852);
nor U2151 (N_2151,N_1844,N_1878);
nand U2152 (N_2152,N_1977,N_1833);
nand U2153 (N_2153,N_1867,N_1933);
and U2154 (N_2154,N_1947,N_1931);
nor U2155 (N_2155,N_1906,N_1893);
nor U2156 (N_2156,N_1822,N_1996);
nand U2157 (N_2157,N_1926,N_1969);
or U2158 (N_2158,N_1955,N_1895);
nor U2159 (N_2159,N_1970,N_1919);
xor U2160 (N_2160,N_1917,N_1974);
nand U2161 (N_2161,N_1949,N_1951);
or U2162 (N_2162,N_1996,N_1823);
xnor U2163 (N_2163,N_1848,N_1856);
nor U2164 (N_2164,N_1800,N_1969);
nand U2165 (N_2165,N_1858,N_1866);
xnor U2166 (N_2166,N_1986,N_1847);
xnor U2167 (N_2167,N_1959,N_1936);
or U2168 (N_2168,N_1955,N_1886);
nand U2169 (N_2169,N_1976,N_1901);
xor U2170 (N_2170,N_1935,N_1937);
or U2171 (N_2171,N_1848,N_1866);
or U2172 (N_2172,N_1910,N_1878);
and U2173 (N_2173,N_1916,N_1907);
xnor U2174 (N_2174,N_1825,N_1896);
nand U2175 (N_2175,N_1886,N_1883);
or U2176 (N_2176,N_1953,N_1921);
nor U2177 (N_2177,N_1911,N_1978);
nor U2178 (N_2178,N_1838,N_1862);
xor U2179 (N_2179,N_1942,N_1894);
xnor U2180 (N_2180,N_1858,N_1845);
and U2181 (N_2181,N_1975,N_1877);
or U2182 (N_2182,N_1838,N_1963);
and U2183 (N_2183,N_1884,N_1920);
or U2184 (N_2184,N_1879,N_1938);
nor U2185 (N_2185,N_1954,N_1864);
and U2186 (N_2186,N_1963,N_1836);
nor U2187 (N_2187,N_1852,N_1821);
or U2188 (N_2188,N_1954,N_1965);
nor U2189 (N_2189,N_1900,N_1942);
nand U2190 (N_2190,N_1914,N_1839);
or U2191 (N_2191,N_1984,N_1863);
or U2192 (N_2192,N_1898,N_1816);
and U2193 (N_2193,N_1802,N_1866);
or U2194 (N_2194,N_1808,N_1915);
xor U2195 (N_2195,N_1880,N_1931);
or U2196 (N_2196,N_1866,N_1880);
nor U2197 (N_2197,N_1950,N_1907);
and U2198 (N_2198,N_1959,N_1978);
nand U2199 (N_2199,N_1841,N_1986);
and U2200 (N_2200,N_2103,N_2178);
and U2201 (N_2201,N_2037,N_2141);
nor U2202 (N_2202,N_2190,N_2100);
xor U2203 (N_2203,N_2187,N_2070);
and U2204 (N_2204,N_2024,N_2195);
or U2205 (N_2205,N_2073,N_2129);
xor U2206 (N_2206,N_2017,N_2076);
or U2207 (N_2207,N_2055,N_2130);
xnor U2208 (N_2208,N_2028,N_2036);
nor U2209 (N_2209,N_2108,N_2163);
and U2210 (N_2210,N_2083,N_2012);
nand U2211 (N_2211,N_2113,N_2044);
or U2212 (N_2212,N_2180,N_2063);
or U2213 (N_2213,N_2046,N_2145);
xnor U2214 (N_2214,N_2112,N_2080);
nand U2215 (N_2215,N_2039,N_2020);
nor U2216 (N_2216,N_2124,N_2142);
and U2217 (N_2217,N_2048,N_2092);
or U2218 (N_2218,N_2116,N_2122);
and U2219 (N_2219,N_2121,N_2167);
and U2220 (N_2220,N_2001,N_2060);
xnor U2221 (N_2221,N_2188,N_2128);
nand U2222 (N_2222,N_2015,N_2027);
xor U2223 (N_2223,N_2157,N_2052);
nor U2224 (N_2224,N_2000,N_2010);
xnor U2225 (N_2225,N_2197,N_2158);
nand U2226 (N_2226,N_2084,N_2031);
nand U2227 (N_2227,N_2185,N_2127);
nand U2228 (N_2228,N_2061,N_2057);
nor U2229 (N_2229,N_2183,N_2101);
and U2230 (N_2230,N_2082,N_2176);
and U2231 (N_2231,N_2096,N_2053);
xnor U2232 (N_2232,N_2035,N_2032);
or U2233 (N_2233,N_2146,N_2072);
or U2234 (N_2234,N_2194,N_2054);
and U2235 (N_2235,N_2090,N_2033);
nor U2236 (N_2236,N_2134,N_2115);
and U2237 (N_2237,N_2182,N_2049);
or U2238 (N_2238,N_2192,N_2114);
nor U2239 (N_2239,N_2013,N_2022);
or U2240 (N_2240,N_2008,N_2136);
and U2241 (N_2241,N_2043,N_2105);
and U2242 (N_2242,N_2109,N_2120);
and U2243 (N_2243,N_2119,N_2034);
or U2244 (N_2244,N_2047,N_2099);
xnor U2245 (N_2245,N_2087,N_2071);
and U2246 (N_2246,N_2179,N_2021);
and U2247 (N_2247,N_2156,N_2093);
and U2248 (N_2248,N_2016,N_2118);
and U2249 (N_2249,N_2152,N_2111);
or U2250 (N_2250,N_2005,N_2170);
nand U2251 (N_2251,N_2155,N_2038);
nor U2252 (N_2252,N_2161,N_2160);
nor U2253 (N_2253,N_2079,N_2097);
and U2254 (N_2254,N_2040,N_2050);
nand U2255 (N_2255,N_2162,N_2198);
and U2256 (N_2256,N_2007,N_2173);
nor U2257 (N_2257,N_2058,N_2125);
xor U2258 (N_2258,N_2117,N_2159);
nand U2259 (N_2259,N_2110,N_2154);
nor U2260 (N_2260,N_2069,N_2014);
nor U2261 (N_2261,N_2098,N_2177);
nor U2262 (N_2262,N_2009,N_2102);
and U2263 (N_2263,N_2002,N_2067);
nor U2264 (N_2264,N_2151,N_2165);
nand U2265 (N_2265,N_2189,N_2042);
and U2266 (N_2266,N_2186,N_2088);
and U2267 (N_2267,N_2095,N_2003);
nand U2268 (N_2268,N_2107,N_2150);
nand U2269 (N_2269,N_2153,N_2074);
xnor U2270 (N_2270,N_2051,N_2123);
xnor U2271 (N_2271,N_2019,N_2004);
or U2272 (N_2272,N_2174,N_2068);
and U2273 (N_2273,N_2029,N_2089);
and U2274 (N_2274,N_2062,N_2196);
nor U2275 (N_2275,N_2065,N_2056);
nand U2276 (N_2276,N_2140,N_2137);
nor U2277 (N_2277,N_2106,N_2094);
or U2278 (N_2278,N_2149,N_2172);
nand U2279 (N_2279,N_2166,N_2059);
and U2280 (N_2280,N_2045,N_2143);
nor U2281 (N_2281,N_2184,N_2139);
nand U2282 (N_2282,N_2025,N_2011);
nand U2283 (N_2283,N_2018,N_2085);
nor U2284 (N_2284,N_2023,N_2026);
xor U2285 (N_2285,N_2144,N_2077);
xor U2286 (N_2286,N_2164,N_2133);
nand U2287 (N_2287,N_2006,N_2168);
xor U2288 (N_2288,N_2064,N_2199);
or U2289 (N_2289,N_2041,N_2091);
nor U2290 (N_2290,N_2131,N_2147);
or U2291 (N_2291,N_2175,N_2078);
nor U2292 (N_2292,N_2132,N_2138);
and U2293 (N_2293,N_2081,N_2104);
and U2294 (N_2294,N_2191,N_2169);
nor U2295 (N_2295,N_2148,N_2181);
xor U2296 (N_2296,N_2126,N_2075);
and U2297 (N_2297,N_2171,N_2193);
nor U2298 (N_2298,N_2086,N_2135);
or U2299 (N_2299,N_2066,N_2030);
xnor U2300 (N_2300,N_2176,N_2178);
nand U2301 (N_2301,N_2097,N_2082);
xnor U2302 (N_2302,N_2013,N_2071);
nor U2303 (N_2303,N_2096,N_2167);
xor U2304 (N_2304,N_2178,N_2177);
and U2305 (N_2305,N_2176,N_2195);
xnor U2306 (N_2306,N_2188,N_2106);
nand U2307 (N_2307,N_2037,N_2122);
or U2308 (N_2308,N_2063,N_2197);
or U2309 (N_2309,N_2033,N_2159);
xor U2310 (N_2310,N_2041,N_2028);
xor U2311 (N_2311,N_2090,N_2143);
or U2312 (N_2312,N_2012,N_2186);
and U2313 (N_2313,N_2112,N_2097);
nand U2314 (N_2314,N_2089,N_2093);
xnor U2315 (N_2315,N_2004,N_2066);
nand U2316 (N_2316,N_2007,N_2113);
xor U2317 (N_2317,N_2159,N_2068);
nor U2318 (N_2318,N_2011,N_2160);
nor U2319 (N_2319,N_2088,N_2050);
or U2320 (N_2320,N_2016,N_2139);
and U2321 (N_2321,N_2122,N_2097);
nor U2322 (N_2322,N_2007,N_2165);
xnor U2323 (N_2323,N_2060,N_2118);
and U2324 (N_2324,N_2119,N_2035);
nor U2325 (N_2325,N_2164,N_2127);
xnor U2326 (N_2326,N_2155,N_2030);
nand U2327 (N_2327,N_2171,N_2124);
xnor U2328 (N_2328,N_2137,N_2135);
nor U2329 (N_2329,N_2039,N_2048);
and U2330 (N_2330,N_2117,N_2025);
and U2331 (N_2331,N_2171,N_2001);
nor U2332 (N_2332,N_2058,N_2027);
or U2333 (N_2333,N_2090,N_2118);
and U2334 (N_2334,N_2148,N_2143);
or U2335 (N_2335,N_2004,N_2077);
xnor U2336 (N_2336,N_2106,N_2161);
nand U2337 (N_2337,N_2121,N_2120);
xnor U2338 (N_2338,N_2086,N_2185);
xor U2339 (N_2339,N_2125,N_2145);
and U2340 (N_2340,N_2172,N_2064);
and U2341 (N_2341,N_2033,N_2024);
nand U2342 (N_2342,N_2165,N_2096);
nand U2343 (N_2343,N_2059,N_2152);
and U2344 (N_2344,N_2115,N_2027);
nand U2345 (N_2345,N_2092,N_2178);
nor U2346 (N_2346,N_2185,N_2072);
and U2347 (N_2347,N_2114,N_2094);
nor U2348 (N_2348,N_2100,N_2152);
and U2349 (N_2349,N_2068,N_2045);
and U2350 (N_2350,N_2193,N_2099);
and U2351 (N_2351,N_2102,N_2047);
or U2352 (N_2352,N_2034,N_2172);
nand U2353 (N_2353,N_2081,N_2072);
and U2354 (N_2354,N_2189,N_2102);
or U2355 (N_2355,N_2152,N_2160);
nand U2356 (N_2356,N_2033,N_2073);
xnor U2357 (N_2357,N_2196,N_2139);
xnor U2358 (N_2358,N_2080,N_2082);
or U2359 (N_2359,N_2128,N_2006);
or U2360 (N_2360,N_2088,N_2164);
and U2361 (N_2361,N_2021,N_2117);
or U2362 (N_2362,N_2036,N_2120);
xnor U2363 (N_2363,N_2141,N_2159);
nand U2364 (N_2364,N_2096,N_2064);
and U2365 (N_2365,N_2052,N_2033);
xnor U2366 (N_2366,N_2018,N_2015);
nor U2367 (N_2367,N_2197,N_2127);
and U2368 (N_2368,N_2056,N_2123);
and U2369 (N_2369,N_2169,N_2134);
nand U2370 (N_2370,N_2102,N_2021);
xnor U2371 (N_2371,N_2079,N_2198);
or U2372 (N_2372,N_2018,N_2198);
nand U2373 (N_2373,N_2170,N_2188);
xnor U2374 (N_2374,N_2163,N_2140);
and U2375 (N_2375,N_2066,N_2145);
or U2376 (N_2376,N_2175,N_2110);
and U2377 (N_2377,N_2149,N_2168);
xor U2378 (N_2378,N_2018,N_2167);
or U2379 (N_2379,N_2046,N_2070);
or U2380 (N_2380,N_2190,N_2005);
xnor U2381 (N_2381,N_2091,N_2075);
nor U2382 (N_2382,N_2010,N_2113);
and U2383 (N_2383,N_2041,N_2093);
xor U2384 (N_2384,N_2034,N_2150);
nor U2385 (N_2385,N_2017,N_2121);
and U2386 (N_2386,N_2091,N_2085);
nor U2387 (N_2387,N_2025,N_2055);
nor U2388 (N_2388,N_2007,N_2049);
xor U2389 (N_2389,N_2192,N_2106);
nor U2390 (N_2390,N_2126,N_2130);
or U2391 (N_2391,N_2048,N_2131);
or U2392 (N_2392,N_2083,N_2091);
or U2393 (N_2393,N_2194,N_2035);
nor U2394 (N_2394,N_2174,N_2184);
and U2395 (N_2395,N_2062,N_2155);
nor U2396 (N_2396,N_2061,N_2012);
xnor U2397 (N_2397,N_2186,N_2128);
nor U2398 (N_2398,N_2010,N_2014);
nor U2399 (N_2399,N_2014,N_2007);
xnor U2400 (N_2400,N_2329,N_2359);
and U2401 (N_2401,N_2228,N_2285);
xor U2402 (N_2402,N_2335,N_2298);
or U2403 (N_2403,N_2311,N_2302);
xor U2404 (N_2404,N_2206,N_2254);
or U2405 (N_2405,N_2300,N_2290);
xor U2406 (N_2406,N_2327,N_2264);
xor U2407 (N_2407,N_2395,N_2317);
nand U2408 (N_2408,N_2343,N_2266);
xnor U2409 (N_2409,N_2344,N_2340);
nand U2410 (N_2410,N_2309,N_2246);
nor U2411 (N_2411,N_2288,N_2238);
xnor U2412 (N_2412,N_2313,N_2339);
nor U2413 (N_2413,N_2377,N_2357);
nand U2414 (N_2414,N_2349,N_2369);
and U2415 (N_2415,N_2213,N_2379);
nor U2416 (N_2416,N_2223,N_2208);
xnor U2417 (N_2417,N_2323,N_2227);
xnor U2418 (N_2418,N_2203,N_2338);
nand U2419 (N_2419,N_2386,N_2326);
xor U2420 (N_2420,N_2282,N_2381);
and U2421 (N_2421,N_2352,N_2333);
or U2422 (N_2422,N_2371,N_2296);
xnor U2423 (N_2423,N_2281,N_2256);
xor U2424 (N_2424,N_2234,N_2399);
and U2425 (N_2425,N_2244,N_2257);
or U2426 (N_2426,N_2398,N_2319);
xnor U2427 (N_2427,N_2305,N_2269);
and U2428 (N_2428,N_2366,N_2331);
or U2429 (N_2429,N_2372,N_2321);
and U2430 (N_2430,N_2217,N_2219);
nand U2431 (N_2431,N_2378,N_2316);
xnor U2432 (N_2432,N_2358,N_2389);
xnor U2433 (N_2433,N_2235,N_2236);
xnor U2434 (N_2434,N_2363,N_2255);
nor U2435 (N_2435,N_2258,N_2367);
xor U2436 (N_2436,N_2364,N_2240);
nor U2437 (N_2437,N_2283,N_2248);
or U2438 (N_2438,N_2259,N_2355);
nor U2439 (N_2439,N_2376,N_2224);
xnor U2440 (N_2440,N_2273,N_2230);
or U2441 (N_2441,N_2210,N_2265);
and U2442 (N_2442,N_2251,N_2370);
and U2443 (N_2443,N_2216,N_2347);
and U2444 (N_2444,N_2249,N_2293);
xor U2445 (N_2445,N_2297,N_2214);
and U2446 (N_2446,N_2330,N_2229);
nand U2447 (N_2447,N_2375,N_2205);
xor U2448 (N_2448,N_2306,N_2299);
and U2449 (N_2449,N_2303,N_2390);
and U2450 (N_2450,N_2263,N_2289);
xor U2451 (N_2451,N_2384,N_2294);
xnor U2452 (N_2452,N_2292,N_2360);
nor U2453 (N_2453,N_2241,N_2337);
xor U2454 (N_2454,N_2267,N_2304);
nand U2455 (N_2455,N_2325,N_2314);
or U2456 (N_2456,N_2276,N_2200);
xor U2457 (N_2457,N_2345,N_2272);
nor U2458 (N_2458,N_2368,N_2354);
xor U2459 (N_2459,N_2373,N_2271);
or U2460 (N_2460,N_2312,N_2211);
nand U2461 (N_2461,N_2374,N_2270);
and U2462 (N_2462,N_2348,N_2320);
nand U2463 (N_2463,N_2252,N_2231);
nand U2464 (N_2464,N_2392,N_2388);
nor U2465 (N_2465,N_2295,N_2286);
nor U2466 (N_2466,N_2237,N_2382);
nor U2467 (N_2467,N_2361,N_2260);
nand U2468 (N_2468,N_2350,N_2262);
nor U2469 (N_2469,N_2336,N_2346);
nor U2470 (N_2470,N_2274,N_2394);
or U2471 (N_2471,N_2342,N_2222);
nand U2472 (N_2472,N_2387,N_2221);
nand U2473 (N_2473,N_2332,N_2396);
and U2474 (N_2474,N_2383,N_2334);
or U2475 (N_2475,N_2207,N_2279);
or U2476 (N_2476,N_2324,N_2307);
nor U2477 (N_2477,N_2318,N_2287);
xnor U2478 (N_2478,N_2380,N_2362);
xor U2479 (N_2479,N_2397,N_2351);
xnor U2480 (N_2480,N_2385,N_2253);
nand U2481 (N_2481,N_2261,N_2328);
nand U2482 (N_2482,N_2353,N_2308);
nor U2483 (N_2483,N_2277,N_2365);
or U2484 (N_2484,N_2212,N_2393);
xor U2485 (N_2485,N_2209,N_2250);
or U2486 (N_2486,N_2275,N_2291);
xnor U2487 (N_2487,N_2310,N_2284);
xnor U2488 (N_2488,N_2243,N_2201);
nor U2489 (N_2489,N_2204,N_2341);
xnor U2490 (N_2490,N_2233,N_2226);
and U2491 (N_2491,N_2391,N_2245);
xor U2492 (N_2492,N_2322,N_2278);
or U2493 (N_2493,N_2239,N_2315);
nor U2494 (N_2494,N_2215,N_2280);
nand U2495 (N_2495,N_2220,N_2218);
nand U2496 (N_2496,N_2232,N_2356);
and U2497 (N_2497,N_2242,N_2301);
and U2498 (N_2498,N_2202,N_2268);
and U2499 (N_2499,N_2225,N_2247);
and U2500 (N_2500,N_2214,N_2317);
or U2501 (N_2501,N_2292,N_2227);
nor U2502 (N_2502,N_2335,N_2383);
nor U2503 (N_2503,N_2253,N_2316);
and U2504 (N_2504,N_2261,N_2218);
or U2505 (N_2505,N_2245,N_2223);
nor U2506 (N_2506,N_2206,N_2326);
and U2507 (N_2507,N_2388,N_2229);
nand U2508 (N_2508,N_2311,N_2371);
or U2509 (N_2509,N_2266,N_2369);
xor U2510 (N_2510,N_2211,N_2314);
or U2511 (N_2511,N_2363,N_2369);
nand U2512 (N_2512,N_2303,N_2233);
nor U2513 (N_2513,N_2221,N_2362);
nor U2514 (N_2514,N_2228,N_2308);
nor U2515 (N_2515,N_2217,N_2244);
and U2516 (N_2516,N_2351,N_2355);
nand U2517 (N_2517,N_2334,N_2397);
nand U2518 (N_2518,N_2237,N_2335);
or U2519 (N_2519,N_2253,N_2364);
or U2520 (N_2520,N_2210,N_2296);
nor U2521 (N_2521,N_2302,N_2207);
nand U2522 (N_2522,N_2266,N_2264);
nand U2523 (N_2523,N_2295,N_2363);
nand U2524 (N_2524,N_2394,N_2263);
nor U2525 (N_2525,N_2330,N_2392);
or U2526 (N_2526,N_2360,N_2270);
and U2527 (N_2527,N_2245,N_2232);
xor U2528 (N_2528,N_2324,N_2250);
and U2529 (N_2529,N_2252,N_2309);
xor U2530 (N_2530,N_2396,N_2223);
nor U2531 (N_2531,N_2389,N_2308);
nor U2532 (N_2532,N_2275,N_2300);
nand U2533 (N_2533,N_2311,N_2285);
or U2534 (N_2534,N_2279,N_2318);
nor U2535 (N_2535,N_2364,N_2264);
or U2536 (N_2536,N_2307,N_2304);
nor U2537 (N_2537,N_2200,N_2246);
or U2538 (N_2538,N_2210,N_2398);
nor U2539 (N_2539,N_2272,N_2276);
nor U2540 (N_2540,N_2374,N_2308);
and U2541 (N_2541,N_2231,N_2333);
nor U2542 (N_2542,N_2349,N_2384);
or U2543 (N_2543,N_2349,N_2360);
nor U2544 (N_2544,N_2292,N_2205);
or U2545 (N_2545,N_2243,N_2359);
and U2546 (N_2546,N_2393,N_2240);
or U2547 (N_2547,N_2307,N_2228);
xor U2548 (N_2548,N_2216,N_2326);
nor U2549 (N_2549,N_2385,N_2243);
xor U2550 (N_2550,N_2332,N_2351);
or U2551 (N_2551,N_2250,N_2354);
and U2552 (N_2552,N_2218,N_2272);
and U2553 (N_2553,N_2221,N_2333);
or U2554 (N_2554,N_2252,N_2202);
nor U2555 (N_2555,N_2268,N_2382);
or U2556 (N_2556,N_2335,N_2316);
and U2557 (N_2557,N_2230,N_2379);
nand U2558 (N_2558,N_2263,N_2257);
nand U2559 (N_2559,N_2337,N_2374);
and U2560 (N_2560,N_2200,N_2327);
or U2561 (N_2561,N_2267,N_2302);
nor U2562 (N_2562,N_2229,N_2285);
nand U2563 (N_2563,N_2256,N_2377);
nand U2564 (N_2564,N_2322,N_2208);
xor U2565 (N_2565,N_2239,N_2338);
nor U2566 (N_2566,N_2219,N_2312);
xor U2567 (N_2567,N_2386,N_2305);
nor U2568 (N_2568,N_2295,N_2355);
or U2569 (N_2569,N_2205,N_2289);
xor U2570 (N_2570,N_2349,N_2227);
or U2571 (N_2571,N_2237,N_2268);
nor U2572 (N_2572,N_2383,N_2319);
xor U2573 (N_2573,N_2274,N_2344);
nand U2574 (N_2574,N_2235,N_2395);
or U2575 (N_2575,N_2281,N_2366);
nor U2576 (N_2576,N_2312,N_2328);
xor U2577 (N_2577,N_2340,N_2229);
xor U2578 (N_2578,N_2333,N_2385);
nand U2579 (N_2579,N_2219,N_2216);
nor U2580 (N_2580,N_2264,N_2219);
and U2581 (N_2581,N_2246,N_2304);
nor U2582 (N_2582,N_2312,N_2380);
nor U2583 (N_2583,N_2242,N_2259);
xnor U2584 (N_2584,N_2347,N_2316);
or U2585 (N_2585,N_2295,N_2378);
xor U2586 (N_2586,N_2256,N_2202);
nor U2587 (N_2587,N_2396,N_2234);
xnor U2588 (N_2588,N_2336,N_2283);
nor U2589 (N_2589,N_2397,N_2341);
xnor U2590 (N_2590,N_2362,N_2260);
nor U2591 (N_2591,N_2385,N_2319);
and U2592 (N_2592,N_2396,N_2360);
or U2593 (N_2593,N_2251,N_2299);
nor U2594 (N_2594,N_2341,N_2378);
and U2595 (N_2595,N_2286,N_2213);
xor U2596 (N_2596,N_2281,N_2372);
and U2597 (N_2597,N_2226,N_2206);
and U2598 (N_2598,N_2303,N_2364);
or U2599 (N_2599,N_2373,N_2273);
or U2600 (N_2600,N_2459,N_2589);
xnor U2601 (N_2601,N_2576,N_2598);
xnor U2602 (N_2602,N_2444,N_2527);
and U2603 (N_2603,N_2582,N_2522);
and U2604 (N_2604,N_2478,N_2487);
xor U2605 (N_2605,N_2473,N_2420);
nand U2606 (N_2606,N_2418,N_2422);
nand U2607 (N_2607,N_2541,N_2448);
nor U2608 (N_2608,N_2513,N_2560);
nor U2609 (N_2609,N_2403,N_2536);
nand U2610 (N_2610,N_2509,N_2592);
or U2611 (N_2611,N_2421,N_2593);
nand U2612 (N_2612,N_2557,N_2491);
nor U2613 (N_2613,N_2575,N_2558);
and U2614 (N_2614,N_2590,N_2481);
nor U2615 (N_2615,N_2532,N_2409);
xor U2616 (N_2616,N_2432,N_2567);
and U2617 (N_2617,N_2597,N_2428);
and U2618 (N_2618,N_2440,N_2562);
or U2619 (N_2619,N_2534,N_2551);
or U2620 (N_2620,N_2416,N_2460);
nor U2621 (N_2621,N_2484,N_2568);
or U2622 (N_2622,N_2542,N_2407);
and U2623 (N_2623,N_2559,N_2445);
nor U2624 (N_2624,N_2578,N_2539);
and U2625 (N_2625,N_2454,N_2424);
nor U2626 (N_2626,N_2430,N_2492);
or U2627 (N_2627,N_2437,N_2436);
nor U2628 (N_2628,N_2468,N_2431);
xnor U2629 (N_2629,N_2419,N_2434);
nand U2630 (N_2630,N_2449,N_2503);
xnor U2631 (N_2631,N_2417,N_2521);
xor U2632 (N_2632,N_2573,N_2554);
or U2633 (N_2633,N_2599,N_2476);
nand U2634 (N_2634,N_2563,N_2496);
nand U2635 (N_2635,N_2435,N_2564);
nand U2636 (N_2636,N_2498,N_2486);
or U2637 (N_2637,N_2512,N_2585);
and U2638 (N_2638,N_2502,N_2415);
nor U2639 (N_2639,N_2517,N_2553);
nand U2640 (N_2640,N_2406,N_2427);
nand U2641 (N_2641,N_2547,N_2561);
nor U2642 (N_2642,N_2401,N_2402);
nand U2643 (N_2643,N_2556,N_2588);
nor U2644 (N_2644,N_2494,N_2495);
or U2645 (N_2645,N_2543,N_2530);
nand U2646 (N_2646,N_2471,N_2463);
and U2647 (N_2647,N_2456,N_2526);
or U2648 (N_2648,N_2482,N_2574);
nand U2649 (N_2649,N_2523,N_2462);
nand U2650 (N_2650,N_2480,N_2524);
nand U2651 (N_2651,N_2508,N_2501);
nor U2652 (N_2652,N_2587,N_2514);
and U2653 (N_2653,N_2469,N_2472);
or U2654 (N_2654,N_2533,N_2583);
nand U2655 (N_2655,N_2477,N_2555);
nand U2656 (N_2656,N_2595,N_2571);
nand U2657 (N_2657,N_2457,N_2441);
and U2658 (N_2658,N_2520,N_2450);
nor U2659 (N_2659,N_2438,N_2447);
nand U2660 (N_2660,N_2552,N_2475);
and U2661 (N_2661,N_2572,N_2461);
nor U2662 (N_2662,N_2452,N_2584);
nand U2663 (N_2663,N_2466,N_2414);
and U2664 (N_2664,N_2537,N_2548);
and U2665 (N_2665,N_2442,N_2464);
nor U2666 (N_2666,N_2412,N_2538);
nand U2667 (N_2667,N_2413,N_2483);
xnor U2668 (N_2668,N_2485,N_2439);
nor U2669 (N_2669,N_2535,N_2565);
or U2670 (N_2670,N_2493,N_2580);
nor U2671 (N_2671,N_2549,N_2425);
xnor U2672 (N_2672,N_2507,N_2566);
xor U2673 (N_2673,N_2410,N_2499);
and U2674 (N_2674,N_2506,N_2516);
xnor U2675 (N_2675,N_2504,N_2570);
or U2676 (N_2676,N_2451,N_2569);
nand U2677 (N_2677,N_2594,N_2591);
nor U2678 (N_2678,N_2531,N_2511);
and U2679 (N_2679,N_2465,N_2515);
and U2680 (N_2680,N_2545,N_2458);
and U2681 (N_2681,N_2586,N_2488);
nand U2682 (N_2682,N_2529,N_2546);
xor U2683 (N_2683,N_2581,N_2405);
nand U2684 (N_2684,N_2479,N_2497);
or U2685 (N_2685,N_2467,N_2423);
xor U2686 (N_2686,N_2455,N_2426);
nand U2687 (N_2687,N_2470,N_2404);
or U2688 (N_2688,N_2540,N_2528);
and U2689 (N_2689,N_2443,N_2518);
and U2690 (N_2690,N_2489,N_2596);
or U2691 (N_2691,N_2577,N_2411);
or U2692 (N_2692,N_2474,N_2453);
or U2693 (N_2693,N_2429,N_2446);
xnor U2694 (N_2694,N_2433,N_2579);
and U2695 (N_2695,N_2550,N_2544);
nand U2696 (N_2696,N_2519,N_2490);
and U2697 (N_2697,N_2510,N_2525);
or U2698 (N_2698,N_2505,N_2408);
xor U2699 (N_2699,N_2500,N_2400);
and U2700 (N_2700,N_2461,N_2518);
nand U2701 (N_2701,N_2571,N_2502);
and U2702 (N_2702,N_2564,N_2543);
xor U2703 (N_2703,N_2517,N_2480);
and U2704 (N_2704,N_2405,N_2534);
nand U2705 (N_2705,N_2507,N_2542);
and U2706 (N_2706,N_2458,N_2421);
and U2707 (N_2707,N_2483,N_2426);
nand U2708 (N_2708,N_2416,N_2523);
and U2709 (N_2709,N_2551,N_2468);
nand U2710 (N_2710,N_2524,N_2486);
nand U2711 (N_2711,N_2408,N_2562);
or U2712 (N_2712,N_2448,N_2469);
nand U2713 (N_2713,N_2591,N_2464);
and U2714 (N_2714,N_2587,N_2583);
or U2715 (N_2715,N_2485,N_2547);
or U2716 (N_2716,N_2563,N_2527);
nor U2717 (N_2717,N_2478,N_2524);
or U2718 (N_2718,N_2522,N_2481);
nor U2719 (N_2719,N_2452,N_2556);
and U2720 (N_2720,N_2560,N_2474);
and U2721 (N_2721,N_2512,N_2470);
xnor U2722 (N_2722,N_2430,N_2511);
nand U2723 (N_2723,N_2433,N_2494);
and U2724 (N_2724,N_2578,N_2517);
xor U2725 (N_2725,N_2489,N_2480);
nor U2726 (N_2726,N_2455,N_2439);
nor U2727 (N_2727,N_2467,N_2520);
xor U2728 (N_2728,N_2595,N_2433);
nand U2729 (N_2729,N_2483,N_2457);
xor U2730 (N_2730,N_2577,N_2429);
nor U2731 (N_2731,N_2518,N_2493);
nor U2732 (N_2732,N_2539,N_2434);
xor U2733 (N_2733,N_2553,N_2582);
or U2734 (N_2734,N_2549,N_2400);
nor U2735 (N_2735,N_2499,N_2432);
xnor U2736 (N_2736,N_2514,N_2529);
or U2737 (N_2737,N_2551,N_2490);
or U2738 (N_2738,N_2576,N_2438);
nor U2739 (N_2739,N_2563,N_2408);
and U2740 (N_2740,N_2453,N_2466);
nand U2741 (N_2741,N_2548,N_2518);
or U2742 (N_2742,N_2571,N_2532);
xnor U2743 (N_2743,N_2453,N_2582);
nand U2744 (N_2744,N_2581,N_2481);
or U2745 (N_2745,N_2529,N_2528);
nor U2746 (N_2746,N_2473,N_2520);
xnor U2747 (N_2747,N_2568,N_2518);
xor U2748 (N_2748,N_2439,N_2454);
xnor U2749 (N_2749,N_2442,N_2446);
nor U2750 (N_2750,N_2447,N_2501);
xnor U2751 (N_2751,N_2512,N_2488);
nor U2752 (N_2752,N_2419,N_2515);
or U2753 (N_2753,N_2477,N_2589);
xor U2754 (N_2754,N_2406,N_2423);
xor U2755 (N_2755,N_2437,N_2406);
nor U2756 (N_2756,N_2436,N_2507);
or U2757 (N_2757,N_2547,N_2522);
and U2758 (N_2758,N_2424,N_2517);
xnor U2759 (N_2759,N_2480,N_2587);
or U2760 (N_2760,N_2493,N_2401);
nor U2761 (N_2761,N_2580,N_2413);
nor U2762 (N_2762,N_2555,N_2585);
nor U2763 (N_2763,N_2588,N_2535);
xor U2764 (N_2764,N_2497,N_2585);
xnor U2765 (N_2765,N_2555,N_2560);
xnor U2766 (N_2766,N_2410,N_2509);
nor U2767 (N_2767,N_2405,N_2510);
and U2768 (N_2768,N_2544,N_2560);
nor U2769 (N_2769,N_2522,N_2465);
nor U2770 (N_2770,N_2584,N_2499);
nor U2771 (N_2771,N_2417,N_2574);
xor U2772 (N_2772,N_2443,N_2516);
and U2773 (N_2773,N_2473,N_2562);
and U2774 (N_2774,N_2513,N_2545);
or U2775 (N_2775,N_2493,N_2437);
xor U2776 (N_2776,N_2492,N_2549);
or U2777 (N_2777,N_2534,N_2545);
nor U2778 (N_2778,N_2527,N_2418);
xnor U2779 (N_2779,N_2515,N_2508);
xnor U2780 (N_2780,N_2572,N_2466);
nand U2781 (N_2781,N_2457,N_2491);
nor U2782 (N_2782,N_2503,N_2578);
nand U2783 (N_2783,N_2548,N_2527);
xor U2784 (N_2784,N_2413,N_2407);
and U2785 (N_2785,N_2514,N_2580);
nand U2786 (N_2786,N_2404,N_2552);
nor U2787 (N_2787,N_2488,N_2528);
nand U2788 (N_2788,N_2565,N_2444);
xnor U2789 (N_2789,N_2582,N_2485);
xnor U2790 (N_2790,N_2475,N_2567);
and U2791 (N_2791,N_2585,N_2535);
and U2792 (N_2792,N_2512,N_2517);
or U2793 (N_2793,N_2557,N_2462);
and U2794 (N_2794,N_2416,N_2568);
xnor U2795 (N_2795,N_2575,N_2471);
nor U2796 (N_2796,N_2524,N_2488);
nor U2797 (N_2797,N_2465,N_2534);
nor U2798 (N_2798,N_2503,N_2550);
or U2799 (N_2799,N_2593,N_2543);
and U2800 (N_2800,N_2710,N_2786);
nand U2801 (N_2801,N_2658,N_2797);
or U2802 (N_2802,N_2762,N_2611);
and U2803 (N_2803,N_2662,N_2779);
nor U2804 (N_2804,N_2705,N_2600);
or U2805 (N_2805,N_2717,N_2711);
nor U2806 (N_2806,N_2706,N_2722);
and U2807 (N_2807,N_2769,N_2736);
or U2808 (N_2808,N_2663,N_2672);
nand U2809 (N_2809,N_2606,N_2643);
or U2810 (N_2810,N_2798,N_2699);
nand U2811 (N_2811,N_2759,N_2737);
nand U2812 (N_2812,N_2753,N_2703);
or U2813 (N_2813,N_2624,N_2751);
nor U2814 (N_2814,N_2620,N_2681);
nor U2815 (N_2815,N_2721,N_2634);
and U2816 (N_2816,N_2603,N_2716);
and U2817 (N_2817,N_2761,N_2612);
xor U2818 (N_2818,N_2622,N_2765);
nor U2819 (N_2819,N_2757,N_2678);
or U2820 (N_2820,N_2649,N_2646);
and U2821 (N_2821,N_2780,N_2684);
nand U2822 (N_2822,N_2726,N_2775);
xnor U2823 (N_2823,N_2701,N_2636);
xor U2824 (N_2824,N_2641,N_2788);
and U2825 (N_2825,N_2601,N_2627);
or U2826 (N_2826,N_2604,N_2756);
or U2827 (N_2827,N_2685,N_2629);
nor U2828 (N_2828,N_2741,N_2704);
and U2829 (N_2829,N_2693,N_2745);
nand U2830 (N_2830,N_2659,N_2764);
nor U2831 (N_2831,N_2760,N_2795);
nor U2832 (N_2832,N_2771,N_2785);
and U2833 (N_2833,N_2794,N_2719);
xnor U2834 (N_2834,N_2671,N_2748);
nand U2835 (N_2835,N_2694,N_2617);
or U2836 (N_2836,N_2645,N_2731);
nor U2837 (N_2837,N_2639,N_2682);
or U2838 (N_2838,N_2778,N_2730);
xnor U2839 (N_2839,N_2725,N_2792);
nand U2840 (N_2840,N_2735,N_2625);
nor U2841 (N_2841,N_2758,N_2616);
nor U2842 (N_2842,N_2680,N_2770);
nand U2843 (N_2843,N_2708,N_2790);
nor U2844 (N_2844,N_2637,N_2697);
nand U2845 (N_2845,N_2698,N_2644);
and U2846 (N_2846,N_2688,N_2689);
nand U2847 (N_2847,N_2667,N_2690);
and U2848 (N_2848,N_2669,N_2679);
xor U2849 (N_2849,N_2674,N_2618);
nor U2850 (N_2850,N_2783,N_2702);
and U2851 (N_2851,N_2747,N_2640);
nand U2852 (N_2852,N_2740,N_2712);
nand U2853 (N_2853,N_2615,N_2766);
nand U2854 (N_2854,N_2675,N_2631);
xor U2855 (N_2855,N_2687,N_2664);
nor U2856 (N_2856,N_2650,N_2743);
xnor U2857 (N_2857,N_2661,N_2666);
nor U2858 (N_2858,N_2668,N_2665);
or U2859 (N_2859,N_2720,N_2655);
xnor U2860 (N_2860,N_2619,N_2714);
nor U2861 (N_2861,N_2739,N_2749);
nand U2862 (N_2862,N_2709,N_2642);
or U2863 (N_2863,N_2784,N_2754);
nand U2864 (N_2864,N_2791,N_2746);
and U2865 (N_2865,N_2713,N_2676);
nor U2866 (N_2866,N_2610,N_2653);
or U2867 (N_2867,N_2626,N_2718);
nor U2868 (N_2868,N_2605,N_2633);
nand U2869 (N_2869,N_2776,N_2614);
nor U2870 (N_2870,N_2733,N_2632);
xnor U2871 (N_2871,N_2724,N_2648);
and U2872 (N_2872,N_2767,N_2742);
and U2873 (N_2873,N_2652,N_2781);
nor U2874 (N_2874,N_2602,N_2755);
xor U2875 (N_2875,N_2692,N_2707);
nand U2876 (N_2876,N_2777,N_2677);
nand U2877 (N_2877,N_2656,N_2750);
or U2878 (N_2878,N_2799,N_2729);
and U2879 (N_2879,N_2696,N_2628);
xnor U2880 (N_2880,N_2728,N_2793);
xor U2881 (N_2881,N_2651,N_2787);
xnor U2882 (N_2882,N_2673,N_2623);
and U2883 (N_2883,N_2621,N_2638);
nor U2884 (N_2884,N_2683,N_2715);
xor U2885 (N_2885,N_2608,N_2744);
or U2886 (N_2886,N_2654,N_2772);
nand U2887 (N_2887,N_2763,N_2773);
and U2888 (N_2888,N_2700,N_2782);
xor U2889 (N_2889,N_2630,N_2695);
xnor U2890 (N_2890,N_2660,N_2732);
xor U2891 (N_2891,N_2657,N_2686);
xnor U2892 (N_2892,N_2613,N_2647);
nand U2893 (N_2893,N_2670,N_2789);
nand U2894 (N_2894,N_2727,N_2774);
nand U2895 (N_2895,N_2609,N_2768);
xor U2896 (N_2896,N_2752,N_2635);
nand U2897 (N_2897,N_2607,N_2796);
or U2898 (N_2898,N_2738,N_2691);
nand U2899 (N_2899,N_2723,N_2734);
nand U2900 (N_2900,N_2715,N_2786);
and U2901 (N_2901,N_2730,N_2691);
or U2902 (N_2902,N_2731,N_2792);
nor U2903 (N_2903,N_2773,N_2753);
xor U2904 (N_2904,N_2677,N_2642);
xor U2905 (N_2905,N_2612,N_2753);
or U2906 (N_2906,N_2649,N_2698);
and U2907 (N_2907,N_2697,N_2711);
and U2908 (N_2908,N_2744,N_2698);
or U2909 (N_2909,N_2647,N_2753);
nand U2910 (N_2910,N_2628,N_2635);
nand U2911 (N_2911,N_2656,N_2730);
and U2912 (N_2912,N_2616,N_2645);
nand U2913 (N_2913,N_2642,N_2730);
and U2914 (N_2914,N_2780,N_2686);
xnor U2915 (N_2915,N_2630,N_2706);
or U2916 (N_2916,N_2798,N_2716);
nand U2917 (N_2917,N_2716,N_2773);
and U2918 (N_2918,N_2637,N_2734);
nor U2919 (N_2919,N_2663,N_2719);
or U2920 (N_2920,N_2687,N_2688);
or U2921 (N_2921,N_2733,N_2683);
or U2922 (N_2922,N_2731,N_2690);
nor U2923 (N_2923,N_2703,N_2735);
or U2924 (N_2924,N_2643,N_2798);
xor U2925 (N_2925,N_2619,N_2609);
xor U2926 (N_2926,N_2663,N_2660);
and U2927 (N_2927,N_2758,N_2768);
nor U2928 (N_2928,N_2748,N_2682);
or U2929 (N_2929,N_2600,N_2662);
nand U2930 (N_2930,N_2725,N_2784);
nor U2931 (N_2931,N_2626,N_2774);
xor U2932 (N_2932,N_2608,N_2616);
and U2933 (N_2933,N_2796,N_2626);
nor U2934 (N_2934,N_2712,N_2774);
and U2935 (N_2935,N_2643,N_2646);
xor U2936 (N_2936,N_2786,N_2649);
or U2937 (N_2937,N_2698,N_2625);
xnor U2938 (N_2938,N_2622,N_2740);
or U2939 (N_2939,N_2784,N_2605);
and U2940 (N_2940,N_2671,N_2616);
nor U2941 (N_2941,N_2746,N_2726);
or U2942 (N_2942,N_2665,N_2625);
nand U2943 (N_2943,N_2708,N_2717);
and U2944 (N_2944,N_2665,N_2673);
nand U2945 (N_2945,N_2731,N_2683);
xor U2946 (N_2946,N_2744,N_2746);
or U2947 (N_2947,N_2620,N_2695);
nand U2948 (N_2948,N_2790,N_2610);
nor U2949 (N_2949,N_2679,N_2721);
nand U2950 (N_2950,N_2659,N_2669);
nor U2951 (N_2951,N_2723,N_2649);
nand U2952 (N_2952,N_2654,N_2637);
nor U2953 (N_2953,N_2636,N_2643);
xor U2954 (N_2954,N_2753,N_2618);
and U2955 (N_2955,N_2738,N_2698);
nand U2956 (N_2956,N_2692,N_2791);
xor U2957 (N_2957,N_2756,N_2770);
or U2958 (N_2958,N_2754,N_2767);
nor U2959 (N_2959,N_2646,N_2779);
and U2960 (N_2960,N_2651,N_2788);
nor U2961 (N_2961,N_2733,N_2713);
and U2962 (N_2962,N_2648,N_2749);
xnor U2963 (N_2963,N_2697,N_2689);
xnor U2964 (N_2964,N_2655,N_2617);
nand U2965 (N_2965,N_2660,N_2657);
xnor U2966 (N_2966,N_2656,N_2641);
nor U2967 (N_2967,N_2620,N_2646);
nand U2968 (N_2968,N_2642,N_2656);
nand U2969 (N_2969,N_2714,N_2631);
and U2970 (N_2970,N_2768,N_2736);
or U2971 (N_2971,N_2726,N_2732);
and U2972 (N_2972,N_2600,N_2735);
nor U2973 (N_2973,N_2784,N_2790);
nand U2974 (N_2974,N_2681,N_2748);
xnor U2975 (N_2975,N_2643,N_2609);
nand U2976 (N_2976,N_2684,N_2610);
or U2977 (N_2977,N_2615,N_2642);
nor U2978 (N_2978,N_2758,N_2729);
xnor U2979 (N_2979,N_2630,N_2656);
or U2980 (N_2980,N_2704,N_2744);
nor U2981 (N_2981,N_2623,N_2644);
nor U2982 (N_2982,N_2786,N_2609);
nor U2983 (N_2983,N_2706,N_2719);
and U2984 (N_2984,N_2703,N_2707);
and U2985 (N_2985,N_2648,N_2766);
nand U2986 (N_2986,N_2788,N_2708);
or U2987 (N_2987,N_2766,N_2666);
xnor U2988 (N_2988,N_2631,N_2734);
nand U2989 (N_2989,N_2713,N_2603);
or U2990 (N_2990,N_2764,N_2773);
nand U2991 (N_2991,N_2755,N_2653);
or U2992 (N_2992,N_2668,N_2776);
nand U2993 (N_2993,N_2651,N_2724);
and U2994 (N_2994,N_2615,N_2731);
xor U2995 (N_2995,N_2757,N_2600);
nor U2996 (N_2996,N_2681,N_2685);
nand U2997 (N_2997,N_2664,N_2705);
xnor U2998 (N_2998,N_2661,N_2681);
nor U2999 (N_2999,N_2747,N_2731);
or UO_0 (O_0,N_2804,N_2845);
nand UO_1 (O_1,N_2934,N_2929);
nor UO_2 (O_2,N_2881,N_2919);
xor UO_3 (O_3,N_2990,N_2909);
nor UO_4 (O_4,N_2991,N_2925);
nor UO_5 (O_5,N_2817,N_2844);
nand UO_6 (O_6,N_2879,N_2923);
xnor UO_7 (O_7,N_2894,N_2943);
and UO_8 (O_8,N_2808,N_2836);
nor UO_9 (O_9,N_2969,N_2848);
xor UO_10 (O_10,N_2813,N_2889);
or UO_11 (O_11,N_2863,N_2945);
and UO_12 (O_12,N_2865,N_2853);
or UO_13 (O_13,N_2822,N_2801);
xor UO_14 (O_14,N_2873,N_2963);
and UO_15 (O_15,N_2912,N_2847);
nor UO_16 (O_16,N_2818,N_2953);
and UO_17 (O_17,N_2901,N_2922);
or UO_18 (O_18,N_2955,N_2852);
xnor UO_19 (O_19,N_2843,N_2829);
or UO_20 (O_20,N_2918,N_2993);
and UO_21 (O_21,N_2928,N_2957);
xor UO_22 (O_22,N_2867,N_2823);
or UO_23 (O_23,N_2954,N_2968);
nand UO_24 (O_24,N_2959,N_2996);
nand UO_25 (O_25,N_2905,N_2860);
or UO_26 (O_26,N_2897,N_2841);
nand UO_27 (O_27,N_2935,N_2807);
and UO_28 (O_28,N_2936,N_2902);
or UO_29 (O_29,N_2977,N_2885);
and UO_30 (O_30,N_2971,N_2927);
and UO_31 (O_31,N_2978,N_2988);
and UO_32 (O_32,N_2903,N_2877);
nor UO_33 (O_33,N_2962,N_2989);
nand UO_34 (O_34,N_2946,N_2854);
or UO_35 (O_35,N_2944,N_2839);
nand UO_36 (O_36,N_2824,N_2916);
or UO_37 (O_37,N_2811,N_2868);
nand UO_38 (O_38,N_2982,N_2961);
and UO_39 (O_39,N_2900,N_2999);
nor UO_40 (O_40,N_2932,N_2915);
nor UO_41 (O_41,N_2948,N_2883);
nand UO_42 (O_42,N_2896,N_2998);
nor UO_43 (O_43,N_2866,N_2908);
or UO_44 (O_44,N_2964,N_2842);
nand UO_45 (O_45,N_2907,N_2898);
or UO_46 (O_46,N_2956,N_2850);
nor UO_47 (O_47,N_2805,N_2886);
nand UO_48 (O_48,N_2814,N_2892);
nor UO_49 (O_49,N_2802,N_2921);
nor UO_50 (O_50,N_2933,N_2904);
nand UO_51 (O_51,N_2890,N_2970);
or UO_52 (O_52,N_2806,N_2880);
nor UO_53 (O_53,N_2859,N_2983);
nand UO_54 (O_54,N_2941,N_2851);
xor UO_55 (O_55,N_2887,N_2830);
xnor UO_56 (O_56,N_2986,N_2816);
and UO_57 (O_57,N_2975,N_2882);
or UO_58 (O_58,N_2980,N_2888);
nand UO_59 (O_59,N_2893,N_2924);
and UO_60 (O_60,N_2979,N_2895);
nand UO_61 (O_61,N_2828,N_2874);
nor UO_62 (O_62,N_2938,N_2913);
nor UO_63 (O_63,N_2967,N_2840);
and UO_64 (O_64,N_2878,N_2884);
or UO_65 (O_65,N_2870,N_2891);
or UO_66 (O_66,N_2871,N_2920);
xnor UO_67 (O_67,N_2984,N_2862);
or UO_68 (O_68,N_2931,N_2981);
nor UO_69 (O_69,N_2826,N_2858);
nor UO_70 (O_70,N_2869,N_2972);
or UO_71 (O_71,N_2820,N_2875);
nor UO_72 (O_72,N_2951,N_2833);
and UO_73 (O_73,N_2855,N_2876);
nor UO_74 (O_74,N_2809,N_2911);
and UO_75 (O_75,N_2952,N_2947);
xnor UO_76 (O_76,N_2906,N_2917);
and UO_77 (O_77,N_2857,N_2974);
and UO_78 (O_78,N_2930,N_2835);
or UO_79 (O_79,N_2815,N_2899);
and UO_80 (O_80,N_2825,N_2939);
and UO_81 (O_81,N_2965,N_2821);
xnor UO_82 (O_82,N_2810,N_2914);
and UO_83 (O_83,N_2864,N_2966);
xnor UO_84 (O_84,N_2846,N_2995);
or UO_85 (O_85,N_2827,N_2800);
or UO_86 (O_86,N_2832,N_2910);
xnor UO_87 (O_87,N_2994,N_2992);
nand UO_88 (O_88,N_2849,N_2973);
and UO_89 (O_89,N_2872,N_2942);
nor UO_90 (O_90,N_2838,N_2819);
xor UO_91 (O_91,N_2950,N_2803);
and UO_92 (O_92,N_2926,N_2861);
or UO_93 (O_93,N_2856,N_2985);
nor UO_94 (O_94,N_2960,N_2837);
and UO_95 (O_95,N_2958,N_2949);
nand UO_96 (O_96,N_2937,N_2834);
nand UO_97 (O_97,N_2940,N_2831);
nor UO_98 (O_98,N_2997,N_2812);
or UO_99 (O_99,N_2976,N_2987);
xor UO_100 (O_100,N_2974,N_2837);
xor UO_101 (O_101,N_2907,N_2874);
or UO_102 (O_102,N_2842,N_2931);
and UO_103 (O_103,N_2854,N_2851);
nand UO_104 (O_104,N_2879,N_2837);
or UO_105 (O_105,N_2840,N_2944);
or UO_106 (O_106,N_2831,N_2856);
nor UO_107 (O_107,N_2833,N_2814);
or UO_108 (O_108,N_2956,N_2962);
and UO_109 (O_109,N_2912,N_2836);
nand UO_110 (O_110,N_2805,N_2889);
xor UO_111 (O_111,N_2856,N_2879);
nand UO_112 (O_112,N_2827,N_2912);
nand UO_113 (O_113,N_2986,N_2966);
and UO_114 (O_114,N_2810,N_2844);
xnor UO_115 (O_115,N_2915,N_2861);
nor UO_116 (O_116,N_2866,N_2869);
or UO_117 (O_117,N_2928,N_2892);
nand UO_118 (O_118,N_2865,N_2877);
nand UO_119 (O_119,N_2888,N_2819);
xor UO_120 (O_120,N_2923,N_2939);
nor UO_121 (O_121,N_2810,N_2890);
nor UO_122 (O_122,N_2893,N_2871);
or UO_123 (O_123,N_2853,N_2894);
and UO_124 (O_124,N_2848,N_2938);
and UO_125 (O_125,N_2851,N_2965);
nand UO_126 (O_126,N_2879,N_2999);
and UO_127 (O_127,N_2855,N_2819);
xnor UO_128 (O_128,N_2958,N_2847);
xnor UO_129 (O_129,N_2858,N_2930);
nand UO_130 (O_130,N_2857,N_2830);
or UO_131 (O_131,N_2963,N_2800);
nor UO_132 (O_132,N_2837,N_2949);
nor UO_133 (O_133,N_2930,N_2808);
or UO_134 (O_134,N_2912,N_2877);
or UO_135 (O_135,N_2902,N_2823);
nand UO_136 (O_136,N_2946,N_2816);
nor UO_137 (O_137,N_2974,N_2815);
and UO_138 (O_138,N_2974,N_2934);
nor UO_139 (O_139,N_2864,N_2851);
xor UO_140 (O_140,N_2941,N_2933);
or UO_141 (O_141,N_2856,N_2853);
nor UO_142 (O_142,N_2888,N_2912);
xor UO_143 (O_143,N_2852,N_2811);
or UO_144 (O_144,N_2946,N_2867);
nand UO_145 (O_145,N_2860,N_2865);
and UO_146 (O_146,N_2986,N_2909);
and UO_147 (O_147,N_2892,N_2842);
nor UO_148 (O_148,N_2918,N_2803);
nor UO_149 (O_149,N_2920,N_2911);
and UO_150 (O_150,N_2840,N_2931);
nand UO_151 (O_151,N_2933,N_2883);
and UO_152 (O_152,N_2951,N_2991);
xor UO_153 (O_153,N_2886,N_2918);
and UO_154 (O_154,N_2844,N_2962);
nor UO_155 (O_155,N_2910,N_2964);
xor UO_156 (O_156,N_2827,N_2947);
or UO_157 (O_157,N_2876,N_2915);
xor UO_158 (O_158,N_2911,N_2923);
or UO_159 (O_159,N_2908,N_2875);
and UO_160 (O_160,N_2810,N_2858);
and UO_161 (O_161,N_2908,N_2960);
nand UO_162 (O_162,N_2877,N_2878);
xor UO_163 (O_163,N_2809,N_2862);
nand UO_164 (O_164,N_2815,N_2800);
xor UO_165 (O_165,N_2979,N_2980);
nand UO_166 (O_166,N_2953,N_2886);
or UO_167 (O_167,N_2964,N_2947);
or UO_168 (O_168,N_2937,N_2830);
nor UO_169 (O_169,N_2888,N_2941);
nor UO_170 (O_170,N_2855,N_2890);
nor UO_171 (O_171,N_2904,N_2934);
xor UO_172 (O_172,N_2878,N_2851);
and UO_173 (O_173,N_2979,N_2814);
and UO_174 (O_174,N_2823,N_2817);
nor UO_175 (O_175,N_2961,N_2905);
xor UO_176 (O_176,N_2874,N_2806);
xor UO_177 (O_177,N_2940,N_2873);
nand UO_178 (O_178,N_2963,N_2824);
nand UO_179 (O_179,N_2972,N_2958);
and UO_180 (O_180,N_2937,N_2954);
nor UO_181 (O_181,N_2909,N_2970);
or UO_182 (O_182,N_2843,N_2817);
and UO_183 (O_183,N_2805,N_2902);
nor UO_184 (O_184,N_2834,N_2816);
and UO_185 (O_185,N_2844,N_2827);
xnor UO_186 (O_186,N_2905,N_2846);
and UO_187 (O_187,N_2819,N_2928);
xnor UO_188 (O_188,N_2817,N_2869);
or UO_189 (O_189,N_2966,N_2962);
nor UO_190 (O_190,N_2832,N_2970);
nand UO_191 (O_191,N_2840,N_2911);
nand UO_192 (O_192,N_2874,N_2929);
and UO_193 (O_193,N_2917,N_2822);
nand UO_194 (O_194,N_2800,N_2818);
xor UO_195 (O_195,N_2930,N_2981);
or UO_196 (O_196,N_2999,N_2942);
nand UO_197 (O_197,N_2922,N_2999);
and UO_198 (O_198,N_2914,N_2911);
nor UO_199 (O_199,N_2875,N_2818);
xnor UO_200 (O_200,N_2943,N_2873);
and UO_201 (O_201,N_2900,N_2877);
and UO_202 (O_202,N_2974,N_2922);
nor UO_203 (O_203,N_2992,N_2884);
or UO_204 (O_204,N_2955,N_2927);
or UO_205 (O_205,N_2934,N_2931);
xor UO_206 (O_206,N_2841,N_2936);
xor UO_207 (O_207,N_2984,N_2918);
or UO_208 (O_208,N_2846,N_2850);
nand UO_209 (O_209,N_2969,N_2968);
or UO_210 (O_210,N_2849,N_2984);
nand UO_211 (O_211,N_2883,N_2895);
or UO_212 (O_212,N_2877,N_2902);
and UO_213 (O_213,N_2810,N_2881);
or UO_214 (O_214,N_2989,N_2908);
nand UO_215 (O_215,N_2996,N_2904);
and UO_216 (O_216,N_2936,N_2900);
and UO_217 (O_217,N_2867,N_2884);
xor UO_218 (O_218,N_2985,N_2989);
and UO_219 (O_219,N_2830,N_2959);
and UO_220 (O_220,N_2936,N_2824);
nand UO_221 (O_221,N_2838,N_2990);
or UO_222 (O_222,N_2919,N_2837);
nand UO_223 (O_223,N_2904,N_2805);
and UO_224 (O_224,N_2817,N_2847);
nor UO_225 (O_225,N_2888,N_2940);
or UO_226 (O_226,N_2810,N_2828);
and UO_227 (O_227,N_2894,N_2873);
xor UO_228 (O_228,N_2844,N_2932);
and UO_229 (O_229,N_2991,N_2903);
nor UO_230 (O_230,N_2875,N_2883);
or UO_231 (O_231,N_2898,N_2954);
or UO_232 (O_232,N_2844,N_2880);
nand UO_233 (O_233,N_2959,N_2805);
or UO_234 (O_234,N_2942,N_2887);
or UO_235 (O_235,N_2925,N_2934);
and UO_236 (O_236,N_2888,N_2884);
and UO_237 (O_237,N_2853,N_2811);
or UO_238 (O_238,N_2952,N_2880);
nor UO_239 (O_239,N_2808,N_2997);
or UO_240 (O_240,N_2907,N_2850);
nor UO_241 (O_241,N_2938,N_2962);
nor UO_242 (O_242,N_2814,N_2957);
xnor UO_243 (O_243,N_2828,N_2917);
and UO_244 (O_244,N_2806,N_2959);
xor UO_245 (O_245,N_2889,N_2901);
nor UO_246 (O_246,N_2918,N_2822);
xnor UO_247 (O_247,N_2861,N_2896);
xnor UO_248 (O_248,N_2918,N_2860);
nor UO_249 (O_249,N_2815,N_2832);
or UO_250 (O_250,N_2808,N_2957);
xnor UO_251 (O_251,N_2894,N_2954);
or UO_252 (O_252,N_2905,N_2909);
nand UO_253 (O_253,N_2853,N_2852);
xor UO_254 (O_254,N_2863,N_2801);
nor UO_255 (O_255,N_2818,N_2942);
or UO_256 (O_256,N_2962,N_2951);
and UO_257 (O_257,N_2872,N_2915);
nand UO_258 (O_258,N_2902,N_2968);
xnor UO_259 (O_259,N_2882,N_2921);
and UO_260 (O_260,N_2918,N_2881);
nand UO_261 (O_261,N_2938,N_2965);
xnor UO_262 (O_262,N_2850,N_2977);
nor UO_263 (O_263,N_2874,N_2843);
xor UO_264 (O_264,N_2884,N_2807);
and UO_265 (O_265,N_2911,N_2955);
or UO_266 (O_266,N_2837,N_2977);
or UO_267 (O_267,N_2956,N_2901);
nand UO_268 (O_268,N_2825,N_2841);
xnor UO_269 (O_269,N_2832,N_2840);
or UO_270 (O_270,N_2990,N_2952);
and UO_271 (O_271,N_2929,N_2858);
nand UO_272 (O_272,N_2937,N_2852);
or UO_273 (O_273,N_2961,N_2833);
nor UO_274 (O_274,N_2814,N_2930);
nor UO_275 (O_275,N_2984,N_2917);
or UO_276 (O_276,N_2893,N_2916);
nor UO_277 (O_277,N_2827,N_2866);
xor UO_278 (O_278,N_2825,N_2804);
or UO_279 (O_279,N_2976,N_2808);
xnor UO_280 (O_280,N_2901,N_2993);
nor UO_281 (O_281,N_2973,N_2856);
nor UO_282 (O_282,N_2867,N_2997);
nor UO_283 (O_283,N_2877,N_2914);
xnor UO_284 (O_284,N_2829,N_2994);
nor UO_285 (O_285,N_2836,N_2897);
or UO_286 (O_286,N_2833,N_2952);
nor UO_287 (O_287,N_2962,N_2985);
xnor UO_288 (O_288,N_2975,N_2979);
and UO_289 (O_289,N_2917,N_2937);
xnor UO_290 (O_290,N_2845,N_2906);
and UO_291 (O_291,N_2999,N_2910);
and UO_292 (O_292,N_2983,N_2802);
nand UO_293 (O_293,N_2904,N_2824);
xor UO_294 (O_294,N_2968,N_2898);
xnor UO_295 (O_295,N_2866,N_2823);
xnor UO_296 (O_296,N_2824,N_2820);
and UO_297 (O_297,N_2843,N_2977);
and UO_298 (O_298,N_2899,N_2838);
or UO_299 (O_299,N_2937,N_2993);
nor UO_300 (O_300,N_2984,N_2840);
nor UO_301 (O_301,N_2859,N_2873);
xnor UO_302 (O_302,N_2919,N_2974);
and UO_303 (O_303,N_2921,N_2978);
xor UO_304 (O_304,N_2978,N_2923);
nand UO_305 (O_305,N_2971,N_2926);
or UO_306 (O_306,N_2843,N_2971);
nand UO_307 (O_307,N_2968,N_2802);
nor UO_308 (O_308,N_2846,N_2956);
nor UO_309 (O_309,N_2905,N_2882);
nand UO_310 (O_310,N_2837,N_2824);
and UO_311 (O_311,N_2945,N_2946);
nand UO_312 (O_312,N_2996,N_2884);
or UO_313 (O_313,N_2815,N_2852);
or UO_314 (O_314,N_2842,N_2805);
or UO_315 (O_315,N_2897,N_2893);
or UO_316 (O_316,N_2960,N_2893);
nor UO_317 (O_317,N_2921,N_2906);
nor UO_318 (O_318,N_2966,N_2950);
xnor UO_319 (O_319,N_2824,N_2924);
or UO_320 (O_320,N_2894,N_2800);
xor UO_321 (O_321,N_2835,N_2953);
nand UO_322 (O_322,N_2809,N_2878);
nand UO_323 (O_323,N_2804,N_2981);
nand UO_324 (O_324,N_2960,N_2822);
nand UO_325 (O_325,N_2839,N_2902);
and UO_326 (O_326,N_2987,N_2943);
nor UO_327 (O_327,N_2858,N_2955);
nand UO_328 (O_328,N_2946,N_2944);
and UO_329 (O_329,N_2996,N_2893);
and UO_330 (O_330,N_2978,N_2935);
and UO_331 (O_331,N_2982,N_2845);
xor UO_332 (O_332,N_2842,N_2815);
nor UO_333 (O_333,N_2926,N_2948);
xnor UO_334 (O_334,N_2886,N_2824);
nor UO_335 (O_335,N_2808,N_2958);
xor UO_336 (O_336,N_2909,N_2958);
nor UO_337 (O_337,N_2860,N_2954);
nand UO_338 (O_338,N_2879,N_2938);
nor UO_339 (O_339,N_2805,N_2928);
xor UO_340 (O_340,N_2937,N_2877);
xnor UO_341 (O_341,N_2891,N_2841);
or UO_342 (O_342,N_2859,N_2864);
nor UO_343 (O_343,N_2894,N_2849);
nor UO_344 (O_344,N_2818,N_2915);
or UO_345 (O_345,N_2973,N_2995);
nand UO_346 (O_346,N_2845,N_2928);
nor UO_347 (O_347,N_2865,N_2947);
nand UO_348 (O_348,N_2868,N_2829);
and UO_349 (O_349,N_2962,N_2817);
xnor UO_350 (O_350,N_2832,N_2978);
nand UO_351 (O_351,N_2887,N_2915);
xor UO_352 (O_352,N_2954,N_2829);
nor UO_353 (O_353,N_2830,N_2966);
xnor UO_354 (O_354,N_2988,N_2895);
nand UO_355 (O_355,N_2805,N_2863);
and UO_356 (O_356,N_2957,N_2934);
xnor UO_357 (O_357,N_2999,N_2862);
nor UO_358 (O_358,N_2859,N_2906);
nand UO_359 (O_359,N_2891,N_2945);
nor UO_360 (O_360,N_2854,N_2862);
nor UO_361 (O_361,N_2894,N_2920);
nor UO_362 (O_362,N_2990,N_2986);
and UO_363 (O_363,N_2979,N_2873);
nor UO_364 (O_364,N_2907,N_2808);
and UO_365 (O_365,N_2888,N_2817);
nor UO_366 (O_366,N_2943,N_2858);
or UO_367 (O_367,N_2852,N_2895);
and UO_368 (O_368,N_2879,N_2905);
nor UO_369 (O_369,N_2822,N_2818);
and UO_370 (O_370,N_2815,N_2911);
or UO_371 (O_371,N_2889,N_2861);
nor UO_372 (O_372,N_2819,N_2896);
xnor UO_373 (O_373,N_2803,N_2897);
and UO_374 (O_374,N_2950,N_2884);
nor UO_375 (O_375,N_2855,N_2867);
nand UO_376 (O_376,N_2914,N_2991);
nand UO_377 (O_377,N_2916,N_2857);
and UO_378 (O_378,N_2840,N_2852);
nand UO_379 (O_379,N_2934,N_2983);
and UO_380 (O_380,N_2890,N_2949);
xnor UO_381 (O_381,N_2804,N_2862);
xnor UO_382 (O_382,N_2924,N_2922);
nand UO_383 (O_383,N_2903,N_2937);
nor UO_384 (O_384,N_2958,N_2905);
xnor UO_385 (O_385,N_2865,N_2999);
and UO_386 (O_386,N_2852,N_2992);
or UO_387 (O_387,N_2857,N_2950);
xnor UO_388 (O_388,N_2823,N_2996);
nor UO_389 (O_389,N_2951,N_2820);
or UO_390 (O_390,N_2839,N_2854);
nand UO_391 (O_391,N_2874,N_2988);
nand UO_392 (O_392,N_2819,N_2974);
nand UO_393 (O_393,N_2870,N_2909);
nand UO_394 (O_394,N_2809,N_2895);
nor UO_395 (O_395,N_2934,N_2911);
nand UO_396 (O_396,N_2804,N_2946);
and UO_397 (O_397,N_2811,N_2905);
or UO_398 (O_398,N_2994,N_2821);
xnor UO_399 (O_399,N_2835,N_2836);
xor UO_400 (O_400,N_2829,N_2903);
xor UO_401 (O_401,N_2877,N_2870);
or UO_402 (O_402,N_2924,N_2992);
xor UO_403 (O_403,N_2834,N_2820);
or UO_404 (O_404,N_2800,N_2837);
or UO_405 (O_405,N_2914,N_2957);
or UO_406 (O_406,N_2920,N_2967);
nand UO_407 (O_407,N_2909,N_2901);
or UO_408 (O_408,N_2879,N_2934);
nand UO_409 (O_409,N_2867,N_2885);
nand UO_410 (O_410,N_2957,N_2844);
nand UO_411 (O_411,N_2971,N_2956);
xor UO_412 (O_412,N_2843,N_2881);
nor UO_413 (O_413,N_2887,N_2940);
nor UO_414 (O_414,N_2887,N_2897);
nor UO_415 (O_415,N_2819,N_2976);
xnor UO_416 (O_416,N_2969,N_2852);
or UO_417 (O_417,N_2986,N_2869);
nor UO_418 (O_418,N_2870,N_2932);
or UO_419 (O_419,N_2846,N_2847);
nand UO_420 (O_420,N_2808,N_2932);
and UO_421 (O_421,N_2930,N_2969);
nand UO_422 (O_422,N_2875,N_2971);
or UO_423 (O_423,N_2939,N_2940);
nand UO_424 (O_424,N_2833,N_2871);
and UO_425 (O_425,N_2990,N_2803);
or UO_426 (O_426,N_2975,N_2886);
xor UO_427 (O_427,N_2808,N_2838);
xor UO_428 (O_428,N_2974,N_2903);
xnor UO_429 (O_429,N_2832,N_2822);
nor UO_430 (O_430,N_2856,N_2935);
or UO_431 (O_431,N_2856,N_2929);
or UO_432 (O_432,N_2821,N_2857);
nor UO_433 (O_433,N_2865,N_2889);
nand UO_434 (O_434,N_2846,N_2992);
nand UO_435 (O_435,N_2847,N_2801);
nor UO_436 (O_436,N_2990,N_2837);
xor UO_437 (O_437,N_2942,N_2911);
xnor UO_438 (O_438,N_2963,N_2908);
nand UO_439 (O_439,N_2867,N_2859);
nor UO_440 (O_440,N_2967,N_2828);
xor UO_441 (O_441,N_2893,N_2870);
nor UO_442 (O_442,N_2850,N_2938);
xor UO_443 (O_443,N_2957,N_2990);
nand UO_444 (O_444,N_2908,N_2924);
or UO_445 (O_445,N_2979,N_2865);
and UO_446 (O_446,N_2968,N_2946);
nor UO_447 (O_447,N_2916,N_2923);
nor UO_448 (O_448,N_2974,N_2951);
xor UO_449 (O_449,N_2957,N_2871);
and UO_450 (O_450,N_2878,N_2992);
xnor UO_451 (O_451,N_2825,N_2879);
and UO_452 (O_452,N_2889,N_2879);
or UO_453 (O_453,N_2944,N_2829);
nand UO_454 (O_454,N_2828,N_2995);
nand UO_455 (O_455,N_2860,N_2986);
xor UO_456 (O_456,N_2974,N_2830);
and UO_457 (O_457,N_2948,N_2882);
nand UO_458 (O_458,N_2907,N_2938);
nor UO_459 (O_459,N_2979,N_2915);
and UO_460 (O_460,N_2851,N_2859);
nand UO_461 (O_461,N_2967,N_2874);
nor UO_462 (O_462,N_2903,N_2837);
and UO_463 (O_463,N_2805,N_2819);
or UO_464 (O_464,N_2844,N_2979);
xor UO_465 (O_465,N_2841,N_2987);
nand UO_466 (O_466,N_2945,N_2806);
or UO_467 (O_467,N_2832,N_2904);
or UO_468 (O_468,N_2892,N_2964);
nand UO_469 (O_469,N_2991,N_2995);
nand UO_470 (O_470,N_2888,N_2942);
or UO_471 (O_471,N_2906,N_2813);
nand UO_472 (O_472,N_2927,N_2960);
and UO_473 (O_473,N_2963,N_2942);
or UO_474 (O_474,N_2959,N_2970);
xor UO_475 (O_475,N_2902,N_2859);
nand UO_476 (O_476,N_2816,N_2863);
nand UO_477 (O_477,N_2920,N_2837);
nor UO_478 (O_478,N_2899,N_2871);
or UO_479 (O_479,N_2864,N_2978);
xnor UO_480 (O_480,N_2867,N_2950);
and UO_481 (O_481,N_2833,N_2925);
and UO_482 (O_482,N_2841,N_2864);
and UO_483 (O_483,N_2961,N_2835);
nor UO_484 (O_484,N_2839,N_2922);
xor UO_485 (O_485,N_2980,N_2925);
or UO_486 (O_486,N_2910,N_2846);
nor UO_487 (O_487,N_2992,N_2867);
nor UO_488 (O_488,N_2884,N_2974);
nand UO_489 (O_489,N_2892,N_2826);
nor UO_490 (O_490,N_2993,N_2928);
or UO_491 (O_491,N_2808,N_2928);
and UO_492 (O_492,N_2921,N_2801);
and UO_493 (O_493,N_2802,N_2978);
and UO_494 (O_494,N_2871,N_2932);
xnor UO_495 (O_495,N_2998,N_2961);
xnor UO_496 (O_496,N_2863,N_2814);
and UO_497 (O_497,N_2872,N_2892);
or UO_498 (O_498,N_2874,N_2985);
and UO_499 (O_499,N_2990,N_2970);
endmodule