module basic_1500_15000_2000_20_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1237,In_1076);
nand U1 (N_1,In_1122,In_440);
xnor U2 (N_2,In_973,In_886);
nor U3 (N_3,In_801,In_201);
nand U4 (N_4,In_1058,In_741);
nand U5 (N_5,In_926,In_561);
nand U6 (N_6,In_542,In_112);
and U7 (N_7,In_160,In_580);
nand U8 (N_8,In_993,In_228);
nand U9 (N_9,In_1021,In_715);
and U10 (N_10,In_1196,In_1282);
and U11 (N_11,In_1267,In_1294);
or U12 (N_12,In_853,In_53);
and U13 (N_13,In_1264,In_498);
and U14 (N_14,In_121,In_579);
nor U15 (N_15,In_1050,In_383);
xor U16 (N_16,In_1379,In_170);
or U17 (N_17,In_394,In_562);
nor U18 (N_18,In_464,In_502);
nor U19 (N_19,In_279,In_677);
nand U20 (N_20,In_809,In_402);
nor U21 (N_21,In_24,In_1391);
nor U22 (N_22,In_574,In_654);
and U23 (N_23,In_636,In_255);
and U24 (N_24,In_524,In_172);
or U25 (N_25,In_581,In_213);
and U26 (N_26,In_180,In_839);
xnor U27 (N_27,In_164,In_352);
and U28 (N_28,In_1159,In_1182);
nor U29 (N_29,In_601,In_1317);
and U30 (N_30,In_1003,In_612);
xnor U31 (N_31,In_1401,In_28);
nand U32 (N_32,In_882,In_635);
nor U33 (N_33,In_348,In_214);
or U34 (N_34,In_531,In_1092);
or U35 (N_35,In_1252,In_1350);
or U36 (N_36,In_1372,In_1309);
nand U37 (N_37,In_560,In_1449);
nand U38 (N_38,In_1219,In_439);
and U39 (N_39,In_1250,In_902);
nand U40 (N_40,In_567,In_43);
or U41 (N_41,In_659,In_752);
nand U42 (N_42,In_1285,In_400);
nand U43 (N_43,In_1094,In_1130);
and U44 (N_44,In_1157,In_983);
nand U45 (N_45,In_218,In_924);
nand U46 (N_46,In_588,In_624);
nor U47 (N_47,In_1344,In_1007);
or U48 (N_48,In_869,In_1180);
and U49 (N_49,In_821,In_666);
or U50 (N_50,In_235,In_35);
or U51 (N_51,In_1263,In_503);
and U52 (N_52,In_1331,In_1479);
nor U53 (N_53,In_763,In_1240);
nand U54 (N_54,In_1428,In_1451);
and U55 (N_55,In_547,In_97);
nor U56 (N_56,In_1319,In_1189);
nand U57 (N_57,In_951,In_1225);
or U58 (N_58,In_594,In_253);
or U59 (N_59,In_685,In_1367);
and U60 (N_60,In_340,In_1418);
and U61 (N_61,In_205,In_47);
and U62 (N_62,In_906,In_1412);
and U63 (N_63,In_663,In_1275);
or U64 (N_64,In_232,In_1467);
and U65 (N_65,In_974,In_37);
nor U66 (N_66,In_1466,In_1483);
nand U67 (N_67,In_1055,In_1233);
or U68 (N_68,In_700,In_306);
nor U69 (N_69,In_449,In_41);
xnor U70 (N_70,In_534,In_1325);
nor U71 (N_71,In_1380,In_392);
nand U72 (N_72,In_1171,In_1475);
and U73 (N_73,In_835,In_1290);
or U74 (N_74,In_1016,In_703);
or U75 (N_75,In_461,In_1060);
nand U76 (N_76,In_958,In_391);
or U77 (N_77,In_173,In_142);
nor U78 (N_78,In_1232,In_1051);
xnor U79 (N_79,In_852,In_327);
and U80 (N_80,In_146,In_591);
nor U81 (N_81,In_740,In_1400);
nand U82 (N_82,In_810,In_55);
or U83 (N_83,In_442,In_425);
nand U84 (N_84,In_1480,In_1280);
xnor U85 (N_85,In_458,In_589);
or U86 (N_86,In_797,In_686);
nand U87 (N_87,In_713,In_538);
or U88 (N_88,In_1167,In_825);
and U89 (N_89,In_489,In_476);
nor U90 (N_90,In_336,In_631);
or U91 (N_91,In_424,In_488);
nand U92 (N_92,In_1072,In_64);
nor U93 (N_93,In_288,In_280);
and U94 (N_94,In_62,In_1213);
or U95 (N_95,In_275,In_66);
nand U96 (N_96,In_1373,In_381);
or U97 (N_97,In_1463,In_429);
nand U98 (N_98,In_333,In_1408);
and U99 (N_99,In_506,In_59);
or U100 (N_100,In_959,In_908);
xor U101 (N_101,In_246,In_1460);
or U102 (N_102,In_571,In_806);
nor U103 (N_103,In_63,In_1487);
and U104 (N_104,In_698,In_312);
nand U105 (N_105,In_1396,In_1289);
or U106 (N_106,In_1382,In_915);
nand U107 (N_107,In_99,In_229);
nand U108 (N_108,In_1310,In_682);
or U109 (N_109,In_911,In_107);
nand U110 (N_110,In_271,In_161);
nor U111 (N_111,In_154,In_38);
nor U112 (N_112,In_1018,In_423);
nor U113 (N_113,In_578,In_748);
nand U114 (N_114,In_1450,In_947);
or U115 (N_115,In_536,In_840);
xnor U116 (N_116,In_153,In_1015);
nand U117 (N_117,In_241,In_1198);
nor U118 (N_118,In_380,In_625);
nand U119 (N_119,In_360,In_26);
nor U120 (N_120,In_1151,In_215);
nand U121 (N_121,In_4,In_1298);
xor U122 (N_122,In_233,In_1358);
xor U123 (N_123,In_89,In_377);
xor U124 (N_124,In_1312,In_484);
or U125 (N_125,In_614,In_653);
nand U126 (N_126,In_359,In_788);
nand U127 (N_127,In_1438,In_769);
nor U128 (N_128,In_1381,In_830);
nor U129 (N_129,In_1153,In_699);
nand U130 (N_130,In_71,In_927);
nand U131 (N_131,In_971,In_526);
nand U132 (N_132,In_443,In_436);
nand U133 (N_133,In_1357,In_238);
and U134 (N_134,In_1215,In_501);
and U135 (N_135,In_1262,In_1404);
xnor U136 (N_136,In_45,In_1226);
and U137 (N_137,In_687,In_943);
or U138 (N_138,In_249,In_242);
nor U139 (N_139,In_963,In_1395);
nor U140 (N_140,In_986,In_1286);
and U141 (N_141,In_1207,In_660);
xor U142 (N_142,In_912,In_873);
nand U143 (N_143,In_168,In_1394);
nor U144 (N_144,In_1332,In_451);
or U145 (N_145,In_118,In_925);
or U146 (N_146,In_1112,In_1083);
xnor U147 (N_147,In_874,In_1389);
and U148 (N_148,In_1138,In_731);
nor U149 (N_149,In_1097,In_679);
and U150 (N_150,In_1136,In_1370);
or U151 (N_151,In_866,In_495);
or U152 (N_152,In_726,In_899);
and U153 (N_153,In_638,In_468);
and U154 (N_154,In_88,In_34);
nor U155 (N_155,In_15,In_5);
and U156 (N_156,In_353,In_1354);
xnor U157 (N_157,In_262,In_174);
nor U158 (N_158,In_1413,In_395);
xor U159 (N_159,In_1469,In_905);
or U160 (N_160,In_937,In_1340);
and U161 (N_161,In_1301,In_568);
nand U162 (N_162,In_437,In_554);
or U163 (N_163,In_74,In_764);
and U164 (N_164,In_1239,In_387);
nor U165 (N_165,In_1246,In_725);
nor U166 (N_166,In_950,In_895);
nand U167 (N_167,In_655,In_1447);
nor U168 (N_168,In_696,In_692);
nor U169 (N_169,In_244,In_234);
or U170 (N_170,In_616,In_247);
and U171 (N_171,In_1063,In_504);
and U172 (N_172,In_193,In_1407);
and U173 (N_173,In_697,In_847);
or U174 (N_174,In_431,In_1231);
nor U175 (N_175,In_789,In_1496);
nand U176 (N_176,In_220,In_1427);
or U177 (N_177,In_152,In_850);
and U178 (N_178,In_441,In_586);
and U179 (N_179,In_1091,In_1067);
nor U180 (N_180,In_329,In_465);
nand U181 (N_181,In_628,In_206);
or U182 (N_182,In_1293,In_264);
xor U183 (N_183,In_841,In_409);
and U184 (N_184,In_1303,In_1028);
and U185 (N_185,In_1208,In_326);
xor U186 (N_186,In_732,In_1045);
nor U187 (N_187,In_1376,In_289);
nand U188 (N_188,In_888,In_1202);
and U189 (N_189,In_137,In_1353);
nand U190 (N_190,In_1339,In_1123);
nor U191 (N_191,In_1452,In_1295);
nor U192 (N_192,In_1161,In_1070);
and U193 (N_193,In_491,In_401);
nand U194 (N_194,In_1378,In_463);
nand U195 (N_195,In_1305,In_608);
or U196 (N_196,In_122,In_1175);
or U197 (N_197,In_781,In_1361);
or U198 (N_198,In_413,In_1271);
nand U199 (N_199,In_192,In_106);
nand U200 (N_200,In_1000,In_1214);
and U201 (N_201,In_1356,In_661);
xnor U202 (N_202,In_139,In_827);
and U203 (N_203,In_389,In_833);
or U204 (N_204,In_254,In_1048);
and U205 (N_205,In_634,In_68);
nor U206 (N_206,In_683,In_668);
nand U207 (N_207,In_155,In_949);
or U208 (N_208,In_640,In_662);
or U209 (N_209,In_1406,In_1477);
xor U210 (N_210,In_548,In_399);
nand U211 (N_211,In_179,In_119);
nand U212 (N_212,In_1120,In_277);
or U213 (N_213,In_721,In_990);
nor U214 (N_214,In_643,In_1056);
nand U215 (N_215,In_315,In_954);
or U216 (N_216,In_1052,In_157);
nand U217 (N_217,In_1326,In_985);
nor U218 (N_218,In_1169,In_317);
nor U219 (N_219,In_551,In_1149);
nand U220 (N_220,In_197,In_1080);
nand U221 (N_221,In_1465,In_1086);
nor U222 (N_222,In_343,In_273);
xor U223 (N_223,In_863,In_604);
nand U224 (N_224,In_1446,In_276);
or U225 (N_225,In_658,In_573);
nand U226 (N_226,In_783,In_596);
or U227 (N_227,In_76,In_1490);
and U228 (N_228,In_421,In_298);
and U229 (N_229,In_310,In_1435);
and U230 (N_230,In_1088,In_1387);
and U231 (N_231,In_362,In_1492);
nor U232 (N_232,In_1318,In_1106);
or U233 (N_233,In_1314,In_60);
and U234 (N_234,In_1145,In_1456);
nor U235 (N_235,In_975,In_1440);
or U236 (N_236,In_258,In_822);
and U237 (N_237,In_135,In_1069);
or U238 (N_238,In_1012,In_17);
and U239 (N_239,In_1040,In_309);
or U240 (N_240,In_508,In_140);
or U241 (N_241,In_272,In_541);
or U242 (N_242,In_21,In_1118);
and U243 (N_243,In_1075,In_1448);
or U244 (N_244,In_1244,In_528);
xor U245 (N_245,In_646,In_1115);
and U246 (N_246,In_630,In_1436);
xnor U247 (N_247,In_885,In_434);
nor U248 (N_248,In_544,In_566);
or U249 (N_249,In_350,In_1363);
or U250 (N_250,In_188,In_1107);
nand U251 (N_251,In_744,In_1030);
and U252 (N_252,In_545,In_456);
nor U253 (N_253,In_1093,In_811);
nor U254 (N_254,In_42,In_1488);
and U255 (N_255,In_445,In_1316);
and U256 (N_256,In_1422,In_1129);
nor U257 (N_257,In_478,In_2);
nand U258 (N_258,In_607,In_1336);
nor U259 (N_259,In_933,In_1243);
nor U260 (N_260,In_1186,In_1270);
nor U261 (N_261,In_1137,In_30);
nand U262 (N_262,In_1307,In_318);
nand U263 (N_263,In_123,In_1494);
nor U264 (N_264,In_1306,In_1334);
nand U265 (N_265,In_406,In_988);
and U266 (N_266,In_470,In_95);
nor U267 (N_267,In_982,In_962);
and U268 (N_268,In_946,In_1328);
xor U269 (N_269,In_460,In_270);
nor U270 (N_270,In_10,In_323);
and U271 (N_271,In_1064,In_556);
nor U272 (N_272,In_370,In_376);
nor U273 (N_273,In_162,In_1143);
nand U274 (N_274,In_1062,In_760);
nand U275 (N_275,In_1269,In_371);
or U276 (N_276,In_824,In_1061);
nor U277 (N_277,In_104,In_375);
or U278 (N_278,In_584,In_1241);
and U279 (N_279,In_1236,In_710);
nor U280 (N_280,In_519,In_1096);
and U281 (N_281,In_832,In_332);
xnor U282 (N_282,In_1338,In_997);
nand U283 (N_283,In_396,In_1148);
nor U284 (N_284,In_770,In_382);
nand U285 (N_285,In_267,In_970);
xor U286 (N_286,In_743,In_539);
and U287 (N_287,In_8,In_674);
nand U288 (N_288,In_1320,In_284);
nor U289 (N_289,In_848,In_452);
and U290 (N_290,In_991,In_956);
or U291 (N_291,In_1065,In_1304);
xnor U292 (N_292,In_403,In_469);
xnor U293 (N_293,In_311,In_656);
nor U294 (N_294,In_415,In_1499);
nand U295 (N_295,In_115,In_163);
and U296 (N_296,In_230,In_1081);
and U297 (N_297,In_49,In_1265);
and U298 (N_298,In_1368,In_292);
or U299 (N_299,In_819,In_736);
nand U300 (N_300,In_290,In_619);
nor U301 (N_301,In_261,In_1375);
and U302 (N_302,In_1197,In_1119);
nand U303 (N_303,In_149,In_379);
and U304 (N_304,In_945,In_194);
nor U305 (N_305,In_795,In_285);
and U306 (N_306,In_471,In_676);
nand U307 (N_307,In_649,In_918);
nor U308 (N_308,In_404,In_533);
xnor U309 (N_309,In_598,In_776);
nand U310 (N_310,In_1009,In_175);
or U311 (N_311,In_747,In_56);
or U312 (N_312,In_397,In_871);
nand U313 (N_313,In_922,In_1187);
nor U314 (N_314,In_892,In_1194);
nor U315 (N_315,In_87,In_1455);
or U316 (N_316,In_268,In_1433);
nor U317 (N_317,In_1409,In_590);
and U318 (N_318,In_1031,In_1308);
and U319 (N_319,In_691,In_1471);
nor U320 (N_320,In_855,In_535);
or U321 (N_321,In_664,In_936);
and U322 (N_322,In_82,In_46);
or U323 (N_323,In_147,In_729);
or U324 (N_324,In_693,In_678);
or U325 (N_325,In_932,In_921);
nand U326 (N_326,In_369,In_1392);
nand U327 (N_327,In_367,In_938);
or U328 (N_328,In_358,In_1321);
and U329 (N_329,In_314,In_1493);
nand U330 (N_330,In_1013,In_890);
and U331 (N_331,In_1330,In_51);
nor U332 (N_332,In_878,In_1209);
or U333 (N_333,In_393,In_1481);
nand U334 (N_334,In_386,In_645);
or U335 (N_335,In_1417,In_319);
or U336 (N_336,In_1327,In_792);
or U337 (N_337,In_78,In_111);
nor U338 (N_338,In_475,In_1168);
or U339 (N_339,In_812,In_512);
nand U340 (N_340,In_1079,In_225);
nor U341 (N_341,In_1364,In_1287);
nor U342 (N_342,In_1181,In_1385);
and U343 (N_343,In_293,In_72);
nand U344 (N_344,In_1221,In_239);
or U345 (N_345,In_1014,In_1335);
or U346 (N_346,In_1443,In_880);
nand U347 (N_347,In_784,In_320);
or U348 (N_348,In_815,In_485);
nor U349 (N_349,In_704,In_647);
or U350 (N_350,In_1283,In_553);
nand U351 (N_351,In_1360,In_257);
and U352 (N_352,In_1324,In_86);
xnor U353 (N_353,In_1084,In_109);
and U354 (N_354,In_689,In_240);
xor U355 (N_355,In_939,In_928);
nand U356 (N_356,In_1172,In_999);
nand U357 (N_357,In_462,In_416);
or U358 (N_358,In_1104,In_1468);
nor U359 (N_359,In_1152,In_39);
nand U360 (N_360,In_877,In_1008);
and U361 (N_361,In_883,In_1195);
nand U362 (N_362,In_339,In_1017);
nand U363 (N_363,In_669,In_209);
or U364 (N_364,In_373,In_1);
or U365 (N_365,In_181,In_1054);
or U366 (N_366,In_136,In_1497);
nand U367 (N_367,In_116,In_802);
and U368 (N_368,In_117,In_1365);
and U369 (N_369,In_25,In_595);
nor U370 (N_370,In_1371,In_1082);
or U371 (N_371,In_1032,In_221);
nand U372 (N_372,In_808,In_1457);
or U373 (N_373,In_870,In_1205);
or U374 (N_374,In_223,In_510);
xnor U375 (N_375,In_414,In_735);
or U376 (N_376,In_20,In_817);
or U377 (N_377,In_641,In_294);
and U378 (N_378,In_879,In_305);
and U379 (N_379,In_22,In_374);
or U380 (N_380,In_1006,In_1258);
or U381 (N_381,In_361,In_1421);
nand U382 (N_382,In_1473,In_884);
xnor U383 (N_383,In_786,In_486);
xnor U384 (N_384,In_1279,In_477);
nand U385 (N_385,In_411,In_995);
nor U386 (N_386,In_718,In_552);
xnor U387 (N_387,In_65,In_479);
nor U388 (N_388,In_303,In_1484);
nor U389 (N_389,In_1235,In_1087);
nor U390 (N_390,In_1095,In_845);
nor U391 (N_391,In_1053,In_701);
nor U392 (N_392,In_648,In_831);
and U393 (N_393,In_826,In_75);
or U394 (N_394,In_250,In_849);
xnor U395 (N_395,In_961,In_1423);
xor U396 (N_396,In_794,In_347);
or U397 (N_397,In_1333,In_448);
xnor U398 (N_398,In_1255,In_900);
and U399 (N_399,In_1177,In_101);
or U400 (N_400,In_966,In_198);
xnor U401 (N_401,In_1253,In_265);
and U402 (N_402,In_793,In_1109);
nor U403 (N_403,In_520,In_1458);
nand U404 (N_404,In_1453,In_259);
or U405 (N_405,In_245,In_365);
xnor U406 (N_406,In_733,In_1134);
nand U407 (N_407,In_587,In_739);
nor U408 (N_408,In_19,In_868);
nand U409 (N_409,In_1281,In_1284);
or U410 (N_410,In_430,In_838);
or U411 (N_411,In_1128,In_513);
nand U412 (N_412,In_466,In_295);
xor U413 (N_413,In_167,In_1291);
nor U414 (N_414,In_299,In_762);
and U415 (N_415,In_978,In_603);
xnor U416 (N_416,In_728,In_785);
nor U417 (N_417,In_1355,In_521);
and U418 (N_418,In_183,In_858);
or U419 (N_419,In_260,In_1043);
nor U420 (N_420,In_860,In_18);
or U421 (N_421,In_199,In_1323);
and U422 (N_422,In_576,In_837);
or U423 (N_423,In_420,In_190);
or U424 (N_424,In_195,In_211);
and U425 (N_425,In_328,In_1147);
and U426 (N_426,In_1098,In_1261);
and U427 (N_427,In_690,In_722);
and U428 (N_428,In_1170,In_694);
or U429 (N_429,In_1230,In_1437);
xor U430 (N_430,In_120,In_186);
and U431 (N_431,In_976,In_6);
nand U432 (N_432,In_564,In_671);
xor U433 (N_433,In_203,In_405);
nor U434 (N_434,In_818,In_1276);
nor U435 (N_435,In_334,In_550);
nand U436 (N_436,In_308,In_889);
or U437 (N_437,In_345,In_1005);
nand U438 (N_438,In_1251,In_1229);
or U439 (N_439,In_1036,In_1139);
nand U440 (N_440,In_942,In_58);
nand U441 (N_441,In_1211,In_525);
or U442 (N_442,In_929,In_1278);
or U443 (N_443,In_1482,In_861);
xnor U444 (N_444,In_1162,In_9);
and U445 (N_445,In_92,In_569);
and U446 (N_446,In_745,In_517);
nor U447 (N_447,In_31,In_398);
or U448 (N_448,In_427,In_1414);
nand U449 (N_449,In_208,In_844);
xnor U450 (N_450,In_901,In_919);
or U451 (N_451,In_113,In_316);
or U452 (N_452,In_1459,In_1200);
or U453 (N_453,In_633,In_166);
and U454 (N_454,In_1248,In_665);
nand U455 (N_455,In_1210,In_807);
and U456 (N_456,In_130,In_952);
nand U457 (N_457,In_557,In_856);
nor U458 (N_458,In_150,In_158);
or U459 (N_459,In_977,In_1410);
or U460 (N_460,In_1026,In_1131);
and U461 (N_461,In_941,In_1216);
and U462 (N_462,In_1001,In_251);
or U463 (N_463,In_714,In_759);
or U464 (N_464,In_105,In_355);
nand U465 (N_465,In_989,In_313);
and U466 (N_466,In_620,In_138);
and U467 (N_467,In_610,In_287);
nand U468 (N_468,In_1133,In_1224);
nand U469 (N_469,In_1302,In_1126);
xnor U470 (N_470,In_820,In_582);
and U471 (N_471,In_1037,In_307);
and U472 (N_472,In_1292,In_1166);
or U473 (N_473,In_16,In_1204);
nand U474 (N_474,In_304,In_1041);
or U475 (N_475,In_1351,In_1039);
nor U476 (N_476,In_335,In_1445);
nand U477 (N_477,In_1329,In_459);
nand U478 (N_478,In_737,In_492);
nand U479 (N_479,In_438,In_734);
or U480 (N_480,In_768,In_1415);
and U481 (N_481,In_243,In_300);
nor U482 (N_482,In_1135,In_44);
xor U483 (N_483,In_1274,In_621);
nor U484 (N_484,In_708,In_497);
or U485 (N_485,In_412,In_216);
nand U486 (N_486,In_632,In_1156);
or U487 (N_487,In_1117,In_823);
or U488 (N_488,In_772,In_706);
xor U489 (N_489,In_1245,In_499);
nand U490 (N_490,In_865,In_720);
nor U491 (N_491,In_1399,In_90);
nor U492 (N_492,In_1193,In_227);
and U493 (N_493,In_1142,In_337);
or U494 (N_494,In_935,In_1322);
and U495 (N_495,In_1154,In_532);
or U496 (N_496,In_418,In_684);
nand U497 (N_497,In_719,In_1257);
nand U498 (N_498,In_955,In_224);
and U499 (N_499,In_207,In_61);
nand U500 (N_500,In_1454,In_1403);
nor U501 (N_501,In_965,In_368);
nand U502 (N_502,In_1174,In_707);
and U503 (N_503,In_930,In_1090);
nor U504 (N_504,In_887,In_182);
and U505 (N_505,In_602,In_23);
or U506 (N_506,In_617,In_1116);
nor U507 (N_507,In_615,In_1405);
and U508 (N_508,In_126,In_1259);
nand U509 (N_509,In_1495,In_964);
and U510 (N_510,In_572,In_81);
nor U511 (N_511,In_67,In_558);
and U512 (N_512,In_366,In_108);
and U513 (N_513,In_1398,In_750);
nand U514 (N_514,In_148,In_1188);
nand U515 (N_515,In_1374,In_779);
or U516 (N_516,In_1068,In_1206);
nor U517 (N_517,In_842,In_480);
or U518 (N_518,In_1266,In_454);
nand U519 (N_519,In_231,In_1038);
nand U520 (N_520,In_291,In_297);
nor U521 (N_521,In_673,In_1393);
nor U522 (N_522,In_143,In_266);
or U523 (N_523,In_85,In_1110);
and U524 (N_524,In_593,In_296);
nor U525 (N_525,In_344,In_1311);
nor U526 (N_526,In_496,In_522);
or U527 (N_527,In_846,In_27);
or U528 (N_528,In_771,In_618);
nor U529 (N_529,In_1027,In_1173);
or U530 (N_530,In_867,In_252);
or U531 (N_531,In_13,In_944);
nand U532 (N_532,In_226,In_749);
nand U533 (N_533,In_1066,In_1397);
nand U534 (N_534,In_667,In_960);
nand U535 (N_535,In_1288,In_1431);
nor U536 (N_536,In_1247,In_407);
or U537 (N_537,In_914,In_1077);
and U538 (N_538,In_549,In_324);
or U539 (N_539,In_829,In_1299);
nand U540 (N_540,In_1191,In_482);
and U541 (N_541,In_354,In_796);
xnor U542 (N_542,In_171,In_1461);
nand U543 (N_543,In_803,In_1074);
nor U544 (N_544,In_1462,In_3);
xnor U545 (N_545,In_1300,In_992);
or U546 (N_546,In_269,In_1071);
and U547 (N_547,In_875,In_184);
or U548 (N_548,In_891,In_12);
nand U549 (N_549,In_644,In_356);
or U550 (N_550,In_507,In_1089);
or U551 (N_551,In_864,In_727);
nor U552 (N_552,In_800,In_73);
or U553 (N_553,In_494,In_798);
and U554 (N_554,In_1019,In_453);
nor U555 (N_555,In_514,In_1025);
xnor U556 (N_556,In_1165,In_96);
and U557 (N_557,In_876,In_490);
or U558 (N_558,In_1044,In_1124);
and U559 (N_559,In_605,In_474);
nand U560 (N_560,In_191,In_1155);
nand U561 (N_561,In_1029,In_1059);
and U562 (N_562,In_1121,In_263);
nand U563 (N_563,In_537,In_799);
nand U564 (N_564,In_79,In_1046);
or U565 (N_565,In_1268,In_642);
nand U566 (N_566,In_834,In_432);
and U567 (N_567,In_103,In_622);
nor U568 (N_568,In_907,In_1425);
xor U569 (N_569,In_48,In_765);
and U570 (N_570,In_493,In_114);
xor U571 (N_571,In_688,In_652);
nor U572 (N_572,In_1315,In_282);
nor U573 (N_573,In_1430,In_1100);
or U574 (N_574,In_1313,In_1383);
or U575 (N_575,In_1158,In_222);
nor U576 (N_576,In_1419,In_1132);
and U577 (N_577,In_859,In_321);
nand U578 (N_578,In_724,In_934);
xnor U579 (N_579,In_712,In_196);
nand U580 (N_580,In_1343,In_364);
nor U581 (N_581,In_1420,In_705);
and U582 (N_582,In_523,In_349);
or U583 (N_583,In_331,In_898);
nand U584 (N_584,In_330,In_1369);
nand U585 (N_585,In_896,In_388);
or U586 (N_586,In_378,In_1201);
nand U587 (N_587,In_210,In_156);
nor U588 (N_588,In_372,In_816);
and U589 (N_589,In_422,In_773);
and U590 (N_590,In_435,In_144);
nand U591 (N_591,In_505,In_133);
nand U592 (N_592,In_854,In_637);
nor U593 (N_593,In_894,In_917);
nor U594 (N_594,In_1042,In_237);
or U595 (N_595,In_670,In_626);
nor U596 (N_596,In_1078,In_1192);
and U597 (N_597,In_217,In_177);
nand U598 (N_598,In_843,In_1146);
or U599 (N_599,In_29,In_1296);
or U600 (N_600,In_592,In_1256);
nand U601 (N_601,In_127,In_385);
and U602 (N_602,In_248,In_131);
and U603 (N_603,In_923,In_984);
or U604 (N_604,In_657,In_755);
or U605 (N_605,In_1099,In_419);
or U606 (N_606,In_599,In_623);
xnor U607 (N_607,In_169,In_200);
and U608 (N_608,In_1183,In_212);
xnor U609 (N_609,In_851,In_639);
nand U610 (N_610,In_50,In_204);
xnor U611 (N_611,In_555,In_36);
nor U612 (N_612,In_1238,In_836);
nand U613 (N_613,In_1476,In_1002);
or U614 (N_614,In_7,In_1352);
and U615 (N_615,In_1345,In_1424);
or U616 (N_616,In_910,In_1273);
or U617 (N_617,In_627,In_857);
nor U618 (N_618,In_408,In_1491);
xor U619 (N_619,In_675,In_1176);
nand U620 (N_620,In_680,In_278);
or U621 (N_621,In_1341,In_1349);
nand U622 (N_622,In_909,In_70);
and U623 (N_623,In_342,In_473);
nor U624 (N_624,In_1004,In_1472);
nor U625 (N_625,In_1441,In_746);
nor U626 (N_626,In_758,In_1234);
or U627 (N_627,In_948,In_546);
nor U628 (N_628,In_1203,In_57);
nand U629 (N_629,In_609,In_1434);
xnor U630 (N_630,In_433,In_487);
xnor U631 (N_631,In_996,In_530);
nor U632 (N_632,In_681,In_1164);
and U633 (N_633,In_583,In_1185);
or U634 (N_634,In_187,In_1444);
or U635 (N_635,In_518,In_1140);
and U636 (N_636,In_467,In_1402);
or U637 (N_637,In_600,In_1432);
nor U638 (N_638,In_69,In_1478);
or U639 (N_639,In_426,In_1111);
xor U640 (N_640,In_428,In_527);
nand U641 (N_641,In_813,In_322);
nand U642 (N_642,In_695,In_565);
nand U643 (N_643,In_1362,In_1297);
or U644 (N_644,In_1103,In_767);
xnor U645 (N_645,In_189,In_102);
nor U646 (N_646,In_597,In_1470);
or U647 (N_647,In_346,In_145);
nand U648 (N_648,In_93,In_1217);
and U649 (N_649,In_987,In_611);
and U650 (N_650,In_511,In_446);
nor U651 (N_651,In_650,In_1227);
or U652 (N_652,In_1022,In_1249);
and U653 (N_653,In_1073,In_417);
nand U654 (N_654,In_341,In_742);
or U655 (N_655,In_363,In_998);
and U656 (N_656,In_351,In_100);
nand U657 (N_657,In_515,In_577);
or U658 (N_658,In_83,In_165);
and U659 (N_659,In_32,In_457);
and U660 (N_660,In_357,In_450);
xnor U661 (N_661,In_1085,In_1464);
nand U662 (N_662,In_1034,In_957);
xnor U663 (N_663,In_159,In_1047);
nor U664 (N_664,In_1439,In_0);
xnor U665 (N_665,In_94,In_1163);
or U666 (N_666,In_738,In_301);
nor U667 (N_667,In_125,In_1035);
or U668 (N_668,In_969,In_1426);
or U669 (N_669,In_1178,In_730);
nor U670 (N_670,In_1489,In_980);
xor U671 (N_671,In_1212,In_286);
xnor U672 (N_672,In_994,In_711);
nand U673 (N_673,In_968,In_1485);
nor U674 (N_674,In_1160,In_132);
and U675 (N_675,In_516,In_709);
nor U676 (N_676,In_1220,In_753);
nor U677 (N_677,In_1144,In_570);
nand U678 (N_678,In_1390,In_872);
nor U679 (N_679,In_606,In_1254);
or U680 (N_680,In_283,In_791);
nand U681 (N_681,In_723,In_1474);
nand U682 (N_682,In_1442,In_219);
and U683 (N_683,In_1377,In_1049);
xor U684 (N_684,In_1033,In_1114);
and U685 (N_685,In_559,In_1057);
xor U686 (N_686,In_979,In_1125);
or U687 (N_687,In_134,In_1199);
and U688 (N_688,In_903,In_176);
nand U689 (N_689,In_98,In_782);
or U690 (N_690,In_1150,In_274);
nor U691 (N_691,In_972,In_444);
and U692 (N_692,In_920,In_1388);
nor U693 (N_693,In_1272,In_1342);
and U694 (N_694,In_410,In_509);
and U695 (N_695,In_916,In_575);
nand U696 (N_696,In_1141,In_1127);
nor U697 (N_697,In_202,In_500);
and U698 (N_698,In_862,In_651);
nor U699 (N_699,In_904,In_1429);
nor U700 (N_700,In_236,In_931);
nand U701 (N_701,In_1346,In_1101);
and U702 (N_702,In_953,In_893);
nand U703 (N_703,In_1337,In_543);
or U704 (N_704,In_1011,In_613);
nand U705 (N_705,In_761,In_447);
nand U706 (N_706,In_540,In_775);
or U707 (N_707,In_185,In_141);
nor U708 (N_708,In_54,In_1108);
nand U709 (N_709,In_124,In_1102);
nor U710 (N_710,In_756,In_151);
or U711 (N_711,In_1113,In_940);
and U712 (N_712,In_766,In_481);
nor U713 (N_713,In_716,In_483);
or U714 (N_714,In_256,In_1348);
or U715 (N_715,In_629,In_1020);
nor U716 (N_716,In_981,In_754);
and U717 (N_717,In_91,In_14);
nor U718 (N_718,In_563,In_1223);
and U719 (N_719,In_40,In_529);
and U720 (N_720,In_390,In_1416);
nand U721 (N_721,In_1384,In_804);
xor U722 (N_722,In_1277,In_129);
nand U723 (N_723,In_110,In_1347);
xnor U724 (N_724,In_814,In_455);
nand U725 (N_725,In_302,In_281);
nand U726 (N_726,In_1024,In_1366);
nor U727 (N_727,In_1260,In_828);
or U728 (N_728,In_967,In_702);
nand U729 (N_729,In_325,In_757);
nor U730 (N_730,In_77,In_787);
or U731 (N_731,In_33,In_384);
and U732 (N_732,In_1359,In_805);
nor U733 (N_733,In_1105,In_897);
nand U734 (N_734,In_1179,In_881);
xnor U735 (N_735,In_1486,In_790);
and U736 (N_736,In_178,In_751);
nor U737 (N_737,In_1023,In_1228);
nand U738 (N_738,In_585,In_1222);
or U739 (N_739,In_1190,In_672);
and U740 (N_740,In_913,In_128);
nor U741 (N_741,In_1184,In_338);
and U742 (N_742,In_1218,In_52);
nand U743 (N_743,In_780,In_80);
and U744 (N_744,In_1411,In_1386);
nand U745 (N_745,In_717,In_778);
or U746 (N_746,In_472,In_1242);
xor U747 (N_747,In_1498,In_774);
nand U748 (N_748,In_11,In_1010);
nor U749 (N_749,In_777,In_84);
xor U750 (N_750,N_455,N_209);
nand U751 (N_751,N_190,N_676);
nor U752 (N_752,N_31,N_735);
xor U753 (N_753,N_687,N_596);
nand U754 (N_754,N_436,N_524);
nand U755 (N_755,N_278,N_42);
nand U756 (N_756,N_590,N_139);
nor U757 (N_757,N_199,N_639);
and U758 (N_758,N_301,N_247);
nor U759 (N_759,N_371,N_619);
or U760 (N_760,N_38,N_552);
and U761 (N_761,N_239,N_588);
xnor U762 (N_762,N_515,N_352);
xnor U763 (N_763,N_447,N_529);
or U764 (N_764,N_587,N_165);
xor U765 (N_765,N_81,N_12);
and U766 (N_766,N_29,N_547);
nor U767 (N_767,N_305,N_143);
nor U768 (N_768,N_633,N_68);
xor U769 (N_769,N_109,N_140);
or U770 (N_770,N_567,N_579);
xor U771 (N_771,N_655,N_441);
and U772 (N_772,N_742,N_240);
nor U773 (N_773,N_335,N_237);
nand U774 (N_774,N_336,N_218);
nor U775 (N_775,N_673,N_54);
and U776 (N_776,N_453,N_150);
nor U777 (N_777,N_37,N_323);
or U778 (N_778,N_671,N_456);
nand U779 (N_779,N_137,N_520);
nor U780 (N_780,N_193,N_610);
and U781 (N_781,N_608,N_219);
and U782 (N_782,N_228,N_9);
and U783 (N_783,N_325,N_389);
nor U784 (N_784,N_294,N_440);
nand U785 (N_785,N_292,N_248);
nor U786 (N_786,N_347,N_424);
nand U787 (N_787,N_250,N_331);
or U788 (N_788,N_729,N_24);
or U789 (N_789,N_463,N_562);
nor U790 (N_790,N_11,N_327);
or U791 (N_791,N_4,N_312);
or U792 (N_792,N_122,N_614);
nand U793 (N_793,N_123,N_138);
nor U794 (N_794,N_76,N_216);
nand U795 (N_795,N_181,N_206);
and U796 (N_796,N_211,N_465);
nand U797 (N_797,N_377,N_259);
nand U798 (N_798,N_513,N_592);
nand U799 (N_799,N_189,N_556);
and U800 (N_800,N_399,N_207);
or U801 (N_801,N_304,N_19);
nor U802 (N_802,N_665,N_580);
or U803 (N_803,N_656,N_415);
or U804 (N_804,N_50,N_48);
and U805 (N_805,N_249,N_420);
nor U806 (N_806,N_669,N_115);
xnor U807 (N_807,N_285,N_23);
or U808 (N_808,N_417,N_727);
nor U809 (N_809,N_126,N_692);
and U810 (N_810,N_565,N_238);
nand U811 (N_811,N_690,N_706);
or U812 (N_812,N_98,N_721);
and U813 (N_813,N_210,N_689);
nor U814 (N_814,N_177,N_409);
nor U815 (N_815,N_51,N_30);
xnor U816 (N_816,N_523,N_183);
nor U817 (N_817,N_668,N_509);
nor U818 (N_818,N_41,N_376);
xnor U819 (N_819,N_2,N_403);
nand U820 (N_820,N_146,N_675);
and U821 (N_821,N_49,N_253);
or U822 (N_822,N_0,N_222);
and U823 (N_823,N_220,N_315);
and U824 (N_824,N_40,N_468);
nor U825 (N_825,N_493,N_470);
or U826 (N_826,N_229,N_539);
nor U827 (N_827,N_343,N_713);
nand U828 (N_828,N_320,N_395);
or U829 (N_829,N_308,N_73);
or U830 (N_830,N_421,N_540);
or U831 (N_831,N_723,N_637);
nor U832 (N_832,N_145,N_271);
or U833 (N_833,N_235,N_442);
nand U834 (N_834,N_407,N_615);
and U835 (N_835,N_510,N_95);
or U836 (N_836,N_164,N_197);
and U837 (N_837,N_194,N_460);
nor U838 (N_838,N_495,N_629);
nor U839 (N_839,N_367,N_152);
nand U840 (N_840,N_712,N_15);
or U841 (N_841,N_67,N_517);
nand U842 (N_842,N_429,N_476);
nand U843 (N_843,N_494,N_408);
nand U844 (N_844,N_302,N_501);
xnor U845 (N_845,N_276,N_256);
nand U846 (N_846,N_745,N_534);
or U847 (N_847,N_353,N_375);
or U848 (N_848,N_281,N_416);
nor U849 (N_849,N_473,N_471);
and U850 (N_850,N_431,N_560);
or U851 (N_851,N_680,N_79);
nor U852 (N_852,N_22,N_354);
nor U853 (N_853,N_201,N_260);
nand U854 (N_854,N_649,N_575);
and U855 (N_855,N_449,N_322);
nor U856 (N_856,N_487,N_66);
nor U857 (N_857,N_356,N_666);
and U858 (N_858,N_132,N_659);
nand U859 (N_859,N_536,N_173);
xnor U860 (N_860,N_572,N_443);
and U861 (N_861,N_551,N_196);
nor U862 (N_862,N_664,N_382);
or U863 (N_863,N_662,N_591);
or U864 (N_864,N_484,N_191);
and U865 (N_865,N_188,N_215);
or U866 (N_866,N_135,N_341);
and U867 (N_867,N_586,N_383);
nand U868 (N_868,N_459,N_722);
or U869 (N_869,N_412,N_338);
nor U870 (N_870,N_573,N_184);
nor U871 (N_871,N_225,N_477);
or U872 (N_872,N_158,N_446);
nor U873 (N_873,N_332,N_681);
nand U874 (N_874,N_101,N_326);
or U875 (N_875,N_154,N_434);
or U876 (N_876,N_363,N_593);
or U877 (N_877,N_339,N_148);
and U878 (N_878,N_433,N_77);
or U879 (N_879,N_702,N_557);
xor U880 (N_880,N_740,N_728);
or U881 (N_881,N_521,N_627);
nand U882 (N_882,N_651,N_679);
and U883 (N_883,N_75,N_232);
or U884 (N_884,N_461,N_21);
xor U885 (N_885,N_92,N_396);
or U886 (N_886,N_703,N_500);
and U887 (N_887,N_130,N_504);
and U888 (N_888,N_94,N_732);
or U889 (N_889,N_648,N_97);
or U890 (N_890,N_364,N_561);
xor U891 (N_891,N_231,N_718);
nand U892 (N_892,N_233,N_373);
or U893 (N_893,N_111,N_317);
nand U894 (N_894,N_46,N_506);
and U895 (N_895,N_749,N_26);
nor U896 (N_896,N_464,N_604);
nand U897 (N_897,N_310,N_124);
and U898 (N_898,N_444,N_620);
nand U899 (N_899,N_609,N_632);
nand U900 (N_900,N_330,N_58);
nand U901 (N_901,N_518,N_612);
nor U902 (N_902,N_195,N_716);
and U903 (N_903,N_685,N_474);
xor U904 (N_904,N_273,N_693);
nor U905 (N_905,N_170,N_660);
or U906 (N_906,N_284,N_594);
nor U907 (N_907,N_631,N_527);
nand U908 (N_908,N_204,N_102);
nand U909 (N_909,N_63,N_372);
and U910 (N_910,N_569,N_85);
or U911 (N_911,N_475,N_566);
nor U912 (N_912,N_623,N_306);
nor U913 (N_913,N_34,N_617);
nor U914 (N_914,N_160,N_142);
or U915 (N_915,N_652,N_125);
or U916 (N_916,N_741,N_485);
or U917 (N_917,N_466,N_646);
and U918 (N_918,N_87,N_576);
and U919 (N_919,N_704,N_243);
and U920 (N_920,N_411,N_202);
xor U921 (N_921,N_333,N_52);
and U922 (N_922,N_127,N_153);
and U923 (N_923,N_597,N_635);
nor U924 (N_924,N_653,N_172);
nor U925 (N_925,N_583,N_611);
and U926 (N_926,N_496,N_695);
and U927 (N_927,N_70,N_599);
nor U928 (N_928,N_585,N_488);
and U929 (N_929,N_167,N_404);
or U930 (N_930,N_528,N_746);
and U931 (N_931,N_283,N_272);
or U932 (N_932,N_563,N_743);
nand U933 (N_933,N_598,N_93);
nor U934 (N_934,N_548,N_44);
nand U935 (N_935,N_486,N_711);
nor U936 (N_936,N_166,N_602);
or U937 (N_937,N_425,N_589);
nand U938 (N_938,N_267,N_214);
or U939 (N_939,N_419,N_708);
nand U940 (N_940,N_119,N_187);
nor U941 (N_941,N_393,N_112);
nor U942 (N_942,N_630,N_28);
nor U943 (N_943,N_246,N_90);
nor U944 (N_944,N_72,N_236);
nor U945 (N_945,N_295,N_169);
nor U946 (N_946,N_251,N_437);
nand U947 (N_947,N_739,N_147);
and U948 (N_948,N_277,N_185);
nor U949 (N_949,N_600,N_120);
nand U950 (N_950,N_55,N_697);
nand U951 (N_951,N_568,N_525);
or U952 (N_952,N_387,N_141);
and U953 (N_953,N_349,N_672);
or U954 (N_954,N_423,N_227);
nor U955 (N_955,N_293,N_663);
nor U956 (N_956,N_252,N_480);
and U957 (N_957,N_638,N_144);
nand U958 (N_958,N_108,N_719);
and U959 (N_959,N_360,N_526);
xor U960 (N_960,N_674,N_359);
and U961 (N_961,N_554,N_3);
or U962 (N_962,N_625,N_178);
or U963 (N_963,N_469,N_406);
or U964 (N_964,N_133,N_606);
nor U965 (N_965,N_698,N_490);
nor U966 (N_966,N_641,N_291);
nor U967 (N_967,N_726,N_577);
nor U968 (N_968,N_351,N_657);
nand U969 (N_969,N_581,N_368);
nor U970 (N_970,N_747,N_691);
and U971 (N_971,N_186,N_157);
or U972 (N_972,N_532,N_479);
or U973 (N_973,N_56,N_282);
nand U974 (N_974,N_381,N_400);
or U975 (N_975,N_329,N_457);
and U976 (N_976,N_16,N_128);
nor U977 (N_977,N_321,N_365);
nand U978 (N_978,N_162,N_438);
xnor U979 (N_979,N_208,N_319);
or U980 (N_980,N_519,N_234);
or U981 (N_981,N_618,N_388);
or U982 (N_982,N_314,N_47);
nand U983 (N_983,N_155,N_448);
nor U984 (N_984,N_405,N_550);
xor U985 (N_985,N_654,N_161);
or U986 (N_986,N_245,N_45);
nand U987 (N_987,N_450,N_350);
nand U988 (N_988,N_340,N_710);
nand U989 (N_989,N_462,N_748);
and U990 (N_990,N_516,N_91);
and U991 (N_991,N_458,N_221);
and U992 (N_992,N_394,N_263);
nand U993 (N_993,N_334,N_574);
nand U994 (N_994,N_118,N_616);
and U995 (N_995,N_492,N_553);
or U996 (N_996,N_570,N_1);
nand U997 (N_997,N_182,N_131);
nand U998 (N_998,N_83,N_299);
nand U999 (N_999,N_451,N_99);
or U1000 (N_1000,N_715,N_626);
or U1001 (N_1001,N_640,N_503);
and U1002 (N_1002,N_18,N_43);
or U1003 (N_1003,N_483,N_595);
xnor U1004 (N_1004,N_621,N_582);
or U1005 (N_1005,N_736,N_694);
nor U1006 (N_1006,N_255,N_397);
and U1007 (N_1007,N_427,N_426);
xor U1008 (N_1008,N_514,N_543);
xnor U1009 (N_1009,N_176,N_264);
nand U1010 (N_1010,N_174,N_380);
and U1011 (N_1011,N_482,N_262);
and U1012 (N_1012,N_542,N_117);
or U1013 (N_1013,N_603,N_200);
or U1014 (N_1014,N_113,N_318);
and U1015 (N_1015,N_683,N_307);
nor U1016 (N_1016,N_505,N_61);
xor U1017 (N_1017,N_499,N_688);
or U1018 (N_1018,N_677,N_20);
or U1019 (N_1019,N_607,N_390);
or U1020 (N_1020,N_96,N_605);
nand U1021 (N_1021,N_701,N_696);
nand U1022 (N_1022,N_257,N_82);
or U1023 (N_1023,N_362,N_535);
or U1024 (N_1024,N_478,N_14);
nor U1025 (N_1025,N_428,N_13);
nand U1026 (N_1026,N_644,N_422);
nor U1027 (N_1027,N_386,N_544);
and U1028 (N_1028,N_129,N_366);
nand U1029 (N_1029,N_645,N_402);
nor U1030 (N_1030,N_296,N_149);
or U1031 (N_1031,N_667,N_337);
nor U1032 (N_1032,N_498,N_370);
or U1033 (N_1033,N_601,N_261);
nor U1034 (N_1034,N_686,N_324);
nand U1035 (N_1035,N_268,N_511);
or U1036 (N_1036,N_104,N_432);
or U1037 (N_1037,N_89,N_717);
nand U1038 (N_1038,N_643,N_10);
nor U1039 (N_1039,N_65,N_53);
nor U1040 (N_1040,N_297,N_59);
and U1041 (N_1041,N_467,N_5);
or U1042 (N_1042,N_439,N_744);
and U1043 (N_1043,N_401,N_33);
nand U1044 (N_1044,N_378,N_700);
and U1045 (N_1045,N_699,N_720);
nand U1046 (N_1046,N_559,N_642);
and U1047 (N_1047,N_290,N_175);
and U1048 (N_1048,N_622,N_670);
or U1049 (N_1049,N_287,N_555);
xnor U1050 (N_1050,N_578,N_110);
xnor U1051 (N_1051,N_628,N_289);
or U1052 (N_1052,N_39,N_242);
nor U1053 (N_1053,N_163,N_179);
nand U1054 (N_1054,N_545,N_538);
xor U1055 (N_1055,N_647,N_27);
and U1056 (N_1056,N_274,N_57);
xor U1057 (N_1057,N_385,N_430);
and U1058 (N_1058,N_714,N_658);
xnor U1059 (N_1059,N_316,N_270);
or U1060 (N_1060,N_300,N_584);
or U1061 (N_1061,N_180,N_205);
or U1062 (N_1062,N_71,N_391);
or U1063 (N_1063,N_286,N_313);
xor U1064 (N_1064,N_100,N_379);
nand U1065 (N_1065,N_730,N_151);
nand U1066 (N_1066,N_684,N_384);
or U1067 (N_1067,N_32,N_192);
and U1068 (N_1068,N_392,N_558);
or U1069 (N_1069,N_705,N_344);
or U1070 (N_1070,N_346,N_311);
nand U1071 (N_1071,N_624,N_650);
and U1072 (N_1072,N_288,N_682);
xnor U1073 (N_1073,N_266,N_636);
or U1074 (N_1074,N_106,N_709);
nor U1075 (N_1075,N_733,N_345);
xnor U1076 (N_1076,N_134,N_541);
and U1077 (N_1077,N_107,N_435);
or U1078 (N_1078,N_445,N_724);
or U1079 (N_1079,N_481,N_512);
nor U1080 (N_1080,N_203,N_280);
nor U1081 (N_1081,N_223,N_734);
xnor U1082 (N_1082,N_410,N_533);
nor U1083 (N_1083,N_452,N_303);
nand U1084 (N_1084,N_114,N_212);
and U1085 (N_1085,N_678,N_328);
or U1086 (N_1086,N_244,N_171);
or U1087 (N_1087,N_342,N_298);
nor U1088 (N_1088,N_348,N_230);
and U1089 (N_1089,N_265,N_136);
or U1090 (N_1090,N_309,N_198);
and U1091 (N_1091,N_355,N_224);
or U1092 (N_1092,N_74,N_8);
xnor U1093 (N_1093,N_103,N_613);
nor U1094 (N_1094,N_357,N_737);
nand U1095 (N_1095,N_549,N_418);
nor U1096 (N_1096,N_241,N_86);
or U1097 (N_1097,N_6,N_275);
nand U1098 (N_1098,N_537,N_269);
nor U1099 (N_1099,N_80,N_661);
and U1100 (N_1100,N_35,N_62);
or U1101 (N_1101,N_507,N_60);
nand U1102 (N_1102,N_36,N_358);
xor U1103 (N_1103,N_454,N_88);
nand U1104 (N_1104,N_508,N_374);
and U1105 (N_1105,N_226,N_105);
nand U1106 (N_1106,N_254,N_522);
and U1107 (N_1107,N_546,N_502);
nand U1108 (N_1108,N_213,N_564);
nand U1109 (N_1109,N_159,N_84);
and U1110 (N_1110,N_414,N_489);
nor U1111 (N_1111,N_17,N_279);
nor U1112 (N_1112,N_258,N_531);
and U1113 (N_1113,N_69,N_707);
or U1114 (N_1114,N_78,N_530);
nor U1115 (N_1115,N_571,N_491);
xor U1116 (N_1116,N_64,N_217);
and U1117 (N_1117,N_725,N_413);
and U1118 (N_1118,N_634,N_472);
and U1119 (N_1119,N_121,N_7);
or U1120 (N_1120,N_25,N_497);
xnor U1121 (N_1121,N_398,N_116);
and U1122 (N_1122,N_731,N_168);
and U1123 (N_1123,N_738,N_156);
and U1124 (N_1124,N_361,N_369);
nand U1125 (N_1125,N_229,N_472);
or U1126 (N_1126,N_120,N_620);
and U1127 (N_1127,N_667,N_699);
and U1128 (N_1128,N_603,N_356);
nor U1129 (N_1129,N_441,N_65);
xnor U1130 (N_1130,N_25,N_84);
nor U1131 (N_1131,N_305,N_169);
nor U1132 (N_1132,N_103,N_96);
nor U1133 (N_1133,N_244,N_489);
nand U1134 (N_1134,N_358,N_592);
and U1135 (N_1135,N_441,N_20);
and U1136 (N_1136,N_176,N_491);
or U1137 (N_1137,N_381,N_156);
nor U1138 (N_1138,N_661,N_387);
nand U1139 (N_1139,N_516,N_67);
nand U1140 (N_1140,N_616,N_683);
nor U1141 (N_1141,N_104,N_71);
or U1142 (N_1142,N_194,N_662);
nand U1143 (N_1143,N_530,N_135);
nor U1144 (N_1144,N_377,N_111);
or U1145 (N_1145,N_277,N_455);
nor U1146 (N_1146,N_373,N_191);
or U1147 (N_1147,N_348,N_162);
nand U1148 (N_1148,N_549,N_51);
nor U1149 (N_1149,N_54,N_518);
nand U1150 (N_1150,N_651,N_9);
or U1151 (N_1151,N_589,N_678);
nand U1152 (N_1152,N_576,N_682);
nand U1153 (N_1153,N_279,N_348);
nand U1154 (N_1154,N_481,N_52);
or U1155 (N_1155,N_699,N_500);
nor U1156 (N_1156,N_321,N_251);
or U1157 (N_1157,N_153,N_464);
or U1158 (N_1158,N_10,N_280);
nand U1159 (N_1159,N_81,N_503);
nor U1160 (N_1160,N_114,N_475);
nand U1161 (N_1161,N_91,N_597);
nand U1162 (N_1162,N_744,N_448);
and U1163 (N_1163,N_283,N_726);
or U1164 (N_1164,N_53,N_301);
and U1165 (N_1165,N_498,N_301);
and U1166 (N_1166,N_663,N_484);
xnor U1167 (N_1167,N_582,N_214);
and U1168 (N_1168,N_711,N_550);
and U1169 (N_1169,N_99,N_229);
or U1170 (N_1170,N_206,N_667);
xor U1171 (N_1171,N_262,N_749);
nor U1172 (N_1172,N_275,N_23);
xnor U1173 (N_1173,N_86,N_495);
nor U1174 (N_1174,N_120,N_36);
xnor U1175 (N_1175,N_415,N_234);
or U1176 (N_1176,N_290,N_600);
and U1177 (N_1177,N_261,N_59);
nand U1178 (N_1178,N_219,N_96);
and U1179 (N_1179,N_327,N_273);
and U1180 (N_1180,N_630,N_451);
and U1181 (N_1181,N_510,N_535);
and U1182 (N_1182,N_582,N_546);
nand U1183 (N_1183,N_346,N_481);
or U1184 (N_1184,N_116,N_290);
nor U1185 (N_1185,N_464,N_539);
nand U1186 (N_1186,N_283,N_494);
and U1187 (N_1187,N_114,N_178);
xor U1188 (N_1188,N_175,N_99);
or U1189 (N_1189,N_748,N_335);
nand U1190 (N_1190,N_370,N_80);
nor U1191 (N_1191,N_64,N_446);
nor U1192 (N_1192,N_195,N_230);
nor U1193 (N_1193,N_320,N_149);
or U1194 (N_1194,N_308,N_740);
nand U1195 (N_1195,N_418,N_741);
xor U1196 (N_1196,N_469,N_399);
and U1197 (N_1197,N_107,N_87);
nand U1198 (N_1198,N_500,N_380);
nor U1199 (N_1199,N_298,N_196);
nor U1200 (N_1200,N_327,N_132);
nand U1201 (N_1201,N_729,N_672);
nor U1202 (N_1202,N_212,N_125);
or U1203 (N_1203,N_742,N_142);
or U1204 (N_1204,N_526,N_97);
nor U1205 (N_1205,N_637,N_106);
nor U1206 (N_1206,N_230,N_666);
nand U1207 (N_1207,N_265,N_57);
nor U1208 (N_1208,N_509,N_482);
nand U1209 (N_1209,N_541,N_598);
and U1210 (N_1210,N_249,N_98);
xor U1211 (N_1211,N_255,N_458);
xnor U1212 (N_1212,N_403,N_504);
nand U1213 (N_1213,N_356,N_345);
and U1214 (N_1214,N_686,N_37);
and U1215 (N_1215,N_216,N_336);
and U1216 (N_1216,N_335,N_279);
nand U1217 (N_1217,N_216,N_615);
or U1218 (N_1218,N_537,N_323);
or U1219 (N_1219,N_659,N_588);
nand U1220 (N_1220,N_153,N_391);
and U1221 (N_1221,N_607,N_36);
nand U1222 (N_1222,N_467,N_67);
or U1223 (N_1223,N_307,N_608);
and U1224 (N_1224,N_150,N_531);
and U1225 (N_1225,N_110,N_676);
nor U1226 (N_1226,N_563,N_273);
nand U1227 (N_1227,N_706,N_350);
xnor U1228 (N_1228,N_649,N_119);
nor U1229 (N_1229,N_113,N_541);
nand U1230 (N_1230,N_135,N_126);
and U1231 (N_1231,N_19,N_333);
or U1232 (N_1232,N_727,N_247);
nand U1233 (N_1233,N_22,N_389);
or U1234 (N_1234,N_699,N_302);
and U1235 (N_1235,N_308,N_235);
and U1236 (N_1236,N_739,N_72);
or U1237 (N_1237,N_104,N_450);
and U1238 (N_1238,N_118,N_661);
nand U1239 (N_1239,N_706,N_82);
nor U1240 (N_1240,N_542,N_535);
or U1241 (N_1241,N_647,N_208);
nor U1242 (N_1242,N_317,N_267);
nor U1243 (N_1243,N_102,N_313);
and U1244 (N_1244,N_635,N_722);
nand U1245 (N_1245,N_10,N_441);
and U1246 (N_1246,N_507,N_615);
xnor U1247 (N_1247,N_624,N_362);
nand U1248 (N_1248,N_745,N_293);
nand U1249 (N_1249,N_88,N_318);
nor U1250 (N_1250,N_654,N_84);
nor U1251 (N_1251,N_121,N_354);
or U1252 (N_1252,N_426,N_738);
and U1253 (N_1253,N_692,N_231);
nor U1254 (N_1254,N_694,N_3);
and U1255 (N_1255,N_321,N_183);
nand U1256 (N_1256,N_675,N_344);
nor U1257 (N_1257,N_227,N_357);
or U1258 (N_1258,N_107,N_48);
nand U1259 (N_1259,N_732,N_242);
nor U1260 (N_1260,N_265,N_224);
nand U1261 (N_1261,N_311,N_260);
and U1262 (N_1262,N_531,N_647);
nand U1263 (N_1263,N_294,N_166);
nor U1264 (N_1264,N_510,N_698);
xor U1265 (N_1265,N_377,N_667);
and U1266 (N_1266,N_281,N_210);
nand U1267 (N_1267,N_591,N_451);
and U1268 (N_1268,N_326,N_501);
nand U1269 (N_1269,N_107,N_257);
nand U1270 (N_1270,N_423,N_218);
xnor U1271 (N_1271,N_136,N_370);
and U1272 (N_1272,N_590,N_436);
or U1273 (N_1273,N_530,N_144);
xnor U1274 (N_1274,N_324,N_293);
or U1275 (N_1275,N_134,N_743);
nor U1276 (N_1276,N_278,N_459);
and U1277 (N_1277,N_271,N_721);
and U1278 (N_1278,N_279,N_19);
nor U1279 (N_1279,N_232,N_242);
or U1280 (N_1280,N_460,N_520);
and U1281 (N_1281,N_363,N_313);
or U1282 (N_1282,N_279,N_360);
nand U1283 (N_1283,N_367,N_518);
nor U1284 (N_1284,N_142,N_461);
and U1285 (N_1285,N_658,N_483);
nand U1286 (N_1286,N_637,N_595);
nor U1287 (N_1287,N_336,N_275);
and U1288 (N_1288,N_245,N_177);
or U1289 (N_1289,N_366,N_522);
nor U1290 (N_1290,N_433,N_195);
nand U1291 (N_1291,N_554,N_463);
nand U1292 (N_1292,N_605,N_603);
nor U1293 (N_1293,N_711,N_251);
nand U1294 (N_1294,N_319,N_478);
and U1295 (N_1295,N_427,N_113);
nand U1296 (N_1296,N_444,N_141);
and U1297 (N_1297,N_46,N_447);
and U1298 (N_1298,N_738,N_191);
nand U1299 (N_1299,N_280,N_288);
or U1300 (N_1300,N_312,N_59);
or U1301 (N_1301,N_583,N_266);
xnor U1302 (N_1302,N_460,N_357);
and U1303 (N_1303,N_270,N_648);
or U1304 (N_1304,N_591,N_157);
nor U1305 (N_1305,N_651,N_258);
nand U1306 (N_1306,N_157,N_435);
and U1307 (N_1307,N_121,N_695);
nand U1308 (N_1308,N_109,N_160);
nor U1309 (N_1309,N_488,N_45);
or U1310 (N_1310,N_740,N_136);
and U1311 (N_1311,N_685,N_289);
and U1312 (N_1312,N_549,N_568);
or U1313 (N_1313,N_124,N_117);
nand U1314 (N_1314,N_285,N_530);
and U1315 (N_1315,N_8,N_500);
nor U1316 (N_1316,N_686,N_164);
and U1317 (N_1317,N_650,N_588);
or U1318 (N_1318,N_493,N_255);
or U1319 (N_1319,N_511,N_456);
nand U1320 (N_1320,N_111,N_577);
nand U1321 (N_1321,N_599,N_390);
nor U1322 (N_1322,N_720,N_97);
nor U1323 (N_1323,N_695,N_593);
nand U1324 (N_1324,N_84,N_142);
nor U1325 (N_1325,N_467,N_99);
or U1326 (N_1326,N_163,N_129);
or U1327 (N_1327,N_228,N_534);
and U1328 (N_1328,N_553,N_251);
and U1329 (N_1329,N_165,N_337);
nor U1330 (N_1330,N_697,N_132);
and U1331 (N_1331,N_509,N_242);
nand U1332 (N_1332,N_130,N_326);
nor U1333 (N_1333,N_138,N_487);
or U1334 (N_1334,N_332,N_496);
and U1335 (N_1335,N_520,N_719);
and U1336 (N_1336,N_294,N_300);
nor U1337 (N_1337,N_373,N_416);
or U1338 (N_1338,N_477,N_219);
nand U1339 (N_1339,N_666,N_677);
or U1340 (N_1340,N_652,N_698);
nor U1341 (N_1341,N_525,N_201);
nor U1342 (N_1342,N_167,N_35);
or U1343 (N_1343,N_150,N_733);
nor U1344 (N_1344,N_335,N_134);
and U1345 (N_1345,N_445,N_636);
nor U1346 (N_1346,N_89,N_512);
or U1347 (N_1347,N_558,N_191);
and U1348 (N_1348,N_225,N_52);
nor U1349 (N_1349,N_436,N_170);
or U1350 (N_1350,N_82,N_396);
and U1351 (N_1351,N_358,N_238);
xor U1352 (N_1352,N_356,N_708);
nand U1353 (N_1353,N_251,N_44);
and U1354 (N_1354,N_387,N_92);
nor U1355 (N_1355,N_256,N_412);
nand U1356 (N_1356,N_643,N_168);
nor U1357 (N_1357,N_457,N_429);
nand U1358 (N_1358,N_397,N_714);
nor U1359 (N_1359,N_10,N_548);
or U1360 (N_1360,N_705,N_369);
nor U1361 (N_1361,N_143,N_471);
or U1362 (N_1362,N_287,N_451);
nor U1363 (N_1363,N_29,N_41);
nand U1364 (N_1364,N_513,N_402);
or U1365 (N_1365,N_360,N_534);
and U1366 (N_1366,N_259,N_406);
or U1367 (N_1367,N_256,N_170);
nor U1368 (N_1368,N_387,N_134);
nand U1369 (N_1369,N_412,N_113);
or U1370 (N_1370,N_648,N_222);
nor U1371 (N_1371,N_105,N_113);
and U1372 (N_1372,N_22,N_408);
or U1373 (N_1373,N_28,N_256);
or U1374 (N_1374,N_274,N_353);
and U1375 (N_1375,N_565,N_141);
nor U1376 (N_1376,N_38,N_669);
nand U1377 (N_1377,N_524,N_452);
nand U1378 (N_1378,N_649,N_347);
and U1379 (N_1379,N_186,N_711);
xnor U1380 (N_1380,N_494,N_691);
nor U1381 (N_1381,N_592,N_217);
xor U1382 (N_1382,N_211,N_349);
or U1383 (N_1383,N_511,N_17);
or U1384 (N_1384,N_676,N_146);
nor U1385 (N_1385,N_491,N_95);
nor U1386 (N_1386,N_438,N_731);
nor U1387 (N_1387,N_25,N_631);
nand U1388 (N_1388,N_228,N_78);
and U1389 (N_1389,N_92,N_507);
or U1390 (N_1390,N_303,N_523);
nand U1391 (N_1391,N_117,N_196);
xnor U1392 (N_1392,N_664,N_100);
and U1393 (N_1393,N_626,N_31);
or U1394 (N_1394,N_46,N_645);
nor U1395 (N_1395,N_341,N_240);
and U1396 (N_1396,N_369,N_398);
and U1397 (N_1397,N_533,N_462);
xnor U1398 (N_1398,N_269,N_246);
nor U1399 (N_1399,N_732,N_436);
xor U1400 (N_1400,N_150,N_475);
xor U1401 (N_1401,N_104,N_110);
and U1402 (N_1402,N_415,N_576);
nand U1403 (N_1403,N_221,N_464);
or U1404 (N_1404,N_472,N_594);
nor U1405 (N_1405,N_477,N_497);
and U1406 (N_1406,N_361,N_427);
nand U1407 (N_1407,N_580,N_685);
and U1408 (N_1408,N_103,N_177);
nor U1409 (N_1409,N_588,N_556);
and U1410 (N_1410,N_546,N_728);
and U1411 (N_1411,N_667,N_124);
or U1412 (N_1412,N_307,N_494);
nand U1413 (N_1413,N_33,N_171);
or U1414 (N_1414,N_459,N_251);
or U1415 (N_1415,N_51,N_489);
and U1416 (N_1416,N_707,N_314);
nand U1417 (N_1417,N_477,N_464);
and U1418 (N_1418,N_746,N_728);
nor U1419 (N_1419,N_717,N_217);
or U1420 (N_1420,N_216,N_129);
nand U1421 (N_1421,N_653,N_316);
or U1422 (N_1422,N_672,N_185);
nor U1423 (N_1423,N_284,N_230);
xor U1424 (N_1424,N_188,N_641);
nand U1425 (N_1425,N_96,N_144);
and U1426 (N_1426,N_156,N_44);
and U1427 (N_1427,N_359,N_522);
nor U1428 (N_1428,N_533,N_632);
and U1429 (N_1429,N_130,N_594);
nand U1430 (N_1430,N_710,N_405);
nand U1431 (N_1431,N_303,N_24);
xnor U1432 (N_1432,N_710,N_539);
or U1433 (N_1433,N_460,N_344);
or U1434 (N_1434,N_88,N_577);
and U1435 (N_1435,N_737,N_10);
or U1436 (N_1436,N_445,N_401);
and U1437 (N_1437,N_653,N_640);
nand U1438 (N_1438,N_252,N_318);
nor U1439 (N_1439,N_281,N_207);
nand U1440 (N_1440,N_604,N_516);
or U1441 (N_1441,N_324,N_653);
nor U1442 (N_1442,N_457,N_520);
and U1443 (N_1443,N_459,N_144);
nand U1444 (N_1444,N_478,N_380);
nand U1445 (N_1445,N_204,N_433);
or U1446 (N_1446,N_292,N_706);
and U1447 (N_1447,N_485,N_576);
or U1448 (N_1448,N_44,N_694);
nor U1449 (N_1449,N_566,N_628);
and U1450 (N_1450,N_321,N_11);
nor U1451 (N_1451,N_74,N_676);
and U1452 (N_1452,N_604,N_127);
and U1453 (N_1453,N_250,N_204);
and U1454 (N_1454,N_40,N_511);
nand U1455 (N_1455,N_86,N_355);
or U1456 (N_1456,N_119,N_525);
xor U1457 (N_1457,N_533,N_377);
or U1458 (N_1458,N_510,N_129);
or U1459 (N_1459,N_210,N_266);
nand U1460 (N_1460,N_362,N_106);
or U1461 (N_1461,N_108,N_82);
or U1462 (N_1462,N_465,N_392);
nand U1463 (N_1463,N_57,N_706);
xnor U1464 (N_1464,N_621,N_78);
or U1465 (N_1465,N_57,N_302);
xnor U1466 (N_1466,N_251,N_538);
and U1467 (N_1467,N_96,N_266);
or U1468 (N_1468,N_58,N_79);
nor U1469 (N_1469,N_259,N_506);
or U1470 (N_1470,N_706,N_36);
xnor U1471 (N_1471,N_361,N_211);
and U1472 (N_1472,N_441,N_334);
xnor U1473 (N_1473,N_591,N_705);
or U1474 (N_1474,N_242,N_409);
nand U1475 (N_1475,N_639,N_202);
nor U1476 (N_1476,N_3,N_238);
and U1477 (N_1477,N_578,N_547);
nor U1478 (N_1478,N_2,N_396);
and U1479 (N_1479,N_40,N_576);
nor U1480 (N_1480,N_315,N_706);
and U1481 (N_1481,N_618,N_665);
or U1482 (N_1482,N_497,N_298);
or U1483 (N_1483,N_335,N_506);
or U1484 (N_1484,N_589,N_176);
and U1485 (N_1485,N_390,N_179);
xnor U1486 (N_1486,N_224,N_472);
and U1487 (N_1487,N_17,N_419);
nor U1488 (N_1488,N_654,N_353);
or U1489 (N_1489,N_415,N_388);
nor U1490 (N_1490,N_249,N_314);
or U1491 (N_1491,N_367,N_571);
nor U1492 (N_1492,N_623,N_555);
nor U1493 (N_1493,N_165,N_443);
nand U1494 (N_1494,N_436,N_422);
nand U1495 (N_1495,N_491,N_527);
nand U1496 (N_1496,N_494,N_17);
or U1497 (N_1497,N_260,N_108);
or U1498 (N_1498,N_272,N_288);
nor U1499 (N_1499,N_716,N_710);
nor U1500 (N_1500,N_798,N_1112);
nor U1501 (N_1501,N_1261,N_1013);
xnor U1502 (N_1502,N_1285,N_913);
or U1503 (N_1503,N_1037,N_1273);
xor U1504 (N_1504,N_1330,N_957);
nor U1505 (N_1505,N_1304,N_1118);
nor U1506 (N_1506,N_1391,N_1068);
or U1507 (N_1507,N_1196,N_1006);
xor U1508 (N_1508,N_1237,N_859);
nand U1509 (N_1509,N_1349,N_1070);
xnor U1510 (N_1510,N_818,N_1086);
and U1511 (N_1511,N_1369,N_1227);
nor U1512 (N_1512,N_1046,N_1348);
nand U1513 (N_1513,N_899,N_922);
and U1514 (N_1514,N_1413,N_1200);
nand U1515 (N_1515,N_1274,N_858);
nor U1516 (N_1516,N_1033,N_948);
nand U1517 (N_1517,N_829,N_1322);
or U1518 (N_1518,N_1302,N_995);
xnor U1519 (N_1519,N_1448,N_1409);
and U1520 (N_1520,N_935,N_1400);
nor U1521 (N_1521,N_1250,N_941);
nor U1522 (N_1522,N_1028,N_891);
or U1523 (N_1523,N_938,N_838);
nand U1524 (N_1524,N_888,N_999);
nand U1525 (N_1525,N_826,N_783);
nor U1526 (N_1526,N_1219,N_915);
and U1527 (N_1527,N_889,N_1486);
and U1528 (N_1528,N_761,N_1236);
or U1529 (N_1529,N_1073,N_1388);
nand U1530 (N_1530,N_1299,N_994);
nand U1531 (N_1531,N_1089,N_1498);
nand U1532 (N_1532,N_764,N_1120);
xor U1533 (N_1533,N_765,N_1451);
nor U1534 (N_1534,N_1359,N_1380);
and U1535 (N_1535,N_1293,N_794);
or U1536 (N_1536,N_1238,N_1057);
or U1537 (N_1537,N_949,N_1318);
or U1538 (N_1538,N_1184,N_895);
nand U1539 (N_1539,N_1278,N_880);
nor U1540 (N_1540,N_919,N_979);
nor U1541 (N_1541,N_1376,N_1469);
or U1542 (N_1542,N_1263,N_1141);
or U1543 (N_1543,N_930,N_752);
xor U1544 (N_1544,N_1043,N_795);
nand U1545 (N_1545,N_1095,N_1496);
and U1546 (N_1546,N_992,N_836);
nor U1547 (N_1547,N_1379,N_1446);
and U1548 (N_1548,N_1020,N_985);
nor U1549 (N_1549,N_878,N_893);
nand U1550 (N_1550,N_1241,N_1189);
nor U1551 (N_1551,N_821,N_1239);
nor U1552 (N_1552,N_1001,N_1280);
and U1553 (N_1553,N_869,N_1283);
or U1554 (N_1554,N_1143,N_897);
or U1555 (N_1555,N_860,N_1438);
and U1556 (N_1556,N_989,N_1384);
nand U1557 (N_1557,N_1139,N_1030);
nand U1558 (N_1558,N_991,N_879);
or U1559 (N_1559,N_1314,N_1075);
xnor U1560 (N_1560,N_1361,N_1216);
or U1561 (N_1561,N_964,N_753);
nand U1562 (N_1562,N_1114,N_912);
or U1563 (N_1563,N_1385,N_837);
nand U1564 (N_1564,N_1331,N_1425);
xor U1565 (N_1565,N_1150,N_1434);
nand U1566 (N_1566,N_1102,N_1182);
or U1567 (N_1567,N_954,N_825);
nand U1568 (N_1568,N_1419,N_1468);
nor U1569 (N_1569,N_1437,N_1256);
nor U1570 (N_1570,N_1166,N_1105);
nor U1571 (N_1571,N_1190,N_1360);
nand U1572 (N_1572,N_1276,N_873);
and U1573 (N_1573,N_790,N_920);
xor U1574 (N_1574,N_1035,N_892);
and U1575 (N_1575,N_816,N_1092);
and U1576 (N_1576,N_1457,N_1375);
nor U1577 (N_1577,N_1366,N_1115);
nor U1578 (N_1578,N_1465,N_1279);
nor U1579 (N_1579,N_1153,N_819);
xor U1580 (N_1580,N_846,N_1281);
nor U1581 (N_1581,N_1091,N_986);
nor U1582 (N_1582,N_1485,N_1297);
and U1583 (N_1583,N_990,N_1164);
xnor U1584 (N_1584,N_960,N_1106);
and U1585 (N_1585,N_1240,N_1146);
nor U1586 (N_1586,N_1204,N_1155);
nor U1587 (N_1587,N_802,N_1218);
nand U1588 (N_1588,N_1179,N_1300);
xor U1589 (N_1589,N_1144,N_1110);
nor U1590 (N_1590,N_1122,N_1161);
or U1591 (N_1591,N_1074,N_1017);
and U1592 (N_1592,N_1082,N_1039);
and U1593 (N_1593,N_1093,N_1253);
or U1594 (N_1594,N_1014,N_1449);
nor U1595 (N_1595,N_1125,N_1442);
nand U1596 (N_1596,N_759,N_907);
or U1597 (N_1597,N_870,N_1307);
or U1598 (N_1598,N_1334,N_774);
xor U1599 (N_1599,N_1065,N_1209);
nand U1600 (N_1600,N_1480,N_1111);
and U1601 (N_1601,N_1466,N_1337);
and U1602 (N_1602,N_1121,N_1367);
nor U1603 (N_1603,N_796,N_984);
and U1604 (N_1604,N_1056,N_932);
or U1605 (N_1605,N_1390,N_787);
and U1606 (N_1606,N_968,N_1259);
nor U1607 (N_1607,N_939,N_959);
or U1608 (N_1608,N_945,N_1372);
xor U1609 (N_1609,N_996,N_1396);
and U1610 (N_1610,N_1244,N_1152);
xor U1611 (N_1611,N_1381,N_1011);
or U1612 (N_1612,N_1345,N_1067);
nand U1613 (N_1613,N_1397,N_886);
xor U1614 (N_1614,N_1365,N_1026);
nand U1615 (N_1615,N_810,N_1172);
nor U1616 (N_1616,N_1195,N_981);
nand U1617 (N_1617,N_1265,N_1350);
or U1618 (N_1618,N_828,N_1488);
nor U1619 (N_1619,N_987,N_921);
or U1620 (N_1620,N_793,N_1258);
nor U1621 (N_1621,N_1309,N_1185);
nand U1622 (N_1622,N_1126,N_1472);
xnor U1623 (N_1623,N_809,N_758);
nand U1624 (N_1624,N_1374,N_835);
and U1625 (N_1625,N_1176,N_1136);
nand U1626 (N_1626,N_1130,N_824);
and U1627 (N_1627,N_914,N_1078);
or U1628 (N_1628,N_1277,N_1420);
xor U1629 (N_1629,N_1066,N_970);
or U1630 (N_1630,N_843,N_789);
or U1631 (N_1631,N_1233,N_1036);
nand U1632 (N_1632,N_1271,N_1203);
or U1633 (N_1633,N_1205,N_788);
or U1634 (N_1634,N_1217,N_777);
nand U1635 (N_1635,N_1431,N_803);
and U1636 (N_1636,N_910,N_1455);
nand U1637 (N_1637,N_1398,N_1387);
or U1638 (N_1638,N_1363,N_1090);
or U1639 (N_1639,N_1016,N_923);
and U1640 (N_1640,N_1096,N_1193);
or U1641 (N_1641,N_931,N_1290);
nand U1642 (N_1642,N_1022,N_1025);
or U1643 (N_1643,N_1422,N_926);
nor U1644 (N_1644,N_1481,N_1170);
or U1645 (N_1645,N_1497,N_1474);
and U1646 (N_1646,N_1007,N_1358);
and U1647 (N_1647,N_1178,N_1284);
or U1648 (N_1648,N_1412,N_1148);
nand U1649 (N_1649,N_1326,N_855);
nor U1650 (N_1650,N_1429,N_1183);
and U1651 (N_1651,N_1417,N_1127);
nor U1652 (N_1652,N_1042,N_1117);
and U1653 (N_1653,N_1181,N_1351);
and U1654 (N_1654,N_1201,N_1289);
or U1655 (N_1655,N_881,N_937);
nor U1656 (N_1656,N_1230,N_993);
and U1657 (N_1657,N_1058,N_1162);
or U1658 (N_1658,N_1080,N_1247);
nand U1659 (N_1659,N_1432,N_1225);
and U1660 (N_1660,N_1054,N_867);
or U1661 (N_1661,N_1404,N_871);
and U1662 (N_1662,N_799,N_850);
nand U1663 (N_1663,N_1221,N_1407);
and U1664 (N_1664,N_768,N_944);
nand U1665 (N_1665,N_1338,N_1059);
nand U1666 (N_1666,N_847,N_961);
nor U1667 (N_1667,N_952,N_1109);
and U1668 (N_1668,N_1000,N_1352);
nor U1669 (N_1669,N_894,N_946);
xor U1670 (N_1670,N_1186,N_769);
xor U1671 (N_1671,N_1131,N_950);
and U1672 (N_1672,N_1167,N_854);
and U1673 (N_1673,N_844,N_1062);
and U1674 (N_1674,N_973,N_1027);
and U1675 (N_1675,N_969,N_1292);
and U1676 (N_1676,N_751,N_1103);
xnor U1677 (N_1677,N_1248,N_1344);
or U1678 (N_1678,N_1234,N_1034);
or U1679 (N_1679,N_1177,N_766);
and U1680 (N_1680,N_1275,N_1198);
or U1681 (N_1681,N_1083,N_928);
nor U1682 (N_1682,N_1145,N_827);
or U1683 (N_1683,N_1473,N_1113);
nand U1684 (N_1684,N_784,N_1128);
or U1685 (N_1685,N_1202,N_853);
and U1686 (N_1686,N_1441,N_998);
nand U1687 (N_1687,N_1427,N_1430);
xor U1688 (N_1688,N_1264,N_1151);
or U1689 (N_1689,N_1119,N_1116);
and U1690 (N_1690,N_1332,N_1424);
nand U1691 (N_1691,N_909,N_1298);
or U1692 (N_1692,N_1440,N_1050);
and U1693 (N_1693,N_1100,N_815);
or U1694 (N_1694,N_1490,N_1245);
or U1695 (N_1695,N_807,N_975);
xor U1696 (N_1696,N_1408,N_955);
nor U1697 (N_1697,N_1101,N_965);
nand U1698 (N_1698,N_848,N_1072);
or U1699 (N_1699,N_1423,N_1308);
and U1700 (N_1700,N_1211,N_1063);
nand U1701 (N_1701,N_785,N_1060);
nand U1702 (N_1702,N_1333,N_884);
nor U1703 (N_1703,N_1312,N_1257);
or U1704 (N_1704,N_1392,N_1255);
or U1705 (N_1705,N_905,N_1008);
or U1706 (N_1706,N_983,N_780);
or U1707 (N_1707,N_967,N_763);
nand U1708 (N_1708,N_808,N_1077);
or U1709 (N_1709,N_1032,N_800);
or U1710 (N_1710,N_918,N_1142);
nand U1711 (N_1711,N_887,N_1341);
or U1712 (N_1712,N_1210,N_1071);
xnor U1713 (N_1713,N_1123,N_1199);
nand U1714 (N_1714,N_1157,N_1310);
and U1715 (N_1715,N_775,N_755);
xor U1716 (N_1716,N_902,N_805);
or U1717 (N_1717,N_900,N_1320);
xnor U1718 (N_1718,N_1315,N_1012);
nand U1719 (N_1719,N_1452,N_1383);
nor U1720 (N_1720,N_1231,N_1019);
nand U1721 (N_1721,N_1306,N_1499);
nand U1722 (N_1722,N_773,N_754);
nand U1723 (N_1723,N_797,N_1133);
xor U1724 (N_1724,N_1393,N_1243);
nand U1725 (N_1725,N_1305,N_830);
or U1726 (N_1726,N_977,N_767);
or U1727 (N_1727,N_1483,N_804);
nor U1728 (N_1728,N_972,N_1319);
or U1729 (N_1729,N_1364,N_781);
nand U1730 (N_1730,N_1251,N_1395);
or U1731 (N_1731,N_1453,N_1076);
and U1732 (N_1732,N_908,N_1169);
xnor U1733 (N_1733,N_1339,N_1378);
and U1734 (N_1734,N_1187,N_770);
and U1735 (N_1735,N_1098,N_916);
nand U1736 (N_1736,N_1175,N_1303);
nor U1737 (N_1737,N_1084,N_1311);
nand U1738 (N_1738,N_1456,N_1478);
and U1739 (N_1739,N_1489,N_1470);
xor U1740 (N_1740,N_1460,N_1137);
and U1741 (N_1741,N_1444,N_1180);
nand U1742 (N_1742,N_1462,N_933);
nor U1743 (N_1743,N_997,N_792);
nor U1744 (N_1744,N_1229,N_1353);
or U1745 (N_1745,N_1347,N_786);
or U1746 (N_1746,N_982,N_1235);
nand U1747 (N_1747,N_1266,N_1246);
or U1748 (N_1748,N_1149,N_1191);
nand U1749 (N_1749,N_1287,N_1406);
and U1750 (N_1750,N_1433,N_1386);
nand U1751 (N_1751,N_1041,N_1159);
or U1752 (N_1752,N_1291,N_833);
nor U1753 (N_1753,N_951,N_956);
or U1754 (N_1754,N_1108,N_1492);
and U1755 (N_1755,N_1223,N_1254);
xnor U1756 (N_1756,N_1329,N_1371);
nand U1757 (N_1757,N_1476,N_1389);
nor U1758 (N_1758,N_1021,N_1296);
or U1759 (N_1759,N_1416,N_1224);
and U1760 (N_1760,N_934,N_1052);
nand U1761 (N_1761,N_1140,N_1458);
nor U1762 (N_1762,N_1031,N_1192);
nor U1763 (N_1763,N_1138,N_1134);
nand U1764 (N_1764,N_840,N_974);
or U1765 (N_1765,N_1405,N_1435);
or U1766 (N_1766,N_943,N_1079);
nor U1767 (N_1767,N_1242,N_1491);
or U1768 (N_1768,N_1346,N_1160);
nor U1769 (N_1769,N_1282,N_822);
nor U1770 (N_1770,N_1048,N_896);
nor U1771 (N_1771,N_958,N_1464);
and U1772 (N_1772,N_852,N_906);
or U1773 (N_1773,N_1328,N_1321);
and U1774 (N_1774,N_1343,N_863);
nor U1775 (N_1775,N_1212,N_1323);
and U1776 (N_1776,N_756,N_1154);
or U1777 (N_1777,N_841,N_1104);
nand U1778 (N_1778,N_978,N_834);
and U1779 (N_1779,N_988,N_1168);
xnor U1780 (N_1780,N_1415,N_1495);
and U1781 (N_1781,N_1428,N_864);
nor U1782 (N_1782,N_1401,N_1135);
and U1783 (N_1783,N_1207,N_1272);
nor U1784 (N_1784,N_1085,N_806);
nor U1785 (N_1785,N_1439,N_966);
nor U1786 (N_1786,N_1482,N_1023);
and U1787 (N_1787,N_1411,N_1402);
or U1788 (N_1788,N_1171,N_1024);
or U1789 (N_1789,N_1047,N_1260);
xor U1790 (N_1790,N_1010,N_1454);
or U1791 (N_1791,N_1463,N_1094);
and U1792 (N_1792,N_876,N_868);
nand U1793 (N_1793,N_917,N_760);
nand U1794 (N_1794,N_885,N_1222);
nand U1795 (N_1795,N_1206,N_842);
and U1796 (N_1796,N_1368,N_1286);
nor U1797 (N_1797,N_904,N_1124);
xnor U1798 (N_1798,N_1087,N_1295);
nor U1799 (N_1799,N_811,N_772);
and U1800 (N_1800,N_1252,N_1325);
and U1801 (N_1801,N_971,N_1317);
nand U1802 (N_1802,N_1107,N_942);
and U1803 (N_1803,N_976,N_927);
nand U1804 (N_1804,N_1493,N_1294);
nand U1805 (N_1805,N_1213,N_947);
or U1806 (N_1806,N_1471,N_1249);
and U1807 (N_1807,N_940,N_849);
nor U1808 (N_1808,N_1051,N_1262);
xnor U1809 (N_1809,N_1188,N_883);
nor U1810 (N_1810,N_875,N_953);
and U1811 (N_1811,N_839,N_1459);
and U1812 (N_1812,N_1132,N_1335);
and U1813 (N_1813,N_1410,N_962);
or U1814 (N_1814,N_1445,N_1197);
or U1815 (N_1815,N_820,N_779);
nand U1816 (N_1816,N_1156,N_1340);
and U1817 (N_1817,N_1055,N_776);
nor U1818 (N_1818,N_924,N_1194);
or U1819 (N_1819,N_817,N_801);
nor U1820 (N_1820,N_1327,N_1147);
nor U1821 (N_1821,N_1403,N_1450);
or U1822 (N_1822,N_814,N_1354);
nor U1823 (N_1823,N_1362,N_813);
nand U1824 (N_1824,N_1484,N_857);
nor U1825 (N_1825,N_851,N_1081);
nand U1826 (N_1826,N_1228,N_1426);
nor U1827 (N_1827,N_861,N_898);
and U1828 (N_1828,N_903,N_1158);
nand U1829 (N_1829,N_866,N_1174);
nand U1830 (N_1830,N_1061,N_1269);
nor U1831 (N_1831,N_1049,N_1165);
nand U1832 (N_1832,N_936,N_1226);
and U1833 (N_1833,N_1443,N_1088);
and U1834 (N_1834,N_1044,N_1356);
or U1835 (N_1835,N_1267,N_1232);
or U1836 (N_1836,N_980,N_757);
or U1837 (N_1837,N_1447,N_1342);
nand U1838 (N_1838,N_1004,N_1487);
nand U1839 (N_1839,N_1418,N_831);
and U1840 (N_1840,N_1214,N_1324);
nor U1841 (N_1841,N_1173,N_1373);
or U1842 (N_1842,N_882,N_823);
nand U1843 (N_1843,N_872,N_1040);
or U1844 (N_1844,N_1053,N_1045);
and U1845 (N_1845,N_963,N_865);
nand U1846 (N_1846,N_1099,N_1370);
or U1847 (N_1847,N_911,N_1208);
or U1848 (N_1848,N_1009,N_1479);
xor U1849 (N_1849,N_791,N_1029);
nor U1850 (N_1850,N_1436,N_1129);
nand U1851 (N_1851,N_1005,N_1399);
or U1852 (N_1852,N_1069,N_1018);
and U1853 (N_1853,N_762,N_1475);
and U1854 (N_1854,N_812,N_890);
xor U1855 (N_1855,N_771,N_1097);
nor U1856 (N_1856,N_877,N_778);
and U1857 (N_1857,N_750,N_1215);
or U1858 (N_1858,N_901,N_1377);
xnor U1859 (N_1859,N_1015,N_856);
or U1860 (N_1860,N_1268,N_1038);
nand U1861 (N_1861,N_929,N_1002);
nand U1862 (N_1862,N_1270,N_1163);
nor U1863 (N_1863,N_845,N_1414);
nor U1864 (N_1864,N_1477,N_1355);
and U1865 (N_1865,N_1288,N_1336);
nor U1866 (N_1866,N_1064,N_862);
nor U1867 (N_1867,N_1316,N_1461);
nand U1868 (N_1868,N_1313,N_1382);
nand U1869 (N_1869,N_874,N_1003);
nand U1870 (N_1870,N_1494,N_1421);
and U1871 (N_1871,N_1394,N_1301);
and U1872 (N_1872,N_1357,N_925);
or U1873 (N_1873,N_1467,N_782);
or U1874 (N_1874,N_832,N_1220);
nand U1875 (N_1875,N_905,N_1442);
or U1876 (N_1876,N_1106,N_809);
nor U1877 (N_1877,N_1228,N_1085);
and U1878 (N_1878,N_1055,N_832);
nand U1879 (N_1879,N_997,N_1068);
and U1880 (N_1880,N_1102,N_797);
nand U1881 (N_1881,N_837,N_1145);
nand U1882 (N_1882,N_1340,N_1188);
nor U1883 (N_1883,N_954,N_1133);
xnor U1884 (N_1884,N_1402,N_1382);
nand U1885 (N_1885,N_913,N_1304);
nor U1886 (N_1886,N_1148,N_771);
or U1887 (N_1887,N_1285,N_1032);
xor U1888 (N_1888,N_993,N_804);
nand U1889 (N_1889,N_788,N_1216);
or U1890 (N_1890,N_911,N_1485);
nor U1891 (N_1891,N_1375,N_1085);
nand U1892 (N_1892,N_1227,N_911);
or U1893 (N_1893,N_1204,N_936);
nor U1894 (N_1894,N_1265,N_1428);
nor U1895 (N_1895,N_1081,N_841);
or U1896 (N_1896,N_1471,N_1465);
and U1897 (N_1897,N_794,N_1034);
nor U1898 (N_1898,N_985,N_1148);
and U1899 (N_1899,N_1470,N_1176);
nand U1900 (N_1900,N_1006,N_877);
xnor U1901 (N_1901,N_1309,N_1206);
and U1902 (N_1902,N_962,N_807);
or U1903 (N_1903,N_1188,N_1448);
and U1904 (N_1904,N_955,N_1102);
nor U1905 (N_1905,N_1259,N_1409);
nor U1906 (N_1906,N_1043,N_1493);
and U1907 (N_1907,N_824,N_762);
xor U1908 (N_1908,N_1295,N_1271);
and U1909 (N_1909,N_1398,N_1184);
nor U1910 (N_1910,N_1323,N_895);
nand U1911 (N_1911,N_1274,N_1170);
and U1912 (N_1912,N_1332,N_1440);
nand U1913 (N_1913,N_981,N_1360);
and U1914 (N_1914,N_1365,N_946);
nand U1915 (N_1915,N_1124,N_1291);
nand U1916 (N_1916,N_805,N_929);
and U1917 (N_1917,N_914,N_1199);
nand U1918 (N_1918,N_1372,N_1056);
or U1919 (N_1919,N_1151,N_950);
or U1920 (N_1920,N_1183,N_983);
and U1921 (N_1921,N_1391,N_1485);
and U1922 (N_1922,N_1488,N_1279);
nor U1923 (N_1923,N_756,N_1417);
or U1924 (N_1924,N_828,N_1406);
or U1925 (N_1925,N_1395,N_1414);
and U1926 (N_1926,N_970,N_780);
nand U1927 (N_1927,N_1145,N_1314);
nand U1928 (N_1928,N_859,N_1460);
and U1929 (N_1929,N_1009,N_1389);
and U1930 (N_1930,N_1313,N_1352);
nor U1931 (N_1931,N_1303,N_1205);
nand U1932 (N_1932,N_1415,N_1054);
and U1933 (N_1933,N_1328,N_901);
nor U1934 (N_1934,N_968,N_756);
nor U1935 (N_1935,N_1223,N_1198);
nor U1936 (N_1936,N_934,N_1477);
nand U1937 (N_1937,N_868,N_901);
and U1938 (N_1938,N_1083,N_1432);
nor U1939 (N_1939,N_1298,N_868);
and U1940 (N_1940,N_811,N_998);
nand U1941 (N_1941,N_1217,N_946);
nor U1942 (N_1942,N_1027,N_870);
or U1943 (N_1943,N_1230,N_1373);
and U1944 (N_1944,N_1403,N_1387);
nor U1945 (N_1945,N_1027,N_1283);
nor U1946 (N_1946,N_1240,N_1475);
and U1947 (N_1947,N_1446,N_1134);
nor U1948 (N_1948,N_1050,N_1314);
nand U1949 (N_1949,N_1405,N_989);
nand U1950 (N_1950,N_1161,N_1412);
nor U1951 (N_1951,N_1153,N_1099);
xor U1952 (N_1952,N_1177,N_1081);
nand U1953 (N_1953,N_844,N_1231);
nand U1954 (N_1954,N_1027,N_998);
and U1955 (N_1955,N_1401,N_1105);
xor U1956 (N_1956,N_1143,N_1449);
nand U1957 (N_1957,N_831,N_1293);
xnor U1958 (N_1958,N_1253,N_930);
and U1959 (N_1959,N_997,N_1475);
and U1960 (N_1960,N_933,N_1056);
or U1961 (N_1961,N_1427,N_1237);
or U1962 (N_1962,N_1425,N_767);
nor U1963 (N_1963,N_872,N_1440);
and U1964 (N_1964,N_895,N_1463);
nand U1965 (N_1965,N_906,N_934);
nor U1966 (N_1966,N_1253,N_1083);
nor U1967 (N_1967,N_1258,N_1009);
and U1968 (N_1968,N_1459,N_1206);
nor U1969 (N_1969,N_799,N_882);
or U1970 (N_1970,N_978,N_1364);
nor U1971 (N_1971,N_1486,N_1331);
or U1972 (N_1972,N_1030,N_829);
or U1973 (N_1973,N_1401,N_1478);
and U1974 (N_1974,N_792,N_1037);
nand U1975 (N_1975,N_1269,N_826);
and U1976 (N_1976,N_1177,N_1245);
xor U1977 (N_1977,N_875,N_753);
or U1978 (N_1978,N_1211,N_1308);
or U1979 (N_1979,N_1095,N_952);
or U1980 (N_1980,N_1224,N_952);
or U1981 (N_1981,N_1357,N_1438);
nor U1982 (N_1982,N_1142,N_1264);
and U1983 (N_1983,N_761,N_1069);
and U1984 (N_1984,N_1344,N_1478);
and U1985 (N_1985,N_919,N_821);
nand U1986 (N_1986,N_1468,N_1459);
nand U1987 (N_1987,N_1304,N_766);
or U1988 (N_1988,N_816,N_1405);
xnor U1989 (N_1989,N_1007,N_1006);
xor U1990 (N_1990,N_1446,N_1042);
and U1991 (N_1991,N_1183,N_1002);
and U1992 (N_1992,N_1489,N_917);
xor U1993 (N_1993,N_1058,N_777);
and U1994 (N_1994,N_1388,N_1296);
and U1995 (N_1995,N_1161,N_1114);
or U1996 (N_1996,N_1279,N_940);
nand U1997 (N_1997,N_1270,N_1045);
xnor U1998 (N_1998,N_1415,N_919);
xnor U1999 (N_1999,N_935,N_1317);
or U2000 (N_2000,N_853,N_1085);
nor U2001 (N_2001,N_1109,N_945);
and U2002 (N_2002,N_1422,N_1225);
nand U2003 (N_2003,N_937,N_1364);
nand U2004 (N_2004,N_1018,N_883);
nor U2005 (N_2005,N_1073,N_881);
nor U2006 (N_2006,N_1426,N_1059);
xnor U2007 (N_2007,N_1457,N_1314);
xor U2008 (N_2008,N_1276,N_1252);
and U2009 (N_2009,N_846,N_881);
or U2010 (N_2010,N_1428,N_996);
nand U2011 (N_2011,N_1448,N_1325);
and U2012 (N_2012,N_1068,N_1328);
nand U2013 (N_2013,N_1002,N_1132);
nor U2014 (N_2014,N_1095,N_1274);
xnor U2015 (N_2015,N_1178,N_1176);
or U2016 (N_2016,N_1129,N_1015);
nand U2017 (N_2017,N_1036,N_853);
nor U2018 (N_2018,N_909,N_893);
or U2019 (N_2019,N_977,N_794);
nand U2020 (N_2020,N_1225,N_1216);
nor U2021 (N_2021,N_1054,N_751);
or U2022 (N_2022,N_1183,N_1488);
and U2023 (N_2023,N_1077,N_1209);
nand U2024 (N_2024,N_1266,N_1315);
and U2025 (N_2025,N_1186,N_796);
nand U2026 (N_2026,N_837,N_999);
nand U2027 (N_2027,N_896,N_1137);
nand U2028 (N_2028,N_965,N_951);
and U2029 (N_2029,N_1211,N_1364);
xor U2030 (N_2030,N_1443,N_793);
nand U2031 (N_2031,N_963,N_1203);
or U2032 (N_2032,N_1231,N_1211);
and U2033 (N_2033,N_1144,N_1041);
xnor U2034 (N_2034,N_857,N_776);
nand U2035 (N_2035,N_1020,N_1439);
nor U2036 (N_2036,N_1332,N_1309);
nor U2037 (N_2037,N_973,N_1090);
and U2038 (N_2038,N_1148,N_867);
nand U2039 (N_2039,N_983,N_754);
or U2040 (N_2040,N_1098,N_1069);
nand U2041 (N_2041,N_955,N_1153);
or U2042 (N_2042,N_1001,N_1198);
and U2043 (N_2043,N_1312,N_947);
and U2044 (N_2044,N_778,N_1408);
nand U2045 (N_2045,N_772,N_1493);
nand U2046 (N_2046,N_1493,N_821);
or U2047 (N_2047,N_1152,N_794);
and U2048 (N_2048,N_1020,N_1234);
and U2049 (N_2049,N_1213,N_946);
nand U2050 (N_2050,N_814,N_1087);
nand U2051 (N_2051,N_976,N_1332);
or U2052 (N_2052,N_1230,N_1231);
nand U2053 (N_2053,N_1280,N_1245);
or U2054 (N_2054,N_1371,N_1312);
and U2055 (N_2055,N_760,N_1235);
nand U2056 (N_2056,N_883,N_922);
nand U2057 (N_2057,N_996,N_1194);
or U2058 (N_2058,N_1231,N_760);
nor U2059 (N_2059,N_1011,N_867);
and U2060 (N_2060,N_872,N_866);
xor U2061 (N_2061,N_1319,N_837);
or U2062 (N_2062,N_1487,N_838);
and U2063 (N_2063,N_1050,N_826);
xor U2064 (N_2064,N_1129,N_1038);
nand U2065 (N_2065,N_781,N_1138);
nand U2066 (N_2066,N_1223,N_1090);
or U2067 (N_2067,N_1296,N_809);
nor U2068 (N_2068,N_1087,N_767);
and U2069 (N_2069,N_1373,N_923);
or U2070 (N_2070,N_1060,N_938);
nor U2071 (N_2071,N_1234,N_1159);
or U2072 (N_2072,N_1361,N_873);
nor U2073 (N_2073,N_1165,N_1381);
or U2074 (N_2074,N_1460,N_842);
and U2075 (N_2075,N_1028,N_1493);
nand U2076 (N_2076,N_936,N_1397);
xnor U2077 (N_2077,N_980,N_1107);
or U2078 (N_2078,N_1111,N_898);
and U2079 (N_2079,N_1128,N_1208);
or U2080 (N_2080,N_1278,N_838);
nand U2081 (N_2081,N_1065,N_1486);
or U2082 (N_2082,N_1232,N_1046);
and U2083 (N_2083,N_988,N_1347);
nor U2084 (N_2084,N_812,N_886);
or U2085 (N_2085,N_1376,N_1372);
nor U2086 (N_2086,N_754,N_1133);
or U2087 (N_2087,N_1072,N_1386);
nand U2088 (N_2088,N_1192,N_838);
and U2089 (N_2089,N_1117,N_1214);
or U2090 (N_2090,N_1009,N_793);
nor U2091 (N_2091,N_1054,N_825);
nor U2092 (N_2092,N_1413,N_787);
nor U2093 (N_2093,N_1468,N_1221);
or U2094 (N_2094,N_1314,N_1382);
or U2095 (N_2095,N_1072,N_1457);
nand U2096 (N_2096,N_1267,N_841);
xnor U2097 (N_2097,N_1482,N_1181);
nand U2098 (N_2098,N_1144,N_927);
and U2099 (N_2099,N_1411,N_987);
or U2100 (N_2100,N_859,N_1040);
and U2101 (N_2101,N_1030,N_929);
and U2102 (N_2102,N_1194,N_1055);
nand U2103 (N_2103,N_971,N_1473);
or U2104 (N_2104,N_1468,N_996);
and U2105 (N_2105,N_1401,N_1369);
xnor U2106 (N_2106,N_874,N_1087);
nor U2107 (N_2107,N_1400,N_1427);
and U2108 (N_2108,N_1093,N_1361);
or U2109 (N_2109,N_1026,N_1181);
nor U2110 (N_2110,N_752,N_825);
and U2111 (N_2111,N_944,N_1349);
xnor U2112 (N_2112,N_1287,N_1316);
nand U2113 (N_2113,N_1245,N_960);
or U2114 (N_2114,N_964,N_1459);
xor U2115 (N_2115,N_1005,N_754);
nor U2116 (N_2116,N_1125,N_1059);
or U2117 (N_2117,N_1298,N_1103);
nand U2118 (N_2118,N_1277,N_936);
or U2119 (N_2119,N_876,N_1347);
and U2120 (N_2120,N_1234,N_1193);
nand U2121 (N_2121,N_1143,N_1279);
nor U2122 (N_2122,N_1416,N_1186);
nand U2123 (N_2123,N_1280,N_1110);
nor U2124 (N_2124,N_1183,N_1125);
or U2125 (N_2125,N_763,N_1271);
nor U2126 (N_2126,N_1437,N_1001);
or U2127 (N_2127,N_1345,N_914);
or U2128 (N_2128,N_777,N_1307);
or U2129 (N_2129,N_1438,N_757);
xnor U2130 (N_2130,N_1290,N_1040);
nor U2131 (N_2131,N_1365,N_926);
nand U2132 (N_2132,N_1096,N_1344);
nor U2133 (N_2133,N_958,N_940);
or U2134 (N_2134,N_1154,N_912);
nand U2135 (N_2135,N_913,N_1246);
nor U2136 (N_2136,N_832,N_1362);
nand U2137 (N_2137,N_1025,N_1325);
xnor U2138 (N_2138,N_1378,N_894);
nand U2139 (N_2139,N_1117,N_1419);
and U2140 (N_2140,N_1020,N_1091);
nand U2141 (N_2141,N_1005,N_1032);
xnor U2142 (N_2142,N_930,N_992);
or U2143 (N_2143,N_1331,N_954);
xor U2144 (N_2144,N_891,N_1121);
or U2145 (N_2145,N_895,N_898);
nand U2146 (N_2146,N_1303,N_1377);
and U2147 (N_2147,N_1412,N_819);
xnor U2148 (N_2148,N_830,N_1328);
and U2149 (N_2149,N_1143,N_1172);
and U2150 (N_2150,N_1020,N_786);
nor U2151 (N_2151,N_875,N_1405);
or U2152 (N_2152,N_1210,N_1051);
nor U2153 (N_2153,N_1064,N_857);
or U2154 (N_2154,N_1238,N_1457);
nor U2155 (N_2155,N_787,N_1013);
and U2156 (N_2156,N_1204,N_787);
nor U2157 (N_2157,N_1187,N_978);
and U2158 (N_2158,N_1382,N_794);
and U2159 (N_2159,N_1067,N_1104);
nand U2160 (N_2160,N_1476,N_931);
and U2161 (N_2161,N_1264,N_1273);
nor U2162 (N_2162,N_1162,N_1294);
nand U2163 (N_2163,N_1197,N_1394);
and U2164 (N_2164,N_989,N_820);
or U2165 (N_2165,N_1035,N_1194);
nand U2166 (N_2166,N_1157,N_1081);
or U2167 (N_2167,N_919,N_1301);
or U2168 (N_2168,N_1346,N_1074);
or U2169 (N_2169,N_1035,N_1255);
or U2170 (N_2170,N_1406,N_1189);
nand U2171 (N_2171,N_1173,N_1450);
nand U2172 (N_2172,N_904,N_1105);
nor U2173 (N_2173,N_1078,N_1412);
nor U2174 (N_2174,N_882,N_1405);
or U2175 (N_2175,N_775,N_1448);
or U2176 (N_2176,N_1263,N_1271);
and U2177 (N_2177,N_1010,N_1345);
nand U2178 (N_2178,N_802,N_1165);
and U2179 (N_2179,N_1445,N_1162);
nand U2180 (N_2180,N_964,N_927);
xnor U2181 (N_2181,N_1136,N_1376);
nand U2182 (N_2182,N_1220,N_837);
or U2183 (N_2183,N_1101,N_1321);
or U2184 (N_2184,N_978,N_1058);
nor U2185 (N_2185,N_1244,N_1193);
or U2186 (N_2186,N_893,N_1303);
or U2187 (N_2187,N_1441,N_750);
nor U2188 (N_2188,N_1204,N_1306);
and U2189 (N_2189,N_1334,N_1368);
nor U2190 (N_2190,N_790,N_1382);
nand U2191 (N_2191,N_1283,N_1450);
nand U2192 (N_2192,N_1116,N_1335);
and U2193 (N_2193,N_1458,N_1152);
nor U2194 (N_2194,N_1057,N_1345);
nor U2195 (N_2195,N_1093,N_892);
or U2196 (N_2196,N_1024,N_817);
or U2197 (N_2197,N_1213,N_1457);
nor U2198 (N_2198,N_1274,N_864);
and U2199 (N_2199,N_1398,N_1197);
nand U2200 (N_2200,N_1348,N_818);
and U2201 (N_2201,N_1476,N_1302);
xor U2202 (N_2202,N_1183,N_841);
nor U2203 (N_2203,N_1323,N_1444);
nor U2204 (N_2204,N_1498,N_1215);
nand U2205 (N_2205,N_964,N_1210);
nand U2206 (N_2206,N_956,N_966);
nor U2207 (N_2207,N_1118,N_1282);
nand U2208 (N_2208,N_819,N_796);
nor U2209 (N_2209,N_942,N_933);
nand U2210 (N_2210,N_1275,N_1457);
and U2211 (N_2211,N_1409,N_853);
xnor U2212 (N_2212,N_1118,N_1020);
xnor U2213 (N_2213,N_1161,N_938);
and U2214 (N_2214,N_1027,N_1172);
or U2215 (N_2215,N_926,N_1155);
nor U2216 (N_2216,N_1110,N_1281);
and U2217 (N_2217,N_928,N_1449);
xnor U2218 (N_2218,N_884,N_1114);
nor U2219 (N_2219,N_1491,N_1087);
and U2220 (N_2220,N_1440,N_1011);
xnor U2221 (N_2221,N_1303,N_1269);
nand U2222 (N_2222,N_773,N_1115);
nor U2223 (N_2223,N_1241,N_1270);
nor U2224 (N_2224,N_1048,N_946);
nand U2225 (N_2225,N_974,N_1175);
nor U2226 (N_2226,N_1016,N_1376);
and U2227 (N_2227,N_1163,N_769);
or U2228 (N_2228,N_981,N_922);
xor U2229 (N_2229,N_1415,N_1311);
nor U2230 (N_2230,N_962,N_892);
or U2231 (N_2231,N_1084,N_847);
or U2232 (N_2232,N_855,N_1393);
and U2233 (N_2233,N_1328,N_778);
nor U2234 (N_2234,N_1469,N_1446);
or U2235 (N_2235,N_1475,N_950);
or U2236 (N_2236,N_1045,N_1227);
nand U2237 (N_2237,N_1156,N_1136);
nor U2238 (N_2238,N_1451,N_844);
and U2239 (N_2239,N_1481,N_910);
and U2240 (N_2240,N_1200,N_1159);
nand U2241 (N_2241,N_860,N_1352);
nand U2242 (N_2242,N_1446,N_1431);
and U2243 (N_2243,N_845,N_1146);
nor U2244 (N_2244,N_989,N_1239);
or U2245 (N_2245,N_1448,N_1071);
nand U2246 (N_2246,N_1085,N_928);
xor U2247 (N_2247,N_838,N_853);
and U2248 (N_2248,N_965,N_788);
and U2249 (N_2249,N_1058,N_1260);
and U2250 (N_2250,N_1852,N_1789);
nor U2251 (N_2251,N_2044,N_1661);
nor U2252 (N_2252,N_1722,N_1836);
nor U2253 (N_2253,N_1608,N_1683);
or U2254 (N_2254,N_1866,N_1542);
and U2255 (N_2255,N_1856,N_1776);
nor U2256 (N_2256,N_2201,N_2042);
nand U2257 (N_2257,N_1931,N_1923);
xor U2258 (N_2258,N_1927,N_1823);
nor U2259 (N_2259,N_1548,N_2163);
nand U2260 (N_2260,N_2243,N_1687);
or U2261 (N_2261,N_2066,N_1969);
nor U2262 (N_2262,N_1822,N_1582);
xor U2263 (N_2263,N_1863,N_2152);
and U2264 (N_2264,N_1951,N_1587);
nor U2265 (N_2265,N_2135,N_1632);
and U2266 (N_2266,N_2187,N_1524);
nand U2267 (N_2267,N_1790,N_1662);
nand U2268 (N_2268,N_1882,N_1938);
nand U2269 (N_2269,N_1635,N_2249);
nand U2270 (N_2270,N_1623,N_1569);
or U2271 (N_2271,N_1625,N_2200);
nor U2272 (N_2272,N_1619,N_1758);
or U2273 (N_2273,N_1805,N_1685);
or U2274 (N_2274,N_1768,N_1909);
xor U2275 (N_2275,N_1798,N_2079);
and U2276 (N_2276,N_2052,N_1511);
or U2277 (N_2277,N_1679,N_1979);
xnor U2278 (N_2278,N_1804,N_1555);
nand U2279 (N_2279,N_2134,N_2064);
or U2280 (N_2280,N_1967,N_1779);
nand U2281 (N_2281,N_1575,N_1714);
or U2282 (N_2282,N_1638,N_1815);
or U2283 (N_2283,N_2061,N_1868);
and U2284 (N_2284,N_1596,N_2238);
nand U2285 (N_2285,N_1881,N_1601);
nand U2286 (N_2286,N_2221,N_2167);
nor U2287 (N_2287,N_1656,N_1532);
nor U2288 (N_2288,N_2026,N_2231);
nand U2289 (N_2289,N_1978,N_2093);
or U2290 (N_2290,N_1865,N_1915);
nor U2291 (N_2291,N_2192,N_1751);
nand U2292 (N_2292,N_1989,N_2013);
nand U2293 (N_2293,N_1963,N_1810);
nor U2294 (N_2294,N_1535,N_2181);
or U2295 (N_2295,N_2118,N_1669);
nand U2296 (N_2296,N_2233,N_1952);
or U2297 (N_2297,N_1874,N_1795);
nor U2298 (N_2298,N_1585,N_1564);
nor U2299 (N_2299,N_2054,N_1580);
or U2300 (N_2300,N_2119,N_1721);
or U2301 (N_2301,N_1664,N_2127);
nor U2302 (N_2302,N_1750,N_1930);
nand U2303 (N_2303,N_2086,N_1925);
nor U2304 (N_2304,N_2025,N_1743);
xnor U2305 (N_2305,N_2111,N_2043);
or U2306 (N_2306,N_1939,N_1794);
nor U2307 (N_2307,N_1840,N_1787);
or U2308 (N_2308,N_1843,N_2202);
and U2309 (N_2309,N_1870,N_1957);
nand U2310 (N_2310,N_1912,N_1665);
nand U2311 (N_2311,N_2197,N_2145);
nor U2312 (N_2312,N_1616,N_1996);
nand U2313 (N_2313,N_1785,N_1723);
or U2314 (N_2314,N_1579,N_1775);
nor U2315 (N_2315,N_1720,N_2117);
nand U2316 (N_2316,N_1509,N_1657);
nand U2317 (N_2317,N_1913,N_1624);
nand U2318 (N_2318,N_2139,N_2216);
and U2319 (N_2319,N_1695,N_1600);
nor U2320 (N_2320,N_2058,N_1546);
nand U2321 (N_2321,N_2138,N_1816);
xnor U2322 (N_2322,N_2219,N_1835);
nor U2323 (N_2323,N_1604,N_2003);
and U2324 (N_2324,N_1761,N_1910);
nand U2325 (N_2325,N_1936,N_1855);
or U2326 (N_2326,N_1692,N_1641);
nor U2327 (N_2327,N_2188,N_1603);
nand U2328 (N_2328,N_1792,N_1703);
nor U2329 (N_2329,N_1926,N_1598);
xor U2330 (N_2330,N_2039,N_2019);
nor U2331 (N_2331,N_2168,N_1746);
or U2332 (N_2332,N_2091,N_1520);
xnor U2333 (N_2333,N_1534,N_1612);
nand U2334 (N_2334,N_1819,N_2136);
nand U2335 (N_2335,N_1879,N_1999);
and U2336 (N_2336,N_1832,N_2151);
nor U2337 (N_2337,N_1578,N_1588);
and U2338 (N_2338,N_1971,N_1566);
and U2339 (N_2339,N_1607,N_1780);
and U2340 (N_2340,N_1611,N_2171);
and U2341 (N_2341,N_1521,N_1505);
nor U2342 (N_2342,N_1981,N_2012);
and U2343 (N_2343,N_1731,N_1693);
and U2344 (N_2344,N_1892,N_1508);
nand U2345 (N_2345,N_2071,N_2245);
nand U2346 (N_2346,N_1911,N_1988);
and U2347 (N_2347,N_1705,N_1760);
or U2348 (N_2348,N_2063,N_1500);
and U2349 (N_2349,N_2185,N_1965);
or U2350 (N_2350,N_2109,N_2235);
nand U2351 (N_2351,N_1917,N_1771);
nand U2352 (N_2352,N_2072,N_2234);
nor U2353 (N_2353,N_1908,N_2018);
and U2354 (N_2354,N_2080,N_1955);
nand U2355 (N_2355,N_2160,N_2212);
or U2356 (N_2356,N_2107,N_2005);
nand U2357 (N_2357,N_2164,N_1867);
and U2358 (N_2358,N_2149,N_1994);
and U2359 (N_2359,N_2148,N_2030);
nand U2360 (N_2360,N_1735,N_2132);
or U2361 (N_2361,N_2126,N_1956);
and U2362 (N_2362,N_1517,N_2184);
nor U2363 (N_2363,N_1799,N_2236);
xnor U2364 (N_2364,N_2154,N_1992);
nor U2365 (N_2365,N_2011,N_1504);
nand U2366 (N_2366,N_1506,N_1948);
nor U2367 (N_2367,N_1857,N_1976);
nand U2368 (N_2368,N_1529,N_1898);
and U2369 (N_2369,N_1682,N_1554);
or U2370 (N_2370,N_1907,N_1675);
or U2371 (N_2371,N_1968,N_1742);
or U2372 (N_2372,N_1774,N_2244);
nor U2373 (N_2373,N_1518,N_2210);
and U2374 (N_2374,N_1709,N_2170);
nor U2375 (N_2375,N_2240,N_2214);
xor U2376 (N_2376,N_2096,N_1557);
or U2377 (N_2377,N_2015,N_2209);
nand U2378 (N_2378,N_1763,N_2083);
nor U2379 (N_2379,N_2104,N_1839);
nor U2380 (N_2380,N_1561,N_1736);
nor U2381 (N_2381,N_1545,N_1629);
and U2382 (N_2382,N_2116,N_2002);
nor U2383 (N_2383,N_2239,N_1636);
nor U2384 (N_2384,N_2137,N_1523);
or U2385 (N_2385,N_1941,N_1778);
or U2386 (N_2386,N_1552,N_1733);
nand U2387 (N_2387,N_1727,N_2147);
or U2388 (N_2388,N_1536,N_1668);
xnor U2389 (N_2389,N_1618,N_1515);
and U2390 (N_2390,N_2099,N_1929);
nand U2391 (N_2391,N_1858,N_1527);
and U2392 (N_2392,N_1697,N_1614);
nand U2393 (N_2393,N_1688,N_1553);
nand U2394 (N_2394,N_2165,N_2225);
nor U2395 (N_2395,N_1739,N_1655);
nand U2396 (N_2396,N_1689,N_1595);
nand U2397 (N_2397,N_1844,N_2009);
and U2398 (N_2398,N_2237,N_1702);
nor U2399 (N_2399,N_1660,N_1833);
or U2400 (N_2400,N_1560,N_1901);
or U2401 (N_2401,N_2059,N_2194);
xnor U2402 (N_2402,N_2036,N_1762);
nor U2403 (N_2403,N_1872,N_1800);
or U2404 (N_2404,N_2029,N_1627);
nor U2405 (N_2405,N_2112,N_1674);
and U2406 (N_2406,N_2180,N_1617);
nand U2407 (N_2407,N_1772,N_1513);
xnor U2408 (N_2408,N_1550,N_1961);
nand U2409 (N_2409,N_1767,N_1814);
or U2410 (N_2410,N_2041,N_1924);
nor U2411 (N_2411,N_1830,N_1537);
nand U2412 (N_2412,N_1526,N_1900);
nor U2413 (N_2413,N_1549,N_1648);
nor U2414 (N_2414,N_1610,N_1663);
or U2415 (N_2415,N_1701,N_1597);
nand U2416 (N_2416,N_1770,N_1667);
or U2417 (N_2417,N_1748,N_1793);
nor U2418 (N_2418,N_2055,N_2077);
nand U2419 (N_2419,N_1876,N_1574);
and U2420 (N_2420,N_2057,N_1681);
or U2421 (N_2421,N_1543,N_1905);
nand U2422 (N_2422,N_2056,N_1708);
and U2423 (N_2423,N_1841,N_2128);
nand U2424 (N_2424,N_2113,N_1670);
xor U2425 (N_2425,N_2074,N_2046);
and U2426 (N_2426,N_1914,N_1885);
nor U2427 (N_2427,N_1888,N_1713);
nor U2428 (N_2428,N_1686,N_1949);
nand U2429 (N_2429,N_1859,N_2242);
xnor U2430 (N_2430,N_2232,N_2124);
nand U2431 (N_2431,N_1680,N_2172);
xnor U2432 (N_2432,N_1934,N_1920);
and U2433 (N_2433,N_1850,N_1928);
and U2434 (N_2434,N_1943,N_1525);
nor U2435 (N_2435,N_2114,N_1788);
nand U2436 (N_2436,N_1539,N_1747);
nand U2437 (N_2437,N_2204,N_1544);
nand U2438 (N_2438,N_1533,N_2034);
xor U2439 (N_2439,N_1845,N_2199);
xnor U2440 (N_2440,N_2223,N_1541);
and U2441 (N_2441,N_1972,N_1676);
and U2442 (N_2442,N_1710,N_2001);
nand U2443 (N_2443,N_1615,N_2183);
or U2444 (N_2444,N_1706,N_1501);
and U2445 (N_2445,N_1590,N_1950);
and U2446 (N_2446,N_1591,N_2087);
nand U2447 (N_2447,N_2162,N_1922);
nor U2448 (N_2448,N_1983,N_1718);
nand U2449 (N_2449,N_2006,N_1719);
nor U2450 (N_2450,N_1725,N_1824);
or U2451 (N_2451,N_1516,N_1854);
xor U2452 (N_2452,N_1724,N_1820);
and U2453 (N_2453,N_1643,N_1602);
xnor U2454 (N_2454,N_1646,N_1812);
or U2455 (N_2455,N_1609,N_2110);
and U2456 (N_2456,N_1658,N_2174);
xnor U2457 (N_2457,N_1707,N_2203);
nand U2458 (N_2458,N_1887,N_1993);
or U2459 (N_2459,N_2051,N_1884);
and U2460 (N_2460,N_1729,N_1826);
nor U2461 (N_2461,N_1606,N_1985);
nand U2462 (N_2462,N_2218,N_1712);
nor U2463 (N_2463,N_1862,N_1973);
nand U2464 (N_2464,N_1899,N_2198);
and U2465 (N_2465,N_2208,N_1987);
nand U2466 (N_2466,N_1944,N_1842);
and U2467 (N_2467,N_2206,N_2070);
xnor U2468 (N_2468,N_2105,N_1878);
xnor U2469 (N_2469,N_2047,N_2205);
xnor U2470 (N_2470,N_1846,N_1652);
nor U2471 (N_2471,N_1694,N_1984);
nor U2472 (N_2472,N_1869,N_2038);
xnor U2473 (N_2473,N_1570,N_2102);
or U2474 (N_2474,N_1613,N_1903);
or U2475 (N_2475,N_1838,N_2156);
and U2476 (N_2476,N_1797,N_1698);
nor U2477 (N_2477,N_2222,N_2085);
nand U2478 (N_2478,N_2021,N_2241);
nand U2479 (N_2479,N_1519,N_1677);
and U2480 (N_2480,N_2014,N_2040);
nor U2481 (N_2481,N_2207,N_1753);
nand U2482 (N_2482,N_2020,N_1568);
nor U2483 (N_2483,N_1880,N_2226);
nor U2484 (N_2484,N_2065,N_2211);
and U2485 (N_2485,N_2186,N_2022);
and U2486 (N_2486,N_1764,N_1696);
nand U2487 (N_2487,N_1960,N_2246);
nand U2488 (N_2488,N_1847,N_1530);
nor U2489 (N_2489,N_1650,N_1640);
and U2490 (N_2490,N_1730,N_1654);
and U2491 (N_2491,N_1577,N_1673);
nor U2492 (N_2492,N_2196,N_2088);
and U2493 (N_2493,N_1528,N_1726);
or U2494 (N_2494,N_1631,N_2176);
xor U2495 (N_2495,N_2144,N_1808);
nand U2496 (N_2496,N_1558,N_1745);
nor U2497 (N_2497,N_2141,N_1959);
xnor U2498 (N_2498,N_1806,N_1977);
and U2499 (N_2499,N_1576,N_2248);
nor U2500 (N_2500,N_1828,N_1829);
xor U2501 (N_2501,N_1651,N_1796);
or U2502 (N_2502,N_2131,N_1875);
nand U2503 (N_2503,N_1877,N_2035);
xor U2504 (N_2504,N_1918,N_1995);
nand U2505 (N_2505,N_2229,N_2215);
nor U2506 (N_2506,N_1547,N_2017);
and U2507 (N_2507,N_1653,N_2158);
and U2508 (N_2508,N_1734,N_1811);
and U2509 (N_2509,N_2082,N_1818);
xnor U2510 (N_2510,N_1563,N_1630);
and U2511 (N_2511,N_2084,N_1594);
nor U2512 (N_2512,N_1986,N_1860);
nand U2513 (N_2513,N_1873,N_1592);
or U2514 (N_2514,N_1715,N_2173);
or U2515 (N_2515,N_2023,N_1752);
nand U2516 (N_2516,N_2028,N_2217);
or U2517 (N_2517,N_2120,N_1581);
nor U2518 (N_2518,N_2094,N_2060);
nand U2519 (N_2519,N_1769,N_1642);
nand U2520 (N_2520,N_1975,N_1649);
and U2521 (N_2521,N_1781,N_1807);
nor U2522 (N_2522,N_1946,N_2101);
nor U2523 (N_2523,N_1690,N_1633);
nor U2524 (N_2524,N_1933,N_2024);
nand U2525 (N_2525,N_1890,N_1962);
and U2526 (N_2526,N_2166,N_1589);
nand U2527 (N_2527,N_1919,N_1620);
and U2528 (N_2528,N_1813,N_1700);
nand U2529 (N_2529,N_1565,N_1717);
nor U2530 (N_2530,N_1990,N_1906);
nand U2531 (N_2531,N_1571,N_2150);
nor U2532 (N_2532,N_1556,N_1848);
nand U2533 (N_2533,N_2078,N_2075);
and U2534 (N_2534,N_1895,N_1684);
nand U2535 (N_2535,N_2097,N_1759);
or U2536 (N_2536,N_1522,N_2153);
or U2537 (N_2537,N_1621,N_1942);
or U2538 (N_2538,N_2062,N_1757);
nor U2539 (N_2539,N_2016,N_1584);
or U2540 (N_2540,N_2228,N_1782);
and U2541 (N_2541,N_1737,N_1672);
nand U2542 (N_2542,N_1766,N_1886);
nor U2543 (N_2543,N_1834,N_1671);
nand U2544 (N_2544,N_1699,N_2108);
or U2545 (N_2545,N_1970,N_2230);
nand U2546 (N_2546,N_1940,N_1637);
nand U2547 (N_2547,N_1947,N_1861);
nor U2548 (N_2548,N_1711,N_2073);
or U2549 (N_2549,N_1998,N_1954);
or U2550 (N_2550,N_1837,N_1622);
xnor U2551 (N_2551,N_1791,N_1583);
nor U2552 (N_2552,N_2195,N_2098);
nand U2553 (N_2553,N_1510,N_1531);
or U2554 (N_2554,N_2247,N_1514);
nand U2555 (N_2555,N_2146,N_2076);
nand U2556 (N_2556,N_1889,N_2032);
and U2557 (N_2557,N_2068,N_1572);
and U2558 (N_2558,N_1507,N_2115);
or U2559 (N_2559,N_2175,N_1864);
xor U2560 (N_2560,N_1678,N_2031);
xor U2561 (N_2561,N_1644,N_1786);
and U2562 (N_2562,N_1849,N_1512);
nor U2563 (N_2563,N_1801,N_2125);
nand U2564 (N_2564,N_2142,N_1634);
xnor U2565 (N_2565,N_1966,N_2177);
nor U2566 (N_2566,N_2089,N_1871);
nand U2567 (N_2567,N_1851,N_1997);
xnor U2568 (N_2568,N_1777,N_1935);
nor U2569 (N_2569,N_2050,N_2048);
or U2570 (N_2570,N_2133,N_1891);
and U2571 (N_2571,N_1904,N_1626);
nand U2572 (N_2572,N_1896,N_1991);
and U2573 (N_2573,N_1803,N_1628);
or U2574 (N_2574,N_2143,N_2092);
and U2575 (N_2575,N_2191,N_1744);
nand U2576 (N_2576,N_2010,N_2037);
and U2577 (N_2577,N_1666,N_2227);
and U2578 (N_2578,N_1756,N_2178);
or U2579 (N_2579,N_1562,N_1593);
or U2580 (N_2580,N_1974,N_2008);
and U2581 (N_2581,N_1937,N_1738);
and U2582 (N_2582,N_1754,N_1704);
nor U2583 (N_2583,N_2182,N_1817);
nor U2584 (N_2584,N_1749,N_2045);
nand U2585 (N_2585,N_2000,N_1964);
nand U2586 (N_2586,N_1502,N_2007);
nand U2587 (N_2587,N_1945,N_2157);
nand U2588 (N_2588,N_1538,N_2100);
or U2589 (N_2589,N_1755,N_2161);
nor U2590 (N_2590,N_1732,N_2189);
nor U2591 (N_2591,N_2140,N_2049);
or U2592 (N_2592,N_2179,N_1540);
nor U2593 (N_2593,N_2159,N_1599);
and U2594 (N_2594,N_1827,N_2027);
nor U2595 (N_2595,N_2155,N_1639);
xor U2596 (N_2596,N_1980,N_2095);
or U2597 (N_2597,N_2081,N_1645);
or U2598 (N_2598,N_2122,N_2190);
nand U2599 (N_2599,N_1902,N_2193);
and U2600 (N_2600,N_1893,N_1551);
or U2601 (N_2601,N_1659,N_2106);
and U2602 (N_2602,N_1894,N_1716);
nor U2603 (N_2603,N_1802,N_1559);
and U2604 (N_2604,N_1783,N_1825);
nor U2605 (N_2605,N_1897,N_2033);
nand U2606 (N_2606,N_1691,N_1883);
nand U2607 (N_2607,N_1921,N_2123);
and U2608 (N_2608,N_1853,N_1573);
nor U2609 (N_2609,N_1784,N_2053);
nand U2610 (N_2610,N_1740,N_1809);
nor U2611 (N_2611,N_1821,N_2213);
nor U2612 (N_2612,N_2067,N_1586);
nor U2613 (N_2613,N_1605,N_1831);
or U2614 (N_2614,N_1741,N_1728);
or U2615 (N_2615,N_1958,N_1503);
and U2616 (N_2616,N_2069,N_1982);
and U2617 (N_2617,N_1567,N_1932);
or U2618 (N_2618,N_2090,N_1765);
nand U2619 (N_2619,N_2224,N_2169);
nor U2620 (N_2620,N_2129,N_2103);
or U2621 (N_2621,N_2220,N_1953);
nand U2622 (N_2622,N_2004,N_1647);
or U2623 (N_2623,N_2130,N_2121);
nor U2624 (N_2624,N_1773,N_1916);
and U2625 (N_2625,N_2112,N_1522);
and U2626 (N_2626,N_1898,N_2239);
nor U2627 (N_2627,N_1726,N_1965);
and U2628 (N_2628,N_1682,N_1608);
xor U2629 (N_2629,N_1907,N_2052);
nor U2630 (N_2630,N_2046,N_2080);
nand U2631 (N_2631,N_2101,N_1778);
nor U2632 (N_2632,N_1797,N_1881);
nand U2633 (N_2633,N_1922,N_1928);
or U2634 (N_2634,N_2177,N_1576);
and U2635 (N_2635,N_2009,N_1743);
nor U2636 (N_2636,N_1969,N_1943);
and U2637 (N_2637,N_1993,N_1740);
nand U2638 (N_2638,N_1895,N_2126);
xor U2639 (N_2639,N_2182,N_2033);
nand U2640 (N_2640,N_1658,N_1691);
nor U2641 (N_2641,N_1546,N_2152);
and U2642 (N_2642,N_2138,N_1567);
nor U2643 (N_2643,N_1678,N_1712);
nand U2644 (N_2644,N_1539,N_2056);
nand U2645 (N_2645,N_1605,N_1503);
nand U2646 (N_2646,N_2079,N_1685);
nand U2647 (N_2647,N_1516,N_1610);
nor U2648 (N_2648,N_2119,N_2059);
and U2649 (N_2649,N_1535,N_1664);
or U2650 (N_2650,N_2006,N_2100);
or U2651 (N_2651,N_1870,N_1961);
or U2652 (N_2652,N_1569,N_1680);
nand U2653 (N_2653,N_2173,N_1782);
or U2654 (N_2654,N_1526,N_1826);
nor U2655 (N_2655,N_1807,N_1932);
xor U2656 (N_2656,N_2039,N_1592);
xor U2657 (N_2657,N_1551,N_2010);
or U2658 (N_2658,N_1672,N_1581);
xor U2659 (N_2659,N_1659,N_2236);
or U2660 (N_2660,N_1590,N_1516);
or U2661 (N_2661,N_1803,N_2184);
and U2662 (N_2662,N_1664,N_2246);
and U2663 (N_2663,N_1646,N_1643);
or U2664 (N_2664,N_1823,N_1926);
nand U2665 (N_2665,N_1788,N_1508);
or U2666 (N_2666,N_1606,N_1721);
and U2667 (N_2667,N_1692,N_1619);
xnor U2668 (N_2668,N_1625,N_1860);
xnor U2669 (N_2669,N_1510,N_1596);
nor U2670 (N_2670,N_2237,N_1897);
and U2671 (N_2671,N_2157,N_1670);
nor U2672 (N_2672,N_1544,N_1590);
xnor U2673 (N_2673,N_1947,N_1968);
or U2674 (N_2674,N_1694,N_1674);
and U2675 (N_2675,N_2028,N_2125);
or U2676 (N_2676,N_1597,N_1946);
nand U2677 (N_2677,N_1565,N_1808);
xor U2678 (N_2678,N_2092,N_1963);
nand U2679 (N_2679,N_2162,N_1625);
and U2680 (N_2680,N_1537,N_2054);
and U2681 (N_2681,N_1622,N_2172);
nor U2682 (N_2682,N_2008,N_1875);
and U2683 (N_2683,N_1600,N_2153);
or U2684 (N_2684,N_1732,N_1863);
nor U2685 (N_2685,N_1508,N_1695);
nand U2686 (N_2686,N_1876,N_1758);
or U2687 (N_2687,N_2186,N_1540);
and U2688 (N_2688,N_1839,N_1624);
nor U2689 (N_2689,N_1747,N_1723);
and U2690 (N_2690,N_1564,N_2046);
nand U2691 (N_2691,N_1700,N_1933);
nor U2692 (N_2692,N_2047,N_1650);
or U2693 (N_2693,N_1883,N_1831);
or U2694 (N_2694,N_2208,N_1858);
nand U2695 (N_2695,N_2172,N_1626);
nor U2696 (N_2696,N_2070,N_1907);
xor U2697 (N_2697,N_1798,N_2132);
or U2698 (N_2698,N_1666,N_2118);
nor U2699 (N_2699,N_1790,N_1518);
or U2700 (N_2700,N_1583,N_1692);
nor U2701 (N_2701,N_2019,N_2046);
nand U2702 (N_2702,N_1588,N_2219);
nand U2703 (N_2703,N_1711,N_1719);
or U2704 (N_2704,N_2240,N_1543);
and U2705 (N_2705,N_1741,N_1742);
xor U2706 (N_2706,N_2154,N_1990);
or U2707 (N_2707,N_1730,N_1959);
nor U2708 (N_2708,N_2038,N_1719);
nand U2709 (N_2709,N_1838,N_2202);
or U2710 (N_2710,N_2178,N_1616);
nor U2711 (N_2711,N_1505,N_1969);
and U2712 (N_2712,N_1979,N_1830);
and U2713 (N_2713,N_1790,N_1516);
or U2714 (N_2714,N_1528,N_1882);
nand U2715 (N_2715,N_2060,N_2246);
or U2716 (N_2716,N_1779,N_1815);
xor U2717 (N_2717,N_1962,N_2222);
and U2718 (N_2718,N_1655,N_1765);
nand U2719 (N_2719,N_1576,N_2178);
nand U2720 (N_2720,N_1681,N_2082);
nand U2721 (N_2721,N_1923,N_1555);
xor U2722 (N_2722,N_2174,N_2236);
nand U2723 (N_2723,N_2111,N_1899);
nor U2724 (N_2724,N_1756,N_1796);
xnor U2725 (N_2725,N_1559,N_1570);
nor U2726 (N_2726,N_2096,N_2073);
nand U2727 (N_2727,N_1667,N_1810);
or U2728 (N_2728,N_1611,N_1589);
xnor U2729 (N_2729,N_1563,N_1561);
xor U2730 (N_2730,N_2045,N_1660);
and U2731 (N_2731,N_1547,N_1766);
nand U2732 (N_2732,N_1879,N_1641);
and U2733 (N_2733,N_1533,N_1846);
nor U2734 (N_2734,N_1580,N_2161);
nor U2735 (N_2735,N_2145,N_1689);
nor U2736 (N_2736,N_2244,N_2088);
or U2737 (N_2737,N_1825,N_2057);
and U2738 (N_2738,N_1762,N_1547);
and U2739 (N_2739,N_2160,N_1875);
nor U2740 (N_2740,N_2107,N_1996);
nand U2741 (N_2741,N_2039,N_1907);
nand U2742 (N_2742,N_1710,N_1634);
nor U2743 (N_2743,N_1620,N_2104);
nor U2744 (N_2744,N_1859,N_1839);
or U2745 (N_2745,N_1624,N_1846);
nand U2746 (N_2746,N_2029,N_2231);
xnor U2747 (N_2747,N_1802,N_1832);
and U2748 (N_2748,N_1725,N_1656);
or U2749 (N_2749,N_1520,N_2148);
or U2750 (N_2750,N_2167,N_2126);
nand U2751 (N_2751,N_2079,N_1895);
nand U2752 (N_2752,N_1626,N_1680);
xor U2753 (N_2753,N_1702,N_1868);
nand U2754 (N_2754,N_1539,N_1639);
or U2755 (N_2755,N_1906,N_1709);
and U2756 (N_2756,N_2160,N_1933);
xor U2757 (N_2757,N_1930,N_2085);
nor U2758 (N_2758,N_2098,N_2016);
and U2759 (N_2759,N_2032,N_1967);
nor U2760 (N_2760,N_1558,N_2179);
xnor U2761 (N_2761,N_2073,N_2118);
or U2762 (N_2762,N_1897,N_2209);
or U2763 (N_2763,N_2090,N_2002);
nand U2764 (N_2764,N_2057,N_2177);
or U2765 (N_2765,N_1946,N_1889);
or U2766 (N_2766,N_1971,N_1767);
nand U2767 (N_2767,N_2025,N_1767);
and U2768 (N_2768,N_1697,N_2225);
or U2769 (N_2769,N_1581,N_1579);
or U2770 (N_2770,N_1852,N_1879);
nor U2771 (N_2771,N_1665,N_1611);
and U2772 (N_2772,N_1690,N_1838);
and U2773 (N_2773,N_1926,N_1542);
nand U2774 (N_2774,N_1730,N_1527);
and U2775 (N_2775,N_1662,N_1695);
nand U2776 (N_2776,N_1611,N_1947);
xnor U2777 (N_2777,N_1504,N_1554);
and U2778 (N_2778,N_1995,N_2192);
and U2779 (N_2779,N_1605,N_1864);
nor U2780 (N_2780,N_1947,N_1928);
and U2781 (N_2781,N_1928,N_1509);
xor U2782 (N_2782,N_2024,N_1599);
nand U2783 (N_2783,N_1685,N_1787);
or U2784 (N_2784,N_1787,N_2009);
nand U2785 (N_2785,N_1632,N_1508);
or U2786 (N_2786,N_2114,N_2226);
or U2787 (N_2787,N_1856,N_2076);
or U2788 (N_2788,N_1655,N_2089);
nor U2789 (N_2789,N_2127,N_1589);
and U2790 (N_2790,N_1930,N_2102);
and U2791 (N_2791,N_1656,N_1880);
or U2792 (N_2792,N_2180,N_1913);
nor U2793 (N_2793,N_2223,N_1570);
or U2794 (N_2794,N_1640,N_1834);
xnor U2795 (N_2795,N_2031,N_1706);
nor U2796 (N_2796,N_1604,N_1918);
nor U2797 (N_2797,N_1939,N_2173);
or U2798 (N_2798,N_2095,N_1907);
and U2799 (N_2799,N_1728,N_1915);
and U2800 (N_2800,N_1528,N_2196);
nor U2801 (N_2801,N_1693,N_2088);
nand U2802 (N_2802,N_2018,N_2094);
nor U2803 (N_2803,N_2222,N_2011);
nor U2804 (N_2804,N_2090,N_1686);
and U2805 (N_2805,N_1787,N_2086);
nor U2806 (N_2806,N_1837,N_1756);
xnor U2807 (N_2807,N_2188,N_1988);
nor U2808 (N_2808,N_1983,N_1878);
and U2809 (N_2809,N_2138,N_1742);
and U2810 (N_2810,N_2247,N_1530);
nand U2811 (N_2811,N_2222,N_1822);
nor U2812 (N_2812,N_1742,N_1966);
or U2813 (N_2813,N_1606,N_2235);
nand U2814 (N_2814,N_2222,N_1846);
and U2815 (N_2815,N_1922,N_1802);
nor U2816 (N_2816,N_2227,N_2156);
and U2817 (N_2817,N_1807,N_1976);
and U2818 (N_2818,N_1593,N_1551);
or U2819 (N_2819,N_2236,N_2233);
or U2820 (N_2820,N_1914,N_2178);
or U2821 (N_2821,N_1546,N_1826);
nor U2822 (N_2822,N_2110,N_1684);
and U2823 (N_2823,N_1635,N_1934);
or U2824 (N_2824,N_1697,N_2054);
nand U2825 (N_2825,N_2193,N_2187);
or U2826 (N_2826,N_2172,N_2173);
nor U2827 (N_2827,N_1800,N_1820);
or U2828 (N_2828,N_2075,N_1586);
or U2829 (N_2829,N_1824,N_1525);
xnor U2830 (N_2830,N_2109,N_2143);
nor U2831 (N_2831,N_1780,N_2154);
nand U2832 (N_2832,N_2174,N_2224);
or U2833 (N_2833,N_2154,N_1889);
nor U2834 (N_2834,N_1863,N_1799);
or U2835 (N_2835,N_2115,N_2103);
xor U2836 (N_2836,N_1707,N_1766);
or U2837 (N_2837,N_1979,N_1771);
nand U2838 (N_2838,N_2242,N_1729);
and U2839 (N_2839,N_1529,N_2130);
and U2840 (N_2840,N_2005,N_2038);
nor U2841 (N_2841,N_2017,N_2211);
nand U2842 (N_2842,N_1726,N_1810);
nand U2843 (N_2843,N_1830,N_2003);
nand U2844 (N_2844,N_1606,N_1960);
and U2845 (N_2845,N_1652,N_1851);
or U2846 (N_2846,N_2075,N_1957);
or U2847 (N_2847,N_2172,N_1521);
nand U2848 (N_2848,N_2239,N_2051);
xnor U2849 (N_2849,N_1586,N_1510);
xnor U2850 (N_2850,N_1999,N_2226);
or U2851 (N_2851,N_2181,N_1594);
and U2852 (N_2852,N_1788,N_2175);
nand U2853 (N_2853,N_1902,N_1522);
and U2854 (N_2854,N_1630,N_2058);
xor U2855 (N_2855,N_1964,N_2159);
nand U2856 (N_2856,N_1882,N_1856);
and U2857 (N_2857,N_1890,N_2149);
nand U2858 (N_2858,N_2058,N_1947);
and U2859 (N_2859,N_2050,N_1633);
and U2860 (N_2860,N_2072,N_1891);
nor U2861 (N_2861,N_2225,N_1516);
or U2862 (N_2862,N_1633,N_2063);
or U2863 (N_2863,N_1857,N_1704);
nor U2864 (N_2864,N_1526,N_2101);
nand U2865 (N_2865,N_1746,N_2068);
or U2866 (N_2866,N_1916,N_1717);
nand U2867 (N_2867,N_1947,N_1723);
xnor U2868 (N_2868,N_2123,N_1591);
or U2869 (N_2869,N_2216,N_2228);
or U2870 (N_2870,N_1924,N_1783);
and U2871 (N_2871,N_1585,N_2103);
nand U2872 (N_2872,N_1617,N_1794);
nand U2873 (N_2873,N_2236,N_1993);
nor U2874 (N_2874,N_1719,N_1805);
xnor U2875 (N_2875,N_1957,N_1919);
xnor U2876 (N_2876,N_2063,N_1712);
xnor U2877 (N_2877,N_1968,N_2029);
and U2878 (N_2878,N_2130,N_1936);
or U2879 (N_2879,N_2091,N_1878);
xor U2880 (N_2880,N_1988,N_1525);
nand U2881 (N_2881,N_1699,N_1822);
and U2882 (N_2882,N_2052,N_2176);
and U2883 (N_2883,N_1518,N_1838);
or U2884 (N_2884,N_1888,N_1986);
or U2885 (N_2885,N_2148,N_1905);
nand U2886 (N_2886,N_2146,N_1722);
nor U2887 (N_2887,N_2140,N_1793);
nor U2888 (N_2888,N_1829,N_1607);
nor U2889 (N_2889,N_2074,N_1981);
xor U2890 (N_2890,N_1875,N_1589);
nor U2891 (N_2891,N_2081,N_1794);
nand U2892 (N_2892,N_1800,N_2119);
or U2893 (N_2893,N_1937,N_2053);
nor U2894 (N_2894,N_2237,N_2071);
and U2895 (N_2895,N_1657,N_2090);
nor U2896 (N_2896,N_1606,N_2188);
xnor U2897 (N_2897,N_1601,N_1683);
nor U2898 (N_2898,N_2195,N_2024);
and U2899 (N_2899,N_1782,N_2207);
and U2900 (N_2900,N_1819,N_1988);
nand U2901 (N_2901,N_2054,N_1713);
nor U2902 (N_2902,N_1644,N_2160);
nor U2903 (N_2903,N_1761,N_2134);
or U2904 (N_2904,N_2066,N_1876);
and U2905 (N_2905,N_1905,N_1685);
nand U2906 (N_2906,N_2152,N_1659);
or U2907 (N_2907,N_1836,N_1568);
nand U2908 (N_2908,N_1591,N_1681);
or U2909 (N_2909,N_1799,N_2165);
or U2910 (N_2910,N_1587,N_1799);
and U2911 (N_2911,N_1794,N_1594);
and U2912 (N_2912,N_1683,N_2178);
xnor U2913 (N_2913,N_2235,N_1756);
nand U2914 (N_2914,N_1743,N_1517);
or U2915 (N_2915,N_2079,N_2197);
nor U2916 (N_2916,N_1992,N_1897);
and U2917 (N_2917,N_1813,N_2001);
or U2918 (N_2918,N_2051,N_1662);
and U2919 (N_2919,N_1987,N_1964);
nand U2920 (N_2920,N_1588,N_2121);
nor U2921 (N_2921,N_2041,N_2244);
and U2922 (N_2922,N_2200,N_1776);
and U2923 (N_2923,N_2202,N_1977);
nor U2924 (N_2924,N_2168,N_2151);
nand U2925 (N_2925,N_2031,N_1680);
and U2926 (N_2926,N_1752,N_1703);
and U2927 (N_2927,N_2084,N_1961);
xnor U2928 (N_2928,N_2158,N_1558);
nand U2929 (N_2929,N_2234,N_1735);
xnor U2930 (N_2930,N_1955,N_2015);
or U2931 (N_2931,N_1952,N_2231);
and U2932 (N_2932,N_1799,N_1699);
xor U2933 (N_2933,N_1599,N_1742);
nand U2934 (N_2934,N_2147,N_1977);
nand U2935 (N_2935,N_1738,N_1859);
nor U2936 (N_2936,N_1682,N_1523);
and U2937 (N_2937,N_1979,N_1793);
nand U2938 (N_2938,N_2154,N_1758);
nand U2939 (N_2939,N_1623,N_1791);
nand U2940 (N_2940,N_2045,N_1612);
nor U2941 (N_2941,N_1561,N_2240);
or U2942 (N_2942,N_1935,N_1583);
nor U2943 (N_2943,N_1847,N_1850);
and U2944 (N_2944,N_1924,N_2088);
or U2945 (N_2945,N_1691,N_1900);
nand U2946 (N_2946,N_1782,N_2054);
and U2947 (N_2947,N_2189,N_2165);
and U2948 (N_2948,N_2119,N_1865);
xor U2949 (N_2949,N_2170,N_2129);
and U2950 (N_2950,N_1845,N_1507);
and U2951 (N_2951,N_2166,N_2109);
nor U2952 (N_2952,N_2097,N_2212);
and U2953 (N_2953,N_1802,N_1745);
nor U2954 (N_2954,N_1690,N_1823);
nor U2955 (N_2955,N_2085,N_1617);
or U2956 (N_2956,N_2098,N_1818);
and U2957 (N_2957,N_1579,N_1951);
nand U2958 (N_2958,N_2005,N_1518);
nand U2959 (N_2959,N_1713,N_1869);
nor U2960 (N_2960,N_1780,N_1687);
xnor U2961 (N_2961,N_1722,N_1885);
nand U2962 (N_2962,N_2162,N_1767);
and U2963 (N_2963,N_1533,N_1575);
nand U2964 (N_2964,N_2008,N_2057);
nor U2965 (N_2965,N_1910,N_1515);
nor U2966 (N_2966,N_1672,N_2158);
nor U2967 (N_2967,N_1617,N_1686);
nor U2968 (N_2968,N_1876,N_1968);
and U2969 (N_2969,N_1532,N_2088);
and U2970 (N_2970,N_1552,N_2151);
nor U2971 (N_2971,N_1928,N_2106);
xnor U2972 (N_2972,N_1609,N_2186);
or U2973 (N_2973,N_1994,N_2187);
nand U2974 (N_2974,N_1816,N_2095);
nor U2975 (N_2975,N_2059,N_1823);
nand U2976 (N_2976,N_2083,N_2097);
or U2977 (N_2977,N_1545,N_1768);
and U2978 (N_2978,N_1954,N_1874);
nor U2979 (N_2979,N_1861,N_2036);
nor U2980 (N_2980,N_2097,N_1932);
nand U2981 (N_2981,N_1654,N_2244);
and U2982 (N_2982,N_1605,N_1916);
and U2983 (N_2983,N_2032,N_1839);
and U2984 (N_2984,N_1863,N_1970);
nand U2985 (N_2985,N_1915,N_1662);
and U2986 (N_2986,N_1669,N_1959);
and U2987 (N_2987,N_1793,N_2173);
xnor U2988 (N_2988,N_1867,N_2086);
and U2989 (N_2989,N_1822,N_1926);
and U2990 (N_2990,N_1644,N_1897);
nor U2991 (N_2991,N_1585,N_2071);
nand U2992 (N_2992,N_1506,N_1963);
nor U2993 (N_2993,N_2004,N_2229);
nand U2994 (N_2994,N_1561,N_1927);
nor U2995 (N_2995,N_1683,N_1725);
and U2996 (N_2996,N_2044,N_2027);
nor U2997 (N_2997,N_1631,N_1655);
nor U2998 (N_2998,N_2171,N_2166);
or U2999 (N_2999,N_2155,N_1537);
xor U3000 (N_3000,N_2435,N_2276);
and U3001 (N_3001,N_2286,N_2260);
nor U3002 (N_3002,N_2253,N_2592);
nor U3003 (N_3003,N_2828,N_2759);
and U3004 (N_3004,N_2375,N_2660);
and U3005 (N_3005,N_2876,N_2443);
nand U3006 (N_3006,N_2781,N_2704);
nor U3007 (N_3007,N_2820,N_2722);
nand U3008 (N_3008,N_2743,N_2401);
and U3009 (N_3009,N_2431,N_2910);
nor U3010 (N_3010,N_2937,N_2279);
and U3011 (N_3011,N_2292,N_2537);
and U3012 (N_3012,N_2985,N_2527);
and U3013 (N_3013,N_2508,N_2888);
or U3014 (N_3014,N_2884,N_2933);
and U3015 (N_3015,N_2418,N_2275);
nor U3016 (N_3016,N_2540,N_2447);
or U3017 (N_3017,N_2277,N_2922);
and U3018 (N_3018,N_2670,N_2434);
or U3019 (N_3019,N_2555,N_2671);
or U3020 (N_3020,N_2998,N_2804);
and U3021 (N_3021,N_2851,N_2341);
and U3022 (N_3022,N_2990,N_2510);
or U3023 (N_3023,N_2261,N_2257);
and U3024 (N_3024,N_2674,N_2805);
and U3025 (N_3025,N_2595,N_2870);
xnor U3026 (N_3026,N_2615,N_2931);
xnor U3027 (N_3027,N_2977,N_2713);
nand U3028 (N_3028,N_2691,N_2474);
and U3029 (N_3029,N_2387,N_2879);
xor U3030 (N_3030,N_2652,N_2733);
xor U3031 (N_3031,N_2865,N_2969);
xnor U3032 (N_3032,N_2367,N_2424);
xor U3033 (N_3033,N_2947,N_2782);
nor U3034 (N_3034,N_2923,N_2329);
nand U3035 (N_3035,N_2873,N_2886);
nor U3036 (N_3036,N_2308,N_2471);
or U3037 (N_3037,N_2402,N_2815);
or U3038 (N_3038,N_2384,N_2525);
xor U3039 (N_3039,N_2609,N_2706);
nand U3040 (N_3040,N_2498,N_2496);
nand U3041 (N_3041,N_2533,N_2897);
and U3042 (N_3042,N_2399,N_2940);
nor U3043 (N_3043,N_2572,N_2895);
and U3044 (N_3044,N_2280,N_2548);
nand U3045 (N_3045,N_2889,N_2757);
xor U3046 (N_3046,N_2874,N_2446);
nand U3047 (N_3047,N_2607,N_2916);
or U3048 (N_3048,N_2349,N_2868);
or U3049 (N_3049,N_2893,N_2974);
or U3050 (N_3050,N_2610,N_2547);
or U3051 (N_3051,N_2846,N_2817);
and U3052 (N_3052,N_2368,N_2386);
or U3053 (N_3053,N_2528,N_2475);
or U3054 (N_3054,N_2681,N_2742);
xor U3055 (N_3055,N_2457,N_2371);
nor U3056 (N_3056,N_2352,N_2642);
xnor U3057 (N_3057,N_2444,N_2307);
or U3058 (N_3058,N_2948,N_2398);
or U3059 (N_3059,N_2882,N_2505);
nor U3060 (N_3060,N_2839,N_2849);
nor U3061 (N_3061,N_2754,N_2677);
nand U3062 (N_3062,N_2536,N_2776);
or U3063 (N_3063,N_2383,N_2966);
and U3064 (N_3064,N_2685,N_2799);
or U3065 (N_3065,N_2669,N_2313);
and U3066 (N_3066,N_2545,N_2321);
nand U3067 (N_3067,N_2661,N_2679);
and U3068 (N_3068,N_2918,N_2506);
and U3069 (N_3069,N_2303,N_2975);
and U3070 (N_3070,N_2943,N_2487);
nor U3071 (N_3071,N_2370,N_2877);
or U3072 (N_3072,N_2278,N_2580);
and U3073 (N_3073,N_2428,N_2574);
xor U3074 (N_3074,N_2252,N_2905);
nand U3075 (N_3075,N_2831,N_2852);
nand U3076 (N_3076,N_2911,N_2251);
nand U3077 (N_3077,N_2978,N_2739);
or U3078 (N_3078,N_2939,N_2550);
nor U3079 (N_3079,N_2779,N_2919);
xnor U3080 (N_3080,N_2684,N_2265);
or U3081 (N_3081,N_2354,N_2535);
or U3082 (N_3082,N_2576,N_2394);
nor U3083 (N_3083,N_2793,N_2456);
or U3084 (N_3084,N_2857,N_2283);
and U3085 (N_3085,N_2591,N_2847);
or U3086 (N_3086,N_2564,N_2494);
nor U3087 (N_3087,N_2723,N_2451);
nor U3088 (N_3088,N_2357,N_2628);
xnor U3089 (N_3089,N_2858,N_2914);
nand U3090 (N_3090,N_2390,N_2732);
and U3091 (N_3091,N_2797,N_2983);
xor U3092 (N_3092,N_2599,N_2833);
and U3093 (N_3093,N_2319,N_2369);
nor U3094 (N_3094,N_2439,N_2478);
xnor U3095 (N_3095,N_2604,N_2921);
xnor U3096 (N_3096,N_2827,N_2663);
or U3097 (N_3097,N_2499,N_2624);
nand U3098 (N_3098,N_2822,N_2302);
nor U3099 (N_3099,N_2710,N_2415);
nor U3100 (N_3100,N_2400,N_2635);
xnor U3101 (N_3101,N_2850,N_2616);
xor U3102 (N_3102,N_2698,N_2790);
and U3103 (N_3103,N_2638,N_2598);
or U3104 (N_3104,N_2271,N_2339);
nor U3105 (N_3105,N_2825,N_2342);
or U3106 (N_3106,N_2760,N_2282);
or U3107 (N_3107,N_2483,N_2539);
and U3108 (N_3108,N_2666,N_2389);
or U3109 (N_3109,N_2938,N_2455);
nor U3110 (N_3110,N_2795,N_2769);
and U3111 (N_3111,N_2408,N_2715);
and U3112 (N_3112,N_2468,N_2584);
nor U3113 (N_3113,N_2423,N_2274);
xor U3114 (N_3114,N_2786,N_2619);
or U3115 (N_3115,N_2951,N_2526);
nor U3116 (N_3116,N_2509,N_2438);
nor U3117 (N_3117,N_2792,N_2737);
or U3118 (N_3118,N_2587,N_2672);
or U3119 (N_3119,N_2814,N_2461);
or U3120 (N_3120,N_2263,N_2345);
xor U3121 (N_3121,N_2773,N_2767);
xnor U3122 (N_3122,N_2891,N_2860);
and U3123 (N_3123,N_2343,N_2801);
nor U3124 (N_3124,N_2785,N_2589);
nand U3125 (N_3125,N_2716,N_2409);
nand U3126 (N_3126,N_2269,N_2359);
and U3127 (N_3127,N_2960,N_2695);
nand U3128 (N_3128,N_2270,N_2824);
and U3129 (N_3129,N_2517,N_2264);
and U3130 (N_3130,N_2521,N_2777);
nor U3131 (N_3131,N_2429,N_2898);
and U3132 (N_3132,N_2440,N_2724);
or U3133 (N_3133,N_2560,N_2376);
or U3134 (N_3134,N_2305,N_2378);
xor U3135 (N_3135,N_2775,N_2950);
nand U3136 (N_3136,N_2899,N_2262);
or U3137 (N_3137,N_2417,N_2411);
or U3138 (N_3138,N_2310,N_2772);
and U3139 (N_3139,N_2784,N_2738);
nand U3140 (N_3140,N_2946,N_2744);
or U3141 (N_3141,N_2291,N_2464);
nand U3142 (N_3142,N_2558,N_2862);
and U3143 (N_3143,N_2331,N_2800);
nand U3144 (N_3144,N_2553,N_2749);
nor U3145 (N_3145,N_2575,N_2682);
nor U3146 (N_3146,N_2594,N_2668);
and U3147 (N_3147,N_2425,N_2323);
nor U3148 (N_3148,N_2747,N_2542);
nand U3149 (N_3149,N_2436,N_2374);
or U3150 (N_3150,N_2845,N_2796);
or U3151 (N_3151,N_2708,N_2654);
or U3152 (N_3152,N_2266,N_2963);
xor U3153 (N_3153,N_2885,N_2485);
nor U3154 (N_3154,N_2569,N_2318);
nor U3155 (N_3155,N_2258,N_2567);
and U3156 (N_3156,N_2309,N_2643);
nand U3157 (N_3157,N_2437,N_2837);
or U3158 (N_3158,N_2541,N_2872);
nor U3159 (N_3159,N_2578,N_2690);
or U3160 (N_3160,N_2452,N_2731);
or U3161 (N_3161,N_2534,N_2328);
or U3162 (N_3162,N_2285,N_2930);
and U3163 (N_3163,N_2491,N_2381);
and U3164 (N_3164,N_2788,N_2887);
or U3165 (N_3165,N_2503,N_2577);
nand U3166 (N_3166,N_2991,N_2693);
or U3167 (N_3167,N_2518,N_2844);
or U3168 (N_3168,N_2377,N_2655);
or U3169 (N_3169,N_2808,N_2848);
xor U3170 (N_3170,N_2284,N_2497);
or U3171 (N_3171,N_2942,N_2433);
nor U3172 (N_3172,N_2763,N_2701);
nand U3173 (N_3173,N_2875,N_2894);
xnor U3174 (N_3174,N_2997,N_2549);
nor U3175 (N_3175,N_2579,N_2636);
or U3176 (N_3176,N_2964,N_2976);
or U3177 (N_3177,N_2501,N_2806);
and U3178 (N_3178,N_2250,N_2970);
and U3179 (N_3179,N_2489,N_2741);
or U3180 (N_3180,N_2372,N_2720);
xor U3181 (N_3181,N_2519,N_2495);
nand U3182 (N_3182,N_2430,N_2532);
or U3183 (N_3183,N_2856,N_2734);
nand U3184 (N_3184,N_2602,N_2397);
xnor U3185 (N_3185,N_2935,N_2687);
and U3186 (N_3186,N_2699,N_2335);
or U3187 (N_3187,N_2707,N_2571);
nand U3188 (N_3188,N_2295,N_2422);
and U3189 (N_3189,N_2753,N_2356);
and U3190 (N_3190,N_2593,N_2662);
nor U3191 (N_3191,N_2794,N_2611);
or U3192 (N_3192,N_2962,N_2696);
nor U3193 (N_3193,N_2648,N_2994);
or U3194 (N_3194,N_2714,N_2813);
nand U3195 (N_3195,N_2630,N_2396);
nor U3196 (N_3196,N_2458,N_2787);
nor U3197 (N_3197,N_2675,N_2954);
or U3198 (N_3198,N_2807,N_2373);
nand U3199 (N_3199,N_2419,N_2859);
nor U3200 (N_3200,N_2765,N_2348);
nand U3201 (N_3201,N_2421,N_2450);
nand U3202 (N_3202,N_2426,N_2256);
and U3203 (N_3203,N_2896,N_2543);
nand U3204 (N_3204,N_2297,N_2758);
nor U3205 (N_3205,N_2404,N_2347);
or U3206 (N_3206,N_2512,N_2255);
and U3207 (N_3207,N_2608,N_2290);
nor U3208 (N_3208,N_2941,N_2816);
and U3209 (N_3209,N_2486,N_2826);
nand U3210 (N_3210,N_2267,N_2834);
or U3211 (N_3211,N_2296,N_2606);
nor U3212 (N_3212,N_2883,N_2633);
and U3213 (N_3213,N_2866,N_2388);
and U3214 (N_3214,N_2466,N_2774);
nor U3215 (N_3215,N_2293,N_2700);
nor U3216 (N_3216,N_2326,N_2351);
nand U3217 (N_3217,N_2459,N_2620);
and U3218 (N_3218,N_2391,N_2557);
and U3219 (N_3219,N_2530,N_2363);
nand U3220 (N_3220,N_2320,N_2554);
xor U3221 (N_3221,N_2987,N_2973);
or U3222 (N_3222,N_2959,N_2465);
or U3223 (N_3223,N_2561,N_2344);
xnor U3224 (N_3224,N_2861,N_2304);
nand U3225 (N_3225,N_2928,N_2657);
and U3226 (N_3226,N_2603,N_2745);
nand U3227 (N_3227,N_2631,N_2812);
nor U3228 (N_3228,N_2819,N_2287);
nor U3229 (N_3229,N_2427,N_2651);
xnor U3230 (N_3230,N_2625,N_2453);
nand U3231 (N_3231,N_2626,N_2366);
and U3232 (N_3232,N_2965,N_2322);
and U3233 (N_3233,N_2712,N_2726);
nor U3234 (N_3234,N_2702,N_2867);
xor U3235 (N_3235,N_2317,N_2907);
nand U3236 (N_3236,N_2717,N_2986);
xnor U3237 (N_3237,N_2993,N_2617);
and U3238 (N_3238,N_2568,N_2337);
xor U3239 (N_3239,N_2334,N_2306);
or U3240 (N_3240,N_2413,N_2614);
and U3241 (N_3241,N_2538,N_2613);
and U3242 (N_3242,N_2904,N_2688);
nor U3243 (N_3243,N_2768,N_2841);
nor U3244 (N_3244,N_2830,N_2705);
nor U3245 (N_3245,N_2752,N_2332);
xor U3246 (N_3246,N_2730,N_2551);
or U3247 (N_3247,N_2906,N_2477);
nand U3248 (N_3248,N_2778,N_2355);
and U3249 (N_3249,N_2721,N_2469);
or U3250 (N_3250,N_2925,N_2880);
nand U3251 (N_3251,N_2522,N_2482);
nor U3252 (N_3252,N_2920,N_2504);
xnor U3253 (N_3253,N_2544,N_2407);
and U3254 (N_3254,N_2520,N_2600);
and U3255 (N_3255,N_2746,N_2460);
or U3256 (N_3256,N_2798,N_2448);
nand U3257 (N_3257,N_2559,N_2936);
and U3258 (N_3258,N_2766,N_2639);
nand U3259 (N_3259,N_2750,N_2573);
nor U3260 (N_3260,N_2420,N_2392);
nand U3261 (N_3261,N_2955,N_2902);
nor U3262 (N_3262,N_2529,N_2629);
xnor U3263 (N_3263,N_2676,N_2982);
xor U3264 (N_3264,N_2944,N_2338);
or U3265 (N_3265,N_2298,N_2645);
and U3266 (N_3266,N_2472,N_2324);
or U3267 (N_3267,N_2484,N_2811);
or U3268 (N_3268,N_2909,N_2838);
nand U3269 (N_3269,N_2912,N_2783);
nand U3270 (N_3270,N_2984,N_2272);
nand U3271 (N_3271,N_2288,N_2729);
and U3272 (N_3272,N_2949,N_2890);
nor U3273 (N_3273,N_2727,N_2597);
and U3274 (N_3274,N_2956,N_2913);
and U3275 (N_3275,N_2596,N_2618);
nor U3276 (N_3276,N_2649,N_2479);
and U3277 (N_3277,N_2694,N_2647);
and U3278 (N_3278,N_2552,N_2582);
nand U3279 (N_3279,N_2988,N_2268);
or U3280 (N_3280,N_2980,N_2315);
or U3281 (N_3281,N_2382,N_2449);
nand U3282 (N_3282,N_2958,N_2473);
and U3283 (N_3283,N_2273,N_2903);
and U3284 (N_3284,N_2832,N_2562);
or U3285 (N_3285,N_2523,N_2673);
nand U3286 (N_3286,N_2842,N_2823);
xnor U3287 (N_3287,N_2294,N_2658);
nand U3288 (N_3288,N_2565,N_2835);
and U3289 (N_3289,N_2590,N_2327);
nand U3290 (N_3290,N_2771,N_2581);
or U3291 (N_3291,N_2454,N_2659);
or U3292 (N_3292,N_2992,N_2863);
and U3293 (N_3293,N_2379,N_2968);
nor U3294 (N_3294,N_2755,N_2864);
nor U3295 (N_3295,N_2445,N_2364);
or U3296 (N_3296,N_2644,N_2653);
nor U3297 (N_3297,N_2637,N_2299);
nor U3298 (N_3298,N_2952,N_2840);
and U3299 (N_3299,N_2476,N_2995);
xor U3300 (N_3300,N_2515,N_2843);
nor U3301 (N_3301,N_2634,N_2583);
and U3302 (N_3302,N_2601,N_2300);
nor U3303 (N_3303,N_2709,N_2281);
nor U3304 (N_3304,N_2829,N_2605);
nand U3305 (N_3305,N_2650,N_2362);
and U3306 (N_3306,N_2513,N_2488);
and U3307 (N_3307,N_2623,N_2405);
or U3308 (N_3308,N_2360,N_2441);
nor U3309 (N_3309,N_2927,N_2719);
or U3310 (N_3310,N_2566,N_2683);
nand U3311 (N_3311,N_2810,N_2802);
or U3312 (N_3312,N_2563,N_2470);
nor U3313 (N_3313,N_2725,N_2770);
nor U3314 (N_3314,N_2361,N_2346);
nand U3315 (N_3315,N_2393,N_2735);
nand U3316 (N_3316,N_2929,N_2981);
nand U3317 (N_3317,N_2908,N_2414);
or U3318 (N_3318,N_2878,N_2301);
xor U3319 (N_3319,N_2312,N_2989);
or U3320 (N_3320,N_2869,N_2646);
xnor U3321 (N_3321,N_2588,N_2395);
or U3322 (N_3322,N_2803,N_2791);
or U3323 (N_3323,N_2748,N_2336);
nor U3324 (N_3324,N_2442,N_2403);
or U3325 (N_3325,N_2546,N_2761);
nor U3326 (N_3326,N_2586,N_2632);
nor U3327 (N_3327,N_2689,N_2531);
nor U3328 (N_3328,N_2330,N_2502);
xor U3329 (N_3329,N_2756,N_2740);
nand U3330 (N_3330,N_2703,N_2917);
or U3331 (N_3331,N_2492,N_2915);
nor U3332 (N_3332,N_2480,N_2736);
nor U3333 (N_3333,N_2340,N_2358);
nor U3334 (N_3334,N_2640,N_2680);
and U3335 (N_3335,N_2353,N_2789);
and U3336 (N_3336,N_2979,N_2516);
and U3337 (N_3337,N_2612,N_2892);
or U3338 (N_3338,N_2945,N_2934);
xor U3339 (N_3339,N_2900,N_2627);
nor U3340 (N_3340,N_2971,N_2762);
nand U3341 (N_3341,N_2621,N_2678);
xor U3342 (N_3342,N_2416,N_2809);
nor U3343 (N_3343,N_2500,N_2728);
xnor U3344 (N_3344,N_2664,N_2467);
or U3345 (N_3345,N_2380,N_2961);
nor U3346 (N_3346,N_2697,N_2507);
and U3347 (N_3347,N_2692,N_2524);
nor U3348 (N_3348,N_2924,N_2259);
and U3349 (N_3349,N_2972,N_2311);
nor U3350 (N_3350,N_2622,N_2490);
nand U3351 (N_3351,N_2350,N_2412);
nand U3352 (N_3352,N_2932,N_2325);
nand U3353 (N_3353,N_2406,N_2316);
nor U3354 (N_3354,N_2901,N_2254);
xnor U3355 (N_3355,N_2854,N_2855);
nand U3356 (N_3356,N_2718,N_2641);
and U3357 (N_3357,N_2289,N_2665);
or U3358 (N_3358,N_2365,N_2711);
nor U3359 (N_3359,N_2493,N_2656);
and U3360 (N_3360,N_2996,N_2953);
or U3361 (N_3361,N_2585,N_2333);
xnor U3362 (N_3362,N_2967,N_2511);
nor U3363 (N_3363,N_2556,N_2514);
and U3364 (N_3364,N_2780,N_2686);
nor U3365 (N_3365,N_2410,N_2462);
nand U3366 (N_3366,N_2764,N_2463);
nand U3367 (N_3367,N_2821,N_2881);
nand U3368 (N_3368,N_2481,N_2999);
xnor U3369 (N_3369,N_2667,N_2432);
and U3370 (N_3370,N_2853,N_2314);
nor U3371 (N_3371,N_2570,N_2385);
nor U3372 (N_3372,N_2751,N_2957);
xor U3373 (N_3373,N_2818,N_2926);
or U3374 (N_3374,N_2836,N_2871);
and U3375 (N_3375,N_2983,N_2612);
nand U3376 (N_3376,N_2604,N_2274);
and U3377 (N_3377,N_2629,N_2333);
and U3378 (N_3378,N_2765,N_2971);
and U3379 (N_3379,N_2733,N_2280);
and U3380 (N_3380,N_2679,N_2493);
or U3381 (N_3381,N_2447,N_2877);
nor U3382 (N_3382,N_2873,N_2803);
and U3383 (N_3383,N_2471,N_2429);
nor U3384 (N_3384,N_2636,N_2368);
or U3385 (N_3385,N_2676,N_2330);
nor U3386 (N_3386,N_2722,N_2801);
xor U3387 (N_3387,N_2778,N_2558);
nor U3388 (N_3388,N_2968,N_2797);
nor U3389 (N_3389,N_2731,N_2455);
and U3390 (N_3390,N_2269,N_2752);
nand U3391 (N_3391,N_2745,N_2429);
xor U3392 (N_3392,N_2448,N_2779);
or U3393 (N_3393,N_2914,N_2806);
xnor U3394 (N_3394,N_2728,N_2465);
nor U3395 (N_3395,N_2718,N_2639);
and U3396 (N_3396,N_2423,N_2338);
and U3397 (N_3397,N_2990,N_2618);
xor U3398 (N_3398,N_2827,N_2523);
nor U3399 (N_3399,N_2457,N_2583);
xor U3400 (N_3400,N_2552,N_2563);
nand U3401 (N_3401,N_2920,N_2677);
nand U3402 (N_3402,N_2880,N_2312);
xor U3403 (N_3403,N_2720,N_2335);
and U3404 (N_3404,N_2516,N_2522);
or U3405 (N_3405,N_2550,N_2267);
or U3406 (N_3406,N_2534,N_2883);
nor U3407 (N_3407,N_2501,N_2787);
or U3408 (N_3408,N_2909,N_2848);
or U3409 (N_3409,N_2749,N_2443);
nand U3410 (N_3410,N_2795,N_2350);
nand U3411 (N_3411,N_2994,N_2487);
nor U3412 (N_3412,N_2496,N_2796);
nor U3413 (N_3413,N_2737,N_2865);
xor U3414 (N_3414,N_2964,N_2291);
nor U3415 (N_3415,N_2659,N_2990);
nor U3416 (N_3416,N_2535,N_2470);
or U3417 (N_3417,N_2736,N_2650);
nor U3418 (N_3418,N_2381,N_2639);
or U3419 (N_3419,N_2960,N_2843);
or U3420 (N_3420,N_2455,N_2480);
nand U3421 (N_3421,N_2701,N_2768);
nand U3422 (N_3422,N_2853,N_2898);
and U3423 (N_3423,N_2782,N_2558);
nand U3424 (N_3424,N_2871,N_2889);
and U3425 (N_3425,N_2849,N_2280);
or U3426 (N_3426,N_2278,N_2906);
or U3427 (N_3427,N_2347,N_2543);
and U3428 (N_3428,N_2269,N_2371);
nand U3429 (N_3429,N_2918,N_2549);
and U3430 (N_3430,N_2547,N_2973);
and U3431 (N_3431,N_2800,N_2556);
and U3432 (N_3432,N_2646,N_2761);
and U3433 (N_3433,N_2465,N_2928);
nand U3434 (N_3434,N_2428,N_2882);
and U3435 (N_3435,N_2567,N_2941);
or U3436 (N_3436,N_2494,N_2718);
nor U3437 (N_3437,N_2667,N_2822);
and U3438 (N_3438,N_2841,N_2809);
and U3439 (N_3439,N_2750,N_2790);
xor U3440 (N_3440,N_2586,N_2946);
xor U3441 (N_3441,N_2262,N_2282);
nor U3442 (N_3442,N_2608,N_2340);
xor U3443 (N_3443,N_2953,N_2412);
nand U3444 (N_3444,N_2379,N_2507);
or U3445 (N_3445,N_2350,N_2324);
nor U3446 (N_3446,N_2650,N_2527);
xor U3447 (N_3447,N_2999,N_2558);
nor U3448 (N_3448,N_2938,N_2505);
or U3449 (N_3449,N_2400,N_2656);
nor U3450 (N_3450,N_2292,N_2689);
or U3451 (N_3451,N_2525,N_2450);
and U3452 (N_3452,N_2617,N_2261);
xor U3453 (N_3453,N_2805,N_2916);
or U3454 (N_3454,N_2820,N_2354);
nor U3455 (N_3455,N_2819,N_2339);
nor U3456 (N_3456,N_2842,N_2409);
and U3457 (N_3457,N_2266,N_2344);
or U3458 (N_3458,N_2425,N_2352);
or U3459 (N_3459,N_2586,N_2311);
or U3460 (N_3460,N_2251,N_2548);
nand U3461 (N_3461,N_2889,N_2608);
nand U3462 (N_3462,N_2808,N_2624);
or U3463 (N_3463,N_2691,N_2995);
and U3464 (N_3464,N_2978,N_2633);
or U3465 (N_3465,N_2869,N_2339);
nand U3466 (N_3466,N_2615,N_2822);
nand U3467 (N_3467,N_2878,N_2353);
or U3468 (N_3468,N_2588,N_2399);
or U3469 (N_3469,N_2534,N_2577);
or U3470 (N_3470,N_2432,N_2756);
nand U3471 (N_3471,N_2852,N_2291);
nor U3472 (N_3472,N_2702,N_2947);
nand U3473 (N_3473,N_2260,N_2538);
nor U3474 (N_3474,N_2875,N_2672);
and U3475 (N_3475,N_2422,N_2309);
nor U3476 (N_3476,N_2693,N_2330);
or U3477 (N_3477,N_2984,N_2530);
or U3478 (N_3478,N_2630,N_2941);
or U3479 (N_3479,N_2308,N_2259);
xnor U3480 (N_3480,N_2543,N_2633);
or U3481 (N_3481,N_2803,N_2611);
nor U3482 (N_3482,N_2440,N_2581);
nor U3483 (N_3483,N_2471,N_2560);
nand U3484 (N_3484,N_2400,N_2938);
and U3485 (N_3485,N_2937,N_2324);
and U3486 (N_3486,N_2870,N_2998);
and U3487 (N_3487,N_2367,N_2521);
nand U3488 (N_3488,N_2762,N_2832);
nand U3489 (N_3489,N_2590,N_2772);
xor U3490 (N_3490,N_2628,N_2866);
nand U3491 (N_3491,N_2346,N_2364);
and U3492 (N_3492,N_2946,N_2585);
nand U3493 (N_3493,N_2638,N_2430);
nand U3494 (N_3494,N_2948,N_2755);
or U3495 (N_3495,N_2698,N_2306);
or U3496 (N_3496,N_2653,N_2460);
and U3497 (N_3497,N_2901,N_2267);
or U3498 (N_3498,N_2723,N_2630);
or U3499 (N_3499,N_2328,N_2689);
and U3500 (N_3500,N_2354,N_2931);
nor U3501 (N_3501,N_2807,N_2283);
nor U3502 (N_3502,N_2289,N_2874);
and U3503 (N_3503,N_2739,N_2449);
nor U3504 (N_3504,N_2457,N_2928);
and U3505 (N_3505,N_2323,N_2421);
nand U3506 (N_3506,N_2954,N_2783);
and U3507 (N_3507,N_2545,N_2643);
nor U3508 (N_3508,N_2695,N_2744);
nor U3509 (N_3509,N_2426,N_2657);
nand U3510 (N_3510,N_2848,N_2641);
or U3511 (N_3511,N_2945,N_2752);
and U3512 (N_3512,N_2757,N_2698);
nand U3513 (N_3513,N_2587,N_2867);
nor U3514 (N_3514,N_2729,N_2798);
and U3515 (N_3515,N_2257,N_2418);
or U3516 (N_3516,N_2360,N_2642);
and U3517 (N_3517,N_2347,N_2322);
and U3518 (N_3518,N_2847,N_2603);
nand U3519 (N_3519,N_2723,N_2801);
nand U3520 (N_3520,N_2887,N_2312);
or U3521 (N_3521,N_2305,N_2793);
or U3522 (N_3522,N_2525,N_2312);
nor U3523 (N_3523,N_2390,N_2639);
nor U3524 (N_3524,N_2346,N_2497);
and U3525 (N_3525,N_2757,N_2566);
and U3526 (N_3526,N_2899,N_2976);
nor U3527 (N_3527,N_2493,N_2851);
xnor U3528 (N_3528,N_2605,N_2768);
or U3529 (N_3529,N_2834,N_2822);
and U3530 (N_3530,N_2936,N_2349);
nand U3531 (N_3531,N_2374,N_2843);
or U3532 (N_3532,N_2961,N_2635);
and U3533 (N_3533,N_2663,N_2922);
and U3534 (N_3534,N_2628,N_2938);
or U3535 (N_3535,N_2847,N_2516);
and U3536 (N_3536,N_2805,N_2510);
nand U3537 (N_3537,N_2338,N_2569);
and U3538 (N_3538,N_2722,N_2321);
nor U3539 (N_3539,N_2722,N_2926);
xnor U3540 (N_3540,N_2568,N_2903);
and U3541 (N_3541,N_2301,N_2757);
nor U3542 (N_3542,N_2515,N_2305);
and U3543 (N_3543,N_2662,N_2420);
nor U3544 (N_3544,N_2659,N_2752);
or U3545 (N_3545,N_2561,N_2285);
and U3546 (N_3546,N_2669,N_2864);
nand U3547 (N_3547,N_2432,N_2842);
or U3548 (N_3548,N_2385,N_2908);
or U3549 (N_3549,N_2775,N_2555);
or U3550 (N_3550,N_2498,N_2993);
or U3551 (N_3551,N_2508,N_2970);
nand U3552 (N_3552,N_2475,N_2339);
nor U3553 (N_3553,N_2969,N_2814);
nand U3554 (N_3554,N_2631,N_2648);
nand U3555 (N_3555,N_2986,N_2345);
xnor U3556 (N_3556,N_2630,N_2780);
and U3557 (N_3557,N_2258,N_2486);
or U3558 (N_3558,N_2856,N_2966);
and U3559 (N_3559,N_2361,N_2635);
and U3560 (N_3560,N_2999,N_2655);
nor U3561 (N_3561,N_2387,N_2847);
xor U3562 (N_3562,N_2547,N_2751);
or U3563 (N_3563,N_2840,N_2380);
nand U3564 (N_3564,N_2374,N_2497);
xnor U3565 (N_3565,N_2978,N_2789);
and U3566 (N_3566,N_2471,N_2884);
or U3567 (N_3567,N_2979,N_2666);
or U3568 (N_3568,N_2670,N_2441);
or U3569 (N_3569,N_2396,N_2876);
nand U3570 (N_3570,N_2793,N_2866);
xnor U3571 (N_3571,N_2389,N_2479);
nand U3572 (N_3572,N_2536,N_2451);
or U3573 (N_3573,N_2787,N_2494);
and U3574 (N_3574,N_2413,N_2415);
nand U3575 (N_3575,N_2608,N_2567);
and U3576 (N_3576,N_2838,N_2276);
and U3577 (N_3577,N_2917,N_2433);
and U3578 (N_3578,N_2965,N_2683);
and U3579 (N_3579,N_2495,N_2360);
nor U3580 (N_3580,N_2576,N_2324);
nor U3581 (N_3581,N_2851,N_2962);
nand U3582 (N_3582,N_2944,N_2677);
xor U3583 (N_3583,N_2701,N_2342);
and U3584 (N_3584,N_2881,N_2704);
nand U3585 (N_3585,N_2808,N_2796);
or U3586 (N_3586,N_2508,N_2430);
and U3587 (N_3587,N_2808,N_2573);
nand U3588 (N_3588,N_2600,N_2992);
nand U3589 (N_3589,N_2582,N_2886);
and U3590 (N_3590,N_2613,N_2716);
nor U3591 (N_3591,N_2649,N_2579);
and U3592 (N_3592,N_2298,N_2478);
and U3593 (N_3593,N_2251,N_2760);
or U3594 (N_3594,N_2295,N_2778);
nand U3595 (N_3595,N_2869,N_2730);
nand U3596 (N_3596,N_2786,N_2867);
and U3597 (N_3597,N_2417,N_2408);
or U3598 (N_3598,N_2350,N_2651);
or U3599 (N_3599,N_2874,N_2935);
nand U3600 (N_3600,N_2927,N_2693);
xnor U3601 (N_3601,N_2913,N_2671);
and U3602 (N_3602,N_2921,N_2816);
nand U3603 (N_3603,N_2926,N_2400);
or U3604 (N_3604,N_2855,N_2446);
xnor U3605 (N_3605,N_2861,N_2802);
and U3606 (N_3606,N_2702,N_2970);
nand U3607 (N_3607,N_2949,N_2732);
nand U3608 (N_3608,N_2726,N_2401);
nand U3609 (N_3609,N_2547,N_2655);
or U3610 (N_3610,N_2533,N_2483);
or U3611 (N_3611,N_2262,N_2821);
and U3612 (N_3612,N_2423,N_2884);
nand U3613 (N_3613,N_2375,N_2423);
and U3614 (N_3614,N_2908,N_2323);
xor U3615 (N_3615,N_2992,N_2733);
nand U3616 (N_3616,N_2343,N_2569);
and U3617 (N_3617,N_2497,N_2896);
or U3618 (N_3618,N_2805,N_2615);
or U3619 (N_3619,N_2991,N_2714);
nand U3620 (N_3620,N_2304,N_2401);
and U3621 (N_3621,N_2811,N_2810);
and U3622 (N_3622,N_2949,N_2362);
nor U3623 (N_3623,N_2438,N_2805);
and U3624 (N_3624,N_2717,N_2425);
nor U3625 (N_3625,N_2473,N_2319);
nand U3626 (N_3626,N_2445,N_2301);
or U3627 (N_3627,N_2554,N_2720);
or U3628 (N_3628,N_2505,N_2732);
nor U3629 (N_3629,N_2452,N_2661);
and U3630 (N_3630,N_2271,N_2847);
xor U3631 (N_3631,N_2614,N_2915);
and U3632 (N_3632,N_2586,N_2481);
and U3633 (N_3633,N_2308,N_2697);
nor U3634 (N_3634,N_2393,N_2621);
or U3635 (N_3635,N_2512,N_2394);
and U3636 (N_3636,N_2973,N_2316);
or U3637 (N_3637,N_2895,N_2914);
or U3638 (N_3638,N_2759,N_2866);
or U3639 (N_3639,N_2583,N_2770);
nand U3640 (N_3640,N_2334,N_2412);
nand U3641 (N_3641,N_2604,N_2419);
or U3642 (N_3642,N_2490,N_2347);
xor U3643 (N_3643,N_2791,N_2388);
nand U3644 (N_3644,N_2404,N_2453);
or U3645 (N_3645,N_2254,N_2509);
and U3646 (N_3646,N_2320,N_2948);
and U3647 (N_3647,N_2913,N_2329);
and U3648 (N_3648,N_2452,N_2440);
nor U3649 (N_3649,N_2732,N_2404);
nand U3650 (N_3650,N_2610,N_2722);
nand U3651 (N_3651,N_2267,N_2712);
nand U3652 (N_3652,N_2561,N_2596);
and U3653 (N_3653,N_2900,N_2540);
xor U3654 (N_3654,N_2784,N_2809);
or U3655 (N_3655,N_2448,N_2424);
nor U3656 (N_3656,N_2764,N_2415);
and U3657 (N_3657,N_2570,N_2402);
xnor U3658 (N_3658,N_2420,N_2395);
nand U3659 (N_3659,N_2927,N_2289);
nor U3660 (N_3660,N_2285,N_2671);
or U3661 (N_3661,N_2465,N_2831);
or U3662 (N_3662,N_2310,N_2942);
nor U3663 (N_3663,N_2729,N_2827);
nand U3664 (N_3664,N_2919,N_2604);
nor U3665 (N_3665,N_2300,N_2775);
or U3666 (N_3666,N_2464,N_2708);
nor U3667 (N_3667,N_2927,N_2797);
nand U3668 (N_3668,N_2786,N_2711);
nand U3669 (N_3669,N_2714,N_2398);
and U3670 (N_3670,N_2560,N_2474);
or U3671 (N_3671,N_2636,N_2733);
nor U3672 (N_3672,N_2570,N_2437);
or U3673 (N_3673,N_2655,N_2957);
and U3674 (N_3674,N_2658,N_2385);
nand U3675 (N_3675,N_2258,N_2325);
or U3676 (N_3676,N_2965,N_2545);
and U3677 (N_3677,N_2337,N_2825);
and U3678 (N_3678,N_2508,N_2403);
and U3679 (N_3679,N_2750,N_2288);
nor U3680 (N_3680,N_2597,N_2415);
and U3681 (N_3681,N_2634,N_2774);
nand U3682 (N_3682,N_2657,N_2613);
or U3683 (N_3683,N_2301,N_2680);
xor U3684 (N_3684,N_2556,N_2320);
nor U3685 (N_3685,N_2921,N_2367);
or U3686 (N_3686,N_2977,N_2299);
nor U3687 (N_3687,N_2272,N_2335);
or U3688 (N_3688,N_2526,N_2442);
nor U3689 (N_3689,N_2914,N_2697);
and U3690 (N_3690,N_2331,N_2982);
nand U3691 (N_3691,N_2333,N_2405);
xor U3692 (N_3692,N_2594,N_2851);
or U3693 (N_3693,N_2352,N_2372);
or U3694 (N_3694,N_2807,N_2510);
nand U3695 (N_3695,N_2282,N_2765);
or U3696 (N_3696,N_2702,N_2429);
or U3697 (N_3697,N_2679,N_2812);
nor U3698 (N_3698,N_2951,N_2433);
and U3699 (N_3699,N_2726,N_2582);
and U3700 (N_3700,N_2442,N_2412);
or U3701 (N_3701,N_2953,N_2267);
and U3702 (N_3702,N_2866,N_2325);
nor U3703 (N_3703,N_2693,N_2282);
nor U3704 (N_3704,N_2708,N_2412);
or U3705 (N_3705,N_2264,N_2398);
and U3706 (N_3706,N_2698,N_2478);
nand U3707 (N_3707,N_2627,N_2447);
nor U3708 (N_3708,N_2794,N_2924);
nor U3709 (N_3709,N_2758,N_2422);
nor U3710 (N_3710,N_2573,N_2259);
nand U3711 (N_3711,N_2803,N_2996);
xnor U3712 (N_3712,N_2437,N_2428);
or U3713 (N_3713,N_2499,N_2998);
nand U3714 (N_3714,N_2430,N_2492);
or U3715 (N_3715,N_2601,N_2786);
nand U3716 (N_3716,N_2336,N_2417);
nand U3717 (N_3717,N_2813,N_2293);
or U3718 (N_3718,N_2852,N_2696);
and U3719 (N_3719,N_2280,N_2630);
and U3720 (N_3720,N_2325,N_2444);
and U3721 (N_3721,N_2416,N_2302);
or U3722 (N_3722,N_2939,N_2927);
nor U3723 (N_3723,N_2810,N_2587);
nand U3724 (N_3724,N_2492,N_2422);
and U3725 (N_3725,N_2454,N_2959);
and U3726 (N_3726,N_2700,N_2490);
and U3727 (N_3727,N_2880,N_2781);
and U3728 (N_3728,N_2601,N_2878);
or U3729 (N_3729,N_2677,N_2821);
or U3730 (N_3730,N_2767,N_2818);
nand U3731 (N_3731,N_2776,N_2614);
nor U3732 (N_3732,N_2906,N_2578);
and U3733 (N_3733,N_2469,N_2447);
or U3734 (N_3734,N_2364,N_2630);
and U3735 (N_3735,N_2888,N_2612);
nand U3736 (N_3736,N_2290,N_2535);
and U3737 (N_3737,N_2797,N_2760);
or U3738 (N_3738,N_2675,N_2256);
xnor U3739 (N_3739,N_2748,N_2502);
nand U3740 (N_3740,N_2504,N_2748);
or U3741 (N_3741,N_2809,N_2295);
or U3742 (N_3742,N_2927,N_2665);
nand U3743 (N_3743,N_2972,N_2260);
or U3744 (N_3744,N_2303,N_2424);
or U3745 (N_3745,N_2276,N_2416);
or U3746 (N_3746,N_2270,N_2360);
nand U3747 (N_3747,N_2817,N_2911);
nand U3748 (N_3748,N_2590,N_2503);
nand U3749 (N_3749,N_2333,N_2982);
and U3750 (N_3750,N_3493,N_3436);
or U3751 (N_3751,N_3642,N_3649);
nor U3752 (N_3752,N_3200,N_3687);
and U3753 (N_3753,N_3094,N_3282);
nor U3754 (N_3754,N_3121,N_3645);
or U3755 (N_3755,N_3636,N_3735);
and U3756 (N_3756,N_3748,N_3290);
nand U3757 (N_3757,N_3044,N_3297);
nand U3758 (N_3758,N_3679,N_3669);
or U3759 (N_3759,N_3003,N_3527);
or U3760 (N_3760,N_3261,N_3575);
or U3761 (N_3761,N_3123,N_3066);
or U3762 (N_3762,N_3439,N_3259);
nor U3763 (N_3763,N_3078,N_3365);
or U3764 (N_3764,N_3035,N_3042);
nand U3765 (N_3765,N_3143,N_3092);
or U3766 (N_3766,N_3271,N_3103);
nand U3767 (N_3767,N_3579,N_3742);
nand U3768 (N_3768,N_3631,N_3445);
or U3769 (N_3769,N_3666,N_3457);
and U3770 (N_3770,N_3516,N_3670);
nor U3771 (N_3771,N_3061,N_3032);
or U3772 (N_3772,N_3058,N_3302);
or U3773 (N_3773,N_3404,N_3084);
nor U3774 (N_3774,N_3437,N_3067);
and U3775 (N_3775,N_3165,N_3415);
and U3776 (N_3776,N_3471,N_3255);
nor U3777 (N_3777,N_3647,N_3624);
nor U3778 (N_3778,N_3623,N_3456);
nand U3779 (N_3779,N_3208,N_3733);
nand U3780 (N_3780,N_3266,N_3586);
and U3781 (N_3781,N_3717,N_3303);
and U3782 (N_3782,N_3225,N_3425);
or U3783 (N_3783,N_3651,N_3611);
xor U3784 (N_3784,N_3336,N_3264);
nand U3785 (N_3785,N_3251,N_3244);
or U3786 (N_3786,N_3479,N_3531);
nor U3787 (N_3787,N_3508,N_3093);
and U3788 (N_3788,N_3263,N_3096);
or U3789 (N_3789,N_3373,N_3024);
or U3790 (N_3790,N_3104,N_3022);
nor U3791 (N_3791,N_3190,N_3332);
and U3792 (N_3792,N_3051,N_3308);
xor U3793 (N_3793,N_3473,N_3227);
and U3794 (N_3794,N_3653,N_3366);
nor U3795 (N_3795,N_3744,N_3343);
and U3796 (N_3796,N_3423,N_3242);
and U3797 (N_3797,N_3671,N_3434);
xor U3798 (N_3798,N_3607,N_3729);
or U3799 (N_3799,N_3345,N_3468);
nor U3800 (N_3800,N_3048,N_3149);
xor U3801 (N_3801,N_3112,N_3464);
nand U3802 (N_3802,N_3069,N_3681);
nor U3803 (N_3803,N_3346,N_3201);
and U3804 (N_3804,N_3416,N_3284);
nor U3805 (N_3805,N_3660,N_3135);
nor U3806 (N_3806,N_3538,N_3128);
and U3807 (N_3807,N_3463,N_3523);
nand U3808 (N_3808,N_3283,N_3406);
nand U3809 (N_3809,N_3617,N_3585);
or U3810 (N_3810,N_3502,N_3378);
and U3811 (N_3811,N_3002,N_3007);
nor U3812 (N_3812,N_3286,N_3004);
and U3813 (N_3813,N_3550,N_3555);
and U3814 (N_3814,N_3257,N_3099);
and U3815 (N_3815,N_3533,N_3221);
nor U3816 (N_3816,N_3388,N_3235);
or U3817 (N_3817,N_3161,N_3402);
and U3818 (N_3818,N_3565,N_3447);
or U3819 (N_3819,N_3719,N_3721);
and U3820 (N_3820,N_3601,N_3041);
or U3821 (N_3821,N_3558,N_3386);
nor U3822 (N_3822,N_3191,N_3610);
nor U3823 (N_3823,N_3151,N_3015);
and U3824 (N_3824,N_3612,N_3029);
nand U3825 (N_3825,N_3139,N_3728);
and U3826 (N_3826,N_3278,N_3148);
nor U3827 (N_3827,N_3699,N_3009);
and U3828 (N_3828,N_3050,N_3339);
nand U3829 (N_3829,N_3424,N_3497);
or U3830 (N_3830,N_3747,N_3134);
or U3831 (N_3831,N_3608,N_3480);
and U3832 (N_3832,N_3548,N_3293);
nor U3833 (N_3833,N_3218,N_3556);
and U3834 (N_3834,N_3299,N_3563);
xor U3835 (N_3835,N_3155,N_3605);
or U3836 (N_3836,N_3432,N_3389);
nand U3837 (N_3837,N_3491,N_3317);
or U3838 (N_3838,N_3391,N_3357);
or U3839 (N_3839,N_3552,N_3226);
nand U3840 (N_3840,N_3458,N_3206);
nand U3841 (N_3841,N_3140,N_3599);
and U3842 (N_3842,N_3509,N_3018);
and U3843 (N_3843,N_3310,N_3247);
nand U3844 (N_3844,N_3011,N_3576);
nor U3845 (N_3845,N_3023,N_3662);
nor U3846 (N_3846,N_3213,N_3364);
nand U3847 (N_3847,N_3202,N_3668);
xnor U3848 (N_3848,N_3709,N_3132);
and U3849 (N_3849,N_3229,N_3499);
and U3850 (N_3850,N_3684,N_3276);
nor U3851 (N_3851,N_3562,N_3539);
nand U3852 (N_3852,N_3064,N_3057);
or U3853 (N_3853,N_3145,N_3622);
nor U3854 (N_3854,N_3354,N_3020);
and U3855 (N_3855,N_3073,N_3138);
nor U3856 (N_3856,N_3420,N_3028);
nor U3857 (N_3857,N_3147,N_3595);
or U3858 (N_3858,N_3697,N_3506);
nor U3859 (N_3859,N_3693,N_3700);
xor U3860 (N_3860,N_3698,N_3708);
or U3861 (N_3861,N_3498,N_3718);
or U3862 (N_3862,N_3187,N_3427);
and U3863 (N_3863,N_3583,N_3535);
and U3864 (N_3864,N_3074,N_3083);
nand U3865 (N_3865,N_3627,N_3426);
or U3866 (N_3866,N_3688,N_3301);
nand U3867 (N_3867,N_3513,N_3342);
xor U3868 (N_3868,N_3216,N_3379);
nand U3869 (N_3869,N_3465,N_3250);
nand U3870 (N_3870,N_3678,N_3108);
nand U3871 (N_3871,N_3566,N_3363);
xor U3872 (N_3872,N_3082,N_3109);
and U3873 (N_3873,N_3285,N_3228);
or U3874 (N_3874,N_3397,N_3325);
nor U3875 (N_3875,N_3484,N_3314);
nor U3876 (N_3876,N_3376,N_3403);
xnor U3877 (N_3877,N_3609,N_3144);
nor U3878 (N_3878,N_3037,N_3287);
nor U3879 (N_3879,N_3316,N_3547);
and U3880 (N_3880,N_3025,N_3635);
nand U3881 (N_3881,N_3163,N_3353);
and U3882 (N_3882,N_3470,N_3300);
nor U3883 (N_3883,N_3455,N_3331);
xor U3884 (N_3884,N_3152,N_3628);
xor U3885 (N_3885,N_3568,N_3127);
nand U3886 (N_3886,N_3478,N_3580);
nand U3887 (N_3887,N_3703,N_3385);
xnor U3888 (N_3888,N_3260,N_3304);
nand U3889 (N_3889,N_3312,N_3160);
nand U3890 (N_3890,N_3210,N_3462);
and U3891 (N_3891,N_3641,N_3292);
nor U3892 (N_3892,N_3722,N_3615);
nor U3893 (N_3893,N_3475,N_3217);
and U3894 (N_3894,N_3536,N_3546);
or U3895 (N_3895,N_3514,N_3168);
or U3896 (N_3896,N_3253,N_3008);
nor U3897 (N_3897,N_3352,N_3344);
nor U3898 (N_3898,N_3534,N_3233);
nor U3899 (N_3899,N_3569,N_3311);
nor U3900 (N_3900,N_3400,N_3162);
or U3901 (N_3901,N_3542,N_3644);
nor U3902 (N_3902,N_3196,N_3249);
or U3903 (N_3903,N_3749,N_3105);
and U3904 (N_3904,N_3665,N_3598);
or U3905 (N_3905,N_3381,N_3421);
nand U3906 (N_3906,N_3474,N_3488);
nand U3907 (N_3907,N_3459,N_3504);
xnor U3908 (N_3908,N_3065,N_3046);
nand U3909 (N_3909,N_3690,N_3731);
or U3910 (N_3910,N_3630,N_3650);
nand U3911 (N_3911,N_3019,N_3492);
nand U3912 (N_3912,N_3730,N_3604);
or U3913 (N_3913,N_3183,N_3347);
and U3914 (N_3914,N_3571,N_3359);
nor U3915 (N_3915,N_3674,N_3000);
nor U3916 (N_3916,N_3382,N_3113);
nand U3917 (N_3917,N_3476,N_3430);
nand U3918 (N_3918,N_3646,N_3095);
or U3919 (N_3919,N_3574,N_3137);
nor U3920 (N_3920,N_3392,N_3477);
nor U3921 (N_3921,N_3116,N_3510);
and U3922 (N_3922,N_3619,N_3172);
and U3923 (N_3923,N_3452,N_3141);
and U3924 (N_3924,N_3340,N_3356);
or U3925 (N_3925,N_3517,N_3330);
nand U3926 (N_3926,N_3413,N_3159);
nor U3927 (N_3927,N_3489,N_3664);
or U3928 (N_3928,N_3106,N_3169);
and U3929 (N_3929,N_3238,N_3237);
and U3930 (N_3930,N_3596,N_3232);
nand U3931 (N_3931,N_3179,N_3068);
or U3932 (N_3932,N_3692,N_3485);
nand U3933 (N_3933,N_3350,N_3387);
or U3934 (N_3934,N_3632,N_3661);
or U3935 (N_3935,N_3245,N_3176);
xnor U3936 (N_3936,N_3383,N_3146);
nand U3937 (N_3937,N_3482,N_3732);
nand U3938 (N_3938,N_3408,N_3265);
and U3939 (N_3939,N_3494,N_3702);
nand U3940 (N_3940,N_3637,N_3648);
nand U3941 (N_3941,N_3736,N_3192);
and U3942 (N_3942,N_3254,N_3659);
nand U3943 (N_3943,N_3043,N_3710);
and U3944 (N_3944,N_3685,N_3189);
nand U3945 (N_3945,N_3587,N_3173);
nand U3946 (N_3946,N_3358,N_3234);
nand U3947 (N_3947,N_3422,N_3184);
nand U3948 (N_3948,N_3560,N_3372);
or U3949 (N_3949,N_3174,N_3001);
or U3950 (N_3950,N_3481,N_3561);
or U3951 (N_3951,N_3100,N_3602);
nand U3952 (N_3952,N_3469,N_3530);
xor U3953 (N_3953,N_3279,N_3031);
nor U3954 (N_3954,N_3472,N_3487);
or U3955 (N_3955,N_3305,N_3272);
and U3956 (N_3956,N_3014,N_3428);
nor U3957 (N_3957,N_3375,N_3501);
and U3958 (N_3958,N_3394,N_3686);
xnor U3959 (N_3959,N_3326,N_3246);
and U3960 (N_3960,N_3496,N_3275);
and U3961 (N_3961,N_3407,N_3440);
and U3962 (N_3962,N_3572,N_3030);
nor U3963 (N_3963,N_3115,N_3417);
nor U3964 (N_3964,N_3089,N_3349);
and U3965 (N_3965,N_3338,N_3435);
and U3966 (N_3966,N_3195,N_3142);
or U3967 (N_3967,N_3180,N_3091);
nand U3968 (N_3968,N_3153,N_3277);
xor U3969 (N_3969,N_3321,N_3578);
or U3970 (N_3970,N_3268,N_3738);
xor U3971 (N_3971,N_3118,N_3157);
and U3972 (N_3972,N_3052,N_3027);
xnor U3973 (N_3973,N_3267,N_3626);
and U3974 (N_3974,N_3097,N_3727);
nor U3975 (N_3975,N_3429,N_3170);
and U3976 (N_3976,N_3682,N_3680);
nand U3977 (N_3977,N_3706,N_3743);
and U3978 (N_3978,N_3274,N_3695);
or U3979 (N_3979,N_3318,N_3655);
nand U3980 (N_3980,N_3291,N_3614);
and U3981 (N_3981,N_3315,N_3131);
nor U3982 (N_3982,N_3212,N_3705);
nor U3983 (N_3983,N_3197,N_3581);
and U3984 (N_3984,N_3038,N_3467);
and U3985 (N_3985,N_3593,N_3449);
nand U3986 (N_3986,N_3460,N_3399);
nand U3987 (N_3987,N_3307,N_3294);
nor U3988 (N_3988,N_3529,N_3088);
nand U3989 (N_3989,N_3652,N_3584);
nand U3990 (N_3990,N_3348,N_3613);
xor U3991 (N_3991,N_3241,N_3553);
and U3992 (N_3992,N_3567,N_3181);
and U3993 (N_3993,N_3518,N_3711);
nand U3994 (N_3994,N_3367,N_3683);
or U3995 (N_3995,N_3133,N_3198);
and U3996 (N_3996,N_3401,N_3324);
nand U3997 (N_3997,N_3746,N_3124);
and U3998 (N_3998,N_3441,N_3039);
nor U3999 (N_3999,N_3570,N_3256);
and U4000 (N_4000,N_3059,N_3588);
or U4001 (N_4001,N_3507,N_3085);
nand U4002 (N_4002,N_3248,N_3616);
or U4003 (N_4003,N_3620,N_3240);
nor U4004 (N_4004,N_3466,N_3111);
and U4005 (N_4005,N_3006,N_3203);
and U4006 (N_4006,N_3712,N_3696);
nand U4007 (N_4007,N_3270,N_3483);
nand U4008 (N_4008,N_3714,N_3384);
xnor U4009 (N_4009,N_3543,N_3040);
nand U4010 (N_4010,N_3745,N_3362);
or U4011 (N_4011,N_3371,N_3656);
or U4012 (N_4012,N_3448,N_3577);
nand U4013 (N_4013,N_3657,N_3182);
or U4014 (N_4014,N_3512,N_3419);
nor U4015 (N_4015,N_3205,N_3438);
and U4016 (N_4016,N_3351,N_3298);
nor U4017 (N_4017,N_3676,N_3269);
and U4018 (N_4018,N_3102,N_3405);
nor U4019 (N_4019,N_3713,N_3689);
or U4020 (N_4020,N_3414,N_3062);
or U4021 (N_4021,N_3126,N_3557);
nor U4022 (N_4022,N_3110,N_3360);
nand U4023 (N_4023,N_3672,N_3258);
and U4024 (N_4024,N_3075,N_3519);
nor U4025 (N_4025,N_3412,N_3211);
nor U4026 (N_4026,N_3117,N_3296);
xnor U4027 (N_4027,N_3230,N_3451);
and U4028 (N_4028,N_3220,N_3734);
and U4029 (N_4029,N_3071,N_3224);
or U4030 (N_4030,N_3590,N_3185);
and U4031 (N_4031,N_3716,N_3167);
nand U4032 (N_4032,N_3390,N_3219);
and U4033 (N_4033,N_3573,N_3418);
and U4034 (N_4034,N_3033,N_3053);
and U4035 (N_4035,N_3629,N_3334);
nand U4036 (N_4036,N_3600,N_3070);
nand U4037 (N_4037,N_3431,N_3280);
or U4038 (N_4038,N_3740,N_3016);
and U4039 (N_4039,N_3072,N_3544);
and U4040 (N_4040,N_3122,N_3520);
and U4041 (N_4041,N_3374,N_3398);
nand U4042 (N_4042,N_3737,N_3329);
xnor U4043 (N_4043,N_3047,N_3076);
or U4044 (N_4044,N_3618,N_3444);
or U4045 (N_4045,N_3724,N_3026);
and U4046 (N_4046,N_3175,N_3154);
nand U4047 (N_4047,N_3704,N_3209);
nor U4048 (N_4048,N_3098,N_3594);
and U4049 (N_4049,N_3120,N_3054);
nor U4050 (N_4050,N_3288,N_3453);
nand U4051 (N_4051,N_3446,N_3355);
nand U4052 (N_4052,N_3522,N_3333);
and U4053 (N_4053,N_3551,N_3540);
and U4054 (N_4054,N_3273,N_3204);
xnor U4055 (N_4055,N_3691,N_3306);
and U4056 (N_4056,N_3320,N_3327);
xnor U4057 (N_4057,N_3136,N_3087);
or U4058 (N_4058,N_3720,N_3638);
and U4059 (N_4059,N_3725,N_3396);
nor U4060 (N_4060,N_3582,N_3081);
nor U4061 (N_4061,N_3036,N_3177);
nor U4062 (N_4062,N_3675,N_3323);
or U4063 (N_4063,N_3049,N_3393);
or U4064 (N_4064,N_3361,N_3701);
or U4065 (N_4065,N_3156,N_3012);
nor U4066 (N_4066,N_3634,N_3597);
nand U4067 (N_4067,N_3673,N_3564);
nand U4068 (N_4068,N_3214,N_3503);
xnor U4069 (N_4069,N_3017,N_3505);
nor U4070 (N_4070,N_3090,N_3335);
nor U4071 (N_4071,N_3454,N_3549);
nand U4072 (N_4072,N_3461,N_3055);
and U4073 (N_4073,N_3541,N_3677);
or U4074 (N_4074,N_3125,N_3521);
nor U4075 (N_4075,N_3319,N_3309);
or U4076 (N_4076,N_3707,N_3341);
xnor U4077 (N_4077,N_3639,N_3164);
and U4078 (N_4078,N_3739,N_3500);
or U4079 (N_4079,N_3486,N_3410);
or U4080 (N_4080,N_3591,N_3199);
nor U4081 (N_4081,N_3289,N_3194);
nand U4082 (N_4082,N_3328,N_3545);
nor U4083 (N_4083,N_3369,N_3231);
xnor U4084 (N_4084,N_3063,N_3490);
and U4085 (N_4085,N_3524,N_3411);
nand U4086 (N_4086,N_3021,N_3045);
and U4087 (N_4087,N_3243,N_3433);
nor U4088 (N_4088,N_3239,N_3150);
nand U4089 (N_4089,N_3129,N_3056);
and U4090 (N_4090,N_3442,N_3079);
nor U4091 (N_4091,N_3726,N_3114);
or U4092 (N_4092,N_3667,N_3295);
xor U4093 (N_4093,N_3409,N_3322);
or U4094 (N_4094,N_3526,N_3715);
and U4095 (N_4095,N_3171,N_3368);
or U4096 (N_4096,N_3223,N_3443);
or U4097 (N_4097,N_3337,N_3589);
or U4098 (N_4098,N_3262,N_3625);
and U4099 (N_4099,N_3119,N_3640);
xnor U4100 (N_4100,N_3511,N_3060);
nand U4101 (N_4101,N_3450,N_3252);
nor U4102 (N_4102,N_3658,N_3178);
xnor U4103 (N_4103,N_3380,N_3186);
or U4104 (N_4104,N_3606,N_3080);
nand U4105 (N_4105,N_3633,N_3215);
or U4106 (N_4106,N_3086,N_3005);
or U4107 (N_4107,N_3663,N_3741);
nor U4108 (N_4108,N_3723,N_3592);
nor U4109 (N_4109,N_3188,N_3525);
nand U4110 (N_4110,N_3158,N_3193);
or U4111 (N_4111,N_3554,N_3515);
and U4112 (N_4112,N_3370,N_3495);
and U4113 (N_4113,N_3077,N_3010);
nand U4114 (N_4114,N_3130,N_3621);
nand U4115 (N_4115,N_3166,N_3034);
or U4116 (N_4116,N_3107,N_3395);
xor U4117 (N_4117,N_3643,N_3101);
and U4118 (N_4118,N_3694,N_3236);
and U4119 (N_4119,N_3207,N_3603);
xnor U4120 (N_4120,N_3013,N_3654);
xor U4121 (N_4121,N_3281,N_3528);
xnor U4122 (N_4122,N_3222,N_3377);
or U4123 (N_4123,N_3313,N_3559);
or U4124 (N_4124,N_3537,N_3532);
xor U4125 (N_4125,N_3488,N_3256);
or U4126 (N_4126,N_3384,N_3274);
or U4127 (N_4127,N_3733,N_3297);
nor U4128 (N_4128,N_3158,N_3610);
nor U4129 (N_4129,N_3550,N_3256);
nand U4130 (N_4130,N_3288,N_3219);
and U4131 (N_4131,N_3150,N_3445);
nand U4132 (N_4132,N_3070,N_3593);
nand U4133 (N_4133,N_3615,N_3478);
nand U4134 (N_4134,N_3555,N_3514);
nor U4135 (N_4135,N_3563,N_3673);
or U4136 (N_4136,N_3708,N_3619);
and U4137 (N_4137,N_3045,N_3447);
and U4138 (N_4138,N_3103,N_3620);
and U4139 (N_4139,N_3489,N_3205);
or U4140 (N_4140,N_3278,N_3540);
nand U4141 (N_4141,N_3093,N_3364);
nand U4142 (N_4142,N_3076,N_3527);
or U4143 (N_4143,N_3607,N_3629);
nand U4144 (N_4144,N_3361,N_3625);
nor U4145 (N_4145,N_3099,N_3740);
and U4146 (N_4146,N_3692,N_3094);
xnor U4147 (N_4147,N_3046,N_3182);
xnor U4148 (N_4148,N_3046,N_3265);
xor U4149 (N_4149,N_3671,N_3447);
and U4150 (N_4150,N_3550,N_3723);
and U4151 (N_4151,N_3531,N_3652);
nor U4152 (N_4152,N_3333,N_3096);
nand U4153 (N_4153,N_3030,N_3293);
or U4154 (N_4154,N_3047,N_3445);
and U4155 (N_4155,N_3690,N_3516);
and U4156 (N_4156,N_3061,N_3259);
or U4157 (N_4157,N_3525,N_3521);
xnor U4158 (N_4158,N_3248,N_3653);
and U4159 (N_4159,N_3009,N_3160);
and U4160 (N_4160,N_3629,N_3713);
nand U4161 (N_4161,N_3149,N_3195);
nor U4162 (N_4162,N_3458,N_3486);
nor U4163 (N_4163,N_3360,N_3681);
nor U4164 (N_4164,N_3023,N_3291);
and U4165 (N_4165,N_3073,N_3017);
nand U4166 (N_4166,N_3274,N_3055);
and U4167 (N_4167,N_3300,N_3624);
nor U4168 (N_4168,N_3458,N_3593);
xnor U4169 (N_4169,N_3107,N_3572);
nor U4170 (N_4170,N_3434,N_3418);
and U4171 (N_4171,N_3297,N_3599);
and U4172 (N_4172,N_3400,N_3270);
or U4173 (N_4173,N_3686,N_3232);
or U4174 (N_4174,N_3320,N_3447);
xor U4175 (N_4175,N_3591,N_3263);
or U4176 (N_4176,N_3592,N_3381);
or U4177 (N_4177,N_3475,N_3730);
or U4178 (N_4178,N_3386,N_3371);
nand U4179 (N_4179,N_3364,N_3250);
xor U4180 (N_4180,N_3473,N_3281);
or U4181 (N_4181,N_3673,N_3280);
nand U4182 (N_4182,N_3063,N_3228);
and U4183 (N_4183,N_3287,N_3352);
nand U4184 (N_4184,N_3393,N_3129);
or U4185 (N_4185,N_3588,N_3262);
and U4186 (N_4186,N_3366,N_3583);
nand U4187 (N_4187,N_3210,N_3713);
xnor U4188 (N_4188,N_3646,N_3148);
and U4189 (N_4189,N_3286,N_3572);
nor U4190 (N_4190,N_3055,N_3548);
nor U4191 (N_4191,N_3481,N_3398);
or U4192 (N_4192,N_3648,N_3276);
and U4193 (N_4193,N_3119,N_3343);
or U4194 (N_4194,N_3203,N_3570);
xnor U4195 (N_4195,N_3664,N_3655);
and U4196 (N_4196,N_3570,N_3593);
nor U4197 (N_4197,N_3579,N_3486);
and U4198 (N_4198,N_3179,N_3066);
nor U4199 (N_4199,N_3067,N_3298);
nor U4200 (N_4200,N_3084,N_3667);
nor U4201 (N_4201,N_3345,N_3327);
nand U4202 (N_4202,N_3671,N_3501);
nor U4203 (N_4203,N_3418,N_3446);
and U4204 (N_4204,N_3211,N_3561);
or U4205 (N_4205,N_3691,N_3411);
or U4206 (N_4206,N_3152,N_3423);
nand U4207 (N_4207,N_3269,N_3586);
nand U4208 (N_4208,N_3376,N_3157);
nor U4209 (N_4209,N_3190,N_3690);
xnor U4210 (N_4210,N_3036,N_3088);
nand U4211 (N_4211,N_3068,N_3528);
nor U4212 (N_4212,N_3249,N_3445);
and U4213 (N_4213,N_3654,N_3105);
or U4214 (N_4214,N_3513,N_3204);
and U4215 (N_4215,N_3714,N_3364);
nor U4216 (N_4216,N_3377,N_3269);
or U4217 (N_4217,N_3069,N_3031);
nand U4218 (N_4218,N_3246,N_3504);
and U4219 (N_4219,N_3394,N_3455);
nor U4220 (N_4220,N_3573,N_3219);
nor U4221 (N_4221,N_3745,N_3009);
nor U4222 (N_4222,N_3331,N_3709);
nor U4223 (N_4223,N_3345,N_3309);
or U4224 (N_4224,N_3665,N_3376);
or U4225 (N_4225,N_3498,N_3061);
nor U4226 (N_4226,N_3448,N_3408);
xnor U4227 (N_4227,N_3048,N_3377);
nand U4228 (N_4228,N_3635,N_3383);
xor U4229 (N_4229,N_3311,N_3328);
nor U4230 (N_4230,N_3057,N_3264);
nor U4231 (N_4231,N_3131,N_3517);
and U4232 (N_4232,N_3115,N_3197);
or U4233 (N_4233,N_3135,N_3461);
or U4234 (N_4234,N_3272,N_3549);
or U4235 (N_4235,N_3459,N_3089);
nor U4236 (N_4236,N_3484,N_3286);
and U4237 (N_4237,N_3440,N_3477);
and U4238 (N_4238,N_3444,N_3239);
nand U4239 (N_4239,N_3187,N_3627);
nand U4240 (N_4240,N_3182,N_3539);
nor U4241 (N_4241,N_3018,N_3268);
nor U4242 (N_4242,N_3201,N_3040);
nor U4243 (N_4243,N_3166,N_3339);
and U4244 (N_4244,N_3522,N_3412);
nand U4245 (N_4245,N_3333,N_3704);
nand U4246 (N_4246,N_3341,N_3235);
nor U4247 (N_4247,N_3144,N_3193);
or U4248 (N_4248,N_3617,N_3477);
xnor U4249 (N_4249,N_3424,N_3529);
nand U4250 (N_4250,N_3665,N_3628);
or U4251 (N_4251,N_3611,N_3365);
nor U4252 (N_4252,N_3042,N_3281);
nand U4253 (N_4253,N_3202,N_3411);
or U4254 (N_4254,N_3711,N_3206);
nand U4255 (N_4255,N_3419,N_3719);
nand U4256 (N_4256,N_3630,N_3242);
nor U4257 (N_4257,N_3263,N_3486);
or U4258 (N_4258,N_3120,N_3143);
xor U4259 (N_4259,N_3681,N_3507);
and U4260 (N_4260,N_3703,N_3379);
or U4261 (N_4261,N_3522,N_3705);
nor U4262 (N_4262,N_3677,N_3438);
and U4263 (N_4263,N_3120,N_3233);
nand U4264 (N_4264,N_3027,N_3194);
or U4265 (N_4265,N_3162,N_3473);
nand U4266 (N_4266,N_3190,N_3465);
or U4267 (N_4267,N_3445,N_3658);
nor U4268 (N_4268,N_3647,N_3744);
xor U4269 (N_4269,N_3435,N_3229);
and U4270 (N_4270,N_3184,N_3362);
nand U4271 (N_4271,N_3624,N_3367);
nor U4272 (N_4272,N_3572,N_3101);
xor U4273 (N_4273,N_3658,N_3036);
and U4274 (N_4274,N_3306,N_3282);
nand U4275 (N_4275,N_3700,N_3334);
or U4276 (N_4276,N_3673,N_3047);
xnor U4277 (N_4277,N_3128,N_3617);
and U4278 (N_4278,N_3207,N_3718);
and U4279 (N_4279,N_3656,N_3749);
nand U4280 (N_4280,N_3156,N_3497);
nand U4281 (N_4281,N_3073,N_3709);
and U4282 (N_4282,N_3365,N_3328);
xnor U4283 (N_4283,N_3454,N_3113);
xnor U4284 (N_4284,N_3282,N_3138);
nand U4285 (N_4285,N_3493,N_3541);
and U4286 (N_4286,N_3133,N_3463);
nand U4287 (N_4287,N_3347,N_3654);
nor U4288 (N_4288,N_3060,N_3068);
and U4289 (N_4289,N_3676,N_3716);
nor U4290 (N_4290,N_3044,N_3640);
nor U4291 (N_4291,N_3272,N_3169);
and U4292 (N_4292,N_3439,N_3383);
nand U4293 (N_4293,N_3451,N_3060);
and U4294 (N_4294,N_3313,N_3561);
and U4295 (N_4295,N_3714,N_3571);
nor U4296 (N_4296,N_3646,N_3378);
nor U4297 (N_4297,N_3186,N_3534);
or U4298 (N_4298,N_3581,N_3694);
or U4299 (N_4299,N_3647,N_3303);
or U4300 (N_4300,N_3010,N_3726);
nor U4301 (N_4301,N_3240,N_3449);
nand U4302 (N_4302,N_3007,N_3378);
nand U4303 (N_4303,N_3088,N_3262);
nor U4304 (N_4304,N_3386,N_3487);
and U4305 (N_4305,N_3603,N_3341);
and U4306 (N_4306,N_3099,N_3747);
or U4307 (N_4307,N_3226,N_3464);
and U4308 (N_4308,N_3539,N_3269);
nor U4309 (N_4309,N_3241,N_3102);
nand U4310 (N_4310,N_3515,N_3739);
xnor U4311 (N_4311,N_3104,N_3167);
nor U4312 (N_4312,N_3269,N_3469);
or U4313 (N_4313,N_3658,N_3465);
or U4314 (N_4314,N_3145,N_3515);
or U4315 (N_4315,N_3456,N_3619);
nand U4316 (N_4316,N_3675,N_3115);
nand U4317 (N_4317,N_3151,N_3020);
and U4318 (N_4318,N_3111,N_3143);
and U4319 (N_4319,N_3435,N_3378);
nor U4320 (N_4320,N_3405,N_3260);
and U4321 (N_4321,N_3389,N_3549);
and U4322 (N_4322,N_3593,N_3516);
nand U4323 (N_4323,N_3332,N_3414);
xor U4324 (N_4324,N_3477,N_3634);
and U4325 (N_4325,N_3287,N_3623);
nor U4326 (N_4326,N_3620,N_3308);
or U4327 (N_4327,N_3003,N_3100);
nor U4328 (N_4328,N_3694,N_3506);
nand U4329 (N_4329,N_3447,N_3614);
nor U4330 (N_4330,N_3398,N_3470);
and U4331 (N_4331,N_3540,N_3577);
or U4332 (N_4332,N_3296,N_3383);
or U4333 (N_4333,N_3379,N_3657);
nand U4334 (N_4334,N_3264,N_3657);
xor U4335 (N_4335,N_3330,N_3058);
and U4336 (N_4336,N_3120,N_3288);
and U4337 (N_4337,N_3589,N_3616);
or U4338 (N_4338,N_3680,N_3389);
nand U4339 (N_4339,N_3435,N_3189);
or U4340 (N_4340,N_3529,N_3392);
or U4341 (N_4341,N_3422,N_3389);
nor U4342 (N_4342,N_3164,N_3338);
xnor U4343 (N_4343,N_3501,N_3483);
nand U4344 (N_4344,N_3669,N_3242);
nand U4345 (N_4345,N_3194,N_3036);
nand U4346 (N_4346,N_3489,N_3534);
and U4347 (N_4347,N_3006,N_3671);
nor U4348 (N_4348,N_3702,N_3707);
and U4349 (N_4349,N_3684,N_3645);
nand U4350 (N_4350,N_3508,N_3164);
nor U4351 (N_4351,N_3137,N_3705);
and U4352 (N_4352,N_3681,N_3011);
nand U4353 (N_4353,N_3268,N_3697);
and U4354 (N_4354,N_3149,N_3086);
nor U4355 (N_4355,N_3395,N_3693);
and U4356 (N_4356,N_3609,N_3415);
or U4357 (N_4357,N_3258,N_3269);
and U4358 (N_4358,N_3036,N_3413);
or U4359 (N_4359,N_3586,N_3102);
and U4360 (N_4360,N_3184,N_3007);
or U4361 (N_4361,N_3537,N_3609);
and U4362 (N_4362,N_3345,N_3435);
and U4363 (N_4363,N_3713,N_3472);
nor U4364 (N_4364,N_3076,N_3110);
xnor U4365 (N_4365,N_3346,N_3135);
or U4366 (N_4366,N_3552,N_3247);
or U4367 (N_4367,N_3198,N_3494);
or U4368 (N_4368,N_3353,N_3090);
nand U4369 (N_4369,N_3722,N_3599);
or U4370 (N_4370,N_3681,N_3096);
and U4371 (N_4371,N_3307,N_3723);
nor U4372 (N_4372,N_3249,N_3201);
and U4373 (N_4373,N_3530,N_3644);
nor U4374 (N_4374,N_3213,N_3224);
and U4375 (N_4375,N_3679,N_3049);
and U4376 (N_4376,N_3077,N_3488);
xnor U4377 (N_4377,N_3727,N_3542);
nand U4378 (N_4378,N_3411,N_3640);
xnor U4379 (N_4379,N_3395,N_3072);
or U4380 (N_4380,N_3746,N_3221);
and U4381 (N_4381,N_3159,N_3359);
nand U4382 (N_4382,N_3112,N_3462);
nand U4383 (N_4383,N_3321,N_3069);
nand U4384 (N_4384,N_3716,N_3639);
nor U4385 (N_4385,N_3208,N_3327);
and U4386 (N_4386,N_3625,N_3075);
and U4387 (N_4387,N_3043,N_3054);
nor U4388 (N_4388,N_3125,N_3195);
nor U4389 (N_4389,N_3167,N_3056);
nor U4390 (N_4390,N_3401,N_3270);
nand U4391 (N_4391,N_3125,N_3420);
or U4392 (N_4392,N_3667,N_3023);
and U4393 (N_4393,N_3736,N_3155);
nand U4394 (N_4394,N_3519,N_3531);
and U4395 (N_4395,N_3376,N_3408);
and U4396 (N_4396,N_3363,N_3083);
nand U4397 (N_4397,N_3362,N_3135);
and U4398 (N_4398,N_3201,N_3647);
nand U4399 (N_4399,N_3292,N_3608);
nand U4400 (N_4400,N_3654,N_3167);
and U4401 (N_4401,N_3163,N_3510);
nand U4402 (N_4402,N_3360,N_3400);
nor U4403 (N_4403,N_3309,N_3465);
or U4404 (N_4404,N_3641,N_3206);
and U4405 (N_4405,N_3236,N_3417);
xnor U4406 (N_4406,N_3587,N_3002);
and U4407 (N_4407,N_3460,N_3232);
nand U4408 (N_4408,N_3621,N_3723);
nor U4409 (N_4409,N_3431,N_3236);
and U4410 (N_4410,N_3555,N_3709);
nand U4411 (N_4411,N_3666,N_3255);
or U4412 (N_4412,N_3282,N_3433);
and U4413 (N_4413,N_3267,N_3523);
xnor U4414 (N_4414,N_3366,N_3625);
nor U4415 (N_4415,N_3505,N_3222);
xor U4416 (N_4416,N_3291,N_3679);
and U4417 (N_4417,N_3259,N_3436);
nor U4418 (N_4418,N_3099,N_3037);
nor U4419 (N_4419,N_3547,N_3598);
and U4420 (N_4420,N_3201,N_3711);
nand U4421 (N_4421,N_3656,N_3000);
nand U4422 (N_4422,N_3476,N_3215);
xnor U4423 (N_4423,N_3706,N_3303);
or U4424 (N_4424,N_3632,N_3155);
nand U4425 (N_4425,N_3527,N_3096);
xnor U4426 (N_4426,N_3070,N_3381);
or U4427 (N_4427,N_3478,N_3688);
or U4428 (N_4428,N_3296,N_3124);
or U4429 (N_4429,N_3343,N_3024);
nand U4430 (N_4430,N_3444,N_3230);
and U4431 (N_4431,N_3613,N_3178);
nor U4432 (N_4432,N_3525,N_3404);
nand U4433 (N_4433,N_3304,N_3196);
nor U4434 (N_4434,N_3391,N_3355);
nor U4435 (N_4435,N_3535,N_3078);
and U4436 (N_4436,N_3426,N_3314);
xnor U4437 (N_4437,N_3383,N_3318);
or U4438 (N_4438,N_3651,N_3431);
nand U4439 (N_4439,N_3538,N_3051);
and U4440 (N_4440,N_3414,N_3300);
or U4441 (N_4441,N_3629,N_3262);
nor U4442 (N_4442,N_3476,N_3352);
or U4443 (N_4443,N_3660,N_3351);
xnor U4444 (N_4444,N_3548,N_3149);
nor U4445 (N_4445,N_3131,N_3345);
xnor U4446 (N_4446,N_3512,N_3548);
nor U4447 (N_4447,N_3270,N_3359);
nor U4448 (N_4448,N_3469,N_3418);
and U4449 (N_4449,N_3441,N_3362);
nand U4450 (N_4450,N_3542,N_3170);
nand U4451 (N_4451,N_3441,N_3620);
xor U4452 (N_4452,N_3533,N_3687);
nand U4453 (N_4453,N_3659,N_3214);
nand U4454 (N_4454,N_3039,N_3745);
and U4455 (N_4455,N_3494,N_3150);
and U4456 (N_4456,N_3017,N_3327);
nand U4457 (N_4457,N_3435,N_3347);
or U4458 (N_4458,N_3184,N_3425);
nor U4459 (N_4459,N_3731,N_3139);
nor U4460 (N_4460,N_3448,N_3200);
or U4461 (N_4461,N_3176,N_3017);
and U4462 (N_4462,N_3530,N_3423);
xor U4463 (N_4463,N_3364,N_3467);
or U4464 (N_4464,N_3441,N_3746);
or U4465 (N_4465,N_3035,N_3019);
and U4466 (N_4466,N_3611,N_3218);
nor U4467 (N_4467,N_3174,N_3307);
and U4468 (N_4468,N_3571,N_3105);
nor U4469 (N_4469,N_3091,N_3513);
and U4470 (N_4470,N_3718,N_3162);
nand U4471 (N_4471,N_3547,N_3315);
and U4472 (N_4472,N_3296,N_3546);
or U4473 (N_4473,N_3473,N_3423);
or U4474 (N_4474,N_3033,N_3072);
nor U4475 (N_4475,N_3583,N_3134);
or U4476 (N_4476,N_3224,N_3133);
nand U4477 (N_4477,N_3241,N_3729);
or U4478 (N_4478,N_3359,N_3062);
nor U4479 (N_4479,N_3423,N_3655);
and U4480 (N_4480,N_3016,N_3219);
or U4481 (N_4481,N_3066,N_3310);
or U4482 (N_4482,N_3120,N_3171);
or U4483 (N_4483,N_3460,N_3576);
nor U4484 (N_4484,N_3326,N_3441);
nor U4485 (N_4485,N_3032,N_3003);
or U4486 (N_4486,N_3597,N_3088);
xor U4487 (N_4487,N_3167,N_3741);
nor U4488 (N_4488,N_3122,N_3615);
and U4489 (N_4489,N_3735,N_3062);
and U4490 (N_4490,N_3027,N_3011);
xnor U4491 (N_4491,N_3440,N_3512);
and U4492 (N_4492,N_3054,N_3145);
and U4493 (N_4493,N_3601,N_3591);
nor U4494 (N_4494,N_3223,N_3284);
nand U4495 (N_4495,N_3368,N_3175);
or U4496 (N_4496,N_3346,N_3690);
and U4497 (N_4497,N_3388,N_3633);
nor U4498 (N_4498,N_3654,N_3016);
nor U4499 (N_4499,N_3517,N_3568);
xor U4500 (N_4500,N_4091,N_4263);
xnor U4501 (N_4501,N_4069,N_4259);
or U4502 (N_4502,N_4114,N_3956);
nand U4503 (N_4503,N_4356,N_4206);
and U4504 (N_4504,N_4137,N_4277);
or U4505 (N_4505,N_4116,N_4299);
nor U4506 (N_4506,N_4350,N_4461);
nand U4507 (N_4507,N_4467,N_4032);
nor U4508 (N_4508,N_3883,N_4360);
xor U4509 (N_4509,N_4110,N_3856);
or U4510 (N_4510,N_4216,N_4045);
or U4511 (N_4511,N_4051,N_3797);
nand U4512 (N_4512,N_4125,N_4298);
and U4513 (N_4513,N_3784,N_3820);
or U4514 (N_4514,N_4381,N_3984);
or U4515 (N_4515,N_4014,N_3950);
nand U4516 (N_4516,N_4370,N_4126);
and U4517 (N_4517,N_3949,N_4468);
or U4518 (N_4518,N_4133,N_3848);
nor U4519 (N_4519,N_3943,N_4330);
nor U4520 (N_4520,N_4455,N_4372);
and U4521 (N_4521,N_4113,N_4065);
xnor U4522 (N_4522,N_4096,N_3990);
and U4523 (N_4523,N_4293,N_3807);
nand U4524 (N_4524,N_4084,N_4417);
and U4525 (N_4525,N_4363,N_3855);
or U4526 (N_4526,N_3983,N_4324);
and U4527 (N_4527,N_4477,N_4101);
nor U4528 (N_4528,N_4175,N_3829);
and U4529 (N_4529,N_3846,N_4345);
nor U4530 (N_4530,N_3996,N_4357);
or U4531 (N_4531,N_3877,N_3960);
and U4532 (N_4532,N_3930,N_4451);
or U4533 (N_4533,N_3945,N_4028);
or U4534 (N_4534,N_4108,N_4378);
or U4535 (N_4535,N_4320,N_4024);
nor U4536 (N_4536,N_4435,N_3886);
nand U4537 (N_4537,N_4207,N_4160);
or U4538 (N_4538,N_4465,N_4411);
nand U4539 (N_4539,N_4013,N_4040);
xor U4540 (N_4540,N_4058,N_3934);
or U4541 (N_4541,N_4005,N_4103);
and U4542 (N_4542,N_4280,N_4176);
nand U4543 (N_4543,N_4443,N_4231);
or U4544 (N_4544,N_3852,N_4161);
nor U4545 (N_4545,N_3922,N_3768);
and U4546 (N_4546,N_4427,N_4082);
or U4547 (N_4547,N_4393,N_3968);
nor U4548 (N_4548,N_3867,N_3786);
xnor U4549 (N_4549,N_4106,N_4361);
nor U4550 (N_4550,N_3915,N_4442);
and U4551 (N_4551,N_4166,N_4202);
or U4552 (N_4552,N_4260,N_3840);
nor U4553 (N_4553,N_4197,N_3770);
nor U4554 (N_4554,N_4056,N_3785);
and U4555 (N_4555,N_4047,N_3892);
nand U4556 (N_4556,N_3760,N_4339);
or U4557 (N_4557,N_3917,N_4475);
and U4558 (N_4558,N_3800,N_4218);
or U4559 (N_4559,N_3799,N_4102);
nor U4560 (N_4560,N_4275,N_4156);
or U4561 (N_4561,N_3961,N_3891);
nor U4562 (N_4562,N_4499,N_4018);
and U4563 (N_4563,N_4323,N_4390);
nor U4564 (N_4564,N_4021,N_4376);
xor U4565 (N_4565,N_3788,N_3783);
xor U4566 (N_4566,N_4067,N_4003);
nand U4567 (N_4567,N_4496,N_4145);
nand U4568 (N_4568,N_4262,N_4087);
nand U4569 (N_4569,N_3780,N_4244);
and U4570 (N_4570,N_4124,N_4071);
nand U4571 (N_4571,N_4495,N_3923);
nand U4572 (N_4572,N_3772,N_3890);
or U4573 (N_4573,N_3970,N_3821);
and U4574 (N_4574,N_4335,N_3913);
xnor U4575 (N_4575,N_4046,N_4131);
xnor U4576 (N_4576,N_4235,N_4070);
and U4577 (N_4577,N_4309,N_4303);
nor U4578 (N_4578,N_3878,N_3812);
xnor U4579 (N_4579,N_4478,N_3920);
nand U4580 (N_4580,N_4012,N_4279);
nor U4581 (N_4581,N_4242,N_3773);
and U4582 (N_4582,N_3909,N_3758);
nor U4583 (N_4583,N_4027,N_4385);
and U4584 (N_4584,N_4484,N_4400);
xnor U4585 (N_4585,N_4191,N_4278);
or U4586 (N_4586,N_4301,N_3837);
nand U4587 (N_4587,N_3824,N_3903);
xor U4588 (N_4588,N_4143,N_4413);
nor U4589 (N_4589,N_4266,N_4420);
xnor U4590 (N_4590,N_4450,N_3981);
nor U4591 (N_4591,N_3888,N_4472);
xor U4592 (N_4592,N_4273,N_3759);
nand U4593 (N_4593,N_4437,N_4256);
nor U4594 (N_4594,N_4097,N_4284);
nand U4595 (N_4595,N_3845,N_4407);
and U4596 (N_4596,N_4354,N_4107);
nand U4597 (N_4597,N_4456,N_4147);
and U4598 (N_4598,N_3929,N_4185);
nor U4599 (N_4599,N_4481,N_4367);
nor U4600 (N_4600,N_4352,N_4000);
or U4601 (N_4601,N_4445,N_4122);
or U4602 (N_4602,N_4422,N_3865);
or U4603 (N_4603,N_4016,N_4130);
and U4604 (N_4604,N_3942,N_4482);
nor U4605 (N_4605,N_3982,N_4395);
nand U4606 (N_4606,N_3782,N_4490);
xnor U4607 (N_4607,N_4048,N_4270);
or U4608 (N_4608,N_4285,N_4483);
nand U4609 (N_4609,N_4076,N_4494);
and U4610 (N_4610,N_3889,N_4312);
or U4611 (N_4611,N_3894,N_4469);
xor U4612 (N_4612,N_4038,N_4139);
and U4613 (N_4613,N_3841,N_4193);
nor U4614 (N_4614,N_4199,N_3963);
nand U4615 (N_4615,N_3766,N_3866);
and U4616 (N_4616,N_3904,N_3844);
or U4617 (N_4617,N_4319,N_3809);
nand U4618 (N_4618,N_3816,N_4062);
nand U4619 (N_4619,N_3964,N_3912);
and U4620 (N_4620,N_3972,N_3969);
nor U4621 (N_4621,N_4389,N_4258);
or U4622 (N_4622,N_4135,N_4022);
or U4623 (N_4623,N_4318,N_4264);
or U4624 (N_4624,N_4037,N_4341);
and U4625 (N_4625,N_3937,N_4008);
or U4626 (N_4626,N_4208,N_4210);
nand U4627 (N_4627,N_4406,N_4439);
xnor U4628 (N_4628,N_4396,N_3801);
xnor U4629 (N_4629,N_4409,N_4243);
nand U4630 (N_4630,N_3973,N_4249);
nor U4631 (N_4631,N_4171,N_4486);
nor U4632 (N_4632,N_4222,N_3965);
and U4633 (N_4633,N_4075,N_4054);
nand U4634 (N_4634,N_4230,N_4060);
and U4635 (N_4635,N_4369,N_4158);
nor U4636 (N_4636,N_4492,N_4010);
and U4637 (N_4637,N_4296,N_4433);
nand U4638 (N_4638,N_3872,N_4321);
or U4639 (N_4639,N_3896,N_3815);
nand U4640 (N_4640,N_4192,N_3900);
or U4641 (N_4641,N_3767,N_4431);
and U4642 (N_4642,N_3908,N_3925);
and U4643 (N_4643,N_4276,N_4204);
nor U4644 (N_4644,N_3880,N_4246);
nor U4645 (N_4645,N_3948,N_4112);
and U4646 (N_4646,N_4064,N_4066);
nor U4647 (N_4647,N_4366,N_4448);
xor U4648 (N_4648,N_4059,N_4247);
xnor U4649 (N_4649,N_4043,N_4223);
and U4650 (N_4650,N_4194,N_4009);
and U4651 (N_4651,N_4155,N_4036);
or U4652 (N_4652,N_4085,N_4294);
nor U4653 (N_4653,N_3864,N_4205);
xnor U4654 (N_4654,N_3762,N_4111);
or U4655 (N_4655,N_3971,N_4408);
nand U4656 (N_4656,N_4384,N_4489);
nor U4657 (N_4657,N_4315,N_4311);
nor U4658 (N_4658,N_4209,N_3860);
nor U4659 (N_4659,N_4136,N_4094);
xor U4660 (N_4660,N_3999,N_3881);
xor U4661 (N_4661,N_4117,N_4228);
or U4662 (N_4662,N_3803,N_4078);
nor U4663 (N_4663,N_4295,N_4282);
and U4664 (N_4664,N_4283,N_3755);
or U4665 (N_4665,N_4353,N_4123);
nand U4666 (N_4666,N_3843,N_4358);
nor U4667 (N_4667,N_4470,N_3763);
or U4668 (N_4668,N_4300,N_4304);
nor U4669 (N_4669,N_3933,N_3850);
or U4670 (N_4670,N_4297,N_3980);
and U4671 (N_4671,N_3884,N_4015);
nand U4672 (N_4672,N_3995,N_4307);
nor U4673 (N_4673,N_4154,N_4100);
or U4674 (N_4674,N_4271,N_4498);
nor U4675 (N_4675,N_3796,N_3869);
or U4676 (N_4676,N_4039,N_4041);
and U4677 (N_4677,N_3870,N_4229);
nor U4678 (N_4678,N_4414,N_4394);
nand U4679 (N_4679,N_4310,N_4444);
nand U4680 (N_4680,N_3826,N_3764);
and U4681 (N_4681,N_4379,N_4164);
nor U4682 (N_4682,N_4375,N_3765);
nand U4683 (N_4683,N_4316,N_4265);
and U4684 (N_4684,N_4188,N_3775);
nand U4685 (N_4685,N_3778,N_3931);
nand U4686 (N_4686,N_4343,N_4261);
and U4687 (N_4687,N_4255,N_4401);
nand U4688 (N_4688,N_3862,N_4426);
nand U4689 (N_4689,N_3998,N_3895);
nor U4690 (N_4690,N_4452,N_4364);
or U4691 (N_4691,N_4165,N_4326);
nor U4692 (N_4692,N_4419,N_4157);
and U4693 (N_4693,N_4460,N_4491);
nand U4694 (N_4694,N_4346,N_4250);
nor U4695 (N_4695,N_4134,N_4337);
nand U4696 (N_4696,N_4221,N_4053);
and U4697 (N_4697,N_4425,N_4121);
nand U4698 (N_4698,N_4274,N_3831);
or U4699 (N_4699,N_4172,N_4377);
and U4700 (N_4700,N_3928,N_4415);
nor U4701 (N_4701,N_3919,N_4127);
nor U4702 (N_4702,N_3827,N_4088);
nand U4703 (N_4703,N_3847,N_4286);
and U4704 (N_4704,N_4092,N_4187);
nand U4705 (N_4705,N_3882,N_4371);
or U4706 (N_4706,N_3811,N_4474);
nor U4707 (N_4707,N_4251,N_4440);
or U4708 (N_4708,N_3994,N_3753);
and U4709 (N_4709,N_3805,N_4167);
nor U4710 (N_4710,N_3958,N_4104);
or U4711 (N_4711,N_4220,N_3914);
and U4712 (N_4712,N_3962,N_4386);
or U4713 (N_4713,N_4327,N_4083);
or U4714 (N_4714,N_4291,N_4093);
or U4715 (N_4715,N_4434,N_3750);
and U4716 (N_4716,N_4257,N_4347);
and U4717 (N_4717,N_4140,N_4336);
xor U4718 (N_4718,N_4129,N_3874);
and U4719 (N_4719,N_4359,N_4267);
and U4720 (N_4720,N_3946,N_4203);
nor U4721 (N_4721,N_3823,N_4333);
nor U4722 (N_4722,N_3769,N_3754);
and U4723 (N_4723,N_3863,N_4179);
xnor U4724 (N_4724,N_4063,N_3810);
nand U4725 (N_4725,N_4488,N_4449);
and U4726 (N_4726,N_3898,N_4153);
nor U4727 (N_4727,N_4368,N_4288);
nor U4728 (N_4728,N_4410,N_4428);
nor U4729 (N_4729,N_3926,N_3951);
xnor U4730 (N_4730,N_3795,N_4493);
xnor U4731 (N_4731,N_4219,N_4466);
or U4732 (N_4732,N_3794,N_4141);
xor U4733 (N_4733,N_4355,N_3771);
or U4734 (N_4734,N_3924,N_4035);
nor U4735 (N_4735,N_4162,N_4148);
or U4736 (N_4736,N_3936,N_3781);
nand U4737 (N_4737,N_4446,N_4186);
nand U4738 (N_4738,N_4240,N_4115);
nand U4739 (N_4739,N_3897,N_4052);
nand U4740 (N_4740,N_4030,N_4099);
nor U4741 (N_4741,N_3804,N_4077);
nor U4742 (N_4742,N_4459,N_4365);
or U4743 (N_4743,N_3879,N_4118);
or U4744 (N_4744,N_4429,N_3871);
or U4745 (N_4745,N_4226,N_4019);
and U4746 (N_4746,N_4001,N_4217);
and U4747 (N_4747,N_3836,N_4349);
and U4748 (N_4748,N_3901,N_4138);
and U4749 (N_4749,N_4380,N_4159);
nor U4750 (N_4750,N_3854,N_4306);
or U4751 (N_4751,N_3851,N_3756);
and U4752 (N_4752,N_4334,N_4232);
xnor U4753 (N_4753,N_4373,N_3791);
or U4754 (N_4754,N_4403,N_4269);
nor U4755 (N_4755,N_3830,N_3947);
xor U4756 (N_4756,N_3938,N_4272);
xor U4757 (N_4757,N_4423,N_4342);
or U4758 (N_4758,N_4149,N_4287);
xnor U4759 (N_4759,N_3991,N_3819);
and U4760 (N_4760,N_4402,N_4195);
nor U4761 (N_4761,N_4142,N_4081);
nor U4762 (N_4762,N_3787,N_3828);
nor U4763 (N_4763,N_3779,N_3822);
and U4764 (N_4764,N_3939,N_4464);
or U4765 (N_4765,N_4029,N_3842);
and U4766 (N_4766,N_4447,N_3774);
nand U4767 (N_4767,N_4055,N_4412);
and U4768 (N_4768,N_4338,N_4163);
or U4769 (N_4769,N_3952,N_4201);
and U4770 (N_4770,N_4239,N_3798);
nor U4771 (N_4771,N_4224,N_4453);
nor U4772 (N_4772,N_3911,N_4236);
or U4773 (N_4773,N_4211,N_3959);
nand U4774 (N_4774,N_4438,N_4080);
nor U4775 (N_4775,N_3978,N_4042);
and U4776 (N_4776,N_4214,N_3987);
nor U4777 (N_4777,N_3953,N_4430);
or U4778 (N_4778,N_4432,N_4281);
or U4779 (N_4779,N_4025,N_3988);
or U4780 (N_4780,N_3833,N_3757);
nor U4781 (N_4781,N_4473,N_4184);
and U4782 (N_4782,N_3853,N_3834);
nand U4783 (N_4783,N_4289,N_4462);
nor U4784 (N_4784,N_4322,N_4476);
nand U4785 (N_4785,N_4302,N_4471);
and U4786 (N_4786,N_4314,N_3992);
and U4787 (N_4787,N_3802,N_4196);
nor U4788 (N_4788,N_3954,N_4317);
nor U4789 (N_4789,N_4023,N_4405);
nor U4790 (N_4790,N_4245,N_3868);
nor U4791 (N_4791,N_3885,N_3979);
or U4792 (N_4792,N_4374,N_4248);
xnor U4793 (N_4793,N_4152,N_4180);
nor U4794 (N_4794,N_3825,N_4007);
or U4795 (N_4795,N_4173,N_3887);
nand U4796 (N_4796,N_3777,N_4325);
nor U4797 (N_4797,N_4057,N_3761);
nand U4798 (N_4798,N_4105,N_3817);
and U4799 (N_4799,N_4098,N_4388);
or U4800 (N_4800,N_4458,N_4198);
nor U4801 (N_4801,N_3918,N_4404);
nor U4802 (N_4802,N_3776,N_4313);
and U4803 (N_4803,N_4418,N_4344);
nor U4804 (N_4804,N_4485,N_3905);
nand U4805 (N_4805,N_3997,N_4421);
nand U4806 (N_4806,N_3975,N_4044);
nand U4807 (N_4807,N_3789,N_4268);
and U4808 (N_4808,N_4050,N_4331);
nand U4809 (N_4809,N_4416,N_4169);
xnor U4810 (N_4810,N_4387,N_4308);
nand U4811 (N_4811,N_4190,N_3857);
and U4812 (N_4812,N_4181,N_3893);
nor U4813 (N_4813,N_3916,N_3910);
nand U4814 (N_4814,N_4254,N_3986);
nor U4815 (N_4815,N_4128,N_3835);
or U4816 (N_4816,N_3808,N_4144);
xnor U4817 (N_4817,N_4328,N_3849);
and U4818 (N_4818,N_3838,N_3832);
or U4819 (N_4819,N_4031,N_4150);
xnor U4820 (N_4820,N_3859,N_3993);
nor U4821 (N_4821,N_4183,N_4362);
and U4822 (N_4822,N_4397,N_4200);
or U4823 (N_4823,N_4089,N_4090);
and U4824 (N_4824,N_4120,N_4479);
nor U4825 (N_4825,N_4079,N_4168);
and U4826 (N_4826,N_3977,N_4441);
or U4827 (N_4827,N_3927,N_3957);
nand U4828 (N_4828,N_4463,N_3818);
nor U4829 (N_4829,N_3813,N_3940);
nor U4830 (N_4830,N_4068,N_4329);
or U4831 (N_4831,N_4233,N_4253);
or U4832 (N_4832,N_3806,N_3989);
or U4833 (N_4833,N_4241,N_4424);
nor U4834 (N_4834,N_3752,N_4189);
or U4835 (N_4835,N_4215,N_3941);
and U4836 (N_4836,N_4305,N_4487);
and U4837 (N_4837,N_3932,N_3944);
nor U4838 (N_4838,N_4480,N_4436);
nor U4839 (N_4839,N_4119,N_4017);
nand U4840 (N_4840,N_4170,N_4033);
nor U4841 (N_4841,N_4174,N_3907);
nor U4842 (N_4842,N_4237,N_4132);
nand U4843 (N_4843,N_3955,N_3935);
and U4844 (N_4844,N_4212,N_4011);
xor U4845 (N_4845,N_4061,N_4072);
nand U4846 (N_4846,N_4073,N_4213);
nor U4847 (N_4847,N_3902,N_3985);
nor U4848 (N_4848,N_3899,N_4234);
or U4849 (N_4849,N_3792,N_4497);
and U4850 (N_4850,N_4398,N_4290);
or U4851 (N_4851,N_3875,N_4109);
or U4852 (N_4852,N_3814,N_4348);
nand U4853 (N_4853,N_4457,N_4151);
nor U4854 (N_4854,N_4146,N_4332);
nand U4855 (N_4855,N_4238,N_4382);
nand U4856 (N_4856,N_3873,N_4034);
nor U4857 (N_4857,N_3793,N_4182);
nor U4858 (N_4858,N_4252,N_3790);
nand U4859 (N_4859,N_4340,N_4074);
nand U4860 (N_4860,N_3967,N_3966);
and U4861 (N_4861,N_4383,N_4020);
nand U4862 (N_4862,N_4392,N_3974);
nand U4863 (N_4863,N_4292,N_4391);
or U4864 (N_4864,N_3751,N_3906);
nor U4865 (N_4865,N_4178,N_4095);
nand U4866 (N_4866,N_4351,N_4006);
and U4867 (N_4867,N_4177,N_4086);
nor U4868 (N_4868,N_4227,N_4049);
or U4869 (N_4869,N_3921,N_4454);
nor U4870 (N_4870,N_3839,N_3976);
nand U4871 (N_4871,N_4004,N_3858);
nand U4872 (N_4872,N_4399,N_4002);
nand U4873 (N_4873,N_3861,N_4026);
nand U4874 (N_4874,N_3876,N_4225);
and U4875 (N_4875,N_3870,N_4213);
or U4876 (N_4876,N_4036,N_4316);
nor U4877 (N_4877,N_4074,N_4247);
xor U4878 (N_4878,N_3850,N_4130);
xor U4879 (N_4879,N_3913,N_3802);
or U4880 (N_4880,N_4417,N_3887);
and U4881 (N_4881,N_4381,N_4279);
nand U4882 (N_4882,N_4052,N_4181);
nand U4883 (N_4883,N_4392,N_4471);
or U4884 (N_4884,N_4416,N_3796);
nand U4885 (N_4885,N_3835,N_4202);
or U4886 (N_4886,N_4403,N_3988);
nand U4887 (N_4887,N_3856,N_4267);
nor U4888 (N_4888,N_4189,N_3839);
or U4889 (N_4889,N_4155,N_3870);
or U4890 (N_4890,N_4373,N_4350);
xor U4891 (N_4891,N_4034,N_3915);
nor U4892 (N_4892,N_4186,N_4085);
and U4893 (N_4893,N_4285,N_4389);
nand U4894 (N_4894,N_4271,N_4363);
xnor U4895 (N_4895,N_4222,N_4033);
or U4896 (N_4896,N_3907,N_4142);
nor U4897 (N_4897,N_4388,N_3937);
or U4898 (N_4898,N_4227,N_4272);
or U4899 (N_4899,N_4080,N_4407);
nor U4900 (N_4900,N_3761,N_4496);
and U4901 (N_4901,N_3926,N_3964);
nand U4902 (N_4902,N_3925,N_3795);
or U4903 (N_4903,N_3791,N_3975);
nand U4904 (N_4904,N_4185,N_3955);
nand U4905 (N_4905,N_4038,N_4280);
and U4906 (N_4906,N_3939,N_3836);
nor U4907 (N_4907,N_4461,N_3905);
or U4908 (N_4908,N_3829,N_4255);
or U4909 (N_4909,N_4151,N_3841);
nand U4910 (N_4910,N_3933,N_3908);
or U4911 (N_4911,N_3962,N_3982);
nand U4912 (N_4912,N_4328,N_4199);
nand U4913 (N_4913,N_3782,N_3984);
or U4914 (N_4914,N_3848,N_4141);
and U4915 (N_4915,N_4353,N_4061);
xor U4916 (N_4916,N_4380,N_4364);
and U4917 (N_4917,N_4485,N_4454);
nand U4918 (N_4918,N_3842,N_4465);
and U4919 (N_4919,N_4148,N_4298);
nand U4920 (N_4920,N_3896,N_3823);
or U4921 (N_4921,N_4308,N_4460);
nor U4922 (N_4922,N_3778,N_3943);
or U4923 (N_4923,N_4359,N_4303);
nand U4924 (N_4924,N_4329,N_3794);
nor U4925 (N_4925,N_3799,N_3889);
and U4926 (N_4926,N_4281,N_4111);
or U4927 (N_4927,N_4364,N_4168);
xor U4928 (N_4928,N_4151,N_4286);
and U4929 (N_4929,N_3890,N_4293);
or U4930 (N_4930,N_4322,N_3920);
and U4931 (N_4931,N_3978,N_3865);
or U4932 (N_4932,N_4070,N_3920);
and U4933 (N_4933,N_4379,N_4423);
nand U4934 (N_4934,N_3902,N_4401);
or U4935 (N_4935,N_4186,N_4369);
nor U4936 (N_4936,N_4370,N_3799);
xor U4937 (N_4937,N_3930,N_3820);
and U4938 (N_4938,N_4304,N_4118);
nand U4939 (N_4939,N_4308,N_4234);
and U4940 (N_4940,N_4289,N_4232);
and U4941 (N_4941,N_3867,N_4162);
nand U4942 (N_4942,N_4447,N_3995);
or U4943 (N_4943,N_4095,N_4492);
nor U4944 (N_4944,N_4268,N_3991);
or U4945 (N_4945,N_4162,N_4363);
nor U4946 (N_4946,N_3923,N_4178);
nor U4947 (N_4947,N_3955,N_4368);
nor U4948 (N_4948,N_3786,N_3933);
or U4949 (N_4949,N_3940,N_4483);
nand U4950 (N_4950,N_4217,N_4130);
or U4951 (N_4951,N_4244,N_4033);
and U4952 (N_4952,N_4091,N_4494);
or U4953 (N_4953,N_3965,N_4054);
nor U4954 (N_4954,N_4149,N_4383);
or U4955 (N_4955,N_4190,N_3819);
xnor U4956 (N_4956,N_4031,N_3830);
xor U4957 (N_4957,N_4161,N_4234);
nand U4958 (N_4958,N_3814,N_4242);
or U4959 (N_4959,N_4231,N_4110);
nand U4960 (N_4960,N_4333,N_4401);
nand U4961 (N_4961,N_3772,N_4362);
nand U4962 (N_4962,N_4363,N_4079);
nor U4963 (N_4963,N_4258,N_4157);
xnor U4964 (N_4964,N_3757,N_3896);
and U4965 (N_4965,N_4347,N_4237);
or U4966 (N_4966,N_4280,N_3891);
or U4967 (N_4967,N_4341,N_4414);
nand U4968 (N_4968,N_4028,N_3815);
xnor U4969 (N_4969,N_3786,N_4012);
or U4970 (N_4970,N_4452,N_4080);
nor U4971 (N_4971,N_4369,N_4394);
or U4972 (N_4972,N_4050,N_4340);
nor U4973 (N_4973,N_3831,N_4401);
nand U4974 (N_4974,N_4391,N_3843);
nor U4975 (N_4975,N_4472,N_4227);
nand U4976 (N_4976,N_4438,N_4468);
or U4977 (N_4977,N_4096,N_4037);
nor U4978 (N_4978,N_4178,N_4324);
xnor U4979 (N_4979,N_4159,N_3894);
or U4980 (N_4980,N_4130,N_3841);
and U4981 (N_4981,N_4442,N_4367);
nor U4982 (N_4982,N_4337,N_4315);
and U4983 (N_4983,N_4178,N_4018);
and U4984 (N_4984,N_3812,N_3868);
nor U4985 (N_4985,N_4266,N_4281);
or U4986 (N_4986,N_4210,N_4276);
and U4987 (N_4987,N_4134,N_3837);
nor U4988 (N_4988,N_3773,N_4478);
nor U4989 (N_4989,N_4129,N_4371);
xnor U4990 (N_4990,N_4038,N_4281);
xor U4991 (N_4991,N_4149,N_4197);
and U4992 (N_4992,N_3913,N_4457);
and U4993 (N_4993,N_3865,N_4248);
and U4994 (N_4994,N_4040,N_3953);
and U4995 (N_4995,N_4491,N_3861);
nor U4996 (N_4996,N_4488,N_4105);
nand U4997 (N_4997,N_4462,N_4219);
and U4998 (N_4998,N_3882,N_4409);
nor U4999 (N_4999,N_4172,N_3772);
nand U5000 (N_5000,N_4436,N_4091);
and U5001 (N_5001,N_4295,N_4353);
or U5002 (N_5002,N_4347,N_4081);
nor U5003 (N_5003,N_4491,N_3871);
and U5004 (N_5004,N_4487,N_4107);
nor U5005 (N_5005,N_3866,N_3907);
xor U5006 (N_5006,N_4290,N_4432);
or U5007 (N_5007,N_4101,N_4440);
nor U5008 (N_5008,N_3837,N_4054);
nand U5009 (N_5009,N_4442,N_4168);
and U5010 (N_5010,N_3997,N_4042);
and U5011 (N_5011,N_3798,N_4156);
nand U5012 (N_5012,N_4426,N_4396);
nand U5013 (N_5013,N_4008,N_4042);
nand U5014 (N_5014,N_4449,N_4408);
nand U5015 (N_5015,N_4381,N_3809);
nand U5016 (N_5016,N_3918,N_4474);
or U5017 (N_5017,N_4136,N_4269);
or U5018 (N_5018,N_4108,N_3973);
nor U5019 (N_5019,N_3813,N_4301);
xor U5020 (N_5020,N_3849,N_4009);
or U5021 (N_5021,N_3871,N_4063);
nor U5022 (N_5022,N_4320,N_4161);
nand U5023 (N_5023,N_4330,N_4025);
nor U5024 (N_5024,N_4003,N_4163);
nand U5025 (N_5025,N_4251,N_4487);
or U5026 (N_5026,N_3771,N_4332);
nor U5027 (N_5027,N_4283,N_4377);
and U5028 (N_5028,N_4030,N_3849);
nor U5029 (N_5029,N_4473,N_3970);
xor U5030 (N_5030,N_4226,N_4415);
nor U5031 (N_5031,N_3870,N_4120);
and U5032 (N_5032,N_4156,N_4024);
or U5033 (N_5033,N_4118,N_4382);
and U5034 (N_5034,N_3803,N_4208);
and U5035 (N_5035,N_4488,N_4382);
xor U5036 (N_5036,N_3849,N_3816);
and U5037 (N_5037,N_4087,N_3763);
or U5038 (N_5038,N_4304,N_4342);
nand U5039 (N_5039,N_4380,N_4265);
nor U5040 (N_5040,N_4176,N_4103);
nand U5041 (N_5041,N_4429,N_4101);
nand U5042 (N_5042,N_3778,N_4322);
or U5043 (N_5043,N_4201,N_3877);
nor U5044 (N_5044,N_4225,N_3813);
or U5045 (N_5045,N_4106,N_3935);
and U5046 (N_5046,N_4492,N_3774);
and U5047 (N_5047,N_4110,N_4270);
or U5048 (N_5048,N_3877,N_4340);
nand U5049 (N_5049,N_4100,N_3797);
nand U5050 (N_5050,N_4035,N_3968);
nand U5051 (N_5051,N_4040,N_3811);
nor U5052 (N_5052,N_4189,N_4227);
xor U5053 (N_5053,N_4322,N_4271);
and U5054 (N_5054,N_4153,N_4294);
and U5055 (N_5055,N_4331,N_4310);
nor U5056 (N_5056,N_4249,N_4029);
and U5057 (N_5057,N_4459,N_4441);
nor U5058 (N_5058,N_4263,N_4088);
and U5059 (N_5059,N_3792,N_4262);
nand U5060 (N_5060,N_4009,N_3860);
nor U5061 (N_5061,N_4140,N_4163);
and U5062 (N_5062,N_4455,N_4244);
xnor U5063 (N_5063,N_4051,N_4300);
and U5064 (N_5064,N_3809,N_4393);
nor U5065 (N_5065,N_4458,N_4097);
nor U5066 (N_5066,N_3907,N_4050);
nand U5067 (N_5067,N_3774,N_4180);
or U5068 (N_5068,N_3860,N_4059);
and U5069 (N_5069,N_4306,N_3803);
or U5070 (N_5070,N_4115,N_4221);
nor U5071 (N_5071,N_4446,N_4033);
or U5072 (N_5072,N_4461,N_4275);
nand U5073 (N_5073,N_4284,N_3846);
nor U5074 (N_5074,N_4321,N_3815);
nand U5075 (N_5075,N_4376,N_4227);
and U5076 (N_5076,N_3870,N_4349);
and U5077 (N_5077,N_4160,N_4420);
nand U5078 (N_5078,N_3785,N_4493);
xor U5079 (N_5079,N_4033,N_4277);
or U5080 (N_5080,N_4403,N_3874);
xor U5081 (N_5081,N_4299,N_4119);
or U5082 (N_5082,N_3754,N_4006);
and U5083 (N_5083,N_4271,N_3949);
xor U5084 (N_5084,N_3770,N_4382);
nor U5085 (N_5085,N_3944,N_4475);
or U5086 (N_5086,N_4052,N_3812);
or U5087 (N_5087,N_4148,N_3936);
nand U5088 (N_5088,N_4129,N_4374);
or U5089 (N_5089,N_4141,N_3859);
nor U5090 (N_5090,N_4406,N_4385);
nor U5091 (N_5091,N_4313,N_4478);
and U5092 (N_5092,N_4070,N_3821);
xnor U5093 (N_5093,N_4431,N_4332);
or U5094 (N_5094,N_3801,N_4495);
xor U5095 (N_5095,N_3897,N_3752);
and U5096 (N_5096,N_3968,N_4396);
nor U5097 (N_5097,N_4177,N_4374);
and U5098 (N_5098,N_4191,N_3755);
or U5099 (N_5099,N_3898,N_4029);
or U5100 (N_5100,N_3828,N_3954);
and U5101 (N_5101,N_4460,N_4242);
nand U5102 (N_5102,N_3814,N_4070);
or U5103 (N_5103,N_4381,N_3907);
nor U5104 (N_5104,N_4302,N_3771);
or U5105 (N_5105,N_4156,N_4442);
nand U5106 (N_5106,N_4160,N_3930);
and U5107 (N_5107,N_3806,N_4281);
nor U5108 (N_5108,N_4333,N_3890);
or U5109 (N_5109,N_3961,N_4479);
nor U5110 (N_5110,N_4075,N_3866);
nand U5111 (N_5111,N_4313,N_3837);
and U5112 (N_5112,N_3844,N_4435);
nor U5113 (N_5113,N_4321,N_4225);
nor U5114 (N_5114,N_4129,N_3888);
and U5115 (N_5115,N_3884,N_4461);
and U5116 (N_5116,N_4035,N_3810);
nand U5117 (N_5117,N_3907,N_4358);
or U5118 (N_5118,N_4433,N_4156);
nor U5119 (N_5119,N_3789,N_4031);
or U5120 (N_5120,N_4333,N_4115);
nor U5121 (N_5121,N_4314,N_4373);
or U5122 (N_5122,N_4302,N_4167);
nand U5123 (N_5123,N_4486,N_4252);
and U5124 (N_5124,N_3931,N_3932);
nor U5125 (N_5125,N_4349,N_4363);
and U5126 (N_5126,N_3994,N_4402);
and U5127 (N_5127,N_3784,N_4230);
and U5128 (N_5128,N_4394,N_4365);
and U5129 (N_5129,N_4009,N_4484);
nand U5130 (N_5130,N_3806,N_4183);
or U5131 (N_5131,N_3783,N_4270);
nand U5132 (N_5132,N_4488,N_4012);
or U5133 (N_5133,N_4459,N_4234);
nand U5134 (N_5134,N_3946,N_4133);
nand U5135 (N_5135,N_4458,N_3860);
or U5136 (N_5136,N_3896,N_4458);
or U5137 (N_5137,N_4193,N_4278);
nor U5138 (N_5138,N_4321,N_4106);
nor U5139 (N_5139,N_3993,N_4063);
and U5140 (N_5140,N_4303,N_4485);
and U5141 (N_5141,N_3759,N_4065);
or U5142 (N_5142,N_4062,N_3783);
nand U5143 (N_5143,N_4265,N_3945);
or U5144 (N_5144,N_4086,N_4029);
or U5145 (N_5145,N_3820,N_3875);
or U5146 (N_5146,N_4289,N_4338);
nand U5147 (N_5147,N_4361,N_4365);
and U5148 (N_5148,N_3805,N_3966);
or U5149 (N_5149,N_4346,N_4499);
or U5150 (N_5150,N_3805,N_4090);
and U5151 (N_5151,N_4030,N_4375);
nand U5152 (N_5152,N_4348,N_4339);
nand U5153 (N_5153,N_3774,N_4254);
or U5154 (N_5154,N_3809,N_4469);
and U5155 (N_5155,N_3771,N_3993);
and U5156 (N_5156,N_4306,N_4248);
or U5157 (N_5157,N_3901,N_4036);
nor U5158 (N_5158,N_4474,N_4093);
and U5159 (N_5159,N_4124,N_4488);
or U5160 (N_5160,N_4013,N_4009);
xor U5161 (N_5161,N_3940,N_4148);
nand U5162 (N_5162,N_4291,N_3868);
and U5163 (N_5163,N_3792,N_4369);
xor U5164 (N_5164,N_4229,N_3864);
and U5165 (N_5165,N_4279,N_4264);
xor U5166 (N_5166,N_3832,N_4270);
nor U5167 (N_5167,N_4462,N_4281);
or U5168 (N_5168,N_4222,N_4447);
nand U5169 (N_5169,N_3999,N_3910);
or U5170 (N_5170,N_4401,N_4197);
and U5171 (N_5171,N_4350,N_4297);
nand U5172 (N_5172,N_3806,N_3996);
or U5173 (N_5173,N_3894,N_4447);
and U5174 (N_5174,N_4246,N_3870);
nand U5175 (N_5175,N_4326,N_4063);
xor U5176 (N_5176,N_4483,N_3949);
nand U5177 (N_5177,N_3863,N_3818);
or U5178 (N_5178,N_4202,N_4216);
or U5179 (N_5179,N_4120,N_4323);
nor U5180 (N_5180,N_4124,N_4088);
and U5181 (N_5181,N_4231,N_4402);
nand U5182 (N_5182,N_4024,N_4387);
xnor U5183 (N_5183,N_4429,N_4001);
xnor U5184 (N_5184,N_4052,N_4186);
nand U5185 (N_5185,N_3813,N_4016);
and U5186 (N_5186,N_3962,N_4164);
nor U5187 (N_5187,N_4079,N_3881);
or U5188 (N_5188,N_4024,N_4332);
nor U5189 (N_5189,N_3785,N_4331);
nand U5190 (N_5190,N_3764,N_4108);
or U5191 (N_5191,N_4171,N_3911);
nand U5192 (N_5192,N_4364,N_4429);
nand U5193 (N_5193,N_4261,N_4000);
or U5194 (N_5194,N_4276,N_4089);
or U5195 (N_5195,N_4183,N_4162);
or U5196 (N_5196,N_3846,N_4029);
nand U5197 (N_5197,N_3874,N_3829);
and U5198 (N_5198,N_3880,N_3929);
or U5199 (N_5199,N_4271,N_3829);
or U5200 (N_5200,N_4352,N_4234);
and U5201 (N_5201,N_3997,N_4473);
nand U5202 (N_5202,N_4323,N_3943);
or U5203 (N_5203,N_4315,N_4303);
nand U5204 (N_5204,N_4459,N_4035);
and U5205 (N_5205,N_4044,N_4328);
nand U5206 (N_5206,N_3945,N_3779);
nor U5207 (N_5207,N_4172,N_4276);
nor U5208 (N_5208,N_3800,N_4034);
nor U5209 (N_5209,N_4231,N_3919);
and U5210 (N_5210,N_4473,N_4276);
nand U5211 (N_5211,N_3994,N_4091);
and U5212 (N_5212,N_4122,N_4361);
nor U5213 (N_5213,N_3943,N_4012);
nand U5214 (N_5214,N_4297,N_4378);
xor U5215 (N_5215,N_3964,N_4022);
nor U5216 (N_5216,N_4257,N_3823);
or U5217 (N_5217,N_4458,N_4432);
and U5218 (N_5218,N_3856,N_4331);
nor U5219 (N_5219,N_4047,N_4144);
or U5220 (N_5220,N_4191,N_4346);
or U5221 (N_5221,N_3936,N_4365);
xor U5222 (N_5222,N_4165,N_4161);
nand U5223 (N_5223,N_4444,N_4098);
or U5224 (N_5224,N_3848,N_4198);
nor U5225 (N_5225,N_4054,N_4280);
nand U5226 (N_5226,N_4463,N_4231);
and U5227 (N_5227,N_4117,N_3867);
nand U5228 (N_5228,N_4488,N_4378);
nor U5229 (N_5229,N_3930,N_4197);
or U5230 (N_5230,N_4381,N_4379);
nor U5231 (N_5231,N_4312,N_3848);
nand U5232 (N_5232,N_4402,N_3977);
nor U5233 (N_5233,N_4301,N_4330);
or U5234 (N_5234,N_4413,N_4067);
nand U5235 (N_5235,N_4306,N_4424);
nand U5236 (N_5236,N_3909,N_4317);
or U5237 (N_5237,N_4257,N_3753);
nand U5238 (N_5238,N_4058,N_3881);
nor U5239 (N_5239,N_4012,N_4157);
and U5240 (N_5240,N_4492,N_3989);
and U5241 (N_5241,N_4288,N_4207);
nand U5242 (N_5242,N_4209,N_4103);
and U5243 (N_5243,N_3808,N_4046);
or U5244 (N_5244,N_3835,N_3981);
xnor U5245 (N_5245,N_4208,N_4249);
or U5246 (N_5246,N_4135,N_4066);
nand U5247 (N_5247,N_4434,N_4003);
nand U5248 (N_5248,N_3779,N_4410);
nor U5249 (N_5249,N_4158,N_3757);
nand U5250 (N_5250,N_5093,N_4649);
or U5251 (N_5251,N_5085,N_5145);
nor U5252 (N_5252,N_5244,N_5177);
and U5253 (N_5253,N_4863,N_4787);
xor U5254 (N_5254,N_4893,N_4883);
nand U5255 (N_5255,N_5105,N_4662);
nand U5256 (N_5256,N_4786,N_5028);
nand U5257 (N_5257,N_5080,N_4792);
nand U5258 (N_5258,N_4679,N_4978);
xor U5259 (N_5259,N_4602,N_5233);
and U5260 (N_5260,N_4714,N_4551);
nand U5261 (N_5261,N_4847,N_4811);
or U5262 (N_5262,N_4754,N_5224);
nor U5263 (N_5263,N_5181,N_4830);
nor U5264 (N_5264,N_4976,N_4848);
or U5265 (N_5265,N_5202,N_5126);
xnor U5266 (N_5266,N_5000,N_4937);
or U5267 (N_5267,N_4755,N_5217);
and U5268 (N_5268,N_5055,N_5130);
nand U5269 (N_5269,N_4885,N_5061);
nor U5270 (N_5270,N_5231,N_4702);
xor U5271 (N_5271,N_4957,N_5109);
nor U5272 (N_5272,N_4985,N_4851);
and U5273 (N_5273,N_4750,N_4615);
and U5274 (N_5274,N_4505,N_5178);
or U5275 (N_5275,N_5154,N_4833);
nand U5276 (N_5276,N_5021,N_4772);
nor U5277 (N_5277,N_4585,N_4546);
xor U5278 (N_5278,N_4928,N_5161);
nor U5279 (N_5279,N_5186,N_4645);
nand U5280 (N_5280,N_5236,N_4866);
and U5281 (N_5281,N_4577,N_4640);
nand U5282 (N_5282,N_4869,N_4859);
and U5283 (N_5283,N_4538,N_4554);
xnor U5284 (N_5284,N_5087,N_5192);
nand U5285 (N_5285,N_5103,N_5114);
and U5286 (N_5286,N_4979,N_4593);
and U5287 (N_5287,N_4823,N_5171);
and U5288 (N_5288,N_5229,N_4803);
and U5289 (N_5289,N_4761,N_5019);
and U5290 (N_5290,N_4712,N_5232);
and U5291 (N_5291,N_5249,N_4718);
nand U5292 (N_5292,N_4793,N_4951);
xnor U5293 (N_5293,N_4599,N_4561);
nor U5294 (N_5294,N_4882,N_4743);
and U5295 (N_5295,N_4832,N_5104);
nand U5296 (N_5296,N_4828,N_4727);
nor U5297 (N_5297,N_5013,N_5043);
nand U5298 (N_5298,N_4661,N_5039);
or U5299 (N_5299,N_5089,N_4784);
nor U5300 (N_5300,N_5174,N_4619);
or U5301 (N_5301,N_4710,N_4766);
nor U5302 (N_5302,N_4958,N_4708);
nand U5303 (N_5303,N_4545,N_4603);
and U5304 (N_5304,N_4665,N_5107);
nand U5305 (N_5305,N_5110,N_4650);
and U5306 (N_5306,N_5245,N_4625);
or U5307 (N_5307,N_4565,N_4687);
nand U5308 (N_5308,N_5094,N_4604);
or U5309 (N_5309,N_5123,N_4524);
nor U5310 (N_5310,N_4699,N_5041);
nand U5311 (N_5311,N_4941,N_4527);
xor U5312 (N_5312,N_4628,N_4808);
nand U5313 (N_5313,N_4529,N_4557);
or U5314 (N_5314,N_5033,N_4873);
and U5315 (N_5315,N_4807,N_4525);
nor U5316 (N_5316,N_4587,N_4919);
or U5317 (N_5317,N_4876,N_4659);
or U5318 (N_5318,N_5050,N_4510);
nand U5319 (N_5319,N_4654,N_4838);
or U5320 (N_5320,N_4757,N_5158);
xor U5321 (N_5321,N_4630,N_4889);
xor U5322 (N_5322,N_5184,N_5149);
and U5323 (N_5323,N_5111,N_4922);
nor U5324 (N_5324,N_4675,N_4553);
and U5325 (N_5325,N_4530,N_4735);
xnor U5326 (N_5326,N_4589,N_5182);
and U5327 (N_5327,N_4834,N_4762);
or U5328 (N_5328,N_4981,N_5185);
and U5329 (N_5329,N_4558,N_4858);
or U5330 (N_5330,N_4908,N_5163);
nand U5331 (N_5331,N_4738,N_4920);
xor U5332 (N_5332,N_4533,N_5214);
nor U5333 (N_5333,N_5137,N_5034);
and U5334 (N_5334,N_4897,N_4657);
or U5335 (N_5335,N_4877,N_5201);
nand U5336 (N_5336,N_4730,N_5120);
and U5337 (N_5337,N_4517,N_4955);
or U5338 (N_5338,N_4676,N_4733);
or U5339 (N_5339,N_5065,N_5219);
or U5340 (N_5340,N_4925,N_5006);
or U5341 (N_5341,N_5070,N_4870);
xor U5342 (N_5342,N_4670,N_4686);
and U5343 (N_5343,N_4963,N_4570);
nor U5344 (N_5344,N_4668,N_5213);
nor U5345 (N_5345,N_5025,N_4672);
nand U5346 (N_5346,N_5058,N_4671);
xor U5347 (N_5347,N_4911,N_4501);
and U5348 (N_5348,N_4669,N_4698);
and U5349 (N_5349,N_4655,N_4658);
and U5350 (N_5350,N_5228,N_4809);
nor U5351 (N_5351,N_5082,N_4818);
xor U5352 (N_5352,N_5012,N_4915);
or U5353 (N_5353,N_4987,N_4998);
nand U5354 (N_5354,N_4566,N_4704);
and U5355 (N_5355,N_5227,N_4875);
or U5356 (N_5356,N_5124,N_4612);
nand U5357 (N_5357,N_4597,N_4990);
and U5358 (N_5358,N_4513,N_4696);
nand U5359 (N_5359,N_4713,N_4556);
nand U5360 (N_5360,N_4917,N_4532);
nor U5361 (N_5361,N_4562,N_4868);
or U5362 (N_5362,N_4732,N_4636);
and U5363 (N_5363,N_4716,N_4829);
or U5364 (N_5364,N_4947,N_4855);
nor U5365 (N_5365,N_5079,N_4550);
xor U5366 (N_5366,N_4503,N_5016);
or U5367 (N_5367,N_4933,N_4779);
nor U5368 (N_5368,N_4506,N_4845);
and U5369 (N_5369,N_4902,N_5125);
nand U5370 (N_5370,N_5169,N_4826);
and U5371 (N_5371,N_5135,N_4707);
nor U5372 (N_5372,N_4664,N_5086);
and U5373 (N_5373,N_5153,N_4610);
nand U5374 (N_5374,N_4663,N_4996);
nor U5375 (N_5375,N_4681,N_5064);
or U5376 (N_5376,N_4886,N_4697);
nor U5377 (N_5377,N_4888,N_4986);
nand U5378 (N_5378,N_5044,N_5196);
nand U5379 (N_5379,N_4677,N_4541);
nor U5380 (N_5380,N_4746,N_4703);
nand U5381 (N_5381,N_4961,N_4680);
nand U5382 (N_5382,N_4880,N_4542);
nand U5383 (N_5383,N_4741,N_5239);
nand U5384 (N_5384,N_5084,N_4798);
or U5385 (N_5385,N_5066,N_5248);
and U5386 (N_5386,N_4683,N_4991);
nand U5387 (N_5387,N_4817,N_5009);
nand U5388 (N_5388,N_4934,N_4853);
nor U5389 (N_5389,N_5129,N_4906);
nor U5390 (N_5390,N_4972,N_4690);
or U5391 (N_5391,N_4768,N_5099);
nor U5392 (N_5392,N_4637,N_4782);
nor U5393 (N_5393,N_4865,N_4765);
nor U5394 (N_5394,N_5029,N_4926);
or U5395 (N_5395,N_4598,N_5203);
xnor U5396 (N_5396,N_5083,N_4887);
and U5397 (N_5397,N_5096,N_4842);
nor U5398 (N_5398,N_4794,N_5197);
and U5399 (N_5399,N_4776,N_4992);
nand U5400 (N_5400,N_4778,N_5140);
nand U5401 (N_5401,N_4652,N_5001);
xor U5402 (N_5402,N_4620,N_4688);
or U5403 (N_5403,N_4999,N_4583);
nor U5404 (N_5404,N_4810,N_4907);
nor U5405 (N_5405,N_5116,N_4753);
xor U5406 (N_5406,N_5026,N_5020);
nand U5407 (N_5407,N_4744,N_5180);
or U5408 (N_5408,N_4959,N_4952);
or U5409 (N_5409,N_4927,N_5212);
nor U5410 (N_5410,N_4633,N_4564);
nor U5411 (N_5411,N_4780,N_4500);
or U5412 (N_5412,N_5030,N_5024);
nor U5413 (N_5413,N_4745,N_4594);
nor U5414 (N_5414,N_5225,N_5234);
nor U5415 (N_5415,N_4984,N_4938);
nand U5416 (N_5416,N_4725,N_4944);
and U5417 (N_5417,N_4854,N_5139);
or U5418 (N_5418,N_4930,N_4783);
or U5419 (N_5419,N_4518,N_4997);
or U5420 (N_5420,N_4841,N_4967);
nor U5421 (N_5421,N_5115,N_4534);
and U5422 (N_5422,N_4606,N_4942);
xnor U5423 (N_5423,N_4820,N_4837);
nand U5424 (N_5424,N_4685,N_4509);
or U5425 (N_5425,N_4971,N_4616);
nand U5426 (N_5426,N_4918,N_4970);
or U5427 (N_5427,N_4571,N_4643);
and U5428 (N_5428,N_4624,N_5146);
and U5429 (N_5429,N_4588,N_4720);
and U5430 (N_5430,N_4579,N_4791);
nand U5431 (N_5431,N_5068,N_4711);
nor U5432 (N_5432,N_5143,N_4614);
nor U5433 (N_5433,N_4578,N_5207);
nand U5434 (N_5434,N_5208,N_4852);
nor U5435 (N_5435,N_4945,N_5052);
and U5436 (N_5436,N_4507,N_5031);
nand U5437 (N_5437,N_4993,N_4567);
xnor U5438 (N_5438,N_4722,N_4822);
nand U5439 (N_5439,N_4804,N_5168);
or U5440 (N_5440,N_5101,N_5241);
nand U5441 (N_5441,N_4795,N_4943);
or U5442 (N_5442,N_4627,N_4969);
and U5443 (N_5443,N_4890,N_4694);
nand U5444 (N_5444,N_5007,N_4693);
nor U5445 (N_5445,N_4805,N_4871);
nand U5446 (N_5446,N_4872,N_5054);
nor U5447 (N_5447,N_4789,N_4512);
and U5448 (N_5448,N_4572,N_4523);
nor U5449 (N_5449,N_4673,N_4946);
nand U5450 (N_5450,N_4611,N_4609);
and U5451 (N_5451,N_5148,N_4773);
nor U5452 (N_5452,N_4796,N_4800);
or U5453 (N_5453,N_5136,N_4935);
nand U5454 (N_5454,N_4514,N_4899);
nand U5455 (N_5455,N_5157,N_5022);
and U5456 (N_5456,N_5060,N_4980);
or U5457 (N_5457,N_5183,N_4641);
and U5458 (N_5458,N_4896,N_4856);
or U5459 (N_5459,N_5206,N_4528);
nand U5460 (N_5460,N_4774,N_5069);
or U5461 (N_5461,N_4892,N_4747);
and U5462 (N_5462,N_4644,N_4715);
or U5463 (N_5463,N_5195,N_4502);
and U5464 (N_5464,N_5073,N_5121);
nor U5465 (N_5465,N_4758,N_4831);
nand U5466 (N_5466,N_5076,N_4543);
nand U5467 (N_5467,N_5205,N_5191);
or U5468 (N_5468,N_5040,N_4634);
and U5469 (N_5469,N_5072,N_4642);
and U5470 (N_5470,N_4751,N_5199);
nor U5471 (N_5471,N_4717,N_5200);
nor U5472 (N_5472,N_5223,N_4989);
nand U5473 (N_5473,N_4660,N_5100);
nor U5474 (N_5474,N_5209,N_4575);
or U5475 (N_5475,N_5023,N_4618);
nand U5476 (N_5476,N_5047,N_4901);
nand U5477 (N_5477,N_5098,N_4891);
and U5478 (N_5478,N_5008,N_4520);
or U5479 (N_5479,N_5071,N_5091);
and U5480 (N_5480,N_4850,N_5048);
or U5481 (N_5481,N_5077,N_4656);
nor U5482 (N_5482,N_5141,N_4522);
nor U5483 (N_5483,N_4909,N_4843);
nand U5484 (N_5484,N_5147,N_4622);
nand U5485 (N_5485,N_4816,N_4736);
xor U5486 (N_5486,N_4626,N_5015);
or U5487 (N_5487,N_5122,N_4595);
nand U5488 (N_5488,N_4540,N_4949);
nor U5489 (N_5489,N_4860,N_4812);
nor U5490 (N_5490,N_5106,N_4775);
nand U5491 (N_5491,N_5002,N_4894);
nor U5492 (N_5492,N_4824,N_4839);
nand U5493 (N_5493,N_4536,N_4623);
nor U5494 (N_5494,N_4874,N_4785);
nor U5495 (N_5495,N_5193,N_4573);
or U5496 (N_5496,N_5198,N_5059);
and U5497 (N_5497,N_4539,N_4849);
and U5498 (N_5498,N_5003,N_5018);
nor U5499 (N_5499,N_5210,N_5051);
nor U5500 (N_5500,N_4988,N_4621);
and U5501 (N_5501,N_4912,N_4548);
xnor U5502 (N_5502,N_5092,N_4764);
nor U5503 (N_5503,N_4631,N_5165);
or U5504 (N_5504,N_4608,N_4726);
nand U5505 (N_5505,N_4881,N_4576);
nor U5506 (N_5506,N_4596,N_5056);
and U5507 (N_5507,N_4983,N_4519);
xor U5508 (N_5508,N_5194,N_4709);
nand U5509 (N_5509,N_4760,N_4749);
nand U5510 (N_5510,N_4613,N_5032);
or U5511 (N_5511,N_5216,N_4884);
nand U5512 (N_5512,N_4695,N_4815);
and U5513 (N_5513,N_4790,N_4799);
nor U5514 (N_5514,N_4737,N_5150);
and U5515 (N_5515,N_5211,N_4974);
or U5516 (N_5516,N_4878,N_4975);
nor U5517 (N_5517,N_4691,N_4777);
nor U5518 (N_5518,N_5176,N_5247);
and U5519 (N_5519,N_4844,N_4605);
nand U5520 (N_5520,N_5238,N_5246);
xnor U5521 (N_5521,N_4728,N_5004);
and U5522 (N_5522,N_4939,N_5243);
or U5523 (N_5523,N_4705,N_4569);
xnor U5524 (N_5524,N_4977,N_5166);
nand U5525 (N_5525,N_4948,N_4580);
and U5526 (N_5526,N_5117,N_5189);
nor U5527 (N_5527,N_5190,N_4617);
xnor U5528 (N_5528,N_5172,N_4929);
and U5529 (N_5529,N_4752,N_4742);
nor U5530 (N_5530,N_4821,N_4653);
and U5531 (N_5531,N_5220,N_5128);
or U5532 (N_5532,N_5011,N_5160);
xnor U5533 (N_5533,N_5159,N_5187);
xor U5534 (N_5534,N_4504,N_4574);
and U5535 (N_5535,N_4731,N_4801);
and U5536 (N_5536,N_5074,N_4590);
nor U5537 (N_5537,N_4916,N_4802);
nand U5538 (N_5538,N_4584,N_5118);
and U5539 (N_5539,N_4684,N_4770);
or U5540 (N_5540,N_5152,N_4682);
nand U5541 (N_5541,N_5155,N_5215);
or U5542 (N_5542,N_4692,N_5037);
nor U5543 (N_5543,N_4813,N_5167);
nor U5544 (N_5544,N_4537,N_4535);
or U5545 (N_5545,N_4763,N_5067);
xnor U5546 (N_5546,N_5088,N_5188);
xor U5547 (N_5547,N_4632,N_5131);
or U5548 (N_5548,N_4648,N_5046);
nor U5549 (N_5549,N_4835,N_5063);
nand U5550 (N_5550,N_5042,N_4953);
and U5551 (N_5551,N_4769,N_5133);
and U5552 (N_5552,N_4547,N_4936);
and U5553 (N_5553,N_5035,N_4995);
nor U5554 (N_5554,N_4582,N_5038);
and U5555 (N_5555,N_4638,N_4559);
nor U5556 (N_5556,N_4739,N_4544);
nor U5557 (N_5557,N_4965,N_4968);
or U5558 (N_5558,N_4910,N_5017);
nand U5559 (N_5559,N_5112,N_5132);
nor U5560 (N_5560,N_4563,N_4788);
nand U5561 (N_5561,N_4857,N_5162);
nor U5562 (N_5562,N_4740,N_4706);
or U5563 (N_5563,N_5078,N_4607);
and U5564 (N_5564,N_4667,N_4827);
or U5565 (N_5565,N_5173,N_5053);
xor U5566 (N_5566,N_4973,N_4771);
nor U5567 (N_5567,N_5156,N_5144);
nor U5568 (N_5568,N_5075,N_4966);
nor U5569 (N_5569,N_5010,N_4862);
or U5570 (N_5570,N_4600,N_5235);
nor U5571 (N_5571,N_4861,N_4552);
or U5572 (N_5572,N_5138,N_4560);
nand U5573 (N_5573,N_4629,N_4836);
nand U5574 (N_5574,N_4982,N_4962);
and U5575 (N_5575,N_5134,N_4921);
and U5576 (N_5576,N_5049,N_4521);
and U5577 (N_5577,N_5218,N_4734);
or U5578 (N_5578,N_4914,N_4964);
nand U5579 (N_5579,N_5036,N_5142);
and U5580 (N_5580,N_4960,N_4903);
and U5581 (N_5581,N_4729,N_4592);
nor U5582 (N_5582,N_5170,N_4719);
nand U5583 (N_5583,N_4581,N_4549);
or U5584 (N_5584,N_5119,N_4950);
xor U5585 (N_5585,N_4864,N_4879);
nand U5586 (N_5586,N_4825,N_5151);
or U5587 (N_5587,N_4806,N_4956);
nor U5588 (N_5588,N_4531,N_4904);
or U5589 (N_5589,N_4924,N_5242);
or U5590 (N_5590,N_5045,N_4840);
or U5591 (N_5591,N_4767,N_4900);
nand U5592 (N_5592,N_5081,N_4701);
xor U5593 (N_5593,N_4721,N_5230);
nand U5594 (N_5594,N_4689,N_4568);
nor U5595 (N_5595,N_4700,N_4932);
or U5596 (N_5596,N_4913,N_4678);
nand U5597 (N_5597,N_4666,N_4905);
nor U5598 (N_5598,N_5127,N_5237);
nor U5599 (N_5599,N_4555,N_4635);
nor U5600 (N_5600,N_4867,N_4846);
or U5601 (N_5601,N_4797,N_4586);
or U5602 (N_5602,N_4646,N_5095);
and U5603 (N_5603,N_4748,N_5027);
xnor U5604 (N_5604,N_5240,N_4923);
nor U5605 (N_5605,N_4651,N_5090);
nand U5606 (N_5606,N_4759,N_4724);
nand U5607 (N_5607,N_4994,N_4723);
nand U5608 (N_5608,N_4756,N_5097);
nand U5609 (N_5609,N_4591,N_4639);
and U5610 (N_5610,N_4647,N_4954);
xnor U5611 (N_5611,N_5226,N_5164);
and U5612 (N_5612,N_5005,N_4898);
nand U5613 (N_5613,N_5222,N_4526);
or U5614 (N_5614,N_4940,N_5179);
and U5615 (N_5615,N_4814,N_4515);
nor U5616 (N_5616,N_4674,N_5062);
and U5617 (N_5617,N_5102,N_4895);
nand U5618 (N_5618,N_4781,N_4601);
xor U5619 (N_5619,N_4511,N_5204);
or U5620 (N_5620,N_5175,N_5221);
nor U5621 (N_5621,N_5057,N_4516);
nor U5622 (N_5622,N_4931,N_5108);
nand U5623 (N_5623,N_4508,N_5113);
and U5624 (N_5624,N_4819,N_5014);
and U5625 (N_5625,N_4556,N_4833);
nor U5626 (N_5626,N_5080,N_4779);
nor U5627 (N_5627,N_4780,N_4950);
and U5628 (N_5628,N_4836,N_4900);
nand U5629 (N_5629,N_4555,N_4767);
xnor U5630 (N_5630,N_4796,N_4541);
xnor U5631 (N_5631,N_5002,N_4821);
and U5632 (N_5632,N_4878,N_4503);
nand U5633 (N_5633,N_4776,N_4679);
and U5634 (N_5634,N_5133,N_4680);
xor U5635 (N_5635,N_5190,N_5037);
or U5636 (N_5636,N_4917,N_4641);
nand U5637 (N_5637,N_4924,N_4867);
nor U5638 (N_5638,N_4796,N_5087);
or U5639 (N_5639,N_4564,N_5218);
nand U5640 (N_5640,N_4790,N_5167);
or U5641 (N_5641,N_4746,N_4920);
and U5642 (N_5642,N_4673,N_4968);
and U5643 (N_5643,N_5168,N_4765);
and U5644 (N_5644,N_4907,N_5078);
and U5645 (N_5645,N_4970,N_4594);
and U5646 (N_5646,N_4613,N_4756);
nand U5647 (N_5647,N_5061,N_5057);
and U5648 (N_5648,N_4811,N_5205);
and U5649 (N_5649,N_4948,N_4917);
and U5650 (N_5650,N_4667,N_4936);
nor U5651 (N_5651,N_4780,N_4999);
xor U5652 (N_5652,N_4810,N_4627);
and U5653 (N_5653,N_4732,N_4923);
and U5654 (N_5654,N_5014,N_4898);
nand U5655 (N_5655,N_4913,N_4655);
nor U5656 (N_5656,N_4697,N_5166);
and U5657 (N_5657,N_5215,N_4899);
or U5658 (N_5658,N_4860,N_4534);
nor U5659 (N_5659,N_4503,N_4749);
or U5660 (N_5660,N_4702,N_4843);
nand U5661 (N_5661,N_4900,N_4857);
nor U5662 (N_5662,N_4831,N_5095);
and U5663 (N_5663,N_5243,N_4592);
nand U5664 (N_5664,N_4648,N_4944);
nor U5665 (N_5665,N_4550,N_5120);
xor U5666 (N_5666,N_4973,N_4672);
xor U5667 (N_5667,N_5113,N_5198);
or U5668 (N_5668,N_4896,N_5249);
nand U5669 (N_5669,N_4535,N_4540);
and U5670 (N_5670,N_4616,N_4857);
or U5671 (N_5671,N_5064,N_5201);
or U5672 (N_5672,N_4645,N_4898);
and U5673 (N_5673,N_4541,N_4758);
nor U5674 (N_5674,N_4804,N_4678);
nor U5675 (N_5675,N_4603,N_4908);
nor U5676 (N_5676,N_4613,N_5073);
and U5677 (N_5677,N_4723,N_4609);
and U5678 (N_5678,N_4543,N_5152);
nor U5679 (N_5679,N_4824,N_4615);
or U5680 (N_5680,N_4801,N_4571);
nor U5681 (N_5681,N_5239,N_4834);
or U5682 (N_5682,N_5134,N_4774);
xnor U5683 (N_5683,N_4994,N_5125);
or U5684 (N_5684,N_4503,N_4734);
nand U5685 (N_5685,N_4965,N_4690);
and U5686 (N_5686,N_4574,N_4704);
nand U5687 (N_5687,N_5050,N_4901);
nor U5688 (N_5688,N_4923,N_5122);
nand U5689 (N_5689,N_5230,N_5175);
and U5690 (N_5690,N_4780,N_5155);
nor U5691 (N_5691,N_4711,N_4732);
and U5692 (N_5692,N_5044,N_4908);
and U5693 (N_5693,N_4915,N_5039);
nand U5694 (N_5694,N_4575,N_4663);
or U5695 (N_5695,N_5175,N_5157);
nor U5696 (N_5696,N_5184,N_4625);
nor U5697 (N_5697,N_4834,N_5031);
nor U5698 (N_5698,N_4913,N_4830);
nor U5699 (N_5699,N_4729,N_5062);
and U5700 (N_5700,N_5180,N_4852);
nand U5701 (N_5701,N_5214,N_5124);
nor U5702 (N_5702,N_4834,N_4897);
nand U5703 (N_5703,N_4706,N_5130);
and U5704 (N_5704,N_4885,N_5241);
nand U5705 (N_5705,N_5017,N_4991);
and U5706 (N_5706,N_5126,N_4785);
nor U5707 (N_5707,N_4975,N_4862);
nor U5708 (N_5708,N_4733,N_4709);
nand U5709 (N_5709,N_5133,N_4861);
and U5710 (N_5710,N_5071,N_5131);
nand U5711 (N_5711,N_5039,N_4842);
or U5712 (N_5712,N_4660,N_4650);
nor U5713 (N_5713,N_4644,N_5238);
and U5714 (N_5714,N_4665,N_4752);
nor U5715 (N_5715,N_4923,N_4965);
xnor U5716 (N_5716,N_4731,N_5141);
nand U5717 (N_5717,N_4614,N_4584);
nor U5718 (N_5718,N_5162,N_4726);
xor U5719 (N_5719,N_4666,N_4748);
nor U5720 (N_5720,N_4657,N_5086);
and U5721 (N_5721,N_5164,N_5002);
nor U5722 (N_5722,N_4765,N_4602);
nand U5723 (N_5723,N_5134,N_4766);
xnor U5724 (N_5724,N_4805,N_5117);
or U5725 (N_5725,N_4742,N_4608);
or U5726 (N_5726,N_4874,N_5024);
nor U5727 (N_5727,N_4656,N_5214);
and U5728 (N_5728,N_4719,N_5063);
or U5729 (N_5729,N_5116,N_5098);
and U5730 (N_5730,N_4890,N_4835);
and U5731 (N_5731,N_4594,N_4534);
and U5732 (N_5732,N_5078,N_5054);
or U5733 (N_5733,N_5032,N_5239);
xor U5734 (N_5734,N_4665,N_4630);
or U5735 (N_5735,N_4693,N_4957);
or U5736 (N_5736,N_4526,N_5184);
or U5737 (N_5737,N_4887,N_5059);
nor U5738 (N_5738,N_4585,N_4760);
nand U5739 (N_5739,N_4986,N_5078);
and U5740 (N_5740,N_5194,N_4744);
or U5741 (N_5741,N_4520,N_4628);
and U5742 (N_5742,N_4732,N_4603);
nand U5743 (N_5743,N_4617,N_4991);
nand U5744 (N_5744,N_5012,N_5101);
nor U5745 (N_5745,N_4644,N_4557);
or U5746 (N_5746,N_5124,N_4734);
and U5747 (N_5747,N_4658,N_4560);
and U5748 (N_5748,N_4549,N_4535);
and U5749 (N_5749,N_4923,N_4645);
nand U5750 (N_5750,N_4941,N_5053);
nand U5751 (N_5751,N_4539,N_4913);
or U5752 (N_5752,N_4743,N_4868);
nor U5753 (N_5753,N_4892,N_4506);
nand U5754 (N_5754,N_4606,N_4680);
and U5755 (N_5755,N_5058,N_5203);
nand U5756 (N_5756,N_4534,N_5151);
nand U5757 (N_5757,N_4881,N_5154);
nor U5758 (N_5758,N_5177,N_4820);
nand U5759 (N_5759,N_4959,N_5222);
and U5760 (N_5760,N_4750,N_5179);
nor U5761 (N_5761,N_4894,N_4652);
or U5762 (N_5762,N_4625,N_4751);
nand U5763 (N_5763,N_4521,N_4856);
nor U5764 (N_5764,N_4678,N_4859);
nor U5765 (N_5765,N_5180,N_4950);
or U5766 (N_5766,N_4880,N_5160);
nor U5767 (N_5767,N_4737,N_4606);
or U5768 (N_5768,N_4971,N_5015);
nand U5769 (N_5769,N_4633,N_4987);
and U5770 (N_5770,N_4740,N_5162);
nand U5771 (N_5771,N_4729,N_4643);
or U5772 (N_5772,N_4599,N_4653);
or U5773 (N_5773,N_4721,N_4792);
and U5774 (N_5774,N_5185,N_4897);
and U5775 (N_5775,N_4748,N_5137);
or U5776 (N_5776,N_5074,N_4671);
and U5777 (N_5777,N_4525,N_5171);
and U5778 (N_5778,N_4570,N_4553);
nand U5779 (N_5779,N_4528,N_4562);
xnor U5780 (N_5780,N_5148,N_4842);
xnor U5781 (N_5781,N_4808,N_5126);
nor U5782 (N_5782,N_5174,N_4517);
nor U5783 (N_5783,N_5156,N_5017);
xnor U5784 (N_5784,N_4891,N_5181);
nor U5785 (N_5785,N_4865,N_5153);
and U5786 (N_5786,N_4897,N_4673);
nand U5787 (N_5787,N_4533,N_5067);
nor U5788 (N_5788,N_4703,N_4730);
or U5789 (N_5789,N_5198,N_4919);
nor U5790 (N_5790,N_4672,N_4543);
or U5791 (N_5791,N_5011,N_4716);
or U5792 (N_5792,N_5148,N_4975);
nor U5793 (N_5793,N_4678,N_4980);
and U5794 (N_5794,N_4541,N_5013);
and U5795 (N_5795,N_4503,N_5176);
nand U5796 (N_5796,N_4671,N_4637);
nand U5797 (N_5797,N_4858,N_4552);
nand U5798 (N_5798,N_4819,N_4750);
and U5799 (N_5799,N_5074,N_4693);
or U5800 (N_5800,N_4904,N_4844);
xnor U5801 (N_5801,N_5159,N_5199);
nand U5802 (N_5802,N_4997,N_5198);
xor U5803 (N_5803,N_5048,N_4708);
nand U5804 (N_5804,N_4729,N_4754);
nand U5805 (N_5805,N_5207,N_4773);
nand U5806 (N_5806,N_5186,N_4623);
xor U5807 (N_5807,N_4783,N_4937);
or U5808 (N_5808,N_5177,N_4680);
or U5809 (N_5809,N_4920,N_5147);
or U5810 (N_5810,N_4683,N_4574);
or U5811 (N_5811,N_4825,N_4933);
xnor U5812 (N_5812,N_5091,N_5151);
or U5813 (N_5813,N_4660,N_4665);
nor U5814 (N_5814,N_5193,N_4944);
or U5815 (N_5815,N_5056,N_5006);
and U5816 (N_5816,N_4585,N_5201);
nand U5817 (N_5817,N_5141,N_4947);
nor U5818 (N_5818,N_4850,N_5155);
and U5819 (N_5819,N_4556,N_5001);
nand U5820 (N_5820,N_4877,N_4720);
nand U5821 (N_5821,N_4900,N_5192);
xnor U5822 (N_5822,N_4984,N_4503);
nand U5823 (N_5823,N_4910,N_4741);
nand U5824 (N_5824,N_5221,N_5145);
or U5825 (N_5825,N_4961,N_5043);
nand U5826 (N_5826,N_4833,N_5242);
nand U5827 (N_5827,N_4540,N_4878);
or U5828 (N_5828,N_5149,N_4903);
and U5829 (N_5829,N_4589,N_5207);
nor U5830 (N_5830,N_4679,N_4728);
nand U5831 (N_5831,N_4580,N_5235);
or U5832 (N_5832,N_4766,N_4925);
and U5833 (N_5833,N_5076,N_4877);
or U5834 (N_5834,N_5101,N_5156);
nor U5835 (N_5835,N_5118,N_4546);
or U5836 (N_5836,N_5024,N_5168);
and U5837 (N_5837,N_5057,N_4820);
or U5838 (N_5838,N_5148,N_4819);
and U5839 (N_5839,N_4922,N_4509);
nand U5840 (N_5840,N_4769,N_5029);
or U5841 (N_5841,N_4848,N_4916);
nand U5842 (N_5842,N_4711,N_4588);
nor U5843 (N_5843,N_5121,N_4915);
and U5844 (N_5844,N_5159,N_5178);
nor U5845 (N_5845,N_4853,N_4506);
or U5846 (N_5846,N_5140,N_4600);
or U5847 (N_5847,N_4500,N_4565);
or U5848 (N_5848,N_5042,N_4709);
nand U5849 (N_5849,N_5068,N_4594);
nor U5850 (N_5850,N_4890,N_4892);
and U5851 (N_5851,N_4660,N_4507);
nor U5852 (N_5852,N_4641,N_4974);
xor U5853 (N_5853,N_4745,N_4780);
or U5854 (N_5854,N_4849,N_5098);
xnor U5855 (N_5855,N_4962,N_4539);
or U5856 (N_5856,N_5130,N_5074);
nand U5857 (N_5857,N_4532,N_4589);
nor U5858 (N_5858,N_4703,N_4754);
nor U5859 (N_5859,N_4720,N_4539);
nand U5860 (N_5860,N_4628,N_4923);
xnor U5861 (N_5861,N_4797,N_5124);
nor U5862 (N_5862,N_4630,N_4704);
nand U5863 (N_5863,N_5009,N_5181);
nor U5864 (N_5864,N_4985,N_4961);
or U5865 (N_5865,N_4744,N_4965);
nand U5866 (N_5866,N_4687,N_5089);
or U5867 (N_5867,N_4672,N_5227);
nor U5868 (N_5868,N_5166,N_4649);
or U5869 (N_5869,N_4998,N_4808);
nor U5870 (N_5870,N_4735,N_4861);
nand U5871 (N_5871,N_4657,N_4778);
xnor U5872 (N_5872,N_5005,N_4569);
nand U5873 (N_5873,N_4518,N_4683);
and U5874 (N_5874,N_4785,N_4642);
xnor U5875 (N_5875,N_5230,N_4682);
and U5876 (N_5876,N_4663,N_4689);
or U5877 (N_5877,N_4740,N_5199);
xor U5878 (N_5878,N_5207,N_5017);
or U5879 (N_5879,N_5217,N_4933);
or U5880 (N_5880,N_5017,N_4716);
xor U5881 (N_5881,N_4939,N_4688);
xnor U5882 (N_5882,N_5021,N_5102);
and U5883 (N_5883,N_5144,N_5177);
and U5884 (N_5884,N_4787,N_4731);
or U5885 (N_5885,N_5080,N_4614);
and U5886 (N_5886,N_5032,N_4811);
and U5887 (N_5887,N_5174,N_4813);
nor U5888 (N_5888,N_4506,N_5163);
or U5889 (N_5889,N_4936,N_5087);
xor U5890 (N_5890,N_4972,N_4876);
xnor U5891 (N_5891,N_4882,N_4539);
and U5892 (N_5892,N_4723,N_5038);
or U5893 (N_5893,N_5235,N_4784);
and U5894 (N_5894,N_5122,N_4791);
and U5895 (N_5895,N_4552,N_4599);
xnor U5896 (N_5896,N_4612,N_5037);
nand U5897 (N_5897,N_4627,N_4681);
nand U5898 (N_5898,N_4672,N_4982);
or U5899 (N_5899,N_4713,N_4869);
xnor U5900 (N_5900,N_4669,N_4502);
nand U5901 (N_5901,N_5151,N_4695);
and U5902 (N_5902,N_4857,N_4942);
nor U5903 (N_5903,N_5126,N_4724);
nor U5904 (N_5904,N_4523,N_5082);
nand U5905 (N_5905,N_4757,N_5098);
xnor U5906 (N_5906,N_4871,N_5084);
and U5907 (N_5907,N_5067,N_4891);
and U5908 (N_5908,N_5203,N_4507);
nand U5909 (N_5909,N_4883,N_5119);
nand U5910 (N_5910,N_4700,N_4552);
nand U5911 (N_5911,N_4829,N_4766);
nor U5912 (N_5912,N_4738,N_4886);
and U5913 (N_5913,N_4915,N_4545);
nor U5914 (N_5914,N_4654,N_4942);
or U5915 (N_5915,N_5073,N_4905);
and U5916 (N_5916,N_4846,N_4539);
and U5917 (N_5917,N_4600,N_5148);
or U5918 (N_5918,N_4872,N_5245);
nand U5919 (N_5919,N_4743,N_4803);
or U5920 (N_5920,N_5177,N_4865);
xor U5921 (N_5921,N_4563,N_4785);
and U5922 (N_5922,N_4693,N_5193);
nand U5923 (N_5923,N_4572,N_5163);
and U5924 (N_5924,N_4622,N_4674);
nand U5925 (N_5925,N_4511,N_4628);
or U5926 (N_5926,N_4534,N_5240);
nand U5927 (N_5927,N_5175,N_5064);
nor U5928 (N_5928,N_5200,N_4617);
and U5929 (N_5929,N_4585,N_5222);
nand U5930 (N_5930,N_4868,N_4961);
nor U5931 (N_5931,N_4705,N_5003);
and U5932 (N_5932,N_4511,N_4793);
or U5933 (N_5933,N_4984,N_5039);
and U5934 (N_5934,N_4561,N_4694);
or U5935 (N_5935,N_4836,N_5190);
nand U5936 (N_5936,N_5225,N_4788);
or U5937 (N_5937,N_4899,N_5055);
and U5938 (N_5938,N_5205,N_4536);
and U5939 (N_5939,N_5174,N_5063);
nor U5940 (N_5940,N_4542,N_4537);
and U5941 (N_5941,N_4530,N_5227);
and U5942 (N_5942,N_4527,N_4953);
and U5943 (N_5943,N_4581,N_5032);
or U5944 (N_5944,N_4766,N_5227);
and U5945 (N_5945,N_4851,N_4783);
and U5946 (N_5946,N_4778,N_4892);
nand U5947 (N_5947,N_4526,N_4731);
nor U5948 (N_5948,N_4525,N_4605);
nor U5949 (N_5949,N_4560,N_5051);
and U5950 (N_5950,N_5001,N_4665);
xnor U5951 (N_5951,N_4571,N_5014);
or U5952 (N_5952,N_4560,N_4975);
or U5953 (N_5953,N_4589,N_5124);
or U5954 (N_5954,N_5013,N_4893);
nor U5955 (N_5955,N_4572,N_4646);
nor U5956 (N_5956,N_4979,N_5042);
nand U5957 (N_5957,N_5117,N_4587);
nor U5958 (N_5958,N_4956,N_4877);
or U5959 (N_5959,N_4923,N_5035);
or U5960 (N_5960,N_4605,N_5072);
xnor U5961 (N_5961,N_4533,N_4587);
nand U5962 (N_5962,N_5227,N_4539);
or U5963 (N_5963,N_4980,N_5140);
and U5964 (N_5964,N_5187,N_4659);
nor U5965 (N_5965,N_4723,N_4762);
nand U5966 (N_5966,N_5065,N_4695);
or U5967 (N_5967,N_4742,N_4552);
or U5968 (N_5968,N_4709,N_5120);
or U5969 (N_5969,N_4798,N_4710);
nor U5970 (N_5970,N_4975,N_4654);
nor U5971 (N_5971,N_4653,N_5081);
nand U5972 (N_5972,N_5138,N_4741);
and U5973 (N_5973,N_4988,N_4619);
nand U5974 (N_5974,N_4993,N_5163);
nand U5975 (N_5975,N_5220,N_4773);
nand U5976 (N_5976,N_4956,N_4769);
xnor U5977 (N_5977,N_4856,N_4949);
and U5978 (N_5978,N_5013,N_4891);
and U5979 (N_5979,N_4808,N_4995);
or U5980 (N_5980,N_4738,N_5216);
or U5981 (N_5981,N_4891,N_5109);
nand U5982 (N_5982,N_4554,N_4600);
nor U5983 (N_5983,N_4698,N_5196);
nand U5984 (N_5984,N_4666,N_5190);
or U5985 (N_5985,N_4638,N_4884);
and U5986 (N_5986,N_4833,N_4707);
nand U5987 (N_5987,N_5178,N_4780);
nor U5988 (N_5988,N_4649,N_4571);
and U5989 (N_5989,N_4503,N_4710);
nor U5990 (N_5990,N_4822,N_4964);
and U5991 (N_5991,N_5215,N_4880);
or U5992 (N_5992,N_5059,N_4657);
or U5993 (N_5993,N_4796,N_4906);
and U5994 (N_5994,N_4675,N_4996);
and U5995 (N_5995,N_5105,N_4832);
and U5996 (N_5996,N_4571,N_5019);
or U5997 (N_5997,N_4701,N_4776);
and U5998 (N_5998,N_4660,N_4758);
nand U5999 (N_5999,N_4787,N_5146);
xnor U6000 (N_6000,N_5486,N_5761);
nand U6001 (N_6001,N_5534,N_5789);
or U6002 (N_6002,N_5353,N_5730);
and U6003 (N_6003,N_5866,N_5937);
nand U6004 (N_6004,N_5646,N_5721);
or U6005 (N_6005,N_5458,N_5258);
nand U6006 (N_6006,N_5599,N_5334);
nor U6007 (N_6007,N_5921,N_5787);
nand U6008 (N_6008,N_5452,N_5467);
nor U6009 (N_6009,N_5352,N_5267);
nor U6010 (N_6010,N_5919,N_5766);
nor U6011 (N_6011,N_5318,N_5728);
and U6012 (N_6012,N_5907,N_5294);
nor U6013 (N_6013,N_5679,N_5429);
or U6014 (N_6014,N_5674,N_5500);
and U6015 (N_6015,N_5417,N_5445);
and U6016 (N_6016,N_5894,N_5282);
xnor U6017 (N_6017,N_5581,N_5925);
nor U6018 (N_6018,N_5924,N_5859);
nor U6019 (N_6019,N_5261,N_5935);
or U6020 (N_6020,N_5427,N_5453);
or U6021 (N_6021,N_5946,N_5831);
or U6022 (N_6022,N_5975,N_5804);
nand U6023 (N_6023,N_5487,N_5468);
nor U6024 (N_6024,N_5607,N_5876);
nor U6025 (N_6025,N_5898,N_5874);
and U6026 (N_6026,N_5600,N_5603);
or U6027 (N_6027,N_5471,N_5477);
xnor U6028 (N_6028,N_5839,N_5271);
or U6029 (N_6029,N_5771,N_5783);
nor U6030 (N_6030,N_5895,N_5531);
or U6031 (N_6031,N_5314,N_5993);
nand U6032 (N_6032,N_5812,N_5462);
nor U6033 (N_6033,N_5684,N_5595);
and U6034 (N_6034,N_5776,N_5338);
and U6035 (N_6035,N_5373,N_5317);
nand U6036 (N_6036,N_5465,N_5760);
and U6037 (N_6037,N_5576,N_5846);
nand U6038 (N_6038,N_5962,N_5662);
nor U6039 (N_6039,N_5914,N_5586);
nor U6040 (N_6040,N_5535,N_5345);
or U6041 (N_6041,N_5902,N_5544);
or U6042 (N_6042,N_5548,N_5801);
nand U6043 (N_6043,N_5396,N_5820);
or U6044 (N_6044,N_5504,N_5428);
or U6045 (N_6045,N_5527,N_5611);
nand U6046 (N_6046,N_5532,N_5568);
and U6047 (N_6047,N_5381,N_5339);
nor U6048 (N_6048,N_5250,N_5718);
xor U6049 (N_6049,N_5525,N_5496);
or U6050 (N_6050,N_5884,N_5751);
xor U6051 (N_6051,N_5631,N_5970);
nor U6052 (N_6052,N_5972,N_5436);
nor U6053 (N_6053,N_5648,N_5606);
nor U6054 (N_6054,N_5779,N_5392);
nor U6055 (N_6055,N_5479,N_5263);
nor U6056 (N_6056,N_5285,N_5998);
nor U6057 (N_6057,N_5514,N_5916);
or U6058 (N_6058,N_5253,N_5802);
or U6059 (N_6059,N_5624,N_5773);
or U6060 (N_6060,N_5419,N_5957);
nor U6061 (N_6061,N_5517,N_5753);
nand U6062 (N_6062,N_5834,N_5908);
nand U6063 (N_6063,N_5357,N_5327);
or U6064 (N_6064,N_5747,N_5347);
or U6065 (N_6065,N_5402,N_5832);
nor U6066 (N_6066,N_5320,N_5841);
and U6067 (N_6067,N_5974,N_5560);
nand U6068 (N_6068,N_5731,N_5494);
xor U6069 (N_6069,N_5750,N_5341);
nor U6070 (N_6070,N_5406,N_5868);
nor U6071 (N_6071,N_5940,N_5954);
nor U6072 (N_6072,N_5980,N_5852);
nand U6073 (N_6073,N_5829,N_5337);
nand U6074 (N_6074,N_5723,N_5572);
nor U6075 (N_6075,N_5764,N_5426);
or U6076 (N_6076,N_5538,N_5948);
and U6077 (N_6077,N_5604,N_5865);
nand U6078 (N_6078,N_5724,N_5552);
nand U6079 (N_6079,N_5609,N_5277);
xor U6080 (N_6080,N_5922,N_5255);
or U6081 (N_6081,N_5322,N_5585);
nand U6082 (N_6082,N_5378,N_5663);
nor U6083 (N_6083,N_5817,N_5823);
and U6084 (N_6084,N_5815,N_5546);
nor U6085 (N_6085,N_5754,N_5509);
nand U6086 (N_6086,N_5635,N_5448);
nor U6087 (N_6087,N_5644,N_5665);
nand U6088 (N_6088,N_5343,N_5302);
and U6089 (N_6089,N_5700,N_5579);
or U6090 (N_6090,N_5470,N_5822);
nand U6091 (N_6091,N_5621,N_5890);
or U6092 (N_6092,N_5694,N_5290);
nor U6093 (N_6093,N_5626,N_5401);
xor U6094 (N_6094,N_5422,N_5391);
nand U6095 (N_6095,N_5573,N_5481);
or U6096 (N_6096,N_5720,N_5668);
or U6097 (N_6097,N_5291,N_5714);
or U6098 (N_6098,N_5519,N_5652);
and U6099 (N_6099,N_5657,N_5778);
nand U6100 (N_6100,N_5870,N_5336);
and U6101 (N_6101,N_5466,N_5254);
or U6102 (N_6102,N_5757,N_5597);
or U6103 (N_6103,N_5814,N_5643);
nand U6104 (N_6104,N_5691,N_5912);
nor U6105 (N_6105,N_5272,N_5686);
nand U6106 (N_6106,N_5386,N_5387);
nor U6107 (N_6107,N_5702,N_5713);
xor U6108 (N_6108,N_5423,N_5601);
nor U6109 (N_6109,N_5257,N_5885);
nor U6110 (N_6110,N_5528,N_5941);
or U6111 (N_6111,N_5797,N_5955);
or U6112 (N_6112,N_5497,N_5639);
nor U6113 (N_6113,N_5301,N_5664);
or U6114 (N_6114,N_5491,N_5268);
nand U6115 (N_6115,N_5412,N_5973);
xnor U6116 (N_6116,N_5855,N_5354);
nor U6117 (N_6117,N_5415,N_5903);
or U6118 (N_6118,N_5440,N_5803);
nor U6119 (N_6119,N_5867,N_5942);
and U6120 (N_6120,N_5276,N_5329);
nor U6121 (N_6121,N_5408,N_5666);
xor U6122 (N_6122,N_5963,N_5325);
or U6123 (N_6123,N_5516,N_5892);
and U6124 (N_6124,N_5443,N_5368);
nor U6125 (N_6125,N_5455,N_5878);
nand U6126 (N_6126,N_5640,N_5360);
xnor U6127 (N_6127,N_5520,N_5602);
and U6128 (N_6128,N_5997,N_5710);
or U6129 (N_6129,N_5274,N_5591);
and U6130 (N_6130,N_5522,N_5616);
nand U6131 (N_6131,N_5541,N_5348);
and U6132 (N_6132,N_5400,N_5542);
nand U6133 (N_6133,N_5340,N_5939);
nand U6134 (N_6134,N_5904,N_5506);
nand U6135 (N_6135,N_5906,N_5698);
nor U6136 (N_6136,N_5252,N_5382);
nand U6137 (N_6137,N_5762,N_5879);
nand U6138 (N_6138,N_5739,N_5550);
or U6139 (N_6139,N_5598,N_5844);
or U6140 (N_6140,N_5807,N_5315);
nor U6141 (N_6141,N_5658,N_5434);
nor U6142 (N_6142,N_5655,N_5513);
nand U6143 (N_6143,N_5781,N_5279);
nor U6144 (N_6144,N_5346,N_5727);
or U6145 (N_6145,N_5351,N_5332);
nand U6146 (N_6146,N_5889,N_5659);
and U6147 (N_6147,N_5960,N_5265);
nor U6148 (N_6148,N_5266,N_5909);
nand U6149 (N_6149,N_5798,N_5888);
nand U6150 (N_6150,N_5370,N_5510);
nor U6151 (N_6151,N_5307,N_5413);
nor U6152 (N_6152,N_5649,N_5424);
and U6153 (N_6153,N_5397,N_5363);
xor U6154 (N_6154,N_5918,N_5669);
and U6155 (N_6155,N_5847,N_5838);
or U6156 (N_6156,N_5953,N_5565);
and U6157 (N_6157,N_5312,N_5310);
nand U6158 (N_6158,N_5505,N_5432);
and U6159 (N_6159,N_5837,N_5881);
nor U6160 (N_6160,N_5769,N_5951);
nor U6161 (N_6161,N_5873,N_5715);
nor U6162 (N_6162,N_5850,N_5701);
nand U6163 (N_6163,N_5326,N_5996);
nor U6164 (N_6164,N_5969,N_5619);
nor U6165 (N_6165,N_5571,N_5660);
nor U6166 (N_6166,N_5641,N_5447);
and U6167 (N_6167,N_5650,N_5705);
nand U6168 (N_6168,N_5435,N_5680);
or U6169 (N_6169,N_5654,N_5316);
nor U6170 (N_6170,N_5883,N_5930);
nor U6171 (N_6171,N_5545,N_5877);
and U6172 (N_6172,N_5275,N_5813);
nor U6173 (N_6173,N_5414,N_5835);
and U6174 (N_6174,N_5683,N_5688);
nor U6175 (N_6175,N_5732,N_5594);
nand U6176 (N_6176,N_5480,N_5526);
and U6177 (N_6177,N_5492,N_5667);
and U6178 (N_6178,N_5697,N_5596);
and U6179 (N_6179,N_5920,N_5809);
and U6180 (N_6180,N_5712,N_5805);
nand U6181 (N_6181,N_5670,N_5896);
nor U6182 (N_6182,N_5956,N_5981);
nor U6183 (N_6183,N_5746,N_5582);
nor U6184 (N_6184,N_5709,N_5741);
and U6185 (N_6185,N_5304,N_5843);
xor U6186 (N_6186,N_5968,N_5826);
xor U6187 (N_6187,N_5882,N_5676);
nand U6188 (N_6188,N_5661,N_5799);
nor U6189 (N_6189,N_5994,N_5482);
xnor U6190 (N_6190,N_5476,N_5938);
nor U6191 (N_6191,N_5886,N_5281);
or U6192 (N_6192,N_5488,N_5344);
nor U6193 (N_6193,N_5431,N_5411);
and U6194 (N_6194,N_5811,N_5444);
nor U6195 (N_6195,N_5449,N_5927);
nor U6196 (N_6196,N_5853,N_5848);
nand U6197 (N_6197,N_5305,N_5861);
nand U6198 (N_6198,N_5965,N_5979);
nand U6199 (N_6199,N_5533,N_5507);
xor U6200 (N_6200,N_5551,N_5840);
nor U6201 (N_6201,N_5398,N_5944);
or U6202 (N_6202,N_5299,N_5264);
nand U6203 (N_6203,N_5377,N_5463);
nand U6204 (N_6204,N_5614,N_5645);
xor U6205 (N_6205,N_5875,N_5342);
nor U6206 (N_6206,N_5899,N_5308);
or U6207 (N_6207,N_5438,N_5540);
nand U6208 (N_6208,N_5399,N_5736);
xnor U6209 (N_6209,N_5690,N_5503);
and U6210 (N_6210,N_5394,N_5259);
and U6211 (N_6211,N_5995,N_5409);
nor U6212 (N_6212,N_5765,N_5355);
or U6213 (N_6213,N_5695,N_5978);
nand U6214 (N_6214,N_5630,N_5923);
or U6215 (N_6215,N_5625,N_5950);
xor U6216 (N_6216,N_5795,N_5543);
nand U6217 (N_6217,N_5749,N_5744);
or U6218 (N_6218,N_5784,N_5763);
nor U6219 (N_6219,N_5917,N_5901);
or U6220 (N_6220,N_5410,N_5557);
and U6221 (N_6221,N_5605,N_5891);
or U6222 (N_6222,N_5359,N_5735);
xor U6223 (N_6223,N_5703,N_5869);
and U6224 (N_6224,N_5459,N_5748);
nor U6225 (N_6225,N_5380,N_5403);
and U6226 (N_6226,N_5623,N_5521);
nor U6227 (N_6227,N_5716,N_5910);
nor U6228 (N_6228,N_5931,N_5537);
and U6229 (N_6229,N_5425,N_5966);
nor U6230 (N_6230,N_5677,N_5722);
nand U6231 (N_6231,N_5785,N_5977);
nor U6232 (N_6232,N_5364,N_5828);
nor U6233 (N_6233,N_5692,N_5260);
or U6234 (N_6234,N_5295,N_5362);
or U6235 (N_6235,N_5366,N_5756);
or U6236 (N_6236,N_5964,N_5593);
or U6237 (N_6237,N_5464,N_5587);
and U6238 (N_6238,N_5439,N_5369);
xor U6239 (N_6239,N_5758,N_5733);
and U6240 (N_6240,N_5478,N_5564);
or U6241 (N_6241,N_5495,N_5856);
nand U6242 (N_6242,N_5303,N_5437);
or U6243 (N_6243,N_5256,N_5986);
nand U6244 (N_6244,N_5622,N_5984);
nor U6245 (N_6245,N_5682,N_5270);
nor U6246 (N_6246,N_5372,N_5793);
or U6247 (N_6247,N_5553,N_5286);
xnor U6248 (N_6248,N_5592,N_5926);
or U6249 (N_6249,N_5508,N_5777);
and U6250 (N_6250,N_5711,N_5755);
nand U6251 (N_6251,N_5985,N_5418);
nand U6252 (N_6252,N_5588,N_5775);
nor U6253 (N_6253,N_5851,N_5880);
nor U6254 (N_6254,N_5794,N_5992);
or U6255 (N_6255,N_5289,N_5499);
nand U6256 (N_6256,N_5780,N_5485);
and U6257 (N_6257,N_5900,N_5292);
xnor U6258 (N_6258,N_5943,N_5772);
and U6259 (N_6259,N_5752,N_5420);
nor U6260 (N_6260,N_5913,N_5864);
nand U6261 (N_6261,N_5999,N_5759);
and U6262 (N_6262,N_5707,N_5945);
nand U6263 (N_6263,N_5678,N_5278);
nand U6264 (N_6264,N_5330,N_5297);
xor U6265 (N_6265,N_5791,N_5383);
or U6266 (N_6266,N_5473,N_5932);
and U6267 (N_6267,N_5335,N_5390);
nor U6268 (N_6268,N_5570,N_5321);
and U6269 (N_6269,N_5450,N_5991);
or U6270 (N_6270,N_5313,N_5566);
nand U6271 (N_6271,N_5726,N_5384);
or U6272 (N_6272,N_5699,N_5498);
nand U6273 (N_6273,N_5349,N_5421);
nor U6274 (N_6274,N_5638,N_5567);
or U6275 (N_6275,N_5293,N_5961);
or U6276 (N_6276,N_5827,N_5687);
and U6277 (N_6277,N_5734,N_5836);
or U6278 (N_6278,N_5284,N_5800);
or U6279 (N_6279,N_5407,N_5502);
nor U6280 (N_6280,N_5633,N_5441);
nand U6281 (N_6281,N_5433,N_5512);
or U6282 (N_6282,N_5983,N_5673);
and U6283 (N_6283,N_5489,N_5331);
nand U6284 (N_6284,N_5627,N_5262);
or U6285 (N_6285,N_5483,N_5928);
nand U6286 (N_6286,N_5636,N_5356);
nor U6287 (N_6287,N_5792,N_5361);
nand U6288 (N_6288,N_5589,N_5474);
nor U6289 (N_6289,N_5460,N_5833);
nor U6290 (N_6290,N_5934,N_5719);
or U6291 (N_6291,N_5949,N_5740);
and U6292 (N_6292,N_5298,N_5849);
or U6293 (N_6293,N_5563,N_5615);
nand U6294 (N_6294,N_5933,N_5457);
nand U6295 (N_6295,N_5283,N_5613);
and U6296 (N_6296,N_5612,N_5887);
or U6297 (N_6297,N_5515,N_5620);
nor U6298 (N_6298,N_5367,N_5562);
nor U6299 (N_6299,N_5893,N_5583);
and U6300 (N_6300,N_5717,N_5743);
or U6301 (N_6301,N_5461,N_5511);
or U6302 (N_6302,N_5704,N_5309);
nor U6303 (N_6303,N_5796,N_5379);
and U6304 (N_6304,N_5810,N_5374);
or U6305 (N_6305,N_5529,N_5617);
xor U6306 (N_6306,N_5501,N_5737);
xor U6307 (N_6307,N_5610,N_5629);
nor U6308 (N_6308,N_5818,N_5971);
or U6309 (N_6309,N_5689,N_5393);
and U6310 (N_6310,N_5915,N_5311);
and U6311 (N_6311,N_5416,N_5905);
or U6312 (N_6312,N_5745,N_5385);
or U6313 (N_6313,N_5988,N_5989);
nor U6314 (N_6314,N_5388,N_5559);
nor U6315 (N_6315,N_5446,N_5539);
nor U6316 (N_6316,N_5816,N_5288);
or U6317 (N_6317,N_5574,N_5269);
nand U6318 (N_6318,N_5872,N_5681);
nor U6319 (N_6319,N_5857,N_5782);
nand U6320 (N_6320,N_5389,N_5929);
and U6321 (N_6321,N_5632,N_5990);
or U6322 (N_6322,N_5371,N_5536);
nor U6323 (N_6323,N_5959,N_5858);
or U6324 (N_6324,N_5790,N_5584);
nand U6325 (N_6325,N_5628,N_5577);
xnor U6326 (N_6326,N_5350,N_5405);
nand U6327 (N_6327,N_5863,N_5845);
and U6328 (N_6328,N_5358,N_5967);
or U6329 (N_6329,N_5558,N_5788);
nor U6330 (N_6330,N_5642,N_5651);
nand U6331 (N_6331,N_5280,N_5842);
or U6332 (N_6332,N_5524,N_5273);
and U6333 (N_6333,N_5442,N_5569);
xnor U6334 (N_6334,N_5333,N_5556);
or U6335 (N_6335,N_5580,N_5819);
nand U6336 (N_6336,N_5806,N_5365);
or U6337 (N_6337,N_5729,N_5675);
nand U6338 (N_6338,N_5738,N_5708);
nor U6339 (N_6339,N_5518,N_5947);
or U6340 (N_6340,N_5490,N_5547);
xor U6341 (N_6341,N_5300,N_5475);
or U6342 (N_6342,N_5830,N_5530);
nand U6343 (N_6343,N_5561,N_5575);
and U6344 (N_6344,N_5871,N_5653);
nor U6345 (N_6345,N_5323,N_5376);
nand U6346 (N_6346,N_5608,N_5618);
and U6347 (N_6347,N_5767,N_5824);
nand U6348 (N_6348,N_5911,N_5555);
or U6349 (N_6349,N_5976,N_5854);
nor U6350 (N_6350,N_5554,N_5770);
nand U6351 (N_6351,N_5696,N_5306);
xor U6352 (N_6352,N_5952,N_5375);
nand U6353 (N_6353,N_5590,N_5469);
xor U6354 (N_6354,N_5958,N_5742);
nor U6355 (N_6355,N_5634,N_5725);
and U6356 (N_6356,N_5768,N_5484);
or U6357 (N_6357,N_5523,N_5549);
nor U6358 (N_6358,N_5637,N_5251);
xnor U6359 (N_6359,N_5685,N_5860);
nand U6360 (N_6360,N_5936,N_5982);
and U6361 (N_6361,N_5472,N_5821);
xor U6362 (N_6362,N_5647,N_5319);
nor U6363 (N_6363,N_5454,N_5578);
nor U6364 (N_6364,N_5862,N_5296);
nor U6365 (N_6365,N_5774,N_5404);
xor U6366 (N_6366,N_5825,N_5493);
nor U6367 (N_6367,N_5672,N_5430);
nand U6368 (N_6368,N_5328,N_5706);
nand U6369 (N_6369,N_5451,N_5287);
xor U6370 (N_6370,N_5987,N_5897);
or U6371 (N_6371,N_5671,N_5324);
nor U6372 (N_6372,N_5808,N_5693);
nand U6373 (N_6373,N_5456,N_5395);
or U6374 (N_6374,N_5786,N_5656);
nand U6375 (N_6375,N_5290,N_5991);
nor U6376 (N_6376,N_5282,N_5632);
or U6377 (N_6377,N_5706,N_5463);
and U6378 (N_6378,N_5438,N_5258);
or U6379 (N_6379,N_5827,N_5977);
or U6380 (N_6380,N_5999,N_5400);
nand U6381 (N_6381,N_5773,N_5665);
xnor U6382 (N_6382,N_5520,N_5609);
nor U6383 (N_6383,N_5993,N_5945);
nor U6384 (N_6384,N_5546,N_5330);
and U6385 (N_6385,N_5295,N_5866);
nand U6386 (N_6386,N_5253,N_5874);
or U6387 (N_6387,N_5882,N_5926);
and U6388 (N_6388,N_5571,N_5383);
or U6389 (N_6389,N_5347,N_5349);
or U6390 (N_6390,N_5731,N_5991);
nor U6391 (N_6391,N_5873,N_5448);
or U6392 (N_6392,N_5963,N_5896);
or U6393 (N_6393,N_5671,N_5510);
and U6394 (N_6394,N_5980,N_5324);
or U6395 (N_6395,N_5486,N_5712);
and U6396 (N_6396,N_5774,N_5548);
or U6397 (N_6397,N_5423,N_5795);
or U6398 (N_6398,N_5724,N_5565);
nor U6399 (N_6399,N_5597,N_5798);
xor U6400 (N_6400,N_5785,N_5852);
or U6401 (N_6401,N_5844,N_5855);
nor U6402 (N_6402,N_5579,N_5273);
nand U6403 (N_6403,N_5621,N_5613);
xnor U6404 (N_6404,N_5349,N_5875);
xnor U6405 (N_6405,N_5782,N_5565);
nor U6406 (N_6406,N_5973,N_5770);
nor U6407 (N_6407,N_5957,N_5625);
and U6408 (N_6408,N_5886,N_5440);
and U6409 (N_6409,N_5308,N_5289);
and U6410 (N_6410,N_5570,N_5390);
xor U6411 (N_6411,N_5958,N_5624);
nand U6412 (N_6412,N_5608,N_5260);
or U6413 (N_6413,N_5880,N_5817);
and U6414 (N_6414,N_5978,N_5693);
nor U6415 (N_6415,N_5367,N_5587);
or U6416 (N_6416,N_5960,N_5464);
and U6417 (N_6417,N_5349,N_5780);
or U6418 (N_6418,N_5923,N_5509);
nand U6419 (N_6419,N_5894,N_5815);
nand U6420 (N_6420,N_5336,N_5666);
nor U6421 (N_6421,N_5485,N_5325);
nand U6422 (N_6422,N_5277,N_5917);
xnor U6423 (N_6423,N_5537,N_5361);
and U6424 (N_6424,N_5275,N_5465);
or U6425 (N_6425,N_5553,N_5669);
nand U6426 (N_6426,N_5859,N_5412);
or U6427 (N_6427,N_5705,N_5371);
and U6428 (N_6428,N_5655,N_5784);
nor U6429 (N_6429,N_5471,N_5707);
nand U6430 (N_6430,N_5798,N_5606);
and U6431 (N_6431,N_5726,N_5445);
or U6432 (N_6432,N_5257,N_5357);
or U6433 (N_6433,N_5443,N_5542);
nand U6434 (N_6434,N_5978,N_5911);
nor U6435 (N_6435,N_5508,N_5801);
nor U6436 (N_6436,N_5266,N_5259);
nand U6437 (N_6437,N_5707,N_5450);
and U6438 (N_6438,N_5750,N_5625);
nand U6439 (N_6439,N_5262,N_5727);
nand U6440 (N_6440,N_5460,N_5861);
nand U6441 (N_6441,N_5403,N_5508);
and U6442 (N_6442,N_5994,N_5945);
and U6443 (N_6443,N_5949,N_5602);
and U6444 (N_6444,N_5719,N_5843);
nor U6445 (N_6445,N_5870,N_5827);
and U6446 (N_6446,N_5928,N_5332);
nor U6447 (N_6447,N_5335,N_5323);
nor U6448 (N_6448,N_5882,N_5649);
or U6449 (N_6449,N_5335,N_5704);
and U6450 (N_6450,N_5644,N_5969);
nor U6451 (N_6451,N_5658,N_5764);
nor U6452 (N_6452,N_5324,N_5605);
and U6453 (N_6453,N_5630,N_5548);
or U6454 (N_6454,N_5377,N_5742);
nor U6455 (N_6455,N_5444,N_5601);
and U6456 (N_6456,N_5341,N_5773);
and U6457 (N_6457,N_5624,N_5631);
or U6458 (N_6458,N_5834,N_5338);
and U6459 (N_6459,N_5319,N_5263);
or U6460 (N_6460,N_5482,N_5724);
and U6461 (N_6461,N_5377,N_5454);
or U6462 (N_6462,N_5484,N_5583);
nand U6463 (N_6463,N_5921,N_5905);
nor U6464 (N_6464,N_5892,N_5660);
nand U6465 (N_6465,N_5847,N_5968);
nand U6466 (N_6466,N_5946,N_5596);
or U6467 (N_6467,N_5712,N_5758);
nor U6468 (N_6468,N_5775,N_5286);
nor U6469 (N_6469,N_5269,N_5338);
and U6470 (N_6470,N_5701,N_5746);
or U6471 (N_6471,N_5430,N_5900);
nor U6472 (N_6472,N_5336,N_5834);
or U6473 (N_6473,N_5561,N_5447);
and U6474 (N_6474,N_5886,N_5640);
or U6475 (N_6475,N_5663,N_5656);
xnor U6476 (N_6476,N_5285,N_5732);
nand U6477 (N_6477,N_5932,N_5872);
or U6478 (N_6478,N_5971,N_5705);
nor U6479 (N_6479,N_5352,N_5274);
nand U6480 (N_6480,N_5359,N_5731);
or U6481 (N_6481,N_5297,N_5761);
or U6482 (N_6482,N_5761,N_5350);
nand U6483 (N_6483,N_5445,N_5537);
or U6484 (N_6484,N_5383,N_5657);
xor U6485 (N_6485,N_5633,N_5314);
and U6486 (N_6486,N_5482,N_5886);
nand U6487 (N_6487,N_5634,N_5463);
and U6488 (N_6488,N_5862,N_5981);
or U6489 (N_6489,N_5454,N_5401);
nand U6490 (N_6490,N_5367,N_5894);
and U6491 (N_6491,N_5472,N_5644);
or U6492 (N_6492,N_5527,N_5415);
nand U6493 (N_6493,N_5567,N_5679);
and U6494 (N_6494,N_5530,N_5714);
nand U6495 (N_6495,N_5945,N_5744);
and U6496 (N_6496,N_5984,N_5266);
nor U6497 (N_6497,N_5505,N_5857);
nor U6498 (N_6498,N_5497,N_5344);
and U6499 (N_6499,N_5290,N_5752);
and U6500 (N_6500,N_5765,N_5531);
xor U6501 (N_6501,N_5315,N_5513);
nor U6502 (N_6502,N_5407,N_5903);
nand U6503 (N_6503,N_5770,N_5250);
and U6504 (N_6504,N_5270,N_5624);
xor U6505 (N_6505,N_5626,N_5890);
nor U6506 (N_6506,N_5745,N_5806);
nor U6507 (N_6507,N_5470,N_5900);
or U6508 (N_6508,N_5544,N_5746);
xor U6509 (N_6509,N_5911,N_5851);
nand U6510 (N_6510,N_5890,N_5372);
xor U6511 (N_6511,N_5841,N_5326);
nor U6512 (N_6512,N_5934,N_5384);
and U6513 (N_6513,N_5549,N_5771);
or U6514 (N_6514,N_5797,N_5908);
xnor U6515 (N_6515,N_5496,N_5758);
nand U6516 (N_6516,N_5547,N_5424);
nand U6517 (N_6517,N_5934,N_5555);
and U6518 (N_6518,N_5443,N_5982);
nand U6519 (N_6519,N_5328,N_5710);
nand U6520 (N_6520,N_5270,N_5414);
or U6521 (N_6521,N_5673,N_5700);
and U6522 (N_6522,N_5905,N_5876);
nand U6523 (N_6523,N_5478,N_5467);
or U6524 (N_6524,N_5879,N_5547);
and U6525 (N_6525,N_5864,N_5578);
and U6526 (N_6526,N_5566,N_5359);
nand U6527 (N_6527,N_5269,N_5905);
nand U6528 (N_6528,N_5730,N_5410);
or U6529 (N_6529,N_5621,N_5297);
and U6530 (N_6530,N_5726,N_5627);
and U6531 (N_6531,N_5254,N_5446);
nand U6532 (N_6532,N_5574,N_5930);
nand U6533 (N_6533,N_5853,N_5298);
and U6534 (N_6534,N_5347,N_5911);
or U6535 (N_6535,N_5732,N_5556);
nand U6536 (N_6536,N_5780,N_5779);
xor U6537 (N_6537,N_5731,N_5651);
and U6538 (N_6538,N_5377,N_5883);
nor U6539 (N_6539,N_5385,N_5723);
nor U6540 (N_6540,N_5973,N_5787);
and U6541 (N_6541,N_5862,N_5933);
xnor U6542 (N_6542,N_5633,N_5637);
and U6543 (N_6543,N_5960,N_5652);
and U6544 (N_6544,N_5859,N_5882);
nor U6545 (N_6545,N_5391,N_5319);
xnor U6546 (N_6546,N_5408,N_5869);
nor U6547 (N_6547,N_5611,N_5668);
nor U6548 (N_6548,N_5728,N_5912);
nor U6549 (N_6549,N_5836,N_5879);
xor U6550 (N_6550,N_5277,N_5663);
nor U6551 (N_6551,N_5397,N_5716);
nand U6552 (N_6552,N_5902,N_5738);
or U6553 (N_6553,N_5261,N_5450);
and U6554 (N_6554,N_5803,N_5961);
nor U6555 (N_6555,N_5695,N_5889);
nand U6556 (N_6556,N_5566,N_5959);
nand U6557 (N_6557,N_5730,N_5555);
nor U6558 (N_6558,N_5757,N_5275);
nand U6559 (N_6559,N_5947,N_5330);
xor U6560 (N_6560,N_5382,N_5706);
xor U6561 (N_6561,N_5470,N_5712);
and U6562 (N_6562,N_5554,N_5677);
or U6563 (N_6563,N_5577,N_5429);
nand U6564 (N_6564,N_5439,N_5366);
or U6565 (N_6565,N_5679,N_5419);
nand U6566 (N_6566,N_5469,N_5365);
nand U6567 (N_6567,N_5985,N_5822);
nor U6568 (N_6568,N_5689,N_5677);
or U6569 (N_6569,N_5271,N_5281);
xnor U6570 (N_6570,N_5750,N_5910);
xor U6571 (N_6571,N_5492,N_5915);
or U6572 (N_6572,N_5317,N_5642);
nor U6573 (N_6573,N_5900,N_5558);
and U6574 (N_6574,N_5683,N_5404);
and U6575 (N_6575,N_5932,N_5265);
or U6576 (N_6576,N_5806,N_5739);
nand U6577 (N_6577,N_5359,N_5282);
xnor U6578 (N_6578,N_5686,N_5921);
and U6579 (N_6579,N_5279,N_5523);
and U6580 (N_6580,N_5731,N_5379);
nor U6581 (N_6581,N_5250,N_5700);
and U6582 (N_6582,N_5859,N_5793);
and U6583 (N_6583,N_5595,N_5371);
nand U6584 (N_6584,N_5415,N_5901);
or U6585 (N_6585,N_5344,N_5555);
and U6586 (N_6586,N_5352,N_5288);
nand U6587 (N_6587,N_5414,N_5754);
nand U6588 (N_6588,N_5677,N_5545);
and U6589 (N_6589,N_5691,N_5791);
nor U6590 (N_6590,N_5568,N_5465);
or U6591 (N_6591,N_5301,N_5964);
nor U6592 (N_6592,N_5445,N_5882);
and U6593 (N_6593,N_5915,N_5626);
or U6594 (N_6594,N_5363,N_5889);
nand U6595 (N_6595,N_5313,N_5685);
and U6596 (N_6596,N_5576,N_5577);
or U6597 (N_6597,N_5918,N_5363);
and U6598 (N_6598,N_5919,N_5912);
nor U6599 (N_6599,N_5687,N_5411);
nor U6600 (N_6600,N_5314,N_5838);
or U6601 (N_6601,N_5490,N_5689);
or U6602 (N_6602,N_5550,N_5322);
nor U6603 (N_6603,N_5403,N_5543);
nand U6604 (N_6604,N_5863,N_5760);
or U6605 (N_6605,N_5638,N_5913);
and U6606 (N_6606,N_5431,N_5943);
nor U6607 (N_6607,N_5641,N_5620);
nand U6608 (N_6608,N_5295,N_5773);
and U6609 (N_6609,N_5895,N_5604);
and U6610 (N_6610,N_5324,N_5682);
nor U6611 (N_6611,N_5811,N_5371);
nand U6612 (N_6612,N_5433,N_5432);
or U6613 (N_6613,N_5482,N_5905);
nand U6614 (N_6614,N_5702,N_5827);
or U6615 (N_6615,N_5956,N_5442);
and U6616 (N_6616,N_5827,N_5286);
or U6617 (N_6617,N_5958,N_5263);
nand U6618 (N_6618,N_5448,N_5441);
or U6619 (N_6619,N_5311,N_5265);
and U6620 (N_6620,N_5293,N_5453);
nand U6621 (N_6621,N_5777,N_5902);
xnor U6622 (N_6622,N_5758,N_5854);
nor U6623 (N_6623,N_5685,N_5983);
or U6624 (N_6624,N_5571,N_5914);
nand U6625 (N_6625,N_5767,N_5682);
xor U6626 (N_6626,N_5306,N_5698);
nand U6627 (N_6627,N_5517,N_5400);
nor U6628 (N_6628,N_5565,N_5667);
and U6629 (N_6629,N_5356,N_5453);
and U6630 (N_6630,N_5892,N_5651);
and U6631 (N_6631,N_5276,N_5940);
and U6632 (N_6632,N_5785,N_5289);
xor U6633 (N_6633,N_5298,N_5372);
and U6634 (N_6634,N_5998,N_5972);
nand U6635 (N_6635,N_5387,N_5330);
and U6636 (N_6636,N_5817,N_5702);
xor U6637 (N_6637,N_5751,N_5367);
and U6638 (N_6638,N_5919,N_5635);
and U6639 (N_6639,N_5992,N_5815);
nand U6640 (N_6640,N_5388,N_5496);
nand U6641 (N_6641,N_5495,N_5358);
and U6642 (N_6642,N_5660,N_5788);
and U6643 (N_6643,N_5828,N_5888);
nor U6644 (N_6644,N_5892,N_5262);
nor U6645 (N_6645,N_5412,N_5906);
and U6646 (N_6646,N_5691,N_5469);
nor U6647 (N_6647,N_5953,N_5945);
nor U6648 (N_6648,N_5594,N_5562);
nor U6649 (N_6649,N_5301,N_5903);
or U6650 (N_6650,N_5333,N_5424);
nand U6651 (N_6651,N_5838,N_5584);
and U6652 (N_6652,N_5791,N_5862);
xnor U6653 (N_6653,N_5514,N_5975);
nor U6654 (N_6654,N_5713,N_5598);
and U6655 (N_6655,N_5470,N_5571);
or U6656 (N_6656,N_5532,N_5373);
nor U6657 (N_6657,N_5329,N_5620);
nand U6658 (N_6658,N_5873,N_5610);
nand U6659 (N_6659,N_5692,N_5661);
nand U6660 (N_6660,N_5623,N_5715);
nand U6661 (N_6661,N_5574,N_5743);
and U6662 (N_6662,N_5259,N_5354);
and U6663 (N_6663,N_5820,N_5876);
or U6664 (N_6664,N_5588,N_5273);
or U6665 (N_6665,N_5551,N_5652);
nand U6666 (N_6666,N_5644,N_5502);
xnor U6667 (N_6667,N_5623,N_5880);
and U6668 (N_6668,N_5971,N_5747);
nand U6669 (N_6669,N_5897,N_5786);
nor U6670 (N_6670,N_5374,N_5918);
xnor U6671 (N_6671,N_5529,N_5345);
or U6672 (N_6672,N_5580,N_5791);
nor U6673 (N_6673,N_5570,N_5687);
nor U6674 (N_6674,N_5939,N_5846);
and U6675 (N_6675,N_5491,N_5251);
nand U6676 (N_6676,N_5283,N_5708);
nand U6677 (N_6677,N_5892,N_5718);
and U6678 (N_6678,N_5452,N_5932);
nand U6679 (N_6679,N_5931,N_5377);
or U6680 (N_6680,N_5457,N_5311);
or U6681 (N_6681,N_5881,N_5411);
or U6682 (N_6682,N_5855,N_5439);
nand U6683 (N_6683,N_5768,N_5791);
nor U6684 (N_6684,N_5553,N_5605);
nand U6685 (N_6685,N_5328,N_5289);
or U6686 (N_6686,N_5552,N_5275);
and U6687 (N_6687,N_5736,N_5540);
nor U6688 (N_6688,N_5376,N_5469);
nor U6689 (N_6689,N_5339,N_5795);
or U6690 (N_6690,N_5974,N_5579);
nand U6691 (N_6691,N_5394,N_5485);
or U6692 (N_6692,N_5819,N_5408);
and U6693 (N_6693,N_5863,N_5280);
or U6694 (N_6694,N_5912,N_5555);
or U6695 (N_6695,N_5752,N_5487);
and U6696 (N_6696,N_5530,N_5688);
nand U6697 (N_6697,N_5900,N_5506);
or U6698 (N_6698,N_5638,N_5394);
nor U6699 (N_6699,N_5721,N_5296);
and U6700 (N_6700,N_5781,N_5738);
nor U6701 (N_6701,N_5551,N_5941);
and U6702 (N_6702,N_5409,N_5711);
nor U6703 (N_6703,N_5284,N_5946);
and U6704 (N_6704,N_5687,N_5305);
nor U6705 (N_6705,N_5994,N_5459);
and U6706 (N_6706,N_5939,N_5911);
nor U6707 (N_6707,N_5827,N_5329);
xor U6708 (N_6708,N_5627,N_5958);
nor U6709 (N_6709,N_5430,N_5966);
nand U6710 (N_6710,N_5802,N_5878);
xnor U6711 (N_6711,N_5612,N_5574);
nor U6712 (N_6712,N_5910,N_5631);
nand U6713 (N_6713,N_5714,N_5760);
xor U6714 (N_6714,N_5250,N_5561);
nor U6715 (N_6715,N_5820,N_5264);
and U6716 (N_6716,N_5958,N_5944);
and U6717 (N_6717,N_5455,N_5492);
xnor U6718 (N_6718,N_5909,N_5735);
and U6719 (N_6719,N_5779,N_5764);
and U6720 (N_6720,N_5778,N_5264);
nand U6721 (N_6721,N_5850,N_5847);
xor U6722 (N_6722,N_5850,N_5693);
and U6723 (N_6723,N_5872,N_5690);
nor U6724 (N_6724,N_5540,N_5548);
and U6725 (N_6725,N_5666,N_5766);
nor U6726 (N_6726,N_5810,N_5422);
and U6727 (N_6727,N_5648,N_5628);
nor U6728 (N_6728,N_5941,N_5796);
nand U6729 (N_6729,N_5631,N_5596);
or U6730 (N_6730,N_5250,N_5423);
nor U6731 (N_6731,N_5859,N_5609);
nand U6732 (N_6732,N_5296,N_5372);
and U6733 (N_6733,N_5581,N_5556);
nand U6734 (N_6734,N_5950,N_5864);
or U6735 (N_6735,N_5908,N_5845);
nor U6736 (N_6736,N_5357,N_5371);
xnor U6737 (N_6737,N_5357,N_5339);
and U6738 (N_6738,N_5499,N_5448);
and U6739 (N_6739,N_5933,N_5668);
or U6740 (N_6740,N_5559,N_5845);
or U6741 (N_6741,N_5535,N_5913);
and U6742 (N_6742,N_5869,N_5733);
or U6743 (N_6743,N_5825,N_5359);
or U6744 (N_6744,N_5947,N_5942);
or U6745 (N_6745,N_5672,N_5425);
and U6746 (N_6746,N_5305,N_5546);
nor U6747 (N_6747,N_5889,N_5313);
and U6748 (N_6748,N_5499,N_5808);
or U6749 (N_6749,N_5622,N_5764);
and U6750 (N_6750,N_6381,N_6382);
nand U6751 (N_6751,N_6130,N_6697);
or U6752 (N_6752,N_6417,N_6566);
nand U6753 (N_6753,N_6675,N_6407);
or U6754 (N_6754,N_6258,N_6559);
xor U6755 (N_6755,N_6578,N_6028);
or U6756 (N_6756,N_6183,N_6469);
or U6757 (N_6757,N_6474,N_6124);
nand U6758 (N_6758,N_6403,N_6097);
or U6759 (N_6759,N_6590,N_6058);
or U6760 (N_6760,N_6207,N_6351);
nor U6761 (N_6761,N_6193,N_6681);
nor U6762 (N_6762,N_6109,N_6427);
nor U6763 (N_6763,N_6485,N_6588);
or U6764 (N_6764,N_6747,N_6635);
nand U6765 (N_6765,N_6375,N_6245);
nand U6766 (N_6766,N_6569,N_6303);
nand U6767 (N_6767,N_6378,N_6227);
or U6768 (N_6768,N_6576,N_6323);
or U6769 (N_6769,N_6198,N_6437);
and U6770 (N_6770,N_6338,N_6110);
nand U6771 (N_6771,N_6367,N_6545);
or U6772 (N_6772,N_6528,N_6271);
and U6773 (N_6773,N_6254,N_6431);
or U6774 (N_6774,N_6636,N_6579);
and U6775 (N_6775,N_6076,N_6422);
nor U6776 (N_6776,N_6455,N_6025);
nor U6777 (N_6777,N_6293,N_6242);
xnor U6778 (N_6778,N_6464,N_6599);
or U6779 (N_6779,N_6461,N_6621);
nor U6780 (N_6780,N_6401,N_6359);
and U6781 (N_6781,N_6530,N_6283);
nand U6782 (N_6782,N_6399,N_6036);
nor U6783 (N_6783,N_6415,N_6612);
nor U6784 (N_6784,N_6581,N_6302);
or U6785 (N_6785,N_6192,N_6572);
or U6786 (N_6786,N_6190,N_6660);
or U6787 (N_6787,N_6249,N_6389);
or U6788 (N_6788,N_6372,N_6045);
or U6789 (N_6789,N_6223,N_6252);
or U6790 (N_6790,N_6208,N_6584);
and U6791 (N_6791,N_6487,N_6472);
and U6792 (N_6792,N_6720,N_6240);
nand U6793 (N_6793,N_6695,N_6347);
and U6794 (N_6794,N_6537,N_6529);
nand U6795 (N_6795,N_6444,N_6535);
and U6796 (N_6796,N_6554,N_6682);
xor U6797 (N_6797,N_6524,N_6292);
nand U6798 (N_6798,N_6212,N_6613);
xnor U6799 (N_6799,N_6744,N_6247);
nand U6800 (N_6800,N_6103,N_6011);
nor U6801 (N_6801,N_6035,N_6706);
nor U6802 (N_6802,N_6170,N_6536);
or U6803 (N_6803,N_6120,N_6672);
nor U6804 (N_6804,N_6585,N_6335);
or U6805 (N_6805,N_6248,N_6506);
and U6806 (N_6806,N_6690,N_6711);
nor U6807 (N_6807,N_6256,N_6322);
nor U6808 (N_6808,N_6459,N_6265);
nor U6809 (N_6809,N_6155,N_6330);
nor U6810 (N_6810,N_6504,N_6484);
and U6811 (N_6811,N_6195,N_6326);
or U6812 (N_6812,N_6231,N_6619);
nand U6813 (N_6813,N_6083,N_6424);
nand U6814 (N_6814,N_6057,N_6220);
nand U6815 (N_6815,N_6387,N_6062);
nor U6816 (N_6816,N_6650,N_6362);
nor U6817 (N_6817,N_6366,N_6709);
or U6818 (N_6818,N_6287,N_6436);
or U6819 (N_6819,N_6040,N_6148);
nand U6820 (N_6820,N_6409,N_6065);
xnor U6821 (N_6821,N_6646,N_6270);
and U6822 (N_6822,N_6331,N_6199);
nor U6823 (N_6823,N_6311,N_6441);
nand U6824 (N_6824,N_6556,N_6204);
nor U6825 (N_6825,N_6435,N_6294);
and U6826 (N_6826,N_6416,N_6216);
nand U6827 (N_6827,N_6080,N_6186);
and U6828 (N_6828,N_6488,N_6047);
xnor U6829 (N_6829,N_6676,N_6099);
nand U6830 (N_6830,N_6289,N_6230);
nor U6831 (N_6831,N_6066,N_6667);
or U6832 (N_6832,N_6527,N_6604);
and U6833 (N_6833,N_6607,N_6070);
and U6834 (N_6834,N_6087,N_6470);
or U6835 (N_6835,N_6340,N_6319);
nor U6836 (N_6836,N_6722,N_6560);
nand U6837 (N_6837,N_6582,N_6726);
nand U6838 (N_6838,N_6390,N_6151);
nand U6839 (N_6839,N_6670,N_6732);
and U6840 (N_6840,N_6200,N_6262);
nand U6841 (N_6841,N_6073,N_6606);
nand U6842 (N_6842,N_6438,N_6593);
or U6843 (N_6843,N_6015,N_6244);
or U6844 (N_6844,N_6081,N_6475);
nand U6845 (N_6845,N_6312,N_6005);
nand U6846 (N_6846,N_6564,N_6514);
nor U6847 (N_6847,N_6222,N_6668);
nor U6848 (N_6848,N_6735,N_6356);
and U6849 (N_6849,N_6145,N_6558);
nor U6850 (N_6850,N_6046,N_6703);
nor U6851 (N_6851,N_6632,N_6101);
or U6852 (N_6852,N_6707,N_6091);
and U6853 (N_6853,N_6385,N_6666);
nor U6854 (N_6854,N_6215,N_6396);
nor U6855 (N_6855,N_6146,N_6563);
nor U6856 (N_6856,N_6386,N_6327);
xor U6857 (N_6857,N_6136,N_6689);
nor U6858 (N_6858,N_6384,N_6662);
nand U6859 (N_6859,N_6609,N_6337);
nor U6860 (N_6860,N_6532,N_6180);
or U6861 (N_6861,N_6392,N_6197);
nand U6862 (N_6862,N_6079,N_6539);
nand U6863 (N_6863,N_6586,N_6365);
nor U6864 (N_6864,N_6157,N_6377);
or U6865 (N_6865,N_6596,N_6022);
or U6866 (N_6866,N_6112,N_6738);
xnor U6867 (N_6867,N_6360,N_6051);
nand U6868 (N_6868,N_6526,N_6024);
xor U6869 (N_6869,N_6510,N_6261);
nand U6870 (N_6870,N_6241,N_6020);
nor U6871 (N_6871,N_6277,N_6633);
xor U6872 (N_6872,N_6259,N_6404);
and U6873 (N_6873,N_6297,N_6368);
and U6874 (N_6874,N_6654,N_6658);
and U6875 (N_6875,N_6276,N_6250);
nand U6876 (N_6876,N_6480,N_6116);
or U6877 (N_6877,N_6631,N_6458);
or U6878 (N_6878,N_6394,N_6234);
nand U6879 (N_6879,N_6742,N_6267);
nor U6880 (N_6880,N_6665,N_6421);
nor U6881 (N_6881,N_6205,N_6627);
nor U6882 (N_6882,N_6023,N_6402);
and U6883 (N_6883,N_6476,N_6466);
nand U6884 (N_6884,N_6640,N_6555);
nand U6885 (N_6885,N_6161,N_6072);
xnor U6886 (N_6886,N_6511,N_6692);
or U6887 (N_6887,N_6339,N_6521);
nand U6888 (N_6888,N_6229,N_6489);
nor U6889 (N_6889,N_6168,N_6178);
nand U6890 (N_6890,N_6280,N_6746);
and U6891 (N_6891,N_6669,N_6219);
nand U6892 (N_6892,N_6055,N_6092);
nand U6893 (N_6893,N_6067,N_6184);
and U6894 (N_6894,N_6557,N_6473);
nand U6895 (N_6895,N_6042,N_6181);
nand U6896 (N_6896,N_6500,N_6121);
and U6897 (N_6897,N_6740,N_6001);
and U6898 (N_6898,N_6063,N_6704);
nor U6899 (N_6899,N_6352,N_6721);
nand U6900 (N_6900,N_6357,N_6160);
nor U6901 (N_6901,N_6291,N_6446);
and U6902 (N_6902,N_6411,N_6034);
nand U6903 (N_6903,N_6592,N_6638);
nor U6904 (N_6904,N_6038,N_6725);
and U6905 (N_6905,N_6054,N_6460);
xor U6906 (N_6906,N_6236,N_6541);
nor U6907 (N_6907,N_6418,N_6508);
nor U6908 (N_6908,N_6630,N_6224);
nand U6909 (N_6909,N_6739,N_6718);
nor U6910 (N_6910,N_6320,N_6004);
nand U6911 (N_6911,N_6696,N_6678);
nand U6912 (N_6912,N_6567,N_6232);
and U6913 (N_6913,N_6251,N_6730);
nand U6914 (N_6914,N_6501,N_6114);
nand U6915 (N_6915,N_6263,N_6053);
nand U6916 (N_6916,N_6479,N_6295);
and U6917 (N_6917,N_6429,N_6071);
and U6918 (N_6918,N_6693,N_6334);
and U6919 (N_6919,N_6454,N_6393);
and U6920 (N_6920,N_6448,N_6445);
nand U6921 (N_6921,N_6715,N_6552);
nor U6922 (N_6922,N_6305,N_6321);
and U6923 (N_6923,N_6450,N_6573);
xnor U6924 (N_6924,N_6492,N_6648);
xor U6925 (N_6925,N_6481,N_6434);
nand U6926 (N_6926,N_6187,N_6174);
xor U6927 (N_6927,N_6611,N_6210);
or U6928 (N_6928,N_6243,N_6749);
and U6929 (N_6929,N_6674,N_6061);
nand U6930 (N_6930,N_6716,N_6026);
nand U6931 (N_6931,N_6502,N_6452);
nand U6932 (N_6932,N_6094,N_6310);
or U6933 (N_6933,N_6000,N_6509);
xnor U6934 (N_6934,N_6565,N_6086);
or U6935 (N_6935,N_6483,N_6708);
nor U6936 (N_6936,N_6534,N_6084);
nand U6937 (N_6937,N_6477,N_6680);
and U6938 (N_6938,N_6380,N_6106);
and U6939 (N_6939,N_6068,N_6354);
nand U6940 (N_6940,N_6017,N_6497);
xor U6941 (N_6941,N_6123,N_6614);
nand U6942 (N_6942,N_6538,N_6202);
or U6943 (N_6943,N_6423,N_6315);
nand U6944 (N_6944,N_6561,N_6296);
and U6945 (N_6945,N_6165,N_6175);
and U6946 (N_6946,N_6218,N_6085);
or U6947 (N_6947,N_6495,N_6089);
nand U6948 (N_6948,N_6655,N_6717);
nand U6949 (N_6949,N_6714,N_6088);
nor U6950 (N_6950,N_6237,N_6498);
xor U6951 (N_6951,N_6007,N_6043);
or U6952 (N_6952,N_6491,N_6128);
xor U6953 (N_6953,N_6406,N_6144);
and U6954 (N_6954,N_6284,N_6133);
and U6955 (N_6955,N_6603,N_6443);
nor U6956 (N_6956,N_6333,N_6052);
nand U6957 (N_6957,N_6553,N_6622);
xor U6958 (N_6958,N_6275,N_6343);
nor U6959 (N_6959,N_6542,N_6142);
nor U6960 (N_6960,N_6041,N_6257);
or U6961 (N_6961,N_6132,N_6615);
nand U6962 (N_6962,N_6143,N_6713);
and U6963 (N_6963,N_6138,N_6719);
and U6964 (N_6964,N_6139,N_6269);
nand U6965 (N_6965,N_6016,N_6652);
or U6966 (N_6966,N_6030,N_6449);
nand U6967 (N_6967,N_6728,N_6286);
and U6968 (N_6968,N_6685,N_6313);
xnor U6969 (N_6969,N_6624,N_6253);
or U6970 (N_6970,N_6268,N_6008);
and U6971 (N_6971,N_6478,N_6580);
or U6972 (N_6972,N_6644,N_6414);
nand U6973 (N_6973,N_6374,N_6264);
or U6974 (N_6974,N_6117,N_6570);
and U6975 (N_6975,N_6637,N_6686);
xor U6976 (N_6976,N_6169,N_6568);
nor U6977 (N_6977,N_6353,N_6507);
nor U6978 (N_6978,N_6664,N_6741);
nor U6979 (N_6979,N_6468,N_6300);
nand U6980 (N_6980,N_6548,N_6358);
or U6981 (N_6981,N_6671,N_6048);
or U6982 (N_6982,N_6629,N_6162);
xnor U6983 (N_6983,N_6141,N_6442);
nand U6984 (N_6984,N_6167,N_6684);
and U6985 (N_6985,N_6661,N_6663);
nor U6986 (N_6986,N_6107,N_6413);
xor U6987 (N_6987,N_6724,N_6486);
nand U6988 (N_6988,N_6517,N_6641);
and U6989 (N_6989,N_6639,N_6285);
nor U6990 (N_6990,N_6577,N_6597);
xor U6991 (N_6991,N_6104,N_6433);
nor U6992 (N_6992,N_6598,N_6490);
nor U6993 (N_6993,N_6350,N_6523);
and U6994 (N_6994,N_6355,N_6395);
nor U6995 (N_6995,N_6499,N_6456);
nand U6996 (N_6996,N_6032,N_6096);
and U6997 (N_6997,N_6274,N_6102);
or U6998 (N_6998,N_6688,N_6656);
nor U6999 (N_6999,N_6075,N_6345);
nor U7000 (N_7000,N_6074,N_6290);
nor U7001 (N_7001,N_6095,N_6308);
nor U7002 (N_7002,N_6298,N_6591);
or U7003 (N_7003,N_6125,N_6628);
or U7004 (N_7004,N_6018,N_6108);
nand U7005 (N_7005,N_6462,N_6003);
nor U7006 (N_7006,N_6172,N_6594);
or U7007 (N_7007,N_6515,N_6683);
nand U7008 (N_7008,N_6059,N_6031);
and U7009 (N_7009,N_6213,N_6616);
nand U7010 (N_7010,N_6583,N_6453);
nor U7011 (N_7011,N_6617,N_6533);
nand U7012 (N_7012,N_6060,N_6137);
nand U7013 (N_7013,N_6013,N_6519);
xnor U7014 (N_7014,N_6518,N_6077);
nor U7015 (N_7015,N_6610,N_6225);
nand U7016 (N_7016,N_6316,N_6221);
nor U7017 (N_7017,N_6194,N_6348);
nand U7018 (N_7018,N_6279,N_6729);
and U7019 (N_7019,N_6164,N_6451);
or U7020 (N_7020,N_6388,N_6505);
and U7021 (N_7021,N_6019,N_6159);
nor U7022 (N_7022,N_6496,N_6679);
or U7023 (N_7023,N_6589,N_6467);
nor U7024 (N_7024,N_6620,N_6182);
or U7025 (N_7025,N_6156,N_6705);
nand U7026 (N_7026,N_6645,N_6154);
or U7027 (N_7027,N_6516,N_6379);
nand U7028 (N_7028,N_6605,N_6173);
and U7029 (N_7029,N_6135,N_6188);
and U7030 (N_7030,N_6400,N_6428);
or U7031 (N_7031,N_6158,N_6673);
xor U7032 (N_7032,N_6282,N_6299);
and U7033 (N_7033,N_6196,N_6642);
xnor U7034 (N_7034,N_6736,N_6027);
nand U7035 (N_7035,N_6332,N_6371);
nand U7036 (N_7036,N_6152,N_6342);
and U7037 (N_7037,N_6214,N_6364);
nor U7038 (N_7038,N_6512,N_6238);
nor U7039 (N_7039,N_6209,N_6734);
nand U7040 (N_7040,N_6543,N_6344);
nand U7041 (N_7041,N_6463,N_6513);
nor U7042 (N_7042,N_6049,N_6177);
nor U7043 (N_7043,N_6702,N_6447);
nand U7044 (N_7044,N_6677,N_6307);
nand U7045 (N_7045,N_6587,N_6147);
nand U7046 (N_7046,N_6425,N_6439);
or U7047 (N_7047,N_6064,N_6440);
nand U7048 (N_7048,N_6540,N_6012);
and U7049 (N_7049,N_6206,N_6550);
and U7050 (N_7050,N_6069,N_6273);
nor U7051 (N_7051,N_6126,N_6260);
nor U7052 (N_7052,N_6176,N_6191);
or U7053 (N_7053,N_6601,N_6266);
and U7054 (N_7054,N_6712,N_6185);
and U7055 (N_7055,N_6412,N_6602);
and U7056 (N_7056,N_6657,N_6226);
nor U7057 (N_7057,N_6118,N_6699);
and U7058 (N_7058,N_6329,N_6571);
and U7059 (N_7059,N_6626,N_6608);
xnor U7060 (N_7060,N_6363,N_6090);
nand U7061 (N_7061,N_6278,N_6115);
nand U7062 (N_7062,N_6361,N_6288);
xor U7063 (N_7063,N_6408,N_6239);
nor U7064 (N_7064,N_6525,N_6082);
and U7065 (N_7065,N_6119,N_6687);
or U7066 (N_7066,N_6050,N_6098);
nor U7067 (N_7067,N_6482,N_6643);
nand U7068 (N_7068,N_6748,N_6398);
nor U7069 (N_7069,N_6228,N_6056);
nor U7070 (N_7070,N_6150,N_6745);
and U7071 (N_7071,N_6134,N_6457);
or U7072 (N_7072,N_6010,N_6651);
and U7073 (N_7073,N_6625,N_6021);
and U7074 (N_7074,N_6430,N_6163);
or U7075 (N_7075,N_6113,N_6211);
and U7076 (N_7076,N_6179,N_6217);
and U7077 (N_7077,N_6691,N_6100);
and U7078 (N_7078,N_6009,N_6600);
and U7079 (N_7079,N_6595,N_6369);
xor U7080 (N_7080,N_6419,N_6006);
xnor U7081 (N_7081,N_6649,N_6618);
nand U7082 (N_7082,N_6710,N_6127);
nor U7083 (N_7083,N_6149,N_6314);
and U7084 (N_7084,N_6391,N_6551);
or U7085 (N_7085,N_6698,N_6531);
nand U7086 (N_7086,N_6304,N_6544);
nor U7087 (N_7087,N_6122,N_6272);
or U7088 (N_7088,N_6301,N_6731);
and U7089 (N_7089,N_6341,N_6432);
nor U7090 (N_7090,N_6410,N_6723);
nand U7091 (N_7091,N_6153,N_6493);
or U7092 (N_7092,N_6465,N_6743);
xnor U7093 (N_7093,N_6336,N_6317);
xor U7094 (N_7094,N_6700,N_6325);
or U7095 (N_7095,N_6129,N_6093);
or U7096 (N_7096,N_6078,N_6562);
and U7097 (N_7097,N_6547,N_6397);
or U7098 (N_7098,N_6522,N_6346);
xnor U7099 (N_7099,N_6166,N_6471);
nor U7100 (N_7100,N_6171,N_6111);
nand U7101 (N_7101,N_6494,N_6233);
nand U7102 (N_7102,N_6029,N_6694);
or U7103 (N_7103,N_6246,N_6255);
nand U7104 (N_7104,N_6383,N_6044);
and U7105 (N_7105,N_6131,N_6014);
or U7106 (N_7106,N_6503,N_6189);
or U7107 (N_7107,N_6701,N_6370);
and U7108 (N_7108,N_6376,N_6653);
or U7109 (N_7109,N_6235,N_6037);
nand U7110 (N_7110,N_6373,N_6203);
nand U7111 (N_7111,N_6647,N_6105);
nor U7112 (N_7112,N_6623,N_6546);
nand U7113 (N_7113,N_6201,N_6306);
and U7114 (N_7114,N_6039,N_6309);
or U7115 (N_7115,N_6659,N_6574);
and U7116 (N_7116,N_6634,N_6328);
nor U7117 (N_7117,N_6033,N_6349);
and U7118 (N_7118,N_6420,N_6140);
nor U7119 (N_7119,N_6405,N_6281);
nand U7120 (N_7120,N_6318,N_6737);
and U7121 (N_7121,N_6002,N_6520);
nand U7122 (N_7122,N_6324,N_6549);
or U7123 (N_7123,N_6575,N_6426);
nor U7124 (N_7124,N_6733,N_6727);
and U7125 (N_7125,N_6696,N_6326);
and U7126 (N_7126,N_6192,N_6230);
xnor U7127 (N_7127,N_6530,N_6200);
and U7128 (N_7128,N_6605,N_6416);
and U7129 (N_7129,N_6289,N_6648);
nor U7130 (N_7130,N_6692,N_6121);
nand U7131 (N_7131,N_6260,N_6205);
and U7132 (N_7132,N_6214,N_6152);
nand U7133 (N_7133,N_6238,N_6498);
xnor U7134 (N_7134,N_6340,N_6260);
nor U7135 (N_7135,N_6599,N_6051);
or U7136 (N_7136,N_6689,N_6550);
nor U7137 (N_7137,N_6519,N_6681);
nor U7138 (N_7138,N_6084,N_6651);
nand U7139 (N_7139,N_6363,N_6508);
nand U7140 (N_7140,N_6551,N_6223);
nor U7141 (N_7141,N_6237,N_6597);
nand U7142 (N_7142,N_6173,N_6098);
and U7143 (N_7143,N_6332,N_6405);
or U7144 (N_7144,N_6601,N_6081);
nand U7145 (N_7145,N_6168,N_6511);
nor U7146 (N_7146,N_6668,N_6301);
or U7147 (N_7147,N_6250,N_6619);
nor U7148 (N_7148,N_6384,N_6589);
nand U7149 (N_7149,N_6598,N_6330);
nand U7150 (N_7150,N_6225,N_6062);
and U7151 (N_7151,N_6070,N_6640);
nor U7152 (N_7152,N_6543,N_6032);
xor U7153 (N_7153,N_6396,N_6659);
and U7154 (N_7154,N_6415,N_6004);
nor U7155 (N_7155,N_6551,N_6670);
and U7156 (N_7156,N_6648,N_6575);
or U7157 (N_7157,N_6424,N_6033);
or U7158 (N_7158,N_6247,N_6163);
xor U7159 (N_7159,N_6679,N_6211);
or U7160 (N_7160,N_6449,N_6571);
and U7161 (N_7161,N_6057,N_6722);
or U7162 (N_7162,N_6623,N_6209);
and U7163 (N_7163,N_6524,N_6707);
and U7164 (N_7164,N_6675,N_6296);
nand U7165 (N_7165,N_6692,N_6260);
nand U7166 (N_7166,N_6146,N_6550);
or U7167 (N_7167,N_6629,N_6503);
or U7168 (N_7168,N_6714,N_6207);
or U7169 (N_7169,N_6223,N_6563);
nand U7170 (N_7170,N_6582,N_6677);
nor U7171 (N_7171,N_6427,N_6673);
nor U7172 (N_7172,N_6112,N_6649);
nor U7173 (N_7173,N_6712,N_6470);
and U7174 (N_7174,N_6329,N_6660);
nand U7175 (N_7175,N_6300,N_6644);
or U7176 (N_7176,N_6334,N_6679);
and U7177 (N_7177,N_6088,N_6296);
and U7178 (N_7178,N_6745,N_6147);
and U7179 (N_7179,N_6735,N_6087);
nor U7180 (N_7180,N_6699,N_6397);
or U7181 (N_7181,N_6333,N_6322);
nand U7182 (N_7182,N_6283,N_6376);
or U7183 (N_7183,N_6039,N_6441);
or U7184 (N_7184,N_6285,N_6001);
and U7185 (N_7185,N_6414,N_6544);
or U7186 (N_7186,N_6198,N_6597);
or U7187 (N_7187,N_6151,N_6509);
xnor U7188 (N_7188,N_6493,N_6110);
and U7189 (N_7189,N_6487,N_6040);
nor U7190 (N_7190,N_6098,N_6016);
nand U7191 (N_7191,N_6098,N_6015);
nand U7192 (N_7192,N_6084,N_6422);
nand U7193 (N_7193,N_6097,N_6720);
nor U7194 (N_7194,N_6193,N_6658);
xnor U7195 (N_7195,N_6627,N_6626);
nor U7196 (N_7196,N_6447,N_6078);
nand U7197 (N_7197,N_6436,N_6291);
nand U7198 (N_7198,N_6437,N_6330);
or U7199 (N_7199,N_6341,N_6311);
xnor U7200 (N_7200,N_6617,N_6594);
or U7201 (N_7201,N_6434,N_6348);
and U7202 (N_7202,N_6550,N_6557);
xnor U7203 (N_7203,N_6316,N_6715);
and U7204 (N_7204,N_6099,N_6092);
nor U7205 (N_7205,N_6299,N_6033);
or U7206 (N_7206,N_6669,N_6243);
nand U7207 (N_7207,N_6236,N_6694);
nand U7208 (N_7208,N_6602,N_6148);
nor U7209 (N_7209,N_6118,N_6318);
or U7210 (N_7210,N_6023,N_6544);
and U7211 (N_7211,N_6298,N_6109);
or U7212 (N_7212,N_6046,N_6064);
nand U7213 (N_7213,N_6589,N_6514);
nor U7214 (N_7214,N_6014,N_6702);
and U7215 (N_7215,N_6330,N_6133);
or U7216 (N_7216,N_6637,N_6519);
xor U7217 (N_7217,N_6369,N_6281);
or U7218 (N_7218,N_6687,N_6156);
nor U7219 (N_7219,N_6563,N_6469);
and U7220 (N_7220,N_6584,N_6159);
or U7221 (N_7221,N_6421,N_6743);
or U7222 (N_7222,N_6714,N_6681);
nor U7223 (N_7223,N_6295,N_6710);
nor U7224 (N_7224,N_6228,N_6512);
xor U7225 (N_7225,N_6700,N_6336);
nand U7226 (N_7226,N_6100,N_6273);
or U7227 (N_7227,N_6741,N_6512);
xor U7228 (N_7228,N_6145,N_6602);
or U7229 (N_7229,N_6350,N_6333);
nand U7230 (N_7230,N_6118,N_6422);
and U7231 (N_7231,N_6161,N_6412);
nor U7232 (N_7232,N_6075,N_6495);
nand U7233 (N_7233,N_6135,N_6335);
nor U7234 (N_7234,N_6551,N_6005);
nor U7235 (N_7235,N_6067,N_6657);
xnor U7236 (N_7236,N_6130,N_6669);
and U7237 (N_7237,N_6349,N_6452);
nor U7238 (N_7238,N_6730,N_6100);
and U7239 (N_7239,N_6137,N_6522);
nand U7240 (N_7240,N_6047,N_6126);
or U7241 (N_7241,N_6519,N_6061);
nand U7242 (N_7242,N_6406,N_6188);
or U7243 (N_7243,N_6148,N_6071);
xor U7244 (N_7244,N_6717,N_6596);
nor U7245 (N_7245,N_6429,N_6723);
nor U7246 (N_7246,N_6275,N_6062);
nor U7247 (N_7247,N_6410,N_6145);
or U7248 (N_7248,N_6748,N_6463);
nand U7249 (N_7249,N_6658,N_6620);
nand U7250 (N_7250,N_6557,N_6654);
nand U7251 (N_7251,N_6357,N_6741);
and U7252 (N_7252,N_6299,N_6478);
nand U7253 (N_7253,N_6168,N_6030);
nor U7254 (N_7254,N_6589,N_6123);
nor U7255 (N_7255,N_6617,N_6226);
nor U7256 (N_7256,N_6040,N_6077);
or U7257 (N_7257,N_6650,N_6593);
nor U7258 (N_7258,N_6704,N_6019);
or U7259 (N_7259,N_6228,N_6083);
nand U7260 (N_7260,N_6603,N_6358);
nor U7261 (N_7261,N_6624,N_6361);
or U7262 (N_7262,N_6469,N_6672);
nor U7263 (N_7263,N_6167,N_6142);
xor U7264 (N_7264,N_6550,N_6003);
nor U7265 (N_7265,N_6332,N_6103);
or U7266 (N_7266,N_6287,N_6045);
nand U7267 (N_7267,N_6664,N_6612);
nand U7268 (N_7268,N_6058,N_6117);
nand U7269 (N_7269,N_6723,N_6121);
xor U7270 (N_7270,N_6018,N_6029);
nor U7271 (N_7271,N_6595,N_6493);
nand U7272 (N_7272,N_6161,N_6699);
nand U7273 (N_7273,N_6086,N_6225);
nor U7274 (N_7274,N_6514,N_6289);
or U7275 (N_7275,N_6619,N_6262);
and U7276 (N_7276,N_6709,N_6612);
or U7277 (N_7277,N_6190,N_6023);
and U7278 (N_7278,N_6207,N_6456);
or U7279 (N_7279,N_6327,N_6230);
nor U7280 (N_7280,N_6507,N_6485);
nor U7281 (N_7281,N_6655,N_6592);
nor U7282 (N_7282,N_6468,N_6650);
nor U7283 (N_7283,N_6691,N_6620);
nand U7284 (N_7284,N_6187,N_6666);
and U7285 (N_7285,N_6202,N_6611);
or U7286 (N_7286,N_6550,N_6125);
nor U7287 (N_7287,N_6337,N_6075);
nor U7288 (N_7288,N_6046,N_6251);
or U7289 (N_7289,N_6627,N_6252);
or U7290 (N_7290,N_6207,N_6712);
or U7291 (N_7291,N_6598,N_6074);
nand U7292 (N_7292,N_6209,N_6004);
nor U7293 (N_7293,N_6198,N_6347);
and U7294 (N_7294,N_6674,N_6262);
nand U7295 (N_7295,N_6032,N_6661);
nor U7296 (N_7296,N_6506,N_6228);
nor U7297 (N_7297,N_6424,N_6055);
or U7298 (N_7298,N_6153,N_6662);
xor U7299 (N_7299,N_6034,N_6740);
nor U7300 (N_7300,N_6467,N_6273);
or U7301 (N_7301,N_6100,N_6248);
nand U7302 (N_7302,N_6256,N_6282);
or U7303 (N_7303,N_6648,N_6257);
xnor U7304 (N_7304,N_6331,N_6673);
nor U7305 (N_7305,N_6673,N_6670);
nor U7306 (N_7306,N_6310,N_6464);
and U7307 (N_7307,N_6070,N_6198);
nor U7308 (N_7308,N_6574,N_6049);
and U7309 (N_7309,N_6043,N_6530);
nor U7310 (N_7310,N_6020,N_6630);
nor U7311 (N_7311,N_6084,N_6349);
nand U7312 (N_7312,N_6603,N_6513);
nor U7313 (N_7313,N_6654,N_6443);
nor U7314 (N_7314,N_6325,N_6575);
nand U7315 (N_7315,N_6497,N_6564);
nor U7316 (N_7316,N_6358,N_6242);
and U7317 (N_7317,N_6535,N_6206);
and U7318 (N_7318,N_6382,N_6220);
nor U7319 (N_7319,N_6661,N_6210);
nor U7320 (N_7320,N_6606,N_6213);
and U7321 (N_7321,N_6175,N_6514);
nand U7322 (N_7322,N_6540,N_6631);
nor U7323 (N_7323,N_6054,N_6669);
nor U7324 (N_7324,N_6071,N_6449);
and U7325 (N_7325,N_6581,N_6141);
nor U7326 (N_7326,N_6269,N_6001);
and U7327 (N_7327,N_6650,N_6387);
xnor U7328 (N_7328,N_6675,N_6189);
and U7329 (N_7329,N_6122,N_6315);
and U7330 (N_7330,N_6656,N_6744);
or U7331 (N_7331,N_6203,N_6726);
nor U7332 (N_7332,N_6685,N_6156);
nor U7333 (N_7333,N_6294,N_6207);
and U7334 (N_7334,N_6611,N_6264);
or U7335 (N_7335,N_6083,N_6303);
nand U7336 (N_7336,N_6124,N_6475);
and U7337 (N_7337,N_6251,N_6014);
and U7338 (N_7338,N_6162,N_6747);
and U7339 (N_7339,N_6278,N_6310);
xor U7340 (N_7340,N_6455,N_6587);
nor U7341 (N_7341,N_6601,N_6749);
nor U7342 (N_7342,N_6206,N_6498);
or U7343 (N_7343,N_6083,N_6556);
nor U7344 (N_7344,N_6189,N_6459);
nor U7345 (N_7345,N_6062,N_6696);
nor U7346 (N_7346,N_6141,N_6447);
nand U7347 (N_7347,N_6392,N_6298);
nor U7348 (N_7348,N_6653,N_6482);
or U7349 (N_7349,N_6304,N_6089);
or U7350 (N_7350,N_6304,N_6734);
xnor U7351 (N_7351,N_6122,N_6104);
and U7352 (N_7352,N_6093,N_6640);
nor U7353 (N_7353,N_6215,N_6330);
nor U7354 (N_7354,N_6156,N_6365);
or U7355 (N_7355,N_6190,N_6548);
nor U7356 (N_7356,N_6429,N_6408);
nand U7357 (N_7357,N_6406,N_6453);
or U7358 (N_7358,N_6618,N_6674);
or U7359 (N_7359,N_6154,N_6075);
nor U7360 (N_7360,N_6598,N_6561);
nor U7361 (N_7361,N_6142,N_6502);
nor U7362 (N_7362,N_6228,N_6294);
or U7363 (N_7363,N_6494,N_6155);
or U7364 (N_7364,N_6310,N_6593);
nor U7365 (N_7365,N_6225,N_6383);
and U7366 (N_7366,N_6089,N_6474);
xor U7367 (N_7367,N_6580,N_6024);
nor U7368 (N_7368,N_6164,N_6554);
nor U7369 (N_7369,N_6375,N_6448);
nor U7370 (N_7370,N_6394,N_6047);
or U7371 (N_7371,N_6742,N_6699);
nor U7372 (N_7372,N_6022,N_6424);
or U7373 (N_7373,N_6670,N_6284);
nand U7374 (N_7374,N_6316,N_6188);
nand U7375 (N_7375,N_6292,N_6085);
or U7376 (N_7376,N_6588,N_6672);
nand U7377 (N_7377,N_6619,N_6551);
or U7378 (N_7378,N_6465,N_6495);
nor U7379 (N_7379,N_6295,N_6127);
nand U7380 (N_7380,N_6326,N_6617);
or U7381 (N_7381,N_6128,N_6552);
nor U7382 (N_7382,N_6009,N_6251);
or U7383 (N_7383,N_6435,N_6481);
and U7384 (N_7384,N_6185,N_6027);
and U7385 (N_7385,N_6431,N_6163);
xor U7386 (N_7386,N_6004,N_6028);
nand U7387 (N_7387,N_6218,N_6304);
nor U7388 (N_7388,N_6433,N_6152);
or U7389 (N_7389,N_6444,N_6090);
xor U7390 (N_7390,N_6164,N_6383);
nor U7391 (N_7391,N_6742,N_6272);
nor U7392 (N_7392,N_6511,N_6469);
nor U7393 (N_7393,N_6544,N_6084);
and U7394 (N_7394,N_6573,N_6329);
nand U7395 (N_7395,N_6703,N_6517);
and U7396 (N_7396,N_6216,N_6655);
nand U7397 (N_7397,N_6114,N_6512);
and U7398 (N_7398,N_6598,N_6372);
xor U7399 (N_7399,N_6213,N_6581);
or U7400 (N_7400,N_6513,N_6069);
nor U7401 (N_7401,N_6373,N_6422);
nand U7402 (N_7402,N_6737,N_6725);
nand U7403 (N_7403,N_6586,N_6482);
nand U7404 (N_7404,N_6291,N_6581);
xor U7405 (N_7405,N_6178,N_6555);
nor U7406 (N_7406,N_6398,N_6407);
or U7407 (N_7407,N_6093,N_6651);
xnor U7408 (N_7408,N_6157,N_6131);
nor U7409 (N_7409,N_6249,N_6138);
xnor U7410 (N_7410,N_6528,N_6220);
or U7411 (N_7411,N_6683,N_6285);
or U7412 (N_7412,N_6688,N_6139);
and U7413 (N_7413,N_6577,N_6579);
and U7414 (N_7414,N_6248,N_6519);
xnor U7415 (N_7415,N_6237,N_6126);
or U7416 (N_7416,N_6686,N_6291);
and U7417 (N_7417,N_6628,N_6709);
and U7418 (N_7418,N_6560,N_6095);
nor U7419 (N_7419,N_6520,N_6197);
nor U7420 (N_7420,N_6077,N_6583);
and U7421 (N_7421,N_6012,N_6315);
or U7422 (N_7422,N_6100,N_6027);
or U7423 (N_7423,N_6412,N_6528);
nor U7424 (N_7424,N_6341,N_6359);
nand U7425 (N_7425,N_6421,N_6163);
or U7426 (N_7426,N_6572,N_6253);
nor U7427 (N_7427,N_6323,N_6008);
nor U7428 (N_7428,N_6340,N_6358);
nor U7429 (N_7429,N_6415,N_6032);
nand U7430 (N_7430,N_6562,N_6466);
nor U7431 (N_7431,N_6302,N_6065);
or U7432 (N_7432,N_6685,N_6651);
nor U7433 (N_7433,N_6266,N_6717);
or U7434 (N_7434,N_6559,N_6707);
nand U7435 (N_7435,N_6332,N_6203);
and U7436 (N_7436,N_6622,N_6353);
and U7437 (N_7437,N_6656,N_6282);
nor U7438 (N_7438,N_6363,N_6695);
xnor U7439 (N_7439,N_6166,N_6233);
nand U7440 (N_7440,N_6478,N_6219);
or U7441 (N_7441,N_6613,N_6165);
xor U7442 (N_7442,N_6742,N_6605);
nor U7443 (N_7443,N_6213,N_6641);
and U7444 (N_7444,N_6322,N_6604);
and U7445 (N_7445,N_6211,N_6577);
or U7446 (N_7446,N_6036,N_6221);
nand U7447 (N_7447,N_6006,N_6390);
nor U7448 (N_7448,N_6204,N_6301);
nor U7449 (N_7449,N_6300,N_6320);
nand U7450 (N_7450,N_6382,N_6059);
and U7451 (N_7451,N_6625,N_6122);
and U7452 (N_7452,N_6080,N_6380);
nor U7453 (N_7453,N_6470,N_6343);
and U7454 (N_7454,N_6475,N_6702);
or U7455 (N_7455,N_6749,N_6090);
nand U7456 (N_7456,N_6140,N_6545);
xnor U7457 (N_7457,N_6648,N_6517);
xor U7458 (N_7458,N_6262,N_6128);
nand U7459 (N_7459,N_6168,N_6707);
nand U7460 (N_7460,N_6544,N_6283);
nand U7461 (N_7461,N_6362,N_6063);
and U7462 (N_7462,N_6614,N_6227);
nor U7463 (N_7463,N_6617,N_6512);
or U7464 (N_7464,N_6021,N_6742);
and U7465 (N_7465,N_6633,N_6441);
and U7466 (N_7466,N_6259,N_6116);
and U7467 (N_7467,N_6128,N_6329);
and U7468 (N_7468,N_6496,N_6477);
nor U7469 (N_7469,N_6637,N_6423);
or U7470 (N_7470,N_6448,N_6676);
nor U7471 (N_7471,N_6484,N_6551);
nand U7472 (N_7472,N_6596,N_6282);
and U7473 (N_7473,N_6501,N_6404);
nand U7474 (N_7474,N_6526,N_6732);
nand U7475 (N_7475,N_6434,N_6178);
and U7476 (N_7476,N_6725,N_6397);
xor U7477 (N_7477,N_6070,N_6538);
nor U7478 (N_7478,N_6747,N_6665);
nor U7479 (N_7479,N_6386,N_6118);
nor U7480 (N_7480,N_6161,N_6055);
and U7481 (N_7481,N_6526,N_6722);
nand U7482 (N_7482,N_6736,N_6364);
and U7483 (N_7483,N_6666,N_6321);
and U7484 (N_7484,N_6127,N_6655);
or U7485 (N_7485,N_6533,N_6574);
nor U7486 (N_7486,N_6105,N_6115);
and U7487 (N_7487,N_6108,N_6283);
nand U7488 (N_7488,N_6626,N_6140);
and U7489 (N_7489,N_6435,N_6469);
nand U7490 (N_7490,N_6631,N_6595);
nand U7491 (N_7491,N_6375,N_6635);
or U7492 (N_7492,N_6472,N_6583);
nor U7493 (N_7493,N_6048,N_6635);
nor U7494 (N_7494,N_6441,N_6479);
xor U7495 (N_7495,N_6539,N_6046);
nand U7496 (N_7496,N_6514,N_6222);
nor U7497 (N_7497,N_6536,N_6293);
nor U7498 (N_7498,N_6575,N_6002);
nor U7499 (N_7499,N_6632,N_6580);
nor U7500 (N_7500,N_6841,N_6932);
or U7501 (N_7501,N_7150,N_7142);
or U7502 (N_7502,N_7247,N_7061);
and U7503 (N_7503,N_7078,N_7235);
nor U7504 (N_7504,N_6783,N_7361);
nand U7505 (N_7505,N_7221,N_6938);
nand U7506 (N_7506,N_7376,N_7046);
or U7507 (N_7507,N_6795,N_6982);
and U7508 (N_7508,N_7284,N_7126);
or U7509 (N_7509,N_7302,N_6945);
or U7510 (N_7510,N_6865,N_7050);
nand U7511 (N_7511,N_6862,N_7122);
nor U7512 (N_7512,N_6825,N_6993);
and U7513 (N_7513,N_7269,N_7196);
and U7514 (N_7514,N_6782,N_7353);
nor U7515 (N_7515,N_6844,N_7044);
nor U7516 (N_7516,N_7365,N_7114);
nor U7517 (N_7517,N_7384,N_6920);
or U7518 (N_7518,N_7370,N_6870);
nand U7519 (N_7519,N_7256,N_7392);
and U7520 (N_7520,N_6959,N_7230);
or U7521 (N_7521,N_7319,N_7482);
and U7522 (N_7522,N_7424,N_6793);
nand U7523 (N_7523,N_7464,N_7296);
nand U7524 (N_7524,N_7032,N_6917);
nand U7525 (N_7525,N_7074,N_6986);
nor U7526 (N_7526,N_7314,N_6878);
nand U7527 (N_7527,N_7250,N_6815);
nor U7528 (N_7528,N_6985,N_7469);
nor U7529 (N_7529,N_7194,N_7245);
nand U7530 (N_7530,N_7372,N_7106);
nor U7531 (N_7531,N_7335,N_6944);
nor U7532 (N_7532,N_7233,N_7283);
nor U7533 (N_7533,N_6757,N_7060);
xor U7534 (N_7534,N_7393,N_7251);
or U7535 (N_7535,N_7022,N_7421);
and U7536 (N_7536,N_7079,N_7434);
nor U7537 (N_7537,N_7495,N_7192);
nand U7538 (N_7538,N_7068,N_7058);
xor U7539 (N_7539,N_7394,N_7193);
nand U7540 (N_7540,N_6758,N_7331);
xor U7541 (N_7541,N_7317,N_6752);
nand U7542 (N_7542,N_7410,N_7189);
nand U7543 (N_7543,N_7163,N_6765);
nor U7544 (N_7544,N_6873,N_6886);
or U7545 (N_7545,N_7213,N_7186);
nand U7546 (N_7546,N_7322,N_7379);
nand U7547 (N_7547,N_7128,N_7087);
nor U7548 (N_7548,N_7075,N_7414);
and U7549 (N_7549,N_7095,N_7131);
nand U7550 (N_7550,N_7404,N_6933);
and U7551 (N_7551,N_7030,N_7459);
nor U7552 (N_7552,N_6869,N_7497);
nand U7553 (N_7553,N_7318,N_7264);
nand U7554 (N_7554,N_7155,N_7214);
xnor U7555 (N_7555,N_7344,N_7279);
nor U7556 (N_7556,N_6810,N_7432);
xnor U7557 (N_7557,N_7368,N_6981);
and U7558 (N_7558,N_7282,N_7208);
or U7559 (N_7559,N_6805,N_6883);
nor U7560 (N_7560,N_6891,N_6750);
or U7561 (N_7561,N_6949,N_6832);
and U7562 (N_7562,N_7453,N_6973);
nand U7563 (N_7563,N_6848,N_6950);
nor U7564 (N_7564,N_7458,N_7490);
nand U7565 (N_7565,N_7113,N_6846);
nor U7566 (N_7566,N_7132,N_7456);
and U7567 (N_7567,N_7057,N_6858);
and U7568 (N_7568,N_6845,N_6751);
nor U7569 (N_7569,N_7146,N_6868);
or U7570 (N_7570,N_7172,N_7499);
nand U7571 (N_7571,N_7270,N_6799);
xor U7572 (N_7572,N_6953,N_7003);
or U7573 (N_7573,N_7134,N_7378);
or U7574 (N_7574,N_6818,N_7492);
or U7575 (N_7575,N_7124,N_7120);
or U7576 (N_7576,N_7479,N_7305);
nor U7577 (N_7577,N_7417,N_6759);
nand U7578 (N_7578,N_7449,N_6927);
or U7579 (N_7579,N_7455,N_6905);
nor U7580 (N_7580,N_7397,N_7367);
and U7581 (N_7581,N_6879,N_6764);
nand U7582 (N_7582,N_6866,N_7339);
nand U7583 (N_7583,N_7219,N_7280);
or U7584 (N_7584,N_7374,N_6937);
nor U7585 (N_7585,N_7486,N_7349);
and U7586 (N_7586,N_7211,N_7445);
xnor U7587 (N_7587,N_7175,N_7109);
nor U7588 (N_7588,N_7439,N_7203);
and U7589 (N_7589,N_6930,N_7165);
nand U7590 (N_7590,N_6943,N_7170);
nand U7591 (N_7591,N_7473,N_7364);
nand U7592 (N_7592,N_7152,N_6761);
nor U7593 (N_7593,N_7162,N_6874);
and U7594 (N_7594,N_7419,N_7225);
and U7595 (N_7595,N_7138,N_7090);
and U7596 (N_7596,N_7487,N_6753);
or U7597 (N_7597,N_6786,N_7156);
nor U7598 (N_7598,N_7045,N_7064);
and U7599 (N_7599,N_7014,N_7369);
and U7600 (N_7600,N_7043,N_7422);
and U7601 (N_7601,N_6888,N_7307);
or U7602 (N_7602,N_7098,N_6952);
nor U7603 (N_7603,N_6901,N_6894);
nand U7604 (N_7604,N_6822,N_7048);
nor U7605 (N_7605,N_7004,N_6881);
nand U7606 (N_7606,N_7388,N_6895);
or U7607 (N_7607,N_6833,N_7199);
nor U7608 (N_7608,N_7051,N_7005);
and U7609 (N_7609,N_6990,N_6942);
nand U7610 (N_7610,N_7412,N_7129);
or U7611 (N_7611,N_6871,N_6899);
and U7612 (N_7612,N_7047,N_7105);
xor U7613 (N_7613,N_7143,N_7085);
and U7614 (N_7614,N_7038,N_7164);
and U7615 (N_7615,N_6908,N_7431);
nand U7616 (N_7616,N_7351,N_7201);
or U7617 (N_7617,N_7340,N_6859);
nor U7618 (N_7618,N_6987,N_6853);
nand U7619 (N_7619,N_7321,N_7053);
nand U7620 (N_7620,N_7236,N_7415);
nand U7621 (N_7621,N_7182,N_7290);
nand U7622 (N_7622,N_7285,N_6762);
and U7623 (N_7623,N_7447,N_7080);
and U7624 (N_7624,N_7333,N_6787);
nand U7625 (N_7625,N_7463,N_7423);
and U7626 (N_7626,N_7466,N_7273);
nand U7627 (N_7627,N_6790,N_7151);
xnor U7628 (N_7628,N_6850,N_6922);
xnor U7629 (N_7629,N_6978,N_6893);
nor U7630 (N_7630,N_6966,N_6970);
nand U7631 (N_7631,N_6897,N_7418);
and U7632 (N_7632,N_7108,N_6926);
nand U7633 (N_7633,N_7145,N_7442);
nand U7634 (N_7634,N_6963,N_7386);
and U7635 (N_7635,N_6813,N_7117);
xnor U7636 (N_7636,N_7493,N_7357);
nand U7637 (N_7637,N_7116,N_6808);
or U7638 (N_7638,N_7382,N_6974);
nor U7639 (N_7639,N_7259,N_6941);
xnor U7640 (N_7640,N_7405,N_7293);
or U7641 (N_7641,N_6931,N_7013);
xnor U7642 (N_7642,N_7119,N_7012);
xor U7643 (N_7643,N_7347,N_6968);
or U7644 (N_7644,N_7470,N_6837);
nand U7645 (N_7645,N_6915,N_7222);
nand U7646 (N_7646,N_7480,N_7020);
nor U7647 (N_7647,N_6766,N_7308);
nor U7648 (N_7648,N_7026,N_7083);
and U7649 (N_7649,N_7402,N_7246);
nand U7650 (N_7650,N_6756,N_7169);
nand U7651 (N_7651,N_7437,N_6872);
or U7652 (N_7652,N_6887,N_6977);
nand U7653 (N_7653,N_7292,N_6877);
nor U7654 (N_7654,N_6817,N_6889);
nand U7655 (N_7655,N_7248,N_6957);
and U7656 (N_7656,N_7006,N_7063);
nand U7657 (N_7657,N_7297,N_7309);
or U7658 (N_7658,N_7157,N_6775);
or U7659 (N_7659,N_7103,N_7077);
nor U7660 (N_7660,N_6754,N_6827);
nor U7661 (N_7661,N_7016,N_6847);
or U7662 (N_7662,N_7149,N_6820);
or U7663 (N_7663,N_7457,N_6979);
nand U7664 (N_7664,N_7240,N_7252);
nor U7665 (N_7665,N_7179,N_7244);
nand U7666 (N_7666,N_7115,N_7190);
nand U7667 (N_7667,N_6856,N_6914);
nor U7668 (N_7668,N_7034,N_6851);
and U7669 (N_7669,N_7107,N_7158);
nand U7670 (N_7670,N_6773,N_6778);
and U7671 (N_7671,N_7183,N_7346);
nor U7672 (N_7672,N_7271,N_7135);
and U7673 (N_7673,N_7065,N_6999);
nor U7674 (N_7674,N_6967,N_7220);
or U7675 (N_7675,N_7121,N_6961);
nand U7676 (N_7676,N_7491,N_6983);
or U7677 (N_7677,N_6780,N_7413);
nand U7678 (N_7678,N_7380,N_6826);
nor U7679 (N_7679,N_7450,N_7461);
xor U7680 (N_7680,N_7072,N_7304);
and U7681 (N_7681,N_7133,N_7033);
or U7682 (N_7682,N_6956,N_6884);
xor U7683 (N_7683,N_7066,N_7411);
nand U7684 (N_7684,N_6940,N_7167);
or U7685 (N_7685,N_7427,N_7180);
nor U7686 (N_7686,N_7433,N_6836);
or U7687 (N_7687,N_7112,N_6767);
or U7688 (N_7688,N_7147,N_6791);
nand U7689 (N_7689,N_7471,N_6829);
xor U7690 (N_7690,N_7359,N_7184);
or U7691 (N_7691,N_7478,N_6924);
or U7692 (N_7692,N_6928,N_6760);
nand U7693 (N_7693,N_7130,N_7477);
nand U7694 (N_7694,N_7036,N_6876);
or U7695 (N_7695,N_7387,N_7281);
and U7696 (N_7696,N_6835,N_7300);
nand U7697 (N_7697,N_7452,N_7462);
nand U7698 (N_7698,N_6800,N_7336);
and U7699 (N_7699,N_7049,N_7390);
nor U7700 (N_7700,N_6902,N_7276);
and U7701 (N_7701,N_7081,N_7327);
and U7702 (N_7702,N_7375,N_7315);
nand U7703 (N_7703,N_6911,N_7311);
nand U7704 (N_7704,N_6936,N_7015);
nor U7705 (N_7705,N_7325,N_7377);
xor U7706 (N_7706,N_7323,N_7355);
xnor U7707 (N_7707,N_7084,N_6935);
nor U7708 (N_7708,N_6984,N_6925);
or U7709 (N_7709,N_7021,N_7239);
or U7710 (N_7710,N_7277,N_7139);
or U7711 (N_7711,N_7268,N_6838);
nor U7712 (N_7712,N_7088,N_7338);
nand U7713 (N_7713,N_7403,N_7154);
xor U7714 (N_7714,N_7056,N_7227);
nor U7715 (N_7715,N_6809,N_7354);
nand U7716 (N_7716,N_7254,N_7241);
xnor U7717 (N_7717,N_7260,N_6814);
nand U7718 (N_7718,N_7207,N_6890);
nand U7719 (N_7719,N_7195,N_7185);
and U7720 (N_7720,N_7391,N_7001);
xnor U7721 (N_7721,N_7018,N_6976);
nor U7722 (N_7722,N_6900,N_6802);
and U7723 (N_7723,N_6992,N_6830);
nor U7724 (N_7724,N_7011,N_7223);
nor U7725 (N_7725,N_6991,N_6807);
or U7726 (N_7726,N_7104,N_6896);
nor U7727 (N_7727,N_6801,N_7330);
xor U7728 (N_7728,N_7485,N_6972);
and U7729 (N_7729,N_6792,N_6763);
nand U7730 (N_7730,N_7481,N_7144);
nand U7731 (N_7731,N_6946,N_7266);
or U7732 (N_7732,N_7118,N_7215);
xnor U7733 (N_7733,N_7316,N_7031);
nand U7734 (N_7734,N_7262,N_6997);
nor U7735 (N_7735,N_6916,N_7301);
or U7736 (N_7736,N_6823,N_6785);
or U7737 (N_7737,N_7430,N_7204);
nand U7738 (N_7738,N_7234,N_7420);
nand U7739 (N_7739,N_6770,N_7363);
nor U7740 (N_7740,N_6919,N_7401);
and U7741 (N_7741,N_7249,N_6860);
nor U7742 (N_7742,N_6885,N_6768);
and U7743 (N_7743,N_7253,N_7009);
and U7744 (N_7744,N_6875,N_7099);
or U7745 (N_7745,N_7489,N_6852);
or U7746 (N_7746,N_7089,N_7127);
nor U7747 (N_7747,N_7035,N_7332);
nand U7748 (N_7748,N_6965,N_7298);
nor U7749 (N_7749,N_7062,N_7069);
or U7750 (N_7750,N_7029,N_7472);
nand U7751 (N_7751,N_7476,N_6995);
nor U7752 (N_7752,N_7100,N_7289);
nor U7753 (N_7753,N_7019,N_7288);
or U7754 (N_7754,N_7178,N_6923);
nor U7755 (N_7755,N_7295,N_7263);
and U7756 (N_7756,N_7362,N_7243);
nor U7757 (N_7757,N_7082,N_7177);
nor U7758 (N_7758,N_7070,N_7426);
nor U7759 (N_7759,N_7028,N_7460);
or U7760 (N_7760,N_7341,N_7443);
nor U7761 (N_7761,N_7409,N_7475);
nand U7762 (N_7762,N_7425,N_7086);
xnor U7763 (N_7763,N_6784,N_6788);
nand U7764 (N_7764,N_6777,N_6892);
nor U7765 (N_7765,N_6910,N_7352);
and U7766 (N_7766,N_7153,N_6996);
nand U7767 (N_7767,N_6939,N_7454);
or U7768 (N_7768,N_7174,N_7496);
nor U7769 (N_7769,N_6951,N_7039);
nand U7770 (N_7770,N_7188,N_6988);
and U7771 (N_7771,N_7111,N_6839);
nand U7772 (N_7772,N_6772,N_7176);
xnor U7773 (N_7773,N_7400,N_6796);
nand U7774 (N_7774,N_6904,N_7373);
or U7775 (N_7775,N_6824,N_7326);
nor U7776 (N_7776,N_7451,N_7218);
or U7777 (N_7777,N_7438,N_7209);
xor U7778 (N_7778,N_7498,N_7007);
nand U7779 (N_7779,N_6828,N_6994);
xnor U7780 (N_7780,N_7435,N_6840);
nand U7781 (N_7781,N_7017,N_7125);
nand U7782 (N_7782,N_7312,N_6779);
nor U7783 (N_7783,N_7303,N_6960);
and U7784 (N_7784,N_7294,N_7041);
nand U7785 (N_7785,N_6789,N_7395);
and U7786 (N_7786,N_7101,N_7212);
or U7787 (N_7787,N_7059,N_7343);
nand U7788 (N_7788,N_6958,N_7440);
and U7789 (N_7789,N_6771,N_7093);
and U7790 (N_7790,N_7141,N_7299);
and U7791 (N_7791,N_6834,N_6794);
or U7792 (N_7792,N_6804,N_7097);
and U7793 (N_7793,N_6929,N_7008);
nor U7794 (N_7794,N_7483,N_7474);
nand U7795 (N_7795,N_7024,N_7187);
nor U7796 (N_7796,N_7267,N_7073);
nand U7797 (N_7797,N_7446,N_7231);
xor U7798 (N_7798,N_7441,N_6909);
nor U7799 (N_7799,N_7025,N_7436);
nand U7800 (N_7800,N_7052,N_7076);
nand U7801 (N_7801,N_7287,N_7040);
nand U7802 (N_7802,N_7348,N_6964);
xnor U7803 (N_7803,N_7448,N_6855);
and U7804 (N_7804,N_7160,N_7027);
nand U7805 (N_7805,N_7275,N_6816);
xnor U7806 (N_7806,N_7398,N_7342);
and U7807 (N_7807,N_7054,N_6831);
nand U7808 (N_7808,N_7306,N_7310);
nand U7809 (N_7809,N_7313,N_7224);
nor U7810 (N_7810,N_7488,N_6861);
or U7811 (N_7811,N_7102,N_6755);
nor U7812 (N_7812,N_7173,N_7161);
nor U7813 (N_7813,N_7096,N_7444);
nor U7814 (N_7814,N_7261,N_7210);
or U7815 (N_7815,N_6948,N_6934);
nand U7816 (N_7816,N_7042,N_7094);
and U7817 (N_7817,N_6918,N_7345);
or U7818 (N_7818,N_6998,N_6797);
and U7819 (N_7819,N_6821,N_7371);
nor U7820 (N_7820,N_6954,N_7206);
or U7821 (N_7821,N_7328,N_7228);
xor U7822 (N_7822,N_7123,N_7202);
nand U7823 (N_7823,N_7484,N_6842);
or U7824 (N_7824,N_6798,N_7197);
nand U7825 (N_7825,N_7255,N_7200);
or U7826 (N_7826,N_7238,N_7092);
xnor U7827 (N_7827,N_7416,N_7037);
and U7828 (N_7828,N_7329,N_6913);
nand U7829 (N_7829,N_7265,N_7191);
xnor U7830 (N_7830,N_7429,N_6774);
and U7831 (N_7831,N_7205,N_7494);
nand U7832 (N_7832,N_7171,N_6921);
and U7833 (N_7833,N_7159,N_6849);
nand U7834 (N_7834,N_7399,N_7385);
or U7835 (N_7835,N_7010,N_7278);
or U7836 (N_7836,N_7140,N_7334);
or U7837 (N_7837,N_6903,N_7337);
or U7838 (N_7838,N_6947,N_7148);
or U7839 (N_7839,N_6843,N_7366);
nor U7840 (N_7840,N_7226,N_7383);
nor U7841 (N_7841,N_6912,N_7237);
or U7842 (N_7842,N_7406,N_6769);
nor U7843 (N_7843,N_6980,N_6857);
nor U7844 (N_7844,N_6806,N_7356);
and U7845 (N_7845,N_7000,N_6906);
and U7846 (N_7846,N_6803,N_7468);
nand U7847 (N_7847,N_6880,N_6898);
nand U7848 (N_7848,N_6975,N_7465);
xor U7849 (N_7849,N_7217,N_7467);
nand U7850 (N_7850,N_6955,N_7110);
or U7851 (N_7851,N_7198,N_7181);
nand U7852 (N_7852,N_7258,N_7229);
xnor U7853 (N_7853,N_6819,N_7428);
nand U7854 (N_7854,N_6882,N_7324);
and U7855 (N_7855,N_7055,N_7360);
nand U7856 (N_7856,N_6854,N_7137);
or U7857 (N_7857,N_7023,N_7071);
nand U7858 (N_7858,N_6867,N_7067);
or U7859 (N_7859,N_7291,N_7381);
nand U7860 (N_7860,N_7396,N_7257);
nor U7861 (N_7861,N_6776,N_7389);
nor U7862 (N_7862,N_6962,N_7358);
nand U7863 (N_7863,N_6863,N_7407);
nand U7864 (N_7864,N_7216,N_7242);
and U7865 (N_7865,N_7232,N_7286);
and U7866 (N_7866,N_7350,N_7408);
or U7867 (N_7867,N_6907,N_7274);
nor U7868 (N_7868,N_7002,N_7272);
and U7869 (N_7869,N_7091,N_6989);
or U7870 (N_7870,N_7136,N_6812);
nor U7871 (N_7871,N_7168,N_7166);
nor U7872 (N_7872,N_6864,N_6781);
or U7873 (N_7873,N_6971,N_6811);
or U7874 (N_7874,N_6969,N_7320);
or U7875 (N_7875,N_7250,N_6995);
or U7876 (N_7876,N_6909,N_7041);
and U7877 (N_7877,N_6890,N_7053);
nor U7878 (N_7878,N_7206,N_7257);
xor U7879 (N_7879,N_6828,N_7433);
nand U7880 (N_7880,N_7013,N_7235);
nor U7881 (N_7881,N_6932,N_6825);
nand U7882 (N_7882,N_6953,N_7034);
or U7883 (N_7883,N_7332,N_6757);
and U7884 (N_7884,N_7291,N_7214);
or U7885 (N_7885,N_7213,N_7098);
nor U7886 (N_7886,N_6897,N_7098);
xor U7887 (N_7887,N_7195,N_7147);
or U7888 (N_7888,N_7117,N_7413);
or U7889 (N_7889,N_7379,N_7108);
nand U7890 (N_7890,N_7298,N_7046);
and U7891 (N_7891,N_7202,N_7415);
or U7892 (N_7892,N_7251,N_7347);
nor U7893 (N_7893,N_7208,N_7285);
nor U7894 (N_7894,N_7330,N_6829);
nand U7895 (N_7895,N_7464,N_7098);
or U7896 (N_7896,N_7485,N_6916);
xnor U7897 (N_7897,N_6794,N_7379);
and U7898 (N_7898,N_6770,N_7061);
or U7899 (N_7899,N_7259,N_7315);
nor U7900 (N_7900,N_7427,N_6906);
nand U7901 (N_7901,N_7210,N_7159);
and U7902 (N_7902,N_6945,N_6999);
and U7903 (N_7903,N_6993,N_7420);
nand U7904 (N_7904,N_7452,N_7350);
nand U7905 (N_7905,N_7395,N_7462);
nand U7906 (N_7906,N_7056,N_7247);
or U7907 (N_7907,N_7340,N_7288);
nor U7908 (N_7908,N_7280,N_7216);
or U7909 (N_7909,N_7375,N_7123);
and U7910 (N_7910,N_6840,N_7477);
or U7911 (N_7911,N_6957,N_6924);
nor U7912 (N_7912,N_7095,N_6931);
nor U7913 (N_7913,N_7084,N_7211);
xor U7914 (N_7914,N_7145,N_6831);
and U7915 (N_7915,N_7140,N_6847);
or U7916 (N_7916,N_7173,N_7477);
nand U7917 (N_7917,N_7440,N_7468);
xnor U7918 (N_7918,N_7068,N_6884);
nor U7919 (N_7919,N_7342,N_6895);
and U7920 (N_7920,N_7345,N_7282);
and U7921 (N_7921,N_6922,N_7230);
xor U7922 (N_7922,N_7313,N_7283);
xor U7923 (N_7923,N_7322,N_7227);
or U7924 (N_7924,N_7122,N_7181);
nor U7925 (N_7925,N_7368,N_7260);
and U7926 (N_7926,N_7347,N_6780);
nor U7927 (N_7927,N_7255,N_7106);
nand U7928 (N_7928,N_7362,N_7023);
and U7929 (N_7929,N_7031,N_7421);
or U7930 (N_7930,N_6979,N_7034);
or U7931 (N_7931,N_7177,N_7466);
and U7932 (N_7932,N_6945,N_7406);
and U7933 (N_7933,N_7162,N_7101);
or U7934 (N_7934,N_7286,N_7411);
nor U7935 (N_7935,N_7177,N_6791);
and U7936 (N_7936,N_7022,N_7126);
nand U7937 (N_7937,N_6969,N_7238);
xnor U7938 (N_7938,N_6990,N_6873);
or U7939 (N_7939,N_7342,N_7492);
nor U7940 (N_7940,N_7479,N_7104);
nand U7941 (N_7941,N_6961,N_7081);
or U7942 (N_7942,N_7052,N_6880);
nor U7943 (N_7943,N_6815,N_6936);
nor U7944 (N_7944,N_7303,N_7469);
nand U7945 (N_7945,N_7190,N_7040);
nor U7946 (N_7946,N_7012,N_6950);
and U7947 (N_7947,N_6945,N_7368);
xnor U7948 (N_7948,N_7247,N_6834);
or U7949 (N_7949,N_7397,N_6973);
nand U7950 (N_7950,N_7271,N_7320);
nor U7951 (N_7951,N_6780,N_6830);
nor U7952 (N_7952,N_7247,N_6999);
nand U7953 (N_7953,N_7032,N_6968);
nand U7954 (N_7954,N_7246,N_7490);
and U7955 (N_7955,N_7280,N_7017);
or U7956 (N_7956,N_7006,N_6802);
xor U7957 (N_7957,N_7157,N_7014);
and U7958 (N_7958,N_7165,N_6835);
or U7959 (N_7959,N_6825,N_7290);
or U7960 (N_7960,N_7388,N_7143);
or U7961 (N_7961,N_7148,N_7419);
xor U7962 (N_7962,N_7320,N_7025);
nor U7963 (N_7963,N_7244,N_7270);
nand U7964 (N_7964,N_6866,N_7234);
nor U7965 (N_7965,N_7228,N_7413);
nor U7966 (N_7966,N_7116,N_7287);
and U7967 (N_7967,N_7195,N_7482);
or U7968 (N_7968,N_7089,N_7390);
and U7969 (N_7969,N_7033,N_6858);
nand U7970 (N_7970,N_7129,N_7085);
or U7971 (N_7971,N_7139,N_7370);
nand U7972 (N_7972,N_7365,N_7059);
xor U7973 (N_7973,N_7235,N_6792);
nor U7974 (N_7974,N_7229,N_7422);
nand U7975 (N_7975,N_7371,N_7080);
or U7976 (N_7976,N_7032,N_6840);
and U7977 (N_7977,N_6953,N_7215);
or U7978 (N_7978,N_6980,N_7210);
and U7979 (N_7979,N_6893,N_6858);
or U7980 (N_7980,N_6789,N_6847);
nand U7981 (N_7981,N_7321,N_6931);
nand U7982 (N_7982,N_7171,N_7458);
or U7983 (N_7983,N_6883,N_6875);
nand U7984 (N_7984,N_6905,N_7161);
nand U7985 (N_7985,N_7465,N_7095);
xor U7986 (N_7986,N_7434,N_6896);
or U7987 (N_7987,N_7432,N_6990);
nand U7988 (N_7988,N_7132,N_7443);
or U7989 (N_7989,N_7396,N_6834);
nand U7990 (N_7990,N_7110,N_7382);
and U7991 (N_7991,N_7421,N_6882);
xnor U7992 (N_7992,N_7031,N_6966);
xnor U7993 (N_7993,N_6930,N_6752);
and U7994 (N_7994,N_7299,N_7058);
or U7995 (N_7995,N_7188,N_7265);
and U7996 (N_7996,N_7382,N_6900);
nor U7997 (N_7997,N_7222,N_6896);
nand U7998 (N_7998,N_6942,N_7222);
or U7999 (N_7999,N_7362,N_7071);
nand U8000 (N_8000,N_7484,N_7113);
or U8001 (N_8001,N_7157,N_6934);
and U8002 (N_8002,N_7075,N_7230);
xnor U8003 (N_8003,N_6891,N_7246);
or U8004 (N_8004,N_7370,N_7250);
nand U8005 (N_8005,N_7246,N_6895);
nor U8006 (N_8006,N_7490,N_6983);
and U8007 (N_8007,N_7287,N_6822);
nand U8008 (N_8008,N_7293,N_7121);
nor U8009 (N_8009,N_7433,N_7322);
or U8010 (N_8010,N_7375,N_7043);
or U8011 (N_8011,N_7298,N_7094);
or U8012 (N_8012,N_7281,N_6794);
nor U8013 (N_8013,N_6828,N_7348);
nand U8014 (N_8014,N_6956,N_7344);
and U8015 (N_8015,N_6858,N_6978);
nand U8016 (N_8016,N_6859,N_7137);
or U8017 (N_8017,N_6810,N_7174);
or U8018 (N_8018,N_6862,N_6952);
nor U8019 (N_8019,N_7049,N_7169);
xor U8020 (N_8020,N_7460,N_7448);
nand U8021 (N_8021,N_7399,N_6981);
and U8022 (N_8022,N_6971,N_7304);
and U8023 (N_8023,N_6806,N_7419);
and U8024 (N_8024,N_6820,N_6793);
nor U8025 (N_8025,N_7151,N_6773);
nand U8026 (N_8026,N_6842,N_7188);
or U8027 (N_8027,N_6972,N_7427);
nand U8028 (N_8028,N_6767,N_7428);
or U8029 (N_8029,N_7255,N_6790);
xnor U8030 (N_8030,N_7183,N_6968);
or U8031 (N_8031,N_6987,N_6928);
nand U8032 (N_8032,N_7433,N_7021);
nand U8033 (N_8033,N_7086,N_7044);
and U8034 (N_8034,N_7326,N_6793);
nor U8035 (N_8035,N_7005,N_6931);
and U8036 (N_8036,N_7264,N_6954);
and U8037 (N_8037,N_7210,N_6933);
nand U8038 (N_8038,N_7100,N_7036);
and U8039 (N_8039,N_7204,N_6810);
and U8040 (N_8040,N_7168,N_6998);
nor U8041 (N_8041,N_7430,N_7148);
or U8042 (N_8042,N_7226,N_7348);
and U8043 (N_8043,N_7279,N_6846);
nand U8044 (N_8044,N_7452,N_7117);
nor U8045 (N_8045,N_7033,N_7037);
or U8046 (N_8046,N_7270,N_6782);
and U8047 (N_8047,N_7144,N_6774);
or U8048 (N_8048,N_7176,N_6858);
and U8049 (N_8049,N_6889,N_7125);
and U8050 (N_8050,N_7160,N_7387);
xor U8051 (N_8051,N_7281,N_6797);
nand U8052 (N_8052,N_7101,N_7183);
nand U8053 (N_8053,N_7013,N_7033);
or U8054 (N_8054,N_7123,N_7093);
xor U8055 (N_8055,N_7203,N_6827);
xnor U8056 (N_8056,N_7428,N_7014);
or U8057 (N_8057,N_7097,N_6769);
or U8058 (N_8058,N_7314,N_6975);
or U8059 (N_8059,N_7120,N_7272);
and U8060 (N_8060,N_7070,N_6809);
or U8061 (N_8061,N_7048,N_7045);
or U8062 (N_8062,N_6855,N_6882);
or U8063 (N_8063,N_7316,N_6969);
nor U8064 (N_8064,N_7195,N_7297);
and U8065 (N_8065,N_7181,N_7350);
nor U8066 (N_8066,N_7272,N_7090);
xnor U8067 (N_8067,N_7478,N_6782);
nor U8068 (N_8068,N_7248,N_7469);
and U8069 (N_8069,N_6953,N_7017);
nor U8070 (N_8070,N_7422,N_7322);
and U8071 (N_8071,N_6970,N_7369);
and U8072 (N_8072,N_6835,N_7095);
or U8073 (N_8073,N_6882,N_6921);
nand U8074 (N_8074,N_7462,N_6774);
and U8075 (N_8075,N_7229,N_7085);
and U8076 (N_8076,N_7219,N_6994);
and U8077 (N_8077,N_7348,N_7408);
xor U8078 (N_8078,N_7044,N_7468);
or U8079 (N_8079,N_7428,N_7234);
or U8080 (N_8080,N_6860,N_7356);
nor U8081 (N_8081,N_6966,N_7300);
and U8082 (N_8082,N_6842,N_6885);
nor U8083 (N_8083,N_6922,N_7241);
nand U8084 (N_8084,N_7052,N_7333);
xnor U8085 (N_8085,N_7289,N_6754);
nand U8086 (N_8086,N_6926,N_7221);
nand U8087 (N_8087,N_6831,N_6984);
or U8088 (N_8088,N_7287,N_7022);
nand U8089 (N_8089,N_7242,N_7277);
and U8090 (N_8090,N_7321,N_7329);
or U8091 (N_8091,N_6995,N_6840);
nand U8092 (N_8092,N_6834,N_7035);
nor U8093 (N_8093,N_6751,N_7143);
nand U8094 (N_8094,N_6979,N_7277);
nand U8095 (N_8095,N_7152,N_7352);
nand U8096 (N_8096,N_7373,N_7355);
nand U8097 (N_8097,N_6917,N_6987);
and U8098 (N_8098,N_7407,N_7339);
and U8099 (N_8099,N_6799,N_7077);
or U8100 (N_8100,N_7223,N_7356);
or U8101 (N_8101,N_7061,N_7056);
nor U8102 (N_8102,N_7477,N_7246);
nor U8103 (N_8103,N_6848,N_7383);
nand U8104 (N_8104,N_7499,N_6904);
nor U8105 (N_8105,N_7052,N_6993);
xor U8106 (N_8106,N_7221,N_6912);
nand U8107 (N_8107,N_7161,N_6799);
or U8108 (N_8108,N_6977,N_7142);
nand U8109 (N_8109,N_7302,N_7180);
or U8110 (N_8110,N_7118,N_7252);
nand U8111 (N_8111,N_7315,N_7470);
or U8112 (N_8112,N_7251,N_7034);
and U8113 (N_8113,N_7177,N_6957);
nand U8114 (N_8114,N_7261,N_6930);
nor U8115 (N_8115,N_7383,N_7173);
or U8116 (N_8116,N_7359,N_7158);
nor U8117 (N_8117,N_7296,N_7290);
nand U8118 (N_8118,N_7310,N_7254);
nor U8119 (N_8119,N_6880,N_6926);
and U8120 (N_8120,N_7357,N_7227);
nor U8121 (N_8121,N_6888,N_6806);
nand U8122 (N_8122,N_7160,N_7183);
xnor U8123 (N_8123,N_7289,N_6986);
and U8124 (N_8124,N_6848,N_6814);
nand U8125 (N_8125,N_7191,N_7257);
and U8126 (N_8126,N_7356,N_7083);
nor U8127 (N_8127,N_6922,N_6753);
or U8128 (N_8128,N_6997,N_7435);
or U8129 (N_8129,N_6750,N_7187);
nand U8130 (N_8130,N_7023,N_7200);
nor U8131 (N_8131,N_7089,N_7479);
or U8132 (N_8132,N_7313,N_7450);
or U8133 (N_8133,N_7234,N_7069);
nand U8134 (N_8134,N_6949,N_7326);
and U8135 (N_8135,N_6925,N_7354);
nand U8136 (N_8136,N_7356,N_7070);
nand U8137 (N_8137,N_6878,N_7146);
nor U8138 (N_8138,N_7262,N_7109);
nand U8139 (N_8139,N_6759,N_6896);
or U8140 (N_8140,N_7305,N_7144);
and U8141 (N_8141,N_7183,N_6857);
or U8142 (N_8142,N_7072,N_7094);
or U8143 (N_8143,N_7325,N_6816);
or U8144 (N_8144,N_6990,N_7207);
or U8145 (N_8145,N_7112,N_6910);
nor U8146 (N_8146,N_7271,N_7308);
and U8147 (N_8147,N_6758,N_7440);
xor U8148 (N_8148,N_7311,N_7493);
or U8149 (N_8149,N_6762,N_7171);
or U8150 (N_8150,N_7101,N_7452);
and U8151 (N_8151,N_6970,N_7493);
or U8152 (N_8152,N_7427,N_7491);
or U8153 (N_8153,N_7309,N_7244);
nand U8154 (N_8154,N_7191,N_7134);
nand U8155 (N_8155,N_7068,N_7361);
nand U8156 (N_8156,N_7003,N_7258);
or U8157 (N_8157,N_6992,N_7397);
nor U8158 (N_8158,N_7001,N_7430);
nand U8159 (N_8159,N_7014,N_7168);
and U8160 (N_8160,N_7203,N_7298);
nor U8161 (N_8161,N_6900,N_7147);
nor U8162 (N_8162,N_6865,N_7273);
and U8163 (N_8163,N_6923,N_7195);
nor U8164 (N_8164,N_7481,N_6889);
and U8165 (N_8165,N_7392,N_7162);
or U8166 (N_8166,N_7272,N_7456);
nor U8167 (N_8167,N_6805,N_7167);
nor U8168 (N_8168,N_6808,N_6816);
nand U8169 (N_8169,N_6751,N_7185);
nor U8170 (N_8170,N_6766,N_7307);
xor U8171 (N_8171,N_6823,N_6759);
nand U8172 (N_8172,N_7234,N_7052);
nor U8173 (N_8173,N_6888,N_6946);
xnor U8174 (N_8174,N_6812,N_7353);
xor U8175 (N_8175,N_7088,N_7308);
or U8176 (N_8176,N_6881,N_7224);
or U8177 (N_8177,N_7229,N_7481);
xnor U8178 (N_8178,N_6837,N_7044);
nor U8179 (N_8179,N_6943,N_7212);
or U8180 (N_8180,N_7074,N_7174);
nand U8181 (N_8181,N_6841,N_7342);
nand U8182 (N_8182,N_6819,N_7455);
nand U8183 (N_8183,N_6835,N_6984);
nor U8184 (N_8184,N_7368,N_6889);
and U8185 (N_8185,N_7311,N_7237);
or U8186 (N_8186,N_6929,N_7401);
xnor U8187 (N_8187,N_7417,N_7084);
and U8188 (N_8188,N_7222,N_6926);
or U8189 (N_8189,N_7465,N_7423);
nand U8190 (N_8190,N_6929,N_7016);
or U8191 (N_8191,N_6916,N_7256);
or U8192 (N_8192,N_7252,N_7173);
or U8193 (N_8193,N_7471,N_7389);
and U8194 (N_8194,N_7013,N_7199);
and U8195 (N_8195,N_6994,N_7231);
and U8196 (N_8196,N_7254,N_7111);
xnor U8197 (N_8197,N_7068,N_7134);
nor U8198 (N_8198,N_7479,N_7278);
nor U8199 (N_8199,N_6993,N_7154);
nor U8200 (N_8200,N_7344,N_6874);
nand U8201 (N_8201,N_6843,N_7433);
and U8202 (N_8202,N_7240,N_7268);
and U8203 (N_8203,N_6838,N_7443);
and U8204 (N_8204,N_7408,N_7115);
nor U8205 (N_8205,N_7205,N_7167);
or U8206 (N_8206,N_6985,N_7129);
or U8207 (N_8207,N_7222,N_7075);
nor U8208 (N_8208,N_6984,N_6897);
or U8209 (N_8209,N_6958,N_7362);
nand U8210 (N_8210,N_7323,N_7359);
nor U8211 (N_8211,N_7084,N_7243);
or U8212 (N_8212,N_7214,N_7422);
and U8213 (N_8213,N_6795,N_7100);
or U8214 (N_8214,N_7268,N_7113);
nand U8215 (N_8215,N_7029,N_7125);
nand U8216 (N_8216,N_7271,N_6964);
and U8217 (N_8217,N_7072,N_7389);
and U8218 (N_8218,N_7248,N_6842);
nor U8219 (N_8219,N_7147,N_6792);
and U8220 (N_8220,N_7000,N_7076);
or U8221 (N_8221,N_7133,N_6891);
nor U8222 (N_8222,N_6971,N_7491);
nor U8223 (N_8223,N_7309,N_7363);
xor U8224 (N_8224,N_7387,N_6755);
xnor U8225 (N_8225,N_6893,N_6807);
or U8226 (N_8226,N_7445,N_7373);
nor U8227 (N_8227,N_7395,N_7293);
nor U8228 (N_8228,N_6954,N_7418);
or U8229 (N_8229,N_6771,N_7327);
nor U8230 (N_8230,N_7265,N_6934);
nor U8231 (N_8231,N_6873,N_7174);
xnor U8232 (N_8232,N_7433,N_7047);
or U8233 (N_8233,N_7196,N_6903);
or U8234 (N_8234,N_7277,N_7099);
or U8235 (N_8235,N_7083,N_7138);
and U8236 (N_8236,N_7351,N_7219);
or U8237 (N_8237,N_6894,N_7177);
nand U8238 (N_8238,N_7091,N_7011);
nor U8239 (N_8239,N_7313,N_7361);
nor U8240 (N_8240,N_7414,N_6875);
and U8241 (N_8241,N_6912,N_7280);
nor U8242 (N_8242,N_7333,N_6755);
nand U8243 (N_8243,N_6863,N_6950);
and U8244 (N_8244,N_7251,N_6880);
nand U8245 (N_8245,N_6795,N_7031);
and U8246 (N_8246,N_7229,N_6910);
and U8247 (N_8247,N_7171,N_6790);
xnor U8248 (N_8248,N_7462,N_6980);
nand U8249 (N_8249,N_6859,N_6988);
or U8250 (N_8250,N_7989,N_7976);
nor U8251 (N_8251,N_7723,N_8167);
or U8252 (N_8252,N_7858,N_8216);
or U8253 (N_8253,N_7582,N_8146);
and U8254 (N_8254,N_7519,N_7835);
nand U8255 (N_8255,N_8032,N_7837);
and U8256 (N_8256,N_7521,N_7774);
and U8257 (N_8257,N_7939,N_7893);
nand U8258 (N_8258,N_7662,N_8188);
nand U8259 (N_8259,N_8190,N_7897);
and U8260 (N_8260,N_7794,N_7879);
xor U8261 (N_8261,N_7504,N_7623);
and U8262 (N_8262,N_7556,N_7742);
nor U8263 (N_8263,N_8244,N_7969);
nand U8264 (N_8264,N_7531,N_8053);
and U8265 (N_8265,N_7945,N_7666);
nand U8266 (N_8266,N_7627,N_7926);
and U8267 (N_8267,N_7831,N_7741);
nand U8268 (N_8268,N_8033,N_8018);
xnor U8269 (N_8269,N_7753,N_7875);
xor U8270 (N_8270,N_7889,N_8173);
or U8271 (N_8271,N_8208,N_7910);
nand U8272 (N_8272,N_7944,N_7718);
and U8273 (N_8273,N_7609,N_8223);
and U8274 (N_8274,N_8103,N_7980);
nand U8275 (N_8275,N_8236,N_7721);
xnor U8276 (N_8276,N_7796,N_8095);
nand U8277 (N_8277,N_7909,N_8054);
nand U8278 (N_8278,N_8084,N_8028);
or U8279 (N_8279,N_7901,N_7757);
nor U8280 (N_8280,N_7560,N_7524);
nor U8281 (N_8281,N_7847,N_8149);
xnor U8282 (N_8282,N_7870,N_7682);
nor U8283 (N_8283,N_7615,N_7553);
or U8284 (N_8284,N_8125,N_8038);
and U8285 (N_8285,N_8011,N_7888);
and U8286 (N_8286,N_7848,N_7839);
xnor U8287 (N_8287,N_8090,N_8221);
nor U8288 (N_8288,N_7624,N_7932);
nor U8289 (N_8289,N_7728,N_7523);
and U8290 (N_8290,N_8062,N_7978);
nor U8291 (N_8291,N_8227,N_8243);
or U8292 (N_8292,N_7746,N_7731);
nor U8293 (N_8293,N_7604,N_7584);
nand U8294 (N_8294,N_7622,N_7898);
and U8295 (N_8295,N_7878,N_7800);
nand U8296 (N_8296,N_8220,N_8222);
nor U8297 (N_8297,N_7679,N_8120);
or U8298 (N_8298,N_7549,N_7915);
nor U8299 (N_8299,N_8166,N_7594);
or U8300 (N_8300,N_7561,N_8073);
or U8301 (N_8301,N_8114,N_7791);
or U8302 (N_8302,N_8080,N_7613);
nand U8303 (N_8303,N_7507,N_8193);
and U8304 (N_8304,N_7591,N_7992);
and U8305 (N_8305,N_7924,N_7844);
or U8306 (N_8306,N_8217,N_7743);
nand U8307 (N_8307,N_7670,N_7798);
and U8308 (N_8308,N_8031,N_8007);
nand U8309 (N_8309,N_8214,N_7687);
nand U8310 (N_8310,N_7656,N_7784);
or U8311 (N_8311,N_7542,N_7955);
nor U8312 (N_8312,N_8002,N_7936);
or U8313 (N_8313,N_8218,N_8237);
xnor U8314 (N_8314,N_7612,N_7614);
or U8315 (N_8315,N_8112,N_7678);
xor U8316 (N_8316,N_7639,N_7942);
or U8317 (N_8317,N_7845,N_7628);
and U8318 (N_8318,N_7533,N_7994);
or U8319 (N_8319,N_7676,N_7896);
nor U8320 (N_8320,N_7812,N_7651);
or U8321 (N_8321,N_8065,N_8207);
nor U8322 (N_8322,N_7587,N_8170);
nor U8323 (N_8323,N_7877,N_7669);
or U8324 (N_8324,N_7506,N_7933);
nand U8325 (N_8325,N_7593,N_7778);
and U8326 (N_8326,N_8093,N_8088);
nor U8327 (N_8327,N_7668,N_7551);
nor U8328 (N_8328,N_7857,N_7706);
and U8329 (N_8329,N_7620,N_7738);
and U8330 (N_8330,N_8196,N_7546);
nor U8331 (N_8331,N_7547,N_8025);
and U8332 (N_8332,N_7704,N_8091);
and U8333 (N_8333,N_8159,N_7868);
nor U8334 (N_8334,N_7640,N_7647);
nor U8335 (N_8335,N_8119,N_7807);
or U8336 (N_8336,N_7780,N_7540);
nand U8337 (N_8337,N_7577,N_7502);
xnor U8338 (N_8338,N_7766,N_7811);
nand U8339 (N_8339,N_7658,N_7759);
nor U8340 (N_8340,N_7641,N_7708);
nor U8341 (N_8341,N_8104,N_7683);
nor U8342 (N_8342,N_8132,N_7971);
xor U8343 (N_8343,N_7694,N_7650);
and U8344 (N_8344,N_7618,N_7821);
or U8345 (N_8345,N_7816,N_7948);
or U8346 (N_8346,N_8141,N_8009);
nor U8347 (N_8347,N_8010,N_8013);
and U8348 (N_8348,N_7884,N_8020);
nand U8349 (N_8349,N_7664,N_7636);
and U8350 (N_8350,N_7792,N_7714);
and U8351 (N_8351,N_8206,N_7903);
and U8352 (N_8352,N_8179,N_7581);
nor U8353 (N_8353,N_7552,N_7625);
or U8354 (N_8354,N_7712,N_7733);
or U8355 (N_8355,N_7817,N_7815);
nor U8356 (N_8356,N_7566,N_7779);
nor U8357 (N_8357,N_8061,N_7619);
nor U8358 (N_8358,N_8136,N_8246);
or U8359 (N_8359,N_7867,N_8134);
nor U8360 (N_8360,N_7536,N_7520);
or U8361 (N_8361,N_7674,N_7751);
and U8362 (N_8362,N_8044,N_8154);
and U8363 (N_8363,N_7554,N_8239);
nand U8364 (N_8364,N_8029,N_8004);
nand U8365 (N_8365,N_7840,N_8245);
nor U8366 (N_8366,N_7834,N_7979);
nor U8367 (N_8367,N_8015,N_8139);
and U8368 (N_8368,N_8169,N_8022);
and U8369 (N_8369,N_8107,N_7735);
nor U8370 (N_8370,N_7538,N_8242);
nor U8371 (N_8371,N_7974,N_7863);
nand U8372 (N_8372,N_8128,N_7541);
nor U8373 (N_8373,N_8185,N_7701);
or U8374 (N_8374,N_7770,N_8005);
nor U8375 (N_8375,N_7637,N_7958);
nor U8376 (N_8376,N_7904,N_8201);
nand U8377 (N_8377,N_7927,N_8186);
and U8378 (N_8378,N_8086,N_7528);
nor U8379 (N_8379,N_7667,N_8123);
and U8380 (N_8380,N_7599,N_7886);
or U8381 (N_8381,N_7890,N_8016);
nand U8382 (N_8382,N_7539,N_7852);
or U8383 (N_8383,N_7607,N_8209);
or U8384 (N_8384,N_8041,N_7929);
or U8385 (N_8385,N_7930,N_7999);
nand U8386 (N_8386,N_8161,N_7765);
nand U8387 (N_8387,N_8059,N_7805);
and U8388 (N_8388,N_8226,N_7653);
and U8389 (N_8389,N_8232,N_7987);
xor U8390 (N_8390,N_8233,N_8230);
nor U8391 (N_8391,N_7588,N_7657);
or U8392 (N_8392,N_7940,N_7854);
nand U8393 (N_8393,N_7754,N_7700);
and U8394 (N_8394,N_7596,N_7876);
nand U8395 (N_8395,N_7830,N_7899);
nand U8396 (N_8396,N_8130,N_7855);
and U8397 (N_8397,N_8017,N_7570);
or U8398 (N_8398,N_7710,N_8126);
or U8399 (N_8399,N_7516,N_8249);
or U8400 (N_8400,N_8203,N_8105);
or U8401 (N_8401,N_8213,N_7938);
xor U8402 (N_8402,N_8064,N_8021);
and U8403 (N_8403,N_8072,N_7672);
nand U8404 (N_8404,N_7906,N_7829);
nand U8405 (N_8405,N_8116,N_7725);
and U8406 (N_8406,N_7762,N_8008);
and U8407 (N_8407,N_7768,N_7913);
and U8408 (N_8408,N_7995,N_7510);
xor U8409 (N_8409,N_7822,N_7900);
and U8410 (N_8410,N_7874,N_7610);
or U8411 (N_8411,N_7922,N_7871);
and U8412 (N_8412,N_7761,N_8058);
or U8413 (N_8413,N_7564,N_7842);
xnor U8414 (N_8414,N_7902,N_7732);
or U8415 (N_8415,N_8162,N_7727);
nand U8416 (N_8416,N_7786,N_8122);
or U8417 (N_8417,N_7959,N_7826);
or U8418 (N_8418,N_7632,N_8078);
or U8419 (N_8419,N_8199,N_7764);
and U8420 (N_8420,N_7745,N_7730);
nor U8421 (N_8421,N_8121,N_7684);
or U8422 (N_8422,N_7951,N_8197);
nor U8423 (N_8423,N_7887,N_7962);
and U8424 (N_8424,N_7643,N_7644);
or U8425 (N_8425,N_7843,N_7841);
or U8426 (N_8426,N_7782,N_8047);
and U8427 (N_8427,N_7716,N_7724);
nor U8428 (N_8428,N_7983,N_8133);
nor U8429 (N_8429,N_7693,N_7908);
or U8430 (N_8430,N_7646,N_7680);
and U8431 (N_8431,N_7565,N_8049);
nor U8432 (N_8432,N_8202,N_7977);
or U8433 (N_8433,N_7824,N_8063);
nor U8434 (N_8434,N_7905,N_8048);
nand U8435 (N_8435,N_7760,N_7861);
and U8436 (N_8436,N_7853,N_7990);
nand U8437 (N_8437,N_8195,N_7525);
nor U8438 (N_8438,N_8157,N_8148);
and U8439 (N_8439,N_7634,N_8229);
nor U8440 (N_8440,N_7655,N_7814);
nor U8441 (N_8441,N_7513,N_8165);
nand U8442 (N_8442,N_7544,N_7691);
and U8443 (N_8443,N_7997,N_8037);
xnor U8444 (N_8444,N_7616,N_7773);
or U8445 (N_8445,N_8211,N_7788);
xnor U8446 (N_8446,N_7921,N_7946);
nand U8447 (N_8447,N_7602,N_8164);
or U8448 (N_8448,N_8156,N_7801);
or U8449 (N_8449,N_7937,N_7785);
or U8450 (N_8450,N_7850,N_7752);
nand U8451 (N_8451,N_8057,N_7715);
nor U8452 (N_8452,N_7920,N_7749);
or U8453 (N_8453,N_7720,N_7763);
nor U8454 (N_8454,N_8142,N_8176);
nand U8455 (N_8455,N_7550,N_8231);
xnor U8456 (N_8456,N_7512,N_7856);
and U8457 (N_8457,N_8068,N_7597);
nand U8458 (N_8458,N_7568,N_7777);
or U8459 (N_8459,N_7892,N_7827);
nand U8460 (N_8460,N_7663,N_8163);
nor U8461 (N_8461,N_7864,N_8098);
and U8462 (N_8462,N_7836,N_8234);
nor U8463 (N_8463,N_7648,N_7916);
or U8464 (N_8464,N_7756,N_7608);
xor U8465 (N_8465,N_8094,N_7739);
or U8466 (N_8466,N_8085,N_7500);
nor U8467 (N_8467,N_7558,N_8192);
or U8468 (N_8468,N_7660,N_7880);
or U8469 (N_8469,N_8129,N_8099);
nor U8470 (N_8470,N_7820,N_7505);
and U8471 (N_8471,N_7789,N_7517);
nand U8472 (N_8472,N_7895,N_7804);
nand U8473 (N_8473,N_7567,N_7705);
xnor U8474 (N_8474,N_7803,N_8155);
nor U8475 (N_8475,N_8212,N_8117);
nor U8476 (N_8476,N_8240,N_7661);
nor U8477 (N_8477,N_7818,N_7917);
nand U8478 (N_8478,N_7767,N_7569);
or U8479 (N_8479,N_7862,N_7967);
or U8480 (N_8480,N_7960,N_8238);
and U8481 (N_8481,N_7873,N_8039);
nand U8482 (N_8482,N_7849,N_8069);
xor U8483 (N_8483,N_7793,N_7585);
xnor U8484 (N_8484,N_7589,N_7645);
or U8485 (N_8485,N_8168,N_7988);
and U8486 (N_8486,N_8060,N_7649);
nor U8487 (N_8487,N_8110,N_8082);
and U8488 (N_8488,N_8014,N_7966);
xnor U8489 (N_8489,N_8182,N_8200);
nand U8490 (N_8490,N_8131,N_7996);
nor U8491 (N_8491,N_8067,N_7697);
and U8492 (N_8492,N_8180,N_8111);
xor U8493 (N_8493,N_7686,N_8036);
nor U8494 (N_8494,N_7642,N_8046);
or U8495 (N_8495,N_7695,N_8106);
nand U8496 (N_8496,N_7809,N_8172);
nor U8497 (N_8497,N_7882,N_7522);
or U8498 (N_8498,N_8205,N_8089);
nor U8499 (N_8499,N_7630,N_7529);
and U8500 (N_8500,N_8143,N_8215);
nor U8501 (N_8501,N_7734,N_7957);
nand U8502 (N_8502,N_8144,N_8006);
and U8503 (N_8503,N_7621,N_8204);
and U8504 (N_8504,N_7729,N_8151);
or U8505 (N_8505,N_7514,N_8152);
xnor U8506 (N_8506,N_7703,N_7783);
or U8507 (N_8507,N_8135,N_7709);
nor U8508 (N_8508,N_7776,N_7947);
nor U8509 (N_8509,N_7772,N_7696);
nor U8510 (N_8510,N_7555,N_7881);
nor U8511 (N_8511,N_7583,N_8079);
nor U8512 (N_8512,N_7769,N_7677);
nor U8513 (N_8513,N_7563,N_7671);
nor U8514 (N_8514,N_7534,N_7956);
xnor U8515 (N_8515,N_7673,N_7787);
and U8516 (N_8516,N_8118,N_7952);
nor U8517 (N_8517,N_7869,N_7737);
xnor U8518 (N_8518,N_7846,N_7802);
and U8519 (N_8519,N_7865,N_7699);
nor U8520 (N_8520,N_7690,N_8224);
nor U8521 (N_8521,N_7931,N_7559);
nand U8522 (N_8522,N_8070,N_7573);
xor U8523 (N_8523,N_8075,N_7574);
xor U8524 (N_8524,N_8153,N_8100);
or U8525 (N_8525,N_7717,N_7685);
and U8526 (N_8526,N_8050,N_7629);
nand U8527 (N_8527,N_7736,N_7747);
nand U8528 (N_8528,N_8074,N_7631);
and U8529 (N_8529,N_7823,N_7617);
nand U8530 (N_8530,N_7813,N_7681);
or U8531 (N_8531,N_8184,N_8087);
or U8532 (N_8532,N_8235,N_8071);
or U8533 (N_8533,N_7509,N_8027);
nand U8534 (N_8534,N_7975,N_8191);
nand U8535 (N_8535,N_7659,N_7635);
nand U8536 (N_8536,N_8171,N_8035);
nand U8537 (N_8537,N_7605,N_7557);
and U8538 (N_8538,N_7543,N_7527);
nand U8539 (N_8539,N_7771,N_7711);
and U8540 (N_8540,N_8019,N_7968);
nand U8541 (N_8541,N_8109,N_7744);
xor U8542 (N_8542,N_7508,N_7526);
nand U8543 (N_8543,N_7511,N_7501);
and U8544 (N_8544,N_7885,N_7982);
or U8545 (N_8545,N_8127,N_7919);
or U8546 (N_8546,N_7503,N_7950);
xnor U8547 (N_8547,N_7790,N_7740);
nand U8548 (N_8548,N_7590,N_7925);
or U8549 (N_8549,N_7912,N_8030);
or U8550 (N_8550,N_7949,N_8001);
or U8551 (N_8551,N_7665,N_7964);
nor U8552 (N_8552,N_8081,N_8024);
nor U8553 (N_8553,N_7859,N_7981);
and U8554 (N_8554,N_7838,N_7586);
or U8555 (N_8555,N_7943,N_7985);
nor U8556 (N_8556,N_7575,N_8056);
and U8557 (N_8557,N_7675,N_8138);
nand U8558 (N_8558,N_8034,N_7580);
and U8559 (N_8559,N_7935,N_7928);
xnor U8560 (N_8560,N_7810,N_7578);
nand U8561 (N_8561,N_7598,N_8042);
and U8562 (N_8562,N_7883,N_8175);
and U8563 (N_8563,N_7518,N_8219);
nor U8564 (N_8564,N_7941,N_7689);
or U8565 (N_8565,N_7611,N_7973);
nor U8566 (N_8566,N_7965,N_8210);
nor U8567 (N_8567,N_7515,N_8096);
and U8568 (N_8568,N_7722,N_7595);
nand U8569 (N_8569,N_7998,N_7750);
nand U8570 (N_8570,N_7972,N_7633);
and U8571 (N_8571,N_7963,N_7984);
and U8572 (N_8572,N_7808,N_7532);
nand U8573 (N_8573,N_7799,N_7698);
nor U8574 (N_8574,N_7548,N_7991);
or U8575 (N_8575,N_7851,N_7833);
or U8576 (N_8576,N_8177,N_7872);
or U8577 (N_8577,N_7970,N_7719);
or U8578 (N_8578,N_8178,N_8248);
nand U8579 (N_8579,N_7781,N_7832);
nor U8580 (N_8580,N_7923,N_7545);
nor U8581 (N_8581,N_7571,N_7535);
nand U8582 (N_8582,N_8183,N_7713);
nand U8583 (N_8583,N_7592,N_8101);
nand U8584 (N_8584,N_7726,N_8076);
or U8585 (N_8585,N_7866,N_7688);
and U8586 (N_8586,N_7828,N_8187);
or U8587 (N_8587,N_7748,N_7626);
nand U8588 (N_8588,N_8115,N_8140);
xor U8589 (N_8589,N_8097,N_7579);
and U8590 (N_8590,N_8012,N_7600);
nor U8591 (N_8591,N_7961,N_7652);
nor U8592 (N_8592,N_7954,N_7537);
nand U8593 (N_8593,N_8066,N_8225);
xnor U8594 (N_8594,N_8003,N_8194);
nor U8595 (N_8595,N_8241,N_8000);
nand U8596 (N_8596,N_7993,N_8045);
and U8597 (N_8597,N_7572,N_7797);
nor U8598 (N_8598,N_7825,N_7806);
xor U8599 (N_8599,N_7638,N_7911);
xnor U8600 (N_8600,N_7654,N_8158);
xor U8601 (N_8601,N_8051,N_7562);
or U8602 (N_8602,N_8147,N_7986);
nand U8603 (N_8603,N_8092,N_8181);
or U8604 (N_8604,N_8102,N_7758);
and U8605 (N_8605,N_7755,N_7918);
or U8606 (N_8606,N_7775,N_7953);
or U8607 (N_8607,N_7934,N_8124);
and U8608 (N_8608,N_8052,N_7907);
or U8609 (N_8609,N_7692,N_8228);
nand U8610 (N_8610,N_8113,N_7860);
nor U8611 (N_8611,N_8137,N_7707);
or U8612 (N_8612,N_8108,N_8189);
nor U8613 (N_8613,N_8160,N_7702);
or U8614 (N_8614,N_8055,N_8247);
nor U8615 (N_8615,N_8023,N_8043);
and U8616 (N_8616,N_7601,N_8026);
xor U8617 (N_8617,N_8150,N_8040);
and U8618 (N_8618,N_7819,N_8145);
and U8619 (N_8619,N_7795,N_7914);
nor U8620 (N_8620,N_7606,N_7530);
nand U8621 (N_8621,N_7576,N_7894);
or U8622 (N_8622,N_8198,N_7891);
nand U8623 (N_8623,N_8083,N_8077);
nor U8624 (N_8624,N_8174,N_7603);
or U8625 (N_8625,N_8075,N_8080);
nand U8626 (N_8626,N_7962,N_7668);
nor U8627 (N_8627,N_8124,N_8106);
or U8628 (N_8628,N_8187,N_7846);
or U8629 (N_8629,N_8209,N_8208);
and U8630 (N_8630,N_8167,N_8207);
and U8631 (N_8631,N_8216,N_8198);
xnor U8632 (N_8632,N_8042,N_7827);
xor U8633 (N_8633,N_8199,N_8077);
nand U8634 (N_8634,N_7987,N_7691);
nand U8635 (N_8635,N_8112,N_7970);
nand U8636 (N_8636,N_7878,N_7683);
or U8637 (N_8637,N_7926,N_7894);
xnor U8638 (N_8638,N_7625,N_8151);
xnor U8639 (N_8639,N_8123,N_7686);
xor U8640 (N_8640,N_7818,N_7890);
and U8641 (N_8641,N_7647,N_8197);
xnor U8642 (N_8642,N_7832,N_7661);
nand U8643 (N_8643,N_7766,N_7694);
nand U8644 (N_8644,N_7825,N_7888);
nor U8645 (N_8645,N_7677,N_7921);
nand U8646 (N_8646,N_7508,N_8231);
nor U8647 (N_8647,N_7989,N_7621);
nor U8648 (N_8648,N_7902,N_8048);
nor U8649 (N_8649,N_7693,N_7656);
xnor U8650 (N_8650,N_7659,N_8019);
nor U8651 (N_8651,N_8025,N_7947);
or U8652 (N_8652,N_7814,N_8093);
nand U8653 (N_8653,N_7727,N_7783);
nand U8654 (N_8654,N_7819,N_7666);
nand U8655 (N_8655,N_7653,N_7544);
xnor U8656 (N_8656,N_7676,N_7679);
or U8657 (N_8657,N_8017,N_7800);
xor U8658 (N_8658,N_7676,N_7840);
nor U8659 (N_8659,N_8229,N_7720);
nand U8660 (N_8660,N_7550,N_8072);
nor U8661 (N_8661,N_8038,N_7856);
nor U8662 (N_8662,N_8241,N_7827);
nand U8663 (N_8663,N_8219,N_7684);
nand U8664 (N_8664,N_7895,N_8190);
nor U8665 (N_8665,N_7686,N_7655);
and U8666 (N_8666,N_7793,N_7712);
nor U8667 (N_8667,N_7885,N_7758);
or U8668 (N_8668,N_7820,N_8199);
xor U8669 (N_8669,N_7964,N_8044);
and U8670 (N_8670,N_7529,N_7746);
nand U8671 (N_8671,N_7664,N_7771);
and U8672 (N_8672,N_8137,N_7916);
nand U8673 (N_8673,N_7551,N_7737);
nand U8674 (N_8674,N_7717,N_7810);
and U8675 (N_8675,N_7940,N_8184);
nor U8676 (N_8676,N_7768,N_8148);
nor U8677 (N_8677,N_7546,N_8120);
or U8678 (N_8678,N_8187,N_7682);
and U8679 (N_8679,N_8010,N_7818);
nor U8680 (N_8680,N_7649,N_8185);
nor U8681 (N_8681,N_8173,N_7991);
and U8682 (N_8682,N_8139,N_8171);
xor U8683 (N_8683,N_7645,N_7717);
nor U8684 (N_8684,N_8042,N_8201);
nand U8685 (N_8685,N_7591,N_7764);
and U8686 (N_8686,N_7537,N_7561);
nor U8687 (N_8687,N_7955,N_7659);
nor U8688 (N_8688,N_8182,N_7518);
nor U8689 (N_8689,N_7895,N_7812);
nand U8690 (N_8690,N_7910,N_8050);
nand U8691 (N_8691,N_7849,N_7717);
or U8692 (N_8692,N_8023,N_8161);
nor U8693 (N_8693,N_8214,N_7847);
or U8694 (N_8694,N_7600,N_8202);
and U8695 (N_8695,N_7671,N_7979);
and U8696 (N_8696,N_8093,N_8060);
nor U8697 (N_8697,N_7911,N_8159);
nand U8698 (N_8698,N_8205,N_8016);
or U8699 (N_8699,N_7998,N_7717);
and U8700 (N_8700,N_8112,N_8190);
nor U8701 (N_8701,N_7874,N_8229);
or U8702 (N_8702,N_7718,N_7516);
and U8703 (N_8703,N_7529,N_8238);
nor U8704 (N_8704,N_7697,N_7878);
or U8705 (N_8705,N_7544,N_7561);
nor U8706 (N_8706,N_7670,N_7682);
nor U8707 (N_8707,N_7838,N_7638);
nand U8708 (N_8708,N_7998,N_8008);
or U8709 (N_8709,N_8222,N_7504);
xnor U8710 (N_8710,N_7879,N_7771);
xor U8711 (N_8711,N_8211,N_8065);
nand U8712 (N_8712,N_7809,N_8058);
and U8713 (N_8713,N_7559,N_7712);
nor U8714 (N_8714,N_7678,N_8188);
nand U8715 (N_8715,N_7815,N_7973);
nand U8716 (N_8716,N_7824,N_7608);
and U8717 (N_8717,N_8182,N_7520);
xnor U8718 (N_8718,N_7528,N_8207);
and U8719 (N_8719,N_8031,N_7757);
and U8720 (N_8720,N_7650,N_7568);
and U8721 (N_8721,N_7938,N_7799);
and U8722 (N_8722,N_7888,N_7620);
or U8723 (N_8723,N_8237,N_8124);
or U8724 (N_8724,N_7714,N_7772);
nand U8725 (N_8725,N_8131,N_8143);
and U8726 (N_8726,N_7988,N_7569);
and U8727 (N_8727,N_7808,N_8004);
nor U8728 (N_8728,N_8055,N_8079);
nand U8729 (N_8729,N_7690,N_7763);
or U8730 (N_8730,N_7594,N_7655);
xnor U8731 (N_8731,N_7687,N_8025);
nor U8732 (N_8732,N_7796,N_7518);
nand U8733 (N_8733,N_8214,N_7871);
and U8734 (N_8734,N_7931,N_8036);
and U8735 (N_8735,N_7889,N_7686);
nand U8736 (N_8736,N_7932,N_7873);
nor U8737 (N_8737,N_7597,N_8014);
and U8738 (N_8738,N_8015,N_7906);
or U8739 (N_8739,N_8021,N_8015);
nand U8740 (N_8740,N_7724,N_7886);
nor U8741 (N_8741,N_7724,N_7961);
xor U8742 (N_8742,N_8003,N_7603);
nor U8743 (N_8743,N_7626,N_7541);
xnor U8744 (N_8744,N_7575,N_7876);
or U8745 (N_8745,N_7836,N_7788);
and U8746 (N_8746,N_7607,N_7836);
nand U8747 (N_8747,N_7540,N_8031);
nor U8748 (N_8748,N_7944,N_7634);
xnor U8749 (N_8749,N_7819,N_8163);
and U8750 (N_8750,N_7987,N_7939);
nand U8751 (N_8751,N_7796,N_7887);
nor U8752 (N_8752,N_8249,N_7600);
nand U8753 (N_8753,N_7523,N_8043);
nor U8754 (N_8754,N_8035,N_8111);
or U8755 (N_8755,N_7758,N_7509);
or U8756 (N_8756,N_7967,N_7813);
nor U8757 (N_8757,N_7996,N_7972);
nor U8758 (N_8758,N_8110,N_7838);
nand U8759 (N_8759,N_7802,N_7728);
and U8760 (N_8760,N_7859,N_8008);
xor U8761 (N_8761,N_7687,N_8183);
or U8762 (N_8762,N_8030,N_7689);
or U8763 (N_8763,N_8126,N_7533);
and U8764 (N_8764,N_7599,N_7950);
xor U8765 (N_8765,N_7874,N_7617);
or U8766 (N_8766,N_7844,N_7974);
and U8767 (N_8767,N_7541,N_7832);
or U8768 (N_8768,N_8247,N_8097);
nand U8769 (N_8769,N_7587,N_8242);
nand U8770 (N_8770,N_8101,N_8150);
nand U8771 (N_8771,N_7729,N_8145);
xor U8772 (N_8772,N_7704,N_7640);
nand U8773 (N_8773,N_7877,N_7918);
nand U8774 (N_8774,N_7556,N_8118);
xor U8775 (N_8775,N_7984,N_7935);
or U8776 (N_8776,N_7740,N_7565);
or U8777 (N_8777,N_7889,N_7986);
xor U8778 (N_8778,N_7782,N_7564);
or U8779 (N_8779,N_7755,N_7963);
and U8780 (N_8780,N_8154,N_7766);
xor U8781 (N_8781,N_7571,N_7527);
nand U8782 (N_8782,N_7640,N_7917);
nor U8783 (N_8783,N_7508,N_7922);
or U8784 (N_8784,N_7607,N_7955);
nand U8785 (N_8785,N_7982,N_8189);
and U8786 (N_8786,N_8134,N_8083);
or U8787 (N_8787,N_7721,N_8043);
nor U8788 (N_8788,N_8243,N_7904);
or U8789 (N_8789,N_7967,N_7972);
and U8790 (N_8790,N_7706,N_7895);
and U8791 (N_8791,N_7692,N_8243);
and U8792 (N_8792,N_8105,N_8108);
nor U8793 (N_8793,N_7929,N_7648);
or U8794 (N_8794,N_7713,N_8130);
or U8795 (N_8795,N_7691,N_8050);
and U8796 (N_8796,N_7863,N_7777);
or U8797 (N_8797,N_7823,N_7549);
xor U8798 (N_8798,N_7600,N_7854);
nand U8799 (N_8799,N_7754,N_8199);
nand U8800 (N_8800,N_8092,N_8073);
nand U8801 (N_8801,N_7876,N_7817);
nor U8802 (N_8802,N_8033,N_7802);
or U8803 (N_8803,N_7864,N_7983);
nand U8804 (N_8804,N_7517,N_7614);
nand U8805 (N_8805,N_8184,N_7917);
or U8806 (N_8806,N_8240,N_8090);
xor U8807 (N_8807,N_8042,N_8143);
nand U8808 (N_8808,N_7707,N_7622);
xor U8809 (N_8809,N_8076,N_7619);
and U8810 (N_8810,N_8092,N_7822);
nor U8811 (N_8811,N_7714,N_7851);
and U8812 (N_8812,N_7683,N_8142);
nand U8813 (N_8813,N_7975,N_8052);
and U8814 (N_8814,N_7701,N_7587);
and U8815 (N_8815,N_7783,N_7829);
nand U8816 (N_8816,N_8002,N_8210);
nor U8817 (N_8817,N_7662,N_7881);
and U8818 (N_8818,N_7768,N_8119);
nor U8819 (N_8819,N_7598,N_7972);
nor U8820 (N_8820,N_7769,N_7796);
and U8821 (N_8821,N_8204,N_7833);
or U8822 (N_8822,N_7978,N_8017);
nor U8823 (N_8823,N_7716,N_8124);
nor U8824 (N_8824,N_7838,N_7860);
nand U8825 (N_8825,N_7970,N_7853);
nor U8826 (N_8826,N_7927,N_7982);
or U8827 (N_8827,N_8161,N_7760);
and U8828 (N_8828,N_7583,N_7837);
or U8829 (N_8829,N_7896,N_7673);
nor U8830 (N_8830,N_7731,N_8018);
nor U8831 (N_8831,N_7916,N_7816);
or U8832 (N_8832,N_7756,N_8005);
or U8833 (N_8833,N_7703,N_7720);
or U8834 (N_8834,N_7749,N_7959);
and U8835 (N_8835,N_7619,N_7890);
nor U8836 (N_8836,N_8211,N_7796);
nand U8837 (N_8837,N_7798,N_7611);
xnor U8838 (N_8838,N_7992,N_7610);
nor U8839 (N_8839,N_7594,N_8145);
and U8840 (N_8840,N_7545,N_8144);
or U8841 (N_8841,N_8232,N_7598);
nor U8842 (N_8842,N_7859,N_8202);
xor U8843 (N_8843,N_7554,N_7552);
nor U8844 (N_8844,N_7727,N_7860);
or U8845 (N_8845,N_8037,N_8128);
nand U8846 (N_8846,N_7538,N_8162);
or U8847 (N_8847,N_7902,N_7953);
or U8848 (N_8848,N_7623,N_7518);
nor U8849 (N_8849,N_8008,N_7633);
nand U8850 (N_8850,N_7985,N_7899);
xnor U8851 (N_8851,N_8094,N_7818);
xor U8852 (N_8852,N_7592,N_7826);
xnor U8853 (N_8853,N_7602,N_7750);
or U8854 (N_8854,N_8243,N_8142);
nand U8855 (N_8855,N_7768,N_7546);
nand U8856 (N_8856,N_7725,N_7789);
xor U8857 (N_8857,N_7517,N_8047);
or U8858 (N_8858,N_8007,N_7764);
and U8859 (N_8859,N_7704,N_7618);
nand U8860 (N_8860,N_8081,N_7764);
and U8861 (N_8861,N_7593,N_8237);
nand U8862 (N_8862,N_7962,N_7598);
and U8863 (N_8863,N_7992,N_8028);
and U8864 (N_8864,N_7548,N_7648);
nor U8865 (N_8865,N_7581,N_8098);
nor U8866 (N_8866,N_7911,N_7707);
or U8867 (N_8867,N_7656,N_7646);
nand U8868 (N_8868,N_8119,N_8043);
and U8869 (N_8869,N_8125,N_7594);
nor U8870 (N_8870,N_8166,N_7979);
nand U8871 (N_8871,N_8062,N_8132);
nor U8872 (N_8872,N_7907,N_7701);
or U8873 (N_8873,N_8071,N_8249);
and U8874 (N_8874,N_8219,N_7574);
or U8875 (N_8875,N_7546,N_8186);
xor U8876 (N_8876,N_8044,N_7803);
nor U8877 (N_8877,N_8049,N_7705);
and U8878 (N_8878,N_7658,N_7775);
nand U8879 (N_8879,N_7758,N_7809);
xnor U8880 (N_8880,N_7506,N_7514);
nand U8881 (N_8881,N_7515,N_7972);
nand U8882 (N_8882,N_7521,N_8038);
and U8883 (N_8883,N_7917,N_7655);
nor U8884 (N_8884,N_7880,N_7829);
xor U8885 (N_8885,N_8083,N_7527);
nor U8886 (N_8886,N_7652,N_8116);
xnor U8887 (N_8887,N_7766,N_7730);
or U8888 (N_8888,N_7602,N_7968);
and U8889 (N_8889,N_7697,N_7577);
or U8890 (N_8890,N_8197,N_7585);
nand U8891 (N_8891,N_8094,N_8081);
and U8892 (N_8892,N_8072,N_7631);
nor U8893 (N_8893,N_7883,N_8052);
and U8894 (N_8894,N_7834,N_7970);
nand U8895 (N_8895,N_8135,N_8190);
nand U8896 (N_8896,N_7801,N_7931);
or U8897 (N_8897,N_7796,N_8143);
nand U8898 (N_8898,N_7835,N_7669);
nor U8899 (N_8899,N_7553,N_8146);
nand U8900 (N_8900,N_7600,N_7721);
nand U8901 (N_8901,N_8180,N_8000);
or U8902 (N_8902,N_7837,N_7615);
or U8903 (N_8903,N_7914,N_7559);
nor U8904 (N_8904,N_7535,N_8197);
or U8905 (N_8905,N_7830,N_8211);
and U8906 (N_8906,N_7728,N_8042);
nor U8907 (N_8907,N_7817,N_7973);
and U8908 (N_8908,N_7809,N_7964);
xnor U8909 (N_8909,N_7894,N_7679);
nand U8910 (N_8910,N_7830,N_8145);
xnor U8911 (N_8911,N_7527,N_7568);
nand U8912 (N_8912,N_8082,N_8243);
and U8913 (N_8913,N_8022,N_7503);
or U8914 (N_8914,N_7624,N_7944);
nor U8915 (N_8915,N_8089,N_7691);
and U8916 (N_8916,N_7961,N_8229);
or U8917 (N_8917,N_7667,N_7772);
xor U8918 (N_8918,N_8151,N_7685);
or U8919 (N_8919,N_7522,N_7851);
nor U8920 (N_8920,N_7800,N_7864);
nand U8921 (N_8921,N_7865,N_7575);
or U8922 (N_8922,N_7666,N_7922);
or U8923 (N_8923,N_7918,N_7911);
or U8924 (N_8924,N_7710,N_8027);
or U8925 (N_8925,N_7664,N_7852);
nor U8926 (N_8926,N_7929,N_8188);
nand U8927 (N_8927,N_7868,N_8181);
and U8928 (N_8928,N_8010,N_7648);
or U8929 (N_8929,N_7765,N_7593);
and U8930 (N_8930,N_7848,N_7552);
xor U8931 (N_8931,N_7968,N_7656);
or U8932 (N_8932,N_7504,N_7946);
xnor U8933 (N_8933,N_7517,N_7703);
nand U8934 (N_8934,N_7517,N_8083);
nor U8935 (N_8935,N_8072,N_7856);
and U8936 (N_8936,N_7963,N_8238);
nand U8937 (N_8937,N_7575,N_7506);
nand U8938 (N_8938,N_7814,N_7792);
nand U8939 (N_8939,N_8062,N_8053);
nor U8940 (N_8940,N_7893,N_8230);
nor U8941 (N_8941,N_8239,N_7995);
xor U8942 (N_8942,N_8026,N_8083);
or U8943 (N_8943,N_7675,N_8089);
nor U8944 (N_8944,N_8114,N_8193);
nor U8945 (N_8945,N_7587,N_7538);
nand U8946 (N_8946,N_8227,N_7661);
nor U8947 (N_8947,N_7972,N_7820);
nor U8948 (N_8948,N_7987,N_7722);
nand U8949 (N_8949,N_8106,N_7659);
xor U8950 (N_8950,N_7860,N_8111);
and U8951 (N_8951,N_8098,N_8109);
xnor U8952 (N_8952,N_8015,N_7527);
nor U8953 (N_8953,N_7849,N_7781);
or U8954 (N_8954,N_7740,N_8202);
nand U8955 (N_8955,N_8220,N_7987);
and U8956 (N_8956,N_8167,N_7606);
and U8957 (N_8957,N_7896,N_7761);
nor U8958 (N_8958,N_8033,N_7909);
nor U8959 (N_8959,N_7675,N_7925);
or U8960 (N_8960,N_8112,N_8135);
nor U8961 (N_8961,N_7552,N_7720);
nor U8962 (N_8962,N_8205,N_7928);
or U8963 (N_8963,N_7719,N_7658);
or U8964 (N_8964,N_7859,N_7554);
or U8965 (N_8965,N_8095,N_7611);
or U8966 (N_8966,N_7594,N_8142);
or U8967 (N_8967,N_7877,N_8101);
nor U8968 (N_8968,N_8014,N_8075);
nor U8969 (N_8969,N_8138,N_7577);
and U8970 (N_8970,N_7826,N_7502);
or U8971 (N_8971,N_8245,N_7720);
nor U8972 (N_8972,N_8102,N_7680);
and U8973 (N_8973,N_7765,N_8020);
or U8974 (N_8974,N_7870,N_7777);
nor U8975 (N_8975,N_7973,N_7672);
or U8976 (N_8976,N_7726,N_7882);
or U8977 (N_8977,N_7880,N_7515);
nor U8978 (N_8978,N_7607,N_8076);
or U8979 (N_8979,N_7693,N_7510);
nand U8980 (N_8980,N_8165,N_7565);
xor U8981 (N_8981,N_7796,N_8198);
nor U8982 (N_8982,N_7546,N_8032);
or U8983 (N_8983,N_7648,N_8046);
nor U8984 (N_8984,N_8222,N_7711);
xnor U8985 (N_8985,N_7629,N_8076);
xor U8986 (N_8986,N_7571,N_7525);
and U8987 (N_8987,N_8024,N_8180);
nor U8988 (N_8988,N_8044,N_8164);
or U8989 (N_8989,N_8137,N_7946);
and U8990 (N_8990,N_7615,N_8183);
or U8991 (N_8991,N_7646,N_8227);
nand U8992 (N_8992,N_7603,N_7552);
and U8993 (N_8993,N_8135,N_7518);
nor U8994 (N_8994,N_7698,N_7717);
nand U8995 (N_8995,N_8223,N_7569);
and U8996 (N_8996,N_7527,N_7691);
nor U8997 (N_8997,N_7747,N_8073);
and U8998 (N_8998,N_7591,N_7528);
and U8999 (N_8999,N_7724,N_7657);
or U9000 (N_9000,N_8880,N_8730);
nand U9001 (N_9001,N_8892,N_8536);
nor U9002 (N_9002,N_8311,N_8985);
nor U9003 (N_9003,N_8390,N_8821);
nand U9004 (N_9004,N_8849,N_8703);
nor U9005 (N_9005,N_8796,N_8261);
xnor U9006 (N_9006,N_8498,N_8296);
or U9007 (N_9007,N_8523,N_8722);
and U9008 (N_9008,N_8607,N_8287);
nor U9009 (N_9009,N_8344,N_8857);
nand U9010 (N_9010,N_8733,N_8956);
nand U9011 (N_9011,N_8830,N_8527);
nand U9012 (N_9012,N_8548,N_8391);
or U9013 (N_9013,N_8786,N_8621);
nor U9014 (N_9014,N_8451,N_8824);
and U9015 (N_9015,N_8575,N_8915);
and U9016 (N_9016,N_8931,N_8445);
nand U9017 (N_9017,N_8411,N_8468);
and U9018 (N_9018,N_8834,N_8590);
nor U9019 (N_9019,N_8691,N_8528);
and U9020 (N_9020,N_8677,N_8283);
nand U9021 (N_9021,N_8347,N_8917);
or U9022 (N_9022,N_8401,N_8842);
or U9023 (N_9023,N_8362,N_8480);
nor U9024 (N_9024,N_8508,N_8255);
nor U9025 (N_9025,N_8663,N_8841);
and U9026 (N_9026,N_8476,N_8592);
or U9027 (N_9027,N_8585,N_8647);
nor U9028 (N_9028,N_8970,N_8534);
nor U9029 (N_9029,N_8509,N_8701);
nand U9030 (N_9030,N_8884,N_8304);
nor U9031 (N_9031,N_8823,N_8763);
or U9032 (N_9032,N_8544,N_8826);
nand U9033 (N_9033,N_8692,N_8573);
nor U9034 (N_9034,N_8455,N_8955);
nor U9035 (N_9035,N_8952,N_8962);
nand U9036 (N_9036,N_8790,N_8872);
nand U9037 (N_9037,N_8765,N_8943);
or U9038 (N_9038,N_8470,N_8812);
nand U9039 (N_9039,N_8695,N_8811);
nor U9040 (N_9040,N_8993,N_8557);
nor U9041 (N_9041,N_8555,N_8697);
nor U9042 (N_9042,N_8650,N_8937);
and U9043 (N_9043,N_8282,N_8665);
or U9044 (N_9044,N_8297,N_8268);
xnor U9045 (N_9045,N_8804,N_8443);
xnor U9046 (N_9046,N_8537,N_8761);
or U9047 (N_9047,N_8949,N_8721);
nand U9048 (N_9048,N_8351,N_8335);
nand U9049 (N_9049,N_8632,N_8977);
xnor U9050 (N_9050,N_8807,N_8623);
or U9051 (N_9051,N_8800,N_8314);
nor U9052 (N_9052,N_8403,N_8641);
nand U9053 (N_9053,N_8518,N_8405);
or U9054 (N_9054,N_8628,N_8615);
nor U9055 (N_9055,N_8373,N_8364);
and U9056 (N_9056,N_8904,N_8618);
nor U9057 (N_9057,N_8348,N_8899);
nand U9058 (N_9058,N_8419,N_8979);
nor U9059 (N_9059,N_8930,N_8612);
nand U9060 (N_9060,N_8846,N_8617);
xnor U9061 (N_9061,N_8700,N_8376);
or U9062 (N_9062,N_8770,N_8400);
xnor U9063 (N_9063,N_8978,N_8291);
and U9064 (N_9064,N_8777,N_8549);
xnor U9065 (N_9065,N_8630,N_8504);
nand U9066 (N_9066,N_8803,N_8859);
nor U9067 (N_9067,N_8748,N_8572);
nor U9068 (N_9068,N_8689,N_8467);
or U9069 (N_9069,N_8731,N_8906);
and U9070 (N_9070,N_8781,N_8942);
or U9071 (N_9071,N_8600,N_8698);
nor U9072 (N_9072,N_8622,N_8472);
nor U9073 (N_9073,N_8512,N_8254);
or U9074 (N_9074,N_8810,N_8975);
nor U9075 (N_9075,N_8659,N_8764);
or U9076 (N_9076,N_8881,N_8945);
or U9077 (N_9077,N_8901,N_8588);
xor U9078 (N_9078,N_8798,N_8624);
or U9079 (N_9079,N_8564,N_8683);
or U9080 (N_9080,N_8936,N_8421);
nand U9081 (N_9081,N_8656,N_8744);
nor U9082 (N_9082,N_8896,N_8374);
nor U9083 (N_9083,N_8346,N_8870);
nor U9084 (N_9084,N_8717,N_8305);
and U9085 (N_9085,N_8513,N_8642);
nor U9086 (N_9086,N_8613,N_8619);
nand U9087 (N_9087,N_8379,N_8666);
and U9088 (N_9088,N_8569,N_8960);
nand U9089 (N_9089,N_8449,N_8320);
nor U9090 (N_9090,N_8558,N_8843);
or U9091 (N_9091,N_8797,N_8357);
nand U9092 (N_9092,N_8394,N_8384);
nor U9093 (N_9093,N_8599,N_8990);
xnor U9094 (N_9094,N_8827,N_8535);
nor U9095 (N_9095,N_8516,N_8771);
or U9096 (N_9096,N_8933,N_8370);
nor U9097 (N_9097,N_8345,N_8462);
nand U9098 (N_9098,N_8319,N_8385);
and U9099 (N_9099,N_8383,N_8999);
or U9100 (N_9100,N_8889,N_8490);
nor U9101 (N_9101,N_8290,N_8487);
xnor U9102 (N_9102,N_8505,N_8660);
and U9103 (N_9103,N_8340,N_8271);
and U9104 (N_9104,N_8920,N_8678);
nor U9105 (N_9105,N_8844,N_8969);
xor U9106 (N_9106,N_8277,N_8724);
nor U9107 (N_9107,N_8773,N_8483);
or U9108 (N_9108,N_8597,N_8668);
xnor U9109 (N_9109,N_8308,N_8946);
or U9110 (N_9110,N_8300,N_8629);
or U9111 (N_9111,N_8414,N_8716);
nand U9112 (N_9112,N_8778,N_8785);
nand U9113 (N_9113,N_8669,N_8372);
nor U9114 (N_9114,N_8735,N_8637);
and U9115 (N_9115,N_8301,N_8402);
xor U9116 (N_9116,N_8316,N_8732);
nand U9117 (N_9117,N_8958,N_8482);
nor U9118 (N_9118,N_8435,N_8742);
xor U9119 (N_9119,N_8540,N_8822);
xnor U9120 (N_9120,N_8986,N_8725);
and U9121 (N_9121,N_8727,N_8634);
or U9122 (N_9122,N_8448,N_8654);
nand U9123 (N_9123,N_8416,N_8309);
nor U9124 (N_9124,N_8438,N_8336);
or U9125 (N_9125,N_8649,N_8329);
or U9126 (N_9126,N_8550,N_8926);
and U9127 (N_9127,N_8802,N_8444);
and U9128 (N_9128,N_8782,N_8878);
or U9129 (N_9129,N_8753,N_8941);
or U9130 (N_9130,N_8801,N_8871);
or U9131 (N_9131,N_8963,N_8829);
nor U9132 (N_9132,N_8503,N_8358);
nor U9133 (N_9133,N_8938,N_8762);
or U9134 (N_9134,N_8552,N_8586);
and U9135 (N_9135,N_8974,N_8746);
or U9136 (N_9136,N_8602,N_8371);
nand U9137 (N_9137,N_8295,N_8350);
nor U9138 (N_9138,N_8886,N_8664);
nor U9139 (N_9139,N_8489,N_8767);
nand U9140 (N_9140,N_8813,N_8521);
and U9141 (N_9141,N_8948,N_8614);
or U9142 (N_9142,N_8966,N_8428);
and U9143 (N_9143,N_8601,N_8363);
and U9144 (N_9144,N_8627,N_8837);
xor U9145 (N_9145,N_8808,N_8574);
and U9146 (N_9146,N_8356,N_8758);
nor U9147 (N_9147,N_8595,N_8288);
and U9148 (N_9148,N_8299,N_8995);
nor U9149 (N_9149,N_8820,N_8934);
and U9150 (N_9150,N_8638,N_8852);
or U9151 (N_9151,N_8631,N_8780);
and U9152 (N_9152,N_8582,N_8606);
and U9153 (N_9153,N_8737,N_8519);
and U9154 (N_9154,N_8479,N_8833);
or U9155 (N_9155,N_8863,N_8431);
nand U9156 (N_9156,N_8578,N_8968);
or U9157 (N_9157,N_8420,N_8662);
nor U9158 (N_9158,N_8988,N_8752);
or U9159 (N_9159,N_8825,N_8532);
and U9160 (N_9160,N_8708,N_8253);
nor U9161 (N_9161,N_8893,N_8322);
and U9162 (N_9162,N_8747,N_8991);
or U9163 (N_9163,N_8422,N_8667);
nand U9164 (N_9164,N_8729,N_8911);
nand U9165 (N_9165,N_8787,N_8603);
nand U9166 (N_9166,N_8567,N_8760);
nand U9167 (N_9167,N_8858,N_8835);
nor U9168 (N_9168,N_8789,N_8581);
nor U9169 (N_9169,N_8559,N_8954);
nand U9170 (N_9170,N_8965,N_8424);
nor U9171 (N_9171,N_8561,N_8398);
nand U9172 (N_9172,N_8743,N_8989);
xor U9173 (N_9173,N_8369,N_8263);
and U9174 (N_9174,N_8452,N_8457);
xor U9175 (N_9175,N_8570,N_8556);
nand U9176 (N_9176,N_8658,N_8755);
and U9177 (N_9177,N_8961,N_8869);
nand U9178 (N_9178,N_8341,N_8593);
nor U9179 (N_9179,N_8705,N_8332);
nand U9180 (N_9180,N_8276,N_8973);
nor U9181 (N_9181,N_8339,N_8895);
nor U9182 (N_9182,N_8262,N_8699);
and U9183 (N_9183,N_8657,N_8325);
nand U9184 (N_9184,N_8888,N_8831);
or U9185 (N_9185,N_8382,N_8909);
or U9186 (N_9186,N_8980,N_8323);
nor U9187 (N_9187,N_8809,N_8851);
nand U9188 (N_9188,N_8776,N_8873);
or U9189 (N_9189,N_8694,N_8684);
or U9190 (N_9190,N_8333,N_8475);
nand U9191 (N_9191,N_8494,N_8343);
nor U9192 (N_9192,N_8759,N_8427);
nand U9193 (N_9193,N_8604,N_8571);
or U9194 (N_9194,N_8784,N_8805);
nand U9195 (N_9195,N_8792,N_8696);
nor U9196 (N_9196,N_8935,N_8473);
and U9197 (N_9197,N_8832,N_8693);
or U9198 (N_9198,N_8736,N_8298);
nand U9199 (N_9199,N_8486,N_8441);
nor U9200 (N_9200,N_8496,N_8608);
and U9201 (N_9201,N_8326,N_8576);
or U9202 (N_9202,N_8655,N_8531);
or U9203 (N_9203,N_8524,N_8779);
nand U9204 (N_9204,N_8616,N_8580);
nor U9205 (N_9205,N_8688,N_8853);
nand U9206 (N_9206,N_8653,N_8542);
nor U9207 (N_9207,N_8375,N_8266);
nor U9208 (N_9208,N_8404,N_8506);
and U9209 (N_9209,N_8815,N_8442);
or U9210 (N_9210,N_8750,N_8367);
or U9211 (N_9211,N_8415,N_8563);
or U9212 (N_9212,N_8690,N_8676);
or U9213 (N_9213,N_8543,N_8610);
xor U9214 (N_9214,N_8992,N_8719);
and U9215 (N_9215,N_8799,N_8738);
nand U9216 (N_9216,N_8587,N_8284);
or U9217 (N_9217,N_8817,N_8636);
nand U9218 (N_9218,N_8754,N_8710);
or U9219 (N_9219,N_8495,N_8547);
xnor U9220 (N_9220,N_8436,N_8591);
nand U9221 (N_9221,N_8366,N_8950);
nand U9222 (N_9222,N_8897,N_8269);
nand U9223 (N_9223,N_8791,N_8806);
nor U9224 (N_9224,N_8568,N_8429);
and U9225 (N_9225,N_8740,N_8426);
xnor U9226 (N_9226,N_8640,N_8940);
or U9227 (N_9227,N_8397,N_8605);
or U9228 (N_9228,N_8947,N_8353);
and U9229 (N_9229,N_8440,N_8996);
and U9230 (N_9230,N_8517,N_8868);
nand U9231 (N_9231,N_8775,N_8279);
and U9232 (N_9232,N_8685,N_8944);
nand U9233 (N_9233,N_8596,N_8551);
or U9234 (N_9234,N_8471,N_8741);
and U9235 (N_9235,N_8598,N_8407);
and U9236 (N_9236,N_8274,N_8877);
nand U9237 (N_9237,N_8499,N_8959);
and U9238 (N_9238,N_8439,N_8739);
and U9239 (N_9239,N_8987,N_8432);
nor U9240 (N_9240,N_8515,N_8997);
nand U9241 (N_9241,N_8360,N_8646);
and U9242 (N_9242,N_8795,N_8355);
nand U9243 (N_9243,N_8929,N_8458);
or U9244 (N_9244,N_8294,N_8611);
nand U9245 (N_9245,N_8919,N_8334);
and U9246 (N_9246,N_8460,N_8713);
and U9247 (N_9247,N_8259,N_8625);
nor U9248 (N_9248,N_8313,N_8768);
nand U9249 (N_9249,N_8981,N_8365);
or U9250 (N_9250,N_8546,N_8644);
nand U9251 (N_9251,N_8887,N_8756);
xor U9252 (N_9252,N_8545,N_8387);
or U9253 (N_9253,N_8533,N_8839);
xnor U9254 (N_9254,N_8406,N_8273);
nor U9255 (N_9255,N_8794,N_8256);
xnor U9256 (N_9256,N_8984,N_8459);
or U9257 (N_9257,N_8749,N_8718);
and U9258 (N_9258,N_8310,N_8891);
and U9259 (N_9259,N_8285,N_8328);
nor U9260 (N_9260,N_8399,N_8876);
nor U9261 (N_9261,N_8715,N_8643);
and U9262 (N_9262,N_8315,N_8894);
nand U9263 (N_9263,N_8270,N_8417);
nand U9264 (N_9264,N_8908,N_8306);
and U9265 (N_9265,N_8928,N_8258);
nor U9266 (N_9266,N_8652,N_8265);
nand U9267 (N_9267,N_8447,N_8418);
and U9268 (N_9268,N_8502,N_8712);
or U9269 (N_9269,N_8951,N_8478);
or U9270 (N_9270,N_8264,N_8251);
or U9271 (N_9271,N_8850,N_8885);
and U9272 (N_9272,N_8539,N_8395);
and U9273 (N_9273,N_8349,N_8324);
or U9274 (N_9274,N_8648,N_8845);
nor U9275 (N_9275,N_8393,N_8312);
and U9276 (N_9276,N_8267,N_8932);
xor U9277 (N_9277,N_8354,N_8711);
nand U9278 (N_9278,N_8983,N_8620);
or U9279 (N_9279,N_8307,N_8454);
and U9280 (N_9280,N_8957,N_8425);
nand U9281 (N_9281,N_8635,N_8566);
and U9282 (N_9282,N_8879,N_8882);
nor U9283 (N_9283,N_8766,N_8774);
xor U9284 (N_9284,N_8529,N_8964);
and U9285 (N_9285,N_8900,N_8862);
nor U9286 (N_9286,N_8651,N_8673);
or U9287 (N_9287,N_8783,N_8412);
and U9288 (N_9288,N_8840,N_8589);
and U9289 (N_9289,N_8709,N_8672);
xnor U9290 (N_9290,N_8318,N_8816);
or U9291 (N_9291,N_8914,N_8953);
and U9292 (N_9292,N_8772,N_8286);
nor U9293 (N_9293,N_8745,N_8679);
or U9294 (N_9294,N_8302,N_8446);
or U9295 (N_9295,N_8331,N_8507);
and U9296 (N_9296,N_8702,N_8898);
nand U9297 (N_9297,N_8706,N_8481);
and U9298 (N_9298,N_8492,N_8994);
and U9299 (N_9299,N_8707,N_8982);
nand U9300 (N_9300,N_8437,N_8463);
nor U9301 (N_9301,N_8485,N_8413);
nand U9302 (N_9302,N_8626,N_8814);
nand U9303 (N_9303,N_8793,N_8865);
nand U9304 (N_9304,N_8303,N_8594);
or U9305 (N_9305,N_8510,N_8565);
nand U9306 (N_9306,N_8861,N_8562);
and U9307 (N_9307,N_8338,N_8864);
and U9308 (N_9308,N_8337,N_8674);
nor U9309 (N_9309,N_8874,N_8728);
and U9310 (N_9310,N_8866,N_8609);
xnor U9311 (N_9311,N_8723,N_8916);
or U9312 (N_9312,N_8396,N_8939);
nand U9313 (N_9313,N_8769,N_8292);
and U9314 (N_9314,N_8456,N_8726);
xnor U9315 (N_9315,N_8560,N_8280);
and U9316 (N_9316,N_8686,N_8681);
nor U9317 (N_9317,N_8670,N_8584);
or U9318 (N_9318,N_8359,N_8520);
or U9319 (N_9319,N_8912,N_8491);
nand U9320 (N_9320,N_8890,N_8967);
and U9321 (N_9321,N_8327,N_8477);
or U9322 (N_9322,N_8704,N_8461);
or U9323 (N_9323,N_8522,N_8579);
nor U9324 (N_9324,N_8847,N_8819);
nor U9325 (N_9325,N_8860,N_8918);
and U9326 (N_9326,N_8828,N_8720);
nor U9327 (N_9327,N_8583,N_8924);
nand U9328 (N_9328,N_8464,N_8927);
xor U9329 (N_9329,N_8466,N_8925);
nor U9330 (N_9330,N_8388,N_8921);
or U9331 (N_9331,N_8818,N_8633);
or U9332 (N_9332,N_8433,N_8317);
nand U9333 (N_9333,N_8905,N_8493);
or U9334 (N_9334,N_8321,N_8484);
or U9335 (N_9335,N_8361,N_8856);
or U9336 (N_9336,N_8903,N_8675);
or U9337 (N_9337,N_8553,N_8577);
nor U9338 (N_9338,N_8788,N_8381);
nand U9339 (N_9339,N_8453,N_8902);
nor U9340 (N_9340,N_8867,N_8410);
and U9341 (N_9341,N_8500,N_8278);
and U9342 (N_9342,N_8250,N_8687);
xor U9343 (N_9343,N_8971,N_8751);
xnor U9344 (N_9344,N_8511,N_8514);
xor U9345 (N_9345,N_8639,N_8836);
nand U9346 (N_9346,N_8378,N_8734);
and U9347 (N_9347,N_8910,N_8554);
and U9348 (N_9348,N_8392,N_8377);
and U9349 (N_9349,N_8293,N_8469);
and U9350 (N_9350,N_8525,N_8913);
nand U9351 (N_9351,N_8998,N_8538);
nand U9352 (N_9352,N_8883,N_8474);
xor U9353 (N_9353,N_8838,N_8423);
nor U9354 (N_9354,N_8342,N_8281);
nor U9355 (N_9355,N_8352,N_8923);
and U9356 (N_9356,N_8976,N_8855);
nand U9357 (N_9357,N_8289,N_8330);
nand U9358 (N_9358,N_8430,N_8380);
nor U9359 (N_9359,N_8386,N_8257);
xor U9360 (N_9360,N_8530,N_8680);
or U9361 (N_9361,N_8526,N_8671);
and U9362 (N_9362,N_8757,N_8501);
and U9363 (N_9363,N_8450,N_8972);
or U9364 (N_9364,N_8260,N_8275);
nor U9365 (N_9365,N_8661,N_8389);
nand U9366 (N_9366,N_8488,N_8252);
nand U9367 (N_9367,N_8434,N_8922);
or U9368 (N_9368,N_8645,N_8408);
nor U9369 (N_9369,N_8497,N_8682);
and U9370 (N_9370,N_8907,N_8848);
nor U9371 (N_9371,N_8409,N_8714);
nor U9372 (N_9372,N_8875,N_8272);
or U9373 (N_9373,N_8465,N_8541);
nor U9374 (N_9374,N_8854,N_8368);
nor U9375 (N_9375,N_8816,N_8636);
xnor U9376 (N_9376,N_8507,N_8393);
xnor U9377 (N_9377,N_8279,N_8760);
xor U9378 (N_9378,N_8338,N_8372);
nand U9379 (N_9379,N_8691,N_8860);
nor U9380 (N_9380,N_8638,N_8933);
xor U9381 (N_9381,N_8473,N_8750);
nor U9382 (N_9382,N_8911,N_8918);
nand U9383 (N_9383,N_8645,N_8444);
or U9384 (N_9384,N_8542,N_8744);
nand U9385 (N_9385,N_8697,N_8623);
or U9386 (N_9386,N_8687,N_8583);
and U9387 (N_9387,N_8723,N_8601);
or U9388 (N_9388,N_8336,N_8746);
or U9389 (N_9389,N_8688,N_8861);
and U9390 (N_9390,N_8269,N_8376);
or U9391 (N_9391,N_8379,N_8604);
nand U9392 (N_9392,N_8258,N_8278);
nor U9393 (N_9393,N_8847,N_8544);
xnor U9394 (N_9394,N_8445,N_8900);
and U9395 (N_9395,N_8350,N_8940);
nand U9396 (N_9396,N_8994,N_8301);
or U9397 (N_9397,N_8943,N_8915);
and U9398 (N_9398,N_8488,N_8442);
and U9399 (N_9399,N_8569,N_8937);
nand U9400 (N_9400,N_8907,N_8710);
xnor U9401 (N_9401,N_8586,N_8711);
and U9402 (N_9402,N_8663,N_8591);
or U9403 (N_9403,N_8831,N_8980);
nand U9404 (N_9404,N_8288,N_8336);
nor U9405 (N_9405,N_8681,N_8435);
or U9406 (N_9406,N_8932,N_8372);
or U9407 (N_9407,N_8861,N_8770);
and U9408 (N_9408,N_8779,N_8827);
nor U9409 (N_9409,N_8622,N_8704);
and U9410 (N_9410,N_8972,N_8782);
nor U9411 (N_9411,N_8561,N_8944);
nand U9412 (N_9412,N_8377,N_8741);
xor U9413 (N_9413,N_8613,N_8965);
or U9414 (N_9414,N_8909,N_8549);
xnor U9415 (N_9415,N_8564,N_8322);
nand U9416 (N_9416,N_8481,N_8523);
or U9417 (N_9417,N_8733,N_8759);
nor U9418 (N_9418,N_8721,N_8432);
or U9419 (N_9419,N_8294,N_8942);
nand U9420 (N_9420,N_8321,N_8651);
nor U9421 (N_9421,N_8411,N_8823);
nand U9422 (N_9422,N_8885,N_8309);
and U9423 (N_9423,N_8264,N_8352);
or U9424 (N_9424,N_8720,N_8695);
nand U9425 (N_9425,N_8965,N_8415);
nand U9426 (N_9426,N_8685,N_8590);
and U9427 (N_9427,N_8528,N_8794);
or U9428 (N_9428,N_8683,N_8626);
nor U9429 (N_9429,N_8825,N_8657);
nor U9430 (N_9430,N_8853,N_8714);
nand U9431 (N_9431,N_8454,N_8487);
nand U9432 (N_9432,N_8381,N_8611);
and U9433 (N_9433,N_8697,N_8362);
nor U9434 (N_9434,N_8479,N_8787);
nor U9435 (N_9435,N_8431,N_8855);
nand U9436 (N_9436,N_8357,N_8466);
nand U9437 (N_9437,N_8269,N_8490);
and U9438 (N_9438,N_8973,N_8836);
and U9439 (N_9439,N_8988,N_8906);
xnor U9440 (N_9440,N_8462,N_8620);
nor U9441 (N_9441,N_8337,N_8905);
nor U9442 (N_9442,N_8845,N_8381);
xnor U9443 (N_9443,N_8374,N_8449);
and U9444 (N_9444,N_8682,N_8903);
or U9445 (N_9445,N_8541,N_8429);
and U9446 (N_9446,N_8429,N_8387);
nor U9447 (N_9447,N_8715,N_8910);
nor U9448 (N_9448,N_8309,N_8704);
xor U9449 (N_9449,N_8755,N_8535);
or U9450 (N_9450,N_8665,N_8527);
nand U9451 (N_9451,N_8879,N_8348);
nand U9452 (N_9452,N_8719,N_8753);
xnor U9453 (N_9453,N_8397,N_8362);
and U9454 (N_9454,N_8962,N_8569);
nor U9455 (N_9455,N_8539,N_8316);
nand U9456 (N_9456,N_8962,N_8920);
or U9457 (N_9457,N_8656,N_8498);
xnor U9458 (N_9458,N_8261,N_8813);
or U9459 (N_9459,N_8381,N_8775);
or U9460 (N_9460,N_8948,N_8421);
or U9461 (N_9461,N_8316,N_8778);
nor U9462 (N_9462,N_8700,N_8631);
nor U9463 (N_9463,N_8457,N_8256);
nor U9464 (N_9464,N_8904,N_8368);
nand U9465 (N_9465,N_8603,N_8492);
or U9466 (N_9466,N_8995,N_8910);
or U9467 (N_9467,N_8662,N_8749);
nand U9468 (N_9468,N_8744,N_8345);
and U9469 (N_9469,N_8688,N_8514);
xor U9470 (N_9470,N_8723,N_8540);
and U9471 (N_9471,N_8675,N_8900);
nor U9472 (N_9472,N_8866,N_8626);
nand U9473 (N_9473,N_8579,N_8966);
nand U9474 (N_9474,N_8384,N_8715);
and U9475 (N_9475,N_8702,N_8498);
nor U9476 (N_9476,N_8786,N_8816);
or U9477 (N_9477,N_8699,N_8878);
or U9478 (N_9478,N_8708,N_8748);
nand U9479 (N_9479,N_8526,N_8817);
and U9480 (N_9480,N_8370,N_8994);
nand U9481 (N_9481,N_8721,N_8870);
nor U9482 (N_9482,N_8857,N_8614);
nor U9483 (N_9483,N_8825,N_8999);
nor U9484 (N_9484,N_8257,N_8675);
nand U9485 (N_9485,N_8726,N_8721);
and U9486 (N_9486,N_8295,N_8710);
and U9487 (N_9487,N_8784,N_8709);
nand U9488 (N_9488,N_8610,N_8734);
or U9489 (N_9489,N_8345,N_8844);
and U9490 (N_9490,N_8388,N_8649);
or U9491 (N_9491,N_8634,N_8914);
nor U9492 (N_9492,N_8919,N_8867);
nand U9493 (N_9493,N_8862,N_8515);
and U9494 (N_9494,N_8800,N_8297);
nand U9495 (N_9495,N_8547,N_8872);
or U9496 (N_9496,N_8809,N_8446);
nand U9497 (N_9497,N_8289,N_8986);
and U9498 (N_9498,N_8712,N_8325);
and U9499 (N_9499,N_8495,N_8713);
nor U9500 (N_9500,N_8884,N_8927);
or U9501 (N_9501,N_8363,N_8821);
and U9502 (N_9502,N_8963,N_8308);
or U9503 (N_9503,N_8917,N_8890);
nand U9504 (N_9504,N_8536,N_8667);
nand U9505 (N_9505,N_8831,N_8623);
nor U9506 (N_9506,N_8654,N_8544);
nand U9507 (N_9507,N_8421,N_8978);
nor U9508 (N_9508,N_8390,N_8311);
or U9509 (N_9509,N_8520,N_8659);
and U9510 (N_9510,N_8555,N_8444);
and U9511 (N_9511,N_8935,N_8276);
and U9512 (N_9512,N_8779,N_8417);
and U9513 (N_9513,N_8886,N_8300);
and U9514 (N_9514,N_8915,N_8462);
nor U9515 (N_9515,N_8470,N_8292);
nor U9516 (N_9516,N_8852,N_8907);
nand U9517 (N_9517,N_8308,N_8703);
nor U9518 (N_9518,N_8645,N_8415);
or U9519 (N_9519,N_8491,N_8780);
nor U9520 (N_9520,N_8471,N_8355);
nor U9521 (N_9521,N_8710,N_8634);
nand U9522 (N_9522,N_8597,N_8516);
or U9523 (N_9523,N_8994,N_8717);
or U9524 (N_9524,N_8989,N_8967);
nand U9525 (N_9525,N_8437,N_8454);
nor U9526 (N_9526,N_8435,N_8467);
or U9527 (N_9527,N_8870,N_8682);
nand U9528 (N_9528,N_8561,N_8330);
nand U9529 (N_9529,N_8735,N_8740);
nor U9530 (N_9530,N_8459,N_8724);
and U9531 (N_9531,N_8653,N_8940);
nor U9532 (N_9532,N_8538,N_8771);
nor U9533 (N_9533,N_8426,N_8436);
or U9534 (N_9534,N_8578,N_8569);
xor U9535 (N_9535,N_8977,N_8978);
nor U9536 (N_9536,N_8261,N_8532);
nor U9537 (N_9537,N_8620,N_8785);
nand U9538 (N_9538,N_8801,N_8507);
or U9539 (N_9539,N_8433,N_8811);
nor U9540 (N_9540,N_8830,N_8576);
and U9541 (N_9541,N_8877,N_8661);
nor U9542 (N_9542,N_8607,N_8747);
xnor U9543 (N_9543,N_8939,N_8570);
or U9544 (N_9544,N_8369,N_8903);
and U9545 (N_9545,N_8832,N_8769);
or U9546 (N_9546,N_8865,N_8624);
nor U9547 (N_9547,N_8615,N_8463);
or U9548 (N_9548,N_8296,N_8702);
nor U9549 (N_9549,N_8979,N_8888);
and U9550 (N_9550,N_8841,N_8438);
and U9551 (N_9551,N_8401,N_8623);
nand U9552 (N_9552,N_8274,N_8978);
or U9553 (N_9553,N_8897,N_8457);
and U9554 (N_9554,N_8573,N_8417);
nand U9555 (N_9555,N_8462,N_8831);
or U9556 (N_9556,N_8314,N_8605);
and U9557 (N_9557,N_8871,N_8363);
or U9558 (N_9558,N_8938,N_8518);
and U9559 (N_9559,N_8642,N_8348);
nor U9560 (N_9560,N_8480,N_8804);
nand U9561 (N_9561,N_8613,N_8660);
and U9562 (N_9562,N_8973,N_8756);
nand U9563 (N_9563,N_8986,N_8579);
and U9564 (N_9564,N_8537,N_8487);
nor U9565 (N_9565,N_8283,N_8698);
nand U9566 (N_9566,N_8601,N_8965);
xor U9567 (N_9567,N_8500,N_8269);
nor U9568 (N_9568,N_8758,N_8313);
or U9569 (N_9569,N_8255,N_8536);
or U9570 (N_9570,N_8912,N_8901);
or U9571 (N_9571,N_8492,N_8928);
nor U9572 (N_9572,N_8342,N_8267);
xor U9573 (N_9573,N_8598,N_8267);
or U9574 (N_9574,N_8865,N_8353);
or U9575 (N_9575,N_8366,N_8654);
nor U9576 (N_9576,N_8536,N_8993);
nand U9577 (N_9577,N_8565,N_8548);
nand U9578 (N_9578,N_8255,N_8296);
nor U9579 (N_9579,N_8374,N_8579);
xor U9580 (N_9580,N_8503,N_8736);
or U9581 (N_9581,N_8314,N_8349);
xor U9582 (N_9582,N_8383,N_8425);
or U9583 (N_9583,N_8714,N_8811);
nor U9584 (N_9584,N_8658,N_8360);
nand U9585 (N_9585,N_8573,N_8420);
nand U9586 (N_9586,N_8727,N_8376);
nand U9587 (N_9587,N_8503,N_8588);
nor U9588 (N_9588,N_8472,N_8872);
and U9589 (N_9589,N_8405,N_8640);
xor U9590 (N_9590,N_8278,N_8966);
and U9591 (N_9591,N_8424,N_8494);
nand U9592 (N_9592,N_8498,N_8847);
and U9593 (N_9593,N_8318,N_8499);
or U9594 (N_9594,N_8639,N_8439);
nand U9595 (N_9595,N_8286,N_8604);
nor U9596 (N_9596,N_8322,N_8850);
or U9597 (N_9597,N_8734,N_8274);
or U9598 (N_9598,N_8696,N_8623);
nor U9599 (N_9599,N_8341,N_8796);
nor U9600 (N_9600,N_8515,N_8575);
nand U9601 (N_9601,N_8682,N_8677);
nor U9602 (N_9602,N_8851,N_8972);
and U9603 (N_9603,N_8959,N_8699);
nand U9604 (N_9604,N_8624,N_8907);
nand U9605 (N_9605,N_8300,N_8675);
or U9606 (N_9606,N_8578,N_8886);
nor U9607 (N_9607,N_8803,N_8919);
nor U9608 (N_9608,N_8309,N_8467);
nor U9609 (N_9609,N_8345,N_8761);
or U9610 (N_9610,N_8824,N_8510);
nor U9611 (N_9611,N_8710,N_8927);
or U9612 (N_9612,N_8632,N_8506);
nand U9613 (N_9613,N_8680,N_8672);
and U9614 (N_9614,N_8779,N_8324);
nand U9615 (N_9615,N_8785,N_8504);
nand U9616 (N_9616,N_8560,N_8604);
nor U9617 (N_9617,N_8319,N_8445);
or U9618 (N_9618,N_8865,N_8600);
and U9619 (N_9619,N_8293,N_8949);
nor U9620 (N_9620,N_8557,N_8558);
and U9621 (N_9621,N_8499,N_8981);
nand U9622 (N_9622,N_8736,N_8467);
nor U9623 (N_9623,N_8410,N_8383);
nor U9624 (N_9624,N_8897,N_8522);
nor U9625 (N_9625,N_8731,N_8835);
or U9626 (N_9626,N_8593,N_8351);
and U9627 (N_9627,N_8818,N_8827);
nor U9628 (N_9628,N_8948,N_8589);
nand U9629 (N_9629,N_8406,N_8329);
nand U9630 (N_9630,N_8309,N_8825);
nor U9631 (N_9631,N_8792,N_8396);
or U9632 (N_9632,N_8740,N_8916);
and U9633 (N_9633,N_8896,N_8685);
or U9634 (N_9634,N_8966,N_8277);
and U9635 (N_9635,N_8781,N_8435);
or U9636 (N_9636,N_8269,N_8714);
xnor U9637 (N_9637,N_8412,N_8882);
nand U9638 (N_9638,N_8990,N_8465);
and U9639 (N_9639,N_8770,N_8744);
nor U9640 (N_9640,N_8370,N_8710);
or U9641 (N_9641,N_8509,N_8718);
nor U9642 (N_9642,N_8492,N_8409);
and U9643 (N_9643,N_8743,N_8476);
or U9644 (N_9644,N_8983,N_8549);
or U9645 (N_9645,N_8279,N_8370);
nor U9646 (N_9646,N_8743,N_8316);
nand U9647 (N_9647,N_8908,N_8856);
xor U9648 (N_9648,N_8402,N_8414);
or U9649 (N_9649,N_8533,N_8884);
or U9650 (N_9650,N_8808,N_8750);
and U9651 (N_9651,N_8269,N_8524);
nor U9652 (N_9652,N_8624,N_8653);
nor U9653 (N_9653,N_8329,N_8829);
and U9654 (N_9654,N_8352,N_8356);
xor U9655 (N_9655,N_8471,N_8668);
nand U9656 (N_9656,N_8903,N_8648);
xnor U9657 (N_9657,N_8435,N_8762);
or U9658 (N_9658,N_8808,N_8328);
and U9659 (N_9659,N_8907,N_8340);
nand U9660 (N_9660,N_8612,N_8770);
nand U9661 (N_9661,N_8527,N_8379);
nand U9662 (N_9662,N_8312,N_8300);
nor U9663 (N_9663,N_8792,N_8891);
or U9664 (N_9664,N_8624,N_8826);
xor U9665 (N_9665,N_8432,N_8771);
nor U9666 (N_9666,N_8365,N_8611);
nand U9667 (N_9667,N_8999,N_8693);
nand U9668 (N_9668,N_8829,N_8263);
or U9669 (N_9669,N_8377,N_8647);
and U9670 (N_9670,N_8366,N_8927);
or U9671 (N_9671,N_8883,N_8353);
nor U9672 (N_9672,N_8800,N_8708);
nand U9673 (N_9673,N_8439,N_8792);
and U9674 (N_9674,N_8602,N_8535);
nor U9675 (N_9675,N_8917,N_8492);
nand U9676 (N_9676,N_8783,N_8340);
nor U9677 (N_9677,N_8584,N_8449);
nand U9678 (N_9678,N_8267,N_8762);
xnor U9679 (N_9679,N_8903,N_8557);
nor U9680 (N_9680,N_8996,N_8980);
and U9681 (N_9681,N_8690,N_8411);
nand U9682 (N_9682,N_8310,N_8633);
or U9683 (N_9683,N_8736,N_8654);
nand U9684 (N_9684,N_8360,N_8604);
or U9685 (N_9685,N_8675,N_8623);
nor U9686 (N_9686,N_8969,N_8519);
xnor U9687 (N_9687,N_8929,N_8500);
or U9688 (N_9688,N_8842,N_8600);
or U9689 (N_9689,N_8953,N_8683);
nand U9690 (N_9690,N_8989,N_8993);
or U9691 (N_9691,N_8311,N_8377);
or U9692 (N_9692,N_8325,N_8312);
or U9693 (N_9693,N_8781,N_8671);
nand U9694 (N_9694,N_8659,N_8971);
or U9695 (N_9695,N_8888,N_8476);
nor U9696 (N_9696,N_8549,N_8563);
or U9697 (N_9697,N_8318,N_8746);
nand U9698 (N_9698,N_8495,N_8993);
or U9699 (N_9699,N_8758,N_8377);
nor U9700 (N_9700,N_8286,N_8624);
and U9701 (N_9701,N_8705,N_8925);
nand U9702 (N_9702,N_8393,N_8374);
nand U9703 (N_9703,N_8432,N_8755);
xnor U9704 (N_9704,N_8453,N_8717);
nor U9705 (N_9705,N_8577,N_8353);
xnor U9706 (N_9706,N_8412,N_8601);
and U9707 (N_9707,N_8803,N_8643);
xor U9708 (N_9708,N_8293,N_8838);
xnor U9709 (N_9709,N_8281,N_8917);
and U9710 (N_9710,N_8259,N_8982);
and U9711 (N_9711,N_8522,N_8568);
xor U9712 (N_9712,N_8772,N_8290);
xor U9713 (N_9713,N_8589,N_8733);
and U9714 (N_9714,N_8855,N_8583);
nand U9715 (N_9715,N_8612,N_8580);
and U9716 (N_9716,N_8351,N_8418);
and U9717 (N_9717,N_8631,N_8969);
nor U9718 (N_9718,N_8540,N_8968);
nor U9719 (N_9719,N_8923,N_8752);
nor U9720 (N_9720,N_8429,N_8878);
nor U9721 (N_9721,N_8951,N_8567);
and U9722 (N_9722,N_8279,N_8522);
or U9723 (N_9723,N_8606,N_8301);
and U9724 (N_9724,N_8599,N_8305);
nand U9725 (N_9725,N_8768,N_8850);
or U9726 (N_9726,N_8581,N_8476);
nor U9727 (N_9727,N_8773,N_8302);
and U9728 (N_9728,N_8716,N_8326);
nand U9729 (N_9729,N_8509,N_8419);
xor U9730 (N_9730,N_8774,N_8480);
or U9731 (N_9731,N_8331,N_8684);
and U9732 (N_9732,N_8736,N_8942);
nand U9733 (N_9733,N_8361,N_8616);
nor U9734 (N_9734,N_8872,N_8344);
nor U9735 (N_9735,N_8847,N_8983);
xor U9736 (N_9736,N_8848,N_8973);
and U9737 (N_9737,N_8769,N_8391);
or U9738 (N_9738,N_8493,N_8388);
nor U9739 (N_9739,N_8878,N_8768);
and U9740 (N_9740,N_8647,N_8595);
nor U9741 (N_9741,N_8538,N_8409);
and U9742 (N_9742,N_8916,N_8994);
and U9743 (N_9743,N_8641,N_8444);
nor U9744 (N_9744,N_8823,N_8517);
nand U9745 (N_9745,N_8895,N_8525);
and U9746 (N_9746,N_8825,N_8793);
nor U9747 (N_9747,N_8918,N_8317);
or U9748 (N_9748,N_8996,N_8947);
or U9749 (N_9749,N_8647,N_8410);
and U9750 (N_9750,N_9427,N_9661);
or U9751 (N_9751,N_9469,N_9313);
nor U9752 (N_9752,N_9348,N_9139);
or U9753 (N_9753,N_9000,N_9172);
nor U9754 (N_9754,N_9578,N_9401);
and U9755 (N_9755,N_9691,N_9108);
or U9756 (N_9756,N_9366,N_9402);
and U9757 (N_9757,N_9193,N_9529);
xor U9758 (N_9758,N_9373,N_9555);
or U9759 (N_9759,N_9600,N_9018);
nor U9760 (N_9760,N_9695,N_9470);
nand U9761 (N_9761,N_9531,N_9296);
xor U9762 (N_9762,N_9560,N_9004);
nor U9763 (N_9763,N_9533,N_9293);
nor U9764 (N_9764,N_9449,N_9713);
nor U9765 (N_9765,N_9404,N_9039);
or U9766 (N_9766,N_9323,N_9011);
or U9767 (N_9767,N_9385,N_9336);
nor U9768 (N_9768,N_9071,N_9681);
and U9769 (N_9769,N_9213,N_9331);
xor U9770 (N_9770,N_9637,N_9181);
or U9771 (N_9771,N_9105,N_9477);
or U9772 (N_9772,N_9662,N_9430);
and U9773 (N_9773,N_9716,N_9437);
or U9774 (N_9774,N_9590,N_9475);
nor U9775 (N_9775,N_9307,N_9527);
nor U9776 (N_9776,N_9692,N_9092);
or U9777 (N_9777,N_9489,N_9727);
nor U9778 (N_9778,N_9288,N_9610);
xor U9779 (N_9779,N_9704,N_9142);
xnor U9780 (N_9780,N_9585,N_9122);
nand U9781 (N_9781,N_9270,N_9262);
or U9782 (N_9782,N_9002,N_9552);
and U9783 (N_9783,N_9619,N_9514);
nor U9784 (N_9784,N_9518,N_9110);
nor U9785 (N_9785,N_9079,N_9743);
and U9786 (N_9786,N_9542,N_9144);
or U9787 (N_9787,N_9370,N_9526);
nor U9788 (N_9788,N_9070,N_9241);
or U9789 (N_9789,N_9549,N_9553);
or U9790 (N_9790,N_9257,N_9403);
or U9791 (N_9791,N_9249,N_9033);
and U9792 (N_9792,N_9606,N_9685);
and U9793 (N_9793,N_9170,N_9633);
nor U9794 (N_9794,N_9146,N_9147);
or U9795 (N_9795,N_9157,N_9318);
or U9796 (N_9796,N_9672,N_9273);
nand U9797 (N_9797,N_9412,N_9048);
and U9798 (N_9798,N_9525,N_9705);
and U9799 (N_9799,N_9368,N_9644);
nand U9800 (N_9800,N_9279,N_9007);
or U9801 (N_9801,N_9722,N_9568);
xor U9802 (N_9802,N_9617,N_9179);
and U9803 (N_9803,N_9454,N_9145);
nor U9804 (N_9804,N_9614,N_9392);
and U9805 (N_9805,N_9010,N_9203);
or U9806 (N_9806,N_9452,N_9223);
nor U9807 (N_9807,N_9493,N_9180);
or U9808 (N_9808,N_9586,N_9584);
and U9809 (N_9809,N_9410,N_9636);
nor U9810 (N_9810,N_9503,N_9308);
nor U9811 (N_9811,N_9679,N_9053);
or U9812 (N_9812,N_9558,N_9740);
or U9813 (N_9813,N_9113,N_9730);
nand U9814 (N_9814,N_9624,N_9572);
nand U9815 (N_9815,N_9134,N_9258);
nand U9816 (N_9816,N_9453,N_9450);
nand U9817 (N_9817,N_9320,N_9457);
nor U9818 (N_9818,N_9745,N_9299);
nor U9819 (N_9819,N_9665,N_9564);
or U9820 (N_9820,N_9339,N_9428);
nor U9821 (N_9821,N_9546,N_9065);
and U9822 (N_9822,N_9066,N_9420);
xnor U9823 (N_9823,N_9265,N_9522);
nor U9824 (N_9824,N_9562,N_9710);
nor U9825 (N_9825,N_9579,N_9380);
and U9826 (N_9826,N_9358,N_9461);
and U9827 (N_9827,N_9153,N_9673);
nand U9828 (N_9828,N_9658,N_9400);
nand U9829 (N_9829,N_9720,N_9354);
xnor U9830 (N_9830,N_9379,N_9229);
and U9831 (N_9831,N_9398,N_9399);
nand U9832 (N_9832,N_9137,N_9741);
xnor U9833 (N_9833,N_9352,N_9311);
nor U9834 (N_9834,N_9228,N_9678);
xor U9835 (N_9835,N_9524,N_9280);
nor U9836 (N_9836,N_9292,N_9343);
nand U9837 (N_9837,N_9301,N_9587);
and U9838 (N_9838,N_9728,N_9523);
nor U9839 (N_9839,N_9576,N_9244);
and U9840 (N_9840,N_9473,N_9266);
nand U9841 (N_9841,N_9657,N_9029);
nand U9842 (N_9842,N_9310,N_9267);
xnor U9843 (N_9843,N_9084,N_9231);
nor U9844 (N_9844,N_9391,N_9544);
and U9845 (N_9845,N_9459,N_9729);
nand U9846 (N_9846,N_9715,N_9281);
nor U9847 (N_9847,N_9407,N_9719);
or U9848 (N_9848,N_9506,N_9441);
nand U9849 (N_9849,N_9243,N_9054);
and U9850 (N_9850,N_9599,N_9341);
or U9851 (N_9851,N_9442,N_9357);
or U9852 (N_9852,N_9748,N_9162);
xnor U9853 (N_9853,N_9375,N_9082);
or U9854 (N_9854,N_9736,N_9702);
or U9855 (N_9855,N_9364,N_9487);
or U9856 (N_9856,N_9471,N_9464);
xor U9857 (N_9857,N_9306,N_9565);
and U9858 (N_9858,N_9239,N_9643);
nand U9859 (N_9859,N_9090,N_9169);
xnor U9860 (N_9860,N_9235,N_9389);
nor U9861 (N_9861,N_9628,N_9448);
or U9862 (N_9862,N_9641,N_9264);
and U9863 (N_9863,N_9197,N_9294);
or U9864 (N_9864,N_9666,N_9012);
and U9865 (N_9865,N_9693,N_9220);
nand U9866 (N_9866,N_9663,N_9116);
nor U9867 (N_9867,N_9259,N_9688);
nand U9868 (N_9868,N_9612,N_9246);
xor U9869 (N_9869,N_9595,N_9278);
or U9870 (N_9870,N_9133,N_9256);
or U9871 (N_9871,N_9100,N_9653);
nor U9872 (N_9872,N_9683,N_9117);
nor U9873 (N_9873,N_9676,N_9156);
or U9874 (N_9874,N_9682,N_9515);
nand U9875 (N_9875,N_9342,N_9335);
nand U9876 (N_9876,N_9047,N_9019);
or U9877 (N_9877,N_9164,N_9630);
nor U9878 (N_9878,N_9508,N_9030);
nand U9879 (N_9879,N_9240,N_9739);
nor U9880 (N_9880,N_9645,N_9290);
and U9881 (N_9881,N_9186,N_9351);
nor U9882 (N_9882,N_9059,N_9201);
or U9883 (N_9883,N_9419,N_9096);
xnor U9884 (N_9884,N_9609,N_9232);
xor U9885 (N_9885,N_9397,N_9001);
nor U9886 (N_9886,N_9534,N_9058);
nand U9887 (N_9887,N_9488,N_9723);
and U9888 (N_9888,N_9214,N_9119);
xnor U9889 (N_9889,N_9605,N_9381);
or U9890 (N_9890,N_9126,N_9009);
nor U9891 (N_9891,N_9149,N_9492);
xnor U9892 (N_9892,N_9594,N_9087);
nor U9893 (N_9893,N_9634,N_9481);
nor U9894 (N_9894,N_9286,N_9543);
nand U9895 (N_9895,N_9659,N_9226);
nor U9896 (N_9896,N_9225,N_9349);
and U9897 (N_9897,N_9447,N_9639);
nor U9898 (N_9898,N_9414,N_9497);
or U9899 (N_9899,N_9569,N_9406);
nand U9900 (N_9900,N_9677,N_9625);
or U9901 (N_9901,N_9174,N_9490);
and U9902 (N_9902,N_9284,N_9629);
nand U9903 (N_9903,N_9106,N_9694);
nor U9904 (N_9904,N_9148,N_9509);
nand U9905 (N_9905,N_9275,N_9498);
nand U9906 (N_9906,N_9080,N_9405);
nand U9907 (N_9907,N_9216,N_9188);
nand U9908 (N_9908,N_9123,N_9615);
and U9909 (N_9909,N_9387,N_9178);
or U9910 (N_9910,N_9025,N_9104);
xnor U9911 (N_9911,N_9283,N_9417);
or U9912 (N_9912,N_9438,N_9218);
nand U9913 (N_9913,N_9334,N_9640);
nand U9914 (N_9914,N_9046,N_9698);
and U9915 (N_9915,N_9749,N_9020);
or U9916 (N_9916,N_9222,N_9230);
and U9917 (N_9917,N_9287,N_9177);
nor U9918 (N_9918,N_9697,N_9652);
nand U9919 (N_9919,N_9022,N_9217);
nand U9920 (N_9920,N_9486,N_9329);
or U9921 (N_9921,N_9035,N_9289);
nor U9922 (N_9922,N_9418,N_9344);
nand U9923 (N_9923,N_9424,N_9260);
nand U9924 (N_9924,N_9166,N_9725);
xnor U9925 (N_9925,N_9496,N_9227);
and U9926 (N_9926,N_9160,N_9253);
and U9927 (N_9927,N_9191,N_9250);
and U9928 (N_9928,N_9581,N_9456);
xnor U9929 (N_9929,N_9171,N_9300);
and U9930 (N_9930,N_9150,N_9502);
and U9931 (N_9931,N_9604,N_9127);
nand U9932 (N_9932,N_9717,N_9194);
and U9933 (N_9933,N_9107,N_9056);
or U9934 (N_9934,N_9049,N_9130);
xnor U9935 (N_9935,N_9315,N_9583);
and U9936 (N_9936,N_9532,N_9413);
nor U9937 (N_9937,N_9362,N_9034);
nor U9938 (N_9938,N_9537,N_9591);
or U9939 (N_9939,N_9045,N_9394);
or U9940 (N_9940,N_9460,N_9069);
and U9941 (N_9941,N_9638,N_9173);
or U9942 (N_9942,N_9043,N_9089);
or U9943 (N_9943,N_9507,N_9738);
and U9944 (N_9944,N_9541,N_9669);
nand U9945 (N_9945,N_9480,N_9557);
nand U9946 (N_9946,N_9667,N_9062);
nor U9947 (N_9947,N_9131,N_9545);
nand U9948 (N_9948,N_9501,N_9718);
nor U9949 (N_9949,N_9233,N_9482);
nor U9950 (N_9950,N_9369,N_9512);
nor U9951 (N_9951,N_9073,N_9535);
or U9952 (N_9952,N_9621,N_9094);
xnor U9953 (N_9953,N_9211,N_9689);
nor U9954 (N_9954,N_9176,N_9550);
nor U9955 (N_9955,N_9703,N_9361);
and U9956 (N_9956,N_9302,N_9592);
xor U9957 (N_9957,N_9124,N_9714);
xor U9958 (N_9958,N_9712,N_9350);
nand U9959 (N_9959,N_9234,N_9395);
and U9960 (N_9960,N_9003,N_9209);
or U9961 (N_9961,N_9282,N_9309);
or U9962 (N_9962,N_9478,N_9190);
nor U9963 (N_9963,N_9731,N_9408);
xor U9964 (N_9964,N_9014,N_9024);
nor U9965 (N_9965,N_9013,N_9451);
xnor U9966 (N_9966,N_9242,N_9642);
or U9967 (N_9967,N_9224,N_9626);
and U9968 (N_9968,N_9031,N_9271);
nand U9969 (N_9969,N_9330,N_9660);
nor U9970 (N_9970,N_9304,N_9155);
nand U9971 (N_9971,N_9429,N_9206);
nor U9972 (N_9972,N_9023,N_9063);
nor U9973 (N_9973,N_9026,N_9050);
or U9974 (N_9974,N_9015,N_9589);
nand U9975 (N_9975,N_9163,N_9483);
nand U9976 (N_9976,N_9363,N_9648);
or U9977 (N_9977,N_9340,N_9434);
nand U9978 (N_9978,N_9319,N_9747);
and U9979 (N_9979,N_9091,N_9511);
xnor U9980 (N_9980,N_9680,N_9516);
and U9981 (N_9981,N_9588,N_9409);
xor U9982 (N_9982,N_9548,N_9654);
nor U9983 (N_9983,N_9620,N_9247);
and U9984 (N_9984,N_9044,N_9382);
nand U9985 (N_9985,N_9495,N_9316);
nor U9986 (N_9986,N_9466,N_9517);
nand U9987 (N_9987,N_9165,N_9251);
nand U9988 (N_9988,N_9706,N_9083);
and U9989 (N_9989,N_9566,N_9603);
nand U9990 (N_9990,N_9465,N_9601);
and U9991 (N_9991,N_9112,N_9699);
nor U9992 (N_9992,N_9102,N_9237);
nor U9993 (N_9993,N_9154,N_9462);
nor U9994 (N_9994,N_9274,N_9199);
and U9995 (N_9995,N_9198,N_9221);
and U9996 (N_9996,N_9151,N_9109);
xnor U9997 (N_9997,N_9425,N_9491);
and U9998 (N_9998,N_9443,N_9494);
nor U9999 (N_9999,N_9118,N_9690);
nor U10000 (N_10000,N_9285,N_9005);
nand U10001 (N_10001,N_9093,N_9081);
xnor U10002 (N_10002,N_9378,N_9184);
nor U10003 (N_10003,N_9128,N_9359);
xnor U10004 (N_10004,N_9333,N_9554);
nor U10005 (N_10005,N_9205,N_9575);
and U10006 (N_10006,N_9426,N_9167);
nand U10007 (N_10007,N_9159,N_9248);
and U10008 (N_10008,N_9036,N_9530);
and U10009 (N_10009,N_9536,N_9076);
nand U10010 (N_10010,N_9563,N_9458);
or U10011 (N_10011,N_9120,N_9067);
nand U10012 (N_10012,N_9708,N_9303);
xor U10013 (N_10013,N_9721,N_9028);
and U10014 (N_10014,N_9686,N_9115);
nand U10015 (N_10015,N_9061,N_9185);
or U10016 (N_10016,N_9152,N_9655);
and U10017 (N_10017,N_9709,N_9746);
nand U10018 (N_10018,N_9269,N_9041);
nand U10019 (N_10019,N_9650,N_9103);
nand U10020 (N_10020,N_9161,N_9396);
nand U10021 (N_10021,N_9440,N_9295);
and U10022 (N_10022,N_9390,N_9631);
nand U10023 (N_10023,N_9276,N_9700);
or U10024 (N_10024,N_9136,N_9618);
nand U10025 (N_10025,N_9416,N_9353);
nand U10026 (N_10026,N_9016,N_9519);
nand U10027 (N_10027,N_9168,N_9101);
nand U10028 (N_10028,N_9421,N_9360);
nor U10029 (N_10029,N_9332,N_9141);
or U10030 (N_10030,N_9060,N_9182);
nor U10031 (N_10031,N_9632,N_9476);
nand U10032 (N_10032,N_9125,N_9696);
and U10033 (N_10033,N_9272,N_9098);
xor U10034 (N_10034,N_9038,N_9707);
nand U10035 (N_10035,N_9338,N_9593);
nor U10036 (N_10036,N_9074,N_9263);
nand U10037 (N_10037,N_9613,N_9189);
nor U10038 (N_10038,N_9345,N_9551);
nor U10039 (N_10039,N_9439,N_9021);
nand U10040 (N_10040,N_9472,N_9192);
nand U10041 (N_10041,N_9322,N_9556);
and U10042 (N_10042,N_9355,N_9737);
and U10043 (N_10043,N_9732,N_9187);
and U10044 (N_10044,N_9305,N_9611);
nor U10045 (N_10045,N_9602,N_9510);
or U10046 (N_10046,N_9734,N_9479);
xor U10047 (N_10047,N_9726,N_9422);
and U10048 (N_10048,N_9356,N_9337);
xnor U10049 (N_10049,N_9393,N_9196);
or U10050 (N_10050,N_9647,N_9255);
nor U10051 (N_10051,N_9540,N_9468);
nor U10052 (N_10052,N_9383,N_9183);
and U10053 (N_10053,N_9671,N_9236);
nor U10054 (N_10054,N_9596,N_9365);
nor U10055 (N_10055,N_9377,N_9651);
and U10056 (N_10056,N_9622,N_9347);
xor U10057 (N_10057,N_9254,N_9277);
or U10058 (N_10058,N_9656,N_9684);
nand U10059 (N_10059,N_9432,N_9055);
and U10060 (N_10060,N_9135,N_9500);
nor U10061 (N_10061,N_9724,N_9032);
and U10062 (N_10062,N_9068,N_9121);
or U10063 (N_10063,N_9064,N_9607);
nor U10064 (N_10064,N_9075,N_9571);
nor U10065 (N_10065,N_9111,N_9561);
or U10066 (N_10066,N_9623,N_9085);
or U10067 (N_10067,N_9314,N_9268);
xnor U10068 (N_10068,N_9436,N_9095);
nand U10069 (N_10069,N_9674,N_9312);
or U10070 (N_10070,N_9415,N_9325);
nor U10071 (N_10071,N_9735,N_9504);
or U10072 (N_10072,N_9321,N_9327);
nand U10073 (N_10073,N_9520,N_9467);
and U10074 (N_10074,N_9646,N_9212);
and U10075 (N_10075,N_9097,N_9372);
or U10076 (N_10076,N_9298,N_9474);
or U10077 (N_10077,N_9077,N_9573);
and U10078 (N_10078,N_9687,N_9582);
nor U10079 (N_10079,N_9143,N_9616);
and U10080 (N_10080,N_9324,N_9559);
and U10081 (N_10081,N_9042,N_9388);
nand U10082 (N_10082,N_9202,N_9513);
or U10083 (N_10083,N_9326,N_9574);
nand U10084 (N_10084,N_9598,N_9297);
or U10085 (N_10085,N_9132,N_9200);
nand U10086 (N_10086,N_9078,N_9742);
or U10087 (N_10087,N_9210,N_9175);
or U10088 (N_10088,N_9037,N_9208);
or U10089 (N_10089,N_9328,N_9423);
nor U10090 (N_10090,N_9580,N_9446);
and U10091 (N_10091,N_9649,N_9670);
nor U10092 (N_10092,N_9367,N_9521);
and U10093 (N_10093,N_9431,N_9701);
or U10094 (N_10094,N_9017,N_9261);
or U10095 (N_10095,N_9057,N_9346);
nor U10096 (N_10096,N_9138,N_9140);
nor U10097 (N_10097,N_9499,N_9744);
or U10098 (N_10098,N_9088,N_9051);
or U10099 (N_10099,N_9114,N_9445);
and U10100 (N_10100,N_9219,N_9635);
xor U10101 (N_10101,N_9570,N_9384);
or U10102 (N_10102,N_9733,N_9376);
and U10103 (N_10103,N_9252,N_9245);
and U10104 (N_10104,N_9538,N_9040);
xor U10105 (N_10105,N_9528,N_9158);
nor U10106 (N_10106,N_9052,N_9072);
nand U10107 (N_10107,N_9597,N_9577);
nor U10108 (N_10108,N_9608,N_9547);
nand U10109 (N_10109,N_9668,N_9433);
xnor U10110 (N_10110,N_9711,N_9567);
and U10111 (N_10111,N_9291,N_9371);
and U10112 (N_10112,N_9664,N_9485);
nor U10113 (N_10113,N_9675,N_9129);
or U10114 (N_10114,N_9317,N_9411);
and U10115 (N_10115,N_9215,N_9008);
nor U10116 (N_10116,N_9455,N_9539);
and U10117 (N_10117,N_9006,N_9207);
or U10118 (N_10118,N_9435,N_9505);
and U10119 (N_10119,N_9027,N_9204);
nor U10120 (N_10120,N_9099,N_9374);
or U10121 (N_10121,N_9484,N_9463);
and U10122 (N_10122,N_9086,N_9238);
and U10123 (N_10123,N_9195,N_9386);
and U10124 (N_10124,N_9444,N_9627);
nor U10125 (N_10125,N_9150,N_9241);
xnor U10126 (N_10126,N_9195,N_9510);
and U10127 (N_10127,N_9235,N_9627);
and U10128 (N_10128,N_9036,N_9263);
nand U10129 (N_10129,N_9202,N_9535);
and U10130 (N_10130,N_9214,N_9060);
and U10131 (N_10131,N_9021,N_9015);
nor U10132 (N_10132,N_9663,N_9353);
nand U10133 (N_10133,N_9231,N_9644);
and U10134 (N_10134,N_9253,N_9629);
nor U10135 (N_10135,N_9139,N_9574);
or U10136 (N_10136,N_9604,N_9704);
or U10137 (N_10137,N_9727,N_9228);
nand U10138 (N_10138,N_9149,N_9442);
nand U10139 (N_10139,N_9448,N_9011);
nor U10140 (N_10140,N_9314,N_9537);
xnor U10141 (N_10141,N_9207,N_9092);
nor U10142 (N_10142,N_9642,N_9310);
and U10143 (N_10143,N_9413,N_9013);
nand U10144 (N_10144,N_9321,N_9427);
xor U10145 (N_10145,N_9267,N_9416);
and U10146 (N_10146,N_9572,N_9400);
nand U10147 (N_10147,N_9296,N_9334);
nor U10148 (N_10148,N_9336,N_9432);
or U10149 (N_10149,N_9058,N_9323);
nor U10150 (N_10150,N_9585,N_9642);
nor U10151 (N_10151,N_9148,N_9725);
nand U10152 (N_10152,N_9140,N_9182);
and U10153 (N_10153,N_9172,N_9218);
nand U10154 (N_10154,N_9697,N_9524);
nand U10155 (N_10155,N_9096,N_9522);
nand U10156 (N_10156,N_9432,N_9389);
nor U10157 (N_10157,N_9226,N_9540);
nand U10158 (N_10158,N_9494,N_9621);
or U10159 (N_10159,N_9340,N_9717);
or U10160 (N_10160,N_9209,N_9728);
nand U10161 (N_10161,N_9231,N_9555);
xnor U10162 (N_10162,N_9681,N_9558);
nor U10163 (N_10163,N_9339,N_9542);
nand U10164 (N_10164,N_9379,N_9476);
nor U10165 (N_10165,N_9039,N_9036);
or U10166 (N_10166,N_9227,N_9702);
and U10167 (N_10167,N_9352,N_9545);
xnor U10168 (N_10168,N_9329,N_9663);
and U10169 (N_10169,N_9337,N_9454);
nor U10170 (N_10170,N_9248,N_9040);
or U10171 (N_10171,N_9316,N_9494);
or U10172 (N_10172,N_9226,N_9078);
or U10173 (N_10173,N_9578,N_9309);
xor U10174 (N_10174,N_9540,N_9104);
xor U10175 (N_10175,N_9566,N_9572);
nand U10176 (N_10176,N_9026,N_9672);
xor U10177 (N_10177,N_9024,N_9018);
and U10178 (N_10178,N_9676,N_9511);
nor U10179 (N_10179,N_9678,N_9376);
and U10180 (N_10180,N_9475,N_9196);
nand U10181 (N_10181,N_9612,N_9400);
nand U10182 (N_10182,N_9343,N_9539);
nor U10183 (N_10183,N_9585,N_9745);
nand U10184 (N_10184,N_9589,N_9033);
or U10185 (N_10185,N_9230,N_9169);
nand U10186 (N_10186,N_9365,N_9676);
and U10187 (N_10187,N_9062,N_9277);
xnor U10188 (N_10188,N_9318,N_9111);
and U10189 (N_10189,N_9528,N_9097);
nand U10190 (N_10190,N_9211,N_9132);
nand U10191 (N_10191,N_9736,N_9344);
or U10192 (N_10192,N_9612,N_9592);
or U10193 (N_10193,N_9558,N_9409);
nand U10194 (N_10194,N_9454,N_9516);
xnor U10195 (N_10195,N_9578,N_9533);
nor U10196 (N_10196,N_9236,N_9204);
nor U10197 (N_10197,N_9667,N_9158);
nor U10198 (N_10198,N_9285,N_9422);
and U10199 (N_10199,N_9520,N_9240);
nand U10200 (N_10200,N_9471,N_9642);
nand U10201 (N_10201,N_9559,N_9179);
and U10202 (N_10202,N_9104,N_9389);
nand U10203 (N_10203,N_9247,N_9545);
xnor U10204 (N_10204,N_9031,N_9284);
nor U10205 (N_10205,N_9198,N_9328);
nor U10206 (N_10206,N_9041,N_9510);
nand U10207 (N_10207,N_9603,N_9538);
nor U10208 (N_10208,N_9630,N_9429);
nand U10209 (N_10209,N_9574,N_9167);
and U10210 (N_10210,N_9748,N_9605);
nor U10211 (N_10211,N_9733,N_9326);
and U10212 (N_10212,N_9700,N_9619);
and U10213 (N_10213,N_9487,N_9547);
nor U10214 (N_10214,N_9049,N_9218);
nand U10215 (N_10215,N_9423,N_9300);
or U10216 (N_10216,N_9547,N_9158);
and U10217 (N_10217,N_9011,N_9467);
nor U10218 (N_10218,N_9165,N_9355);
or U10219 (N_10219,N_9634,N_9496);
xnor U10220 (N_10220,N_9710,N_9157);
or U10221 (N_10221,N_9063,N_9499);
and U10222 (N_10222,N_9394,N_9355);
nor U10223 (N_10223,N_9510,N_9349);
or U10224 (N_10224,N_9503,N_9249);
and U10225 (N_10225,N_9101,N_9098);
nand U10226 (N_10226,N_9741,N_9215);
nor U10227 (N_10227,N_9069,N_9356);
nor U10228 (N_10228,N_9696,N_9063);
and U10229 (N_10229,N_9098,N_9463);
nand U10230 (N_10230,N_9288,N_9484);
xnor U10231 (N_10231,N_9422,N_9029);
xor U10232 (N_10232,N_9448,N_9589);
and U10233 (N_10233,N_9041,N_9121);
nor U10234 (N_10234,N_9466,N_9518);
nand U10235 (N_10235,N_9330,N_9580);
and U10236 (N_10236,N_9495,N_9480);
nand U10237 (N_10237,N_9132,N_9597);
or U10238 (N_10238,N_9739,N_9052);
xnor U10239 (N_10239,N_9335,N_9403);
or U10240 (N_10240,N_9172,N_9337);
and U10241 (N_10241,N_9659,N_9649);
nor U10242 (N_10242,N_9494,N_9349);
and U10243 (N_10243,N_9056,N_9297);
or U10244 (N_10244,N_9482,N_9445);
nand U10245 (N_10245,N_9026,N_9351);
nor U10246 (N_10246,N_9605,N_9637);
and U10247 (N_10247,N_9468,N_9472);
nand U10248 (N_10248,N_9410,N_9147);
nand U10249 (N_10249,N_9091,N_9303);
or U10250 (N_10250,N_9121,N_9335);
nor U10251 (N_10251,N_9356,N_9360);
nand U10252 (N_10252,N_9477,N_9466);
nand U10253 (N_10253,N_9440,N_9524);
nand U10254 (N_10254,N_9662,N_9107);
nand U10255 (N_10255,N_9710,N_9326);
and U10256 (N_10256,N_9249,N_9065);
nor U10257 (N_10257,N_9217,N_9567);
and U10258 (N_10258,N_9520,N_9431);
and U10259 (N_10259,N_9002,N_9366);
or U10260 (N_10260,N_9291,N_9397);
and U10261 (N_10261,N_9185,N_9311);
xnor U10262 (N_10262,N_9687,N_9131);
and U10263 (N_10263,N_9710,N_9586);
and U10264 (N_10264,N_9588,N_9343);
nand U10265 (N_10265,N_9018,N_9142);
or U10266 (N_10266,N_9269,N_9039);
nand U10267 (N_10267,N_9512,N_9622);
nor U10268 (N_10268,N_9425,N_9317);
and U10269 (N_10269,N_9145,N_9249);
nand U10270 (N_10270,N_9024,N_9609);
and U10271 (N_10271,N_9551,N_9433);
and U10272 (N_10272,N_9094,N_9220);
xor U10273 (N_10273,N_9194,N_9367);
xnor U10274 (N_10274,N_9211,N_9266);
nor U10275 (N_10275,N_9329,N_9414);
nor U10276 (N_10276,N_9311,N_9161);
and U10277 (N_10277,N_9584,N_9616);
nand U10278 (N_10278,N_9143,N_9408);
and U10279 (N_10279,N_9444,N_9018);
or U10280 (N_10280,N_9450,N_9055);
xnor U10281 (N_10281,N_9536,N_9264);
nor U10282 (N_10282,N_9248,N_9654);
nand U10283 (N_10283,N_9745,N_9133);
and U10284 (N_10284,N_9573,N_9447);
or U10285 (N_10285,N_9639,N_9025);
or U10286 (N_10286,N_9648,N_9376);
xor U10287 (N_10287,N_9389,N_9631);
nand U10288 (N_10288,N_9481,N_9534);
xnor U10289 (N_10289,N_9045,N_9105);
nor U10290 (N_10290,N_9479,N_9371);
and U10291 (N_10291,N_9023,N_9499);
nor U10292 (N_10292,N_9695,N_9542);
nor U10293 (N_10293,N_9364,N_9507);
or U10294 (N_10294,N_9057,N_9637);
nand U10295 (N_10295,N_9124,N_9580);
or U10296 (N_10296,N_9441,N_9091);
xnor U10297 (N_10297,N_9221,N_9705);
nand U10298 (N_10298,N_9100,N_9647);
nor U10299 (N_10299,N_9419,N_9012);
or U10300 (N_10300,N_9057,N_9409);
nand U10301 (N_10301,N_9593,N_9330);
xnor U10302 (N_10302,N_9116,N_9382);
nor U10303 (N_10303,N_9069,N_9355);
nor U10304 (N_10304,N_9073,N_9724);
and U10305 (N_10305,N_9644,N_9602);
xnor U10306 (N_10306,N_9584,N_9141);
and U10307 (N_10307,N_9506,N_9251);
or U10308 (N_10308,N_9695,N_9498);
xnor U10309 (N_10309,N_9069,N_9024);
and U10310 (N_10310,N_9412,N_9326);
nand U10311 (N_10311,N_9611,N_9298);
nand U10312 (N_10312,N_9728,N_9215);
and U10313 (N_10313,N_9603,N_9667);
or U10314 (N_10314,N_9397,N_9241);
nand U10315 (N_10315,N_9466,N_9627);
or U10316 (N_10316,N_9340,N_9192);
xor U10317 (N_10317,N_9164,N_9588);
nor U10318 (N_10318,N_9526,N_9531);
and U10319 (N_10319,N_9642,N_9425);
nor U10320 (N_10320,N_9141,N_9616);
nor U10321 (N_10321,N_9743,N_9654);
and U10322 (N_10322,N_9607,N_9042);
xor U10323 (N_10323,N_9381,N_9488);
or U10324 (N_10324,N_9413,N_9255);
nor U10325 (N_10325,N_9626,N_9312);
and U10326 (N_10326,N_9442,N_9331);
nor U10327 (N_10327,N_9335,N_9402);
nor U10328 (N_10328,N_9024,N_9335);
or U10329 (N_10329,N_9155,N_9406);
and U10330 (N_10330,N_9085,N_9408);
nand U10331 (N_10331,N_9086,N_9385);
and U10332 (N_10332,N_9748,N_9045);
and U10333 (N_10333,N_9069,N_9092);
and U10334 (N_10334,N_9524,N_9516);
nand U10335 (N_10335,N_9557,N_9723);
nor U10336 (N_10336,N_9006,N_9290);
nand U10337 (N_10337,N_9386,N_9227);
nor U10338 (N_10338,N_9165,N_9613);
nand U10339 (N_10339,N_9482,N_9084);
nand U10340 (N_10340,N_9307,N_9552);
nand U10341 (N_10341,N_9533,N_9374);
nand U10342 (N_10342,N_9709,N_9576);
nand U10343 (N_10343,N_9622,N_9054);
nand U10344 (N_10344,N_9227,N_9239);
and U10345 (N_10345,N_9590,N_9435);
nor U10346 (N_10346,N_9578,N_9300);
or U10347 (N_10347,N_9202,N_9707);
and U10348 (N_10348,N_9544,N_9128);
nor U10349 (N_10349,N_9647,N_9297);
and U10350 (N_10350,N_9703,N_9663);
and U10351 (N_10351,N_9027,N_9211);
and U10352 (N_10352,N_9508,N_9662);
nor U10353 (N_10353,N_9383,N_9701);
and U10354 (N_10354,N_9066,N_9418);
or U10355 (N_10355,N_9446,N_9545);
xor U10356 (N_10356,N_9424,N_9382);
and U10357 (N_10357,N_9144,N_9290);
nor U10358 (N_10358,N_9634,N_9139);
xor U10359 (N_10359,N_9346,N_9331);
and U10360 (N_10360,N_9326,N_9148);
and U10361 (N_10361,N_9674,N_9284);
or U10362 (N_10362,N_9565,N_9272);
nand U10363 (N_10363,N_9461,N_9477);
and U10364 (N_10364,N_9419,N_9661);
nand U10365 (N_10365,N_9672,N_9034);
nand U10366 (N_10366,N_9214,N_9256);
nand U10367 (N_10367,N_9026,N_9293);
nand U10368 (N_10368,N_9382,N_9611);
and U10369 (N_10369,N_9507,N_9485);
nor U10370 (N_10370,N_9505,N_9462);
nand U10371 (N_10371,N_9278,N_9677);
nand U10372 (N_10372,N_9745,N_9714);
or U10373 (N_10373,N_9561,N_9485);
and U10374 (N_10374,N_9722,N_9519);
nand U10375 (N_10375,N_9169,N_9149);
xor U10376 (N_10376,N_9274,N_9574);
nand U10377 (N_10377,N_9098,N_9721);
and U10378 (N_10378,N_9295,N_9444);
or U10379 (N_10379,N_9211,N_9301);
nand U10380 (N_10380,N_9739,N_9038);
nor U10381 (N_10381,N_9556,N_9459);
xor U10382 (N_10382,N_9328,N_9152);
nand U10383 (N_10383,N_9426,N_9595);
or U10384 (N_10384,N_9338,N_9075);
nor U10385 (N_10385,N_9040,N_9259);
or U10386 (N_10386,N_9322,N_9734);
and U10387 (N_10387,N_9108,N_9565);
or U10388 (N_10388,N_9713,N_9101);
or U10389 (N_10389,N_9648,N_9143);
nor U10390 (N_10390,N_9462,N_9106);
nand U10391 (N_10391,N_9257,N_9568);
and U10392 (N_10392,N_9447,N_9058);
xnor U10393 (N_10393,N_9407,N_9554);
nand U10394 (N_10394,N_9559,N_9286);
and U10395 (N_10395,N_9542,N_9406);
nor U10396 (N_10396,N_9641,N_9493);
nand U10397 (N_10397,N_9019,N_9089);
or U10398 (N_10398,N_9415,N_9095);
and U10399 (N_10399,N_9390,N_9374);
or U10400 (N_10400,N_9326,N_9517);
or U10401 (N_10401,N_9145,N_9261);
or U10402 (N_10402,N_9511,N_9631);
or U10403 (N_10403,N_9724,N_9175);
nor U10404 (N_10404,N_9226,N_9165);
nor U10405 (N_10405,N_9291,N_9055);
or U10406 (N_10406,N_9189,N_9530);
and U10407 (N_10407,N_9546,N_9141);
nand U10408 (N_10408,N_9099,N_9394);
and U10409 (N_10409,N_9572,N_9583);
nor U10410 (N_10410,N_9408,N_9529);
nand U10411 (N_10411,N_9577,N_9203);
nor U10412 (N_10412,N_9485,N_9569);
xnor U10413 (N_10413,N_9671,N_9679);
and U10414 (N_10414,N_9082,N_9177);
nand U10415 (N_10415,N_9559,N_9588);
nand U10416 (N_10416,N_9324,N_9690);
and U10417 (N_10417,N_9497,N_9222);
or U10418 (N_10418,N_9562,N_9480);
or U10419 (N_10419,N_9531,N_9393);
nand U10420 (N_10420,N_9380,N_9426);
and U10421 (N_10421,N_9019,N_9158);
nand U10422 (N_10422,N_9428,N_9417);
or U10423 (N_10423,N_9238,N_9330);
or U10424 (N_10424,N_9348,N_9725);
or U10425 (N_10425,N_9422,N_9352);
and U10426 (N_10426,N_9340,N_9255);
nor U10427 (N_10427,N_9099,N_9599);
and U10428 (N_10428,N_9059,N_9003);
nand U10429 (N_10429,N_9503,N_9238);
or U10430 (N_10430,N_9293,N_9671);
nor U10431 (N_10431,N_9102,N_9723);
nor U10432 (N_10432,N_9638,N_9424);
and U10433 (N_10433,N_9191,N_9557);
nand U10434 (N_10434,N_9518,N_9477);
and U10435 (N_10435,N_9549,N_9514);
and U10436 (N_10436,N_9623,N_9474);
nor U10437 (N_10437,N_9647,N_9011);
and U10438 (N_10438,N_9481,N_9485);
or U10439 (N_10439,N_9477,N_9451);
or U10440 (N_10440,N_9709,N_9241);
nor U10441 (N_10441,N_9312,N_9060);
or U10442 (N_10442,N_9465,N_9433);
nand U10443 (N_10443,N_9384,N_9478);
nor U10444 (N_10444,N_9109,N_9635);
nor U10445 (N_10445,N_9699,N_9093);
nand U10446 (N_10446,N_9603,N_9745);
or U10447 (N_10447,N_9096,N_9710);
and U10448 (N_10448,N_9268,N_9035);
nand U10449 (N_10449,N_9239,N_9269);
xnor U10450 (N_10450,N_9172,N_9394);
nor U10451 (N_10451,N_9581,N_9105);
nand U10452 (N_10452,N_9675,N_9257);
nor U10453 (N_10453,N_9459,N_9228);
or U10454 (N_10454,N_9323,N_9605);
and U10455 (N_10455,N_9626,N_9373);
or U10456 (N_10456,N_9459,N_9221);
nand U10457 (N_10457,N_9564,N_9316);
and U10458 (N_10458,N_9492,N_9520);
and U10459 (N_10459,N_9210,N_9115);
nor U10460 (N_10460,N_9262,N_9397);
and U10461 (N_10461,N_9188,N_9403);
nor U10462 (N_10462,N_9019,N_9132);
or U10463 (N_10463,N_9306,N_9025);
and U10464 (N_10464,N_9243,N_9118);
nand U10465 (N_10465,N_9388,N_9237);
nor U10466 (N_10466,N_9252,N_9450);
or U10467 (N_10467,N_9695,N_9244);
and U10468 (N_10468,N_9117,N_9615);
nor U10469 (N_10469,N_9468,N_9682);
xnor U10470 (N_10470,N_9254,N_9553);
nand U10471 (N_10471,N_9674,N_9111);
nor U10472 (N_10472,N_9275,N_9732);
xor U10473 (N_10473,N_9277,N_9221);
nor U10474 (N_10474,N_9628,N_9461);
and U10475 (N_10475,N_9198,N_9461);
and U10476 (N_10476,N_9297,N_9587);
and U10477 (N_10477,N_9526,N_9573);
or U10478 (N_10478,N_9595,N_9378);
nand U10479 (N_10479,N_9614,N_9165);
or U10480 (N_10480,N_9013,N_9609);
and U10481 (N_10481,N_9550,N_9436);
nand U10482 (N_10482,N_9369,N_9695);
nand U10483 (N_10483,N_9115,N_9110);
and U10484 (N_10484,N_9572,N_9506);
nor U10485 (N_10485,N_9538,N_9726);
nor U10486 (N_10486,N_9215,N_9209);
nand U10487 (N_10487,N_9383,N_9429);
xor U10488 (N_10488,N_9539,N_9500);
and U10489 (N_10489,N_9139,N_9181);
nand U10490 (N_10490,N_9395,N_9563);
and U10491 (N_10491,N_9012,N_9613);
nand U10492 (N_10492,N_9314,N_9072);
nand U10493 (N_10493,N_9135,N_9120);
or U10494 (N_10494,N_9173,N_9627);
and U10495 (N_10495,N_9557,N_9057);
nand U10496 (N_10496,N_9278,N_9181);
or U10497 (N_10497,N_9449,N_9310);
nor U10498 (N_10498,N_9611,N_9381);
and U10499 (N_10499,N_9405,N_9583);
and U10500 (N_10500,N_9907,N_9775);
or U10501 (N_10501,N_10425,N_10118);
nor U10502 (N_10502,N_10103,N_9946);
nand U10503 (N_10503,N_10081,N_10332);
and U10504 (N_10504,N_10001,N_10349);
xnor U10505 (N_10505,N_10056,N_10069);
or U10506 (N_10506,N_10356,N_10419);
or U10507 (N_10507,N_9931,N_10057);
or U10508 (N_10508,N_10386,N_9882);
nand U10509 (N_10509,N_9761,N_10454);
and U10510 (N_10510,N_10208,N_9956);
or U10511 (N_10511,N_9861,N_10113);
nor U10512 (N_10512,N_10443,N_9800);
and U10513 (N_10513,N_9763,N_9881);
and U10514 (N_10514,N_9901,N_10011);
and U10515 (N_10515,N_10231,N_10275);
nand U10516 (N_10516,N_9754,N_9913);
nor U10517 (N_10517,N_10068,N_10211);
nor U10518 (N_10518,N_10437,N_10064);
nor U10519 (N_10519,N_10390,N_10105);
or U10520 (N_10520,N_9985,N_9834);
and U10521 (N_10521,N_10247,N_9828);
and U10522 (N_10522,N_10201,N_10190);
nor U10523 (N_10523,N_10092,N_10097);
or U10524 (N_10524,N_10300,N_10492);
nand U10525 (N_10525,N_10235,N_10071);
xnor U10526 (N_10526,N_9918,N_10304);
and U10527 (N_10527,N_9768,N_9900);
nor U10528 (N_10528,N_10246,N_10418);
and U10529 (N_10529,N_9887,N_10311);
nor U10530 (N_10530,N_10164,N_9787);
nand U10531 (N_10531,N_10217,N_10104);
or U10532 (N_10532,N_10416,N_9976);
nor U10533 (N_10533,N_10361,N_10421);
nor U10534 (N_10534,N_10041,N_10233);
or U10535 (N_10535,N_10370,N_10373);
nor U10536 (N_10536,N_10471,N_9904);
xnor U10537 (N_10537,N_10396,N_10176);
or U10538 (N_10538,N_10261,N_10030);
or U10539 (N_10539,N_10406,N_10274);
or U10540 (N_10540,N_10009,N_10456);
nor U10541 (N_10541,N_9826,N_10444);
nand U10542 (N_10542,N_10021,N_9999);
or U10543 (N_10543,N_10474,N_9806);
nand U10544 (N_10544,N_9893,N_10120);
and U10545 (N_10545,N_9879,N_9943);
or U10546 (N_10546,N_9850,N_10210);
and U10547 (N_10547,N_10207,N_9909);
and U10548 (N_10548,N_10273,N_10499);
nand U10549 (N_10549,N_9797,N_10015);
nand U10550 (N_10550,N_9932,N_9903);
or U10551 (N_10551,N_10445,N_10496);
and U10552 (N_10552,N_10381,N_9849);
nand U10553 (N_10553,N_10293,N_10144);
nand U10554 (N_10554,N_9812,N_10163);
or U10555 (N_10555,N_10412,N_10091);
nor U10556 (N_10556,N_10366,N_10408);
nand U10557 (N_10557,N_9770,N_10153);
nor U10558 (N_10558,N_9854,N_10331);
and U10559 (N_10559,N_9944,N_9979);
or U10560 (N_10560,N_10379,N_10225);
or U10561 (N_10561,N_10491,N_9824);
xor U10562 (N_10562,N_10321,N_10382);
and U10563 (N_10563,N_10214,N_10158);
or U10564 (N_10564,N_10199,N_9786);
and U10565 (N_10565,N_10435,N_9841);
nor U10566 (N_10566,N_10295,N_10348);
nor U10567 (N_10567,N_10297,N_10162);
nor U10568 (N_10568,N_9859,N_10289);
or U10569 (N_10569,N_9928,N_9912);
and U10570 (N_10570,N_10268,N_9872);
nor U10571 (N_10571,N_10050,N_10218);
nor U10572 (N_10572,N_10060,N_9891);
or U10573 (N_10573,N_10291,N_10065);
nand U10574 (N_10574,N_10354,N_9837);
xnor U10575 (N_10575,N_10122,N_9839);
nand U10576 (N_10576,N_9815,N_10039);
and U10577 (N_10577,N_9791,N_9752);
and U10578 (N_10578,N_10448,N_9781);
or U10579 (N_10579,N_9813,N_9750);
and U10580 (N_10580,N_10249,N_10334);
and U10581 (N_10581,N_9778,N_10326);
and U10582 (N_10582,N_10478,N_10481);
and U10583 (N_10583,N_10154,N_10085);
and U10584 (N_10584,N_10417,N_10371);
xnor U10585 (N_10585,N_9984,N_9858);
nor U10586 (N_10586,N_10132,N_9751);
and U10587 (N_10587,N_10219,N_9764);
nor U10588 (N_10588,N_10137,N_10107);
or U10589 (N_10589,N_9766,N_9832);
nor U10590 (N_10590,N_10161,N_10155);
or U10591 (N_10591,N_9848,N_9899);
nand U10592 (N_10592,N_10033,N_10380);
or U10593 (N_10593,N_10242,N_10243);
and U10594 (N_10594,N_9794,N_10049);
nand U10595 (N_10595,N_9762,N_9923);
or U10596 (N_10596,N_10288,N_10362);
or U10597 (N_10597,N_10303,N_9941);
or U10598 (N_10598,N_10283,N_9936);
nor U10599 (N_10599,N_10135,N_10357);
nand U10600 (N_10600,N_9771,N_10455);
xor U10601 (N_10601,N_10125,N_9990);
or U10602 (N_10602,N_9811,N_9830);
and U10603 (N_10603,N_10160,N_10200);
nand U10604 (N_10604,N_9788,N_9980);
and U10605 (N_10605,N_10313,N_10424);
nor U10606 (N_10606,N_10465,N_10131);
nor U10607 (N_10607,N_10184,N_10094);
or U10608 (N_10608,N_9895,N_9880);
xor U10609 (N_10609,N_10173,N_9961);
or U10610 (N_10610,N_10466,N_10377);
and U10611 (N_10611,N_10213,N_10195);
nor U10612 (N_10612,N_10494,N_9935);
xnor U10613 (N_10613,N_10262,N_10407);
xor U10614 (N_10614,N_9974,N_9802);
nor U10615 (N_10615,N_9962,N_9846);
nand U10616 (N_10616,N_10401,N_9983);
xor U10617 (N_10617,N_10266,N_9878);
and U10618 (N_10618,N_10272,N_10278);
or U10619 (N_10619,N_10309,N_10359);
or U10620 (N_10620,N_9845,N_10358);
nor U10621 (N_10621,N_9793,N_10487);
or U10622 (N_10622,N_10051,N_9869);
nor U10623 (N_10623,N_10338,N_10329);
and U10624 (N_10624,N_9842,N_10254);
nand U10625 (N_10625,N_10328,N_10388);
or U10626 (N_10626,N_9809,N_10281);
or U10627 (N_10627,N_10336,N_10447);
nor U10628 (N_10628,N_10442,N_10223);
and U10629 (N_10629,N_10251,N_10096);
nand U10630 (N_10630,N_9982,N_9772);
or U10631 (N_10631,N_10292,N_9840);
and U10632 (N_10632,N_10182,N_9897);
and U10633 (N_10633,N_9853,N_10397);
nand U10634 (N_10634,N_10138,N_10115);
nand U10635 (N_10635,N_10013,N_9939);
nand U10636 (N_10636,N_9992,N_10151);
or U10637 (N_10637,N_10433,N_10183);
or U10638 (N_10638,N_9917,N_9942);
or U10639 (N_10639,N_9908,N_9987);
and U10640 (N_10640,N_9902,N_9951);
or U10641 (N_10641,N_10157,N_9873);
and U10642 (N_10642,N_10469,N_9922);
or U10643 (N_10643,N_10367,N_9890);
nand U10644 (N_10644,N_10308,N_10186);
nand U10645 (N_10645,N_10053,N_10024);
or U10646 (N_10646,N_10026,N_10119);
nand U10647 (N_10647,N_10178,N_10044);
nor U10648 (N_10648,N_10102,N_10229);
xnor U10649 (N_10649,N_9831,N_10341);
xnor U10650 (N_10650,N_10260,N_10414);
and U10651 (N_10651,N_10175,N_10286);
or U10652 (N_10652,N_9905,N_10485);
or U10653 (N_10653,N_9822,N_9993);
nand U10654 (N_10654,N_9915,N_10016);
xnor U10655 (N_10655,N_10345,N_10296);
or U10656 (N_10656,N_9814,N_9798);
or U10657 (N_10657,N_10073,N_9953);
nor U10658 (N_10658,N_10098,N_9776);
xnor U10659 (N_10659,N_9949,N_10344);
nor U10660 (N_10660,N_10325,N_10270);
or U10661 (N_10661,N_10127,N_10038);
and U10662 (N_10662,N_9838,N_10383);
xor U10663 (N_10663,N_10238,N_10314);
nand U10664 (N_10664,N_9792,N_10083);
nor U10665 (N_10665,N_10449,N_10043);
nor U10666 (N_10666,N_10196,N_10411);
nor U10667 (N_10667,N_10269,N_10028);
and U10668 (N_10668,N_10434,N_9801);
xor U10669 (N_10669,N_10022,N_10369);
nand U10670 (N_10670,N_10181,N_10475);
or U10671 (N_10671,N_10340,N_10074);
nand U10672 (N_10672,N_9972,N_10267);
nand U10673 (N_10673,N_10299,N_10258);
and U10674 (N_10674,N_9906,N_10143);
and U10675 (N_10675,N_10025,N_9894);
and U10676 (N_10676,N_10076,N_10228);
nand U10677 (N_10677,N_9777,N_10042);
and U10678 (N_10678,N_10446,N_10368);
or U10679 (N_10679,N_10405,N_10128);
nor U10680 (N_10680,N_10240,N_10106);
or U10681 (N_10681,N_10215,N_9938);
and U10682 (N_10682,N_10318,N_10439);
xor U10683 (N_10683,N_10384,N_9948);
nand U10684 (N_10684,N_10222,N_10188);
nor U10685 (N_10685,N_10280,N_9952);
nor U10686 (N_10686,N_10145,N_9898);
nor U10687 (N_10687,N_10265,N_9991);
nor U10688 (N_10688,N_10453,N_9844);
xor U10689 (N_10689,N_9924,N_9966);
nand U10690 (N_10690,N_9964,N_9865);
and U10691 (N_10691,N_10312,N_9876);
nand U10692 (N_10692,N_9988,N_9919);
and U10693 (N_10693,N_9796,N_10259);
nand U10694 (N_10694,N_10110,N_10169);
xor U10695 (N_10695,N_10470,N_10093);
xnor U10696 (N_10696,N_9947,N_10029);
xnor U10697 (N_10697,N_10090,N_10187);
or U10698 (N_10698,N_10263,N_10316);
and U10699 (N_10699,N_10264,N_9833);
nand U10700 (N_10700,N_10376,N_10440);
nor U10701 (N_10701,N_10070,N_10237);
nand U10702 (N_10702,N_9916,N_9963);
nor U10703 (N_10703,N_10393,N_9989);
or U10704 (N_10704,N_10017,N_9755);
nand U10705 (N_10705,N_10398,N_10046);
nor U10706 (N_10706,N_10462,N_10241);
or U10707 (N_10707,N_9866,N_10194);
nand U10708 (N_10708,N_10306,N_9860);
nand U10709 (N_10709,N_10488,N_10484);
nor U10710 (N_10710,N_10279,N_10450);
and U10711 (N_10711,N_10226,N_10121);
and U10712 (N_10712,N_10375,N_10476);
nor U10713 (N_10713,N_9790,N_10239);
xor U10714 (N_10714,N_10430,N_10490);
nor U10715 (N_10715,N_10374,N_10431);
nor U10716 (N_10716,N_10084,N_9757);
or U10717 (N_10717,N_10134,N_10198);
nand U10718 (N_10718,N_9875,N_10018);
xor U10719 (N_10719,N_10052,N_10032);
nor U10720 (N_10720,N_10146,N_9934);
nand U10721 (N_10721,N_10253,N_10031);
nor U10722 (N_10722,N_10342,N_10006);
and U10723 (N_10723,N_10463,N_10350);
nand U10724 (N_10724,N_9847,N_10403);
and U10725 (N_10725,N_9779,N_9825);
nand U10726 (N_10726,N_10477,N_10497);
and U10727 (N_10727,N_10395,N_10034);
and U10728 (N_10728,N_10271,N_10245);
and U10729 (N_10729,N_10480,N_10324);
and U10730 (N_10730,N_10346,N_10467);
nand U10731 (N_10731,N_10165,N_10495);
and U10732 (N_10732,N_10482,N_9877);
nor U10733 (N_10733,N_10202,N_10078);
and U10734 (N_10734,N_10483,N_9920);
nor U10735 (N_10735,N_9975,N_10413);
nand U10736 (N_10736,N_9753,N_9821);
nand U10737 (N_10737,N_10192,N_10436);
nor U10738 (N_10738,N_10330,N_10045);
nand U10739 (N_10739,N_10458,N_10012);
and U10740 (N_10740,N_10197,N_10355);
and U10741 (N_10741,N_10061,N_9756);
xnor U10742 (N_10742,N_9886,N_9958);
or U10743 (N_10743,N_10205,N_10075);
and U10744 (N_10744,N_10037,N_9971);
or U10745 (N_10745,N_10489,N_10360);
and U10746 (N_10746,N_10473,N_10220);
and U10747 (N_10747,N_10333,N_9871);
xnor U10748 (N_10748,N_10156,N_10111);
and U10749 (N_10749,N_10101,N_9765);
nor U10750 (N_10750,N_10117,N_10493);
nor U10751 (N_10751,N_10000,N_10422);
nand U10752 (N_10752,N_9864,N_10167);
or U10753 (N_10753,N_10123,N_10077);
nor U10754 (N_10754,N_10428,N_9965);
and U10755 (N_10755,N_9959,N_9892);
and U10756 (N_10756,N_10339,N_10129);
nor U10757 (N_10757,N_10319,N_10148);
nand U10758 (N_10758,N_10343,N_9836);
and U10759 (N_10759,N_9820,N_10019);
xor U10760 (N_10760,N_10352,N_9883);
nor U10761 (N_10761,N_10172,N_10317);
and U10762 (N_10762,N_9957,N_10007);
or U10763 (N_10763,N_9767,N_9785);
nor U10764 (N_10764,N_9855,N_10140);
xor U10765 (N_10765,N_10392,N_10464);
and U10766 (N_10766,N_10285,N_10452);
and U10767 (N_10767,N_9994,N_10185);
or U10768 (N_10768,N_10461,N_10438);
nor U10769 (N_10769,N_9888,N_10124);
nor U10770 (N_10770,N_10365,N_10058);
nor U10771 (N_10771,N_10166,N_10353);
nor U10772 (N_10772,N_10472,N_10193);
xor U10773 (N_10773,N_10114,N_10002);
nand U10774 (N_10774,N_9874,N_10116);
nand U10775 (N_10775,N_10150,N_9759);
nor U10776 (N_10776,N_10179,N_9852);
nand U10777 (N_10777,N_9870,N_9996);
or U10778 (N_10778,N_9818,N_10048);
nand U10779 (N_10779,N_10402,N_10180);
and U10780 (N_10780,N_10126,N_10415);
and U10781 (N_10781,N_10088,N_10305);
nor U10782 (N_10782,N_10204,N_9803);
xor U10783 (N_10783,N_10389,N_9827);
nor U10784 (N_10784,N_10335,N_10005);
and U10785 (N_10785,N_10191,N_10072);
nor U10786 (N_10786,N_9863,N_9929);
or U10787 (N_10787,N_10027,N_10212);
xnor U10788 (N_10788,N_10036,N_10327);
nand U10789 (N_10789,N_10099,N_9896);
nand U10790 (N_10790,N_10040,N_10203);
or U10791 (N_10791,N_10079,N_9783);
and U10792 (N_10792,N_10159,N_10423);
and U10793 (N_10793,N_9926,N_10250);
and U10794 (N_10794,N_10420,N_10244);
or U10795 (N_10795,N_10136,N_10276);
or U10796 (N_10796,N_9795,N_9955);
nand U10797 (N_10797,N_9807,N_10378);
or U10798 (N_10798,N_10014,N_10351);
xor U10799 (N_10799,N_9789,N_10468);
xnor U10800 (N_10800,N_10498,N_10089);
and U10801 (N_10801,N_10320,N_9911);
nor U10802 (N_10802,N_10248,N_10147);
and U10803 (N_10803,N_10086,N_9998);
or U10804 (N_10804,N_10059,N_10174);
nor U10805 (N_10805,N_10236,N_9856);
and U10806 (N_10806,N_10429,N_9808);
nor U10807 (N_10807,N_10451,N_10294);
xor U10808 (N_10808,N_9970,N_10055);
nor U10809 (N_10809,N_9819,N_9782);
or U10810 (N_10810,N_9758,N_10323);
nand U10811 (N_10811,N_9910,N_10302);
and U10812 (N_10812,N_10307,N_9805);
or U10813 (N_10813,N_10287,N_9930);
xnor U10814 (N_10814,N_10023,N_9967);
nand U10815 (N_10815,N_10277,N_9940);
and U10816 (N_10816,N_10257,N_10168);
xnor U10817 (N_10817,N_10149,N_10170);
or U10818 (N_10818,N_10385,N_10141);
nand U10819 (N_10819,N_10171,N_10206);
nor U10820 (N_10820,N_10457,N_10035);
nand U10821 (N_10821,N_10010,N_10139);
or U10822 (N_10822,N_9804,N_9995);
nor U10823 (N_10823,N_9889,N_9760);
and U10824 (N_10824,N_10230,N_9914);
xnor U10825 (N_10825,N_10460,N_9986);
or U10826 (N_10826,N_9810,N_9784);
or U10827 (N_10827,N_9954,N_10062);
nor U10828 (N_10828,N_10337,N_9997);
nor U10829 (N_10829,N_10152,N_9843);
nand U10830 (N_10830,N_10142,N_10054);
or U10831 (N_10831,N_9925,N_9829);
and U10832 (N_10832,N_10426,N_10095);
or U10833 (N_10833,N_9921,N_9773);
nand U10834 (N_10834,N_10216,N_9868);
or U10835 (N_10835,N_10008,N_10363);
and U10836 (N_10836,N_10047,N_10004);
nor U10837 (N_10837,N_10322,N_10066);
nor U10838 (N_10838,N_10189,N_10227);
and U10839 (N_10839,N_10432,N_10479);
or U10840 (N_10840,N_9978,N_10109);
and U10841 (N_10841,N_10256,N_10232);
or U10842 (N_10842,N_9862,N_10298);
xnor U10843 (N_10843,N_10290,N_10209);
xnor U10844 (N_10844,N_9933,N_10391);
nand U10845 (N_10845,N_9851,N_10459);
and U10846 (N_10846,N_9799,N_10224);
and U10847 (N_10847,N_9817,N_10082);
nor U10848 (N_10848,N_10087,N_10347);
or U10849 (N_10849,N_9927,N_10221);
or U10850 (N_10850,N_9816,N_9977);
nor U10851 (N_10851,N_10108,N_9857);
or U10852 (N_10852,N_10003,N_9885);
and U10853 (N_10853,N_9968,N_9774);
nor U10854 (N_10854,N_9937,N_9835);
and U10855 (N_10855,N_9973,N_10284);
or U10856 (N_10856,N_10427,N_10486);
or U10857 (N_10857,N_9823,N_9960);
nor U10858 (N_10858,N_10410,N_10394);
and U10859 (N_10859,N_10399,N_9884);
or U10860 (N_10860,N_10080,N_10404);
nand U10861 (N_10861,N_10400,N_10282);
nor U10862 (N_10862,N_9769,N_9969);
nand U10863 (N_10863,N_9945,N_10020);
or U10864 (N_10864,N_10177,N_10234);
and U10865 (N_10865,N_10387,N_10112);
nor U10866 (N_10866,N_9981,N_10441);
or U10867 (N_10867,N_9950,N_10372);
nand U10868 (N_10868,N_10063,N_9867);
or U10869 (N_10869,N_10301,N_10255);
nor U10870 (N_10870,N_10364,N_10310);
nor U10871 (N_10871,N_10409,N_10252);
nand U10872 (N_10872,N_10130,N_10100);
and U10873 (N_10873,N_10315,N_10067);
xnor U10874 (N_10874,N_9780,N_10133);
or U10875 (N_10875,N_9901,N_9989);
and U10876 (N_10876,N_10370,N_10291);
and U10877 (N_10877,N_9770,N_10466);
or U10878 (N_10878,N_10348,N_10144);
and U10879 (N_10879,N_9969,N_9907);
nor U10880 (N_10880,N_10469,N_10194);
and U10881 (N_10881,N_9782,N_10136);
nor U10882 (N_10882,N_9935,N_10220);
nor U10883 (N_10883,N_10256,N_9786);
or U10884 (N_10884,N_10368,N_10071);
nor U10885 (N_10885,N_10041,N_9799);
xnor U10886 (N_10886,N_10372,N_10271);
nor U10887 (N_10887,N_9843,N_10472);
or U10888 (N_10888,N_9993,N_9881);
and U10889 (N_10889,N_9804,N_10141);
and U10890 (N_10890,N_10119,N_10181);
and U10891 (N_10891,N_9852,N_10373);
nand U10892 (N_10892,N_9868,N_9810);
or U10893 (N_10893,N_9940,N_10072);
and U10894 (N_10894,N_10164,N_10079);
or U10895 (N_10895,N_10332,N_9811);
xor U10896 (N_10896,N_10327,N_10040);
nand U10897 (N_10897,N_9983,N_10348);
nand U10898 (N_10898,N_10219,N_10456);
or U10899 (N_10899,N_10478,N_10326);
xnor U10900 (N_10900,N_10238,N_9842);
or U10901 (N_10901,N_10421,N_10424);
and U10902 (N_10902,N_10092,N_10400);
nand U10903 (N_10903,N_9769,N_10282);
and U10904 (N_10904,N_10262,N_9762);
and U10905 (N_10905,N_9903,N_10436);
nand U10906 (N_10906,N_10374,N_9910);
nor U10907 (N_10907,N_10123,N_10458);
and U10908 (N_10908,N_10104,N_10442);
and U10909 (N_10909,N_10233,N_10241);
or U10910 (N_10910,N_10382,N_10073);
or U10911 (N_10911,N_10386,N_9767);
or U10912 (N_10912,N_10492,N_9764);
nand U10913 (N_10913,N_10396,N_10056);
nand U10914 (N_10914,N_10327,N_10397);
nand U10915 (N_10915,N_9928,N_10154);
or U10916 (N_10916,N_10237,N_10045);
and U10917 (N_10917,N_10159,N_10486);
nor U10918 (N_10918,N_10040,N_10433);
and U10919 (N_10919,N_9939,N_10065);
or U10920 (N_10920,N_9799,N_10268);
or U10921 (N_10921,N_10016,N_10237);
and U10922 (N_10922,N_9976,N_10338);
or U10923 (N_10923,N_10361,N_10088);
nor U10924 (N_10924,N_10331,N_10293);
nand U10925 (N_10925,N_9990,N_10236);
and U10926 (N_10926,N_10478,N_10391);
xor U10927 (N_10927,N_10227,N_10117);
or U10928 (N_10928,N_10348,N_10368);
xnor U10929 (N_10929,N_10347,N_10453);
nand U10930 (N_10930,N_10144,N_10146);
nor U10931 (N_10931,N_10451,N_10156);
nor U10932 (N_10932,N_10193,N_10247);
nand U10933 (N_10933,N_10281,N_9852);
nor U10934 (N_10934,N_10028,N_10410);
and U10935 (N_10935,N_9826,N_10206);
or U10936 (N_10936,N_9992,N_10047);
nand U10937 (N_10937,N_10367,N_10016);
xnor U10938 (N_10938,N_10300,N_10028);
nand U10939 (N_10939,N_10134,N_10068);
nand U10940 (N_10940,N_9990,N_10373);
nand U10941 (N_10941,N_9790,N_10105);
xor U10942 (N_10942,N_9778,N_10420);
nand U10943 (N_10943,N_10184,N_10485);
nand U10944 (N_10944,N_9883,N_10244);
and U10945 (N_10945,N_10166,N_10213);
nand U10946 (N_10946,N_10260,N_10242);
and U10947 (N_10947,N_9970,N_10115);
nand U10948 (N_10948,N_9933,N_10104);
or U10949 (N_10949,N_9898,N_9980);
and U10950 (N_10950,N_9993,N_10050);
and U10951 (N_10951,N_10388,N_9894);
and U10952 (N_10952,N_10311,N_9852);
nand U10953 (N_10953,N_10300,N_10240);
and U10954 (N_10954,N_9935,N_10008);
and U10955 (N_10955,N_10191,N_10402);
nor U10956 (N_10956,N_10373,N_9867);
or U10957 (N_10957,N_10416,N_10009);
xnor U10958 (N_10958,N_10479,N_10226);
nor U10959 (N_10959,N_10053,N_10434);
and U10960 (N_10960,N_10353,N_9910);
nand U10961 (N_10961,N_9930,N_10140);
and U10962 (N_10962,N_10323,N_9905);
nor U10963 (N_10963,N_9867,N_10481);
nand U10964 (N_10964,N_10316,N_10470);
and U10965 (N_10965,N_10139,N_10389);
and U10966 (N_10966,N_10403,N_9831);
nor U10967 (N_10967,N_9866,N_10185);
nand U10968 (N_10968,N_10378,N_10414);
or U10969 (N_10969,N_10422,N_10070);
nor U10970 (N_10970,N_10104,N_10324);
and U10971 (N_10971,N_10377,N_10401);
nor U10972 (N_10972,N_10162,N_9818);
nor U10973 (N_10973,N_10394,N_10004);
nor U10974 (N_10974,N_10494,N_10019);
nand U10975 (N_10975,N_10334,N_9964);
or U10976 (N_10976,N_10105,N_10134);
nand U10977 (N_10977,N_9962,N_10428);
or U10978 (N_10978,N_9834,N_9924);
or U10979 (N_10979,N_10305,N_10036);
nand U10980 (N_10980,N_10202,N_10161);
and U10981 (N_10981,N_9946,N_10133);
nor U10982 (N_10982,N_9793,N_10412);
nand U10983 (N_10983,N_10159,N_9786);
and U10984 (N_10984,N_10151,N_10412);
or U10985 (N_10985,N_10237,N_9782);
and U10986 (N_10986,N_9905,N_10089);
nand U10987 (N_10987,N_9857,N_9935);
or U10988 (N_10988,N_9798,N_10390);
or U10989 (N_10989,N_10061,N_9919);
and U10990 (N_10990,N_10295,N_9765);
nand U10991 (N_10991,N_10279,N_10135);
and U10992 (N_10992,N_9990,N_10046);
or U10993 (N_10993,N_9915,N_10210);
nand U10994 (N_10994,N_10459,N_10007);
or U10995 (N_10995,N_10038,N_10160);
and U10996 (N_10996,N_9773,N_9849);
xnor U10997 (N_10997,N_9853,N_9811);
nor U10998 (N_10998,N_10455,N_10259);
xnor U10999 (N_10999,N_10377,N_10008);
nor U11000 (N_11000,N_10294,N_10318);
nor U11001 (N_11001,N_10329,N_10060);
or U11002 (N_11002,N_10039,N_9917);
and U11003 (N_11003,N_10475,N_10130);
nor U11004 (N_11004,N_9796,N_10072);
nor U11005 (N_11005,N_9952,N_10209);
nand U11006 (N_11006,N_9974,N_10276);
xor U11007 (N_11007,N_10078,N_10349);
or U11008 (N_11008,N_10455,N_10292);
or U11009 (N_11009,N_9958,N_9781);
nor U11010 (N_11010,N_10171,N_10282);
nand U11011 (N_11011,N_9856,N_10340);
or U11012 (N_11012,N_10255,N_10351);
nor U11013 (N_11013,N_10122,N_9836);
and U11014 (N_11014,N_10157,N_10107);
xor U11015 (N_11015,N_9900,N_10350);
and U11016 (N_11016,N_10194,N_10009);
nand U11017 (N_11017,N_9981,N_10242);
xnor U11018 (N_11018,N_9857,N_10280);
and U11019 (N_11019,N_9906,N_10235);
nand U11020 (N_11020,N_10209,N_10274);
or U11021 (N_11021,N_10098,N_10363);
or U11022 (N_11022,N_10021,N_10276);
nand U11023 (N_11023,N_10247,N_10166);
nand U11024 (N_11024,N_9995,N_10307);
and U11025 (N_11025,N_10147,N_10445);
and U11026 (N_11026,N_10215,N_10087);
nand U11027 (N_11027,N_10279,N_9844);
nand U11028 (N_11028,N_9890,N_9918);
nand U11029 (N_11029,N_10376,N_10112);
or U11030 (N_11030,N_10228,N_9760);
nand U11031 (N_11031,N_10453,N_10490);
and U11032 (N_11032,N_10003,N_10321);
nor U11033 (N_11033,N_9987,N_10485);
nor U11034 (N_11034,N_10191,N_9813);
or U11035 (N_11035,N_10281,N_10463);
and U11036 (N_11036,N_10423,N_9899);
and U11037 (N_11037,N_10433,N_10238);
and U11038 (N_11038,N_10444,N_10395);
and U11039 (N_11039,N_9876,N_9875);
nor U11040 (N_11040,N_10242,N_10329);
and U11041 (N_11041,N_10470,N_10006);
nor U11042 (N_11042,N_10329,N_10275);
nor U11043 (N_11043,N_10033,N_10090);
and U11044 (N_11044,N_9960,N_10209);
xor U11045 (N_11045,N_10048,N_10071);
and U11046 (N_11046,N_10432,N_10289);
or U11047 (N_11047,N_10056,N_10482);
nand U11048 (N_11048,N_10125,N_10377);
nor U11049 (N_11049,N_10060,N_10302);
or U11050 (N_11050,N_10184,N_10307);
or U11051 (N_11051,N_10159,N_9778);
and U11052 (N_11052,N_10117,N_9807);
or U11053 (N_11053,N_10249,N_9982);
nand U11054 (N_11054,N_10329,N_10296);
and U11055 (N_11055,N_10227,N_10347);
and U11056 (N_11056,N_10056,N_10348);
or U11057 (N_11057,N_10240,N_10299);
nand U11058 (N_11058,N_10330,N_10167);
nor U11059 (N_11059,N_10317,N_10251);
xnor U11060 (N_11060,N_10352,N_9781);
or U11061 (N_11061,N_10429,N_9916);
or U11062 (N_11062,N_10144,N_10159);
nor U11063 (N_11063,N_10468,N_9823);
or U11064 (N_11064,N_10112,N_10235);
and U11065 (N_11065,N_10135,N_10499);
nor U11066 (N_11066,N_10072,N_10283);
nor U11067 (N_11067,N_10189,N_9779);
nor U11068 (N_11068,N_10169,N_10390);
nor U11069 (N_11069,N_9770,N_10070);
or U11070 (N_11070,N_10242,N_10349);
xnor U11071 (N_11071,N_10493,N_10334);
nor U11072 (N_11072,N_9993,N_9871);
and U11073 (N_11073,N_10286,N_10303);
xnor U11074 (N_11074,N_10179,N_9900);
or U11075 (N_11075,N_9951,N_10085);
or U11076 (N_11076,N_9958,N_10289);
and U11077 (N_11077,N_9856,N_10298);
or U11078 (N_11078,N_10029,N_10481);
or U11079 (N_11079,N_9753,N_9884);
nor U11080 (N_11080,N_9883,N_10393);
or U11081 (N_11081,N_9858,N_10114);
or U11082 (N_11082,N_10146,N_9844);
and U11083 (N_11083,N_10391,N_10016);
nand U11084 (N_11084,N_9949,N_10487);
nor U11085 (N_11085,N_10007,N_10067);
or U11086 (N_11086,N_10030,N_10461);
xnor U11087 (N_11087,N_10390,N_10342);
nand U11088 (N_11088,N_9866,N_10357);
xnor U11089 (N_11089,N_9865,N_10098);
nand U11090 (N_11090,N_10318,N_10297);
xor U11091 (N_11091,N_9837,N_9822);
and U11092 (N_11092,N_9834,N_9917);
and U11093 (N_11093,N_9957,N_10030);
xnor U11094 (N_11094,N_10041,N_10243);
or U11095 (N_11095,N_9942,N_10417);
or U11096 (N_11096,N_10403,N_9776);
xnor U11097 (N_11097,N_10205,N_9929);
and U11098 (N_11098,N_9820,N_10384);
and U11099 (N_11099,N_10183,N_10170);
or U11100 (N_11100,N_10028,N_9952);
xor U11101 (N_11101,N_10362,N_9930);
nor U11102 (N_11102,N_10065,N_9888);
nor U11103 (N_11103,N_10093,N_9872);
nand U11104 (N_11104,N_10413,N_10298);
nor U11105 (N_11105,N_10335,N_10187);
and U11106 (N_11106,N_10462,N_9779);
and U11107 (N_11107,N_10449,N_10462);
and U11108 (N_11108,N_9940,N_9985);
nand U11109 (N_11109,N_10405,N_10004);
xnor U11110 (N_11110,N_9802,N_9848);
or U11111 (N_11111,N_9785,N_9981);
or U11112 (N_11112,N_10121,N_9920);
nand U11113 (N_11113,N_9892,N_10324);
and U11114 (N_11114,N_9929,N_10222);
xnor U11115 (N_11115,N_10390,N_10029);
xnor U11116 (N_11116,N_10384,N_10363);
or U11117 (N_11117,N_9773,N_10237);
or U11118 (N_11118,N_10205,N_10121);
xnor U11119 (N_11119,N_10229,N_10224);
or U11120 (N_11120,N_10280,N_9968);
nand U11121 (N_11121,N_9849,N_9775);
or U11122 (N_11122,N_10459,N_10199);
xnor U11123 (N_11123,N_10485,N_10391);
or U11124 (N_11124,N_9963,N_10497);
nand U11125 (N_11125,N_10346,N_9989);
nand U11126 (N_11126,N_10204,N_9766);
nand U11127 (N_11127,N_10354,N_9992);
and U11128 (N_11128,N_10467,N_10399);
and U11129 (N_11129,N_10001,N_10382);
nand U11130 (N_11130,N_10398,N_10197);
and U11131 (N_11131,N_10154,N_10286);
and U11132 (N_11132,N_9755,N_10375);
or U11133 (N_11133,N_9961,N_10266);
or U11134 (N_11134,N_10310,N_10388);
nor U11135 (N_11135,N_9936,N_10364);
xor U11136 (N_11136,N_9897,N_10248);
xnor U11137 (N_11137,N_9839,N_10171);
or U11138 (N_11138,N_10345,N_9890);
or U11139 (N_11139,N_9760,N_9807);
nor U11140 (N_11140,N_9976,N_10319);
or U11141 (N_11141,N_10059,N_10216);
nor U11142 (N_11142,N_10433,N_10349);
nand U11143 (N_11143,N_9789,N_10370);
and U11144 (N_11144,N_10217,N_9816);
nor U11145 (N_11145,N_10473,N_10015);
xor U11146 (N_11146,N_10241,N_9769);
and U11147 (N_11147,N_10246,N_9970);
or U11148 (N_11148,N_10079,N_9899);
nand U11149 (N_11149,N_9983,N_10085);
nand U11150 (N_11150,N_9751,N_10448);
or U11151 (N_11151,N_10486,N_10198);
nor U11152 (N_11152,N_10464,N_10099);
and U11153 (N_11153,N_10163,N_10327);
nor U11154 (N_11154,N_10026,N_10134);
nand U11155 (N_11155,N_10213,N_10075);
and U11156 (N_11156,N_10048,N_9957);
nand U11157 (N_11157,N_10267,N_10061);
and U11158 (N_11158,N_10018,N_9970);
nor U11159 (N_11159,N_10339,N_10393);
and U11160 (N_11160,N_10386,N_10212);
and U11161 (N_11161,N_9842,N_10044);
nand U11162 (N_11162,N_9790,N_9917);
or U11163 (N_11163,N_10393,N_10167);
or U11164 (N_11164,N_10225,N_10193);
or U11165 (N_11165,N_9996,N_9979);
nor U11166 (N_11166,N_10166,N_9995);
and U11167 (N_11167,N_9890,N_9875);
nand U11168 (N_11168,N_9754,N_9759);
nor U11169 (N_11169,N_10318,N_10109);
xor U11170 (N_11170,N_10291,N_9912);
nand U11171 (N_11171,N_10139,N_10011);
nand U11172 (N_11172,N_9785,N_9885);
nor U11173 (N_11173,N_10329,N_10098);
and U11174 (N_11174,N_9791,N_10023);
nand U11175 (N_11175,N_10026,N_10314);
nor U11176 (N_11176,N_10346,N_9966);
xnor U11177 (N_11177,N_10129,N_10303);
and U11178 (N_11178,N_10190,N_10187);
nor U11179 (N_11179,N_10162,N_9804);
nand U11180 (N_11180,N_10258,N_9882);
and U11181 (N_11181,N_10278,N_9972);
or U11182 (N_11182,N_10243,N_10163);
or U11183 (N_11183,N_9820,N_10321);
nor U11184 (N_11184,N_9900,N_9838);
or U11185 (N_11185,N_10442,N_9802);
nor U11186 (N_11186,N_9839,N_10230);
and U11187 (N_11187,N_10007,N_9914);
nor U11188 (N_11188,N_10027,N_9912);
nor U11189 (N_11189,N_9950,N_9895);
nand U11190 (N_11190,N_9965,N_10028);
nand U11191 (N_11191,N_10320,N_10177);
nor U11192 (N_11192,N_10415,N_9932);
nor U11193 (N_11193,N_9780,N_10404);
nand U11194 (N_11194,N_10415,N_10458);
nor U11195 (N_11195,N_9929,N_10210);
and U11196 (N_11196,N_10183,N_10179);
xor U11197 (N_11197,N_10082,N_9916);
nand U11198 (N_11198,N_9813,N_9877);
or U11199 (N_11199,N_10414,N_10131);
and U11200 (N_11200,N_10035,N_10239);
or U11201 (N_11201,N_9819,N_10074);
and U11202 (N_11202,N_10041,N_10180);
or U11203 (N_11203,N_10222,N_9903);
nand U11204 (N_11204,N_9807,N_10432);
and U11205 (N_11205,N_9918,N_10323);
nand U11206 (N_11206,N_9956,N_10138);
and U11207 (N_11207,N_10102,N_9827);
or U11208 (N_11208,N_10319,N_10258);
or U11209 (N_11209,N_10281,N_9822);
and U11210 (N_11210,N_9852,N_10456);
xnor U11211 (N_11211,N_9760,N_10095);
and U11212 (N_11212,N_9957,N_9837);
xnor U11213 (N_11213,N_10300,N_10339);
and U11214 (N_11214,N_9846,N_10441);
and U11215 (N_11215,N_9964,N_10412);
nor U11216 (N_11216,N_10351,N_10479);
and U11217 (N_11217,N_9894,N_9978);
or U11218 (N_11218,N_9882,N_10046);
or U11219 (N_11219,N_10258,N_10445);
nor U11220 (N_11220,N_10079,N_10137);
and U11221 (N_11221,N_10091,N_10219);
xnor U11222 (N_11222,N_10273,N_10218);
nor U11223 (N_11223,N_9856,N_9776);
nor U11224 (N_11224,N_10396,N_9823);
nor U11225 (N_11225,N_10205,N_10352);
and U11226 (N_11226,N_9863,N_10308);
nand U11227 (N_11227,N_10116,N_9780);
nor U11228 (N_11228,N_9901,N_10090);
nand U11229 (N_11229,N_10393,N_10281);
nor U11230 (N_11230,N_10297,N_10253);
or U11231 (N_11231,N_10119,N_10268);
nand U11232 (N_11232,N_9787,N_9781);
nand U11233 (N_11233,N_10416,N_10314);
nand U11234 (N_11234,N_10466,N_10168);
or U11235 (N_11235,N_9955,N_10359);
nand U11236 (N_11236,N_9904,N_9852);
nand U11237 (N_11237,N_10118,N_10475);
and U11238 (N_11238,N_9913,N_10451);
nand U11239 (N_11239,N_10344,N_10031);
and U11240 (N_11240,N_9882,N_10123);
nand U11241 (N_11241,N_10344,N_10098);
or U11242 (N_11242,N_10225,N_10260);
nand U11243 (N_11243,N_10389,N_9859);
and U11244 (N_11244,N_10108,N_10361);
and U11245 (N_11245,N_9946,N_10343);
and U11246 (N_11246,N_10422,N_9792);
nor U11247 (N_11247,N_10373,N_9820);
or U11248 (N_11248,N_9824,N_10295);
and U11249 (N_11249,N_10167,N_9868);
nand U11250 (N_11250,N_10726,N_10850);
nor U11251 (N_11251,N_10952,N_10993);
or U11252 (N_11252,N_11149,N_11186);
and U11253 (N_11253,N_10748,N_10608);
and U11254 (N_11254,N_10692,N_10628);
or U11255 (N_11255,N_10684,N_11178);
nand U11256 (N_11256,N_10507,N_10553);
nor U11257 (N_11257,N_11130,N_10916);
nand U11258 (N_11258,N_10731,N_10764);
and U11259 (N_11259,N_11029,N_11013);
xnor U11260 (N_11260,N_11227,N_10574);
or U11261 (N_11261,N_11069,N_11117);
nand U11262 (N_11262,N_10554,N_10552);
xnor U11263 (N_11263,N_10898,N_11153);
xor U11264 (N_11264,N_10905,N_10638);
xor U11265 (N_11265,N_10822,N_11123);
nand U11266 (N_11266,N_11049,N_10754);
nor U11267 (N_11267,N_10832,N_11216);
or U11268 (N_11268,N_10788,N_10977);
xor U11269 (N_11269,N_10947,N_11067);
or U11270 (N_11270,N_11134,N_10654);
or U11271 (N_11271,N_11062,N_11147);
xor U11272 (N_11272,N_10837,N_11143);
nand U11273 (N_11273,N_10680,N_11071);
and U11274 (N_11274,N_10596,N_11107);
nor U11275 (N_11275,N_10941,N_10547);
nor U11276 (N_11276,N_10845,N_10529);
nor U11277 (N_11277,N_10694,N_11129);
xnor U11278 (N_11278,N_10716,N_11128);
or U11279 (N_11279,N_10683,N_11089);
nand U11280 (N_11280,N_11002,N_10972);
and U11281 (N_11281,N_10917,N_11116);
and U11282 (N_11282,N_11198,N_10755);
nand U11283 (N_11283,N_11213,N_10923);
xnor U11284 (N_11284,N_10909,N_10899);
nand U11285 (N_11285,N_10734,N_11088);
xor U11286 (N_11286,N_11166,N_10970);
nor U11287 (N_11287,N_10718,N_10636);
or U11288 (N_11288,N_10802,N_10777);
xnor U11289 (N_11289,N_10519,N_10906);
and U11290 (N_11290,N_10512,N_10620);
nor U11291 (N_11291,N_10843,N_10518);
or U11292 (N_11292,N_10880,N_10690);
xor U11293 (N_11293,N_10665,N_10752);
nor U11294 (N_11294,N_10723,N_10650);
or U11295 (N_11295,N_11025,N_11161);
or U11296 (N_11296,N_10924,N_10659);
nor U11297 (N_11297,N_11032,N_10773);
or U11298 (N_11298,N_11023,N_10876);
and U11299 (N_11299,N_10908,N_11103);
or U11300 (N_11300,N_11093,N_10869);
or U11301 (N_11301,N_10535,N_10696);
and U11302 (N_11302,N_11036,N_10522);
nand U11303 (N_11303,N_10576,N_10767);
or U11304 (N_11304,N_10921,N_11090);
xnor U11305 (N_11305,N_10804,N_11192);
nor U11306 (N_11306,N_10691,N_10846);
nor U11307 (N_11307,N_11208,N_10634);
nand U11308 (N_11308,N_10724,N_10893);
and U11309 (N_11309,N_11200,N_10737);
xnor U11310 (N_11310,N_11185,N_11115);
and U11311 (N_11311,N_10791,N_10939);
xor U11312 (N_11312,N_11160,N_10673);
nand U11313 (N_11313,N_10819,N_11211);
and U11314 (N_11314,N_11188,N_11196);
xnor U11315 (N_11315,N_10581,N_10931);
and U11316 (N_11316,N_11110,N_11060);
and U11317 (N_11317,N_10672,N_10753);
nand U11318 (N_11318,N_10514,N_10763);
and U11319 (N_11319,N_11068,N_10541);
or U11320 (N_11320,N_10818,N_11114);
nand U11321 (N_11321,N_10999,N_10859);
or U11322 (N_11322,N_11207,N_10833);
nor U11323 (N_11323,N_11054,N_10885);
and U11324 (N_11324,N_11073,N_10844);
and U11325 (N_11325,N_11174,N_11173);
or U11326 (N_11326,N_10635,N_10558);
or U11327 (N_11327,N_11236,N_10681);
and U11328 (N_11328,N_10536,N_10935);
and U11329 (N_11329,N_10912,N_10897);
and U11330 (N_11330,N_10772,N_10569);
nor U11331 (N_11331,N_11096,N_10639);
or U11332 (N_11332,N_10984,N_10983);
nor U11333 (N_11333,N_10761,N_10936);
xnor U11334 (N_11334,N_10820,N_10873);
xor U11335 (N_11335,N_11039,N_10814);
nor U11336 (N_11336,N_11187,N_10711);
xnor U11337 (N_11337,N_10511,N_10652);
and U11338 (N_11338,N_10858,N_10913);
or U11339 (N_11339,N_10591,N_10625);
nand U11340 (N_11340,N_11124,N_10544);
nand U11341 (N_11341,N_10875,N_10828);
nand U11342 (N_11342,N_11119,N_11183);
nand U11343 (N_11343,N_10594,N_10851);
or U11344 (N_11344,N_10823,N_10821);
or U11345 (N_11345,N_10521,N_10870);
nor U11346 (N_11346,N_10728,N_11095);
nor U11347 (N_11347,N_10901,N_11182);
xnor U11348 (N_11348,N_10903,N_10747);
nor U11349 (N_11349,N_10915,N_10733);
and U11350 (N_11350,N_11136,N_11004);
nand U11351 (N_11351,N_10611,N_10964);
or U11352 (N_11352,N_11201,N_10686);
nand U11353 (N_11353,N_10550,N_10895);
nand U11354 (N_11354,N_10602,N_10729);
nand U11355 (N_11355,N_10735,N_10907);
nand U11356 (N_11356,N_10701,N_11078);
xnor U11357 (N_11357,N_10528,N_10987);
nand U11358 (N_11358,N_10888,N_11005);
nand U11359 (N_11359,N_10532,N_10978);
xnor U11360 (N_11360,N_10570,N_10838);
and U11361 (N_11361,N_10505,N_11242);
xor U11362 (N_11362,N_11138,N_11214);
and U11363 (N_11363,N_10593,N_10744);
nor U11364 (N_11364,N_11046,N_10586);
or U11365 (N_11365,N_10517,N_10504);
and U11366 (N_11366,N_10891,N_11132);
nand U11367 (N_11367,N_11047,N_10704);
and U11368 (N_11368,N_10920,N_11194);
and U11369 (N_11369,N_11246,N_10644);
nor U11370 (N_11370,N_10633,N_10961);
or U11371 (N_11371,N_11197,N_11168);
and U11372 (N_11372,N_10709,N_10808);
and U11373 (N_11373,N_11191,N_10548);
and U11374 (N_11374,N_10966,N_10693);
or U11375 (N_11375,N_10948,N_10730);
or U11376 (N_11376,N_10982,N_11059);
or U11377 (N_11377,N_10577,N_10661);
or U11378 (N_11378,N_10894,N_10831);
nand U11379 (N_11379,N_10991,N_11063);
or U11380 (N_11380,N_11008,N_11225);
or U11381 (N_11381,N_10623,N_11003);
and U11382 (N_11382,N_10938,N_10979);
or U11383 (N_11383,N_11235,N_10604);
xnor U11384 (N_11384,N_10925,N_10955);
or U11385 (N_11385,N_10572,N_10809);
or U11386 (N_11386,N_11238,N_10933);
or U11387 (N_11387,N_10758,N_10958);
nand U11388 (N_11388,N_10525,N_11131);
and U11389 (N_11389,N_11206,N_10962);
nor U11390 (N_11390,N_10712,N_10877);
nor U11391 (N_11391,N_10688,N_11177);
xor U11392 (N_11392,N_11065,N_10995);
or U11393 (N_11393,N_11048,N_11229);
xor U11394 (N_11394,N_11024,N_10806);
and U11395 (N_11395,N_11195,N_11179);
nand U11396 (N_11396,N_10768,N_10781);
nor U11397 (N_11397,N_10871,N_10674);
nand U11398 (N_11398,N_10649,N_11070);
and U11399 (N_11399,N_11156,N_10539);
and U11400 (N_11400,N_11150,N_10615);
and U11401 (N_11401,N_10957,N_10578);
nor U11402 (N_11402,N_10805,N_11030);
nor U11403 (N_11403,N_10827,N_10813);
or U11404 (N_11404,N_10883,N_11021);
nand U11405 (N_11405,N_10789,N_10516);
or U11406 (N_11406,N_10646,N_10655);
nand U11407 (N_11407,N_10662,N_10657);
and U11408 (N_11408,N_10971,N_10765);
and U11409 (N_11409,N_10904,N_10559);
nand U11410 (N_11410,N_10700,N_11017);
nor U11411 (N_11411,N_10780,N_11012);
and U11412 (N_11412,N_11237,N_11170);
nand U11413 (N_11413,N_11244,N_11220);
nor U11414 (N_11414,N_10515,N_10727);
nand U11415 (N_11415,N_11239,N_10595);
or U11416 (N_11416,N_10956,N_10703);
nor U11417 (N_11417,N_11106,N_10699);
nand U11418 (N_11418,N_10862,N_10841);
or U11419 (N_11419,N_10616,N_10798);
nor U11420 (N_11420,N_10563,N_11218);
nor U11421 (N_11421,N_10695,N_11072);
and U11422 (N_11422,N_10946,N_10713);
nand U11423 (N_11423,N_10992,N_10756);
nand U11424 (N_11424,N_10617,N_10857);
and U11425 (N_11425,N_11076,N_10951);
nor U11426 (N_11426,N_10524,N_11109);
nand U11427 (N_11427,N_10679,N_10531);
nor U11428 (N_11428,N_11248,N_10775);
or U11429 (N_11429,N_10836,N_10597);
nand U11430 (N_11430,N_10751,N_10868);
or U11431 (N_11431,N_11180,N_10782);
nor U11432 (N_11432,N_10799,N_10668);
and U11433 (N_11433,N_10865,N_11204);
or U11434 (N_11434,N_10998,N_10797);
nand U11435 (N_11435,N_10863,N_11152);
and U11436 (N_11436,N_11027,N_10551);
nor U11437 (N_11437,N_10682,N_10878);
and U11438 (N_11438,N_10896,N_10826);
and U11439 (N_11439,N_11233,N_10705);
or U11440 (N_11440,N_11241,N_10592);
xnor U11441 (N_11441,N_10526,N_10603);
xor U11442 (N_11442,N_10940,N_10835);
or U11443 (N_11443,N_10557,N_11077);
and U11444 (N_11444,N_10612,N_10509);
nand U11445 (N_11445,N_10932,N_10583);
nand U11446 (N_11446,N_11155,N_10549);
nand U11447 (N_11447,N_10934,N_10879);
nor U11448 (N_11448,N_10825,N_10842);
or U11449 (N_11449,N_10783,N_10757);
nor U11450 (N_11450,N_11037,N_10629);
or U11451 (N_11451,N_11135,N_10839);
nor U11452 (N_11452,N_10508,N_10817);
xor U11453 (N_11453,N_10506,N_10543);
nor U11454 (N_11454,N_11243,N_10658);
xnor U11455 (N_11455,N_10520,N_11112);
nand U11456 (N_11456,N_10601,N_10969);
nand U11457 (N_11457,N_11104,N_11041);
nand U11458 (N_11458,N_11097,N_10588);
or U11459 (N_11459,N_10965,N_10954);
or U11460 (N_11460,N_11121,N_11042);
and U11461 (N_11461,N_10619,N_10555);
and U11462 (N_11462,N_10803,N_11190);
and U11463 (N_11463,N_10990,N_10985);
or U11464 (N_11464,N_11175,N_10627);
nor U11465 (N_11465,N_10584,N_10847);
and U11466 (N_11466,N_10632,N_11040);
and U11467 (N_11467,N_10937,N_10725);
nand U11468 (N_11468,N_10647,N_11105);
and U11469 (N_11469,N_10779,N_11165);
xor U11470 (N_11470,N_10560,N_11189);
or U11471 (N_11471,N_11169,N_10786);
and U11472 (N_11472,N_10527,N_11234);
nand U11473 (N_11473,N_10943,N_10538);
xor U11474 (N_11474,N_11159,N_10864);
xnor U11475 (N_11475,N_11001,N_10562);
and U11476 (N_11476,N_10759,N_11101);
or U11477 (N_11477,N_11141,N_10922);
nand U11478 (N_11478,N_10959,N_11052);
nand U11479 (N_11479,N_10975,N_11154);
nand U11480 (N_11480,N_10942,N_10776);
or U11481 (N_11481,N_10708,N_10929);
xor U11482 (N_11482,N_10784,N_10571);
nor U11483 (N_11483,N_10762,N_10919);
or U11484 (N_11484,N_10834,N_10914);
and U11485 (N_11485,N_11011,N_10613);
xor U11486 (N_11486,N_10660,N_11184);
nor U11487 (N_11487,N_10736,N_11083);
nand U11488 (N_11488,N_10793,N_10927);
nand U11489 (N_11489,N_10542,N_10886);
or U11490 (N_11490,N_10926,N_10963);
nand U11491 (N_11491,N_11028,N_10787);
nand U11492 (N_11492,N_11064,N_10537);
nand U11493 (N_11493,N_10771,N_10967);
and U11494 (N_11494,N_10545,N_11018);
and U11495 (N_11495,N_11061,N_11099);
nor U11496 (N_11496,N_11140,N_10648);
and U11497 (N_11497,N_10643,N_11056);
nand U11498 (N_11498,N_10651,N_10860);
and U11499 (N_11499,N_10645,N_10669);
xnor U11500 (N_11500,N_10714,N_11228);
and U11501 (N_11501,N_11232,N_10815);
or U11502 (N_11502,N_10740,N_10830);
or U11503 (N_11503,N_10950,N_11014);
nand U11504 (N_11504,N_11120,N_10607);
xor U11505 (N_11505,N_10567,N_10760);
nor U11506 (N_11506,N_10953,N_10579);
xor U11507 (N_11507,N_10530,N_10949);
nand U11508 (N_11508,N_11145,N_11249);
or U11509 (N_11509,N_10605,N_10867);
nor U11510 (N_11510,N_10546,N_10989);
and U11511 (N_11511,N_10848,N_11075);
xnor U11512 (N_11512,N_11158,N_10996);
nor U11513 (N_11513,N_11035,N_10732);
xnor U11514 (N_11514,N_10575,N_10974);
nand U11515 (N_11515,N_10774,N_10503);
and U11516 (N_11516,N_10980,N_10698);
xor U11517 (N_11517,N_10853,N_10968);
nor U11518 (N_11518,N_11019,N_11108);
nand U11519 (N_11519,N_11015,N_10670);
nor U11520 (N_11520,N_10722,N_11210);
or U11521 (N_11521,N_10928,N_10866);
xnor U11522 (N_11522,N_11199,N_10710);
nand U11523 (N_11523,N_11034,N_10677);
and U11524 (N_11524,N_10739,N_11146);
nand U11525 (N_11525,N_10882,N_11007);
or U11526 (N_11526,N_11006,N_10944);
nor U11527 (N_11527,N_11205,N_11125);
nand U11528 (N_11528,N_11113,N_10702);
nor U11529 (N_11529,N_10664,N_11086);
xnor U11530 (N_11530,N_11085,N_10568);
nor U11531 (N_11531,N_10855,N_10614);
and U11532 (N_11532,N_11058,N_11137);
nor U11533 (N_11533,N_10561,N_11181);
and U11534 (N_11534,N_11231,N_10981);
or U11535 (N_11535,N_11133,N_10653);
nand U11536 (N_11536,N_11033,N_10687);
or U11537 (N_11537,N_10918,N_10667);
or U11538 (N_11538,N_10534,N_11219);
or U11539 (N_11539,N_10749,N_10640);
and U11540 (N_11540,N_10587,N_11080);
nor U11541 (N_11541,N_10637,N_10540);
nor U11542 (N_11542,N_10631,N_10889);
or U11543 (N_11543,N_11215,N_10884);
nor U11544 (N_11544,N_10854,N_11221);
nand U11545 (N_11545,N_11176,N_10930);
and U11546 (N_11546,N_11139,N_11074);
and U11547 (N_11547,N_11102,N_10618);
nor U11548 (N_11548,N_11226,N_10656);
nor U11549 (N_11549,N_10500,N_10872);
nor U11550 (N_11550,N_10598,N_11223);
nor U11551 (N_11551,N_10887,N_10810);
nand U11552 (N_11552,N_10801,N_10785);
nand U11553 (N_11553,N_11020,N_10675);
and U11554 (N_11554,N_10745,N_10792);
and U11555 (N_11555,N_10816,N_10510);
and U11556 (N_11556,N_11057,N_10973);
or U11557 (N_11557,N_11066,N_11053);
or U11558 (N_11558,N_10720,N_11202);
and U11559 (N_11559,N_10580,N_10666);
nor U11560 (N_11560,N_11100,N_10986);
nand U11561 (N_11561,N_10589,N_10600);
nor U11562 (N_11562,N_11050,N_10582);
nand U11563 (N_11563,N_11172,N_11217);
or U11564 (N_11564,N_10738,N_11111);
nor U11565 (N_11565,N_10742,N_10715);
xnor U11566 (N_11566,N_10707,N_10501);
and U11567 (N_11567,N_11016,N_11045);
nor U11568 (N_11568,N_10719,N_11164);
nand U11569 (N_11569,N_10766,N_11010);
nor U11570 (N_11570,N_11094,N_10852);
nand U11571 (N_11571,N_10663,N_11079);
nor U11572 (N_11572,N_11091,N_10523);
and U11573 (N_11573,N_10721,N_10585);
and U11574 (N_11574,N_11055,N_11222);
or U11575 (N_11575,N_11051,N_11245);
nand U11576 (N_11576,N_11044,N_11022);
and U11577 (N_11577,N_11122,N_10671);
or U11578 (N_11578,N_11203,N_10642);
and U11579 (N_11579,N_11247,N_11127);
nand U11580 (N_11580,N_10890,N_10717);
and U11581 (N_11581,N_10502,N_10945);
nand U11582 (N_11582,N_11087,N_10676);
and U11583 (N_11583,N_11031,N_10900);
xor U11584 (N_11584,N_10606,N_10795);
nand U11585 (N_11585,N_10892,N_10622);
or U11586 (N_11586,N_10812,N_10610);
and U11587 (N_11587,N_10824,N_10796);
nor U11588 (N_11588,N_11142,N_10829);
or U11589 (N_11589,N_11167,N_10811);
nor U11590 (N_11590,N_10599,N_10630);
nand U11591 (N_11591,N_10856,N_11009);
nor U11592 (N_11592,N_10556,N_10902);
or U11593 (N_11593,N_10743,N_10513);
and U11594 (N_11594,N_10988,N_10800);
xor U11595 (N_11595,N_10746,N_10641);
and U11596 (N_11596,N_11151,N_10997);
nor U11597 (N_11597,N_10994,N_10861);
or U11598 (N_11598,N_10769,N_10689);
and U11599 (N_11599,N_10770,N_10564);
nand U11600 (N_11600,N_11240,N_10624);
nand U11601 (N_11601,N_10678,N_11043);
or U11602 (N_11602,N_10960,N_10790);
nor U11603 (N_11603,N_11212,N_11084);
nor U11604 (N_11604,N_10626,N_10807);
or U11605 (N_11605,N_11157,N_11230);
or U11606 (N_11606,N_11098,N_11163);
and U11607 (N_11607,N_10621,N_10697);
or U11608 (N_11608,N_10840,N_10976);
or U11609 (N_11609,N_11148,N_10565);
nand U11610 (N_11610,N_10750,N_11118);
xor U11611 (N_11611,N_11026,N_10685);
or U11612 (N_11612,N_11038,N_10874);
nand U11613 (N_11613,N_11209,N_11162);
or U11614 (N_11614,N_11126,N_11193);
nor U11615 (N_11615,N_10911,N_10794);
nor U11616 (N_11616,N_10778,N_10881);
nand U11617 (N_11617,N_11092,N_10910);
nand U11618 (N_11618,N_11081,N_10706);
xor U11619 (N_11619,N_10849,N_10566);
nor U11620 (N_11620,N_10533,N_10590);
nor U11621 (N_11621,N_10741,N_11224);
xor U11622 (N_11622,N_10609,N_11171);
nand U11623 (N_11623,N_11000,N_11144);
or U11624 (N_11624,N_11082,N_10573);
nand U11625 (N_11625,N_11211,N_10670);
and U11626 (N_11626,N_10883,N_11041);
and U11627 (N_11627,N_10963,N_11206);
nor U11628 (N_11628,N_11091,N_10685);
and U11629 (N_11629,N_10736,N_11174);
nand U11630 (N_11630,N_10644,N_10531);
nor U11631 (N_11631,N_10749,N_10940);
xnor U11632 (N_11632,N_10610,N_10842);
and U11633 (N_11633,N_11015,N_11016);
and U11634 (N_11634,N_10504,N_11003);
nand U11635 (N_11635,N_10901,N_10743);
and U11636 (N_11636,N_10529,N_10885);
and U11637 (N_11637,N_10716,N_11026);
nor U11638 (N_11638,N_11087,N_10742);
xor U11639 (N_11639,N_10500,N_10868);
or U11640 (N_11640,N_10712,N_10550);
or U11641 (N_11641,N_11043,N_10799);
and U11642 (N_11642,N_11149,N_10691);
nor U11643 (N_11643,N_10750,N_10539);
xor U11644 (N_11644,N_11104,N_10712);
xnor U11645 (N_11645,N_10671,N_11182);
xnor U11646 (N_11646,N_11115,N_10740);
nor U11647 (N_11647,N_10978,N_11170);
nand U11648 (N_11648,N_11230,N_11113);
or U11649 (N_11649,N_10579,N_11137);
xnor U11650 (N_11650,N_11056,N_10842);
nand U11651 (N_11651,N_10981,N_10802);
nor U11652 (N_11652,N_11199,N_10518);
nand U11653 (N_11653,N_10987,N_10780);
xor U11654 (N_11654,N_11129,N_11057);
nand U11655 (N_11655,N_10820,N_10961);
or U11656 (N_11656,N_10637,N_11169);
nand U11657 (N_11657,N_11015,N_10960);
xnor U11658 (N_11658,N_10660,N_10741);
and U11659 (N_11659,N_10869,N_10703);
nor U11660 (N_11660,N_11229,N_10669);
or U11661 (N_11661,N_10980,N_10731);
and U11662 (N_11662,N_10632,N_10746);
or U11663 (N_11663,N_11156,N_11053);
or U11664 (N_11664,N_11233,N_10998);
or U11665 (N_11665,N_10753,N_10720);
or U11666 (N_11666,N_11068,N_10965);
or U11667 (N_11667,N_10694,N_10711);
and U11668 (N_11668,N_11045,N_10931);
and U11669 (N_11669,N_10918,N_11011);
or U11670 (N_11670,N_10968,N_10897);
xor U11671 (N_11671,N_11215,N_10636);
and U11672 (N_11672,N_10672,N_10910);
xnor U11673 (N_11673,N_10803,N_10583);
nand U11674 (N_11674,N_11181,N_10843);
nor U11675 (N_11675,N_10911,N_10524);
or U11676 (N_11676,N_10718,N_11169);
or U11677 (N_11677,N_10800,N_11063);
nand U11678 (N_11678,N_10584,N_11089);
or U11679 (N_11679,N_10937,N_10887);
and U11680 (N_11680,N_10975,N_11084);
and U11681 (N_11681,N_11132,N_11236);
xnor U11682 (N_11682,N_10725,N_10777);
nor U11683 (N_11683,N_10563,N_11191);
or U11684 (N_11684,N_10620,N_11186);
nor U11685 (N_11685,N_11137,N_10661);
nor U11686 (N_11686,N_10817,N_10553);
or U11687 (N_11687,N_11204,N_10982);
or U11688 (N_11688,N_11074,N_10852);
nand U11689 (N_11689,N_10999,N_10642);
xnor U11690 (N_11690,N_10551,N_10535);
nand U11691 (N_11691,N_10953,N_10880);
and U11692 (N_11692,N_11235,N_10808);
nor U11693 (N_11693,N_11089,N_10758);
nor U11694 (N_11694,N_10728,N_10664);
and U11695 (N_11695,N_11151,N_10957);
nor U11696 (N_11696,N_10895,N_11145);
nor U11697 (N_11697,N_10897,N_11127);
nor U11698 (N_11698,N_11070,N_10997);
and U11699 (N_11699,N_11064,N_10841);
nand U11700 (N_11700,N_10579,N_10500);
and U11701 (N_11701,N_11043,N_11207);
xor U11702 (N_11702,N_10662,N_10686);
nand U11703 (N_11703,N_11047,N_10800);
and U11704 (N_11704,N_10788,N_10651);
xnor U11705 (N_11705,N_10632,N_10666);
nand U11706 (N_11706,N_10564,N_11053);
or U11707 (N_11707,N_10631,N_10870);
nor U11708 (N_11708,N_10582,N_10688);
nand U11709 (N_11709,N_10708,N_10962);
nand U11710 (N_11710,N_10552,N_11124);
and U11711 (N_11711,N_10685,N_11205);
or U11712 (N_11712,N_10964,N_11085);
and U11713 (N_11713,N_10636,N_10508);
and U11714 (N_11714,N_11046,N_10672);
nor U11715 (N_11715,N_11193,N_10520);
or U11716 (N_11716,N_11057,N_11181);
and U11717 (N_11717,N_11095,N_10542);
or U11718 (N_11718,N_10782,N_10678);
nor U11719 (N_11719,N_10623,N_10861);
or U11720 (N_11720,N_10568,N_10642);
and U11721 (N_11721,N_10527,N_10941);
or U11722 (N_11722,N_11133,N_11060);
xor U11723 (N_11723,N_11224,N_10665);
or U11724 (N_11724,N_10658,N_10530);
nor U11725 (N_11725,N_10579,N_10833);
or U11726 (N_11726,N_11079,N_10871);
and U11727 (N_11727,N_10700,N_10627);
nand U11728 (N_11728,N_10607,N_11030);
or U11729 (N_11729,N_10598,N_10865);
or U11730 (N_11730,N_10960,N_10557);
nor U11731 (N_11731,N_10824,N_10514);
nand U11732 (N_11732,N_11234,N_10917);
or U11733 (N_11733,N_11006,N_11109);
or U11734 (N_11734,N_10520,N_11089);
nand U11735 (N_11735,N_11239,N_10627);
nand U11736 (N_11736,N_10931,N_10739);
nor U11737 (N_11737,N_11170,N_10877);
or U11738 (N_11738,N_11084,N_10730);
and U11739 (N_11739,N_11121,N_10929);
nor U11740 (N_11740,N_10827,N_10655);
nand U11741 (N_11741,N_11029,N_11028);
or U11742 (N_11742,N_10634,N_10588);
nand U11743 (N_11743,N_10893,N_10766);
and U11744 (N_11744,N_10507,N_11188);
nand U11745 (N_11745,N_10940,N_10797);
and U11746 (N_11746,N_11176,N_10877);
and U11747 (N_11747,N_10655,N_10958);
or U11748 (N_11748,N_11129,N_10834);
or U11749 (N_11749,N_11126,N_11222);
or U11750 (N_11750,N_10776,N_10775);
nor U11751 (N_11751,N_10966,N_10731);
and U11752 (N_11752,N_11229,N_11163);
and U11753 (N_11753,N_11049,N_10881);
nor U11754 (N_11754,N_10849,N_11070);
nand U11755 (N_11755,N_11199,N_10552);
or U11756 (N_11756,N_10592,N_11124);
nor U11757 (N_11757,N_10659,N_10949);
and U11758 (N_11758,N_10677,N_10971);
or U11759 (N_11759,N_11047,N_11060);
or U11760 (N_11760,N_10674,N_11144);
nand U11761 (N_11761,N_10970,N_11100);
or U11762 (N_11762,N_11191,N_11074);
xnor U11763 (N_11763,N_10791,N_10999);
nor U11764 (N_11764,N_11117,N_11238);
xnor U11765 (N_11765,N_10669,N_10737);
and U11766 (N_11766,N_10532,N_11069);
and U11767 (N_11767,N_10624,N_11227);
and U11768 (N_11768,N_10567,N_10923);
nor U11769 (N_11769,N_10916,N_10826);
and U11770 (N_11770,N_10625,N_10826);
xor U11771 (N_11771,N_11026,N_10746);
nor U11772 (N_11772,N_10907,N_10893);
xor U11773 (N_11773,N_10948,N_11164);
nand U11774 (N_11774,N_11179,N_10538);
nand U11775 (N_11775,N_10932,N_10829);
nor U11776 (N_11776,N_10954,N_11081);
nand U11777 (N_11777,N_10634,N_10507);
nor U11778 (N_11778,N_10658,N_10984);
nand U11779 (N_11779,N_11024,N_11215);
xor U11780 (N_11780,N_10912,N_11023);
xnor U11781 (N_11781,N_11114,N_11190);
nor U11782 (N_11782,N_11138,N_10900);
and U11783 (N_11783,N_10530,N_10917);
nand U11784 (N_11784,N_11042,N_10951);
nand U11785 (N_11785,N_11207,N_11087);
xor U11786 (N_11786,N_10796,N_10758);
nand U11787 (N_11787,N_10694,N_10910);
nand U11788 (N_11788,N_10766,N_10571);
nand U11789 (N_11789,N_10996,N_10533);
and U11790 (N_11790,N_10596,N_11040);
and U11791 (N_11791,N_10754,N_11039);
nand U11792 (N_11792,N_11059,N_10928);
xor U11793 (N_11793,N_11077,N_10988);
nor U11794 (N_11794,N_11217,N_11179);
nor U11795 (N_11795,N_10720,N_10669);
or U11796 (N_11796,N_10969,N_10776);
and U11797 (N_11797,N_10593,N_10668);
or U11798 (N_11798,N_11002,N_11035);
and U11799 (N_11799,N_10625,N_10638);
nor U11800 (N_11800,N_11114,N_10532);
nor U11801 (N_11801,N_10986,N_10530);
nand U11802 (N_11802,N_10726,N_10937);
and U11803 (N_11803,N_10527,N_10823);
nand U11804 (N_11804,N_10854,N_10866);
nor U11805 (N_11805,N_11238,N_11184);
nor U11806 (N_11806,N_10815,N_11063);
nand U11807 (N_11807,N_10527,N_11091);
nor U11808 (N_11808,N_10911,N_11219);
or U11809 (N_11809,N_10813,N_10647);
or U11810 (N_11810,N_10789,N_11097);
nor U11811 (N_11811,N_10809,N_11104);
or U11812 (N_11812,N_10830,N_10936);
nor U11813 (N_11813,N_10846,N_11202);
or U11814 (N_11814,N_11238,N_11085);
nand U11815 (N_11815,N_10571,N_10782);
nor U11816 (N_11816,N_10956,N_10920);
xor U11817 (N_11817,N_10979,N_11173);
nor U11818 (N_11818,N_10746,N_10680);
nand U11819 (N_11819,N_11211,N_10985);
nand U11820 (N_11820,N_11005,N_10937);
or U11821 (N_11821,N_10854,N_11211);
and U11822 (N_11822,N_11039,N_10577);
xor U11823 (N_11823,N_11066,N_11219);
and U11824 (N_11824,N_11213,N_10780);
nand U11825 (N_11825,N_10566,N_10965);
nand U11826 (N_11826,N_10562,N_10823);
and U11827 (N_11827,N_10753,N_10926);
nand U11828 (N_11828,N_10822,N_10842);
nand U11829 (N_11829,N_10942,N_11065);
nand U11830 (N_11830,N_10823,N_11057);
nor U11831 (N_11831,N_10621,N_10720);
or U11832 (N_11832,N_10602,N_11005);
nor U11833 (N_11833,N_10871,N_10703);
nor U11834 (N_11834,N_10712,N_10949);
or U11835 (N_11835,N_10645,N_10767);
and U11836 (N_11836,N_10943,N_10504);
nand U11837 (N_11837,N_10852,N_11243);
xor U11838 (N_11838,N_10767,N_10567);
or U11839 (N_11839,N_11099,N_10516);
and U11840 (N_11840,N_10881,N_11210);
or U11841 (N_11841,N_11011,N_11015);
or U11842 (N_11842,N_11030,N_10630);
and U11843 (N_11843,N_10881,N_11085);
or U11844 (N_11844,N_10913,N_11098);
nor U11845 (N_11845,N_10787,N_10933);
and U11846 (N_11846,N_11144,N_10787);
xor U11847 (N_11847,N_10702,N_10508);
nand U11848 (N_11848,N_10653,N_10609);
xor U11849 (N_11849,N_10751,N_10760);
nor U11850 (N_11850,N_10819,N_10883);
nor U11851 (N_11851,N_11214,N_11192);
and U11852 (N_11852,N_10972,N_11071);
nor U11853 (N_11853,N_10786,N_11111);
nand U11854 (N_11854,N_10736,N_10918);
or U11855 (N_11855,N_11125,N_10635);
nand U11856 (N_11856,N_10674,N_10712);
xor U11857 (N_11857,N_11041,N_10929);
nand U11858 (N_11858,N_11089,N_10945);
nor U11859 (N_11859,N_11130,N_10631);
nor U11860 (N_11860,N_11116,N_10714);
or U11861 (N_11861,N_10653,N_10930);
or U11862 (N_11862,N_11113,N_11239);
nand U11863 (N_11863,N_11110,N_10576);
and U11864 (N_11864,N_10854,N_10859);
xor U11865 (N_11865,N_11070,N_10759);
xor U11866 (N_11866,N_11029,N_11173);
and U11867 (N_11867,N_10867,N_11194);
or U11868 (N_11868,N_11054,N_10710);
and U11869 (N_11869,N_11225,N_10526);
nand U11870 (N_11870,N_10606,N_11177);
nand U11871 (N_11871,N_10722,N_11016);
nand U11872 (N_11872,N_10599,N_10836);
or U11873 (N_11873,N_10726,N_10574);
or U11874 (N_11874,N_11202,N_10635);
or U11875 (N_11875,N_11007,N_10783);
nor U11876 (N_11876,N_11040,N_10747);
or U11877 (N_11877,N_10589,N_11051);
xor U11878 (N_11878,N_10569,N_11064);
and U11879 (N_11879,N_11236,N_10648);
and U11880 (N_11880,N_10967,N_11122);
and U11881 (N_11881,N_11198,N_11065);
xor U11882 (N_11882,N_10950,N_10906);
and U11883 (N_11883,N_10881,N_11186);
nand U11884 (N_11884,N_11068,N_11021);
nand U11885 (N_11885,N_10782,N_10888);
nor U11886 (N_11886,N_11166,N_10841);
nand U11887 (N_11887,N_10894,N_11050);
nand U11888 (N_11888,N_10668,N_11142);
nand U11889 (N_11889,N_11139,N_11247);
nand U11890 (N_11890,N_11100,N_11151);
or U11891 (N_11891,N_10754,N_10528);
or U11892 (N_11892,N_10873,N_10724);
nand U11893 (N_11893,N_10584,N_10954);
xnor U11894 (N_11894,N_11118,N_10862);
or U11895 (N_11895,N_10552,N_10896);
nor U11896 (N_11896,N_11035,N_11238);
and U11897 (N_11897,N_10852,N_11090);
nor U11898 (N_11898,N_11150,N_10999);
or U11899 (N_11899,N_11029,N_10783);
and U11900 (N_11900,N_10850,N_10928);
nor U11901 (N_11901,N_10578,N_10944);
and U11902 (N_11902,N_11124,N_10782);
xnor U11903 (N_11903,N_11072,N_10650);
and U11904 (N_11904,N_10704,N_10650);
or U11905 (N_11905,N_11223,N_11024);
or U11906 (N_11906,N_10939,N_11242);
or U11907 (N_11907,N_11052,N_11249);
nand U11908 (N_11908,N_10781,N_10897);
nor U11909 (N_11909,N_11212,N_11191);
nand U11910 (N_11910,N_10675,N_11081);
nor U11911 (N_11911,N_10630,N_11240);
nor U11912 (N_11912,N_11001,N_10854);
nor U11913 (N_11913,N_11000,N_10561);
nand U11914 (N_11914,N_10907,N_10715);
nand U11915 (N_11915,N_11029,N_10888);
nand U11916 (N_11916,N_11227,N_10739);
or U11917 (N_11917,N_11143,N_10623);
nor U11918 (N_11918,N_10941,N_10559);
and U11919 (N_11919,N_11147,N_10984);
and U11920 (N_11920,N_11049,N_10589);
nor U11921 (N_11921,N_10568,N_10808);
or U11922 (N_11922,N_11169,N_11171);
nand U11923 (N_11923,N_10998,N_10929);
nand U11924 (N_11924,N_10809,N_10542);
xor U11925 (N_11925,N_11242,N_10605);
xnor U11926 (N_11926,N_10985,N_11207);
nor U11927 (N_11927,N_11225,N_10842);
and U11928 (N_11928,N_10657,N_10546);
or U11929 (N_11929,N_10751,N_10548);
and U11930 (N_11930,N_10753,N_10638);
nor U11931 (N_11931,N_11218,N_10683);
nor U11932 (N_11932,N_10900,N_11072);
and U11933 (N_11933,N_11039,N_10602);
nand U11934 (N_11934,N_10910,N_10803);
xnor U11935 (N_11935,N_10803,N_11202);
and U11936 (N_11936,N_11135,N_10627);
nand U11937 (N_11937,N_10852,N_10677);
nor U11938 (N_11938,N_10953,N_11168);
or U11939 (N_11939,N_10927,N_11036);
or U11940 (N_11940,N_10855,N_10821);
nor U11941 (N_11941,N_10916,N_10787);
or U11942 (N_11942,N_10810,N_10963);
xnor U11943 (N_11943,N_10776,N_11157);
nor U11944 (N_11944,N_10797,N_10513);
or U11945 (N_11945,N_10619,N_10599);
nor U11946 (N_11946,N_10934,N_10993);
nor U11947 (N_11947,N_10557,N_10729);
nand U11948 (N_11948,N_11205,N_10750);
or U11949 (N_11949,N_10811,N_11014);
or U11950 (N_11950,N_10615,N_10990);
nor U11951 (N_11951,N_10963,N_10741);
and U11952 (N_11952,N_10886,N_10597);
nor U11953 (N_11953,N_11041,N_11030);
nor U11954 (N_11954,N_11104,N_11042);
or U11955 (N_11955,N_10758,N_10514);
nand U11956 (N_11956,N_10753,N_10704);
nor U11957 (N_11957,N_11232,N_10891);
xor U11958 (N_11958,N_10576,N_10967);
nor U11959 (N_11959,N_10739,N_10954);
xnor U11960 (N_11960,N_10856,N_10957);
and U11961 (N_11961,N_10524,N_10688);
or U11962 (N_11962,N_11228,N_10839);
nand U11963 (N_11963,N_11010,N_10696);
or U11964 (N_11964,N_10814,N_10602);
or U11965 (N_11965,N_11181,N_11164);
nand U11966 (N_11966,N_11227,N_11060);
nand U11967 (N_11967,N_10726,N_10505);
nor U11968 (N_11968,N_10646,N_10508);
or U11969 (N_11969,N_10933,N_10843);
or U11970 (N_11970,N_10651,N_10525);
nand U11971 (N_11971,N_10503,N_11135);
nor U11972 (N_11972,N_10606,N_10504);
or U11973 (N_11973,N_10609,N_10632);
or U11974 (N_11974,N_11086,N_10833);
or U11975 (N_11975,N_11238,N_10990);
nand U11976 (N_11976,N_11164,N_10660);
or U11977 (N_11977,N_10961,N_10956);
or U11978 (N_11978,N_10780,N_11075);
nand U11979 (N_11979,N_10881,N_11061);
nand U11980 (N_11980,N_11152,N_10537);
or U11981 (N_11981,N_10784,N_10517);
nor U11982 (N_11982,N_11162,N_10562);
or U11983 (N_11983,N_10927,N_10672);
nor U11984 (N_11984,N_11079,N_10905);
nor U11985 (N_11985,N_11145,N_11084);
and U11986 (N_11986,N_11152,N_10624);
nor U11987 (N_11987,N_10613,N_11224);
and U11988 (N_11988,N_11218,N_10921);
nand U11989 (N_11989,N_10733,N_10724);
and U11990 (N_11990,N_10916,N_11221);
and U11991 (N_11991,N_10549,N_11196);
xnor U11992 (N_11992,N_11031,N_10642);
nor U11993 (N_11993,N_10846,N_10630);
or U11994 (N_11994,N_10512,N_10780);
xnor U11995 (N_11995,N_11156,N_10887);
xnor U11996 (N_11996,N_10852,N_10621);
xnor U11997 (N_11997,N_10900,N_10761);
nand U11998 (N_11998,N_10539,N_10740);
or U11999 (N_11999,N_10900,N_10984);
nor U12000 (N_12000,N_11810,N_11445);
or U12001 (N_12001,N_11809,N_11987);
xnor U12002 (N_12002,N_11819,N_11313);
nor U12003 (N_12003,N_11306,N_11264);
nand U12004 (N_12004,N_11553,N_11312);
nor U12005 (N_12005,N_11650,N_11356);
nor U12006 (N_12006,N_11652,N_11865);
nand U12007 (N_12007,N_11887,N_11271);
and U12008 (N_12008,N_11675,N_11354);
or U12009 (N_12009,N_11931,N_11431);
and U12010 (N_12010,N_11473,N_11903);
and U12011 (N_12011,N_11750,N_11404);
and U12012 (N_12012,N_11627,N_11712);
nand U12013 (N_12013,N_11827,N_11894);
nand U12014 (N_12014,N_11695,N_11623);
nand U12015 (N_12015,N_11564,N_11976);
xor U12016 (N_12016,N_11651,N_11765);
nand U12017 (N_12017,N_11807,N_11378);
or U12018 (N_12018,N_11337,N_11783);
nor U12019 (N_12019,N_11332,N_11520);
and U12020 (N_12020,N_11967,N_11983);
or U12021 (N_12021,N_11462,N_11492);
nor U12022 (N_12022,N_11577,N_11795);
or U12023 (N_12023,N_11624,N_11552);
or U12024 (N_12024,N_11329,N_11872);
and U12025 (N_12025,N_11396,N_11472);
and U12026 (N_12026,N_11294,N_11981);
or U12027 (N_12027,N_11679,N_11422);
nor U12028 (N_12028,N_11575,N_11517);
nand U12029 (N_12029,N_11657,N_11556);
or U12030 (N_12030,N_11979,N_11498);
nor U12031 (N_12031,N_11893,N_11779);
and U12032 (N_12032,N_11283,N_11767);
and U12033 (N_12033,N_11468,N_11834);
nor U12034 (N_12034,N_11358,N_11992);
nor U12035 (N_12035,N_11622,N_11371);
and U12036 (N_12036,N_11461,N_11847);
nand U12037 (N_12037,N_11547,N_11942);
and U12038 (N_12038,N_11697,N_11537);
or U12039 (N_12039,N_11780,N_11690);
nand U12040 (N_12040,N_11421,N_11427);
and U12041 (N_12041,N_11853,N_11781);
or U12042 (N_12042,N_11532,N_11459);
and U12043 (N_12043,N_11570,N_11866);
nor U12044 (N_12044,N_11331,N_11720);
or U12045 (N_12045,N_11543,N_11739);
or U12046 (N_12046,N_11822,N_11913);
nor U12047 (N_12047,N_11705,N_11310);
nor U12048 (N_12048,N_11545,N_11862);
nor U12049 (N_12049,N_11429,N_11911);
xor U12050 (N_12050,N_11996,N_11797);
or U12051 (N_12051,N_11565,N_11787);
or U12052 (N_12052,N_11633,N_11531);
and U12053 (N_12053,N_11724,N_11734);
nor U12054 (N_12054,N_11475,N_11267);
nand U12055 (N_12055,N_11261,N_11533);
or U12056 (N_12056,N_11938,N_11508);
and U12057 (N_12057,N_11770,N_11263);
and U12058 (N_12058,N_11602,N_11812);
and U12059 (N_12059,N_11694,N_11258);
or U12060 (N_12060,N_11684,N_11961);
and U12061 (N_12061,N_11325,N_11891);
nor U12062 (N_12062,N_11282,N_11832);
nor U12063 (N_12063,N_11447,N_11709);
and U12064 (N_12064,N_11398,N_11292);
or U12065 (N_12065,N_11688,N_11601);
nor U12066 (N_12066,N_11998,N_11732);
and U12067 (N_12067,N_11760,N_11661);
xnor U12068 (N_12068,N_11890,N_11450);
or U12069 (N_12069,N_11743,N_11405);
and U12070 (N_12070,N_11558,N_11848);
and U12071 (N_12071,N_11907,N_11859);
nor U12072 (N_12072,N_11791,N_11438);
and U12073 (N_12073,N_11265,N_11844);
nand U12074 (N_12074,N_11728,N_11719);
nand U12075 (N_12075,N_11756,N_11584);
xor U12076 (N_12076,N_11495,N_11999);
nand U12077 (N_12077,N_11776,N_11539);
and U12078 (N_12078,N_11933,N_11374);
xor U12079 (N_12079,N_11443,N_11334);
xnor U12080 (N_12080,N_11717,N_11453);
nor U12081 (N_12081,N_11595,N_11917);
nand U12082 (N_12082,N_11272,N_11746);
and U12083 (N_12083,N_11710,N_11723);
nand U12084 (N_12084,N_11617,N_11293);
nor U12085 (N_12085,N_11274,N_11660);
nor U12086 (N_12086,N_11658,N_11954);
and U12087 (N_12087,N_11278,N_11689);
nor U12088 (N_12088,N_11729,N_11649);
or U12089 (N_12089,N_11401,N_11796);
and U12090 (N_12090,N_11437,N_11359);
nor U12091 (N_12091,N_11388,N_11403);
and U12092 (N_12092,N_11351,N_11342);
nand U12093 (N_12093,N_11432,N_11480);
or U12094 (N_12094,N_11433,N_11350);
nand U12095 (N_12095,N_11386,N_11837);
or U12096 (N_12096,N_11380,N_11940);
and U12097 (N_12097,N_11395,N_11557);
or U12098 (N_12098,N_11586,N_11522);
nor U12099 (N_12099,N_11693,N_11687);
and U12100 (N_12100,N_11511,N_11730);
and U12101 (N_12101,N_11490,N_11944);
nor U12102 (N_12102,N_11927,N_11609);
nor U12103 (N_12103,N_11410,N_11659);
or U12104 (N_12104,N_11873,N_11250);
nand U12105 (N_12105,N_11766,N_11288);
or U12106 (N_12106,N_11471,N_11470);
or U12107 (N_12107,N_11731,N_11973);
nor U12108 (N_12108,N_11953,N_11618);
nand U12109 (N_12109,N_11528,N_11774);
and U12110 (N_12110,N_11527,N_11343);
nand U12111 (N_12111,N_11318,N_11928);
and U12112 (N_12112,N_11676,N_11497);
and U12113 (N_12113,N_11888,N_11482);
nor U12114 (N_12114,N_11467,N_11854);
or U12115 (N_12115,N_11727,N_11871);
nand U12116 (N_12116,N_11889,N_11786);
and U12117 (N_12117,N_11307,N_11408);
xor U12118 (N_12118,N_11266,N_11639);
nor U12119 (N_12119,N_11273,N_11711);
or U12120 (N_12120,N_11930,N_11270);
and U12121 (N_12121,N_11883,N_11785);
or U12122 (N_12122,N_11792,N_11458);
nor U12123 (N_12123,N_11745,N_11372);
or U12124 (N_12124,N_11773,N_11455);
nand U12125 (N_12125,N_11607,N_11858);
nand U12126 (N_12126,N_11424,N_11663);
nand U12127 (N_12127,N_11525,N_11985);
nor U12128 (N_12128,N_11524,N_11379);
or U12129 (N_12129,N_11302,N_11397);
and U12130 (N_12130,N_11852,N_11965);
nor U12131 (N_12131,N_11625,N_11608);
or U12132 (N_12132,N_11662,N_11841);
nor U12133 (N_12133,N_11665,N_11576);
nor U12134 (N_12134,N_11414,N_11777);
nor U12135 (N_12135,N_11778,N_11594);
nor U12136 (N_12136,N_11549,N_11604);
or U12137 (N_12137,N_11997,N_11389);
and U12138 (N_12138,N_11559,N_11925);
xnor U12139 (N_12139,N_11857,N_11934);
nor U12140 (N_12140,N_11835,N_11434);
nand U12141 (N_12141,N_11346,N_11707);
and U12142 (N_12142,N_11978,N_11571);
and U12143 (N_12143,N_11964,N_11896);
nand U12144 (N_12144,N_11631,N_11691);
xor U12145 (N_12145,N_11823,N_11700);
nand U12146 (N_12146,N_11301,N_11648);
nor U12147 (N_12147,N_11988,N_11817);
and U12148 (N_12148,N_11845,N_11790);
and U12149 (N_12149,N_11920,N_11674);
nor U12150 (N_12150,N_11647,N_11260);
or U12151 (N_12151,N_11441,N_11326);
nor U12152 (N_12152,N_11840,N_11642);
and U12153 (N_12153,N_11352,N_11824);
or U12154 (N_12154,N_11335,N_11534);
nor U12155 (N_12155,N_11514,N_11668);
and U12156 (N_12156,N_11451,N_11587);
nor U12157 (N_12157,N_11741,N_11400);
xnor U12158 (N_12158,N_11339,N_11360);
nand U12159 (N_12159,N_11805,N_11505);
and U12160 (N_12160,N_11982,N_11813);
nor U12161 (N_12161,N_11308,N_11753);
xor U12162 (N_12162,N_11995,N_11794);
nand U12163 (N_12163,N_11348,N_11503);
and U12164 (N_12164,N_11423,N_11507);
nand U12165 (N_12165,N_11875,N_11643);
and U12166 (N_12166,N_11755,N_11950);
or U12167 (N_12167,N_11521,N_11966);
nor U12168 (N_12168,N_11555,N_11276);
or U12169 (N_12169,N_11673,N_11828);
nor U12170 (N_12170,N_11744,N_11692);
xnor U12171 (N_12171,N_11603,N_11993);
nand U12172 (N_12172,N_11383,N_11365);
and U12173 (N_12173,N_11736,N_11653);
or U12174 (N_12174,N_11628,N_11415);
nor U12175 (N_12175,N_11962,N_11513);
nor U12176 (N_12176,N_11910,N_11580);
or U12177 (N_12177,N_11937,N_11821);
nand U12178 (N_12178,N_11990,N_11377);
nor U12179 (N_12179,N_11784,N_11314);
xor U12180 (N_12180,N_11892,N_11298);
nor U12181 (N_12181,N_11478,N_11678);
or U12182 (N_12182,N_11632,N_11818);
nand U12183 (N_12183,N_11814,N_11904);
and U12184 (N_12184,N_11884,N_11290);
nor U12185 (N_12185,N_11941,N_11958);
nor U12186 (N_12186,N_11926,N_11898);
xnor U12187 (N_12187,N_11936,N_11757);
nand U12188 (N_12188,N_11820,N_11672);
nand U12189 (N_12189,N_11991,N_11614);
and U12190 (N_12190,N_11304,N_11879);
xor U12191 (N_12191,N_11843,N_11929);
or U12192 (N_12192,N_11484,N_11634);
and U12193 (N_12193,N_11535,N_11519);
or U12194 (N_12194,N_11764,N_11959);
xor U12195 (N_12195,N_11782,N_11469);
and U12196 (N_12196,N_11749,N_11385);
or U12197 (N_12197,N_11563,N_11456);
xor U12198 (N_12198,N_11444,N_11680);
and U12199 (N_12199,N_11476,N_11322);
nor U12200 (N_12200,N_11948,N_11949);
or U12201 (N_12201,N_11567,N_11338);
or U12202 (N_12202,N_11994,N_11486);
nor U12203 (N_12203,N_11590,N_11568);
and U12204 (N_12204,N_11636,N_11426);
and U12205 (N_12205,N_11295,N_11804);
and U12206 (N_12206,N_11382,N_11952);
nor U12207 (N_12207,N_11353,N_11621);
xor U12208 (N_12208,N_11391,N_11986);
or U12209 (N_12209,N_11387,N_11772);
and U12210 (N_12210,N_11425,N_11542);
nand U12211 (N_12211,N_11921,N_11466);
nor U12212 (N_12212,N_11488,N_11375);
or U12213 (N_12213,N_11641,N_11251);
nand U12214 (N_12214,N_11368,N_11487);
nor U12215 (N_12215,N_11943,N_11955);
nand U12216 (N_12216,N_11611,N_11666);
xor U12217 (N_12217,N_11355,N_11698);
nand U12218 (N_12218,N_11912,N_11815);
xor U12219 (N_12219,N_11935,N_11561);
and U12220 (N_12220,N_11341,N_11579);
and U12221 (N_12221,N_11706,N_11256);
or U12222 (N_12222,N_11956,N_11864);
or U12223 (N_12223,N_11363,N_11446);
or U12224 (N_12224,N_11763,N_11914);
or U12225 (N_12225,N_11754,N_11578);
or U12226 (N_12226,N_11932,N_11860);
nor U12227 (N_12227,N_11855,N_11737);
xor U12228 (N_12228,N_11902,N_11394);
nand U12229 (N_12229,N_11646,N_11900);
and U12230 (N_12230,N_11253,N_11876);
nand U12231 (N_12231,N_11489,N_11257);
or U12232 (N_12232,N_11874,N_11340);
or U12233 (N_12233,N_11946,N_11554);
xor U12234 (N_12234,N_11849,N_11369);
or U12235 (N_12235,N_11742,N_11980);
or U12236 (N_12236,N_11589,N_11771);
nand U12237 (N_12237,N_11850,N_11515);
or U12238 (N_12238,N_11977,N_11886);
and U12239 (N_12239,N_11596,N_11619);
nor U12240 (N_12240,N_11867,N_11330);
nand U12241 (N_12241,N_11297,N_11440);
and U12242 (N_12242,N_11381,N_11530);
or U12243 (N_12243,N_11775,N_11877);
xor U12244 (N_12244,N_11504,N_11916);
nor U12245 (N_12245,N_11409,N_11494);
and U12246 (N_12246,N_11275,N_11262);
nor U12247 (N_12247,N_11905,N_11442);
nand U12248 (N_12248,N_11882,N_11918);
nand U12249 (N_12249,N_11605,N_11474);
or U12250 (N_12250,N_11726,N_11477);
nand U12251 (N_12251,N_11699,N_11960);
or U12252 (N_12252,N_11825,N_11529);
nor U12253 (N_12253,N_11670,N_11512);
xnor U12254 (N_12254,N_11357,N_11829);
nor U12255 (N_12255,N_11868,N_11816);
and U12256 (N_12256,N_11544,N_11550);
nor U12257 (N_12257,N_11838,N_11481);
nor U12258 (N_12258,N_11600,N_11523);
nand U12259 (N_12259,N_11291,N_11402);
nand U12260 (N_12260,N_11768,N_11656);
nand U12261 (N_12261,N_11345,N_11430);
or U12262 (N_12262,N_11572,N_11588);
nor U12263 (N_12263,N_11566,N_11501);
or U12264 (N_12264,N_11485,N_11573);
nand U12265 (N_12265,N_11317,N_11452);
or U12266 (N_12266,N_11491,N_11885);
or U12267 (N_12267,N_11897,N_11963);
nor U12268 (N_12268,N_11861,N_11808);
or U12269 (N_12269,N_11721,N_11702);
nand U12270 (N_12270,N_11610,N_11393);
or U12271 (N_12271,N_11616,N_11384);
nor U12272 (N_12272,N_11364,N_11915);
or U12273 (N_12273,N_11863,N_11412);
nand U12274 (N_12274,N_11683,N_11599);
xnor U12275 (N_12275,N_11418,N_11733);
xnor U12276 (N_12276,N_11947,N_11738);
xnor U12277 (N_12277,N_11793,N_11899);
nand U12278 (N_12278,N_11439,N_11655);
nor U12279 (N_12279,N_11671,N_11644);
nor U12280 (N_12280,N_11289,N_11972);
and U12281 (N_12281,N_11344,N_11957);
or U12282 (N_12282,N_11323,N_11349);
or U12283 (N_12283,N_11798,N_11831);
nor U12284 (N_12284,N_11895,N_11939);
or U12285 (N_12285,N_11309,N_11800);
nor U12286 (N_12286,N_11551,N_11637);
nand U12287 (N_12287,N_11613,N_11638);
and U12288 (N_12288,N_11399,N_11305);
or U12289 (N_12289,N_11316,N_11333);
or U12290 (N_12290,N_11436,N_11591);
or U12291 (N_12291,N_11851,N_11908);
and U12292 (N_12292,N_11984,N_11806);
or U12293 (N_12293,N_11615,N_11320);
nor U12294 (N_12294,N_11448,N_11255);
and U12295 (N_12295,N_11463,N_11361);
and U12296 (N_12296,N_11376,N_11465);
nor U12297 (N_12297,N_11716,N_11669);
and U12298 (N_12298,N_11923,N_11420);
and U12299 (N_12299,N_11725,N_11536);
nand U12300 (N_12300,N_11906,N_11285);
nand U12301 (N_12301,N_11681,N_11704);
nor U12302 (N_12302,N_11696,N_11502);
or U12303 (N_12303,N_11801,N_11703);
xor U12304 (N_12304,N_11626,N_11296);
and U12305 (N_12305,N_11259,N_11583);
nand U12306 (N_12306,N_11464,N_11975);
and U12307 (N_12307,N_11799,N_11924);
and U12308 (N_12308,N_11748,N_11518);
or U12309 (N_12309,N_11284,N_11449);
and U12310 (N_12310,N_11509,N_11336);
nand U12311 (N_12311,N_11803,N_11880);
or U12312 (N_12312,N_11826,N_11560);
and U12313 (N_12313,N_11496,N_11759);
nand U12314 (N_12314,N_11390,N_11321);
nor U12315 (N_12315,N_11546,N_11856);
nand U12316 (N_12316,N_11416,N_11752);
and U12317 (N_12317,N_11367,N_11833);
and U12318 (N_12318,N_11582,N_11319);
nand U12319 (N_12319,N_11254,N_11645);
xor U12320 (N_12320,N_11919,N_11846);
and U12321 (N_12321,N_11802,N_11878);
nor U12322 (N_12322,N_11324,N_11277);
and U12323 (N_12323,N_11901,N_11612);
and U12324 (N_12324,N_11406,N_11479);
or U12325 (N_12325,N_11969,N_11686);
nand U12326 (N_12326,N_11677,N_11735);
xor U12327 (N_12327,N_11842,N_11635);
and U12328 (N_12328,N_11722,N_11280);
nand U12329 (N_12329,N_11548,N_11909);
or U12330 (N_12330,N_11606,N_11870);
nand U12331 (N_12331,N_11685,N_11510);
or U12332 (N_12332,N_11493,N_11300);
nand U12333 (N_12333,N_11373,N_11788);
or U12334 (N_12334,N_11968,N_11411);
xnor U12335 (N_12335,N_11714,N_11881);
or U12336 (N_12336,N_11279,N_11740);
nor U12337 (N_12337,N_11974,N_11419);
nor U12338 (N_12338,N_11362,N_11597);
xor U12339 (N_12339,N_11407,N_11789);
and U12340 (N_12340,N_11581,N_11989);
and U12341 (N_12341,N_11598,N_11311);
nand U12342 (N_12342,N_11413,N_11328);
nor U12343 (N_12343,N_11435,N_11417);
or U12344 (N_12344,N_11569,N_11315);
xnor U12345 (N_12345,N_11869,N_11327);
or U12346 (N_12346,N_11747,N_11281);
nand U12347 (N_12347,N_11971,N_11839);
nor U12348 (N_12348,N_11713,N_11299);
nand U12349 (N_12349,N_11366,N_11836);
nand U12350 (N_12350,N_11347,N_11460);
nor U12351 (N_12351,N_11667,N_11252);
or U12352 (N_12352,N_11428,N_11303);
or U12353 (N_12353,N_11682,N_11830);
xor U12354 (N_12354,N_11945,N_11286);
nand U12355 (N_12355,N_11392,N_11701);
nand U12356 (N_12356,N_11499,N_11269);
and U12357 (N_12357,N_11457,N_11592);
or U12358 (N_12358,N_11287,N_11506);
xnor U12359 (N_12359,N_11540,N_11715);
and U12360 (N_12360,N_11574,N_11708);
nor U12361 (N_12361,N_11483,N_11922);
or U12362 (N_12362,N_11762,N_11370);
or U12363 (N_12363,N_11268,N_11811);
and U12364 (N_12364,N_11654,N_11526);
nor U12365 (N_12365,N_11718,N_11593);
nor U12366 (N_12366,N_11761,N_11640);
nor U12367 (N_12367,N_11585,N_11951);
nand U12368 (N_12368,N_11630,N_11769);
or U12369 (N_12369,N_11500,N_11541);
or U12370 (N_12370,N_11751,N_11620);
nand U12371 (N_12371,N_11629,N_11516);
and U12372 (N_12372,N_11970,N_11758);
or U12373 (N_12373,N_11664,N_11562);
and U12374 (N_12374,N_11538,N_11454);
xnor U12375 (N_12375,N_11744,N_11418);
and U12376 (N_12376,N_11372,N_11625);
nor U12377 (N_12377,N_11998,N_11408);
xor U12378 (N_12378,N_11551,N_11523);
and U12379 (N_12379,N_11541,N_11972);
and U12380 (N_12380,N_11462,N_11968);
xnor U12381 (N_12381,N_11958,N_11738);
or U12382 (N_12382,N_11378,N_11251);
and U12383 (N_12383,N_11622,N_11649);
or U12384 (N_12384,N_11697,N_11301);
or U12385 (N_12385,N_11889,N_11624);
xnor U12386 (N_12386,N_11807,N_11743);
or U12387 (N_12387,N_11327,N_11834);
or U12388 (N_12388,N_11588,N_11560);
and U12389 (N_12389,N_11713,N_11749);
or U12390 (N_12390,N_11520,N_11913);
nor U12391 (N_12391,N_11642,N_11333);
or U12392 (N_12392,N_11254,N_11801);
nor U12393 (N_12393,N_11644,N_11705);
nand U12394 (N_12394,N_11754,N_11539);
nor U12395 (N_12395,N_11400,N_11331);
xnor U12396 (N_12396,N_11650,N_11968);
xor U12397 (N_12397,N_11648,N_11842);
nor U12398 (N_12398,N_11685,N_11333);
nand U12399 (N_12399,N_11731,N_11318);
and U12400 (N_12400,N_11259,N_11275);
nand U12401 (N_12401,N_11595,N_11717);
nor U12402 (N_12402,N_11720,N_11354);
or U12403 (N_12403,N_11319,N_11279);
nand U12404 (N_12404,N_11574,N_11569);
nand U12405 (N_12405,N_11681,N_11341);
nor U12406 (N_12406,N_11843,N_11298);
nor U12407 (N_12407,N_11610,N_11639);
nor U12408 (N_12408,N_11616,N_11912);
nor U12409 (N_12409,N_11555,N_11778);
nand U12410 (N_12410,N_11986,N_11572);
nand U12411 (N_12411,N_11618,N_11252);
or U12412 (N_12412,N_11419,N_11672);
nand U12413 (N_12413,N_11445,N_11290);
or U12414 (N_12414,N_11563,N_11495);
and U12415 (N_12415,N_11485,N_11826);
or U12416 (N_12416,N_11464,N_11446);
nand U12417 (N_12417,N_11897,N_11626);
and U12418 (N_12418,N_11254,N_11250);
nand U12419 (N_12419,N_11272,N_11333);
and U12420 (N_12420,N_11858,N_11620);
and U12421 (N_12421,N_11562,N_11536);
and U12422 (N_12422,N_11629,N_11575);
nor U12423 (N_12423,N_11951,N_11656);
nor U12424 (N_12424,N_11948,N_11964);
nand U12425 (N_12425,N_11630,N_11794);
nand U12426 (N_12426,N_11254,N_11683);
nand U12427 (N_12427,N_11995,N_11473);
or U12428 (N_12428,N_11846,N_11309);
nand U12429 (N_12429,N_11861,N_11917);
nand U12430 (N_12430,N_11288,N_11779);
nor U12431 (N_12431,N_11445,N_11937);
or U12432 (N_12432,N_11272,N_11779);
nand U12433 (N_12433,N_11907,N_11819);
and U12434 (N_12434,N_11488,N_11789);
and U12435 (N_12435,N_11669,N_11682);
nor U12436 (N_12436,N_11764,N_11709);
nor U12437 (N_12437,N_11684,N_11595);
or U12438 (N_12438,N_11966,N_11286);
and U12439 (N_12439,N_11420,N_11809);
and U12440 (N_12440,N_11257,N_11629);
or U12441 (N_12441,N_11377,N_11888);
or U12442 (N_12442,N_11527,N_11335);
and U12443 (N_12443,N_11452,N_11928);
nor U12444 (N_12444,N_11839,N_11764);
xnor U12445 (N_12445,N_11798,N_11641);
nor U12446 (N_12446,N_11343,N_11858);
and U12447 (N_12447,N_11553,N_11756);
or U12448 (N_12448,N_11676,N_11993);
and U12449 (N_12449,N_11843,N_11918);
or U12450 (N_12450,N_11846,N_11739);
nand U12451 (N_12451,N_11914,N_11459);
nand U12452 (N_12452,N_11980,N_11971);
xor U12453 (N_12453,N_11468,N_11261);
and U12454 (N_12454,N_11682,N_11975);
nor U12455 (N_12455,N_11508,N_11568);
nand U12456 (N_12456,N_11741,N_11270);
and U12457 (N_12457,N_11602,N_11756);
nand U12458 (N_12458,N_11385,N_11531);
xor U12459 (N_12459,N_11970,N_11586);
xnor U12460 (N_12460,N_11372,N_11287);
and U12461 (N_12461,N_11370,N_11818);
and U12462 (N_12462,N_11401,N_11755);
nor U12463 (N_12463,N_11644,N_11376);
nand U12464 (N_12464,N_11629,N_11774);
nand U12465 (N_12465,N_11469,N_11831);
nand U12466 (N_12466,N_11452,N_11808);
or U12467 (N_12467,N_11968,N_11957);
or U12468 (N_12468,N_11255,N_11607);
and U12469 (N_12469,N_11940,N_11630);
or U12470 (N_12470,N_11921,N_11859);
or U12471 (N_12471,N_11318,N_11376);
xor U12472 (N_12472,N_11921,N_11517);
xnor U12473 (N_12473,N_11649,N_11713);
nand U12474 (N_12474,N_11642,N_11507);
xnor U12475 (N_12475,N_11540,N_11721);
or U12476 (N_12476,N_11597,N_11988);
and U12477 (N_12477,N_11739,N_11492);
nand U12478 (N_12478,N_11657,N_11934);
xor U12479 (N_12479,N_11699,N_11673);
and U12480 (N_12480,N_11535,N_11254);
nand U12481 (N_12481,N_11363,N_11281);
and U12482 (N_12482,N_11639,N_11555);
or U12483 (N_12483,N_11963,N_11852);
or U12484 (N_12484,N_11463,N_11304);
nand U12485 (N_12485,N_11382,N_11482);
or U12486 (N_12486,N_11423,N_11342);
or U12487 (N_12487,N_11913,N_11911);
nand U12488 (N_12488,N_11970,N_11672);
nand U12489 (N_12489,N_11502,N_11495);
nor U12490 (N_12490,N_11251,N_11566);
nand U12491 (N_12491,N_11623,N_11919);
and U12492 (N_12492,N_11668,N_11937);
nor U12493 (N_12493,N_11302,N_11496);
or U12494 (N_12494,N_11660,N_11294);
and U12495 (N_12495,N_11450,N_11477);
xor U12496 (N_12496,N_11669,N_11273);
nand U12497 (N_12497,N_11581,N_11347);
or U12498 (N_12498,N_11895,N_11962);
nand U12499 (N_12499,N_11705,N_11313);
xor U12500 (N_12500,N_11399,N_11594);
nand U12501 (N_12501,N_11643,N_11547);
nand U12502 (N_12502,N_11670,N_11658);
and U12503 (N_12503,N_11742,N_11434);
and U12504 (N_12504,N_11905,N_11254);
nor U12505 (N_12505,N_11958,N_11325);
nand U12506 (N_12506,N_11643,N_11803);
nand U12507 (N_12507,N_11863,N_11843);
nand U12508 (N_12508,N_11469,N_11444);
nor U12509 (N_12509,N_11458,N_11619);
nor U12510 (N_12510,N_11820,N_11576);
nand U12511 (N_12511,N_11593,N_11569);
and U12512 (N_12512,N_11350,N_11708);
xor U12513 (N_12513,N_11527,N_11732);
nor U12514 (N_12514,N_11680,N_11701);
nand U12515 (N_12515,N_11972,N_11814);
nor U12516 (N_12516,N_11564,N_11501);
nor U12517 (N_12517,N_11618,N_11375);
and U12518 (N_12518,N_11298,N_11419);
or U12519 (N_12519,N_11982,N_11596);
and U12520 (N_12520,N_11693,N_11868);
nor U12521 (N_12521,N_11913,N_11647);
and U12522 (N_12522,N_11732,N_11492);
nor U12523 (N_12523,N_11549,N_11278);
and U12524 (N_12524,N_11495,N_11828);
nand U12525 (N_12525,N_11835,N_11285);
nand U12526 (N_12526,N_11274,N_11962);
and U12527 (N_12527,N_11912,N_11832);
nand U12528 (N_12528,N_11571,N_11472);
nor U12529 (N_12529,N_11543,N_11565);
and U12530 (N_12530,N_11585,N_11390);
or U12531 (N_12531,N_11538,N_11257);
nand U12532 (N_12532,N_11410,N_11251);
nor U12533 (N_12533,N_11513,N_11611);
nor U12534 (N_12534,N_11535,N_11410);
xnor U12535 (N_12535,N_11370,N_11518);
nand U12536 (N_12536,N_11363,N_11934);
or U12537 (N_12537,N_11375,N_11661);
nor U12538 (N_12538,N_11428,N_11596);
nand U12539 (N_12539,N_11255,N_11650);
and U12540 (N_12540,N_11263,N_11304);
xnor U12541 (N_12541,N_11448,N_11603);
nor U12542 (N_12542,N_11259,N_11305);
nor U12543 (N_12543,N_11338,N_11900);
nor U12544 (N_12544,N_11948,N_11702);
and U12545 (N_12545,N_11543,N_11362);
nand U12546 (N_12546,N_11259,N_11635);
or U12547 (N_12547,N_11970,N_11489);
or U12548 (N_12548,N_11571,N_11622);
xnor U12549 (N_12549,N_11630,N_11297);
and U12550 (N_12550,N_11883,N_11904);
nand U12551 (N_12551,N_11449,N_11294);
or U12552 (N_12552,N_11772,N_11974);
nor U12553 (N_12553,N_11856,N_11305);
nand U12554 (N_12554,N_11683,N_11299);
nor U12555 (N_12555,N_11600,N_11507);
or U12556 (N_12556,N_11631,N_11304);
nand U12557 (N_12557,N_11331,N_11350);
nand U12558 (N_12558,N_11265,N_11330);
nor U12559 (N_12559,N_11960,N_11623);
or U12560 (N_12560,N_11823,N_11388);
nand U12561 (N_12561,N_11634,N_11967);
xnor U12562 (N_12562,N_11266,N_11724);
or U12563 (N_12563,N_11617,N_11971);
nor U12564 (N_12564,N_11402,N_11412);
or U12565 (N_12565,N_11449,N_11887);
or U12566 (N_12566,N_11466,N_11720);
and U12567 (N_12567,N_11458,N_11700);
nand U12568 (N_12568,N_11758,N_11620);
nor U12569 (N_12569,N_11770,N_11257);
nand U12570 (N_12570,N_11298,N_11361);
nor U12571 (N_12571,N_11566,N_11932);
nand U12572 (N_12572,N_11467,N_11435);
nand U12573 (N_12573,N_11278,N_11594);
or U12574 (N_12574,N_11785,N_11652);
or U12575 (N_12575,N_11834,N_11524);
xor U12576 (N_12576,N_11909,N_11433);
or U12577 (N_12577,N_11588,N_11795);
xnor U12578 (N_12578,N_11419,N_11429);
and U12579 (N_12579,N_11331,N_11518);
xor U12580 (N_12580,N_11268,N_11800);
xnor U12581 (N_12581,N_11452,N_11902);
nand U12582 (N_12582,N_11990,N_11743);
or U12583 (N_12583,N_11281,N_11389);
or U12584 (N_12584,N_11516,N_11495);
or U12585 (N_12585,N_11460,N_11976);
or U12586 (N_12586,N_11661,N_11573);
and U12587 (N_12587,N_11432,N_11897);
nand U12588 (N_12588,N_11405,N_11286);
nand U12589 (N_12589,N_11299,N_11977);
and U12590 (N_12590,N_11501,N_11437);
xor U12591 (N_12591,N_11704,N_11508);
nor U12592 (N_12592,N_11265,N_11487);
nand U12593 (N_12593,N_11593,N_11755);
nor U12594 (N_12594,N_11682,N_11568);
nand U12595 (N_12595,N_11538,N_11767);
or U12596 (N_12596,N_11926,N_11796);
and U12597 (N_12597,N_11932,N_11664);
and U12598 (N_12598,N_11445,N_11830);
nand U12599 (N_12599,N_11940,N_11511);
xnor U12600 (N_12600,N_11441,N_11672);
or U12601 (N_12601,N_11720,N_11965);
or U12602 (N_12602,N_11553,N_11262);
and U12603 (N_12603,N_11902,N_11399);
nor U12604 (N_12604,N_11262,N_11421);
xor U12605 (N_12605,N_11579,N_11647);
and U12606 (N_12606,N_11417,N_11433);
nand U12607 (N_12607,N_11252,N_11518);
nand U12608 (N_12608,N_11915,N_11349);
nor U12609 (N_12609,N_11284,N_11534);
nor U12610 (N_12610,N_11537,N_11422);
xor U12611 (N_12611,N_11286,N_11798);
and U12612 (N_12612,N_11738,N_11833);
or U12613 (N_12613,N_11689,N_11373);
and U12614 (N_12614,N_11444,N_11858);
xor U12615 (N_12615,N_11564,N_11259);
or U12616 (N_12616,N_11641,N_11693);
or U12617 (N_12617,N_11809,N_11292);
and U12618 (N_12618,N_11376,N_11631);
nand U12619 (N_12619,N_11880,N_11806);
nand U12620 (N_12620,N_11746,N_11700);
or U12621 (N_12621,N_11544,N_11760);
nand U12622 (N_12622,N_11819,N_11845);
xor U12623 (N_12623,N_11671,N_11869);
nand U12624 (N_12624,N_11273,N_11846);
xor U12625 (N_12625,N_11451,N_11642);
xor U12626 (N_12626,N_11682,N_11912);
and U12627 (N_12627,N_11402,N_11289);
nand U12628 (N_12628,N_11414,N_11615);
or U12629 (N_12629,N_11845,N_11536);
nor U12630 (N_12630,N_11302,N_11537);
nand U12631 (N_12631,N_11275,N_11680);
and U12632 (N_12632,N_11825,N_11747);
and U12633 (N_12633,N_11465,N_11257);
and U12634 (N_12634,N_11780,N_11304);
nand U12635 (N_12635,N_11858,N_11932);
and U12636 (N_12636,N_11572,N_11999);
nor U12637 (N_12637,N_11491,N_11808);
nor U12638 (N_12638,N_11477,N_11585);
nand U12639 (N_12639,N_11780,N_11480);
nor U12640 (N_12640,N_11939,N_11676);
nor U12641 (N_12641,N_11572,N_11810);
and U12642 (N_12642,N_11431,N_11765);
or U12643 (N_12643,N_11939,N_11418);
nand U12644 (N_12644,N_11545,N_11546);
nor U12645 (N_12645,N_11603,N_11535);
xnor U12646 (N_12646,N_11539,N_11308);
nand U12647 (N_12647,N_11356,N_11914);
and U12648 (N_12648,N_11829,N_11917);
xor U12649 (N_12649,N_11487,N_11351);
nand U12650 (N_12650,N_11264,N_11314);
nand U12651 (N_12651,N_11434,N_11926);
nor U12652 (N_12652,N_11569,N_11414);
xnor U12653 (N_12653,N_11917,N_11324);
nor U12654 (N_12654,N_11465,N_11721);
nor U12655 (N_12655,N_11562,N_11784);
nand U12656 (N_12656,N_11765,N_11840);
or U12657 (N_12657,N_11682,N_11862);
nor U12658 (N_12658,N_11326,N_11697);
or U12659 (N_12659,N_11328,N_11862);
nor U12660 (N_12660,N_11684,N_11612);
xnor U12661 (N_12661,N_11273,N_11959);
or U12662 (N_12662,N_11400,N_11265);
nor U12663 (N_12663,N_11388,N_11498);
nand U12664 (N_12664,N_11580,N_11835);
nand U12665 (N_12665,N_11587,N_11946);
or U12666 (N_12666,N_11749,N_11496);
nand U12667 (N_12667,N_11704,N_11439);
or U12668 (N_12668,N_11889,N_11614);
nor U12669 (N_12669,N_11492,N_11769);
and U12670 (N_12670,N_11764,N_11749);
xor U12671 (N_12671,N_11695,N_11611);
or U12672 (N_12672,N_11252,N_11731);
nor U12673 (N_12673,N_11692,N_11899);
and U12674 (N_12674,N_11319,N_11843);
and U12675 (N_12675,N_11520,N_11962);
nand U12676 (N_12676,N_11267,N_11839);
nand U12677 (N_12677,N_11637,N_11343);
and U12678 (N_12678,N_11599,N_11713);
nand U12679 (N_12679,N_11766,N_11811);
and U12680 (N_12680,N_11672,N_11515);
or U12681 (N_12681,N_11368,N_11829);
and U12682 (N_12682,N_11288,N_11355);
nor U12683 (N_12683,N_11485,N_11933);
or U12684 (N_12684,N_11684,N_11745);
or U12685 (N_12685,N_11886,N_11513);
nor U12686 (N_12686,N_11356,N_11577);
nor U12687 (N_12687,N_11880,N_11592);
nand U12688 (N_12688,N_11776,N_11866);
nand U12689 (N_12689,N_11277,N_11620);
nor U12690 (N_12690,N_11475,N_11854);
or U12691 (N_12691,N_11944,N_11668);
or U12692 (N_12692,N_11302,N_11777);
nor U12693 (N_12693,N_11295,N_11320);
xnor U12694 (N_12694,N_11306,N_11417);
nor U12695 (N_12695,N_11334,N_11920);
nor U12696 (N_12696,N_11496,N_11256);
and U12697 (N_12697,N_11451,N_11619);
xnor U12698 (N_12698,N_11641,N_11521);
nand U12699 (N_12699,N_11841,N_11681);
or U12700 (N_12700,N_11379,N_11496);
and U12701 (N_12701,N_11487,N_11300);
and U12702 (N_12702,N_11562,N_11773);
or U12703 (N_12703,N_11799,N_11774);
and U12704 (N_12704,N_11529,N_11753);
and U12705 (N_12705,N_11449,N_11572);
or U12706 (N_12706,N_11823,N_11495);
or U12707 (N_12707,N_11669,N_11778);
nor U12708 (N_12708,N_11500,N_11814);
xnor U12709 (N_12709,N_11603,N_11327);
nor U12710 (N_12710,N_11660,N_11819);
nand U12711 (N_12711,N_11668,N_11342);
and U12712 (N_12712,N_11294,N_11633);
nor U12713 (N_12713,N_11462,N_11907);
xnor U12714 (N_12714,N_11621,N_11872);
nand U12715 (N_12715,N_11468,N_11630);
nor U12716 (N_12716,N_11828,N_11655);
or U12717 (N_12717,N_11710,N_11473);
nor U12718 (N_12718,N_11994,N_11648);
nor U12719 (N_12719,N_11512,N_11522);
nor U12720 (N_12720,N_11457,N_11623);
or U12721 (N_12721,N_11812,N_11989);
and U12722 (N_12722,N_11567,N_11954);
or U12723 (N_12723,N_11309,N_11905);
nor U12724 (N_12724,N_11604,N_11913);
nor U12725 (N_12725,N_11545,N_11678);
or U12726 (N_12726,N_11262,N_11474);
and U12727 (N_12727,N_11363,N_11300);
nand U12728 (N_12728,N_11693,N_11452);
nor U12729 (N_12729,N_11744,N_11388);
and U12730 (N_12730,N_11575,N_11343);
xor U12731 (N_12731,N_11980,N_11303);
or U12732 (N_12732,N_11951,N_11655);
xnor U12733 (N_12733,N_11940,N_11743);
nor U12734 (N_12734,N_11938,N_11866);
and U12735 (N_12735,N_11606,N_11497);
nand U12736 (N_12736,N_11451,N_11325);
or U12737 (N_12737,N_11820,N_11588);
nand U12738 (N_12738,N_11722,N_11919);
and U12739 (N_12739,N_11815,N_11421);
and U12740 (N_12740,N_11253,N_11426);
or U12741 (N_12741,N_11919,N_11962);
nand U12742 (N_12742,N_11621,N_11334);
or U12743 (N_12743,N_11383,N_11677);
and U12744 (N_12744,N_11579,N_11274);
nand U12745 (N_12745,N_11533,N_11474);
and U12746 (N_12746,N_11811,N_11635);
xor U12747 (N_12747,N_11588,N_11389);
nand U12748 (N_12748,N_11796,N_11860);
nor U12749 (N_12749,N_11956,N_11640);
and U12750 (N_12750,N_12587,N_12714);
or U12751 (N_12751,N_12327,N_12466);
or U12752 (N_12752,N_12566,N_12238);
and U12753 (N_12753,N_12163,N_12440);
or U12754 (N_12754,N_12319,N_12116);
nand U12755 (N_12755,N_12222,N_12356);
and U12756 (N_12756,N_12366,N_12124);
and U12757 (N_12757,N_12737,N_12670);
nand U12758 (N_12758,N_12530,N_12479);
or U12759 (N_12759,N_12224,N_12552);
or U12760 (N_12760,N_12653,N_12660);
and U12761 (N_12761,N_12394,N_12209);
nor U12762 (N_12762,N_12656,N_12353);
nand U12763 (N_12763,N_12623,N_12457);
nand U12764 (N_12764,N_12627,N_12279);
nand U12765 (N_12765,N_12599,N_12326);
nor U12766 (N_12766,N_12151,N_12459);
nor U12767 (N_12767,N_12174,N_12452);
nor U12768 (N_12768,N_12518,N_12484);
or U12769 (N_12769,N_12684,N_12683);
or U12770 (N_12770,N_12519,N_12536);
and U12771 (N_12771,N_12483,N_12244);
nand U12772 (N_12772,N_12748,N_12503);
and U12773 (N_12773,N_12490,N_12139);
or U12774 (N_12774,N_12525,N_12091);
and U12775 (N_12775,N_12314,N_12245);
xor U12776 (N_12776,N_12060,N_12411);
or U12777 (N_12777,N_12720,N_12210);
nor U12778 (N_12778,N_12137,N_12056);
nor U12779 (N_12779,N_12239,N_12157);
and U12780 (N_12780,N_12223,N_12702);
nand U12781 (N_12781,N_12333,N_12383);
xnor U12782 (N_12782,N_12213,N_12711);
nor U12783 (N_12783,N_12251,N_12300);
nand U12784 (N_12784,N_12712,N_12078);
or U12785 (N_12785,N_12260,N_12634);
nand U12786 (N_12786,N_12571,N_12414);
xor U12787 (N_12787,N_12351,N_12334);
nand U12788 (N_12788,N_12572,N_12087);
and U12789 (N_12789,N_12665,N_12299);
and U12790 (N_12790,N_12134,N_12008);
nand U12791 (N_12791,N_12183,N_12232);
or U12792 (N_12792,N_12680,N_12123);
nor U12793 (N_12793,N_12724,N_12674);
or U12794 (N_12794,N_12731,N_12713);
nand U12795 (N_12795,N_12565,N_12497);
nor U12796 (N_12796,N_12036,N_12092);
and U12797 (N_12797,N_12603,N_12598);
nor U12798 (N_12798,N_12585,N_12025);
nor U12799 (N_12799,N_12359,N_12147);
and U12800 (N_12800,N_12551,N_12102);
or U12801 (N_12801,N_12371,N_12622);
or U12802 (N_12802,N_12425,N_12258);
nand U12803 (N_12803,N_12318,N_12156);
xor U12804 (N_12804,N_12246,N_12203);
and U12805 (N_12805,N_12038,N_12654);
nand U12806 (N_12806,N_12591,N_12482);
xnor U12807 (N_12807,N_12478,N_12372);
and U12808 (N_12808,N_12013,N_12403);
nand U12809 (N_12809,N_12419,N_12377);
nand U12810 (N_12810,N_12690,N_12494);
or U12811 (N_12811,N_12271,N_12256);
xnor U12812 (N_12812,N_12114,N_12584);
or U12813 (N_12813,N_12563,N_12301);
nand U12814 (N_12814,N_12336,N_12589);
nand U12815 (N_12815,N_12172,N_12605);
or U12816 (N_12816,N_12586,N_12241);
nand U12817 (N_12817,N_12168,N_12272);
nand U12818 (N_12818,N_12216,N_12645);
or U12819 (N_12819,N_12000,N_12606);
nand U12820 (N_12820,N_12662,N_12669);
nand U12821 (N_12821,N_12625,N_12220);
xnor U12822 (N_12822,N_12167,N_12495);
nor U12823 (N_12823,N_12588,N_12335);
and U12824 (N_12824,N_12264,N_12707);
xnor U12825 (N_12825,N_12728,N_12595);
nand U12826 (N_12826,N_12066,N_12171);
and U12827 (N_12827,N_12744,N_12706);
or U12828 (N_12828,N_12109,N_12590);
xor U12829 (N_12829,N_12568,N_12447);
or U12830 (N_12830,N_12397,N_12095);
xor U12831 (N_12831,N_12541,N_12212);
nand U12832 (N_12832,N_12685,N_12570);
nor U12833 (N_12833,N_12199,N_12019);
and U12834 (N_12834,N_12026,N_12321);
and U12835 (N_12835,N_12057,N_12323);
or U12836 (N_12836,N_12053,N_12655);
nor U12837 (N_12837,N_12320,N_12369);
and U12838 (N_12838,N_12010,N_12396);
or U12839 (N_12839,N_12030,N_12405);
nand U12840 (N_12840,N_12636,N_12436);
nand U12841 (N_12841,N_12122,N_12449);
xor U12842 (N_12842,N_12144,N_12557);
nand U12843 (N_12843,N_12108,N_12170);
nand U12844 (N_12844,N_12154,N_12069);
or U12845 (N_12845,N_12128,N_12149);
nor U12846 (N_12846,N_12024,N_12666);
xnor U12847 (N_12847,N_12675,N_12637);
xnor U12848 (N_12848,N_12499,N_12138);
nand U12849 (N_12849,N_12727,N_12671);
nor U12850 (N_12850,N_12578,N_12677);
nand U12851 (N_12851,N_12464,N_12288);
nor U12852 (N_12852,N_12221,N_12158);
or U12853 (N_12853,N_12225,N_12045);
or U12854 (N_12854,N_12522,N_12415);
and U12855 (N_12855,N_12746,N_12364);
or U12856 (N_12856,N_12088,N_12237);
and U12857 (N_12857,N_12190,N_12658);
xnor U12858 (N_12858,N_12663,N_12041);
and U12859 (N_12859,N_12249,N_12145);
and U12860 (N_12860,N_12455,N_12701);
nor U12861 (N_12861,N_12480,N_12446);
and U12862 (N_12862,N_12474,N_12579);
nand U12863 (N_12863,N_12597,N_12614);
or U12864 (N_12864,N_12621,N_12352);
nand U12865 (N_12865,N_12341,N_12194);
and U12866 (N_12866,N_12534,N_12016);
nand U12867 (N_12867,N_12079,N_12136);
nand U12868 (N_12868,N_12009,N_12097);
or U12869 (N_12869,N_12063,N_12186);
and U12870 (N_12870,N_12179,N_12560);
xnor U12871 (N_12871,N_12491,N_12506);
nor U12872 (N_12872,N_12442,N_12242);
and U12873 (N_12873,N_12098,N_12559);
xor U12874 (N_12874,N_12704,N_12460);
or U12875 (N_12875,N_12650,N_12725);
nand U12876 (N_12876,N_12287,N_12094);
nand U12877 (N_12877,N_12281,N_12197);
nor U12878 (N_12878,N_12517,N_12234);
or U12879 (N_12879,N_12076,N_12006);
or U12880 (N_12880,N_12740,N_12062);
nand U12881 (N_12881,N_12023,N_12120);
nor U12882 (N_12882,N_12472,N_12280);
nand U12883 (N_12883,N_12526,N_12343);
or U12884 (N_12884,N_12747,N_12125);
xnor U12885 (N_12885,N_12404,N_12421);
nor U12886 (N_12886,N_12127,N_12523);
nor U12887 (N_12887,N_12718,N_12428);
xor U12888 (N_12888,N_12236,N_12620);
or U12889 (N_12889,N_12601,N_12409);
or U12890 (N_12890,N_12015,N_12514);
nand U12891 (N_12891,N_12513,N_12035);
or U12892 (N_12892,N_12561,N_12741);
nor U12893 (N_12893,N_12148,N_12354);
or U12894 (N_12894,N_12569,N_12667);
or U12895 (N_12895,N_12705,N_12412);
or U12896 (N_12896,N_12500,N_12002);
and U12897 (N_12897,N_12227,N_12233);
or U12898 (N_12898,N_12073,N_12119);
xnor U12899 (N_12899,N_12535,N_12337);
nor U12900 (N_12900,N_12043,N_12161);
or U12901 (N_12901,N_12304,N_12577);
xnor U12902 (N_12902,N_12202,N_12681);
or U12903 (N_12903,N_12730,N_12450);
and U12904 (N_12904,N_12608,N_12435);
nor U12905 (N_12905,N_12059,N_12611);
xnor U12906 (N_12906,N_12735,N_12485);
or U12907 (N_12907,N_12538,N_12292);
and U12908 (N_12908,N_12722,N_12291);
or U12909 (N_12909,N_12528,N_12182);
nor U12910 (N_12910,N_12070,N_12185);
and U12911 (N_12911,N_12481,N_12039);
xnor U12912 (N_12912,N_12709,N_12020);
or U12913 (N_12913,N_12574,N_12261);
nand U12914 (N_12914,N_12742,N_12150);
and U12915 (N_12915,N_12520,N_12391);
nor U12916 (N_12916,N_12378,N_12324);
nor U12917 (N_12917,N_12434,N_12592);
xor U12918 (N_12918,N_12061,N_12708);
and U12919 (N_12919,N_12255,N_12355);
nor U12920 (N_12920,N_12229,N_12505);
xnor U12921 (N_12921,N_12562,N_12527);
nor U12922 (N_12922,N_12386,N_12099);
xnor U12923 (N_12923,N_12005,N_12338);
or U12924 (N_12924,N_12311,N_12177);
nor U12925 (N_12925,N_12198,N_12159);
or U12926 (N_12926,N_12376,N_12107);
xor U12927 (N_12927,N_12529,N_12676);
nand U12928 (N_12928,N_12721,N_12286);
and U12929 (N_12929,N_12382,N_12370);
and U12930 (N_12930,N_12090,N_12470);
or U12931 (N_12931,N_12027,N_12454);
or U12932 (N_12932,N_12248,N_12498);
and U12933 (N_12933,N_12263,N_12465);
or U12934 (N_12934,N_12646,N_12384);
and U12935 (N_12935,N_12423,N_12379);
nand U12936 (N_12936,N_12389,N_12651);
or U12937 (N_12937,N_12630,N_12668);
nor U12938 (N_12938,N_12130,N_12739);
nand U12939 (N_12939,N_12080,N_12710);
nor U12940 (N_12940,N_12349,N_12439);
nand U12941 (N_12941,N_12407,N_12451);
nor U12942 (N_12942,N_12253,N_12101);
or U12943 (N_12943,N_12188,N_12029);
nand U12944 (N_12944,N_12432,N_12184);
nor U12945 (N_12945,N_12247,N_12420);
and U12946 (N_12946,N_12678,N_12325);
nor U12947 (N_12947,N_12112,N_12211);
or U12948 (N_12948,N_12697,N_12100);
and U12949 (N_12949,N_12118,N_12294);
xor U12950 (N_12950,N_12406,N_12192);
and U12951 (N_12951,N_12339,N_12594);
or U12952 (N_12952,N_12141,N_12208);
or U12953 (N_12953,N_12516,N_12607);
nor U12954 (N_12954,N_12072,N_12135);
nor U12955 (N_12955,N_12049,N_12315);
and U12956 (N_12956,N_12165,N_12558);
or U12957 (N_12957,N_12306,N_12152);
nor U12958 (N_12958,N_12084,N_12374);
xnor U12959 (N_12959,N_12347,N_12723);
and U12960 (N_12960,N_12430,N_12042);
and U12961 (N_12961,N_12082,N_12071);
xnor U12962 (N_12962,N_12302,N_12508);
xor U12963 (N_12963,N_12537,N_12745);
nor U12964 (N_12964,N_12433,N_12738);
or U12965 (N_12965,N_12290,N_12254);
nor U12966 (N_12966,N_12546,N_12007);
nor U12967 (N_12967,N_12583,N_12240);
and U12968 (N_12968,N_12047,N_12226);
nor U12969 (N_12969,N_12657,N_12331);
nand U12970 (N_12970,N_12257,N_12031);
nand U12971 (N_12971,N_12673,N_12596);
nand U12972 (N_12972,N_12295,N_12664);
and U12973 (N_12973,N_12357,N_12052);
xor U12974 (N_12974,N_12126,N_12160);
xor U12975 (N_12975,N_12231,N_12618);
or U12976 (N_12976,N_12215,N_12417);
or U12977 (N_12977,N_12316,N_12093);
nor U12978 (N_12978,N_12330,N_12462);
and U12979 (N_12979,N_12077,N_12313);
nand U12980 (N_12980,N_12283,N_12162);
nor U12981 (N_12981,N_12032,N_12547);
nor U12982 (N_12982,N_12489,N_12749);
and U12983 (N_12983,N_12582,N_12539);
and U12984 (N_12984,N_12613,N_12661);
nand U12985 (N_12985,N_12471,N_12543);
and U12986 (N_12986,N_12553,N_12413);
and U12987 (N_12987,N_12317,N_12243);
nor U12988 (N_12988,N_12687,N_12729);
and U12989 (N_12989,N_12629,N_12328);
and U12990 (N_12990,N_12204,N_12081);
or U12991 (N_12991,N_12219,N_12422);
nor U12992 (N_12992,N_12269,N_12133);
or U12993 (N_12993,N_12488,N_12003);
nand U12994 (N_12994,N_12703,N_12140);
nor U12995 (N_12995,N_12549,N_12395);
nor U12996 (N_12996,N_12619,N_12350);
and U12997 (N_12997,N_12217,N_12228);
nor U12998 (N_12998,N_12265,N_12401);
nand U12999 (N_12999,N_12187,N_12166);
nand U13000 (N_13000,N_12146,N_12554);
xnor U13001 (N_13001,N_12715,N_12461);
nand U13002 (N_13002,N_12524,N_12293);
xnor U13003 (N_13003,N_12278,N_12688);
and U13004 (N_13004,N_12437,N_12429);
nand U13005 (N_13005,N_12410,N_12682);
nand U13006 (N_13006,N_12544,N_12473);
nor U13007 (N_13007,N_12115,N_12103);
or U13008 (N_13008,N_12282,N_12632);
nand U13009 (N_13009,N_12033,N_12626);
and U13010 (N_13010,N_12085,N_12453);
xnor U13011 (N_13011,N_12493,N_12507);
or U13012 (N_13012,N_12178,N_12196);
nand U13013 (N_13013,N_12445,N_12262);
nand U13014 (N_13014,N_12131,N_12733);
or U13015 (N_13015,N_12207,N_12610);
nor U13016 (N_13016,N_12067,N_12113);
nor U13017 (N_13017,N_12298,N_12700);
nor U13018 (N_13018,N_12380,N_12443);
or U13019 (N_13019,N_12096,N_12694);
and U13020 (N_13020,N_12051,N_12487);
nand U13021 (N_13021,N_12046,N_12652);
nor U13022 (N_13022,N_12548,N_12180);
or U13023 (N_13023,N_12512,N_12693);
nor U13024 (N_13024,N_12468,N_12270);
xor U13025 (N_13025,N_12106,N_12322);
or U13026 (N_13026,N_12312,N_12521);
or U13027 (N_13027,N_12573,N_12201);
or U13028 (N_13028,N_12424,N_12361);
or U13029 (N_13029,N_12696,N_12624);
or U13030 (N_13030,N_12344,N_12089);
nand U13031 (N_13031,N_12310,N_12075);
and U13032 (N_13032,N_12475,N_12285);
and U13033 (N_13033,N_12486,N_12307);
nand U13034 (N_13034,N_12346,N_12054);
nand U13035 (N_13035,N_12289,N_12385);
or U13036 (N_13036,N_12679,N_12532);
nor U13037 (N_13037,N_12416,N_12510);
or U13038 (N_13038,N_12719,N_12164);
or U13039 (N_13039,N_12575,N_12533);
and U13040 (N_13040,N_12218,N_12064);
xor U13041 (N_13041,N_12362,N_12305);
and U13042 (N_13042,N_12155,N_12550);
nand U13043 (N_13043,N_12639,N_12068);
nand U13044 (N_13044,N_12441,N_12252);
nand U13045 (N_13045,N_12476,N_12360);
nor U13046 (N_13046,N_12050,N_12205);
and U13047 (N_13047,N_12644,N_12176);
xor U13048 (N_13048,N_12332,N_12504);
and U13049 (N_13049,N_12345,N_12086);
and U13050 (N_13050,N_12542,N_12153);
nor U13051 (N_13051,N_12399,N_12531);
nor U13052 (N_13052,N_12277,N_12580);
and U13053 (N_13053,N_12250,N_12274);
nor U13054 (N_13054,N_12408,N_12612);
nand U13055 (N_13055,N_12275,N_12104);
and U13056 (N_13056,N_12048,N_12117);
or U13057 (N_13057,N_12686,N_12129);
and U13058 (N_13058,N_12477,N_12398);
and U13059 (N_13059,N_12193,N_12309);
nand U13060 (N_13060,N_12173,N_12649);
nor U13061 (N_13061,N_12392,N_12132);
nor U13062 (N_13062,N_12022,N_12111);
xnor U13063 (N_13063,N_12438,N_12736);
nor U13064 (N_13064,N_12593,N_12635);
or U13065 (N_13065,N_12235,N_12267);
nand U13066 (N_13066,N_12017,N_12540);
nand U13067 (N_13067,N_12175,N_12659);
nor U13068 (N_13068,N_12492,N_12444);
nand U13069 (N_13069,N_12648,N_12600);
and U13070 (N_13070,N_12367,N_12609);
or U13071 (N_13071,N_12284,N_12555);
or U13072 (N_13072,N_12647,N_12373);
and U13073 (N_13073,N_12058,N_12400);
nand U13074 (N_13074,N_12469,N_12368);
nor U13075 (N_13075,N_12640,N_12689);
nor U13076 (N_13076,N_12456,N_12342);
nand U13077 (N_13077,N_12083,N_12699);
nor U13078 (N_13078,N_12259,N_12191);
nor U13079 (N_13079,N_12509,N_12044);
nand U13080 (N_13080,N_12268,N_12230);
nand U13081 (N_13081,N_12340,N_12638);
or U13082 (N_13082,N_12616,N_12458);
and U13083 (N_13083,N_12717,N_12308);
nand U13084 (N_13084,N_12695,N_12581);
nor U13085 (N_13085,N_12200,N_12716);
or U13086 (N_13086,N_12556,N_12515);
or U13087 (N_13087,N_12037,N_12381);
nor U13088 (N_13088,N_12427,N_12358);
nor U13089 (N_13089,N_12375,N_12142);
nand U13090 (N_13090,N_12034,N_12567);
or U13091 (N_13091,N_12273,N_12463);
nor U13092 (N_13092,N_12169,N_12021);
nand U13093 (N_13093,N_12363,N_12643);
nor U13094 (N_13094,N_12431,N_12743);
and U13095 (N_13095,N_12502,N_12388);
xor U13096 (N_13096,N_12181,N_12576);
or U13097 (N_13097,N_12206,N_12266);
nand U13098 (N_13098,N_12018,N_12012);
or U13099 (N_13099,N_12672,N_12001);
or U13100 (N_13100,N_12496,N_12303);
nand U13101 (N_13101,N_12467,N_12393);
nor U13102 (N_13102,N_12604,N_12692);
and U13103 (N_13103,N_12011,N_12426);
xor U13104 (N_13104,N_12040,N_12004);
or U13105 (N_13105,N_12602,N_12276);
or U13106 (N_13106,N_12387,N_12121);
and U13107 (N_13107,N_12296,N_12564);
and U13108 (N_13108,N_12014,N_12631);
and U13109 (N_13109,N_12055,N_12329);
nand U13110 (N_13110,N_12065,N_12189);
and U13111 (N_13111,N_12214,N_12726);
nand U13112 (N_13112,N_12511,N_12105);
nand U13113 (N_13113,N_12732,N_12418);
or U13114 (N_13114,N_12641,N_12074);
nand U13115 (N_13115,N_12734,N_12617);
or U13116 (N_13116,N_12348,N_12028);
or U13117 (N_13117,N_12143,N_12615);
and U13118 (N_13118,N_12698,N_12545);
nor U13119 (N_13119,N_12365,N_12195);
xnor U13120 (N_13120,N_12633,N_12501);
nand U13121 (N_13121,N_12390,N_12110);
xnor U13122 (N_13122,N_12628,N_12642);
nand U13123 (N_13123,N_12402,N_12448);
or U13124 (N_13124,N_12691,N_12297);
nand U13125 (N_13125,N_12308,N_12239);
nand U13126 (N_13126,N_12009,N_12246);
and U13127 (N_13127,N_12574,N_12184);
and U13128 (N_13128,N_12103,N_12124);
nor U13129 (N_13129,N_12296,N_12089);
nand U13130 (N_13130,N_12437,N_12346);
and U13131 (N_13131,N_12232,N_12184);
nor U13132 (N_13132,N_12586,N_12453);
xor U13133 (N_13133,N_12264,N_12686);
nor U13134 (N_13134,N_12129,N_12228);
xor U13135 (N_13135,N_12432,N_12433);
and U13136 (N_13136,N_12417,N_12735);
nand U13137 (N_13137,N_12194,N_12084);
nor U13138 (N_13138,N_12638,N_12151);
nor U13139 (N_13139,N_12231,N_12196);
nand U13140 (N_13140,N_12409,N_12374);
nor U13141 (N_13141,N_12596,N_12112);
or U13142 (N_13142,N_12119,N_12222);
nand U13143 (N_13143,N_12068,N_12486);
and U13144 (N_13144,N_12496,N_12232);
nand U13145 (N_13145,N_12199,N_12028);
nand U13146 (N_13146,N_12609,N_12282);
xnor U13147 (N_13147,N_12201,N_12435);
or U13148 (N_13148,N_12422,N_12443);
and U13149 (N_13149,N_12614,N_12080);
and U13150 (N_13150,N_12692,N_12662);
and U13151 (N_13151,N_12595,N_12148);
or U13152 (N_13152,N_12613,N_12308);
or U13153 (N_13153,N_12339,N_12560);
and U13154 (N_13154,N_12597,N_12225);
xor U13155 (N_13155,N_12367,N_12480);
and U13156 (N_13156,N_12597,N_12664);
or U13157 (N_13157,N_12692,N_12441);
nand U13158 (N_13158,N_12289,N_12042);
or U13159 (N_13159,N_12239,N_12368);
and U13160 (N_13160,N_12580,N_12392);
xor U13161 (N_13161,N_12590,N_12432);
or U13162 (N_13162,N_12657,N_12592);
and U13163 (N_13163,N_12081,N_12386);
or U13164 (N_13164,N_12179,N_12427);
nand U13165 (N_13165,N_12700,N_12576);
nand U13166 (N_13166,N_12214,N_12577);
nand U13167 (N_13167,N_12662,N_12418);
nand U13168 (N_13168,N_12687,N_12727);
or U13169 (N_13169,N_12725,N_12368);
nand U13170 (N_13170,N_12198,N_12720);
or U13171 (N_13171,N_12010,N_12255);
nor U13172 (N_13172,N_12437,N_12533);
nor U13173 (N_13173,N_12632,N_12208);
or U13174 (N_13174,N_12418,N_12293);
nor U13175 (N_13175,N_12367,N_12287);
nand U13176 (N_13176,N_12559,N_12042);
and U13177 (N_13177,N_12674,N_12270);
or U13178 (N_13178,N_12696,N_12013);
nand U13179 (N_13179,N_12733,N_12663);
and U13180 (N_13180,N_12596,N_12453);
nand U13181 (N_13181,N_12446,N_12721);
or U13182 (N_13182,N_12314,N_12391);
xnor U13183 (N_13183,N_12288,N_12217);
nor U13184 (N_13184,N_12264,N_12311);
nor U13185 (N_13185,N_12258,N_12131);
nand U13186 (N_13186,N_12039,N_12290);
or U13187 (N_13187,N_12400,N_12674);
nand U13188 (N_13188,N_12569,N_12711);
xnor U13189 (N_13189,N_12161,N_12587);
nand U13190 (N_13190,N_12157,N_12275);
or U13191 (N_13191,N_12627,N_12053);
nand U13192 (N_13192,N_12125,N_12261);
xor U13193 (N_13193,N_12636,N_12707);
or U13194 (N_13194,N_12432,N_12021);
or U13195 (N_13195,N_12110,N_12346);
or U13196 (N_13196,N_12489,N_12168);
nor U13197 (N_13197,N_12647,N_12576);
nand U13198 (N_13198,N_12566,N_12699);
nor U13199 (N_13199,N_12499,N_12006);
and U13200 (N_13200,N_12231,N_12659);
nor U13201 (N_13201,N_12413,N_12665);
nand U13202 (N_13202,N_12290,N_12032);
and U13203 (N_13203,N_12674,N_12378);
nand U13204 (N_13204,N_12216,N_12072);
nand U13205 (N_13205,N_12212,N_12409);
or U13206 (N_13206,N_12102,N_12245);
and U13207 (N_13207,N_12539,N_12588);
or U13208 (N_13208,N_12654,N_12473);
nand U13209 (N_13209,N_12479,N_12585);
nor U13210 (N_13210,N_12376,N_12058);
and U13211 (N_13211,N_12250,N_12476);
nand U13212 (N_13212,N_12595,N_12090);
nor U13213 (N_13213,N_12701,N_12525);
and U13214 (N_13214,N_12038,N_12714);
and U13215 (N_13215,N_12642,N_12676);
nor U13216 (N_13216,N_12573,N_12265);
nand U13217 (N_13217,N_12629,N_12457);
and U13218 (N_13218,N_12655,N_12500);
and U13219 (N_13219,N_12273,N_12326);
nand U13220 (N_13220,N_12236,N_12041);
nand U13221 (N_13221,N_12036,N_12023);
or U13222 (N_13222,N_12349,N_12069);
nor U13223 (N_13223,N_12434,N_12189);
and U13224 (N_13224,N_12551,N_12123);
nand U13225 (N_13225,N_12441,N_12342);
and U13226 (N_13226,N_12215,N_12299);
or U13227 (N_13227,N_12306,N_12292);
or U13228 (N_13228,N_12576,N_12649);
nor U13229 (N_13229,N_12657,N_12198);
or U13230 (N_13230,N_12153,N_12535);
and U13231 (N_13231,N_12540,N_12525);
nand U13232 (N_13232,N_12038,N_12022);
and U13233 (N_13233,N_12144,N_12503);
nand U13234 (N_13234,N_12627,N_12402);
nor U13235 (N_13235,N_12317,N_12462);
xor U13236 (N_13236,N_12456,N_12336);
nand U13237 (N_13237,N_12402,N_12366);
nor U13238 (N_13238,N_12295,N_12251);
xor U13239 (N_13239,N_12703,N_12272);
nor U13240 (N_13240,N_12534,N_12114);
or U13241 (N_13241,N_12158,N_12123);
and U13242 (N_13242,N_12315,N_12473);
xnor U13243 (N_13243,N_12152,N_12370);
nand U13244 (N_13244,N_12543,N_12740);
nor U13245 (N_13245,N_12098,N_12568);
xnor U13246 (N_13246,N_12376,N_12348);
nor U13247 (N_13247,N_12639,N_12360);
and U13248 (N_13248,N_12263,N_12331);
or U13249 (N_13249,N_12646,N_12674);
nand U13250 (N_13250,N_12732,N_12099);
nand U13251 (N_13251,N_12511,N_12713);
nor U13252 (N_13252,N_12429,N_12052);
and U13253 (N_13253,N_12400,N_12708);
and U13254 (N_13254,N_12147,N_12492);
xnor U13255 (N_13255,N_12552,N_12080);
or U13256 (N_13256,N_12314,N_12550);
and U13257 (N_13257,N_12240,N_12727);
nor U13258 (N_13258,N_12146,N_12307);
and U13259 (N_13259,N_12310,N_12430);
nor U13260 (N_13260,N_12057,N_12544);
nand U13261 (N_13261,N_12035,N_12461);
xor U13262 (N_13262,N_12531,N_12509);
and U13263 (N_13263,N_12420,N_12441);
nand U13264 (N_13264,N_12024,N_12478);
and U13265 (N_13265,N_12547,N_12700);
or U13266 (N_13266,N_12674,N_12283);
nand U13267 (N_13267,N_12749,N_12676);
or U13268 (N_13268,N_12294,N_12221);
nand U13269 (N_13269,N_12014,N_12006);
nand U13270 (N_13270,N_12548,N_12670);
and U13271 (N_13271,N_12217,N_12165);
or U13272 (N_13272,N_12722,N_12155);
and U13273 (N_13273,N_12475,N_12268);
nor U13274 (N_13274,N_12431,N_12560);
and U13275 (N_13275,N_12703,N_12599);
nor U13276 (N_13276,N_12398,N_12662);
and U13277 (N_13277,N_12540,N_12375);
or U13278 (N_13278,N_12319,N_12422);
nor U13279 (N_13279,N_12566,N_12350);
xnor U13280 (N_13280,N_12710,N_12564);
nor U13281 (N_13281,N_12418,N_12171);
or U13282 (N_13282,N_12724,N_12721);
nor U13283 (N_13283,N_12357,N_12615);
xnor U13284 (N_13284,N_12738,N_12188);
or U13285 (N_13285,N_12461,N_12051);
and U13286 (N_13286,N_12607,N_12206);
and U13287 (N_13287,N_12654,N_12017);
or U13288 (N_13288,N_12633,N_12306);
or U13289 (N_13289,N_12263,N_12558);
nor U13290 (N_13290,N_12160,N_12239);
and U13291 (N_13291,N_12241,N_12242);
and U13292 (N_13292,N_12465,N_12445);
nor U13293 (N_13293,N_12502,N_12198);
and U13294 (N_13294,N_12304,N_12449);
or U13295 (N_13295,N_12296,N_12325);
xnor U13296 (N_13296,N_12517,N_12432);
or U13297 (N_13297,N_12463,N_12354);
nand U13298 (N_13298,N_12745,N_12027);
and U13299 (N_13299,N_12031,N_12314);
nand U13300 (N_13300,N_12527,N_12490);
nor U13301 (N_13301,N_12444,N_12647);
or U13302 (N_13302,N_12431,N_12154);
or U13303 (N_13303,N_12257,N_12161);
and U13304 (N_13304,N_12421,N_12407);
or U13305 (N_13305,N_12666,N_12042);
nor U13306 (N_13306,N_12564,N_12423);
nor U13307 (N_13307,N_12042,N_12359);
and U13308 (N_13308,N_12599,N_12261);
xor U13309 (N_13309,N_12406,N_12320);
nand U13310 (N_13310,N_12471,N_12385);
nor U13311 (N_13311,N_12175,N_12412);
nand U13312 (N_13312,N_12015,N_12719);
nand U13313 (N_13313,N_12131,N_12341);
and U13314 (N_13314,N_12608,N_12360);
nor U13315 (N_13315,N_12501,N_12429);
or U13316 (N_13316,N_12519,N_12206);
nand U13317 (N_13317,N_12701,N_12351);
nand U13318 (N_13318,N_12719,N_12563);
and U13319 (N_13319,N_12709,N_12163);
or U13320 (N_13320,N_12584,N_12558);
or U13321 (N_13321,N_12505,N_12333);
nor U13322 (N_13322,N_12298,N_12211);
nor U13323 (N_13323,N_12671,N_12036);
nand U13324 (N_13324,N_12084,N_12686);
xor U13325 (N_13325,N_12593,N_12265);
nor U13326 (N_13326,N_12676,N_12275);
nand U13327 (N_13327,N_12329,N_12292);
nand U13328 (N_13328,N_12441,N_12483);
and U13329 (N_13329,N_12526,N_12474);
nand U13330 (N_13330,N_12016,N_12699);
and U13331 (N_13331,N_12284,N_12725);
nor U13332 (N_13332,N_12244,N_12065);
nand U13333 (N_13333,N_12402,N_12729);
nor U13334 (N_13334,N_12058,N_12601);
or U13335 (N_13335,N_12322,N_12123);
or U13336 (N_13336,N_12227,N_12335);
nor U13337 (N_13337,N_12284,N_12174);
nand U13338 (N_13338,N_12649,N_12157);
nor U13339 (N_13339,N_12249,N_12034);
nand U13340 (N_13340,N_12616,N_12581);
nand U13341 (N_13341,N_12347,N_12521);
nand U13342 (N_13342,N_12633,N_12015);
nor U13343 (N_13343,N_12489,N_12312);
nor U13344 (N_13344,N_12328,N_12480);
or U13345 (N_13345,N_12042,N_12637);
nand U13346 (N_13346,N_12351,N_12089);
xor U13347 (N_13347,N_12696,N_12444);
nand U13348 (N_13348,N_12427,N_12233);
and U13349 (N_13349,N_12736,N_12348);
and U13350 (N_13350,N_12747,N_12036);
or U13351 (N_13351,N_12063,N_12159);
and U13352 (N_13352,N_12282,N_12430);
xnor U13353 (N_13353,N_12487,N_12433);
nand U13354 (N_13354,N_12308,N_12498);
nand U13355 (N_13355,N_12309,N_12297);
nand U13356 (N_13356,N_12267,N_12312);
xor U13357 (N_13357,N_12701,N_12121);
nor U13358 (N_13358,N_12013,N_12441);
nand U13359 (N_13359,N_12211,N_12153);
or U13360 (N_13360,N_12375,N_12287);
and U13361 (N_13361,N_12677,N_12313);
nor U13362 (N_13362,N_12028,N_12549);
and U13363 (N_13363,N_12650,N_12682);
xnor U13364 (N_13364,N_12336,N_12211);
and U13365 (N_13365,N_12651,N_12445);
or U13366 (N_13366,N_12688,N_12652);
or U13367 (N_13367,N_12437,N_12729);
nor U13368 (N_13368,N_12512,N_12459);
or U13369 (N_13369,N_12185,N_12080);
and U13370 (N_13370,N_12611,N_12641);
and U13371 (N_13371,N_12062,N_12173);
nand U13372 (N_13372,N_12474,N_12570);
or U13373 (N_13373,N_12577,N_12372);
xor U13374 (N_13374,N_12728,N_12329);
nand U13375 (N_13375,N_12011,N_12253);
or U13376 (N_13376,N_12634,N_12628);
nor U13377 (N_13377,N_12261,N_12329);
and U13378 (N_13378,N_12046,N_12170);
nand U13379 (N_13379,N_12320,N_12404);
or U13380 (N_13380,N_12339,N_12526);
nor U13381 (N_13381,N_12672,N_12217);
xnor U13382 (N_13382,N_12516,N_12432);
xnor U13383 (N_13383,N_12725,N_12058);
nand U13384 (N_13384,N_12413,N_12039);
nor U13385 (N_13385,N_12721,N_12685);
or U13386 (N_13386,N_12686,N_12350);
nor U13387 (N_13387,N_12040,N_12690);
nor U13388 (N_13388,N_12129,N_12716);
nor U13389 (N_13389,N_12084,N_12141);
nand U13390 (N_13390,N_12362,N_12519);
or U13391 (N_13391,N_12591,N_12059);
xor U13392 (N_13392,N_12447,N_12368);
nor U13393 (N_13393,N_12569,N_12579);
nand U13394 (N_13394,N_12502,N_12037);
or U13395 (N_13395,N_12441,N_12215);
nand U13396 (N_13396,N_12407,N_12447);
nand U13397 (N_13397,N_12705,N_12028);
or U13398 (N_13398,N_12737,N_12711);
or U13399 (N_13399,N_12382,N_12297);
nand U13400 (N_13400,N_12268,N_12713);
nor U13401 (N_13401,N_12559,N_12166);
nand U13402 (N_13402,N_12338,N_12612);
nor U13403 (N_13403,N_12647,N_12408);
xor U13404 (N_13404,N_12417,N_12573);
nor U13405 (N_13405,N_12511,N_12252);
xnor U13406 (N_13406,N_12061,N_12054);
or U13407 (N_13407,N_12723,N_12338);
or U13408 (N_13408,N_12397,N_12272);
or U13409 (N_13409,N_12021,N_12303);
nand U13410 (N_13410,N_12133,N_12434);
nand U13411 (N_13411,N_12180,N_12160);
nand U13412 (N_13412,N_12535,N_12026);
nor U13413 (N_13413,N_12100,N_12062);
and U13414 (N_13414,N_12141,N_12673);
nor U13415 (N_13415,N_12394,N_12185);
xnor U13416 (N_13416,N_12121,N_12392);
nor U13417 (N_13417,N_12052,N_12720);
or U13418 (N_13418,N_12266,N_12484);
nor U13419 (N_13419,N_12699,N_12600);
or U13420 (N_13420,N_12139,N_12625);
or U13421 (N_13421,N_12602,N_12381);
or U13422 (N_13422,N_12092,N_12001);
nand U13423 (N_13423,N_12216,N_12327);
nand U13424 (N_13424,N_12377,N_12667);
nor U13425 (N_13425,N_12677,N_12471);
nand U13426 (N_13426,N_12067,N_12420);
nor U13427 (N_13427,N_12307,N_12708);
and U13428 (N_13428,N_12012,N_12220);
nand U13429 (N_13429,N_12193,N_12389);
nor U13430 (N_13430,N_12173,N_12373);
or U13431 (N_13431,N_12475,N_12021);
nand U13432 (N_13432,N_12246,N_12375);
xor U13433 (N_13433,N_12491,N_12129);
xor U13434 (N_13434,N_12629,N_12403);
xnor U13435 (N_13435,N_12605,N_12397);
xnor U13436 (N_13436,N_12097,N_12110);
and U13437 (N_13437,N_12371,N_12726);
or U13438 (N_13438,N_12438,N_12510);
or U13439 (N_13439,N_12579,N_12400);
nor U13440 (N_13440,N_12063,N_12274);
or U13441 (N_13441,N_12128,N_12404);
and U13442 (N_13442,N_12584,N_12646);
nand U13443 (N_13443,N_12000,N_12434);
or U13444 (N_13444,N_12413,N_12294);
or U13445 (N_13445,N_12217,N_12450);
or U13446 (N_13446,N_12096,N_12021);
or U13447 (N_13447,N_12176,N_12114);
xnor U13448 (N_13448,N_12472,N_12392);
nand U13449 (N_13449,N_12192,N_12667);
nand U13450 (N_13450,N_12493,N_12686);
nor U13451 (N_13451,N_12109,N_12089);
nor U13452 (N_13452,N_12131,N_12076);
nor U13453 (N_13453,N_12301,N_12149);
nor U13454 (N_13454,N_12218,N_12580);
nor U13455 (N_13455,N_12166,N_12067);
nor U13456 (N_13456,N_12362,N_12571);
nor U13457 (N_13457,N_12364,N_12594);
nor U13458 (N_13458,N_12645,N_12310);
or U13459 (N_13459,N_12706,N_12214);
and U13460 (N_13460,N_12275,N_12695);
nor U13461 (N_13461,N_12714,N_12397);
or U13462 (N_13462,N_12466,N_12393);
nor U13463 (N_13463,N_12405,N_12704);
and U13464 (N_13464,N_12141,N_12424);
nor U13465 (N_13465,N_12072,N_12276);
nor U13466 (N_13466,N_12189,N_12343);
and U13467 (N_13467,N_12461,N_12393);
and U13468 (N_13468,N_12362,N_12044);
and U13469 (N_13469,N_12362,N_12724);
xnor U13470 (N_13470,N_12088,N_12416);
and U13471 (N_13471,N_12259,N_12566);
nand U13472 (N_13472,N_12685,N_12553);
nor U13473 (N_13473,N_12013,N_12559);
nor U13474 (N_13474,N_12494,N_12179);
and U13475 (N_13475,N_12308,N_12282);
or U13476 (N_13476,N_12001,N_12117);
and U13477 (N_13477,N_12177,N_12314);
nor U13478 (N_13478,N_12355,N_12448);
or U13479 (N_13479,N_12523,N_12123);
or U13480 (N_13480,N_12027,N_12371);
and U13481 (N_13481,N_12254,N_12189);
nand U13482 (N_13482,N_12094,N_12715);
nand U13483 (N_13483,N_12548,N_12234);
or U13484 (N_13484,N_12664,N_12700);
or U13485 (N_13485,N_12277,N_12366);
or U13486 (N_13486,N_12134,N_12277);
xor U13487 (N_13487,N_12689,N_12376);
and U13488 (N_13488,N_12366,N_12313);
nor U13489 (N_13489,N_12112,N_12135);
or U13490 (N_13490,N_12570,N_12601);
or U13491 (N_13491,N_12477,N_12099);
nor U13492 (N_13492,N_12704,N_12069);
and U13493 (N_13493,N_12592,N_12391);
nand U13494 (N_13494,N_12416,N_12208);
nand U13495 (N_13495,N_12580,N_12296);
or U13496 (N_13496,N_12071,N_12582);
or U13497 (N_13497,N_12746,N_12395);
and U13498 (N_13498,N_12016,N_12437);
and U13499 (N_13499,N_12192,N_12516);
nand U13500 (N_13500,N_13113,N_13331);
and U13501 (N_13501,N_13013,N_12914);
nand U13502 (N_13502,N_13233,N_12807);
or U13503 (N_13503,N_13049,N_13403);
or U13504 (N_13504,N_12883,N_13121);
nand U13505 (N_13505,N_12798,N_12881);
nor U13506 (N_13506,N_13463,N_13185);
and U13507 (N_13507,N_13125,N_13365);
nand U13508 (N_13508,N_13028,N_12931);
and U13509 (N_13509,N_12844,N_13357);
nor U13510 (N_13510,N_13465,N_12759);
xor U13511 (N_13511,N_13257,N_13019);
xnor U13512 (N_13512,N_13399,N_13003);
nand U13513 (N_13513,N_12831,N_13175);
xor U13514 (N_13514,N_13434,N_13372);
or U13515 (N_13515,N_13116,N_12839);
nor U13516 (N_13516,N_13474,N_13203);
or U13517 (N_13517,N_12849,N_13353);
or U13518 (N_13518,N_13010,N_12940);
xnor U13519 (N_13519,N_13249,N_13222);
nand U13520 (N_13520,N_12991,N_13050);
and U13521 (N_13521,N_13297,N_12851);
or U13522 (N_13522,N_12752,N_13084);
nand U13523 (N_13523,N_12949,N_12868);
nand U13524 (N_13524,N_12987,N_13273);
nor U13525 (N_13525,N_13158,N_12898);
xor U13526 (N_13526,N_12767,N_12838);
nand U13527 (N_13527,N_12879,N_13215);
and U13528 (N_13528,N_13371,N_13124);
and U13529 (N_13529,N_12915,N_13339);
xor U13530 (N_13530,N_12869,N_13012);
or U13531 (N_13531,N_13380,N_13088);
xnor U13532 (N_13532,N_13060,N_13422);
nor U13533 (N_13533,N_12775,N_12800);
nand U13534 (N_13534,N_13398,N_13334);
nand U13535 (N_13535,N_13245,N_13412);
nor U13536 (N_13536,N_12997,N_12765);
and U13537 (N_13537,N_12818,N_12825);
or U13538 (N_13538,N_13486,N_12900);
nor U13539 (N_13539,N_13142,N_13234);
nand U13540 (N_13540,N_13497,N_12803);
nor U13541 (N_13541,N_13032,N_12768);
or U13542 (N_13542,N_12787,N_13256);
or U13543 (N_13543,N_13208,N_13082);
nand U13544 (N_13544,N_13355,N_12813);
nand U13545 (N_13545,N_13202,N_13494);
and U13546 (N_13546,N_12964,N_13106);
and U13547 (N_13547,N_12939,N_13345);
nand U13548 (N_13548,N_12791,N_13147);
nand U13549 (N_13549,N_13078,N_13254);
xnor U13550 (N_13550,N_13314,N_13296);
xnor U13551 (N_13551,N_13430,N_12756);
nand U13552 (N_13552,N_13002,N_13467);
and U13553 (N_13553,N_13413,N_13066);
and U13554 (N_13554,N_13235,N_13343);
nand U13555 (N_13555,N_12918,N_13476);
or U13556 (N_13556,N_12941,N_12856);
and U13557 (N_13557,N_13024,N_12967);
or U13558 (N_13558,N_12896,N_13423);
or U13559 (N_13559,N_13166,N_13018);
or U13560 (N_13560,N_13128,N_13445);
nand U13561 (N_13561,N_13146,N_13014);
and U13562 (N_13562,N_13394,N_13431);
or U13563 (N_13563,N_13275,N_13324);
nor U13564 (N_13564,N_13022,N_13362);
and U13565 (N_13565,N_13056,N_12799);
nor U13566 (N_13566,N_12965,N_13200);
nand U13567 (N_13567,N_12801,N_12910);
nand U13568 (N_13568,N_13492,N_13457);
nand U13569 (N_13569,N_13456,N_13098);
nand U13570 (N_13570,N_12859,N_12786);
and U13571 (N_13571,N_13199,N_13135);
nor U13572 (N_13572,N_13144,N_12961);
or U13573 (N_13573,N_12835,N_12929);
and U13574 (N_13574,N_13498,N_12935);
or U13575 (N_13575,N_13183,N_13358);
xor U13576 (N_13576,N_12908,N_12990);
or U13577 (N_13577,N_12836,N_12828);
nand U13578 (N_13578,N_13209,N_12817);
nand U13579 (N_13579,N_13348,N_13310);
and U13580 (N_13580,N_13093,N_13005);
nand U13581 (N_13581,N_13055,N_12814);
nand U13582 (N_13582,N_13157,N_13283);
and U13583 (N_13583,N_13416,N_12976);
nand U13584 (N_13584,N_12995,N_13408);
or U13585 (N_13585,N_13107,N_13409);
and U13586 (N_13586,N_13038,N_13246);
nand U13587 (N_13587,N_13369,N_12823);
nand U13588 (N_13588,N_13193,N_12969);
nand U13589 (N_13589,N_12829,N_12878);
nand U13590 (N_13590,N_13228,N_12834);
nand U13591 (N_13591,N_12764,N_13352);
and U13592 (N_13592,N_12843,N_13090);
or U13593 (N_13593,N_13081,N_13460);
nor U13594 (N_13594,N_13026,N_13286);
and U13595 (N_13595,N_13393,N_13099);
nand U13596 (N_13596,N_12983,N_12771);
or U13597 (N_13597,N_13263,N_12865);
nand U13598 (N_13598,N_13220,N_12947);
xor U13599 (N_13599,N_13360,N_13020);
xnor U13600 (N_13600,N_13258,N_13232);
nand U13601 (N_13601,N_13391,N_12815);
nand U13602 (N_13602,N_13092,N_12959);
xor U13603 (N_13603,N_13328,N_12892);
nor U13604 (N_13604,N_13164,N_13270);
nand U13605 (N_13605,N_12778,N_13268);
nand U13606 (N_13606,N_12755,N_12751);
nor U13607 (N_13607,N_13469,N_13037);
or U13608 (N_13608,N_13036,N_13138);
or U13609 (N_13609,N_13281,N_12862);
nand U13610 (N_13610,N_13397,N_12780);
or U13611 (N_13611,N_13342,N_13405);
nor U13612 (N_13612,N_13426,N_13471);
nand U13613 (N_13613,N_13104,N_12902);
and U13614 (N_13614,N_13453,N_13114);
xor U13615 (N_13615,N_12982,N_12826);
nor U13616 (N_13616,N_12847,N_13145);
nor U13617 (N_13617,N_12797,N_12884);
xnor U13618 (N_13618,N_13279,N_13053);
nand U13619 (N_13619,N_13006,N_13052);
or U13620 (N_13620,N_12962,N_12769);
nand U13621 (N_13621,N_13206,N_12907);
and U13622 (N_13622,N_13087,N_13274);
or U13623 (N_13623,N_12841,N_13194);
nor U13624 (N_13624,N_13390,N_12850);
and U13625 (N_13625,N_13079,N_12812);
nand U13626 (N_13626,N_13155,N_12998);
or U13627 (N_13627,N_12833,N_13221);
nor U13628 (N_13628,N_13051,N_13285);
or U13629 (N_13629,N_12891,N_13289);
nand U13630 (N_13630,N_12760,N_13485);
or U13631 (N_13631,N_13011,N_12880);
xnor U13632 (N_13632,N_12942,N_13337);
nor U13633 (N_13633,N_13095,N_13300);
nor U13634 (N_13634,N_12920,N_13196);
xor U13635 (N_13635,N_13260,N_12928);
nor U13636 (N_13636,N_13265,N_12827);
nand U13637 (N_13637,N_13370,N_13229);
xor U13638 (N_13638,N_13424,N_13311);
nand U13639 (N_13639,N_12779,N_13168);
or U13640 (N_13640,N_12845,N_13217);
nor U13641 (N_13641,N_12972,N_13421);
xor U13642 (N_13642,N_12772,N_12978);
and U13643 (N_13643,N_13284,N_12796);
or U13644 (N_13644,N_13455,N_12870);
and U13645 (N_13645,N_12893,N_13385);
and U13646 (N_13646,N_12840,N_12816);
nand U13647 (N_13647,N_13293,N_13466);
nor U13648 (N_13648,N_13115,N_12770);
xnor U13649 (N_13649,N_12871,N_13216);
and U13650 (N_13650,N_13117,N_13179);
nand U13651 (N_13651,N_12858,N_13187);
nor U13652 (N_13652,N_13475,N_13338);
or U13653 (N_13653,N_12773,N_13459);
or U13654 (N_13654,N_13126,N_13262);
and U13655 (N_13655,N_13015,N_13165);
or U13656 (N_13656,N_13282,N_13080);
nor U13657 (N_13657,N_13483,N_13186);
xor U13658 (N_13658,N_12919,N_12811);
nand U13659 (N_13659,N_13354,N_13302);
xnor U13660 (N_13660,N_13241,N_12977);
and U13661 (N_13661,N_13230,N_13054);
and U13662 (N_13662,N_12963,N_12948);
nor U13663 (N_13663,N_13479,N_13350);
and U13664 (N_13664,N_13131,N_13074);
xnor U13665 (N_13665,N_13150,N_12974);
and U13666 (N_13666,N_13325,N_13103);
or U13667 (N_13667,N_13227,N_13250);
xnor U13668 (N_13668,N_13212,N_13499);
nor U13669 (N_13669,N_12958,N_12857);
or U13670 (N_13670,N_12927,N_13143);
or U13671 (N_13671,N_13004,N_12904);
nand U13672 (N_13672,N_12943,N_13151);
and U13673 (N_13673,N_13491,N_13041);
xnor U13674 (N_13674,N_12992,N_13288);
nor U13675 (N_13675,N_13487,N_13139);
and U13676 (N_13676,N_12852,N_13123);
nand U13677 (N_13677,N_12973,N_13176);
and U13678 (N_13678,N_12877,N_12867);
xnor U13679 (N_13679,N_13410,N_13432);
or U13680 (N_13680,N_13047,N_13490);
xnor U13681 (N_13681,N_13443,N_12750);
nor U13682 (N_13682,N_13366,N_13320);
or U13683 (N_13683,N_13441,N_13259);
and U13684 (N_13684,N_12794,N_13240);
nand U13685 (N_13685,N_13442,N_13048);
xnor U13686 (N_13686,N_12945,N_13468);
nor U13687 (N_13687,N_13321,N_12876);
and U13688 (N_13688,N_13452,N_13253);
or U13689 (N_13689,N_13100,N_12754);
nand U13690 (N_13690,N_13294,N_13428);
nor U13691 (N_13691,N_13153,N_13213);
or U13692 (N_13692,N_12981,N_12916);
and U13693 (N_13693,N_13322,N_13210);
nor U13694 (N_13694,N_13306,N_13458);
nand U13695 (N_13695,N_13025,N_13075);
nand U13696 (N_13696,N_12824,N_13180);
nand U13697 (N_13697,N_13305,N_13007);
and U13698 (N_13698,N_13031,N_13190);
nand U13699 (N_13699,N_13017,N_13386);
nand U13700 (N_13700,N_12854,N_13415);
and U13701 (N_13701,N_12885,N_13272);
and U13702 (N_13702,N_12886,N_13335);
nand U13703 (N_13703,N_12864,N_12951);
or U13704 (N_13704,N_13309,N_13344);
or U13705 (N_13705,N_13198,N_12781);
nand U13706 (N_13706,N_13425,N_13231);
nor U13707 (N_13707,N_12952,N_13069);
and U13708 (N_13708,N_13255,N_13450);
and U13709 (N_13709,N_13349,N_13363);
and U13710 (N_13710,N_13163,N_13112);
nor U13711 (N_13711,N_13182,N_12873);
nor U13712 (N_13712,N_13152,N_12968);
nor U13713 (N_13713,N_13197,N_13361);
and U13714 (N_13714,N_13108,N_13298);
and U13715 (N_13715,N_12846,N_12890);
nor U13716 (N_13716,N_13030,N_13438);
nor U13717 (N_13717,N_12985,N_13067);
and U13718 (N_13718,N_13429,N_13313);
nor U13719 (N_13719,N_13189,N_13096);
and U13720 (N_13720,N_13448,N_13059);
and U13721 (N_13721,N_13029,N_13440);
or U13722 (N_13722,N_13418,N_13000);
nand U13723 (N_13723,N_13046,N_13218);
or U13724 (N_13724,N_13173,N_12777);
or U13725 (N_13725,N_12785,N_13433);
or U13726 (N_13726,N_13111,N_13172);
and U13727 (N_13727,N_12930,N_12894);
and U13728 (N_13728,N_13402,N_13171);
or U13729 (N_13729,N_13470,N_12954);
nand U13730 (N_13730,N_13211,N_12793);
xnor U13731 (N_13731,N_13188,N_13378);
nand U13732 (N_13732,N_13065,N_13336);
nand U13733 (N_13733,N_12795,N_13244);
or U13734 (N_13734,N_12790,N_12955);
xnor U13735 (N_13735,N_12808,N_13243);
or U13736 (N_13736,N_13223,N_13488);
nand U13737 (N_13737,N_13280,N_13071);
nand U13738 (N_13738,N_13027,N_13195);
nand U13739 (N_13739,N_13484,N_13435);
and U13740 (N_13740,N_13473,N_13381);
and U13741 (N_13741,N_12975,N_13383);
or U13742 (N_13742,N_12933,N_13449);
nor U13743 (N_13743,N_13271,N_13478);
nor U13744 (N_13744,N_13446,N_13192);
nor U13745 (N_13745,N_13238,N_13323);
xnor U13746 (N_13746,N_13364,N_13299);
nand U13747 (N_13747,N_13021,N_12895);
and U13748 (N_13748,N_12924,N_12821);
nand U13749 (N_13749,N_13042,N_13436);
xnor U13750 (N_13750,N_13091,N_12788);
nand U13751 (N_13751,N_13148,N_13461);
and U13752 (N_13752,N_13489,N_13267);
and U13753 (N_13753,N_13001,N_12805);
and U13754 (N_13754,N_12986,N_12832);
and U13755 (N_13755,N_13043,N_13057);
or U13756 (N_13756,N_12932,N_13304);
nand U13757 (N_13757,N_13045,N_13137);
nor U13758 (N_13758,N_12783,N_13129);
xor U13759 (N_13759,N_12848,N_13252);
and U13760 (N_13760,N_13033,N_13159);
and U13761 (N_13761,N_12922,N_12837);
and U13762 (N_13762,N_13382,N_13039);
xor U13763 (N_13763,N_13340,N_12861);
and U13764 (N_13764,N_13346,N_12820);
xor U13765 (N_13765,N_12903,N_13451);
and U13766 (N_13766,N_13308,N_13070);
nand U13767 (N_13767,N_12810,N_13292);
nor U13768 (N_13768,N_13444,N_13102);
nand U13769 (N_13769,N_13149,N_13472);
nor U13770 (N_13770,N_13404,N_12766);
nand U13771 (N_13771,N_12996,N_13064);
nand U13772 (N_13772,N_12761,N_13356);
or U13773 (N_13773,N_12937,N_12901);
nand U13774 (N_13774,N_13127,N_13261);
nand U13775 (N_13775,N_13496,N_12762);
nor U13776 (N_13776,N_12957,N_13406);
nor U13777 (N_13777,N_13156,N_13035);
and U13778 (N_13778,N_13395,N_13040);
nand U13779 (N_13779,N_12979,N_13136);
xnor U13780 (N_13780,N_12806,N_13264);
or U13781 (N_13781,N_13332,N_12774);
or U13782 (N_13782,N_13008,N_12888);
nor U13783 (N_13783,N_13407,N_12882);
nand U13784 (N_13784,N_13437,N_13400);
or U13785 (N_13785,N_13247,N_13482);
and U13786 (N_13786,N_13376,N_13411);
nand U13787 (N_13787,N_12789,N_12758);
and U13788 (N_13788,N_12874,N_12875);
nand U13789 (N_13789,N_13118,N_13375);
nand U13790 (N_13790,N_12905,N_13239);
xor U13791 (N_13791,N_13278,N_13009);
nand U13792 (N_13792,N_13277,N_13347);
or U13793 (N_13793,N_13388,N_13477);
and U13794 (N_13794,N_13316,N_13447);
nand U13795 (N_13795,N_13493,N_12763);
xnor U13796 (N_13796,N_12984,N_12830);
nand U13797 (N_13797,N_12988,N_12912);
nor U13798 (N_13798,N_12994,N_13130);
or U13799 (N_13799,N_13464,N_13315);
nand U13800 (N_13800,N_12921,N_13301);
nand U13801 (N_13801,N_13086,N_12776);
nand U13802 (N_13802,N_13105,N_13462);
nand U13803 (N_13803,N_13303,N_13063);
and U13804 (N_13804,N_13439,N_13384);
nand U13805 (N_13805,N_13097,N_13392);
nor U13806 (N_13806,N_12911,N_13225);
nor U13807 (N_13807,N_13226,N_13122);
nor U13808 (N_13808,N_12866,N_12926);
or U13809 (N_13809,N_13120,N_12936);
nor U13810 (N_13810,N_12917,N_13242);
nand U13811 (N_13811,N_12819,N_12950);
and U13812 (N_13812,N_13204,N_12906);
and U13813 (N_13813,N_13248,N_13389);
nand U13814 (N_13814,N_13161,N_13058);
or U13815 (N_13815,N_13224,N_13109);
nor U13816 (N_13816,N_13401,N_12897);
nor U13817 (N_13817,N_13317,N_13184);
nor U13818 (N_13818,N_13016,N_12944);
xor U13819 (N_13819,N_12989,N_13351);
or U13820 (N_13820,N_13367,N_12842);
nand U13821 (N_13821,N_12863,N_12960);
and U13822 (N_13822,N_12971,N_13414);
and U13823 (N_13823,N_12966,N_13205);
or U13824 (N_13824,N_12782,N_13330);
or U13825 (N_13825,N_13201,N_13170);
xnor U13826 (N_13826,N_13276,N_13094);
nand U13827 (N_13827,N_13177,N_12993);
nand U13828 (N_13828,N_13119,N_13141);
or U13829 (N_13829,N_12946,N_13181);
nor U13830 (N_13830,N_13110,N_13167);
nand U13831 (N_13831,N_12757,N_13072);
nand U13832 (N_13832,N_12802,N_13327);
and U13833 (N_13833,N_13089,N_12970);
or U13834 (N_13834,N_13085,N_13480);
and U13835 (N_13835,N_13178,N_12956);
nand U13836 (N_13836,N_13162,N_13237);
or U13837 (N_13837,N_12980,N_13191);
and U13838 (N_13838,N_13236,N_13266);
nand U13839 (N_13839,N_13341,N_13154);
nor U13840 (N_13840,N_12999,N_13379);
or U13841 (N_13841,N_13291,N_13044);
xnor U13842 (N_13842,N_13374,N_13319);
nor U13843 (N_13843,N_13396,N_13269);
xor U13844 (N_13844,N_13312,N_13368);
nor U13845 (N_13845,N_13326,N_13061);
or U13846 (N_13846,N_13134,N_12913);
or U13847 (N_13847,N_12887,N_12899);
nor U13848 (N_13848,N_13140,N_13073);
and U13849 (N_13849,N_13318,N_13207);
and U13850 (N_13850,N_12938,N_13329);
and U13851 (N_13851,N_13417,N_12822);
nor U13852 (N_13852,N_13373,N_13214);
nor U13853 (N_13853,N_13101,N_12872);
and U13854 (N_13854,N_13160,N_13174);
nor U13855 (N_13855,N_12753,N_12809);
or U13856 (N_13856,N_13034,N_13454);
nor U13857 (N_13857,N_12923,N_13295);
nor U13858 (N_13858,N_13133,N_13359);
nand U13859 (N_13859,N_13023,N_13219);
and U13860 (N_13860,N_12804,N_12784);
or U13861 (N_13861,N_13387,N_13251);
nand U13862 (N_13862,N_12853,N_13287);
nor U13863 (N_13863,N_13076,N_12792);
or U13864 (N_13864,N_13077,N_13307);
and U13865 (N_13865,N_12934,N_12909);
nand U13866 (N_13866,N_12953,N_13169);
nand U13867 (N_13867,N_12855,N_13495);
nor U13868 (N_13868,N_13062,N_12889);
or U13869 (N_13869,N_13333,N_13481);
xor U13870 (N_13870,N_12860,N_12925);
or U13871 (N_13871,N_13419,N_13377);
nor U13872 (N_13872,N_13290,N_13132);
xor U13873 (N_13873,N_13427,N_13420);
or U13874 (N_13874,N_13083,N_13068);
nand U13875 (N_13875,N_13472,N_12961);
nor U13876 (N_13876,N_12836,N_13447);
or U13877 (N_13877,N_13205,N_12949);
nor U13878 (N_13878,N_12872,N_13295);
nor U13879 (N_13879,N_12980,N_13445);
or U13880 (N_13880,N_12819,N_13231);
and U13881 (N_13881,N_13456,N_13197);
nor U13882 (N_13882,N_13108,N_13088);
and U13883 (N_13883,N_13461,N_13444);
xnor U13884 (N_13884,N_13392,N_13141);
nand U13885 (N_13885,N_13089,N_12952);
or U13886 (N_13886,N_13023,N_12871);
nand U13887 (N_13887,N_13397,N_13413);
nor U13888 (N_13888,N_12840,N_13413);
nand U13889 (N_13889,N_13024,N_12990);
nand U13890 (N_13890,N_13232,N_12874);
or U13891 (N_13891,N_12859,N_13058);
and U13892 (N_13892,N_13078,N_13011);
nor U13893 (N_13893,N_12881,N_13339);
or U13894 (N_13894,N_13392,N_12836);
nand U13895 (N_13895,N_13147,N_13273);
and U13896 (N_13896,N_13034,N_12949);
nand U13897 (N_13897,N_12823,N_13467);
and U13898 (N_13898,N_12795,N_13398);
and U13899 (N_13899,N_13274,N_13367);
nand U13900 (N_13900,N_13238,N_12947);
nor U13901 (N_13901,N_13115,N_13086);
nor U13902 (N_13902,N_13268,N_13314);
nor U13903 (N_13903,N_13126,N_12942);
or U13904 (N_13904,N_13353,N_12962);
xor U13905 (N_13905,N_13262,N_13471);
nand U13906 (N_13906,N_12854,N_13194);
and U13907 (N_13907,N_13109,N_12859);
nor U13908 (N_13908,N_13167,N_12887);
and U13909 (N_13909,N_13290,N_13198);
nor U13910 (N_13910,N_13259,N_13152);
nor U13911 (N_13911,N_13253,N_13413);
or U13912 (N_13912,N_13001,N_13097);
or U13913 (N_13913,N_12778,N_13378);
or U13914 (N_13914,N_12961,N_13048);
and U13915 (N_13915,N_12899,N_13033);
nor U13916 (N_13916,N_12870,N_12969);
and U13917 (N_13917,N_13412,N_12897);
nor U13918 (N_13918,N_12993,N_13443);
and U13919 (N_13919,N_12984,N_12802);
xnor U13920 (N_13920,N_13243,N_13260);
nor U13921 (N_13921,N_13399,N_13059);
xor U13922 (N_13922,N_12925,N_13113);
or U13923 (N_13923,N_13497,N_12832);
nand U13924 (N_13924,N_13381,N_13235);
nand U13925 (N_13925,N_12822,N_13180);
or U13926 (N_13926,N_13221,N_13060);
nor U13927 (N_13927,N_12899,N_12969);
or U13928 (N_13928,N_13221,N_13137);
nand U13929 (N_13929,N_13430,N_13018);
or U13930 (N_13930,N_12799,N_13395);
or U13931 (N_13931,N_13093,N_13102);
and U13932 (N_13932,N_13325,N_12987);
or U13933 (N_13933,N_13207,N_13386);
nand U13934 (N_13934,N_13205,N_12860);
nor U13935 (N_13935,N_13139,N_13176);
or U13936 (N_13936,N_13350,N_13261);
or U13937 (N_13937,N_13202,N_13353);
nand U13938 (N_13938,N_13266,N_13293);
or U13939 (N_13939,N_13303,N_13337);
and U13940 (N_13940,N_13451,N_13190);
nor U13941 (N_13941,N_13498,N_13139);
nor U13942 (N_13942,N_13064,N_12947);
or U13943 (N_13943,N_13331,N_12976);
and U13944 (N_13944,N_12851,N_12871);
nor U13945 (N_13945,N_12854,N_13378);
nor U13946 (N_13946,N_13328,N_13158);
and U13947 (N_13947,N_12995,N_12967);
or U13948 (N_13948,N_12952,N_13496);
nand U13949 (N_13949,N_12849,N_13355);
and U13950 (N_13950,N_13461,N_12817);
xnor U13951 (N_13951,N_13038,N_13144);
nand U13952 (N_13952,N_13375,N_13373);
and U13953 (N_13953,N_13039,N_12877);
nor U13954 (N_13954,N_13387,N_12751);
xnor U13955 (N_13955,N_12869,N_13042);
nand U13956 (N_13956,N_12797,N_13464);
or U13957 (N_13957,N_13247,N_13230);
nand U13958 (N_13958,N_13221,N_13019);
nand U13959 (N_13959,N_13433,N_13100);
or U13960 (N_13960,N_12952,N_12794);
nor U13961 (N_13961,N_13369,N_12867);
xor U13962 (N_13962,N_12874,N_13063);
nor U13963 (N_13963,N_12927,N_13129);
or U13964 (N_13964,N_13294,N_13004);
nand U13965 (N_13965,N_13373,N_13147);
or U13966 (N_13966,N_13089,N_13443);
nor U13967 (N_13967,N_13261,N_13222);
xnor U13968 (N_13968,N_13454,N_13390);
xnor U13969 (N_13969,N_13319,N_12947);
nor U13970 (N_13970,N_12820,N_12856);
nor U13971 (N_13971,N_12990,N_12947);
xor U13972 (N_13972,N_12783,N_13018);
xnor U13973 (N_13973,N_13019,N_13205);
or U13974 (N_13974,N_12759,N_13199);
xnor U13975 (N_13975,N_13071,N_13126);
xnor U13976 (N_13976,N_13249,N_13419);
nand U13977 (N_13977,N_12905,N_12860);
nand U13978 (N_13978,N_13269,N_13144);
nor U13979 (N_13979,N_13347,N_13069);
nand U13980 (N_13980,N_12860,N_13022);
nand U13981 (N_13981,N_13498,N_13486);
xnor U13982 (N_13982,N_13098,N_12922);
or U13983 (N_13983,N_12781,N_12786);
nor U13984 (N_13984,N_13143,N_13184);
and U13985 (N_13985,N_13492,N_12920);
or U13986 (N_13986,N_12931,N_13382);
or U13987 (N_13987,N_13134,N_13220);
or U13988 (N_13988,N_13419,N_12993);
or U13989 (N_13989,N_13369,N_12939);
or U13990 (N_13990,N_12773,N_13203);
nand U13991 (N_13991,N_12767,N_13076);
nand U13992 (N_13992,N_13085,N_13342);
nor U13993 (N_13993,N_13158,N_13127);
and U13994 (N_13994,N_12907,N_13231);
xnor U13995 (N_13995,N_13435,N_13361);
and U13996 (N_13996,N_13006,N_12778);
nor U13997 (N_13997,N_13167,N_13436);
nor U13998 (N_13998,N_13050,N_13488);
nand U13999 (N_13999,N_13032,N_13291);
or U14000 (N_14000,N_12852,N_13345);
and U14001 (N_14001,N_13242,N_13255);
nor U14002 (N_14002,N_13235,N_12919);
nand U14003 (N_14003,N_12904,N_12870);
nand U14004 (N_14004,N_13132,N_13229);
or U14005 (N_14005,N_13170,N_13479);
nor U14006 (N_14006,N_13175,N_12965);
or U14007 (N_14007,N_13272,N_13193);
or U14008 (N_14008,N_13137,N_13041);
or U14009 (N_14009,N_12770,N_12888);
or U14010 (N_14010,N_13047,N_13384);
or U14011 (N_14011,N_13220,N_13034);
or U14012 (N_14012,N_12897,N_13343);
and U14013 (N_14013,N_12965,N_12873);
or U14014 (N_14014,N_12776,N_13027);
and U14015 (N_14015,N_13128,N_12935);
xnor U14016 (N_14016,N_13413,N_13436);
nand U14017 (N_14017,N_13049,N_13204);
nand U14018 (N_14018,N_13436,N_12959);
nand U14019 (N_14019,N_13215,N_13421);
nand U14020 (N_14020,N_12800,N_13038);
nand U14021 (N_14021,N_13406,N_13176);
nand U14022 (N_14022,N_12959,N_12750);
and U14023 (N_14023,N_13153,N_13173);
nand U14024 (N_14024,N_12757,N_12869);
or U14025 (N_14025,N_13211,N_13260);
nor U14026 (N_14026,N_13148,N_12760);
nand U14027 (N_14027,N_13244,N_12910);
nand U14028 (N_14028,N_13200,N_13440);
or U14029 (N_14029,N_13446,N_13302);
nor U14030 (N_14030,N_12862,N_13041);
and U14031 (N_14031,N_13322,N_13427);
or U14032 (N_14032,N_12886,N_13033);
or U14033 (N_14033,N_12910,N_13321);
or U14034 (N_14034,N_12823,N_13390);
and U14035 (N_14035,N_13171,N_13249);
or U14036 (N_14036,N_13372,N_13454);
nor U14037 (N_14037,N_12986,N_12759);
xnor U14038 (N_14038,N_13283,N_12924);
or U14039 (N_14039,N_13009,N_13242);
nor U14040 (N_14040,N_12961,N_13054);
and U14041 (N_14041,N_13051,N_13361);
nand U14042 (N_14042,N_12837,N_13442);
nor U14043 (N_14043,N_13134,N_13394);
or U14044 (N_14044,N_12773,N_12992);
and U14045 (N_14045,N_13327,N_12996);
and U14046 (N_14046,N_12984,N_13002);
xor U14047 (N_14047,N_13439,N_13310);
or U14048 (N_14048,N_12957,N_13485);
nand U14049 (N_14049,N_13082,N_13099);
nand U14050 (N_14050,N_12945,N_13080);
or U14051 (N_14051,N_12995,N_12768);
or U14052 (N_14052,N_12973,N_13355);
or U14053 (N_14053,N_12948,N_13006);
or U14054 (N_14054,N_13142,N_13079);
or U14055 (N_14055,N_13058,N_12822);
and U14056 (N_14056,N_13189,N_13266);
or U14057 (N_14057,N_13369,N_13138);
xor U14058 (N_14058,N_13431,N_13076);
and U14059 (N_14059,N_13305,N_13006);
or U14060 (N_14060,N_12895,N_12763);
or U14061 (N_14061,N_13365,N_13333);
and U14062 (N_14062,N_12929,N_13119);
or U14063 (N_14063,N_13130,N_13169);
and U14064 (N_14064,N_13255,N_12779);
nor U14065 (N_14065,N_13227,N_13286);
or U14066 (N_14066,N_13379,N_13437);
nor U14067 (N_14067,N_13144,N_12970);
or U14068 (N_14068,N_13410,N_12996);
and U14069 (N_14069,N_13417,N_12857);
and U14070 (N_14070,N_12770,N_12848);
or U14071 (N_14071,N_13145,N_13443);
nand U14072 (N_14072,N_12926,N_13459);
nand U14073 (N_14073,N_13162,N_13312);
nor U14074 (N_14074,N_12909,N_13197);
nand U14075 (N_14075,N_13077,N_13036);
or U14076 (N_14076,N_13415,N_13358);
nor U14077 (N_14077,N_13481,N_13397);
or U14078 (N_14078,N_13388,N_13116);
nor U14079 (N_14079,N_13130,N_13110);
nor U14080 (N_14080,N_13406,N_12817);
nand U14081 (N_14081,N_13391,N_13491);
and U14082 (N_14082,N_12772,N_13452);
or U14083 (N_14083,N_12862,N_13394);
nor U14084 (N_14084,N_12930,N_13013);
nor U14085 (N_14085,N_13299,N_13442);
nor U14086 (N_14086,N_13229,N_13122);
and U14087 (N_14087,N_13485,N_13198);
and U14088 (N_14088,N_12858,N_13335);
nor U14089 (N_14089,N_13110,N_12951);
nand U14090 (N_14090,N_12969,N_13414);
nand U14091 (N_14091,N_13344,N_12962);
nand U14092 (N_14092,N_12881,N_13172);
or U14093 (N_14093,N_12915,N_13300);
nand U14094 (N_14094,N_12887,N_12814);
and U14095 (N_14095,N_13080,N_13228);
nand U14096 (N_14096,N_12779,N_12848);
nand U14097 (N_14097,N_12978,N_13215);
and U14098 (N_14098,N_13182,N_13395);
and U14099 (N_14099,N_13064,N_13144);
xor U14100 (N_14100,N_13416,N_12820);
or U14101 (N_14101,N_13095,N_13191);
nor U14102 (N_14102,N_13096,N_13466);
or U14103 (N_14103,N_12799,N_13387);
and U14104 (N_14104,N_13090,N_13361);
xnor U14105 (N_14105,N_13139,N_12942);
or U14106 (N_14106,N_13446,N_13497);
or U14107 (N_14107,N_12909,N_13052);
and U14108 (N_14108,N_13094,N_13438);
nor U14109 (N_14109,N_13185,N_13335);
nor U14110 (N_14110,N_13391,N_13178);
nor U14111 (N_14111,N_13154,N_13236);
or U14112 (N_14112,N_13276,N_12999);
nand U14113 (N_14113,N_13363,N_13188);
or U14114 (N_14114,N_13082,N_13391);
and U14115 (N_14115,N_12792,N_12767);
or U14116 (N_14116,N_13402,N_12937);
xor U14117 (N_14117,N_13078,N_12773);
or U14118 (N_14118,N_13069,N_13107);
and U14119 (N_14119,N_13051,N_13085);
nand U14120 (N_14120,N_12824,N_12842);
nand U14121 (N_14121,N_13202,N_13034);
nand U14122 (N_14122,N_13349,N_12832);
xnor U14123 (N_14123,N_13404,N_13490);
nand U14124 (N_14124,N_12909,N_12929);
nand U14125 (N_14125,N_13447,N_13267);
nand U14126 (N_14126,N_12850,N_13460);
nor U14127 (N_14127,N_12991,N_12948);
or U14128 (N_14128,N_12766,N_13106);
nand U14129 (N_14129,N_13218,N_12820);
nor U14130 (N_14130,N_12799,N_13335);
or U14131 (N_14131,N_12754,N_12845);
and U14132 (N_14132,N_13073,N_13428);
or U14133 (N_14133,N_12871,N_13185);
nand U14134 (N_14134,N_13412,N_13020);
nand U14135 (N_14135,N_13018,N_13093);
xor U14136 (N_14136,N_13315,N_13152);
nand U14137 (N_14137,N_13221,N_13284);
and U14138 (N_14138,N_13455,N_13223);
nor U14139 (N_14139,N_13095,N_13342);
xor U14140 (N_14140,N_13199,N_12827);
or U14141 (N_14141,N_13230,N_12957);
nor U14142 (N_14142,N_12937,N_13455);
nand U14143 (N_14143,N_13049,N_13272);
nor U14144 (N_14144,N_13201,N_12864);
or U14145 (N_14145,N_13329,N_12772);
or U14146 (N_14146,N_13343,N_12885);
nand U14147 (N_14147,N_13012,N_13471);
nor U14148 (N_14148,N_13396,N_13149);
nand U14149 (N_14149,N_13308,N_13007);
and U14150 (N_14150,N_13313,N_12784);
and U14151 (N_14151,N_12754,N_13110);
and U14152 (N_14152,N_12827,N_13177);
nand U14153 (N_14153,N_13086,N_12929);
nand U14154 (N_14154,N_12984,N_12760);
nor U14155 (N_14155,N_13209,N_13385);
nor U14156 (N_14156,N_13363,N_12760);
or U14157 (N_14157,N_12877,N_12981);
and U14158 (N_14158,N_12925,N_12945);
nor U14159 (N_14159,N_13208,N_13186);
and U14160 (N_14160,N_13289,N_13466);
nor U14161 (N_14161,N_12909,N_12938);
nand U14162 (N_14162,N_13012,N_12975);
nor U14163 (N_14163,N_13076,N_13238);
or U14164 (N_14164,N_13214,N_13391);
xnor U14165 (N_14165,N_12848,N_13408);
and U14166 (N_14166,N_13042,N_13066);
nand U14167 (N_14167,N_13331,N_13370);
or U14168 (N_14168,N_13412,N_12804);
and U14169 (N_14169,N_13064,N_13109);
and U14170 (N_14170,N_13047,N_13213);
nand U14171 (N_14171,N_13332,N_12760);
and U14172 (N_14172,N_13136,N_12937);
nand U14173 (N_14173,N_12903,N_12816);
nor U14174 (N_14174,N_12868,N_12762);
nor U14175 (N_14175,N_12848,N_13279);
nor U14176 (N_14176,N_13421,N_13241);
nor U14177 (N_14177,N_13397,N_13495);
nor U14178 (N_14178,N_13423,N_12809);
nand U14179 (N_14179,N_13082,N_13285);
xor U14180 (N_14180,N_12796,N_12993);
nand U14181 (N_14181,N_13388,N_12938);
and U14182 (N_14182,N_13203,N_13069);
or U14183 (N_14183,N_13301,N_12925);
xor U14184 (N_14184,N_12987,N_13394);
or U14185 (N_14185,N_13012,N_12863);
nand U14186 (N_14186,N_13387,N_13289);
nor U14187 (N_14187,N_13492,N_13346);
xnor U14188 (N_14188,N_13097,N_13042);
nand U14189 (N_14189,N_13211,N_13146);
xor U14190 (N_14190,N_13386,N_12871);
and U14191 (N_14191,N_13293,N_12904);
and U14192 (N_14192,N_12970,N_13094);
nor U14193 (N_14193,N_13080,N_12853);
and U14194 (N_14194,N_13035,N_13480);
and U14195 (N_14195,N_13393,N_13322);
and U14196 (N_14196,N_13454,N_13074);
xor U14197 (N_14197,N_13467,N_13190);
nand U14198 (N_14198,N_13284,N_13248);
nand U14199 (N_14199,N_12941,N_12928);
xor U14200 (N_14200,N_13331,N_13338);
or U14201 (N_14201,N_13281,N_13267);
nor U14202 (N_14202,N_12850,N_13477);
nor U14203 (N_14203,N_13463,N_13079);
nand U14204 (N_14204,N_13109,N_12960);
or U14205 (N_14205,N_12990,N_13075);
xnor U14206 (N_14206,N_13147,N_13087);
nor U14207 (N_14207,N_13203,N_12910);
and U14208 (N_14208,N_13119,N_12753);
nor U14209 (N_14209,N_13244,N_12872);
or U14210 (N_14210,N_13288,N_13480);
and U14211 (N_14211,N_13119,N_12822);
or U14212 (N_14212,N_12903,N_13374);
and U14213 (N_14213,N_13280,N_12981);
and U14214 (N_14214,N_13030,N_12804);
and U14215 (N_14215,N_13387,N_13213);
or U14216 (N_14216,N_13314,N_13180);
nor U14217 (N_14217,N_13415,N_13444);
and U14218 (N_14218,N_12761,N_13221);
nor U14219 (N_14219,N_13491,N_12830);
nor U14220 (N_14220,N_12978,N_12942);
nor U14221 (N_14221,N_12793,N_13021);
nand U14222 (N_14222,N_13310,N_13226);
nor U14223 (N_14223,N_13297,N_13398);
nand U14224 (N_14224,N_12880,N_13005);
nand U14225 (N_14225,N_12971,N_12917);
or U14226 (N_14226,N_13057,N_12865);
nor U14227 (N_14227,N_12949,N_13476);
nor U14228 (N_14228,N_13296,N_13061);
and U14229 (N_14229,N_13058,N_13166);
nor U14230 (N_14230,N_13271,N_13291);
or U14231 (N_14231,N_12905,N_13431);
and U14232 (N_14232,N_13322,N_12862);
nand U14233 (N_14233,N_12817,N_12938);
nor U14234 (N_14234,N_13289,N_12853);
or U14235 (N_14235,N_12978,N_13013);
nand U14236 (N_14236,N_12862,N_12932);
and U14237 (N_14237,N_13231,N_12794);
nand U14238 (N_14238,N_12797,N_12810);
xor U14239 (N_14239,N_12885,N_13253);
or U14240 (N_14240,N_13492,N_13264);
or U14241 (N_14241,N_13430,N_13150);
xnor U14242 (N_14242,N_12751,N_12857);
xnor U14243 (N_14243,N_12799,N_12907);
nor U14244 (N_14244,N_13388,N_13499);
nor U14245 (N_14245,N_13286,N_13347);
and U14246 (N_14246,N_12985,N_13420);
or U14247 (N_14247,N_12863,N_13089);
nor U14248 (N_14248,N_13496,N_13434);
nor U14249 (N_14249,N_13475,N_12784);
xor U14250 (N_14250,N_13872,N_13956);
nor U14251 (N_14251,N_13774,N_13761);
nand U14252 (N_14252,N_13942,N_13522);
and U14253 (N_14253,N_13706,N_13543);
nor U14254 (N_14254,N_13911,N_13574);
or U14255 (N_14255,N_13863,N_14091);
nor U14256 (N_14256,N_14068,N_13675);
and U14257 (N_14257,N_13728,N_14193);
xor U14258 (N_14258,N_14047,N_14229);
nor U14259 (N_14259,N_13925,N_14206);
nand U14260 (N_14260,N_13869,N_14156);
nand U14261 (N_14261,N_14248,N_13739);
nand U14262 (N_14262,N_13998,N_13825);
nor U14263 (N_14263,N_13818,N_13717);
and U14264 (N_14264,N_13832,N_13900);
nor U14265 (N_14265,N_13539,N_13636);
or U14266 (N_14266,N_14028,N_14109);
nand U14267 (N_14267,N_13614,N_13866);
or U14268 (N_14268,N_13947,N_14197);
nor U14269 (N_14269,N_14040,N_13561);
and U14270 (N_14270,N_13784,N_13674);
nand U14271 (N_14271,N_13792,N_13606);
nor U14272 (N_14272,N_14086,N_13898);
or U14273 (N_14273,N_13546,N_14118);
xor U14274 (N_14274,N_13989,N_14112);
nor U14275 (N_14275,N_13723,N_13757);
and U14276 (N_14276,N_14228,N_13782);
or U14277 (N_14277,N_13957,N_13994);
nor U14278 (N_14278,N_14236,N_14191);
nand U14279 (N_14279,N_13908,N_13831);
or U14280 (N_14280,N_13565,N_13875);
nand U14281 (N_14281,N_13977,N_13979);
xor U14282 (N_14282,N_13530,N_13852);
and U14283 (N_14283,N_13807,N_14108);
nor U14284 (N_14284,N_13993,N_13573);
xnor U14285 (N_14285,N_13927,N_13581);
nand U14286 (N_14286,N_14131,N_14064);
nor U14287 (N_14287,N_14085,N_13755);
nand U14288 (N_14288,N_13625,N_14221);
nand U14289 (N_14289,N_13973,N_13524);
and U14290 (N_14290,N_13858,N_14102);
xor U14291 (N_14291,N_13868,N_13634);
or U14292 (N_14292,N_13732,N_13926);
nand U14293 (N_14293,N_13638,N_13748);
or U14294 (N_14294,N_13585,N_14094);
nor U14295 (N_14295,N_14225,N_13859);
nor U14296 (N_14296,N_13809,N_14138);
or U14297 (N_14297,N_14172,N_13735);
nand U14298 (N_14298,N_13895,N_13741);
nand U14299 (N_14299,N_14042,N_14169);
nor U14300 (N_14300,N_13975,N_13824);
and U14301 (N_14301,N_14226,N_13787);
nand U14302 (N_14302,N_13659,N_13929);
nor U14303 (N_14303,N_13579,N_13963);
or U14304 (N_14304,N_14015,N_13621);
or U14305 (N_14305,N_14135,N_14136);
or U14306 (N_14306,N_13523,N_14182);
or U14307 (N_14307,N_13631,N_13948);
xor U14308 (N_14308,N_13856,N_13580);
and U14309 (N_14309,N_14029,N_13589);
and U14310 (N_14310,N_13557,N_13528);
nand U14311 (N_14311,N_13946,N_13878);
and U14312 (N_14312,N_13701,N_13779);
nor U14313 (N_14313,N_14070,N_13600);
or U14314 (N_14314,N_13976,N_13892);
or U14315 (N_14315,N_13608,N_13940);
or U14316 (N_14316,N_14144,N_13867);
and U14317 (N_14317,N_13775,N_13607);
nor U14318 (N_14318,N_13722,N_14008);
or U14319 (N_14319,N_14035,N_14174);
and U14320 (N_14320,N_14049,N_13844);
nand U14321 (N_14321,N_13584,N_13931);
nor U14322 (N_14322,N_14044,N_13990);
and U14323 (N_14323,N_13810,N_14178);
nor U14324 (N_14324,N_14212,N_14159);
nand U14325 (N_14325,N_13952,N_13758);
nor U14326 (N_14326,N_13747,N_13943);
nand U14327 (N_14327,N_13679,N_14087);
or U14328 (N_14328,N_13899,N_13888);
nor U14329 (N_14329,N_13696,N_13536);
xnor U14330 (N_14330,N_14006,N_14184);
and U14331 (N_14331,N_14198,N_13919);
nand U14332 (N_14332,N_14097,N_13798);
nor U14333 (N_14333,N_13647,N_13501);
or U14334 (N_14334,N_13996,N_13808);
nor U14335 (N_14335,N_13924,N_13874);
and U14336 (N_14336,N_13951,N_14146);
nand U14337 (N_14337,N_13713,N_13843);
nand U14338 (N_14338,N_13937,N_13691);
nor U14339 (N_14339,N_13766,N_14020);
nand U14340 (N_14340,N_14058,N_13750);
and U14341 (N_14341,N_13958,N_13520);
nand U14342 (N_14342,N_13511,N_13563);
and U14343 (N_14343,N_14244,N_13666);
nand U14344 (N_14344,N_13710,N_14100);
xor U14345 (N_14345,N_13752,N_14249);
and U14346 (N_14346,N_13683,N_13693);
xor U14347 (N_14347,N_13971,N_13889);
or U14348 (N_14348,N_13802,N_13778);
nor U14349 (N_14349,N_13588,N_14116);
nor U14350 (N_14350,N_13671,N_13829);
nand U14351 (N_14351,N_14151,N_14195);
nand U14352 (N_14352,N_13639,N_14120);
nor U14353 (N_14353,N_13725,N_14066);
nand U14354 (N_14354,N_13862,N_13734);
or U14355 (N_14355,N_14000,N_14217);
nor U14356 (N_14356,N_13605,N_13918);
or U14357 (N_14357,N_13592,N_14187);
nor U14358 (N_14358,N_13883,N_13813);
nand U14359 (N_14359,N_13737,N_14065);
nor U14360 (N_14360,N_14190,N_13887);
nand U14361 (N_14361,N_13845,N_13804);
or U14362 (N_14362,N_13986,N_14063);
and U14363 (N_14363,N_14034,N_14210);
or U14364 (N_14364,N_14067,N_13707);
and U14365 (N_14365,N_13838,N_14204);
and U14366 (N_14366,N_13527,N_13978);
nand U14367 (N_14367,N_13746,N_13780);
nor U14368 (N_14368,N_13500,N_14001);
and U14369 (N_14369,N_13715,N_13944);
xnor U14370 (N_14370,N_13816,N_13566);
and U14371 (N_14371,N_13901,N_14007);
and U14372 (N_14372,N_14243,N_13587);
or U14373 (N_14373,N_14104,N_13799);
xor U14374 (N_14374,N_13533,N_14232);
and U14375 (N_14375,N_14176,N_13984);
xnor U14376 (N_14376,N_13902,N_13591);
and U14377 (N_14377,N_14211,N_14163);
nand U14378 (N_14378,N_13814,N_14219);
nor U14379 (N_14379,N_13950,N_14186);
and U14380 (N_14380,N_13941,N_13783);
and U14381 (N_14381,N_13609,N_14078);
nand U14382 (N_14382,N_13603,N_14117);
nand U14383 (N_14383,N_13697,N_13554);
nor U14384 (N_14384,N_13815,N_13583);
and U14385 (N_14385,N_14164,N_13712);
and U14386 (N_14386,N_13655,N_13969);
and U14387 (N_14387,N_13938,N_14011);
xnor U14388 (N_14388,N_14084,N_13542);
nor U14389 (N_14389,N_14003,N_14059);
nand U14390 (N_14390,N_13823,N_13578);
nor U14391 (N_14391,N_13801,N_13686);
or U14392 (N_14392,N_13537,N_13716);
and U14393 (N_14393,N_14177,N_13525);
and U14394 (N_14394,N_14194,N_13516);
and U14395 (N_14395,N_14074,N_14062);
and U14396 (N_14396,N_13772,N_13916);
nor U14397 (N_14397,N_13652,N_14129);
or U14398 (N_14398,N_13767,N_13645);
and U14399 (N_14399,N_13670,N_13879);
nor U14400 (N_14400,N_14013,N_13893);
and U14401 (N_14401,N_13514,N_13669);
and U14402 (N_14402,N_14072,N_13885);
and U14403 (N_14403,N_13604,N_14180);
nor U14404 (N_14404,N_13934,N_13930);
and U14405 (N_14405,N_13812,N_13833);
and U14406 (N_14406,N_13544,N_13660);
or U14407 (N_14407,N_14173,N_13548);
xor U14408 (N_14408,N_13905,N_13980);
nor U14409 (N_14409,N_13923,N_13754);
nor U14410 (N_14410,N_14231,N_13515);
and U14411 (N_14411,N_13650,N_13654);
nor U14412 (N_14412,N_14081,N_14125);
and U14413 (N_14413,N_13702,N_13982);
nand U14414 (N_14414,N_13932,N_13850);
nor U14415 (N_14415,N_13623,N_13553);
and U14416 (N_14416,N_13531,N_13611);
or U14417 (N_14417,N_13910,N_13826);
or U14418 (N_14418,N_14237,N_14139);
or U14419 (N_14419,N_14012,N_14128);
or U14420 (N_14420,N_13882,N_13896);
and U14421 (N_14421,N_14205,N_13635);
and U14422 (N_14422,N_13820,N_13502);
nand U14423 (N_14423,N_13762,N_13551);
xnor U14424 (N_14424,N_13742,N_13769);
and U14425 (N_14425,N_13847,N_14199);
nor U14426 (N_14426,N_14046,N_13593);
or U14427 (N_14427,N_13740,N_13630);
nor U14428 (N_14428,N_14132,N_13770);
nor U14429 (N_14429,N_13805,N_13835);
or U14430 (N_14430,N_13997,N_13575);
or U14431 (N_14431,N_13673,N_13595);
nor U14432 (N_14432,N_13785,N_14016);
or U14433 (N_14433,N_13828,N_13756);
xor U14434 (N_14434,N_14113,N_13698);
and U14435 (N_14435,N_14073,N_13620);
nand U14436 (N_14436,N_14238,N_13624);
nand U14437 (N_14437,N_13541,N_13796);
or U14438 (N_14438,N_13837,N_13510);
nor U14439 (N_14439,N_14005,N_13550);
or U14440 (N_14440,N_14235,N_13857);
and U14441 (N_14441,N_14216,N_13724);
or U14442 (N_14442,N_14179,N_14083);
nand U14443 (N_14443,N_14166,N_13649);
nor U14444 (N_14444,N_14121,N_14222);
or U14445 (N_14445,N_14030,N_14014);
nand U14446 (N_14446,N_13598,N_13841);
nor U14447 (N_14447,N_13834,N_13526);
nand U14448 (N_14448,N_13864,N_14089);
nand U14449 (N_14449,N_14230,N_14189);
nor U14450 (N_14450,N_13505,N_13800);
or U14451 (N_14451,N_13955,N_13695);
or U14452 (N_14452,N_13983,N_13676);
nor U14453 (N_14453,N_14201,N_14060);
xnor U14454 (N_14454,N_13771,N_13726);
or U14455 (N_14455,N_13953,N_14162);
and U14456 (N_14456,N_14038,N_13615);
or U14457 (N_14457,N_13791,N_13519);
nor U14458 (N_14458,N_13738,N_14092);
or U14459 (N_14459,N_13653,N_14088);
or U14460 (N_14460,N_14054,N_13504);
nand U14461 (N_14461,N_13777,N_14141);
or U14462 (N_14462,N_13661,N_13933);
and U14463 (N_14463,N_13870,N_13904);
and U14464 (N_14464,N_13719,N_14050);
and U14465 (N_14465,N_13981,N_13995);
and U14466 (N_14466,N_13521,N_13909);
nand U14467 (N_14467,N_14127,N_14140);
and U14468 (N_14468,N_13788,N_13729);
nor U14469 (N_14469,N_14202,N_13599);
nor U14470 (N_14470,N_13632,N_13960);
nand U14471 (N_14471,N_13711,N_13836);
nor U14472 (N_14472,N_14200,N_13821);
nand U14473 (N_14473,N_13936,N_14126);
or U14474 (N_14474,N_14082,N_13744);
nor U14475 (N_14475,N_13861,N_14105);
and U14476 (N_14476,N_13518,N_13643);
and U14477 (N_14477,N_13633,N_13939);
xor U14478 (N_14478,N_13602,N_13840);
or U14479 (N_14479,N_14080,N_13610);
xnor U14480 (N_14480,N_13860,N_14053);
nand U14481 (N_14481,N_13751,N_13648);
nand U14482 (N_14482,N_13912,N_13556);
nor U14483 (N_14483,N_13720,N_13687);
or U14484 (N_14484,N_13705,N_13759);
nand U14485 (N_14485,N_13682,N_13733);
or U14486 (N_14486,N_13590,N_13513);
or U14487 (N_14487,N_13992,N_14158);
xor U14488 (N_14488,N_14234,N_13571);
or U14489 (N_14489,N_13954,N_13891);
nor U14490 (N_14490,N_13506,N_13658);
or U14491 (N_14491,N_14134,N_13640);
or U14492 (N_14492,N_14077,N_13577);
or U14493 (N_14493,N_14165,N_13594);
or U14494 (N_14494,N_13517,N_14185);
nand U14495 (N_14495,N_14036,N_14147);
nor U14496 (N_14496,N_14019,N_14137);
and U14497 (N_14497,N_13651,N_13793);
or U14498 (N_14498,N_13663,N_13622);
nor U14499 (N_14499,N_14213,N_14130);
xor U14500 (N_14500,N_13873,N_13806);
and U14501 (N_14501,N_14076,N_14026);
and U14502 (N_14502,N_13545,N_13700);
or U14503 (N_14503,N_13667,N_13914);
nand U14504 (N_14504,N_13677,N_14240);
or U14505 (N_14505,N_13876,N_13877);
and U14506 (N_14506,N_13672,N_13637);
nand U14507 (N_14507,N_14124,N_14037);
nor U14508 (N_14508,N_14214,N_13681);
or U14509 (N_14509,N_13991,N_13959);
xnor U14510 (N_14510,N_14002,N_13968);
or U14511 (N_14511,N_13985,N_13664);
or U14512 (N_14512,N_14018,N_14167);
and U14513 (N_14513,N_13616,N_13532);
nor U14514 (N_14514,N_14096,N_13830);
nand U14515 (N_14515,N_13678,N_13897);
and U14516 (N_14516,N_14107,N_14192);
nand U14517 (N_14517,N_13657,N_14111);
nor U14518 (N_14518,N_13567,N_13743);
xnor U14519 (N_14519,N_13688,N_13881);
nand U14520 (N_14520,N_13974,N_13558);
nor U14521 (N_14521,N_14069,N_13966);
xnor U14522 (N_14522,N_14239,N_13794);
and U14523 (N_14523,N_14052,N_14142);
nor U14524 (N_14524,N_14041,N_13848);
and U14525 (N_14525,N_13763,N_14150);
nor U14526 (N_14526,N_13646,N_13509);
and U14527 (N_14527,N_14079,N_13851);
xnor U14528 (N_14528,N_14023,N_13721);
or U14529 (N_14529,N_13618,N_13753);
and U14530 (N_14530,N_14057,N_14247);
nor U14531 (N_14531,N_13512,N_13708);
nand U14532 (N_14532,N_14145,N_13964);
or U14533 (N_14533,N_14051,N_13855);
and U14534 (N_14534,N_13827,N_13718);
nor U14535 (N_14535,N_14025,N_13795);
nand U14536 (N_14536,N_13928,N_14021);
and U14537 (N_14537,N_14048,N_14242);
and U14538 (N_14538,N_13736,N_13596);
and U14539 (N_14539,N_13570,N_13662);
and U14540 (N_14540,N_14009,N_13803);
or U14541 (N_14541,N_13680,N_13534);
nand U14542 (N_14542,N_14188,N_14175);
nand U14543 (N_14543,N_14024,N_14061);
and U14544 (N_14544,N_13817,N_13641);
nor U14545 (N_14545,N_14033,N_13920);
nor U14546 (N_14546,N_13962,N_13703);
nor U14547 (N_14547,N_14103,N_14101);
and U14548 (N_14548,N_14039,N_13749);
xor U14549 (N_14549,N_13842,N_14099);
nor U14550 (N_14550,N_14032,N_13789);
nand U14551 (N_14551,N_14161,N_14075);
and U14552 (N_14552,N_13768,N_13538);
xor U14553 (N_14553,N_13764,N_13564);
nor U14554 (N_14554,N_13576,N_14055);
or U14555 (N_14555,N_13540,N_13987);
nand U14556 (N_14556,N_13935,N_13913);
nor U14557 (N_14557,N_14071,N_14017);
nand U14558 (N_14558,N_13601,N_13582);
nor U14559 (N_14559,N_14207,N_14093);
and U14560 (N_14560,N_14220,N_14155);
nor U14561 (N_14561,N_14045,N_13572);
or U14562 (N_14562,N_13945,N_13760);
or U14563 (N_14563,N_13529,N_13790);
and U14564 (N_14564,N_14133,N_14170);
xnor U14565 (N_14565,N_14122,N_13822);
and U14566 (N_14566,N_14241,N_14154);
or U14567 (N_14567,N_14027,N_14149);
and U14568 (N_14568,N_13839,N_13626);
xor U14569 (N_14569,N_14148,N_13507);
nand U14570 (N_14570,N_13886,N_13727);
nand U14571 (N_14571,N_14110,N_13562);
xnor U14572 (N_14572,N_14123,N_13699);
nor U14573 (N_14573,N_13922,N_13628);
nor U14574 (N_14574,N_14143,N_14171);
and U14575 (N_14575,N_13745,N_13907);
and U14576 (N_14576,N_13694,N_13781);
xor U14577 (N_14577,N_13961,N_13846);
nor U14578 (N_14578,N_13586,N_13684);
and U14579 (N_14579,N_14227,N_13965);
and U14580 (N_14580,N_14203,N_13617);
or U14581 (N_14581,N_13568,N_13972);
nor U14582 (N_14582,N_13730,N_14043);
nand U14583 (N_14583,N_13921,N_13915);
xnor U14584 (N_14584,N_14209,N_13704);
or U14585 (N_14585,N_13871,N_14022);
or U14586 (N_14586,N_13890,N_14090);
and U14587 (N_14587,N_14004,N_14183);
or U14588 (N_14588,N_13559,N_13644);
or U14589 (N_14589,N_13549,N_13894);
and U14590 (N_14590,N_13560,N_14098);
or U14591 (N_14591,N_13819,N_13642);
or U14592 (N_14592,N_13508,N_13547);
and U14593 (N_14593,N_14031,N_14245);
nor U14594 (N_14594,N_13690,N_13970);
nand U14595 (N_14595,N_13692,N_13849);
nor U14596 (N_14596,N_14215,N_14181);
nor U14597 (N_14597,N_14106,N_13552);
nor U14598 (N_14598,N_14056,N_13629);
or U14599 (N_14599,N_14157,N_13689);
nor U14600 (N_14600,N_13773,N_14114);
nand U14601 (N_14601,N_13627,N_13535);
nor U14602 (N_14602,N_14208,N_13668);
or U14603 (N_14603,N_13597,N_13917);
or U14604 (N_14604,N_14218,N_14119);
nand U14605 (N_14605,N_13988,N_13714);
nor U14606 (N_14606,N_13854,N_14196);
or U14607 (N_14607,N_13613,N_14160);
and U14608 (N_14608,N_13853,N_13765);
and U14609 (N_14609,N_14246,N_14115);
or U14610 (N_14610,N_13656,N_13569);
nor U14611 (N_14611,N_14224,N_13665);
and U14612 (N_14612,N_13999,N_13903);
and U14613 (N_14613,N_13685,N_13555);
and U14614 (N_14614,N_14223,N_14153);
or U14615 (N_14615,N_13776,N_13797);
or U14616 (N_14616,N_13949,N_13811);
nor U14617 (N_14617,N_13786,N_14168);
nand U14618 (N_14618,N_14233,N_13731);
and U14619 (N_14619,N_13906,N_13865);
nor U14620 (N_14620,N_13612,N_13967);
nor U14621 (N_14621,N_13880,N_13884);
nand U14622 (N_14622,N_14095,N_13503);
and U14623 (N_14623,N_13619,N_14152);
nand U14624 (N_14624,N_14010,N_13709);
xor U14625 (N_14625,N_13608,N_13960);
nor U14626 (N_14626,N_13544,N_14053);
nor U14627 (N_14627,N_13776,N_13628);
or U14628 (N_14628,N_13855,N_13644);
and U14629 (N_14629,N_13728,N_14220);
nor U14630 (N_14630,N_13918,N_14188);
and U14631 (N_14631,N_14150,N_13558);
nor U14632 (N_14632,N_13709,N_13608);
and U14633 (N_14633,N_13974,N_13689);
and U14634 (N_14634,N_14127,N_14080);
and U14635 (N_14635,N_14093,N_13955);
and U14636 (N_14636,N_14015,N_14078);
and U14637 (N_14637,N_14152,N_13946);
and U14638 (N_14638,N_14153,N_13736);
nor U14639 (N_14639,N_14016,N_14160);
nand U14640 (N_14640,N_14232,N_13771);
and U14641 (N_14641,N_14023,N_14232);
and U14642 (N_14642,N_13543,N_13685);
and U14643 (N_14643,N_14098,N_13974);
or U14644 (N_14644,N_14019,N_14154);
or U14645 (N_14645,N_14038,N_13840);
nor U14646 (N_14646,N_13628,N_13663);
and U14647 (N_14647,N_13888,N_13637);
and U14648 (N_14648,N_14144,N_14143);
nand U14649 (N_14649,N_13786,N_13689);
or U14650 (N_14650,N_13719,N_14065);
nand U14651 (N_14651,N_13550,N_13625);
nand U14652 (N_14652,N_13942,N_13512);
or U14653 (N_14653,N_13897,N_14056);
or U14654 (N_14654,N_13759,N_14093);
or U14655 (N_14655,N_13992,N_13969);
and U14656 (N_14656,N_14061,N_13587);
nor U14657 (N_14657,N_13543,N_14020);
nand U14658 (N_14658,N_13715,N_13930);
or U14659 (N_14659,N_13611,N_13744);
and U14660 (N_14660,N_14159,N_13915);
and U14661 (N_14661,N_14216,N_13633);
and U14662 (N_14662,N_14016,N_13562);
nand U14663 (N_14663,N_13679,N_14227);
or U14664 (N_14664,N_14152,N_13620);
or U14665 (N_14665,N_13883,N_13870);
nor U14666 (N_14666,N_13699,N_13924);
nand U14667 (N_14667,N_14108,N_13569);
xor U14668 (N_14668,N_13986,N_13857);
xor U14669 (N_14669,N_14210,N_13519);
nand U14670 (N_14670,N_13746,N_14184);
and U14671 (N_14671,N_13788,N_13578);
nand U14672 (N_14672,N_13509,N_14017);
and U14673 (N_14673,N_14096,N_14234);
nor U14674 (N_14674,N_13966,N_13974);
nor U14675 (N_14675,N_14213,N_13576);
nand U14676 (N_14676,N_14163,N_13781);
xor U14677 (N_14677,N_14219,N_13674);
nand U14678 (N_14678,N_14097,N_13919);
and U14679 (N_14679,N_13616,N_13903);
nor U14680 (N_14680,N_13986,N_13649);
nand U14681 (N_14681,N_14055,N_13689);
or U14682 (N_14682,N_13636,N_13600);
nand U14683 (N_14683,N_13983,N_13742);
or U14684 (N_14684,N_14180,N_13576);
nand U14685 (N_14685,N_14101,N_13677);
nand U14686 (N_14686,N_13635,N_13576);
and U14687 (N_14687,N_13796,N_13912);
nand U14688 (N_14688,N_13742,N_14016);
or U14689 (N_14689,N_13662,N_13547);
xor U14690 (N_14690,N_13858,N_13659);
and U14691 (N_14691,N_13741,N_13928);
and U14692 (N_14692,N_13836,N_13763);
xor U14693 (N_14693,N_13976,N_14137);
and U14694 (N_14694,N_13819,N_14208);
nor U14695 (N_14695,N_13710,N_13755);
or U14696 (N_14696,N_13995,N_13693);
nand U14697 (N_14697,N_14210,N_14113);
nor U14698 (N_14698,N_14022,N_13728);
and U14699 (N_14699,N_13970,N_13918);
nand U14700 (N_14700,N_13985,N_14233);
or U14701 (N_14701,N_14171,N_14178);
and U14702 (N_14702,N_14245,N_14236);
nor U14703 (N_14703,N_14056,N_14213);
xnor U14704 (N_14704,N_13755,N_13716);
or U14705 (N_14705,N_13632,N_14229);
nand U14706 (N_14706,N_13808,N_14007);
nand U14707 (N_14707,N_13898,N_14025);
and U14708 (N_14708,N_14084,N_13967);
and U14709 (N_14709,N_13707,N_13720);
nand U14710 (N_14710,N_14079,N_13783);
nor U14711 (N_14711,N_13701,N_13876);
nand U14712 (N_14712,N_13655,N_14218);
or U14713 (N_14713,N_13648,N_13560);
or U14714 (N_14714,N_14238,N_13916);
or U14715 (N_14715,N_13641,N_14213);
or U14716 (N_14716,N_14100,N_13994);
and U14717 (N_14717,N_14174,N_14010);
and U14718 (N_14718,N_13882,N_13743);
and U14719 (N_14719,N_14188,N_14233);
xor U14720 (N_14720,N_13515,N_13941);
and U14721 (N_14721,N_13717,N_14200);
and U14722 (N_14722,N_13641,N_13535);
nor U14723 (N_14723,N_14145,N_13780);
nor U14724 (N_14724,N_13704,N_14165);
or U14725 (N_14725,N_13629,N_13633);
nand U14726 (N_14726,N_13538,N_13974);
nor U14727 (N_14727,N_14103,N_14246);
nor U14728 (N_14728,N_13566,N_13798);
or U14729 (N_14729,N_13955,N_14007);
nand U14730 (N_14730,N_14153,N_13690);
and U14731 (N_14731,N_13789,N_14222);
or U14732 (N_14732,N_13998,N_13710);
and U14733 (N_14733,N_13943,N_13947);
xnor U14734 (N_14734,N_13520,N_13653);
nand U14735 (N_14735,N_13519,N_13990);
and U14736 (N_14736,N_13665,N_13979);
and U14737 (N_14737,N_13792,N_13893);
or U14738 (N_14738,N_13764,N_13863);
xor U14739 (N_14739,N_13593,N_13911);
or U14740 (N_14740,N_14005,N_13578);
or U14741 (N_14741,N_14032,N_13927);
or U14742 (N_14742,N_13659,N_13731);
or U14743 (N_14743,N_14068,N_13732);
or U14744 (N_14744,N_13674,N_13596);
or U14745 (N_14745,N_14022,N_14123);
nand U14746 (N_14746,N_13678,N_14104);
or U14747 (N_14747,N_13640,N_13970);
or U14748 (N_14748,N_13571,N_14243);
nor U14749 (N_14749,N_13545,N_13979);
and U14750 (N_14750,N_13554,N_14052);
and U14751 (N_14751,N_13760,N_14081);
nor U14752 (N_14752,N_14061,N_13595);
and U14753 (N_14753,N_14011,N_13501);
nor U14754 (N_14754,N_13561,N_13758);
nand U14755 (N_14755,N_14237,N_14078);
nand U14756 (N_14756,N_14024,N_13813);
or U14757 (N_14757,N_13710,N_14233);
nor U14758 (N_14758,N_13800,N_14019);
nor U14759 (N_14759,N_13791,N_13784);
nand U14760 (N_14760,N_14106,N_14212);
or U14761 (N_14761,N_14233,N_13979);
nor U14762 (N_14762,N_13707,N_14119);
or U14763 (N_14763,N_13782,N_14201);
nor U14764 (N_14764,N_13623,N_13886);
and U14765 (N_14765,N_14137,N_14204);
xnor U14766 (N_14766,N_13876,N_13619);
nand U14767 (N_14767,N_13572,N_13813);
nor U14768 (N_14768,N_13534,N_13802);
or U14769 (N_14769,N_14243,N_14067);
nor U14770 (N_14770,N_14110,N_13672);
nand U14771 (N_14771,N_14070,N_14038);
or U14772 (N_14772,N_13503,N_13649);
or U14773 (N_14773,N_13754,N_14095);
or U14774 (N_14774,N_13943,N_14100);
nand U14775 (N_14775,N_13500,N_13783);
and U14776 (N_14776,N_13801,N_14188);
xor U14777 (N_14777,N_14154,N_13818);
and U14778 (N_14778,N_13946,N_13945);
or U14779 (N_14779,N_14062,N_13654);
or U14780 (N_14780,N_13806,N_13832);
or U14781 (N_14781,N_13815,N_13579);
xnor U14782 (N_14782,N_13758,N_13603);
nor U14783 (N_14783,N_13776,N_14209);
nor U14784 (N_14784,N_13598,N_13789);
xnor U14785 (N_14785,N_14091,N_14080);
and U14786 (N_14786,N_14205,N_14219);
nor U14787 (N_14787,N_13851,N_13741);
nor U14788 (N_14788,N_13589,N_13615);
or U14789 (N_14789,N_13979,N_13736);
or U14790 (N_14790,N_13671,N_14170);
nor U14791 (N_14791,N_13809,N_13882);
or U14792 (N_14792,N_14017,N_14092);
or U14793 (N_14793,N_13665,N_13945);
nor U14794 (N_14794,N_14093,N_13760);
or U14795 (N_14795,N_13658,N_13970);
or U14796 (N_14796,N_13698,N_14145);
and U14797 (N_14797,N_13621,N_13672);
nor U14798 (N_14798,N_13581,N_14229);
xor U14799 (N_14799,N_14233,N_13653);
nand U14800 (N_14800,N_14228,N_14093);
or U14801 (N_14801,N_13642,N_13871);
nor U14802 (N_14802,N_14248,N_13742);
or U14803 (N_14803,N_14008,N_13893);
and U14804 (N_14804,N_13626,N_13718);
or U14805 (N_14805,N_13593,N_13638);
or U14806 (N_14806,N_14040,N_14221);
xnor U14807 (N_14807,N_13762,N_13509);
or U14808 (N_14808,N_13613,N_13691);
nor U14809 (N_14809,N_13912,N_13688);
nand U14810 (N_14810,N_13528,N_13843);
nor U14811 (N_14811,N_13523,N_14229);
nand U14812 (N_14812,N_13630,N_14231);
and U14813 (N_14813,N_13680,N_13513);
and U14814 (N_14814,N_14112,N_13825);
and U14815 (N_14815,N_14131,N_13720);
nand U14816 (N_14816,N_13742,N_13502);
nor U14817 (N_14817,N_13906,N_13587);
nor U14818 (N_14818,N_13635,N_13933);
and U14819 (N_14819,N_14170,N_14188);
and U14820 (N_14820,N_13722,N_13602);
or U14821 (N_14821,N_13808,N_13686);
or U14822 (N_14822,N_13510,N_13769);
and U14823 (N_14823,N_13527,N_14055);
xor U14824 (N_14824,N_13674,N_13551);
nand U14825 (N_14825,N_13815,N_13626);
nor U14826 (N_14826,N_13692,N_13818);
nand U14827 (N_14827,N_14173,N_14063);
xnor U14828 (N_14828,N_13677,N_14060);
and U14829 (N_14829,N_13718,N_13926);
or U14830 (N_14830,N_14166,N_14217);
xor U14831 (N_14831,N_13803,N_14205);
nor U14832 (N_14832,N_13743,N_13787);
and U14833 (N_14833,N_13914,N_14007);
or U14834 (N_14834,N_14044,N_13889);
or U14835 (N_14835,N_13976,N_14183);
and U14836 (N_14836,N_13928,N_13996);
xnor U14837 (N_14837,N_13587,N_14220);
nand U14838 (N_14838,N_13872,N_13775);
nand U14839 (N_14839,N_13586,N_13725);
or U14840 (N_14840,N_14008,N_14153);
or U14841 (N_14841,N_13636,N_13747);
and U14842 (N_14842,N_13731,N_14104);
nand U14843 (N_14843,N_14044,N_13571);
nor U14844 (N_14844,N_13901,N_13595);
nor U14845 (N_14845,N_14050,N_14162);
xor U14846 (N_14846,N_14104,N_14241);
nand U14847 (N_14847,N_14177,N_13900);
and U14848 (N_14848,N_13785,N_14142);
and U14849 (N_14849,N_13795,N_13999);
and U14850 (N_14850,N_13670,N_13951);
or U14851 (N_14851,N_13952,N_13659);
and U14852 (N_14852,N_14096,N_13767);
and U14853 (N_14853,N_13819,N_13633);
nor U14854 (N_14854,N_13772,N_14173);
and U14855 (N_14855,N_13713,N_13892);
xor U14856 (N_14856,N_13521,N_13965);
nand U14857 (N_14857,N_13688,N_14077);
nand U14858 (N_14858,N_13977,N_13793);
nor U14859 (N_14859,N_13524,N_13900);
and U14860 (N_14860,N_13822,N_13546);
nor U14861 (N_14861,N_13627,N_14197);
nor U14862 (N_14862,N_13852,N_14060);
xnor U14863 (N_14863,N_13978,N_13586);
nor U14864 (N_14864,N_13871,N_13900);
nor U14865 (N_14865,N_13992,N_13621);
or U14866 (N_14866,N_13867,N_13740);
nor U14867 (N_14867,N_14248,N_13754);
nor U14868 (N_14868,N_13547,N_13613);
nand U14869 (N_14869,N_14149,N_13780);
nand U14870 (N_14870,N_13973,N_14139);
or U14871 (N_14871,N_14034,N_13511);
nand U14872 (N_14872,N_13695,N_13919);
and U14873 (N_14873,N_14188,N_13854);
or U14874 (N_14874,N_13615,N_13611);
or U14875 (N_14875,N_13575,N_13865);
or U14876 (N_14876,N_13624,N_14020);
nand U14877 (N_14877,N_14112,N_13501);
xor U14878 (N_14878,N_14171,N_14109);
nand U14879 (N_14879,N_13579,N_13847);
or U14880 (N_14880,N_13923,N_13644);
or U14881 (N_14881,N_13860,N_13693);
or U14882 (N_14882,N_13883,N_13726);
xor U14883 (N_14883,N_13633,N_14118);
nand U14884 (N_14884,N_14170,N_14151);
nor U14885 (N_14885,N_13614,N_13931);
or U14886 (N_14886,N_13887,N_13993);
and U14887 (N_14887,N_13849,N_13937);
nor U14888 (N_14888,N_13714,N_13523);
xor U14889 (N_14889,N_13988,N_13670);
nor U14890 (N_14890,N_13856,N_13786);
nand U14891 (N_14891,N_13777,N_13744);
nand U14892 (N_14892,N_14172,N_13618);
nor U14893 (N_14893,N_13787,N_14212);
or U14894 (N_14894,N_13626,N_13907);
and U14895 (N_14895,N_13523,N_13911);
and U14896 (N_14896,N_14137,N_13584);
nand U14897 (N_14897,N_13903,N_13740);
or U14898 (N_14898,N_13705,N_14166);
and U14899 (N_14899,N_14031,N_13813);
nor U14900 (N_14900,N_13738,N_13683);
nor U14901 (N_14901,N_13822,N_13800);
nand U14902 (N_14902,N_13722,N_13564);
nand U14903 (N_14903,N_14064,N_14084);
nand U14904 (N_14904,N_14244,N_14010);
nor U14905 (N_14905,N_13971,N_14171);
and U14906 (N_14906,N_13580,N_13900);
nand U14907 (N_14907,N_13879,N_13635);
and U14908 (N_14908,N_13645,N_13548);
xnor U14909 (N_14909,N_13708,N_13572);
nor U14910 (N_14910,N_13656,N_13878);
nand U14911 (N_14911,N_13825,N_13975);
or U14912 (N_14912,N_14177,N_13608);
xor U14913 (N_14913,N_13899,N_14168);
nor U14914 (N_14914,N_13816,N_13588);
nand U14915 (N_14915,N_13986,N_14203);
xor U14916 (N_14916,N_14172,N_13982);
xnor U14917 (N_14917,N_14070,N_14051);
nand U14918 (N_14918,N_13700,N_13652);
and U14919 (N_14919,N_13633,N_14175);
nor U14920 (N_14920,N_14128,N_13835);
and U14921 (N_14921,N_14215,N_13570);
and U14922 (N_14922,N_14178,N_14067);
and U14923 (N_14923,N_13936,N_13757);
or U14924 (N_14924,N_14227,N_13838);
xor U14925 (N_14925,N_13753,N_13665);
nand U14926 (N_14926,N_14224,N_13977);
and U14927 (N_14927,N_13765,N_13538);
or U14928 (N_14928,N_13883,N_13917);
nor U14929 (N_14929,N_13666,N_14019);
nand U14930 (N_14930,N_14070,N_13994);
nand U14931 (N_14931,N_13890,N_14135);
or U14932 (N_14932,N_13794,N_13651);
xor U14933 (N_14933,N_14133,N_13915);
nor U14934 (N_14934,N_14189,N_14062);
nand U14935 (N_14935,N_13903,N_14208);
nor U14936 (N_14936,N_14202,N_14234);
and U14937 (N_14937,N_13927,N_13522);
and U14938 (N_14938,N_13715,N_13867);
and U14939 (N_14939,N_13980,N_14021);
xor U14940 (N_14940,N_13991,N_14091);
nand U14941 (N_14941,N_13566,N_13565);
nand U14942 (N_14942,N_13750,N_13526);
or U14943 (N_14943,N_14217,N_14121);
nor U14944 (N_14944,N_14013,N_14168);
or U14945 (N_14945,N_14190,N_13619);
xor U14946 (N_14946,N_14118,N_14034);
nor U14947 (N_14947,N_14027,N_14098);
nor U14948 (N_14948,N_14037,N_13982);
or U14949 (N_14949,N_14109,N_13907);
and U14950 (N_14950,N_13675,N_14201);
nand U14951 (N_14951,N_13830,N_13758);
nand U14952 (N_14952,N_13925,N_13524);
or U14953 (N_14953,N_13591,N_14166);
and U14954 (N_14954,N_14029,N_14076);
and U14955 (N_14955,N_14003,N_14180);
or U14956 (N_14956,N_13817,N_14178);
and U14957 (N_14957,N_14118,N_13808);
or U14958 (N_14958,N_14180,N_13900);
nand U14959 (N_14959,N_14187,N_14100);
nor U14960 (N_14960,N_13637,N_13629);
and U14961 (N_14961,N_13725,N_13758);
and U14962 (N_14962,N_13875,N_13651);
and U14963 (N_14963,N_13671,N_14049);
and U14964 (N_14964,N_13510,N_14204);
nor U14965 (N_14965,N_14204,N_14044);
or U14966 (N_14966,N_13691,N_13579);
xnor U14967 (N_14967,N_13528,N_13891);
nor U14968 (N_14968,N_14224,N_13511);
or U14969 (N_14969,N_13655,N_13716);
nand U14970 (N_14970,N_13666,N_13597);
nand U14971 (N_14971,N_14185,N_13962);
and U14972 (N_14972,N_13798,N_14084);
nor U14973 (N_14973,N_13526,N_14073);
xnor U14974 (N_14974,N_13876,N_13520);
nand U14975 (N_14975,N_13812,N_14028);
and U14976 (N_14976,N_13526,N_13822);
nand U14977 (N_14977,N_14068,N_13938);
nor U14978 (N_14978,N_14046,N_14007);
or U14979 (N_14979,N_14093,N_13752);
xnor U14980 (N_14980,N_13697,N_13989);
nor U14981 (N_14981,N_13668,N_13835);
or U14982 (N_14982,N_13892,N_13640);
and U14983 (N_14983,N_13849,N_13935);
and U14984 (N_14984,N_13678,N_13525);
nor U14985 (N_14985,N_13681,N_14220);
and U14986 (N_14986,N_14009,N_13588);
xnor U14987 (N_14987,N_13749,N_14219);
xnor U14988 (N_14988,N_13580,N_13520);
and U14989 (N_14989,N_13757,N_13599);
nor U14990 (N_14990,N_13901,N_13984);
xor U14991 (N_14991,N_13741,N_13632);
or U14992 (N_14992,N_13747,N_14062);
and U14993 (N_14993,N_13584,N_13693);
or U14994 (N_14994,N_14183,N_13686);
nor U14995 (N_14995,N_14088,N_13985);
nor U14996 (N_14996,N_14148,N_13627);
nand U14997 (N_14997,N_13631,N_13721);
xnor U14998 (N_14998,N_14191,N_13554);
and U14999 (N_14999,N_13552,N_13511);
nor UO_0 (O_0,N_14691,N_14574);
and UO_1 (O_1,N_14257,N_14467);
or UO_2 (O_2,N_14264,N_14939);
nand UO_3 (O_3,N_14267,N_14306);
and UO_4 (O_4,N_14361,N_14923);
xor UO_5 (O_5,N_14671,N_14646);
xnor UO_6 (O_6,N_14366,N_14878);
xor UO_7 (O_7,N_14664,N_14269);
and UO_8 (O_8,N_14511,N_14323);
nand UO_9 (O_9,N_14859,N_14555);
nor UO_10 (O_10,N_14358,N_14405);
or UO_11 (O_11,N_14581,N_14413);
and UO_12 (O_12,N_14732,N_14421);
or UO_13 (O_13,N_14308,N_14698);
and UO_14 (O_14,N_14778,N_14775);
nor UO_15 (O_15,N_14381,N_14596);
or UO_16 (O_16,N_14615,N_14556);
and UO_17 (O_17,N_14475,N_14702);
or UO_18 (O_18,N_14398,N_14779);
or UO_19 (O_19,N_14924,N_14410);
nand UO_20 (O_20,N_14605,N_14334);
or UO_21 (O_21,N_14625,N_14313);
nand UO_22 (O_22,N_14510,N_14521);
nand UO_23 (O_23,N_14966,N_14609);
or UO_24 (O_24,N_14647,N_14342);
nor UO_25 (O_25,N_14639,N_14838);
or UO_26 (O_26,N_14650,N_14331);
and UO_27 (O_27,N_14616,N_14975);
or UO_28 (O_28,N_14635,N_14900);
or UO_29 (O_29,N_14712,N_14478);
nand UO_30 (O_30,N_14570,N_14485);
nor UO_31 (O_31,N_14281,N_14707);
and UO_32 (O_32,N_14294,N_14551);
nand UO_33 (O_33,N_14285,N_14634);
nor UO_34 (O_34,N_14817,N_14663);
or UO_35 (O_35,N_14665,N_14651);
or UO_36 (O_36,N_14364,N_14290);
and UO_37 (O_37,N_14981,N_14872);
and UO_38 (O_38,N_14669,N_14482);
or UO_39 (O_39,N_14465,N_14350);
or UO_40 (O_40,N_14340,N_14881);
and UO_41 (O_41,N_14988,N_14329);
xor UO_42 (O_42,N_14481,N_14662);
nand UO_43 (O_43,N_14268,N_14417);
and UO_44 (O_44,N_14636,N_14642);
nand UO_45 (O_45,N_14491,N_14328);
nor UO_46 (O_46,N_14270,N_14653);
or UO_47 (O_47,N_14254,N_14289);
nand UO_48 (O_48,N_14330,N_14367);
or UO_49 (O_49,N_14470,N_14758);
nor UO_50 (O_50,N_14764,N_14456);
and UO_51 (O_51,N_14517,N_14628);
or UO_52 (O_52,N_14554,N_14565);
nor UO_53 (O_53,N_14837,N_14607);
and UO_54 (O_54,N_14363,N_14567);
xnor UO_55 (O_55,N_14278,N_14529);
or UO_56 (O_56,N_14845,N_14586);
nand UO_57 (O_57,N_14406,N_14479);
nand UO_58 (O_58,N_14487,N_14751);
and UO_59 (O_59,N_14755,N_14575);
nor UO_60 (O_60,N_14537,N_14725);
or UO_61 (O_61,N_14833,N_14718);
nand UO_62 (O_62,N_14566,N_14800);
or UO_63 (O_63,N_14549,N_14291);
or UO_64 (O_64,N_14950,N_14700);
nor UO_65 (O_65,N_14305,N_14640);
or UO_66 (O_66,N_14304,N_14885);
or UO_67 (O_67,N_14962,N_14906);
or UO_68 (O_68,N_14760,N_14969);
or UO_69 (O_69,N_14948,N_14344);
nand UO_70 (O_70,N_14433,N_14284);
and UO_71 (O_71,N_14892,N_14723);
and UO_72 (O_72,N_14250,N_14790);
or UO_73 (O_73,N_14867,N_14385);
or UO_74 (O_74,N_14714,N_14560);
xor UO_75 (O_75,N_14271,N_14438);
and UO_76 (O_76,N_14535,N_14743);
nand UO_77 (O_77,N_14747,N_14875);
nor UO_78 (O_78,N_14690,N_14538);
nand UO_79 (O_79,N_14703,N_14693);
xor UO_80 (O_80,N_14834,N_14641);
or UO_81 (O_81,N_14443,N_14498);
or UO_82 (O_82,N_14695,N_14874);
xnor UO_83 (O_83,N_14757,N_14705);
nand UO_84 (O_84,N_14637,N_14419);
nand UO_85 (O_85,N_14654,N_14766);
nand UO_86 (O_86,N_14337,N_14710);
xor UO_87 (O_87,N_14493,N_14968);
nand UO_88 (O_88,N_14624,N_14970);
nand UO_89 (O_89,N_14896,N_14709);
nor UO_90 (O_90,N_14473,N_14955);
nand UO_91 (O_91,N_14518,N_14721);
nand UO_92 (O_92,N_14391,N_14431);
and UO_93 (O_93,N_14748,N_14412);
and UO_94 (O_94,N_14287,N_14884);
or UO_95 (O_95,N_14883,N_14801);
nor UO_96 (O_96,N_14638,N_14765);
and UO_97 (O_97,N_14861,N_14595);
or UO_98 (O_98,N_14430,N_14315);
xor UO_99 (O_99,N_14610,N_14411);
nand UO_100 (O_100,N_14522,N_14440);
nand UO_101 (O_101,N_14652,N_14719);
nor UO_102 (O_102,N_14426,N_14908);
xor UO_103 (O_103,N_14986,N_14809);
and UO_104 (O_104,N_14375,N_14684);
xor UO_105 (O_105,N_14828,N_14857);
and UO_106 (O_106,N_14869,N_14463);
nor UO_107 (O_107,N_14572,N_14374);
and UO_108 (O_108,N_14820,N_14953);
and UO_109 (O_109,N_14614,N_14873);
nand UO_110 (O_110,N_14339,N_14409);
xnor UO_111 (O_111,N_14677,N_14795);
and UO_112 (O_112,N_14461,N_14840);
nor UO_113 (O_113,N_14357,N_14952);
nor UO_114 (O_114,N_14414,N_14489);
or UO_115 (O_115,N_14797,N_14643);
and UO_116 (O_116,N_14667,N_14882);
or UO_117 (O_117,N_14928,N_14998);
and UO_118 (O_118,N_14633,N_14437);
xor UO_119 (O_119,N_14830,N_14544);
xor UO_120 (O_120,N_14697,N_14769);
xor UO_121 (O_121,N_14320,N_14804);
nand UO_122 (O_122,N_14852,N_14546);
and UO_123 (O_123,N_14648,N_14490);
nor UO_124 (O_124,N_14961,N_14965);
and UO_125 (O_125,N_14984,N_14803);
and UO_126 (O_126,N_14422,N_14325);
nand UO_127 (O_127,N_14387,N_14327);
and UO_128 (O_128,N_14844,N_14656);
or UO_129 (O_129,N_14347,N_14940);
nor UO_130 (O_130,N_14392,N_14571);
and UO_131 (O_131,N_14750,N_14548);
and UO_132 (O_132,N_14523,N_14659);
nand UO_133 (O_133,N_14584,N_14951);
nand UO_134 (O_134,N_14356,N_14746);
nand UO_135 (O_135,N_14369,N_14477);
or UO_136 (O_136,N_14696,N_14520);
nor UO_137 (O_137,N_14827,N_14310);
nor UO_138 (O_138,N_14321,N_14362);
or UO_139 (O_139,N_14726,N_14887);
or UO_140 (O_140,N_14831,N_14853);
or UO_141 (O_141,N_14474,N_14503);
nor UO_142 (O_142,N_14780,N_14938);
or UO_143 (O_143,N_14326,N_14858);
nand UO_144 (O_144,N_14441,N_14259);
nand UO_145 (O_145,N_14569,N_14558);
or UO_146 (O_146,N_14811,N_14927);
or UO_147 (O_147,N_14810,N_14683);
nor UO_148 (O_148,N_14488,N_14850);
and UO_149 (O_149,N_14871,N_14865);
xnor UO_150 (O_150,N_14386,N_14279);
or UO_151 (O_151,N_14911,N_14979);
xnor UO_152 (O_152,N_14715,N_14793);
nor UO_153 (O_153,N_14516,N_14274);
nand UO_154 (O_154,N_14457,N_14423);
nand UO_155 (O_155,N_14262,N_14734);
and UO_156 (O_156,N_14397,N_14316);
and UO_157 (O_157,N_14371,N_14848);
nand UO_158 (O_158,N_14588,N_14622);
nand UO_159 (O_159,N_14785,N_14377);
or UO_160 (O_160,N_14782,N_14949);
nand UO_161 (O_161,N_14352,N_14260);
and UO_162 (O_162,N_14727,N_14956);
nand UO_163 (O_163,N_14436,N_14762);
and UO_164 (O_164,N_14519,N_14672);
and UO_165 (O_165,N_14711,N_14805);
xor UO_166 (O_166,N_14842,N_14349);
and UO_167 (O_167,N_14909,N_14505);
xnor UO_168 (O_168,N_14922,N_14752);
nand UO_169 (O_169,N_14439,N_14891);
nor UO_170 (O_170,N_14644,N_14360);
or UO_171 (O_171,N_14749,N_14370);
nor UO_172 (O_172,N_14620,N_14343);
and UO_173 (O_173,N_14318,N_14314);
and UO_174 (O_174,N_14914,N_14798);
and UO_175 (O_175,N_14252,N_14919);
nand UO_176 (O_176,N_14396,N_14826);
or UO_177 (O_177,N_14997,N_14612);
and UO_178 (O_178,N_14302,N_14445);
and UO_179 (O_179,N_14701,N_14819);
nor UO_180 (O_180,N_14545,N_14598);
or UO_181 (O_181,N_14945,N_14886);
nand UO_182 (O_182,N_14630,N_14447);
nor UO_183 (O_183,N_14288,N_14847);
nor UO_184 (O_184,N_14454,N_14812);
nor UO_185 (O_185,N_14759,N_14736);
or UO_186 (O_186,N_14686,N_14716);
and UO_187 (O_187,N_14332,N_14261);
nor UO_188 (O_188,N_14602,N_14770);
nor UO_189 (O_189,N_14685,N_14983);
and UO_190 (O_190,N_14774,N_14486);
and UO_191 (O_191,N_14855,N_14960);
nor UO_192 (O_192,N_14963,N_14720);
nand UO_193 (O_193,N_14587,N_14553);
or UO_194 (O_194,N_14263,N_14737);
and UO_195 (O_195,N_14256,N_14592);
or UO_196 (O_196,N_14296,N_14832);
nor UO_197 (O_197,N_14585,N_14996);
nand UO_198 (O_198,N_14818,N_14389);
nor UO_199 (O_199,N_14613,N_14462);
or UO_200 (O_200,N_14416,N_14300);
nor UO_201 (O_201,N_14880,N_14678);
and UO_202 (O_202,N_14864,N_14729);
nand UO_203 (O_203,N_14499,N_14687);
nand UO_204 (O_204,N_14617,N_14901);
nand UO_205 (O_205,N_14539,N_14899);
or UO_206 (O_206,N_14995,N_14799);
nor UO_207 (O_207,N_14964,N_14512);
or UO_208 (O_208,N_14925,N_14657);
nand UO_209 (O_209,N_14253,N_14841);
xnor UO_210 (O_210,N_14787,N_14735);
or UO_211 (O_211,N_14724,N_14355);
nand UO_212 (O_212,N_14480,N_14303);
nand UO_213 (O_213,N_14843,N_14335);
nor UO_214 (O_214,N_14929,N_14680);
xnor UO_215 (O_215,N_14824,N_14694);
or UO_216 (O_216,N_14599,N_14890);
or UO_217 (O_217,N_14573,N_14277);
nand UO_218 (O_218,N_14946,N_14415);
nand UO_219 (O_219,N_14492,N_14404);
nand UO_220 (O_220,N_14373,N_14301);
or UO_221 (O_221,N_14382,N_14670);
nor UO_222 (O_222,N_14333,N_14608);
or UO_223 (O_223,N_14495,N_14338);
or UO_224 (O_224,N_14676,N_14982);
or UO_225 (O_225,N_14442,N_14455);
or UO_226 (O_226,N_14806,N_14449);
nand UO_227 (O_227,N_14388,N_14689);
and UO_228 (O_228,N_14744,N_14561);
or UO_229 (O_229,N_14973,N_14295);
and UO_230 (O_230,N_14353,N_14910);
nand UO_231 (O_231,N_14784,N_14679);
and UO_232 (O_232,N_14528,N_14424);
nand UO_233 (O_233,N_14682,N_14655);
and UO_234 (O_234,N_14380,N_14920);
xor UO_235 (O_235,N_14783,N_14282);
or UO_236 (O_236,N_14731,N_14788);
nand UO_237 (O_237,N_14383,N_14856);
nor UO_238 (O_238,N_14851,N_14895);
or UO_239 (O_239,N_14452,N_14854);
and UO_240 (O_240,N_14297,N_14401);
and UO_241 (O_241,N_14513,N_14930);
nand UO_242 (O_242,N_14972,N_14876);
and UO_243 (O_243,N_14276,N_14336);
xnor UO_244 (O_244,N_14976,N_14450);
nor UO_245 (O_245,N_14307,N_14954);
and UO_246 (O_246,N_14298,N_14578);
or UO_247 (O_247,N_14822,N_14286);
nand UO_248 (O_248,N_14400,N_14540);
xnor UO_249 (O_249,N_14403,N_14435);
or UO_250 (O_250,N_14594,N_14311);
xnor UO_251 (O_251,N_14533,N_14425);
and UO_252 (O_252,N_14593,N_14802);
nand UO_253 (O_253,N_14541,N_14547);
xnor UO_254 (O_254,N_14835,N_14524);
or UO_255 (O_255,N_14789,N_14542);
nand UO_256 (O_256,N_14904,N_14597);
or UO_257 (O_257,N_14471,N_14459);
or UO_258 (O_258,N_14293,N_14591);
nand UO_259 (O_259,N_14536,N_14603);
nor UO_260 (O_260,N_14453,N_14319);
and UO_261 (O_261,N_14469,N_14777);
or UO_262 (O_262,N_14564,N_14434);
nand UO_263 (O_263,N_14730,N_14897);
and UO_264 (O_264,N_14395,N_14958);
or UO_265 (O_265,N_14590,N_14621);
nand UO_266 (O_266,N_14974,N_14912);
and UO_267 (O_267,N_14754,N_14476);
nand UO_268 (O_268,N_14589,N_14273);
and UO_269 (O_269,N_14576,N_14629);
nand UO_270 (O_270,N_14530,N_14877);
nor UO_271 (O_271,N_14866,N_14563);
or UO_272 (O_272,N_14807,N_14681);
nand UO_273 (O_273,N_14378,N_14579);
and UO_274 (O_274,N_14552,N_14879);
and UO_275 (O_275,N_14509,N_14991);
nand UO_276 (O_276,N_14265,N_14889);
xnor UO_277 (O_277,N_14913,N_14796);
nor UO_278 (O_278,N_14947,N_14816);
xor UO_279 (O_279,N_14568,N_14526);
xnor UO_280 (O_280,N_14728,N_14557);
xor UO_281 (O_281,N_14534,N_14767);
xor UO_282 (O_282,N_14688,N_14660);
and UO_283 (O_283,N_14934,N_14836);
nand UO_284 (O_284,N_14903,N_14708);
nor UO_285 (O_285,N_14483,N_14661);
and UO_286 (O_286,N_14990,N_14745);
nor UO_287 (O_287,N_14915,N_14507);
nand UO_288 (O_288,N_14781,N_14739);
xor UO_289 (O_289,N_14917,N_14418);
xor UO_290 (O_290,N_14446,N_14863);
and UO_291 (O_291,N_14532,N_14606);
nand UO_292 (O_292,N_14740,N_14829);
nand UO_293 (O_293,N_14444,N_14272);
nor UO_294 (O_294,N_14980,N_14351);
nor UO_295 (O_295,N_14959,N_14791);
nor UO_296 (O_296,N_14673,N_14813);
and UO_297 (O_297,N_14967,N_14792);
nand UO_298 (O_298,N_14645,N_14742);
or UO_299 (O_299,N_14525,N_14985);
nor UO_300 (O_300,N_14738,N_14992);
nand UO_301 (O_301,N_14905,N_14600);
nor UO_302 (O_302,N_14464,N_14408);
and UO_303 (O_303,N_14292,N_14773);
nor UO_304 (O_304,N_14429,N_14849);
xor UO_305 (O_305,N_14500,N_14384);
or UO_306 (O_306,N_14627,N_14756);
and UO_307 (O_307,N_14942,N_14428);
nand UO_308 (O_308,N_14699,N_14994);
xnor UO_309 (O_309,N_14514,N_14393);
or UO_310 (O_310,N_14825,N_14266);
or UO_311 (O_311,N_14317,N_14977);
nor UO_312 (O_312,N_14935,N_14978);
nor UO_313 (O_313,N_14504,N_14666);
nand UO_314 (O_314,N_14931,N_14580);
xnor UO_315 (O_315,N_14379,N_14376);
or UO_316 (O_316,N_14704,N_14618);
nor UO_317 (O_317,N_14280,N_14432);
nand UO_318 (O_318,N_14870,N_14823);
or UO_319 (O_319,N_14502,N_14365);
and UO_320 (O_320,N_14626,N_14506);
nor UO_321 (O_321,N_14354,N_14815);
and UO_322 (O_322,N_14771,N_14846);
and UO_323 (O_323,N_14407,N_14907);
nor UO_324 (O_324,N_14255,N_14936);
or UO_325 (O_325,N_14918,N_14898);
or UO_326 (O_326,N_14448,N_14348);
or UO_327 (O_327,N_14868,N_14839);
or UO_328 (O_328,N_14989,N_14258);
and UO_329 (O_329,N_14559,N_14427);
or UO_330 (O_330,N_14275,N_14390);
nor UO_331 (O_331,N_14706,N_14674);
or UO_332 (O_332,N_14741,N_14860);
or UO_333 (O_333,N_14794,N_14345);
or UO_334 (O_334,N_14394,N_14776);
nand UO_335 (O_335,N_14926,N_14562);
nand UO_336 (O_336,N_14916,N_14692);
or UO_337 (O_337,N_14299,N_14372);
nor UO_338 (O_338,N_14466,N_14993);
nand UO_339 (O_339,N_14468,N_14309);
or UO_340 (O_340,N_14957,N_14312);
or UO_341 (O_341,N_14717,N_14893);
nor UO_342 (O_342,N_14733,N_14619);
or UO_343 (O_343,N_14460,N_14531);
nand UO_344 (O_344,N_14341,N_14888);
nand UO_345 (O_345,N_14987,N_14577);
or UO_346 (O_346,N_14543,N_14527);
nand UO_347 (O_347,N_14251,N_14937);
nor UO_348 (O_348,N_14359,N_14402);
and UO_349 (O_349,N_14582,N_14550);
nand UO_350 (O_350,N_14768,N_14763);
or UO_351 (O_351,N_14894,N_14921);
and UO_352 (O_352,N_14649,N_14583);
and UO_353 (O_353,N_14761,N_14933);
or UO_354 (O_354,N_14722,N_14631);
nand UO_355 (O_355,N_14451,N_14971);
or UO_356 (O_356,N_14753,N_14324);
and UO_357 (O_357,N_14496,N_14472);
nor UO_358 (O_358,N_14713,N_14458);
or UO_359 (O_359,N_14944,N_14675);
or UO_360 (O_360,N_14772,N_14515);
nor UO_361 (O_361,N_14808,N_14501);
and UO_362 (O_362,N_14484,N_14658);
or UO_363 (O_363,N_14814,N_14862);
or UO_364 (O_364,N_14611,N_14346);
nor UO_365 (O_365,N_14601,N_14941);
nand UO_366 (O_366,N_14821,N_14283);
nor UO_367 (O_367,N_14943,N_14322);
nor UO_368 (O_368,N_14668,N_14902);
and UO_369 (O_369,N_14632,N_14368);
nor UO_370 (O_370,N_14623,N_14786);
xor UO_371 (O_371,N_14932,N_14497);
nor UO_372 (O_372,N_14999,N_14399);
xnor UO_373 (O_373,N_14494,N_14420);
nand UO_374 (O_374,N_14604,N_14508);
nor UO_375 (O_375,N_14917,N_14403);
or UO_376 (O_376,N_14615,N_14487);
nor UO_377 (O_377,N_14772,N_14955);
or UO_378 (O_378,N_14529,N_14833);
nor UO_379 (O_379,N_14793,N_14399);
nand UO_380 (O_380,N_14554,N_14459);
nor UO_381 (O_381,N_14390,N_14960);
and UO_382 (O_382,N_14897,N_14928);
xor UO_383 (O_383,N_14349,N_14497);
and UO_384 (O_384,N_14391,N_14258);
or UO_385 (O_385,N_14385,N_14470);
or UO_386 (O_386,N_14747,N_14660);
and UO_387 (O_387,N_14539,N_14995);
nor UO_388 (O_388,N_14343,N_14631);
nor UO_389 (O_389,N_14282,N_14723);
and UO_390 (O_390,N_14819,N_14725);
nand UO_391 (O_391,N_14369,N_14326);
or UO_392 (O_392,N_14866,N_14813);
nand UO_393 (O_393,N_14444,N_14269);
or UO_394 (O_394,N_14460,N_14944);
nor UO_395 (O_395,N_14333,N_14967);
nand UO_396 (O_396,N_14273,N_14462);
nand UO_397 (O_397,N_14491,N_14441);
or UO_398 (O_398,N_14721,N_14496);
or UO_399 (O_399,N_14424,N_14870);
xor UO_400 (O_400,N_14272,N_14381);
and UO_401 (O_401,N_14919,N_14472);
nand UO_402 (O_402,N_14503,N_14285);
or UO_403 (O_403,N_14958,N_14476);
nand UO_404 (O_404,N_14737,N_14897);
nor UO_405 (O_405,N_14968,N_14425);
and UO_406 (O_406,N_14943,N_14496);
and UO_407 (O_407,N_14262,N_14576);
nand UO_408 (O_408,N_14613,N_14918);
nand UO_409 (O_409,N_14537,N_14260);
nand UO_410 (O_410,N_14283,N_14809);
or UO_411 (O_411,N_14573,N_14810);
nor UO_412 (O_412,N_14981,N_14934);
and UO_413 (O_413,N_14940,N_14729);
nand UO_414 (O_414,N_14402,N_14680);
or UO_415 (O_415,N_14834,N_14731);
xor UO_416 (O_416,N_14708,N_14658);
or UO_417 (O_417,N_14470,N_14865);
or UO_418 (O_418,N_14544,N_14716);
nand UO_419 (O_419,N_14539,N_14776);
nor UO_420 (O_420,N_14924,N_14927);
and UO_421 (O_421,N_14360,N_14817);
nand UO_422 (O_422,N_14300,N_14687);
or UO_423 (O_423,N_14585,N_14933);
and UO_424 (O_424,N_14714,N_14554);
nand UO_425 (O_425,N_14284,N_14905);
or UO_426 (O_426,N_14688,N_14537);
nor UO_427 (O_427,N_14431,N_14345);
nand UO_428 (O_428,N_14941,N_14319);
nor UO_429 (O_429,N_14302,N_14658);
xnor UO_430 (O_430,N_14959,N_14459);
or UO_431 (O_431,N_14567,N_14547);
and UO_432 (O_432,N_14864,N_14621);
nor UO_433 (O_433,N_14538,N_14925);
nand UO_434 (O_434,N_14490,N_14543);
nor UO_435 (O_435,N_14400,N_14473);
nand UO_436 (O_436,N_14819,N_14596);
nor UO_437 (O_437,N_14422,N_14667);
or UO_438 (O_438,N_14351,N_14576);
or UO_439 (O_439,N_14360,N_14327);
or UO_440 (O_440,N_14724,N_14420);
xnor UO_441 (O_441,N_14513,N_14322);
or UO_442 (O_442,N_14869,N_14785);
or UO_443 (O_443,N_14672,N_14399);
and UO_444 (O_444,N_14724,N_14573);
xnor UO_445 (O_445,N_14874,N_14994);
nor UO_446 (O_446,N_14974,N_14624);
nor UO_447 (O_447,N_14992,N_14898);
nand UO_448 (O_448,N_14897,N_14291);
nor UO_449 (O_449,N_14690,N_14900);
nand UO_450 (O_450,N_14903,N_14250);
nor UO_451 (O_451,N_14951,N_14733);
or UO_452 (O_452,N_14917,N_14660);
nor UO_453 (O_453,N_14671,N_14882);
nand UO_454 (O_454,N_14581,N_14697);
xnor UO_455 (O_455,N_14746,N_14548);
and UO_456 (O_456,N_14278,N_14382);
and UO_457 (O_457,N_14595,N_14995);
nor UO_458 (O_458,N_14819,N_14638);
nor UO_459 (O_459,N_14372,N_14827);
xnor UO_460 (O_460,N_14757,N_14778);
nor UO_461 (O_461,N_14403,N_14787);
and UO_462 (O_462,N_14481,N_14597);
or UO_463 (O_463,N_14891,N_14343);
and UO_464 (O_464,N_14407,N_14799);
nor UO_465 (O_465,N_14471,N_14258);
or UO_466 (O_466,N_14877,N_14631);
nor UO_467 (O_467,N_14431,N_14981);
nor UO_468 (O_468,N_14437,N_14304);
or UO_469 (O_469,N_14949,N_14969);
nor UO_470 (O_470,N_14351,N_14622);
or UO_471 (O_471,N_14318,N_14870);
or UO_472 (O_472,N_14645,N_14429);
nand UO_473 (O_473,N_14444,N_14359);
or UO_474 (O_474,N_14273,N_14463);
or UO_475 (O_475,N_14871,N_14295);
xor UO_476 (O_476,N_14670,N_14496);
nand UO_477 (O_477,N_14390,N_14886);
or UO_478 (O_478,N_14381,N_14312);
xnor UO_479 (O_479,N_14921,N_14547);
and UO_480 (O_480,N_14851,N_14350);
nor UO_481 (O_481,N_14368,N_14453);
xor UO_482 (O_482,N_14614,N_14888);
and UO_483 (O_483,N_14629,N_14415);
and UO_484 (O_484,N_14808,N_14513);
xnor UO_485 (O_485,N_14606,N_14490);
and UO_486 (O_486,N_14473,N_14721);
nand UO_487 (O_487,N_14949,N_14532);
or UO_488 (O_488,N_14834,N_14646);
nand UO_489 (O_489,N_14261,N_14558);
or UO_490 (O_490,N_14373,N_14333);
and UO_491 (O_491,N_14976,N_14749);
or UO_492 (O_492,N_14691,N_14755);
and UO_493 (O_493,N_14803,N_14548);
and UO_494 (O_494,N_14608,N_14475);
nor UO_495 (O_495,N_14371,N_14805);
nand UO_496 (O_496,N_14895,N_14628);
or UO_497 (O_497,N_14400,N_14396);
nor UO_498 (O_498,N_14328,N_14842);
xor UO_499 (O_499,N_14378,N_14543);
xnor UO_500 (O_500,N_14852,N_14791);
and UO_501 (O_501,N_14390,N_14574);
and UO_502 (O_502,N_14393,N_14780);
or UO_503 (O_503,N_14312,N_14807);
nand UO_504 (O_504,N_14338,N_14745);
nor UO_505 (O_505,N_14683,N_14647);
nand UO_506 (O_506,N_14943,N_14337);
or UO_507 (O_507,N_14296,N_14561);
and UO_508 (O_508,N_14496,N_14622);
xor UO_509 (O_509,N_14266,N_14535);
or UO_510 (O_510,N_14287,N_14980);
nor UO_511 (O_511,N_14775,N_14786);
or UO_512 (O_512,N_14700,N_14252);
nor UO_513 (O_513,N_14460,N_14747);
nor UO_514 (O_514,N_14608,N_14427);
or UO_515 (O_515,N_14758,N_14444);
nor UO_516 (O_516,N_14844,N_14863);
nor UO_517 (O_517,N_14670,N_14842);
nand UO_518 (O_518,N_14902,N_14598);
nand UO_519 (O_519,N_14277,N_14497);
nor UO_520 (O_520,N_14881,N_14912);
nor UO_521 (O_521,N_14791,N_14612);
and UO_522 (O_522,N_14775,N_14696);
nand UO_523 (O_523,N_14824,N_14481);
nor UO_524 (O_524,N_14943,N_14450);
nor UO_525 (O_525,N_14361,N_14664);
and UO_526 (O_526,N_14331,N_14759);
nor UO_527 (O_527,N_14904,N_14386);
nand UO_528 (O_528,N_14318,N_14508);
or UO_529 (O_529,N_14347,N_14715);
xor UO_530 (O_530,N_14507,N_14770);
xnor UO_531 (O_531,N_14977,N_14497);
xnor UO_532 (O_532,N_14931,N_14960);
nand UO_533 (O_533,N_14531,N_14265);
nand UO_534 (O_534,N_14768,N_14817);
or UO_535 (O_535,N_14607,N_14320);
and UO_536 (O_536,N_14458,N_14552);
nand UO_537 (O_537,N_14848,N_14558);
and UO_538 (O_538,N_14685,N_14577);
or UO_539 (O_539,N_14647,N_14777);
or UO_540 (O_540,N_14984,N_14527);
nand UO_541 (O_541,N_14721,N_14911);
nor UO_542 (O_542,N_14421,N_14731);
and UO_543 (O_543,N_14828,N_14770);
and UO_544 (O_544,N_14351,N_14513);
or UO_545 (O_545,N_14327,N_14995);
or UO_546 (O_546,N_14915,N_14252);
or UO_547 (O_547,N_14317,N_14368);
xnor UO_548 (O_548,N_14357,N_14837);
nand UO_549 (O_549,N_14471,N_14769);
nor UO_550 (O_550,N_14641,N_14572);
xor UO_551 (O_551,N_14977,N_14411);
or UO_552 (O_552,N_14706,N_14891);
nand UO_553 (O_553,N_14705,N_14415);
nor UO_554 (O_554,N_14576,N_14903);
nand UO_555 (O_555,N_14869,N_14932);
xnor UO_556 (O_556,N_14770,N_14671);
nor UO_557 (O_557,N_14826,N_14362);
and UO_558 (O_558,N_14987,N_14667);
nand UO_559 (O_559,N_14821,N_14560);
and UO_560 (O_560,N_14375,N_14543);
nor UO_561 (O_561,N_14320,N_14651);
nand UO_562 (O_562,N_14497,N_14972);
or UO_563 (O_563,N_14726,N_14608);
nand UO_564 (O_564,N_14621,N_14394);
and UO_565 (O_565,N_14821,N_14475);
or UO_566 (O_566,N_14774,N_14338);
nor UO_567 (O_567,N_14367,N_14282);
nand UO_568 (O_568,N_14664,N_14535);
xor UO_569 (O_569,N_14752,N_14905);
or UO_570 (O_570,N_14903,N_14945);
nand UO_571 (O_571,N_14859,N_14809);
xor UO_572 (O_572,N_14573,N_14418);
xor UO_573 (O_573,N_14563,N_14676);
and UO_574 (O_574,N_14341,N_14946);
nand UO_575 (O_575,N_14343,N_14746);
nand UO_576 (O_576,N_14805,N_14660);
or UO_577 (O_577,N_14436,N_14855);
and UO_578 (O_578,N_14534,N_14578);
nor UO_579 (O_579,N_14483,N_14285);
nand UO_580 (O_580,N_14479,N_14666);
or UO_581 (O_581,N_14341,N_14681);
and UO_582 (O_582,N_14411,N_14904);
nand UO_583 (O_583,N_14832,N_14473);
and UO_584 (O_584,N_14816,N_14630);
and UO_585 (O_585,N_14390,N_14290);
nor UO_586 (O_586,N_14605,N_14719);
or UO_587 (O_587,N_14972,N_14638);
and UO_588 (O_588,N_14527,N_14360);
nor UO_589 (O_589,N_14377,N_14676);
nand UO_590 (O_590,N_14832,N_14701);
or UO_591 (O_591,N_14772,N_14842);
and UO_592 (O_592,N_14597,N_14404);
nand UO_593 (O_593,N_14311,N_14465);
nor UO_594 (O_594,N_14859,N_14595);
or UO_595 (O_595,N_14766,N_14358);
nor UO_596 (O_596,N_14621,N_14473);
nor UO_597 (O_597,N_14994,N_14370);
xor UO_598 (O_598,N_14854,N_14561);
nor UO_599 (O_599,N_14973,N_14946);
and UO_600 (O_600,N_14506,N_14411);
or UO_601 (O_601,N_14331,N_14344);
xnor UO_602 (O_602,N_14882,N_14799);
or UO_603 (O_603,N_14295,N_14618);
and UO_604 (O_604,N_14989,N_14845);
nor UO_605 (O_605,N_14667,N_14288);
xnor UO_606 (O_606,N_14949,N_14751);
or UO_607 (O_607,N_14613,N_14544);
nand UO_608 (O_608,N_14464,N_14558);
and UO_609 (O_609,N_14557,N_14754);
or UO_610 (O_610,N_14317,N_14625);
nor UO_611 (O_611,N_14923,N_14301);
or UO_612 (O_612,N_14821,N_14930);
nand UO_613 (O_613,N_14746,N_14434);
nand UO_614 (O_614,N_14664,N_14469);
nand UO_615 (O_615,N_14929,N_14730);
and UO_616 (O_616,N_14745,N_14524);
or UO_617 (O_617,N_14324,N_14968);
or UO_618 (O_618,N_14769,N_14259);
and UO_619 (O_619,N_14422,N_14765);
nor UO_620 (O_620,N_14704,N_14324);
xnor UO_621 (O_621,N_14976,N_14878);
and UO_622 (O_622,N_14884,N_14849);
and UO_623 (O_623,N_14555,N_14535);
nand UO_624 (O_624,N_14464,N_14719);
nand UO_625 (O_625,N_14894,N_14312);
and UO_626 (O_626,N_14895,N_14921);
nor UO_627 (O_627,N_14872,N_14947);
or UO_628 (O_628,N_14594,N_14892);
and UO_629 (O_629,N_14544,N_14767);
nand UO_630 (O_630,N_14571,N_14498);
xnor UO_631 (O_631,N_14589,N_14531);
and UO_632 (O_632,N_14843,N_14894);
nand UO_633 (O_633,N_14586,N_14334);
and UO_634 (O_634,N_14716,N_14976);
and UO_635 (O_635,N_14691,N_14951);
nor UO_636 (O_636,N_14662,N_14912);
xor UO_637 (O_637,N_14800,N_14461);
nand UO_638 (O_638,N_14308,N_14808);
and UO_639 (O_639,N_14376,N_14342);
or UO_640 (O_640,N_14467,N_14315);
nor UO_641 (O_641,N_14540,N_14896);
nor UO_642 (O_642,N_14826,N_14381);
and UO_643 (O_643,N_14570,N_14684);
and UO_644 (O_644,N_14489,N_14378);
nand UO_645 (O_645,N_14877,N_14885);
nand UO_646 (O_646,N_14662,N_14638);
xor UO_647 (O_647,N_14823,N_14542);
or UO_648 (O_648,N_14499,N_14747);
and UO_649 (O_649,N_14820,N_14735);
or UO_650 (O_650,N_14781,N_14523);
or UO_651 (O_651,N_14639,N_14276);
nor UO_652 (O_652,N_14891,N_14392);
or UO_653 (O_653,N_14361,N_14800);
nor UO_654 (O_654,N_14746,N_14891);
and UO_655 (O_655,N_14509,N_14548);
and UO_656 (O_656,N_14960,N_14531);
or UO_657 (O_657,N_14650,N_14588);
or UO_658 (O_658,N_14336,N_14930);
and UO_659 (O_659,N_14633,N_14889);
xor UO_660 (O_660,N_14949,N_14367);
xnor UO_661 (O_661,N_14379,N_14785);
and UO_662 (O_662,N_14353,N_14799);
nor UO_663 (O_663,N_14324,N_14283);
nand UO_664 (O_664,N_14425,N_14317);
nor UO_665 (O_665,N_14505,N_14916);
and UO_666 (O_666,N_14387,N_14848);
nor UO_667 (O_667,N_14805,N_14258);
xnor UO_668 (O_668,N_14279,N_14710);
nand UO_669 (O_669,N_14964,N_14686);
and UO_670 (O_670,N_14553,N_14868);
nand UO_671 (O_671,N_14563,N_14959);
or UO_672 (O_672,N_14806,N_14291);
or UO_673 (O_673,N_14832,N_14487);
nor UO_674 (O_674,N_14553,N_14637);
and UO_675 (O_675,N_14811,N_14271);
or UO_676 (O_676,N_14774,N_14547);
xor UO_677 (O_677,N_14261,N_14738);
nor UO_678 (O_678,N_14564,N_14438);
and UO_679 (O_679,N_14513,N_14717);
xor UO_680 (O_680,N_14609,N_14269);
nor UO_681 (O_681,N_14363,N_14922);
nand UO_682 (O_682,N_14891,N_14883);
nand UO_683 (O_683,N_14747,N_14613);
nor UO_684 (O_684,N_14455,N_14866);
and UO_685 (O_685,N_14429,N_14464);
nand UO_686 (O_686,N_14380,N_14739);
nor UO_687 (O_687,N_14277,N_14762);
nand UO_688 (O_688,N_14490,N_14281);
nand UO_689 (O_689,N_14452,N_14487);
nand UO_690 (O_690,N_14996,N_14300);
nor UO_691 (O_691,N_14339,N_14685);
nor UO_692 (O_692,N_14408,N_14942);
nor UO_693 (O_693,N_14830,N_14790);
nor UO_694 (O_694,N_14632,N_14944);
nor UO_695 (O_695,N_14796,N_14621);
and UO_696 (O_696,N_14562,N_14928);
nand UO_697 (O_697,N_14910,N_14253);
nor UO_698 (O_698,N_14514,N_14707);
xnor UO_699 (O_699,N_14717,N_14435);
nor UO_700 (O_700,N_14522,N_14357);
and UO_701 (O_701,N_14670,N_14666);
and UO_702 (O_702,N_14334,N_14359);
or UO_703 (O_703,N_14676,N_14465);
or UO_704 (O_704,N_14734,N_14679);
or UO_705 (O_705,N_14860,N_14560);
nand UO_706 (O_706,N_14760,N_14585);
or UO_707 (O_707,N_14371,N_14440);
nand UO_708 (O_708,N_14555,N_14528);
and UO_709 (O_709,N_14388,N_14971);
nand UO_710 (O_710,N_14632,N_14394);
nor UO_711 (O_711,N_14849,N_14796);
nand UO_712 (O_712,N_14883,N_14712);
nor UO_713 (O_713,N_14935,N_14819);
or UO_714 (O_714,N_14543,N_14452);
xnor UO_715 (O_715,N_14973,N_14427);
nand UO_716 (O_716,N_14448,N_14829);
or UO_717 (O_717,N_14619,N_14893);
nor UO_718 (O_718,N_14651,N_14353);
or UO_719 (O_719,N_14339,N_14543);
and UO_720 (O_720,N_14694,N_14991);
and UO_721 (O_721,N_14813,N_14605);
or UO_722 (O_722,N_14498,N_14513);
nor UO_723 (O_723,N_14535,N_14397);
xor UO_724 (O_724,N_14434,N_14361);
and UO_725 (O_725,N_14759,N_14447);
nand UO_726 (O_726,N_14499,N_14906);
nand UO_727 (O_727,N_14883,N_14320);
or UO_728 (O_728,N_14362,N_14967);
xor UO_729 (O_729,N_14430,N_14784);
or UO_730 (O_730,N_14494,N_14501);
and UO_731 (O_731,N_14910,N_14783);
or UO_732 (O_732,N_14973,N_14572);
or UO_733 (O_733,N_14259,N_14800);
nor UO_734 (O_734,N_14281,N_14793);
or UO_735 (O_735,N_14949,N_14395);
nand UO_736 (O_736,N_14862,N_14251);
nand UO_737 (O_737,N_14508,N_14264);
nor UO_738 (O_738,N_14437,N_14500);
or UO_739 (O_739,N_14484,N_14544);
or UO_740 (O_740,N_14769,N_14828);
or UO_741 (O_741,N_14334,N_14963);
and UO_742 (O_742,N_14537,N_14759);
nor UO_743 (O_743,N_14735,N_14549);
or UO_744 (O_744,N_14354,N_14479);
nor UO_745 (O_745,N_14539,N_14684);
and UO_746 (O_746,N_14615,N_14529);
and UO_747 (O_747,N_14914,N_14652);
and UO_748 (O_748,N_14575,N_14412);
and UO_749 (O_749,N_14873,N_14318);
nor UO_750 (O_750,N_14897,N_14949);
nor UO_751 (O_751,N_14332,N_14419);
and UO_752 (O_752,N_14669,N_14718);
nor UO_753 (O_753,N_14283,N_14764);
or UO_754 (O_754,N_14859,N_14453);
nand UO_755 (O_755,N_14276,N_14295);
nand UO_756 (O_756,N_14322,N_14471);
and UO_757 (O_757,N_14293,N_14334);
and UO_758 (O_758,N_14703,N_14923);
and UO_759 (O_759,N_14987,N_14273);
nor UO_760 (O_760,N_14948,N_14605);
or UO_761 (O_761,N_14355,N_14862);
xor UO_762 (O_762,N_14975,N_14528);
or UO_763 (O_763,N_14880,N_14926);
and UO_764 (O_764,N_14673,N_14590);
nand UO_765 (O_765,N_14683,N_14629);
nand UO_766 (O_766,N_14400,N_14947);
xor UO_767 (O_767,N_14562,N_14828);
nand UO_768 (O_768,N_14964,N_14477);
nand UO_769 (O_769,N_14644,N_14882);
or UO_770 (O_770,N_14296,N_14305);
or UO_771 (O_771,N_14301,N_14417);
nor UO_772 (O_772,N_14644,N_14797);
xnor UO_773 (O_773,N_14876,N_14444);
nor UO_774 (O_774,N_14654,N_14631);
nor UO_775 (O_775,N_14945,N_14597);
and UO_776 (O_776,N_14689,N_14989);
nor UO_777 (O_777,N_14483,N_14701);
and UO_778 (O_778,N_14547,N_14581);
or UO_779 (O_779,N_14639,N_14417);
xnor UO_780 (O_780,N_14666,N_14392);
nand UO_781 (O_781,N_14616,N_14748);
nand UO_782 (O_782,N_14546,N_14565);
nand UO_783 (O_783,N_14822,N_14550);
nor UO_784 (O_784,N_14679,N_14819);
xnor UO_785 (O_785,N_14858,N_14994);
or UO_786 (O_786,N_14749,N_14985);
nand UO_787 (O_787,N_14568,N_14663);
xnor UO_788 (O_788,N_14569,N_14714);
or UO_789 (O_789,N_14322,N_14755);
nor UO_790 (O_790,N_14420,N_14635);
or UO_791 (O_791,N_14344,N_14907);
xnor UO_792 (O_792,N_14459,N_14859);
nor UO_793 (O_793,N_14475,N_14301);
and UO_794 (O_794,N_14878,N_14490);
and UO_795 (O_795,N_14799,N_14826);
nor UO_796 (O_796,N_14557,N_14377);
nor UO_797 (O_797,N_14797,N_14748);
nor UO_798 (O_798,N_14636,N_14635);
nand UO_799 (O_799,N_14648,N_14416);
or UO_800 (O_800,N_14403,N_14369);
nor UO_801 (O_801,N_14293,N_14579);
and UO_802 (O_802,N_14411,N_14939);
nand UO_803 (O_803,N_14900,N_14775);
or UO_804 (O_804,N_14528,N_14348);
or UO_805 (O_805,N_14995,N_14581);
and UO_806 (O_806,N_14816,N_14586);
and UO_807 (O_807,N_14580,N_14330);
or UO_808 (O_808,N_14731,N_14650);
or UO_809 (O_809,N_14828,N_14861);
and UO_810 (O_810,N_14722,N_14419);
xnor UO_811 (O_811,N_14795,N_14665);
and UO_812 (O_812,N_14337,N_14348);
and UO_813 (O_813,N_14941,N_14908);
xor UO_814 (O_814,N_14900,N_14451);
nand UO_815 (O_815,N_14272,N_14940);
nand UO_816 (O_816,N_14699,N_14307);
xor UO_817 (O_817,N_14412,N_14677);
nor UO_818 (O_818,N_14788,N_14866);
nand UO_819 (O_819,N_14432,N_14264);
nor UO_820 (O_820,N_14733,N_14351);
nand UO_821 (O_821,N_14497,N_14627);
xnor UO_822 (O_822,N_14838,N_14480);
xor UO_823 (O_823,N_14623,N_14826);
nor UO_824 (O_824,N_14529,N_14736);
and UO_825 (O_825,N_14277,N_14888);
nand UO_826 (O_826,N_14923,N_14437);
nand UO_827 (O_827,N_14427,N_14442);
nor UO_828 (O_828,N_14331,N_14983);
or UO_829 (O_829,N_14400,N_14378);
xnor UO_830 (O_830,N_14625,N_14698);
or UO_831 (O_831,N_14855,N_14623);
or UO_832 (O_832,N_14498,N_14297);
nand UO_833 (O_833,N_14591,N_14678);
xor UO_834 (O_834,N_14587,N_14305);
and UO_835 (O_835,N_14612,N_14801);
nand UO_836 (O_836,N_14695,N_14691);
nor UO_837 (O_837,N_14711,N_14533);
nand UO_838 (O_838,N_14270,N_14958);
nor UO_839 (O_839,N_14976,N_14288);
or UO_840 (O_840,N_14612,N_14538);
nor UO_841 (O_841,N_14347,N_14919);
nand UO_842 (O_842,N_14910,N_14500);
nand UO_843 (O_843,N_14778,N_14482);
and UO_844 (O_844,N_14274,N_14796);
nand UO_845 (O_845,N_14855,N_14400);
and UO_846 (O_846,N_14698,N_14949);
nor UO_847 (O_847,N_14828,N_14284);
and UO_848 (O_848,N_14444,N_14833);
and UO_849 (O_849,N_14449,N_14336);
nand UO_850 (O_850,N_14826,N_14577);
nor UO_851 (O_851,N_14568,N_14520);
nor UO_852 (O_852,N_14961,N_14604);
or UO_853 (O_853,N_14572,N_14504);
or UO_854 (O_854,N_14718,N_14263);
or UO_855 (O_855,N_14639,N_14530);
nand UO_856 (O_856,N_14472,N_14958);
or UO_857 (O_857,N_14509,N_14638);
nand UO_858 (O_858,N_14290,N_14286);
or UO_859 (O_859,N_14405,N_14284);
or UO_860 (O_860,N_14632,N_14992);
and UO_861 (O_861,N_14522,N_14648);
and UO_862 (O_862,N_14895,N_14524);
xor UO_863 (O_863,N_14542,N_14486);
xnor UO_864 (O_864,N_14643,N_14591);
nand UO_865 (O_865,N_14329,N_14744);
or UO_866 (O_866,N_14847,N_14300);
or UO_867 (O_867,N_14634,N_14452);
and UO_868 (O_868,N_14371,N_14970);
nor UO_869 (O_869,N_14478,N_14675);
nand UO_870 (O_870,N_14504,N_14826);
or UO_871 (O_871,N_14469,N_14785);
nor UO_872 (O_872,N_14989,N_14494);
or UO_873 (O_873,N_14364,N_14599);
and UO_874 (O_874,N_14993,N_14999);
nand UO_875 (O_875,N_14629,N_14688);
xnor UO_876 (O_876,N_14905,N_14620);
nand UO_877 (O_877,N_14533,N_14885);
or UO_878 (O_878,N_14914,N_14409);
or UO_879 (O_879,N_14525,N_14628);
and UO_880 (O_880,N_14830,N_14496);
and UO_881 (O_881,N_14796,N_14295);
and UO_882 (O_882,N_14823,N_14282);
nand UO_883 (O_883,N_14965,N_14632);
nand UO_884 (O_884,N_14547,N_14464);
and UO_885 (O_885,N_14621,N_14711);
nor UO_886 (O_886,N_14364,N_14973);
nor UO_887 (O_887,N_14860,N_14407);
or UO_888 (O_888,N_14484,N_14472);
nand UO_889 (O_889,N_14876,N_14597);
and UO_890 (O_890,N_14457,N_14750);
nor UO_891 (O_891,N_14756,N_14551);
and UO_892 (O_892,N_14784,N_14965);
or UO_893 (O_893,N_14732,N_14273);
nor UO_894 (O_894,N_14323,N_14543);
and UO_895 (O_895,N_14307,N_14616);
xor UO_896 (O_896,N_14394,N_14995);
or UO_897 (O_897,N_14486,N_14866);
and UO_898 (O_898,N_14552,N_14307);
nor UO_899 (O_899,N_14847,N_14851);
or UO_900 (O_900,N_14300,N_14638);
xnor UO_901 (O_901,N_14977,N_14950);
nor UO_902 (O_902,N_14277,N_14676);
nand UO_903 (O_903,N_14693,N_14610);
and UO_904 (O_904,N_14476,N_14711);
nand UO_905 (O_905,N_14323,N_14546);
nand UO_906 (O_906,N_14313,N_14316);
nor UO_907 (O_907,N_14687,N_14424);
or UO_908 (O_908,N_14822,N_14424);
nand UO_909 (O_909,N_14701,N_14990);
nor UO_910 (O_910,N_14759,N_14503);
nor UO_911 (O_911,N_14654,N_14558);
or UO_912 (O_912,N_14618,N_14570);
nor UO_913 (O_913,N_14831,N_14508);
nand UO_914 (O_914,N_14687,N_14955);
nand UO_915 (O_915,N_14329,N_14818);
nand UO_916 (O_916,N_14618,N_14790);
nor UO_917 (O_917,N_14506,N_14857);
nor UO_918 (O_918,N_14823,N_14573);
and UO_919 (O_919,N_14367,N_14975);
nand UO_920 (O_920,N_14832,N_14696);
nor UO_921 (O_921,N_14440,N_14447);
nand UO_922 (O_922,N_14582,N_14459);
nor UO_923 (O_923,N_14740,N_14618);
nand UO_924 (O_924,N_14517,N_14697);
and UO_925 (O_925,N_14663,N_14517);
and UO_926 (O_926,N_14324,N_14806);
or UO_927 (O_927,N_14909,N_14422);
and UO_928 (O_928,N_14274,N_14311);
nor UO_929 (O_929,N_14738,N_14425);
or UO_930 (O_930,N_14829,N_14389);
xor UO_931 (O_931,N_14813,N_14401);
nor UO_932 (O_932,N_14608,N_14699);
nor UO_933 (O_933,N_14479,N_14932);
nor UO_934 (O_934,N_14619,N_14316);
or UO_935 (O_935,N_14981,N_14907);
xor UO_936 (O_936,N_14455,N_14796);
xor UO_937 (O_937,N_14436,N_14985);
nor UO_938 (O_938,N_14566,N_14934);
nand UO_939 (O_939,N_14940,N_14951);
nor UO_940 (O_940,N_14594,N_14536);
or UO_941 (O_941,N_14445,N_14297);
and UO_942 (O_942,N_14756,N_14978);
and UO_943 (O_943,N_14343,N_14412);
nand UO_944 (O_944,N_14718,N_14876);
and UO_945 (O_945,N_14807,N_14714);
or UO_946 (O_946,N_14685,N_14406);
xor UO_947 (O_947,N_14509,N_14255);
and UO_948 (O_948,N_14475,N_14812);
and UO_949 (O_949,N_14759,N_14886);
xnor UO_950 (O_950,N_14379,N_14473);
nand UO_951 (O_951,N_14488,N_14418);
nor UO_952 (O_952,N_14800,N_14671);
or UO_953 (O_953,N_14508,N_14348);
nor UO_954 (O_954,N_14413,N_14580);
or UO_955 (O_955,N_14425,N_14912);
nand UO_956 (O_956,N_14969,N_14620);
and UO_957 (O_957,N_14880,N_14557);
nor UO_958 (O_958,N_14503,N_14964);
and UO_959 (O_959,N_14835,N_14974);
or UO_960 (O_960,N_14512,N_14552);
and UO_961 (O_961,N_14989,N_14284);
nor UO_962 (O_962,N_14995,N_14325);
or UO_963 (O_963,N_14423,N_14396);
and UO_964 (O_964,N_14936,N_14673);
and UO_965 (O_965,N_14609,N_14616);
xor UO_966 (O_966,N_14266,N_14481);
nand UO_967 (O_967,N_14815,N_14347);
nor UO_968 (O_968,N_14631,N_14955);
or UO_969 (O_969,N_14776,N_14590);
or UO_970 (O_970,N_14848,N_14359);
and UO_971 (O_971,N_14491,N_14862);
or UO_972 (O_972,N_14983,N_14305);
nor UO_973 (O_973,N_14967,N_14923);
or UO_974 (O_974,N_14996,N_14954);
nand UO_975 (O_975,N_14572,N_14590);
nand UO_976 (O_976,N_14628,N_14631);
nor UO_977 (O_977,N_14469,N_14296);
and UO_978 (O_978,N_14621,N_14340);
nor UO_979 (O_979,N_14675,N_14858);
or UO_980 (O_980,N_14595,N_14281);
and UO_981 (O_981,N_14579,N_14835);
and UO_982 (O_982,N_14513,N_14770);
nand UO_983 (O_983,N_14855,N_14410);
nand UO_984 (O_984,N_14922,N_14799);
nand UO_985 (O_985,N_14371,N_14872);
nor UO_986 (O_986,N_14795,N_14494);
nor UO_987 (O_987,N_14838,N_14345);
or UO_988 (O_988,N_14345,N_14563);
nand UO_989 (O_989,N_14774,N_14257);
and UO_990 (O_990,N_14742,N_14607);
or UO_991 (O_991,N_14730,N_14674);
nand UO_992 (O_992,N_14761,N_14792);
or UO_993 (O_993,N_14951,N_14847);
and UO_994 (O_994,N_14723,N_14820);
or UO_995 (O_995,N_14513,N_14958);
nor UO_996 (O_996,N_14620,N_14422);
or UO_997 (O_997,N_14831,N_14445);
or UO_998 (O_998,N_14677,N_14897);
nor UO_999 (O_999,N_14426,N_14885);
nand UO_1000 (O_1000,N_14578,N_14916);
and UO_1001 (O_1001,N_14657,N_14471);
xor UO_1002 (O_1002,N_14371,N_14429);
or UO_1003 (O_1003,N_14535,N_14330);
or UO_1004 (O_1004,N_14508,N_14728);
and UO_1005 (O_1005,N_14894,N_14629);
nand UO_1006 (O_1006,N_14408,N_14964);
nand UO_1007 (O_1007,N_14837,N_14633);
nand UO_1008 (O_1008,N_14935,N_14651);
or UO_1009 (O_1009,N_14883,N_14868);
or UO_1010 (O_1010,N_14667,N_14876);
nand UO_1011 (O_1011,N_14616,N_14864);
nand UO_1012 (O_1012,N_14259,N_14422);
xor UO_1013 (O_1013,N_14875,N_14300);
or UO_1014 (O_1014,N_14293,N_14516);
xor UO_1015 (O_1015,N_14407,N_14990);
nand UO_1016 (O_1016,N_14301,N_14395);
nor UO_1017 (O_1017,N_14672,N_14572);
or UO_1018 (O_1018,N_14761,N_14868);
nor UO_1019 (O_1019,N_14616,N_14868);
nor UO_1020 (O_1020,N_14887,N_14666);
nand UO_1021 (O_1021,N_14689,N_14803);
or UO_1022 (O_1022,N_14380,N_14410);
nor UO_1023 (O_1023,N_14876,N_14514);
nand UO_1024 (O_1024,N_14286,N_14985);
nor UO_1025 (O_1025,N_14615,N_14921);
nor UO_1026 (O_1026,N_14822,N_14796);
nor UO_1027 (O_1027,N_14871,N_14337);
nor UO_1028 (O_1028,N_14414,N_14642);
nand UO_1029 (O_1029,N_14534,N_14263);
and UO_1030 (O_1030,N_14342,N_14497);
nand UO_1031 (O_1031,N_14726,N_14266);
nor UO_1032 (O_1032,N_14495,N_14898);
or UO_1033 (O_1033,N_14793,N_14354);
or UO_1034 (O_1034,N_14814,N_14454);
and UO_1035 (O_1035,N_14519,N_14662);
nor UO_1036 (O_1036,N_14608,N_14390);
xnor UO_1037 (O_1037,N_14737,N_14946);
xor UO_1038 (O_1038,N_14371,N_14281);
nand UO_1039 (O_1039,N_14269,N_14522);
nor UO_1040 (O_1040,N_14606,N_14680);
nor UO_1041 (O_1041,N_14842,N_14783);
and UO_1042 (O_1042,N_14389,N_14254);
and UO_1043 (O_1043,N_14788,N_14643);
and UO_1044 (O_1044,N_14840,N_14542);
nor UO_1045 (O_1045,N_14356,N_14928);
or UO_1046 (O_1046,N_14601,N_14420);
or UO_1047 (O_1047,N_14311,N_14914);
or UO_1048 (O_1048,N_14402,N_14656);
and UO_1049 (O_1049,N_14696,N_14641);
nand UO_1050 (O_1050,N_14734,N_14260);
nor UO_1051 (O_1051,N_14647,N_14614);
xnor UO_1052 (O_1052,N_14363,N_14643);
xor UO_1053 (O_1053,N_14382,N_14776);
nand UO_1054 (O_1054,N_14393,N_14500);
and UO_1055 (O_1055,N_14965,N_14588);
nand UO_1056 (O_1056,N_14454,N_14474);
nor UO_1057 (O_1057,N_14838,N_14809);
xor UO_1058 (O_1058,N_14923,N_14743);
or UO_1059 (O_1059,N_14999,N_14574);
nor UO_1060 (O_1060,N_14416,N_14519);
and UO_1061 (O_1061,N_14619,N_14489);
nand UO_1062 (O_1062,N_14563,N_14704);
or UO_1063 (O_1063,N_14741,N_14674);
nor UO_1064 (O_1064,N_14574,N_14689);
nor UO_1065 (O_1065,N_14485,N_14907);
nor UO_1066 (O_1066,N_14560,N_14961);
xnor UO_1067 (O_1067,N_14686,N_14273);
and UO_1068 (O_1068,N_14776,N_14644);
nor UO_1069 (O_1069,N_14971,N_14599);
nor UO_1070 (O_1070,N_14867,N_14387);
nor UO_1071 (O_1071,N_14857,N_14775);
xor UO_1072 (O_1072,N_14501,N_14476);
nand UO_1073 (O_1073,N_14651,N_14809);
nor UO_1074 (O_1074,N_14339,N_14668);
or UO_1075 (O_1075,N_14575,N_14629);
nand UO_1076 (O_1076,N_14447,N_14406);
xnor UO_1077 (O_1077,N_14438,N_14283);
and UO_1078 (O_1078,N_14470,N_14332);
and UO_1079 (O_1079,N_14659,N_14774);
nand UO_1080 (O_1080,N_14828,N_14760);
nand UO_1081 (O_1081,N_14504,N_14337);
and UO_1082 (O_1082,N_14777,N_14787);
nand UO_1083 (O_1083,N_14914,N_14799);
or UO_1084 (O_1084,N_14909,N_14973);
or UO_1085 (O_1085,N_14876,N_14303);
nand UO_1086 (O_1086,N_14402,N_14928);
nor UO_1087 (O_1087,N_14983,N_14542);
nand UO_1088 (O_1088,N_14339,N_14250);
and UO_1089 (O_1089,N_14786,N_14585);
nor UO_1090 (O_1090,N_14636,N_14501);
nand UO_1091 (O_1091,N_14553,N_14856);
nand UO_1092 (O_1092,N_14857,N_14376);
or UO_1093 (O_1093,N_14428,N_14633);
or UO_1094 (O_1094,N_14279,N_14601);
and UO_1095 (O_1095,N_14571,N_14643);
nor UO_1096 (O_1096,N_14976,N_14371);
nand UO_1097 (O_1097,N_14699,N_14374);
xnor UO_1098 (O_1098,N_14994,N_14705);
or UO_1099 (O_1099,N_14512,N_14654);
or UO_1100 (O_1100,N_14268,N_14467);
nand UO_1101 (O_1101,N_14290,N_14869);
and UO_1102 (O_1102,N_14643,N_14498);
or UO_1103 (O_1103,N_14795,N_14797);
nor UO_1104 (O_1104,N_14801,N_14793);
and UO_1105 (O_1105,N_14962,N_14326);
nand UO_1106 (O_1106,N_14375,N_14327);
nor UO_1107 (O_1107,N_14589,N_14580);
nor UO_1108 (O_1108,N_14366,N_14331);
nor UO_1109 (O_1109,N_14684,N_14389);
and UO_1110 (O_1110,N_14693,N_14593);
nor UO_1111 (O_1111,N_14437,N_14426);
or UO_1112 (O_1112,N_14424,N_14842);
or UO_1113 (O_1113,N_14622,N_14456);
nor UO_1114 (O_1114,N_14300,N_14252);
nand UO_1115 (O_1115,N_14788,N_14655);
nand UO_1116 (O_1116,N_14558,N_14723);
and UO_1117 (O_1117,N_14833,N_14346);
and UO_1118 (O_1118,N_14708,N_14674);
and UO_1119 (O_1119,N_14624,N_14278);
nor UO_1120 (O_1120,N_14252,N_14384);
and UO_1121 (O_1121,N_14883,N_14857);
nand UO_1122 (O_1122,N_14396,N_14885);
xor UO_1123 (O_1123,N_14888,N_14780);
and UO_1124 (O_1124,N_14934,N_14437);
nand UO_1125 (O_1125,N_14444,N_14389);
or UO_1126 (O_1126,N_14557,N_14820);
nand UO_1127 (O_1127,N_14462,N_14542);
nand UO_1128 (O_1128,N_14828,N_14807);
nor UO_1129 (O_1129,N_14319,N_14652);
nor UO_1130 (O_1130,N_14789,N_14832);
or UO_1131 (O_1131,N_14357,N_14727);
and UO_1132 (O_1132,N_14444,N_14319);
xnor UO_1133 (O_1133,N_14377,N_14706);
nand UO_1134 (O_1134,N_14764,N_14926);
nor UO_1135 (O_1135,N_14701,N_14271);
xnor UO_1136 (O_1136,N_14620,N_14874);
or UO_1137 (O_1137,N_14780,N_14474);
and UO_1138 (O_1138,N_14327,N_14880);
nand UO_1139 (O_1139,N_14800,N_14377);
and UO_1140 (O_1140,N_14640,N_14683);
nor UO_1141 (O_1141,N_14574,N_14566);
and UO_1142 (O_1142,N_14915,N_14686);
xnor UO_1143 (O_1143,N_14693,N_14972);
nor UO_1144 (O_1144,N_14583,N_14278);
nor UO_1145 (O_1145,N_14510,N_14789);
nor UO_1146 (O_1146,N_14600,N_14373);
and UO_1147 (O_1147,N_14812,N_14294);
nand UO_1148 (O_1148,N_14836,N_14720);
xnor UO_1149 (O_1149,N_14840,N_14442);
nand UO_1150 (O_1150,N_14690,N_14819);
and UO_1151 (O_1151,N_14917,N_14894);
or UO_1152 (O_1152,N_14539,N_14727);
nor UO_1153 (O_1153,N_14968,N_14559);
nor UO_1154 (O_1154,N_14387,N_14870);
and UO_1155 (O_1155,N_14732,N_14418);
nor UO_1156 (O_1156,N_14370,N_14906);
nand UO_1157 (O_1157,N_14587,N_14440);
nor UO_1158 (O_1158,N_14331,N_14746);
xor UO_1159 (O_1159,N_14434,N_14674);
nor UO_1160 (O_1160,N_14843,N_14360);
nor UO_1161 (O_1161,N_14341,N_14385);
or UO_1162 (O_1162,N_14983,N_14699);
nand UO_1163 (O_1163,N_14409,N_14868);
and UO_1164 (O_1164,N_14828,N_14576);
nor UO_1165 (O_1165,N_14473,N_14394);
xnor UO_1166 (O_1166,N_14795,N_14695);
or UO_1167 (O_1167,N_14922,N_14425);
and UO_1168 (O_1168,N_14997,N_14558);
and UO_1169 (O_1169,N_14404,N_14810);
nor UO_1170 (O_1170,N_14443,N_14682);
or UO_1171 (O_1171,N_14800,N_14941);
or UO_1172 (O_1172,N_14487,N_14517);
or UO_1173 (O_1173,N_14549,N_14647);
nand UO_1174 (O_1174,N_14714,N_14903);
or UO_1175 (O_1175,N_14266,N_14501);
nand UO_1176 (O_1176,N_14706,N_14945);
nand UO_1177 (O_1177,N_14833,N_14474);
and UO_1178 (O_1178,N_14503,N_14545);
and UO_1179 (O_1179,N_14512,N_14470);
or UO_1180 (O_1180,N_14535,N_14982);
nand UO_1181 (O_1181,N_14289,N_14265);
nor UO_1182 (O_1182,N_14630,N_14798);
xnor UO_1183 (O_1183,N_14309,N_14445);
or UO_1184 (O_1184,N_14537,N_14313);
nor UO_1185 (O_1185,N_14938,N_14840);
nand UO_1186 (O_1186,N_14924,N_14552);
xnor UO_1187 (O_1187,N_14765,N_14424);
nand UO_1188 (O_1188,N_14310,N_14748);
or UO_1189 (O_1189,N_14463,N_14379);
or UO_1190 (O_1190,N_14957,N_14310);
nor UO_1191 (O_1191,N_14351,N_14936);
nand UO_1192 (O_1192,N_14560,N_14918);
nand UO_1193 (O_1193,N_14712,N_14877);
nor UO_1194 (O_1194,N_14914,N_14706);
or UO_1195 (O_1195,N_14336,N_14570);
nor UO_1196 (O_1196,N_14358,N_14986);
and UO_1197 (O_1197,N_14478,N_14283);
nor UO_1198 (O_1198,N_14628,N_14600);
nor UO_1199 (O_1199,N_14864,N_14655);
nor UO_1200 (O_1200,N_14866,N_14493);
nand UO_1201 (O_1201,N_14341,N_14470);
and UO_1202 (O_1202,N_14878,N_14422);
xor UO_1203 (O_1203,N_14689,N_14785);
nor UO_1204 (O_1204,N_14953,N_14439);
nor UO_1205 (O_1205,N_14305,N_14285);
nand UO_1206 (O_1206,N_14943,N_14334);
and UO_1207 (O_1207,N_14919,N_14961);
nor UO_1208 (O_1208,N_14479,N_14279);
nand UO_1209 (O_1209,N_14355,N_14869);
and UO_1210 (O_1210,N_14912,N_14877);
or UO_1211 (O_1211,N_14472,N_14601);
or UO_1212 (O_1212,N_14964,N_14724);
and UO_1213 (O_1213,N_14261,N_14764);
or UO_1214 (O_1214,N_14490,N_14403);
xor UO_1215 (O_1215,N_14340,N_14882);
or UO_1216 (O_1216,N_14250,N_14315);
nor UO_1217 (O_1217,N_14506,N_14504);
nand UO_1218 (O_1218,N_14468,N_14517);
nor UO_1219 (O_1219,N_14374,N_14588);
nand UO_1220 (O_1220,N_14702,N_14395);
and UO_1221 (O_1221,N_14798,N_14776);
nor UO_1222 (O_1222,N_14486,N_14879);
nand UO_1223 (O_1223,N_14698,N_14674);
nor UO_1224 (O_1224,N_14811,N_14423);
or UO_1225 (O_1225,N_14884,N_14910);
xnor UO_1226 (O_1226,N_14423,N_14925);
and UO_1227 (O_1227,N_14300,N_14517);
nand UO_1228 (O_1228,N_14317,N_14623);
nand UO_1229 (O_1229,N_14859,N_14996);
and UO_1230 (O_1230,N_14858,N_14824);
nor UO_1231 (O_1231,N_14773,N_14481);
or UO_1232 (O_1232,N_14397,N_14741);
and UO_1233 (O_1233,N_14642,N_14560);
nor UO_1234 (O_1234,N_14977,N_14379);
or UO_1235 (O_1235,N_14444,N_14927);
or UO_1236 (O_1236,N_14659,N_14914);
nor UO_1237 (O_1237,N_14329,N_14442);
nand UO_1238 (O_1238,N_14352,N_14991);
and UO_1239 (O_1239,N_14618,N_14341);
or UO_1240 (O_1240,N_14529,N_14292);
xnor UO_1241 (O_1241,N_14874,N_14474);
xnor UO_1242 (O_1242,N_14534,N_14453);
and UO_1243 (O_1243,N_14276,N_14613);
nand UO_1244 (O_1244,N_14384,N_14707);
nor UO_1245 (O_1245,N_14694,N_14723);
nor UO_1246 (O_1246,N_14435,N_14466);
or UO_1247 (O_1247,N_14323,N_14530);
xor UO_1248 (O_1248,N_14376,N_14312);
xnor UO_1249 (O_1249,N_14820,N_14829);
or UO_1250 (O_1250,N_14789,N_14716);
nor UO_1251 (O_1251,N_14556,N_14667);
nor UO_1252 (O_1252,N_14277,N_14976);
or UO_1253 (O_1253,N_14935,N_14660);
nand UO_1254 (O_1254,N_14524,N_14656);
or UO_1255 (O_1255,N_14903,N_14627);
and UO_1256 (O_1256,N_14855,N_14459);
nand UO_1257 (O_1257,N_14834,N_14499);
nand UO_1258 (O_1258,N_14310,N_14558);
nor UO_1259 (O_1259,N_14824,N_14558);
and UO_1260 (O_1260,N_14653,N_14304);
nand UO_1261 (O_1261,N_14384,N_14645);
nand UO_1262 (O_1262,N_14370,N_14303);
nand UO_1263 (O_1263,N_14890,N_14624);
xor UO_1264 (O_1264,N_14675,N_14591);
and UO_1265 (O_1265,N_14501,N_14387);
and UO_1266 (O_1266,N_14346,N_14416);
and UO_1267 (O_1267,N_14355,N_14286);
or UO_1268 (O_1268,N_14295,N_14798);
and UO_1269 (O_1269,N_14319,N_14289);
nor UO_1270 (O_1270,N_14367,N_14301);
nand UO_1271 (O_1271,N_14921,N_14643);
nor UO_1272 (O_1272,N_14752,N_14794);
nand UO_1273 (O_1273,N_14328,N_14998);
xnor UO_1274 (O_1274,N_14845,N_14275);
or UO_1275 (O_1275,N_14529,N_14365);
and UO_1276 (O_1276,N_14998,N_14779);
xnor UO_1277 (O_1277,N_14274,N_14529);
and UO_1278 (O_1278,N_14787,N_14957);
nand UO_1279 (O_1279,N_14368,N_14308);
nor UO_1280 (O_1280,N_14438,N_14897);
nor UO_1281 (O_1281,N_14291,N_14315);
and UO_1282 (O_1282,N_14277,N_14884);
or UO_1283 (O_1283,N_14757,N_14433);
and UO_1284 (O_1284,N_14487,N_14930);
and UO_1285 (O_1285,N_14934,N_14371);
xnor UO_1286 (O_1286,N_14469,N_14894);
or UO_1287 (O_1287,N_14320,N_14816);
nor UO_1288 (O_1288,N_14987,N_14715);
nor UO_1289 (O_1289,N_14829,N_14714);
and UO_1290 (O_1290,N_14703,N_14804);
and UO_1291 (O_1291,N_14706,N_14957);
nor UO_1292 (O_1292,N_14304,N_14810);
nor UO_1293 (O_1293,N_14504,N_14544);
xnor UO_1294 (O_1294,N_14733,N_14722);
or UO_1295 (O_1295,N_14318,N_14274);
nor UO_1296 (O_1296,N_14581,N_14362);
and UO_1297 (O_1297,N_14629,N_14382);
and UO_1298 (O_1298,N_14698,N_14555);
or UO_1299 (O_1299,N_14537,N_14338);
xnor UO_1300 (O_1300,N_14691,N_14702);
xor UO_1301 (O_1301,N_14889,N_14922);
nand UO_1302 (O_1302,N_14792,N_14294);
or UO_1303 (O_1303,N_14862,N_14424);
nand UO_1304 (O_1304,N_14356,N_14579);
or UO_1305 (O_1305,N_14791,N_14790);
nand UO_1306 (O_1306,N_14603,N_14972);
and UO_1307 (O_1307,N_14656,N_14676);
xor UO_1308 (O_1308,N_14914,N_14406);
nand UO_1309 (O_1309,N_14765,N_14561);
nor UO_1310 (O_1310,N_14571,N_14402);
or UO_1311 (O_1311,N_14800,N_14691);
and UO_1312 (O_1312,N_14424,N_14864);
or UO_1313 (O_1313,N_14374,N_14635);
nand UO_1314 (O_1314,N_14600,N_14775);
or UO_1315 (O_1315,N_14356,N_14775);
or UO_1316 (O_1316,N_14545,N_14790);
nand UO_1317 (O_1317,N_14501,N_14367);
or UO_1318 (O_1318,N_14351,N_14440);
nand UO_1319 (O_1319,N_14580,N_14451);
or UO_1320 (O_1320,N_14776,N_14277);
and UO_1321 (O_1321,N_14357,N_14970);
or UO_1322 (O_1322,N_14342,N_14833);
nor UO_1323 (O_1323,N_14275,N_14266);
and UO_1324 (O_1324,N_14656,N_14935);
and UO_1325 (O_1325,N_14904,N_14485);
or UO_1326 (O_1326,N_14398,N_14272);
xnor UO_1327 (O_1327,N_14472,N_14756);
xor UO_1328 (O_1328,N_14469,N_14967);
xor UO_1329 (O_1329,N_14965,N_14314);
and UO_1330 (O_1330,N_14305,N_14559);
and UO_1331 (O_1331,N_14568,N_14331);
or UO_1332 (O_1332,N_14472,N_14316);
nor UO_1333 (O_1333,N_14857,N_14366);
nand UO_1334 (O_1334,N_14655,N_14751);
or UO_1335 (O_1335,N_14331,N_14520);
or UO_1336 (O_1336,N_14498,N_14796);
nor UO_1337 (O_1337,N_14873,N_14867);
xnor UO_1338 (O_1338,N_14834,N_14992);
nor UO_1339 (O_1339,N_14995,N_14536);
or UO_1340 (O_1340,N_14821,N_14577);
xnor UO_1341 (O_1341,N_14297,N_14686);
or UO_1342 (O_1342,N_14490,N_14762);
nor UO_1343 (O_1343,N_14310,N_14556);
or UO_1344 (O_1344,N_14816,N_14578);
nor UO_1345 (O_1345,N_14462,N_14595);
nor UO_1346 (O_1346,N_14640,N_14485);
and UO_1347 (O_1347,N_14343,N_14795);
nand UO_1348 (O_1348,N_14910,N_14455);
or UO_1349 (O_1349,N_14769,N_14654);
xor UO_1350 (O_1350,N_14758,N_14814);
or UO_1351 (O_1351,N_14840,N_14400);
and UO_1352 (O_1352,N_14692,N_14552);
and UO_1353 (O_1353,N_14562,N_14919);
or UO_1354 (O_1354,N_14642,N_14521);
and UO_1355 (O_1355,N_14709,N_14847);
or UO_1356 (O_1356,N_14544,N_14605);
or UO_1357 (O_1357,N_14294,N_14496);
nand UO_1358 (O_1358,N_14413,N_14433);
nand UO_1359 (O_1359,N_14506,N_14963);
nor UO_1360 (O_1360,N_14752,N_14626);
xor UO_1361 (O_1361,N_14445,N_14258);
or UO_1362 (O_1362,N_14774,N_14552);
nand UO_1363 (O_1363,N_14285,N_14677);
nand UO_1364 (O_1364,N_14583,N_14745);
xor UO_1365 (O_1365,N_14395,N_14251);
and UO_1366 (O_1366,N_14564,N_14301);
or UO_1367 (O_1367,N_14778,N_14972);
nor UO_1368 (O_1368,N_14293,N_14534);
nand UO_1369 (O_1369,N_14782,N_14655);
xnor UO_1370 (O_1370,N_14394,N_14987);
or UO_1371 (O_1371,N_14524,N_14335);
xor UO_1372 (O_1372,N_14708,N_14524);
or UO_1373 (O_1373,N_14857,N_14448);
or UO_1374 (O_1374,N_14622,N_14396);
and UO_1375 (O_1375,N_14799,N_14757);
nor UO_1376 (O_1376,N_14294,N_14489);
nor UO_1377 (O_1377,N_14838,N_14716);
nor UO_1378 (O_1378,N_14528,N_14856);
nand UO_1379 (O_1379,N_14919,N_14599);
nand UO_1380 (O_1380,N_14667,N_14693);
and UO_1381 (O_1381,N_14994,N_14402);
and UO_1382 (O_1382,N_14320,N_14751);
nand UO_1383 (O_1383,N_14883,N_14678);
nor UO_1384 (O_1384,N_14562,N_14849);
xnor UO_1385 (O_1385,N_14893,N_14298);
nand UO_1386 (O_1386,N_14996,N_14755);
nor UO_1387 (O_1387,N_14677,N_14481);
and UO_1388 (O_1388,N_14959,N_14522);
nand UO_1389 (O_1389,N_14720,N_14587);
nand UO_1390 (O_1390,N_14420,N_14957);
nand UO_1391 (O_1391,N_14322,N_14835);
nor UO_1392 (O_1392,N_14664,N_14728);
nor UO_1393 (O_1393,N_14608,N_14520);
nand UO_1394 (O_1394,N_14972,N_14460);
and UO_1395 (O_1395,N_14597,N_14475);
and UO_1396 (O_1396,N_14508,N_14833);
nand UO_1397 (O_1397,N_14897,N_14736);
nand UO_1398 (O_1398,N_14252,N_14371);
or UO_1399 (O_1399,N_14265,N_14864);
nand UO_1400 (O_1400,N_14592,N_14388);
or UO_1401 (O_1401,N_14449,N_14750);
or UO_1402 (O_1402,N_14508,N_14378);
nor UO_1403 (O_1403,N_14262,N_14479);
or UO_1404 (O_1404,N_14644,N_14902);
and UO_1405 (O_1405,N_14652,N_14904);
xor UO_1406 (O_1406,N_14272,N_14846);
and UO_1407 (O_1407,N_14315,N_14670);
nor UO_1408 (O_1408,N_14909,N_14512);
and UO_1409 (O_1409,N_14982,N_14482);
nand UO_1410 (O_1410,N_14963,N_14590);
and UO_1411 (O_1411,N_14547,N_14721);
or UO_1412 (O_1412,N_14438,N_14972);
or UO_1413 (O_1413,N_14321,N_14370);
nor UO_1414 (O_1414,N_14740,N_14346);
nand UO_1415 (O_1415,N_14700,N_14387);
nor UO_1416 (O_1416,N_14848,N_14461);
nor UO_1417 (O_1417,N_14345,N_14472);
nand UO_1418 (O_1418,N_14265,N_14312);
and UO_1419 (O_1419,N_14969,N_14296);
nor UO_1420 (O_1420,N_14507,N_14700);
or UO_1421 (O_1421,N_14462,N_14523);
nand UO_1422 (O_1422,N_14843,N_14979);
xor UO_1423 (O_1423,N_14513,N_14367);
xor UO_1424 (O_1424,N_14973,N_14493);
nor UO_1425 (O_1425,N_14945,N_14648);
xnor UO_1426 (O_1426,N_14908,N_14611);
nor UO_1427 (O_1427,N_14837,N_14639);
nor UO_1428 (O_1428,N_14982,N_14979);
or UO_1429 (O_1429,N_14753,N_14804);
and UO_1430 (O_1430,N_14945,N_14735);
nand UO_1431 (O_1431,N_14451,N_14510);
and UO_1432 (O_1432,N_14922,N_14251);
nor UO_1433 (O_1433,N_14285,N_14819);
and UO_1434 (O_1434,N_14269,N_14337);
or UO_1435 (O_1435,N_14651,N_14360);
and UO_1436 (O_1436,N_14335,N_14684);
nand UO_1437 (O_1437,N_14349,N_14700);
or UO_1438 (O_1438,N_14622,N_14526);
or UO_1439 (O_1439,N_14990,N_14252);
nor UO_1440 (O_1440,N_14994,N_14889);
and UO_1441 (O_1441,N_14915,N_14875);
and UO_1442 (O_1442,N_14555,N_14837);
or UO_1443 (O_1443,N_14467,N_14748);
nand UO_1444 (O_1444,N_14492,N_14402);
nand UO_1445 (O_1445,N_14856,N_14609);
or UO_1446 (O_1446,N_14542,N_14683);
nand UO_1447 (O_1447,N_14920,N_14997);
or UO_1448 (O_1448,N_14327,N_14304);
nand UO_1449 (O_1449,N_14538,N_14339);
xor UO_1450 (O_1450,N_14420,N_14454);
nor UO_1451 (O_1451,N_14434,N_14982);
nand UO_1452 (O_1452,N_14658,N_14600);
nand UO_1453 (O_1453,N_14894,N_14906);
and UO_1454 (O_1454,N_14867,N_14665);
or UO_1455 (O_1455,N_14276,N_14433);
nand UO_1456 (O_1456,N_14983,N_14368);
nand UO_1457 (O_1457,N_14587,N_14747);
nand UO_1458 (O_1458,N_14787,N_14751);
nand UO_1459 (O_1459,N_14931,N_14789);
nand UO_1460 (O_1460,N_14668,N_14655);
nor UO_1461 (O_1461,N_14317,N_14849);
or UO_1462 (O_1462,N_14791,N_14870);
or UO_1463 (O_1463,N_14847,N_14624);
and UO_1464 (O_1464,N_14379,N_14663);
or UO_1465 (O_1465,N_14634,N_14962);
nor UO_1466 (O_1466,N_14888,N_14679);
nand UO_1467 (O_1467,N_14477,N_14735);
nand UO_1468 (O_1468,N_14891,N_14930);
or UO_1469 (O_1469,N_14775,N_14633);
xor UO_1470 (O_1470,N_14567,N_14309);
nor UO_1471 (O_1471,N_14253,N_14713);
nand UO_1472 (O_1472,N_14692,N_14641);
nand UO_1473 (O_1473,N_14526,N_14486);
or UO_1474 (O_1474,N_14605,N_14405);
nand UO_1475 (O_1475,N_14325,N_14329);
nand UO_1476 (O_1476,N_14478,N_14394);
or UO_1477 (O_1477,N_14485,N_14326);
and UO_1478 (O_1478,N_14827,N_14566);
and UO_1479 (O_1479,N_14559,N_14343);
or UO_1480 (O_1480,N_14745,N_14604);
nor UO_1481 (O_1481,N_14700,N_14511);
xor UO_1482 (O_1482,N_14412,N_14375);
or UO_1483 (O_1483,N_14288,N_14301);
and UO_1484 (O_1484,N_14447,N_14612);
nand UO_1485 (O_1485,N_14401,N_14863);
or UO_1486 (O_1486,N_14761,N_14264);
nor UO_1487 (O_1487,N_14941,N_14250);
xnor UO_1488 (O_1488,N_14707,N_14873);
xor UO_1489 (O_1489,N_14365,N_14568);
nand UO_1490 (O_1490,N_14900,N_14492);
or UO_1491 (O_1491,N_14556,N_14567);
or UO_1492 (O_1492,N_14478,N_14887);
nor UO_1493 (O_1493,N_14614,N_14916);
nor UO_1494 (O_1494,N_14830,N_14508);
nand UO_1495 (O_1495,N_14792,N_14832);
and UO_1496 (O_1496,N_14752,N_14300);
xor UO_1497 (O_1497,N_14396,N_14424);
nor UO_1498 (O_1498,N_14776,N_14668);
or UO_1499 (O_1499,N_14930,N_14560);
and UO_1500 (O_1500,N_14278,N_14575);
or UO_1501 (O_1501,N_14600,N_14784);
or UO_1502 (O_1502,N_14960,N_14569);
and UO_1503 (O_1503,N_14944,N_14310);
xnor UO_1504 (O_1504,N_14855,N_14540);
nor UO_1505 (O_1505,N_14719,N_14626);
xor UO_1506 (O_1506,N_14740,N_14460);
nor UO_1507 (O_1507,N_14421,N_14629);
and UO_1508 (O_1508,N_14729,N_14299);
nor UO_1509 (O_1509,N_14764,N_14491);
and UO_1510 (O_1510,N_14887,N_14886);
nand UO_1511 (O_1511,N_14822,N_14321);
and UO_1512 (O_1512,N_14340,N_14500);
or UO_1513 (O_1513,N_14734,N_14314);
nor UO_1514 (O_1514,N_14655,N_14522);
nor UO_1515 (O_1515,N_14927,N_14867);
or UO_1516 (O_1516,N_14711,N_14309);
nand UO_1517 (O_1517,N_14842,N_14853);
xnor UO_1518 (O_1518,N_14521,N_14983);
nand UO_1519 (O_1519,N_14281,N_14805);
nor UO_1520 (O_1520,N_14272,N_14375);
nor UO_1521 (O_1521,N_14572,N_14708);
nor UO_1522 (O_1522,N_14519,N_14774);
or UO_1523 (O_1523,N_14615,N_14510);
and UO_1524 (O_1524,N_14332,N_14382);
xor UO_1525 (O_1525,N_14591,N_14299);
and UO_1526 (O_1526,N_14897,N_14579);
nand UO_1527 (O_1527,N_14304,N_14655);
or UO_1528 (O_1528,N_14453,N_14748);
or UO_1529 (O_1529,N_14427,N_14685);
and UO_1530 (O_1530,N_14389,N_14951);
and UO_1531 (O_1531,N_14972,N_14576);
nor UO_1532 (O_1532,N_14280,N_14391);
nor UO_1533 (O_1533,N_14403,N_14355);
nand UO_1534 (O_1534,N_14299,N_14437);
or UO_1535 (O_1535,N_14953,N_14769);
nor UO_1536 (O_1536,N_14510,N_14594);
or UO_1537 (O_1537,N_14398,N_14978);
or UO_1538 (O_1538,N_14370,N_14585);
nor UO_1539 (O_1539,N_14890,N_14422);
and UO_1540 (O_1540,N_14837,N_14461);
or UO_1541 (O_1541,N_14820,N_14799);
or UO_1542 (O_1542,N_14920,N_14950);
and UO_1543 (O_1543,N_14622,N_14589);
nand UO_1544 (O_1544,N_14322,N_14767);
nor UO_1545 (O_1545,N_14523,N_14453);
nand UO_1546 (O_1546,N_14766,N_14294);
nor UO_1547 (O_1547,N_14737,N_14660);
and UO_1548 (O_1548,N_14725,N_14904);
nor UO_1549 (O_1549,N_14649,N_14279);
and UO_1550 (O_1550,N_14384,N_14893);
or UO_1551 (O_1551,N_14600,N_14320);
nand UO_1552 (O_1552,N_14801,N_14649);
or UO_1553 (O_1553,N_14731,N_14518);
and UO_1554 (O_1554,N_14313,N_14331);
and UO_1555 (O_1555,N_14349,N_14910);
nor UO_1556 (O_1556,N_14540,N_14792);
nand UO_1557 (O_1557,N_14597,N_14422);
nor UO_1558 (O_1558,N_14851,N_14691);
and UO_1559 (O_1559,N_14969,N_14321);
nor UO_1560 (O_1560,N_14904,N_14807);
nor UO_1561 (O_1561,N_14349,N_14643);
nor UO_1562 (O_1562,N_14971,N_14493);
or UO_1563 (O_1563,N_14472,N_14896);
and UO_1564 (O_1564,N_14397,N_14742);
nor UO_1565 (O_1565,N_14911,N_14919);
and UO_1566 (O_1566,N_14659,N_14539);
nor UO_1567 (O_1567,N_14505,N_14305);
and UO_1568 (O_1568,N_14391,N_14333);
or UO_1569 (O_1569,N_14508,N_14253);
or UO_1570 (O_1570,N_14826,N_14931);
and UO_1571 (O_1571,N_14404,N_14261);
or UO_1572 (O_1572,N_14304,N_14251);
nand UO_1573 (O_1573,N_14780,N_14255);
nand UO_1574 (O_1574,N_14951,N_14889);
or UO_1575 (O_1575,N_14910,N_14917);
or UO_1576 (O_1576,N_14471,N_14352);
nand UO_1577 (O_1577,N_14770,N_14775);
nand UO_1578 (O_1578,N_14277,N_14297);
or UO_1579 (O_1579,N_14951,N_14752);
or UO_1580 (O_1580,N_14724,N_14692);
nand UO_1581 (O_1581,N_14669,N_14454);
nor UO_1582 (O_1582,N_14975,N_14999);
nand UO_1583 (O_1583,N_14919,N_14493);
nor UO_1584 (O_1584,N_14473,N_14354);
nor UO_1585 (O_1585,N_14966,N_14328);
nand UO_1586 (O_1586,N_14601,N_14841);
nor UO_1587 (O_1587,N_14493,N_14397);
nand UO_1588 (O_1588,N_14861,N_14484);
or UO_1589 (O_1589,N_14900,N_14414);
and UO_1590 (O_1590,N_14261,N_14886);
and UO_1591 (O_1591,N_14832,N_14803);
and UO_1592 (O_1592,N_14577,N_14358);
xor UO_1593 (O_1593,N_14623,N_14782);
xnor UO_1594 (O_1594,N_14406,N_14337);
nor UO_1595 (O_1595,N_14961,N_14834);
and UO_1596 (O_1596,N_14286,N_14798);
and UO_1597 (O_1597,N_14986,N_14864);
nand UO_1598 (O_1598,N_14690,N_14933);
nand UO_1599 (O_1599,N_14413,N_14599);
or UO_1600 (O_1600,N_14570,N_14576);
or UO_1601 (O_1601,N_14672,N_14968);
nor UO_1602 (O_1602,N_14735,N_14907);
and UO_1603 (O_1603,N_14924,N_14878);
nor UO_1604 (O_1604,N_14933,N_14793);
and UO_1605 (O_1605,N_14492,N_14670);
nor UO_1606 (O_1606,N_14568,N_14702);
nand UO_1607 (O_1607,N_14403,N_14689);
nor UO_1608 (O_1608,N_14262,N_14870);
nor UO_1609 (O_1609,N_14843,N_14326);
nor UO_1610 (O_1610,N_14704,N_14468);
or UO_1611 (O_1611,N_14745,N_14849);
nor UO_1612 (O_1612,N_14255,N_14661);
nor UO_1613 (O_1613,N_14741,N_14828);
nor UO_1614 (O_1614,N_14615,N_14551);
nor UO_1615 (O_1615,N_14451,N_14905);
or UO_1616 (O_1616,N_14506,N_14332);
and UO_1617 (O_1617,N_14482,N_14602);
and UO_1618 (O_1618,N_14498,N_14770);
and UO_1619 (O_1619,N_14353,N_14797);
nor UO_1620 (O_1620,N_14691,N_14872);
nand UO_1621 (O_1621,N_14984,N_14392);
and UO_1622 (O_1622,N_14401,N_14817);
xor UO_1623 (O_1623,N_14854,N_14476);
nor UO_1624 (O_1624,N_14701,N_14788);
nand UO_1625 (O_1625,N_14349,N_14470);
or UO_1626 (O_1626,N_14491,N_14521);
and UO_1627 (O_1627,N_14641,N_14654);
nor UO_1628 (O_1628,N_14883,N_14851);
or UO_1629 (O_1629,N_14269,N_14251);
xor UO_1630 (O_1630,N_14535,N_14532);
or UO_1631 (O_1631,N_14992,N_14465);
and UO_1632 (O_1632,N_14320,N_14531);
nand UO_1633 (O_1633,N_14438,N_14747);
nand UO_1634 (O_1634,N_14557,N_14730);
and UO_1635 (O_1635,N_14335,N_14489);
nand UO_1636 (O_1636,N_14509,N_14804);
xor UO_1637 (O_1637,N_14876,N_14417);
xor UO_1638 (O_1638,N_14633,N_14789);
and UO_1639 (O_1639,N_14677,N_14595);
nor UO_1640 (O_1640,N_14898,N_14722);
nand UO_1641 (O_1641,N_14574,N_14301);
xnor UO_1642 (O_1642,N_14743,N_14802);
nand UO_1643 (O_1643,N_14650,N_14550);
or UO_1644 (O_1644,N_14932,N_14791);
or UO_1645 (O_1645,N_14272,N_14285);
nor UO_1646 (O_1646,N_14430,N_14497);
nor UO_1647 (O_1647,N_14314,N_14651);
or UO_1648 (O_1648,N_14700,N_14338);
or UO_1649 (O_1649,N_14449,N_14611);
and UO_1650 (O_1650,N_14693,N_14478);
nand UO_1651 (O_1651,N_14889,N_14849);
nor UO_1652 (O_1652,N_14937,N_14829);
nor UO_1653 (O_1653,N_14516,N_14712);
or UO_1654 (O_1654,N_14379,N_14721);
and UO_1655 (O_1655,N_14849,N_14475);
nand UO_1656 (O_1656,N_14732,N_14929);
or UO_1657 (O_1657,N_14880,N_14515);
nand UO_1658 (O_1658,N_14271,N_14868);
or UO_1659 (O_1659,N_14459,N_14639);
xnor UO_1660 (O_1660,N_14688,N_14338);
nor UO_1661 (O_1661,N_14669,N_14674);
nand UO_1662 (O_1662,N_14480,N_14681);
nor UO_1663 (O_1663,N_14250,N_14654);
and UO_1664 (O_1664,N_14647,N_14925);
xor UO_1665 (O_1665,N_14892,N_14473);
or UO_1666 (O_1666,N_14936,N_14343);
nand UO_1667 (O_1667,N_14632,N_14706);
nor UO_1668 (O_1668,N_14699,N_14418);
or UO_1669 (O_1669,N_14870,N_14736);
nand UO_1670 (O_1670,N_14869,N_14509);
nor UO_1671 (O_1671,N_14297,N_14632);
and UO_1672 (O_1672,N_14365,N_14591);
nand UO_1673 (O_1673,N_14328,N_14949);
and UO_1674 (O_1674,N_14736,N_14906);
nor UO_1675 (O_1675,N_14370,N_14528);
nand UO_1676 (O_1676,N_14900,N_14944);
and UO_1677 (O_1677,N_14872,N_14519);
nand UO_1678 (O_1678,N_14477,N_14675);
nand UO_1679 (O_1679,N_14678,N_14652);
xor UO_1680 (O_1680,N_14444,N_14600);
nor UO_1681 (O_1681,N_14418,N_14293);
and UO_1682 (O_1682,N_14854,N_14745);
and UO_1683 (O_1683,N_14461,N_14269);
or UO_1684 (O_1684,N_14427,N_14887);
nor UO_1685 (O_1685,N_14785,N_14864);
nor UO_1686 (O_1686,N_14723,N_14889);
or UO_1687 (O_1687,N_14626,N_14990);
and UO_1688 (O_1688,N_14634,N_14421);
xnor UO_1689 (O_1689,N_14251,N_14614);
nand UO_1690 (O_1690,N_14312,N_14821);
and UO_1691 (O_1691,N_14890,N_14902);
nor UO_1692 (O_1692,N_14675,N_14383);
nand UO_1693 (O_1693,N_14996,N_14397);
nor UO_1694 (O_1694,N_14250,N_14587);
nor UO_1695 (O_1695,N_14950,N_14266);
nor UO_1696 (O_1696,N_14812,N_14327);
nor UO_1697 (O_1697,N_14406,N_14601);
nand UO_1698 (O_1698,N_14687,N_14366);
xnor UO_1699 (O_1699,N_14314,N_14555);
and UO_1700 (O_1700,N_14950,N_14587);
and UO_1701 (O_1701,N_14661,N_14303);
and UO_1702 (O_1702,N_14568,N_14335);
and UO_1703 (O_1703,N_14550,N_14384);
and UO_1704 (O_1704,N_14617,N_14441);
nand UO_1705 (O_1705,N_14564,N_14882);
xor UO_1706 (O_1706,N_14935,N_14698);
nand UO_1707 (O_1707,N_14387,N_14697);
nand UO_1708 (O_1708,N_14948,N_14582);
nand UO_1709 (O_1709,N_14653,N_14705);
nand UO_1710 (O_1710,N_14339,N_14432);
and UO_1711 (O_1711,N_14536,N_14544);
nor UO_1712 (O_1712,N_14880,N_14798);
or UO_1713 (O_1713,N_14711,N_14457);
and UO_1714 (O_1714,N_14878,N_14856);
nand UO_1715 (O_1715,N_14612,N_14601);
and UO_1716 (O_1716,N_14555,N_14541);
nor UO_1717 (O_1717,N_14941,N_14600);
or UO_1718 (O_1718,N_14760,N_14539);
xor UO_1719 (O_1719,N_14494,N_14383);
xnor UO_1720 (O_1720,N_14613,N_14724);
nor UO_1721 (O_1721,N_14436,N_14586);
nand UO_1722 (O_1722,N_14494,N_14783);
nor UO_1723 (O_1723,N_14531,N_14396);
nor UO_1724 (O_1724,N_14334,N_14538);
and UO_1725 (O_1725,N_14396,N_14601);
nand UO_1726 (O_1726,N_14855,N_14626);
nor UO_1727 (O_1727,N_14535,N_14867);
xor UO_1728 (O_1728,N_14953,N_14467);
or UO_1729 (O_1729,N_14676,N_14967);
and UO_1730 (O_1730,N_14819,N_14484);
or UO_1731 (O_1731,N_14724,N_14517);
nand UO_1732 (O_1732,N_14830,N_14522);
nand UO_1733 (O_1733,N_14263,N_14255);
nand UO_1734 (O_1734,N_14736,N_14615);
nor UO_1735 (O_1735,N_14651,N_14646);
and UO_1736 (O_1736,N_14953,N_14541);
nand UO_1737 (O_1737,N_14981,N_14308);
nand UO_1738 (O_1738,N_14995,N_14974);
nand UO_1739 (O_1739,N_14428,N_14546);
and UO_1740 (O_1740,N_14382,N_14496);
or UO_1741 (O_1741,N_14367,N_14290);
xor UO_1742 (O_1742,N_14836,N_14252);
or UO_1743 (O_1743,N_14781,N_14491);
nor UO_1744 (O_1744,N_14267,N_14658);
nor UO_1745 (O_1745,N_14604,N_14825);
xor UO_1746 (O_1746,N_14589,N_14986);
nand UO_1747 (O_1747,N_14395,N_14346);
or UO_1748 (O_1748,N_14959,N_14269);
or UO_1749 (O_1749,N_14704,N_14543);
and UO_1750 (O_1750,N_14976,N_14741);
xnor UO_1751 (O_1751,N_14501,N_14463);
nor UO_1752 (O_1752,N_14808,N_14926);
or UO_1753 (O_1753,N_14479,N_14816);
or UO_1754 (O_1754,N_14899,N_14835);
and UO_1755 (O_1755,N_14547,N_14314);
nor UO_1756 (O_1756,N_14343,N_14833);
nand UO_1757 (O_1757,N_14667,N_14646);
and UO_1758 (O_1758,N_14378,N_14257);
or UO_1759 (O_1759,N_14551,N_14309);
nand UO_1760 (O_1760,N_14670,N_14770);
nor UO_1761 (O_1761,N_14569,N_14529);
nand UO_1762 (O_1762,N_14859,N_14934);
nor UO_1763 (O_1763,N_14895,N_14265);
and UO_1764 (O_1764,N_14620,N_14978);
or UO_1765 (O_1765,N_14554,N_14988);
xnor UO_1766 (O_1766,N_14744,N_14419);
nand UO_1767 (O_1767,N_14386,N_14970);
and UO_1768 (O_1768,N_14891,N_14691);
nor UO_1769 (O_1769,N_14919,N_14768);
and UO_1770 (O_1770,N_14907,N_14628);
nor UO_1771 (O_1771,N_14523,N_14394);
nor UO_1772 (O_1772,N_14631,N_14501);
and UO_1773 (O_1773,N_14607,N_14741);
or UO_1774 (O_1774,N_14808,N_14622);
or UO_1775 (O_1775,N_14383,N_14491);
nor UO_1776 (O_1776,N_14899,N_14455);
nor UO_1777 (O_1777,N_14697,N_14291);
and UO_1778 (O_1778,N_14944,N_14957);
xor UO_1779 (O_1779,N_14629,N_14488);
xnor UO_1780 (O_1780,N_14406,N_14837);
and UO_1781 (O_1781,N_14316,N_14612);
and UO_1782 (O_1782,N_14689,N_14815);
and UO_1783 (O_1783,N_14406,N_14761);
nor UO_1784 (O_1784,N_14928,N_14732);
nand UO_1785 (O_1785,N_14931,N_14735);
nand UO_1786 (O_1786,N_14959,N_14628);
and UO_1787 (O_1787,N_14678,N_14668);
or UO_1788 (O_1788,N_14394,N_14341);
or UO_1789 (O_1789,N_14931,N_14470);
nor UO_1790 (O_1790,N_14354,N_14416);
nor UO_1791 (O_1791,N_14517,N_14974);
nand UO_1792 (O_1792,N_14414,N_14912);
nor UO_1793 (O_1793,N_14684,N_14521);
or UO_1794 (O_1794,N_14444,N_14589);
nor UO_1795 (O_1795,N_14964,N_14405);
and UO_1796 (O_1796,N_14676,N_14597);
nor UO_1797 (O_1797,N_14266,N_14422);
xor UO_1798 (O_1798,N_14580,N_14343);
and UO_1799 (O_1799,N_14660,N_14877);
and UO_1800 (O_1800,N_14923,N_14614);
nor UO_1801 (O_1801,N_14825,N_14424);
and UO_1802 (O_1802,N_14455,N_14417);
or UO_1803 (O_1803,N_14696,N_14569);
nor UO_1804 (O_1804,N_14710,N_14411);
and UO_1805 (O_1805,N_14958,N_14670);
nand UO_1806 (O_1806,N_14827,N_14626);
or UO_1807 (O_1807,N_14857,N_14355);
and UO_1808 (O_1808,N_14375,N_14443);
nand UO_1809 (O_1809,N_14333,N_14549);
and UO_1810 (O_1810,N_14671,N_14880);
nor UO_1811 (O_1811,N_14327,N_14704);
or UO_1812 (O_1812,N_14882,N_14507);
nor UO_1813 (O_1813,N_14895,N_14902);
nor UO_1814 (O_1814,N_14641,N_14976);
xor UO_1815 (O_1815,N_14338,N_14576);
and UO_1816 (O_1816,N_14983,N_14377);
and UO_1817 (O_1817,N_14580,N_14932);
nor UO_1818 (O_1818,N_14831,N_14903);
nor UO_1819 (O_1819,N_14695,N_14386);
nor UO_1820 (O_1820,N_14942,N_14530);
nor UO_1821 (O_1821,N_14531,N_14637);
nand UO_1822 (O_1822,N_14885,N_14918);
and UO_1823 (O_1823,N_14560,N_14409);
nand UO_1824 (O_1824,N_14355,N_14452);
nor UO_1825 (O_1825,N_14714,N_14618);
nand UO_1826 (O_1826,N_14856,N_14745);
or UO_1827 (O_1827,N_14518,N_14872);
and UO_1828 (O_1828,N_14267,N_14811);
nor UO_1829 (O_1829,N_14299,N_14880);
and UO_1830 (O_1830,N_14469,N_14500);
and UO_1831 (O_1831,N_14993,N_14271);
nand UO_1832 (O_1832,N_14277,N_14906);
or UO_1833 (O_1833,N_14392,N_14504);
nor UO_1834 (O_1834,N_14794,N_14392);
nor UO_1835 (O_1835,N_14872,N_14692);
xnor UO_1836 (O_1836,N_14552,N_14939);
nor UO_1837 (O_1837,N_14680,N_14413);
and UO_1838 (O_1838,N_14871,N_14855);
nor UO_1839 (O_1839,N_14955,N_14352);
and UO_1840 (O_1840,N_14694,N_14786);
nor UO_1841 (O_1841,N_14845,N_14916);
nand UO_1842 (O_1842,N_14351,N_14396);
or UO_1843 (O_1843,N_14895,N_14794);
nor UO_1844 (O_1844,N_14751,N_14252);
nand UO_1845 (O_1845,N_14439,N_14601);
or UO_1846 (O_1846,N_14816,N_14908);
nand UO_1847 (O_1847,N_14438,N_14504);
xnor UO_1848 (O_1848,N_14761,N_14691);
nand UO_1849 (O_1849,N_14499,N_14670);
xor UO_1850 (O_1850,N_14486,N_14872);
nor UO_1851 (O_1851,N_14427,N_14889);
xnor UO_1852 (O_1852,N_14952,N_14435);
nor UO_1853 (O_1853,N_14718,N_14978);
nor UO_1854 (O_1854,N_14500,N_14355);
and UO_1855 (O_1855,N_14501,N_14642);
and UO_1856 (O_1856,N_14285,N_14820);
nor UO_1857 (O_1857,N_14780,N_14746);
and UO_1858 (O_1858,N_14250,N_14937);
xnor UO_1859 (O_1859,N_14286,N_14722);
xor UO_1860 (O_1860,N_14519,N_14816);
and UO_1861 (O_1861,N_14738,N_14703);
nand UO_1862 (O_1862,N_14549,N_14608);
nor UO_1863 (O_1863,N_14636,N_14536);
and UO_1864 (O_1864,N_14953,N_14949);
and UO_1865 (O_1865,N_14498,N_14275);
nor UO_1866 (O_1866,N_14634,N_14979);
nand UO_1867 (O_1867,N_14264,N_14457);
nand UO_1868 (O_1868,N_14890,N_14745);
or UO_1869 (O_1869,N_14344,N_14299);
or UO_1870 (O_1870,N_14766,N_14650);
and UO_1871 (O_1871,N_14751,N_14542);
nand UO_1872 (O_1872,N_14766,N_14397);
nor UO_1873 (O_1873,N_14883,N_14600);
and UO_1874 (O_1874,N_14774,N_14286);
xor UO_1875 (O_1875,N_14423,N_14776);
or UO_1876 (O_1876,N_14716,N_14464);
and UO_1877 (O_1877,N_14290,N_14665);
nor UO_1878 (O_1878,N_14799,N_14654);
and UO_1879 (O_1879,N_14930,N_14929);
and UO_1880 (O_1880,N_14289,N_14676);
or UO_1881 (O_1881,N_14517,N_14274);
and UO_1882 (O_1882,N_14967,N_14635);
and UO_1883 (O_1883,N_14277,N_14376);
nor UO_1884 (O_1884,N_14672,N_14552);
nand UO_1885 (O_1885,N_14721,N_14776);
nand UO_1886 (O_1886,N_14373,N_14864);
nor UO_1887 (O_1887,N_14299,N_14825);
or UO_1888 (O_1888,N_14379,N_14950);
and UO_1889 (O_1889,N_14391,N_14544);
xnor UO_1890 (O_1890,N_14549,N_14361);
nand UO_1891 (O_1891,N_14670,N_14387);
nand UO_1892 (O_1892,N_14306,N_14660);
nand UO_1893 (O_1893,N_14336,N_14985);
or UO_1894 (O_1894,N_14698,N_14772);
xnor UO_1895 (O_1895,N_14981,N_14722);
and UO_1896 (O_1896,N_14423,N_14524);
nand UO_1897 (O_1897,N_14668,N_14375);
xnor UO_1898 (O_1898,N_14818,N_14702);
xor UO_1899 (O_1899,N_14826,N_14299);
and UO_1900 (O_1900,N_14846,N_14775);
and UO_1901 (O_1901,N_14756,N_14693);
nand UO_1902 (O_1902,N_14262,N_14991);
and UO_1903 (O_1903,N_14285,N_14335);
and UO_1904 (O_1904,N_14687,N_14514);
or UO_1905 (O_1905,N_14803,N_14971);
or UO_1906 (O_1906,N_14771,N_14753);
nor UO_1907 (O_1907,N_14495,N_14744);
nor UO_1908 (O_1908,N_14309,N_14326);
nor UO_1909 (O_1909,N_14955,N_14818);
nand UO_1910 (O_1910,N_14670,N_14767);
and UO_1911 (O_1911,N_14433,N_14902);
and UO_1912 (O_1912,N_14621,N_14402);
and UO_1913 (O_1913,N_14902,N_14968);
nor UO_1914 (O_1914,N_14852,N_14901);
nor UO_1915 (O_1915,N_14652,N_14280);
nor UO_1916 (O_1916,N_14840,N_14768);
nand UO_1917 (O_1917,N_14584,N_14299);
and UO_1918 (O_1918,N_14841,N_14427);
and UO_1919 (O_1919,N_14791,N_14927);
nor UO_1920 (O_1920,N_14296,N_14991);
nand UO_1921 (O_1921,N_14800,N_14775);
and UO_1922 (O_1922,N_14727,N_14612);
and UO_1923 (O_1923,N_14715,N_14341);
nand UO_1924 (O_1924,N_14266,N_14316);
xor UO_1925 (O_1925,N_14277,N_14712);
xor UO_1926 (O_1926,N_14485,N_14374);
nand UO_1927 (O_1927,N_14833,N_14476);
and UO_1928 (O_1928,N_14907,N_14944);
or UO_1929 (O_1929,N_14742,N_14746);
xnor UO_1930 (O_1930,N_14799,N_14366);
or UO_1931 (O_1931,N_14603,N_14283);
nand UO_1932 (O_1932,N_14258,N_14972);
or UO_1933 (O_1933,N_14991,N_14965);
or UO_1934 (O_1934,N_14547,N_14536);
nor UO_1935 (O_1935,N_14309,N_14963);
and UO_1936 (O_1936,N_14630,N_14462);
and UO_1937 (O_1937,N_14848,N_14929);
nor UO_1938 (O_1938,N_14469,N_14951);
or UO_1939 (O_1939,N_14567,N_14781);
or UO_1940 (O_1940,N_14554,N_14978);
nand UO_1941 (O_1941,N_14448,N_14893);
and UO_1942 (O_1942,N_14361,N_14660);
xor UO_1943 (O_1943,N_14659,N_14696);
nand UO_1944 (O_1944,N_14723,N_14507);
or UO_1945 (O_1945,N_14416,N_14657);
or UO_1946 (O_1946,N_14511,N_14753);
or UO_1947 (O_1947,N_14435,N_14591);
or UO_1948 (O_1948,N_14496,N_14495);
nor UO_1949 (O_1949,N_14899,N_14638);
or UO_1950 (O_1950,N_14956,N_14862);
xor UO_1951 (O_1951,N_14814,N_14263);
xor UO_1952 (O_1952,N_14476,N_14401);
and UO_1953 (O_1953,N_14702,N_14279);
nand UO_1954 (O_1954,N_14616,N_14771);
and UO_1955 (O_1955,N_14374,N_14970);
and UO_1956 (O_1956,N_14369,N_14670);
and UO_1957 (O_1957,N_14453,N_14349);
nand UO_1958 (O_1958,N_14743,N_14525);
and UO_1959 (O_1959,N_14740,N_14602);
or UO_1960 (O_1960,N_14348,N_14856);
and UO_1961 (O_1961,N_14709,N_14966);
nand UO_1962 (O_1962,N_14818,N_14584);
nor UO_1963 (O_1963,N_14448,N_14983);
or UO_1964 (O_1964,N_14422,N_14406);
or UO_1965 (O_1965,N_14571,N_14506);
or UO_1966 (O_1966,N_14491,N_14353);
and UO_1967 (O_1967,N_14581,N_14544);
nor UO_1968 (O_1968,N_14511,N_14780);
nor UO_1969 (O_1969,N_14955,N_14529);
or UO_1970 (O_1970,N_14517,N_14956);
or UO_1971 (O_1971,N_14532,N_14784);
nand UO_1972 (O_1972,N_14807,N_14980);
nor UO_1973 (O_1973,N_14299,N_14842);
or UO_1974 (O_1974,N_14435,N_14935);
nand UO_1975 (O_1975,N_14711,N_14572);
and UO_1976 (O_1976,N_14757,N_14998);
or UO_1977 (O_1977,N_14432,N_14991);
nor UO_1978 (O_1978,N_14348,N_14801);
nor UO_1979 (O_1979,N_14720,N_14451);
or UO_1980 (O_1980,N_14956,N_14524);
and UO_1981 (O_1981,N_14561,N_14886);
nor UO_1982 (O_1982,N_14801,N_14693);
and UO_1983 (O_1983,N_14926,N_14258);
and UO_1984 (O_1984,N_14746,N_14789);
and UO_1985 (O_1985,N_14857,N_14327);
nand UO_1986 (O_1986,N_14842,N_14990);
and UO_1987 (O_1987,N_14801,N_14863);
and UO_1988 (O_1988,N_14710,N_14651);
nand UO_1989 (O_1989,N_14279,N_14773);
nor UO_1990 (O_1990,N_14650,N_14575);
xnor UO_1991 (O_1991,N_14782,N_14557);
nor UO_1992 (O_1992,N_14485,N_14980);
nand UO_1993 (O_1993,N_14574,N_14319);
and UO_1994 (O_1994,N_14578,N_14284);
nand UO_1995 (O_1995,N_14927,N_14963);
and UO_1996 (O_1996,N_14972,N_14825);
or UO_1997 (O_1997,N_14328,N_14401);
or UO_1998 (O_1998,N_14934,N_14858);
nand UO_1999 (O_1999,N_14622,N_14969);
endmodule