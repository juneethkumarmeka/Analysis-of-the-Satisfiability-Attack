module basic_500_3000_500_30_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_210,In_452);
nand U1 (N_1,In_60,In_248);
or U2 (N_2,In_486,In_381);
or U3 (N_3,In_327,In_464);
nor U4 (N_4,In_445,In_296);
or U5 (N_5,In_304,In_402);
or U6 (N_6,In_328,In_130);
and U7 (N_7,In_498,In_140);
nor U8 (N_8,In_433,In_474);
or U9 (N_9,In_305,In_90);
nor U10 (N_10,In_212,In_404);
nand U11 (N_11,In_367,In_182);
xor U12 (N_12,In_384,In_75);
or U13 (N_13,In_164,In_320);
and U14 (N_14,In_66,In_11);
and U15 (N_15,In_256,In_123);
nand U16 (N_16,In_370,In_176);
and U17 (N_17,In_293,In_205);
nand U18 (N_18,In_266,In_326);
nor U19 (N_19,In_349,In_400);
and U20 (N_20,In_110,In_442);
and U21 (N_21,In_218,In_59);
or U22 (N_22,In_382,In_309);
and U23 (N_23,In_280,In_149);
nand U24 (N_24,In_343,In_314);
nand U25 (N_25,In_50,In_12);
xor U26 (N_26,In_481,In_128);
nor U27 (N_27,In_431,In_156);
nor U28 (N_28,In_335,In_67);
and U29 (N_29,In_412,In_117);
or U30 (N_30,In_261,In_341);
and U31 (N_31,In_19,In_145);
and U32 (N_32,In_245,In_365);
xnor U33 (N_33,In_23,In_71);
or U34 (N_34,In_83,In_70);
nor U35 (N_35,In_397,In_17);
or U36 (N_36,In_371,In_4);
and U37 (N_37,In_153,In_268);
xnor U38 (N_38,In_480,In_73);
and U39 (N_39,In_306,In_16);
or U40 (N_40,In_143,In_58);
nand U41 (N_41,In_134,In_3);
nand U42 (N_42,In_279,In_62);
nor U43 (N_43,In_129,In_426);
nor U44 (N_44,In_340,In_286);
xor U45 (N_45,In_72,In_411);
or U46 (N_46,In_438,In_109);
or U47 (N_47,In_312,In_232);
nand U48 (N_48,In_186,In_177);
nor U49 (N_49,In_291,In_81);
nor U50 (N_50,In_420,In_479);
nand U51 (N_51,In_389,In_394);
nand U52 (N_52,In_100,In_220);
xor U53 (N_53,In_355,In_251);
nand U54 (N_54,In_54,In_234);
or U55 (N_55,In_409,In_250);
and U56 (N_56,In_278,In_263);
nor U57 (N_57,In_388,In_357);
or U58 (N_58,In_133,In_347);
nand U59 (N_59,In_275,In_471);
nand U60 (N_60,In_387,In_132);
or U61 (N_61,In_437,In_424);
nor U62 (N_62,In_175,In_353);
or U63 (N_63,In_47,In_354);
nor U64 (N_64,In_1,In_368);
nor U65 (N_65,In_206,In_316);
xnor U66 (N_66,In_336,In_484);
nand U67 (N_67,In_141,In_489);
nor U68 (N_68,In_473,In_152);
nand U69 (N_69,In_274,In_85);
nor U70 (N_70,In_138,In_462);
nor U71 (N_71,In_77,In_399);
or U72 (N_72,In_364,In_151);
and U73 (N_73,In_300,In_262);
nand U74 (N_74,In_475,In_324);
nand U75 (N_75,In_289,In_254);
nand U76 (N_76,In_61,In_159);
nand U77 (N_77,In_491,In_162);
nor U78 (N_78,In_242,In_361);
nor U79 (N_79,In_284,In_375);
or U80 (N_80,In_160,In_416);
nor U81 (N_81,In_377,In_376);
xnor U82 (N_82,In_43,In_202);
nor U83 (N_83,In_122,In_216);
and U84 (N_84,In_69,In_403);
xor U85 (N_85,In_302,In_239);
nor U86 (N_86,In_13,In_449);
nor U87 (N_87,In_84,In_200);
nand U88 (N_88,In_86,In_344);
nand U89 (N_89,In_476,In_22);
nand U90 (N_90,In_450,In_292);
and U91 (N_91,In_32,In_222);
nand U92 (N_92,In_112,In_319);
and U93 (N_93,In_482,In_163);
or U94 (N_94,In_135,In_42);
or U95 (N_95,In_435,In_187);
and U96 (N_96,In_391,In_421);
nand U97 (N_97,In_9,In_271);
and U98 (N_98,In_252,In_374);
nor U99 (N_99,In_283,In_45);
and U100 (N_100,N_34,In_217);
or U101 (N_101,In_315,In_459);
or U102 (N_102,N_33,N_65);
nor U103 (N_103,N_59,In_267);
nand U104 (N_104,N_87,In_229);
or U105 (N_105,N_93,In_178);
or U106 (N_106,In_258,In_429);
or U107 (N_107,In_104,In_166);
nand U108 (N_108,In_427,In_385);
or U109 (N_109,In_401,N_37);
and U110 (N_110,N_82,In_310);
and U111 (N_111,In_269,N_4);
or U112 (N_112,In_244,In_287);
xor U113 (N_113,In_398,In_10);
and U114 (N_114,In_246,In_236);
nand U115 (N_115,In_103,In_101);
nand U116 (N_116,N_94,In_80);
nor U117 (N_117,In_430,In_49);
and U118 (N_118,N_78,In_499);
nor U119 (N_119,N_66,N_41);
or U120 (N_120,N_58,In_494);
and U121 (N_121,In_333,N_53);
xor U122 (N_122,In_114,In_64);
nand U123 (N_123,In_76,N_23);
nor U124 (N_124,In_249,In_334);
or U125 (N_125,N_86,N_69);
and U126 (N_126,N_36,In_224);
nor U127 (N_127,N_46,In_243);
and U128 (N_128,In_440,In_55);
and U129 (N_129,In_139,In_35);
nor U130 (N_130,N_12,N_45);
nand U131 (N_131,In_18,In_63);
or U132 (N_132,In_225,In_276);
nor U133 (N_133,In_443,In_40);
or U134 (N_134,In_161,In_2);
nor U135 (N_135,In_99,In_28);
nand U136 (N_136,N_14,In_195);
and U137 (N_137,In_157,N_99);
nand U138 (N_138,In_406,In_339);
xor U139 (N_139,In_192,In_25);
or U140 (N_140,In_209,In_201);
nand U141 (N_141,In_115,In_348);
xnor U142 (N_142,In_392,In_360);
nor U143 (N_143,In_38,In_208);
nor U144 (N_144,N_7,N_90);
and U145 (N_145,N_83,In_5);
or U146 (N_146,In_193,N_0);
or U147 (N_147,N_3,In_463);
and U148 (N_148,In_94,In_317);
nand U149 (N_149,In_57,In_172);
or U150 (N_150,In_238,N_10);
nand U151 (N_151,In_264,In_277);
nor U152 (N_152,In_359,In_41);
or U153 (N_153,N_50,N_61);
or U154 (N_154,In_181,In_329);
and U155 (N_155,In_227,In_155);
nor U156 (N_156,In_457,In_386);
nand U157 (N_157,In_167,In_492);
or U158 (N_158,In_31,In_247);
xnor U159 (N_159,In_179,In_257);
and U160 (N_160,N_13,In_350);
and U161 (N_161,In_282,In_456);
nand U162 (N_162,In_230,In_235);
and U163 (N_163,In_95,N_71);
or U164 (N_164,In_418,In_211);
nor U165 (N_165,In_171,In_46);
xor U166 (N_166,In_121,In_165);
and U167 (N_167,In_288,In_154);
nand U168 (N_168,N_80,In_495);
nor U169 (N_169,In_342,N_55);
and U170 (N_170,In_33,In_96);
nor U171 (N_171,In_131,In_472);
nand U172 (N_172,N_39,In_307);
nand U173 (N_173,In_118,In_226);
nor U174 (N_174,In_15,In_441);
and U175 (N_175,In_26,In_39);
nand U176 (N_176,In_469,N_74);
and U177 (N_177,N_26,N_56);
and U178 (N_178,In_183,N_73);
xor U179 (N_179,In_219,In_383);
nand U180 (N_180,In_414,In_199);
xor U181 (N_181,In_273,In_228);
or U182 (N_182,In_322,In_147);
or U183 (N_183,In_444,In_108);
nand U184 (N_184,In_337,In_146);
or U185 (N_185,N_22,In_373);
nor U186 (N_186,N_1,In_150);
or U187 (N_187,N_88,In_170);
nor U188 (N_188,In_191,In_30);
xor U189 (N_189,In_126,N_48);
nor U190 (N_190,N_89,In_272);
nand U191 (N_191,In_423,N_96);
nor U192 (N_192,In_410,In_144);
or U193 (N_193,In_51,In_148);
nand U194 (N_194,In_113,In_318);
nor U195 (N_195,In_231,In_417);
nor U196 (N_196,In_56,In_7);
and U197 (N_197,N_9,In_408);
or U198 (N_198,N_52,In_79);
or U199 (N_199,N_64,In_203);
or U200 (N_200,In_378,N_125);
or U201 (N_201,In_413,N_110);
nor U202 (N_202,In_169,In_36);
nand U203 (N_203,N_137,N_196);
or U204 (N_204,N_126,N_138);
and U205 (N_205,N_167,In_197);
and U206 (N_206,In_173,In_14);
and U207 (N_207,N_95,In_92);
and U208 (N_208,N_146,In_298);
nor U209 (N_209,In_487,In_483);
or U210 (N_210,N_109,N_116);
nor U211 (N_211,N_32,In_20);
or U212 (N_212,N_120,N_57);
and U213 (N_213,N_67,In_93);
and U214 (N_214,N_147,N_152);
nor U215 (N_215,N_2,In_127);
or U216 (N_216,In_297,In_447);
nand U217 (N_217,In_116,N_124);
and U218 (N_218,N_114,N_148);
nand U219 (N_219,N_166,N_176);
or U220 (N_220,In_439,In_102);
nand U221 (N_221,In_460,In_380);
nor U222 (N_222,N_15,N_113);
or U223 (N_223,In_270,N_144);
or U224 (N_224,In_338,In_255);
or U225 (N_225,N_81,In_253);
and U226 (N_226,N_111,N_101);
nor U227 (N_227,N_118,N_195);
nor U228 (N_228,In_390,N_75);
and U229 (N_229,In_37,In_0);
nand U230 (N_230,In_265,In_330);
nor U231 (N_231,N_102,In_419);
nand U232 (N_232,In_290,In_496);
or U233 (N_233,N_131,In_393);
and U234 (N_234,In_260,N_30);
xor U235 (N_235,In_436,N_60);
nand U236 (N_236,N_158,In_120);
nand U237 (N_237,N_97,In_356);
or U238 (N_238,In_89,In_395);
nand U239 (N_239,N_100,In_27);
nand U240 (N_240,In_207,In_52);
or U241 (N_241,N_24,N_178);
and U242 (N_242,N_172,In_465);
nor U243 (N_243,In_68,N_145);
nand U244 (N_244,N_191,In_455);
nand U245 (N_245,In_454,In_281);
or U246 (N_246,In_405,N_157);
nor U247 (N_247,N_159,In_106);
and U248 (N_248,N_135,N_54);
nor U249 (N_249,N_6,N_108);
and U250 (N_250,In_237,In_34);
xnor U251 (N_251,N_171,N_162);
nor U252 (N_252,N_168,N_121);
and U253 (N_253,In_345,In_346);
nand U254 (N_254,In_485,In_451);
or U255 (N_255,In_497,N_112);
nor U256 (N_256,In_88,In_308);
or U257 (N_257,N_175,N_170);
and U258 (N_258,In_98,N_19);
nor U259 (N_259,In_490,N_184);
nand U260 (N_260,In_240,N_185);
nand U261 (N_261,N_142,N_130);
nand U262 (N_262,N_197,In_142);
nand U263 (N_263,N_105,N_11);
nand U264 (N_264,N_141,In_214);
nor U265 (N_265,N_163,N_77);
or U266 (N_266,N_179,In_351);
nand U267 (N_267,N_91,N_193);
nor U268 (N_268,In_223,In_466);
and U269 (N_269,N_8,N_183);
nor U270 (N_270,In_311,N_76);
or U271 (N_271,In_422,N_199);
xnor U272 (N_272,In_301,In_323);
or U273 (N_273,N_198,In_313);
or U274 (N_274,In_105,N_98);
nand U275 (N_275,N_62,In_24);
or U276 (N_276,In_198,In_488);
and U277 (N_277,N_154,In_358);
nand U278 (N_278,N_5,N_134);
and U279 (N_279,N_139,In_434);
nand U280 (N_280,In_458,In_366);
and U281 (N_281,N_106,In_137);
nor U282 (N_282,In_294,N_156);
nand U283 (N_283,In_352,N_35);
and U284 (N_284,N_16,In_158);
nor U285 (N_285,In_107,In_6);
or U286 (N_286,N_28,N_136);
nor U287 (N_287,In_204,In_493);
nand U288 (N_288,N_17,In_124);
and U289 (N_289,N_173,In_194);
xor U290 (N_290,N_20,In_432);
and U291 (N_291,N_72,N_169);
or U292 (N_292,In_321,N_68);
xnor U293 (N_293,In_259,In_233);
nand U294 (N_294,N_85,N_31);
or U295 (N_295,In_8,N_180);
xnor U296 (N_296,In_379,N_127);
or U297 (N_297,N_40,In_332);
nor U298 (N_298,N_164,N_155);
or U299 (N_299,In_48,In_363);
and U300 (N_300,In_82,N_216);
nor U301 (N_301,N_269,N_265);
nand U302 (N_302,N_243,N_293);
and U303 (N_303,In_470,N_149);
xor U304 (N_304,N_234,N_211);
or U305 (N_305,N_189,N_242);
and U306 (N_306,N_241,N_279);
nand U307 (N_307,N_208,N_217);
or U308 (N_308,N_119,N_294);
or U309 (N_309,N_133,N_233);
and U310 (N_310,N_186,In_21);
nor U311 (N_311,N_298,N_283);
or U312 (N_312,N_249,N_104);
xnor U313 (N_313,In_221,In_303);
or U314 (N_314,In_125,N_255);
and U315 (N_315,N_285,N_273);
xnor U316 (N_316,N_25,N_299);
or U317 (N_317,N_297,In_299);
or U318 (N_318,N_264,N_160);
nand U319 (N_319,N_219,N_271);
or U320 (N_320,N_103,N_246);
and U321 (N_321,N_115,N_128);
and U322 (N_322,N_272,N_51);
and U323 (N_323,N_181,In_295);
nand U324 (N_324,N_225,N_220);
nor U325 (N_325,N_280,In_478);
xnor U326 (N_326,N_92,N_276);
nor U327 (N_327,N_231,N_84);
nor U328 (N_328,N_213,In_189);
nor U329 (N_329,N_218,N_232);
nor U330 (N_330,N_221,In_362);
or U331 (N_331,N_222,N_245);
or U332 (N_332,N_256,N_79);
nor U333 (N_333,N_267,N_212);
or U334 (N_334,In_111,N_47);
nor U335 (N_335,N_227,N_44);
xor U336 (N_336,N_257,N_239);
nor U337 (N_337,N_200,N_165);
nor U338 (N_338,N_295,N_268);
and U339 (N_339,N_190,N_182);
or U340 (N_340,N_18,N_203);
nand U341 (N_341,N_206,In_174);
and U342 (N_342,In_168,N_274);
nand U343 (N_343,N_261,N_204);
nor U344 (N_344,In_29,N_122);
and U345 (N_345,N_150,N_174);
and U346 (N_346,In_428,N_214);
xor U347 (N_347,N_260,N_290);
xnor U348 (N_348,In_44,N_123);
nor U349 (N_349,N_188,N_132);
or U350 (N_350,N_235,N_129);
or U351 (N_351,N_177,N_202);
and U352 (N_352,N_151,In_467);
nor U353 (N_353,N_289,N_240);
xnor U354 (N_354,N_70,N_194);
and U355 (N_355,In_325,In_119);
or U356 (N_356,N_27,In_185);
or U357 (N_357,In_74,N_266);
nand U358 (N_358,In_196,N_43);
and U359 (N_359,In_136,N_237);
or U360 (N_360,N_250,N_238);
nor U361 (N_361,N_282,N_236);
or U362 (N_362,In_213,N_192);
nand U363 (N_363,In_241,N_278);
nor U364 (N_364,In_453,N_63);
nand U365 (N_365,In_446,N_140);
nor U366 (N_366,N_38,N_226);
nand U367 (N_367,N_262,N_277);
nand U368 (N_368,In_448,N_286);
xor U369 (N_369,N_153,In_215);
and U370 (N_370,N_275,In_468);
nor U371 (N_371,N_296,N_117);
xor U372 (N_372,N_210,N_107);
or U373 (N_373,N_244,N_292);
nand U374 (N_374,N_259,N_248);
nor U375 (N_375,N_253,In_97);
nor U376 (N_376,N_201,In_425);
and U377 (N_377,N_224,In_369);
nand U378 (N_378,N_258,N_281);
nand U379 (N_379,N_247,N_251);
and U380 (N_380,In_407,N_223);
or U381 (N_381,In_285,N_252);
nor U382 (N_382,N_215,N_29);
or U383 (N_383,N_284,In_87);
or U384 (N_384,In_91,In_78);
or U385 (N_385,N_209,In_331);
or U386 (N_386,N_42,In_372);
and U387 (N_387,N_291,In_396);
or U388 (N_388,N_270,N_287);
and U389 (N_389,In_461,N_143);
and U390 (N_390,N_161,In_477);
and U391 (N_391,N_230,N_228);
nor U392 (N_392,N_288,In_184);
xor U393 (N_393,N_49,N_263);
nand U394 (N_394,In_180,In_65);
xnor U395 (N_395,In_190,N_187);
nor U396 (N_396,In_188,N_229);
and U397 (N_397,N_254,N_205);
and U398 (N_398,N_21,In_53);
xor U399 (N_399,N_207,In_415);
nand U400 (N_400,N_357,N_330);
nor U401 (N_401,N_343,N_344);
nor U402 (N_402,N_310,N_308);
and U403 (N_403,N_389,N_394);
nor U404 (N_404,N_335,N_395);
nor U405 (N_405,N_320,N_307);
nor U406 (N_406,N_334,N_353);
and U407 (N_407,N_355,N_350);
or U408 (N_408,N_372,N_370);
nand U409 (N_409,N_393,N_329);
and U410 (N_410,N_374,N_348);
nor U411 (N_411,N_323,N_332);
and U412 (N_412,N_301,N_382);
xor U413 (N_413,N_352,N_302);
or U414 (N_414,N_309,N_311);
nand U415 (N_415,N_333,N_397);
nor U416 (N_416,N_387,N_327);
xor U417 (N_417,N_303,N_378);
or U418 (N_418,N_398,N_364);
nor U419 (N_419,N_306,N_347);
nor U420 (N_420,N_321,N_354);
nand U421 (N_421,N_388,N_319);
and U422 (N_422,N_375,N_304);
or U423 (N_423,N_358,N_300);
or U424 (N_424,N_346,N_324);
nor U425 (N_425,N_381,N_384);
nand U426 (N_426,N_326,N_315);
or U427 (N_427,N_318,N_386);
and U428 (N_428,N_396,N_383);
and U429 (N_429,N_369,N_345);
and U430 (N_430,N_341,N_392);
xor U431 (N_431,N_376,N_366);
xnor U432 (N_432,N_305,N_377);
nor U433 (N_433,N_360,N_328);
nor U434 (N_434,N_339,N_390);
nor U435 (N_435,N_316,N_361);
nor U436 (N_436,N_362,N_356);
and U437 (N_437,N_359,N_391);
or U438 (N_438,N_367,N_325);
xnor U439 (N_439,N_379,N_337);
nor U440 (N_440,N_351,N_317);
nor U441 (N_441,N_399,N_314);
nand U442 (N_442,N_312,N_336);
and U443 (N_443,N_338,N_380);
and U444 (N_444,N_363,N_371);
xnor U445 (N_445,N_385,N_322);
xor U446 (N_446,N_365,N_349);
nand U447 (N_447,N_331,N_368);
nand U448 (N_448,N_340,N_342);
xnor U449 (N_449,N_373,N_313);
and U450 (N_450,N_383,N_304);
nor U451 (N_451,N_367,N_395);
xor U452 (N_452,N_317,N_326);
nor U453 (N_453,N_313,N_368);
nand U454 (N_454,N_303,N_390);
nand U455 (N_455,N_398,N_370);
xor U456 (N_456,N_301,N_365);
or U457 (N_457,N_372,N_368);
and U458 (N_458,N_352,N_392);
nor U459 (N_459,N_329,N_302);
and U460 (N_460,N_311,N_393);
and U461 (N_461,N_360,N_346);
and U462 (N_462,N_318,N_378);
nand U463 (N_463,N_399,N_318);
nand U464 (N_464,N_353,N_303);
nor U465 (N_465,N_315,N_384);
nand U466 (N_466,N_338,N_361);
and U467 (N_467,N_362,N_390);
or U468 (N_468,N_337,N_361);
or U469 (N_469,N_348,N_307);
nand U470 (N_470,N_325,N_338);
nor U471 (N_471,N_378,N_312);
nor U472 (N_472,N_391,N_385);
nand U473 (N_473,N_380,N_302);
or U474 (N_474,N_327,N_350);
nor U475 (N_475,N_364,N_389);
nand U476 (N_476,N_337,N_376);
and U477 (N_477,N_394,N_378);
and U478 (N_478,N_314,N_374);
or U479 (N_479,N_337,N_325);
nor U480 (N_480,N_323,N_354);
xnor U481 (N_481,N_392,N_315);
or U482 (N_482,N_323,N_377);
nand U483 (N_483,N_307,N_323);
or U484 (N_484,N_375,N_340);
nand U485 (N_485,N_370,N_340);
nand U486 (N_486,N_371,N_336);
and U487 (N_487,N_354,N_349);
xor U488 (N_488,N_332,N_342);
or U489 (N_489,N_312,N_367);
or U490 (N_490,N_302,N_316);
nor U491 (N_491,N_327,N_328);
and U492 (N_492,N_309,N_337);
nor U493 (N_493,N_304,N_362);
or U494 (N_494,N_383,N_381);
nor U495 (N_495,N_392,N_300);
nand U496 (N_496,N_365,N_364);
nand U497 (N_497,N_328,N_308);
nor U498 (N_498,N_318,N_385);
nor U499 (N_499,N_361,N_393);
or U500 (N_500,N_483,N_403);
xor U501 (N_501,N_430,N_480);
or U502 (N_502,N_453,N_493);
or U503 (N_503,N_405,N_438);
nor U504 (N_504,N_425,N_489);
or U505 (N_505,N_432,N_441);
xnor U506 (N_506,N_478,N_461);
and U507 (N_507,N_427,N_408);
or U508 (N_508,N_467,N_463);
nor U509 (N_509,N_440,N_473);
nand U510 (N_510,N_486,N_423);
or U511 (N_511,N_499,N_419);
nor U512 (N_512,N_429,N_457);
nor U513 (N_513,N_455,N_417);
nor U514 (N_514,N_404,N_449);
or U515 (N_515,N_412,N_436);
nand U516 (N_516,N_495,N_435);
nor U517 (N_517,N_420,N_444);
nand U518 (N_518,N_418,N_487);
and U519 (N_519,N_410,N_496);
and U520 (N_520,N_459,N_465);
nand U521 (N_521,N_426,N_454);
nand U522 (N_522,N_460,N_470);
nand U523 (N_523,N_481,N_433);
nand U524 (N_524,N_450,N_456);
nand U525 (N_525,N_476,N_422);
nor U526 (N_526,N_409,N_402);
nand U527 (N_527,N_492,N_498);
xnor U528 (N_528,N_475,N_445);
xnor U529 (N_529,N_407,N_415);
or U530 (N_530,N_416,N_400);
nor U531 (N_531,N_411,N_431);
or U532 (N_532,N_413,N_448);
or U533 (N_533,N_494,N_434);
nand U534 (N_534,N_421,N_484);
nand U535 (N_535,N_443,N_442);
nand U536 (N_536,N_401,N_477);
nand U537 (N_537,N_479,N_462);
and U538 (N_538,N_439,N_490);
and U539 (N_539,N_452,N_466);
or U540 (N_540,N_464,N_488);
nand U541 (N_541,N_414,N_497);
nand U542 (N_542,N_437,N_406);
nand U543 (N_543,N_447,N_446);
nand U544 (N_544,N_474,N_458);
xor U545 (N_545,N_471,N_424);
nor U546 (N_546,N_472,N_482);
nor U547 (N_547,N_485,N_469);
nor U548 (N_548,N_451,N_468);
and U549 (N_549,N_491,N_428);
or U550 (N_550,N_496,N_424);
or U551 (N_551,N_422,N_420);
nor U552 (N_552,N_464,N_463);
and U553 (N_553,N_458,N_471);
xor U554 (N_554,N_492,N_494);
xnor U555 (N_555,N_493,N_439);
and U556 (N_556,N_477,N_480);
nor U557 (N_557,N_413,N_441);
nor U558 (N_558,N_435,N_464);
and U559 (N_559,N_451,N_495);
nor U560 (N_560,N_445,N_486);
and U561 (N_561,N_483,N_402);
nor U562 (N_562,N_490,N_434);
xor U563 (N_563,N_437,N_464);
and U564 (N_564,N_426,N_407);
or U565 (N_565,N_408,N_448);
nand U566 (N_566,N_434,N_431);
nand U567 (N_567,N_456,N_498);
or U568 (N_568,N_427,N_445);
nor U569 (N_569,N_470,N_418);
xor U570 (N_570,N_476,N_494);
or U571 (N_571,N_407,N_484);
and U572 (N_572,N_402,N_457);
and U573 (N_573,N_494,N_436);
or U574 (N_574,N_412,N_492);
and U575 (N_575,N_410,N_427);
nand U576 (N_576,N_498,N_450);
xnor U577 (N_577,N_495,N_406);
or U578 (N_578,N_438,N_435);
and U579 (N_579,N_459,N_470);
or U580 (N_580,N_498,N_433);
nand U581 (N_581,N_465,N_472);
or U582 (N_582,N_413,N_466);
and U583 (N_583,N_453,N_449);
and U584 (N_584,N_444,N_405);
or U585 (N_585,N_448,N_466);
xnor U586 (N_586,N_496,N_434);
or U587 (N_587,N_441,N_499);
nor U588 (N_588,N_447,N_443);
or U589 (N_589,N_446,N_440);
or U590 (N_590,N_438,N_471);
nor U591 (N_591,N_477,N_476);
and U592 (N_592,N_453,N_406);
nand U593 (N_593,N_468,N_466);
nand U594 (N_594,N_444,N_461);
nor U595 (N_595,N_454,N_436);
xnor U596 (N_596,N_471,N_491);
xor U597 (N_597,N_403,N_405);
nand U598 (N_598,N_437,N_474);
and U599 (N_599,N_442,N_448);
nor U600 (N_600,N_594,N_551);
and U601 (N_601,N_549,N_590);
xor U602 (N_602,N_524,N_514);
nor U603 (N_603,N_577,N_592);
and U604 (N_604,N_520,N_521);
or U605 (N_605,N_599,N_579);
nand U606 (N_606,N_571,N_540);
or U607 (N_607,N_554,N_563);
nand U608 (N_608,N_593,N_582);
nand U609 (N_609,N_509,N_531);
and U610 (N_610,N_576,N_552);
nor U611 (N_611,N_534,N_591);
nand U612 (N_612,N_532,N_556);
xnor U613 (N_613,N_589,N_544);
or U614 (N_614,N_557,N_567);
nor U615 (N_615,N_518,N_536);
nand U616 (N_616,N_501,N_538);
or U617 (N_617,N_580,N_596);
nand U618 (N_618,N_513,N_512);
and U619 (N_619,N_510,N_528);
nand U620 (N_620,N_530,N_539);
xor U621 (N_621,N_598,N_595);
nand U622 (N_622,N_533,N_535);
nor U623 (N_623,N_517,N_525);
or U624 (N_624,N_585,N_553);
xor U625 (N_625,N_566,N_555);
or U626 (N_626,N_565,N_541);
and U627 (N_627,N_503,N_561);
and U628 (N_628,N_507,N_574);
nand U629 (N_629,N_515,N_570);
nor U630 (N_630,N_581,N_527);
nand U631 (N_631,N_526,N_558);
xor U632 (N_632,N_559,N_562);
nor U633 (N_633,N_564,N_537);
or U634 (N_634,N_511,N_543);
nor U635 (N_635,N_568,N_584);
nand U636 (N_636,N_578,N_597);
and U637 (N_637,N_529,N_587);
nor U638 (N_638,N_516,N_500);
nor U639 (N_639,N_505,N_519);
nor U640 (N_640,N_550,N_560);
or U641 (N_641,N_502,N_522);
and U642 (N_642,N_583,N_545);
nand U643 (N_643,N_542,N_588);
nor U644 (N_644,N_508,N_523);
or U645 (N_645,N_575,N_506);
or U646 (N_646,N_569,N_504);
nand U647 (N_647,N_548,N_547);
and U648 (N_648,N_586,N_573);
or U649 (N_649,N_572,N_546);
nand U650 (N_650,N_587,N_536);
or U651 (N_651,N_528,N_554);
nand U652 (N_652,N_598,N_528);
or U653 (N_653,N_549,N_531);
xor U654 (N_654,N_514,N_516);
nand U655 (N_655,N_552,N_596);
and U656 (N_656,N_543,N_590);
nand U657 (N_657,N_589,N_502);
or U658 (N_658,N_548,N_553);
and U659 (N_659,N_558,N_523);
and U660 (N_660,N_526,N_519);
or U661 (N_661,N_553,N_524);
nand U662 (N_662,N_528,N_535);
nand U663 (N_663,N_534,N_515);
xnor U664 (N_664,N_537,N_590);
or U665 (N_665,N_551,N_592);
nand U666 (N_666,N_524,N_579);
nor U667 (N_667,N_514,N_527);
and U668 (N_668,N_521,N_503);
or U669 (N_669,N_531,N_565);
nand U670 (N_670,N_557,N_544);
xor U671 (N_671,N_582,N_579);
nor U672 (N_672,N_596,N_564);
nor U673 (N_673,N_523,N_593);
nand U674 (N_674,N_510,N_505);
nor U675 (N_675,N_560,N_508);
and U676 (N_676,N_560,N_500);
and U677 (N_677,N_512,N_551);
nand U678 (N_678,N_514,N_566);
or U679 (N_679,N_532,N_579);
nand U680 (N_680,N_593,N_561);
nand U681 (N_681,N_586,N_507);
and U682 (N_682,N_580,N_568);
xnor U683 (N_683,N_512,N_599);
or U684 (N_684,N_573,N_548);
nand U685 (N_685,N_556,N_505);
and U686 (N_686,N_504,N_559);
and U687 (N_687,N_505,N_598);
xnor U688 (N_688,N_549,N_534);
or U689 (N_689,N_538,N_521);
nor U690 (N_690,N_548,N_522);
nand U691 (N_691,N_516,N_571);
nand U692 (N_692,N_591,N_563);
nand U693 (N_693,N_531,N_539);
and U694 (N_694,N_567,N_597);
or U695 (N_695,N_587,N_553);
xor U696 (N_696,N_504,N_578);
nor U697 (N_697,N_556,N_530);
nand U698 (N_698,N_519,N_503);
nand U699 (N_699,N_576,N_529);
nand U700 (N_700,N_629,N_691);
nand U701 (N_701,N_679,N_607);
nor U702 (N_702,N_602,N_615);
and U703 (N_703,N_671,N_613);
nand U704 (N_704,N_648,N_653);
or U705 (N_705,N_689,N_684);
nand U706 (N_706,N_611,N_635);
nand U707 (N_707,N_654,N_634);
and U708 (N_708,N_670,N_668);
nand U709 (N_709,N_675,N_601);
or U710 (N_710,N_626,N_622);
xor U711 (N_711,N_688,N_612);
or U712 (N_712,N_683,N_680);
or U713 (N_713,N_604,N_621);
nor U714 (N_714,N_674,N_661);
nand U715 (N_715,N_678,N_644);
nor U716 (N_716,N_633,N_672);
and U717 (N_717,N_637,N_697);
or U718 (N_718,N_657,N_686);
nor U719 (N_719,N_610,N_656);
or U720 (N_720,N_681,N_642);
or U721 (N_721,N_650,N_699);
nor U722 (N_722,N_630,N_696);
or U723 (N_723,N_631,N_669);
nand U724 (N_724,N_690,N_645);
nor U725 (N_725,N_608,N_687);
xnor U726 (N_726,N_625,N_609);
xor U727 (N_727,N_659,N_618);
nor U728 (N_728,N_664,N_651);
or U729 (N_729,N_692,N_658);
xor U730 (N_730,N_603,N_655);
nor U731 (N_731,N_695,N_652);
nor U732 (N_732,N_649,N_663);
nor U733 (N_733,N_673,N_617);
xor U734 (N_734,N_639,N_676);
and U735 (N_735,N_665,N_600);
and U736 (N_736,N_698,N_666);
nor U737 (N_737,N_614,N_636);
or U738 (N_738,N_667,N_694);
nor U739 (N_739,N_624,N_619);
nand U740 (N_740,N_693,N_632);
or U741 (N_741,N_647,N_662);
and U742 (N_742,N_605,N_646);
nor U743 (N_743,N_623,N_643);
nand U744 (N_744,N_620,N_616);
or U745 (N_745,N_641,N_627);
or U746 (N_746,N_660,N_638);
or U747 (N_747,N_682,N_677);
nand U748 (N_748,N_685,N_628);
or U749 (N_749,N_640,N_606);
xor U750 (N_750,N_677,N_650);
nor U751 (N_751,N_609,N_666);
nor U752 (N_752,N_665,N_603);
and U753 (N_753,N_668,N_623);
and U754 (N_754,N_611,N_610);
nor U755 (N_755,N_688,N_625);
nor U756 (N_756,N_650,N_604);
or U757 (N_757,N_644,N_602);
nand U758 (N_758,N_670,N_671);
nor U759 (N_759,N_674,N_659);
and U760 (N_760,N_612,N_679);
and U761 (N_761,N_670,N_655);
nor U762 (N_762,N_689,N_624);
xor U763 (N_763,N_605,N_604);
nand U764 (N_764,N_610,N_663);
nor U765 (N_765,N_682,N_650);
or U766 (N_766,N_670,N_648);
or U767 (N_767,N_692,N_671);
or U768 (N_768,N_651,N_694);
or U769 (N_769,N_626,N_642);
nor U770 (N_770,N_685,N_648);
and U771 (N_771,N_695,N_624);
nand U772 (N_772,N_663,N_667);
or U773 (N_773,N_641,N_672);
and U774 (N_774,N_654,N_669);
nor U775 (N_775,N_690,N_607);
and U776 (N_776,N_686,N_667);
and U777 (N_777,N_669,N_634);
nor U778 (N_778,N_632,N_660);
nor U779 (N_779,N_634,N_689);
nor U780 (N_780,N_670,N_647);
nand U781 (N_781,N_604,N_623);
and U782 (N_782,N_680,N_690);
nand U783 (N_783,N_618,N_602);
and U784 (N_784,N_673,N_693);
nand U785 (N_785,N_654,N_693);
nor U786 (N_786,N_696,N_675);
xnor U787 (N_787,N_687,N_618);
and U788 (N_788,N_625,N_636);
nand U789 (N_789,N_627,N_685);
nor U790 (N_790,N_606,N_668);
and U791 (N_791,N_676,N_638);
nand U792 (N_792,N_633,N_622);
and U793 (N_793,N_672,N_685);
or U794 (N_794,N_634,N_681);
nor U795 (N_795,N_698,N_633);
or U796 (N_796,N_689,N_671);
nand U797 (N_797,N_667,N_680);
nor U798 (N_798,N_605,N_616);
nor U799 (N_799,N_670,N_689);
nand U800 (N_800,N_788,N_708);
or U801 (N_801,N_764,N_769);
nor U802 (N_802,N_796,N_710);
nand U803 (N_803,N_706,N_720);
nand U804 (N_804,N_768,N_721);
xor U805 (N_805,N_741,N_715);
or U806 (N_806,N_739,N_753);
nor U807 (N_807,N_732,N_789);
xor U808 (N_808,N_723,N_733);
nand U809 (N_809,N_709,N_773);
or U810 (N_810,N_762,N_747);
nand U811 (N_811,N_791,N_726);
nor U812 (N_812,N_783,N_750);
or U813 (N_813,N_765,N_734);
and U814 (N_814,N_775,N_763);
or U815 (N_815,N_751,N_759);
nor U816 (N_816,N_798,N_738);
or U817 (N_817,N_787,N_774);
or U818 (N_818,N_776,N_785);
nor U819 (N_819,N_758,N_746);
nand U820 (N_820,N_722,N_761);
nand U821 (N_821,N_729,N_737);
or U822 (N_822,N_711,N_767);
or U823 (N_823,N_730,N_755);
xor U824 (N_824,N_700,N_756);
and U825 (N_825,N_795,N_712);
or U826 (N_826,N_731,N_777);
or U827 (N_827,N_704,N_717);
or U828 (N_828,N_748,N_744);
nand U829 (N_829,N_772,N_782);
or U830 (N_830,N_779,N_760);
or U831 (N_831,N_740,N_794);
nand U832 (N_832,N_754,N_703);
or U833 (N_833,N_736,N_771);
and U834 (N_834,N_702,N_714);
or U835 (N_835,N_793,N_713);
and U836 (N_836,N_770,N_797);
nand U837 (N_837,N_799,N_743);
nand U838 (N_838,N_727,N_752);
or U839 (N_839,N_728,N_705);
or U840 (N_840,N_701,N_742);
xnor U841 (N_841,N_792,N_781);
nor U842 (N_842,N_735,N_790);
nand U843 (N_843,N_757,N_724);
nand U844 (N_844,N_718,N_780);
and U845 (N_845,N_707,N_745);
nor U846 (N_846,N_719,N_784);
nor U847 (N_847,N_716,N_725);
or U848 (N_848,N_786,N_766);
nand U849 (N_849,N_749,N_778);
or U850 (N_850,N_780,N_728);
or U851 (N_851,N_776,N_779);
or U852 (N_852,N_771,N_739);
and U853 (N_853,N_723,N_736);
nand U854 (N_854,N_742,N_781);
xnor U855 (N_855,N_774,N_720);
or U856 (N_856,N_713,N_738);
xor U857 (N_857,N_706,N_722);
nand U858 (N_858,N_758,N_729);
xnor U859 (N_859,N_775,N_774);
xnor U860 (N_860,N_707,N_779);
and U861 (N_861,N_778,N_754);
nand U862 (N_862,N_753,N_754);
or U863 (N_863,N_711,N_760);
nand U864 (N_864,N_764,N_773);
nor U865 (N_865,N_743,N_735);
nor U866 (N_866,N_765,N_790);
or U867 (N_867,N_762,N_700);
nor U868 (N_868,N_757,N_707);
or U869 (N_869,N_712,N_744);
or U870 (N_870,N_777,N_783);
and U871 (N_871,N_729,N_752);
or U872 (N_872,N_720,N_784);
nor U873 (N_873,N_792,N_766);
nor U874 (N_874,N_745,N_747);
and U875 (N_875,N_727,N_709);
xor U876 (N_876,N_731,N_745);
nand U877 (N_877,N_752,N_786);
or U878 (N_878,N_783,N_707);
and U879 (N_879,N_799,N_759);
or U880 (N_880,N_724,N_775);
nand U881 (N_881,N_751,N_778);
nor U882 (N_882,N_760,N_700);
xor U883 (N_883,N_797,N_752);
nor U884 (N_884,N_719,N_701);
or U885 (N_885,N_790,N_737);
and U886 (N_886,N_746,N_753);
and U887 (N_887,N_730,N_792);
and U888 (N_888,N_779,N_770);
xor U889 (N_889,N_734,N_776);
xnor U890 (N_890,N_705,N_746);
and U891 (N_891,N_722,N_750);
nand U892 (N_892,N_737,N_728);
and U893 (N_893,N_795,N_793);
nand U894 (N_894,N_770,N_757);
or U895 (N_895,N_726,N_735);
nand U896 (N_896,N_792,N_732);
nor U897 (N_897,N_734,N_709);
nand U898 (N_898,N_764,N_775);
nand U899 (N_899,N_792,N_785);
and U900 (N_900,N_886,N_848);
or U901 (N_901,N_835,N_803);
and U902 (N_902,N_895,N_821);
nand U903 (N_903,N_869,N_873);
nor U904 (N_904,N_825,N_832);
and U905 (N_905,N_871,N_884);
nor U906 (N_906,N_809,N_804);
xnor U907 (N_907,N_898,N_889);
nand U908 (N_908,N_813,N_875);
and U909 (N_909,N_823,N_838);
or U910 (N_910,N_807,N_841);
nor U911 (N_911,N_896,N_801);
nand U912 (N_912,N_874,N_893);
or U913 (N_913,N_858,N_888);
and U914 (N_914,N_877,N_855);
or U915 (N_915,N_817,N_826);
nand U916 (N_916,N_856,N_882);
nand U917 (N_917,N_881,N_846);
nand U918 (N_918,N_853,N_899);
nor U919 (N_919,N_843,N_819);
nor U920 (N_920,N_865,N_830);
or U921 (N_921,N_811,N_876);
nor U922 (N_922,N_879,N_851);
nand U923 (N_923,N_867,N_836);
or U924 (N_924,N_860,N_827);
nor U925 (N_925,N_828,N_862);
or U926 (N_926,N_878,N_822);
and U927 (N_927,N_872,N_837);
or U928 (N_928,N_844,N_842);
nor U929 (N_929,N_897,N_870);
and U930 (N_930,N_847,N_863);
or U931 (N_931,N_894,N_812);
nand U932 (N_932,N_820,N_891);
nor U933 (N_933,N_866,N_805);
and U934 (N_934,N_883,N_814);
or U935 (N_935,N_806,N_852);
or U936 (N_936,N_859,N_849);
or U937 (N_937,N_833,N_845);
and U938 (N_938,N_892,N_864);
or U939 (N_939,N_887,N_818);
nand U940 (N_940,N_816,N_824);
and U941 (N_941,N_857,N_868);
xor U942 (N_942,N_808,N_810);
nand U943 (N_943,N_890,N_839);
or U944 (N_944,N_854,N_861);
nand U945 (N_945,N_850,N_885);
and U946 (N_946,N_800,N_834);
nand U947 (N_947,N_880,N_829);
nand U948 (N_948,N_831,N_802);
nor U949 (N_949,N_840,N_815);
nand U950 (N_950,N_806,N_858);
nor U951 (N_951,N_878,N_855);
nor U952 (N_952,N_819,N_897);
nor U953 (N_953,N_815,N_813);
nand U954 (N_954,N_808,N_893);
xor U955 (N_955,N_869,N_883);
and U956 (N_956,N_863,N_822);
nand U957 (N_957,N_869,N_801);
nand U958 (N_958,N_845,N_860);
nand U959 (N_959,N_823,N_875);
and U960 (N_960,N_883,N_874);
and U961 (N_961,N_828,N_818);
and U962 (N_962,N_805,N_807);
and U963 (N_963,N_832,N_859);
nand U964 (N_964,N_853,N_836);
nor U965 (N_965,N_881,N_847);
nand U966 (N_966,N_817,N_899);
nand U967 (N_967,N_898,N_823);
or U968 (N_968,N_844,N_878);
nor U969 (N_969,N_887,N_831);
xnor U970 (N_970,N_869,N_805);
or U971 (N_971,N_803,N_841);
or U972 (N_972,N_839,N_868);
nand U973 (N_973,N_888,N_897);
or U974 (N_974,N_883,N_838);
and U975 (N_975,N_806,N_859);
or U976 (N_976,N_831,N_881);
nor U977 (N_977,N_849,N_833);
and U978 (N_978,N_875,N_889);
nor U979 (N_979,N_814,N_864);
nand U980 (N_980,N_862,N_879);
nor U981 (N_981,N_875,N_800);
nor U982 (N_982,N_859,N_851);
nand U983 (N_983,N_873,N_851);
nand U984 (N_984,N_811,N_861);
and U985 (N_985,N_863,N_816);
or U986 (N_986,N_811,N_828);
xor U987 (N_987,N_801,N_860);
nor U988 (N_988,N_874,N_895);
or U989 (N_989,N_889,N_854);
xnor U990 (N_990,N_813,N_850);
and U991 (N_991,N_862,N_805);
nor U992 (N_992,N_862,N_873);
and U993 (N_993,N_812,N_863);
xnor U994 (N_994,N_846,N_894);
or U995 (N_995,N_876,N_835);
or U996 (N_996,N_808,N_852);
nand U997 (N_997,N_820,N_813);
and U998 (N_998,N_853,N_866);
or U999 (N_999,N_804,N_887);
or U1000 (N_1000,N_996,N_900);
nor U1001 (N_1001,N_903,N_954);
nand U1002 (N_1002,N_978,N_918);
and U1003 (N_1003,N_985,N_979);
xor U1004 (N_1004,N_955,N_916);
xor U1005 (N_1005,N_910,N_959);
or U1006 (N_1006,N_957,N_975);
nor U1007 (N_1007,N_971,N_968);
nor U1008 (N_1008,N_961,N_924);
and U1009 (N_1009,N_904,N_913);
nand U1010 (N_1010,N_911,N_983);
nand U1011 (N_1011,N_984,N_938);
nand U1012 (N_1012,N_993,N_952);
nor U1013 (N_1013,N_970,N_998);
and U1014 (N_1014,N_986,N_927);
nor U1015 (N_1015,N_974,N_966);
nand U1016 (N_1016,N_973,N_935);
xnor U1017 (N_1017,N_944,N_997);
and U1018 (N_1018,N_914,N_969);
and U1019 (N_1019,N_992,N_990);
xnor U1020 (N_1020,N_980,N_922);
or U1021 (N_1021,N_951,N_994);
nor U1022 (N_1022,N_923,N_962);
nand U1023 (N_1023,N_929,N_930);
nand U1024 (N_1024,N_921,N_981);
nand U1025 (N_1025,N_917,N_989);
xnor U1026 (N_1026,N_939,N_912);
nand U1027 (N_1027,N_909,N_931);
nor U1028 (N_1028,N_934,N_919);
xor U1029 (N_1029,N_995,N_947);
nand U1030 (N_1030,N_991,N_976);
nor U1031 (N_1031,N_977,N_982);
and U1032 (N_1032,N_928,N_965);
xnor U1033 (N_1033,N_907,N_925);
nand U1034 (N_1034,N_963,N_972);
or U1035 (N_1035,N_901,N_940);
nor U1036 (N_1036,N_946,N_942);
nor U1037 (N_1037,N_964,N_906);
or U1038 (N_1038,N_902,N_960);
nand U1039 (N_1039,N_945,N_988);
nand U1040 (N_1040,N_933,N_948);
nand U1041 (N_1041,N_905,N_915);
xor U1042 (N_1042,N_950,N_920);
or U1043 (N_1043,N_936,N_999);
nand U1044 (N_1044,N_953,N_949);
or U1045 (N_1045,N_967,N_908);
nor U1046 (N_1046,N_941,N_956);
nand U1047 (N_1047,N_958,N_932);
nor U1048 (N_1048,N_937,N_926);
nor U1049 (N_1049,N_987,N_943);
or U1050 (N_1050,N_971,N_992);
xor U1051 (N_1051,N_922,N_926);
nor U1052 (N_1052,N_938,N_942);
and U1053 (N_1053,N_984,N_997);
nand U1054 (N_1054,N_948,N_984);
nor U1055 (N_1055,N_938,N_963);
and U1056 (N_1056,N_953,N_996);
nor U1057 (N_1057,N_923,N_989);
or U1058 (N_1058,N_962,N_909);
nand U1059 (N_1059,N_923,N_901);
nand U1060 (N_1060,N_919,N_969);
or U1061 (N_1061,N_991,N_989);
nor U1062 (N_1062,N_935,N_957);
or U1063 (N_1063,N_957,N_991);
nand U1064 (N_1064,N_972,N_932);
and U1065 (N_1065,N_927,N_979);
nor U1066 (N_1066,N_925,N_982);
nor U1067 (N_1067,N_903,N_971);
or U1068 (N_1068,N_938,N_901);
or U1069 (N_1069,N_925,N_943);
nor U1070 (N_1070,N_983,N_967);
nor U1071 (N_1071,N_989,N_941);
or U1072 (N_1072,N_958,N_910);
xor U1073 (N_1073,N_928,N_978);
and U1074 (N_1074,N_918,N_992);
or U1075 (N_1075,N_906,N_910);
nand U1076 (N_1076,N_930,N_952);
or U1077 (N_1077,N_932,N_926);
nand U1078 (N_1078,N_906,N_905);
or U1079 (N_1079,N_968,N_900);
or U1080 (N_1080,N_943,N_970);
or U1081 (N_1081,N_943,N_938);
nor U1082 (N_1082,N_928,N_911);
nor U1083 (N_1083,N_921,N_958);
and U1084 (N_1084,N_967,N_978);
or U1085 (N_1085,N_975,N_950);
or U1086 (N_1086,N_979,N_971);
nand U1087 (N_1087,N_995,N_915);
and U1088 (N_1088,N_986,N_926);
nand U1089 (N_1089,N_960,N_937);
or U1090 (N_1090,N_967,N_975);
or U1091 (N_1091,N_906,N_900);
xor U1092 (N_1092,N_986,N_905);
and U1093 (N_1093,N_907,N_910);
nor U1094 (N_1094,N_967,N_971);
nor U1095 (N_1095,N_900,N_936);
nand U1096 (N_1096,N_909,N_968);
nor U1097 (N_1097,N_983,N_938);
and U1098 (N_1098,N_924,N_933);
nor U1099 (N_1099,N_961,N_975);
nand U1100 (N_1100,N_1027,N_1002);
and U1101 (N_1101,N_1035,N_1092);
nand U1102 (N_1102,N_1028,N_1080);
and U1103 (N_1103,N_1090,N_1094);
and U1104 (N_1104,N_1099,N_1054);
nand U1105 (N_1105,N_1072,N_1087);
or U1106 (N_1106,N_1075,N_1019);
and U1107 (N_1107,N_1040,N_1030);
and U1108 (N_1108,N_1073,N_1005);
xnor U1109 (N_1109,N_1031,N_1007);
nand U1110 (N_1110,N_1064,N_1025);
nand U1111 (N_1111,N_1061,N_1088);
nor U1112 (N_1112,N_1041,N_1017);
nor U1113 (N_1113,N_1009,N_1071);
xnor U1114 (N_1114,N_1068,N_1023);
nor U1115 (N_1115,N_1086,N_1037);
or U1116 (N_1116,N_1096,N_1039);
nor U1117 (N_1117,N_1059,N_1015);
xnor U1118 (N_1118,N_1000,N_1042);
nor U1119 (N_1119,N_1006,N_1029);
or U1120 (N_1120,N_1052,N_1018);
or U1121 (N_1121,N_1003,N_1022);
nor U1122 (N_1122,N_1008,N_1043);
nand U1123 (N_1123,N_1026,N_1091);
xor U1124 (N_1124,N_1069,N_1014);
xnor U1125 (N_1125,N_1077,N_1057);
xnor U1126 (N_1126,N_1033,N_1060);
or U1127 (N_1127,N_1047,N_1066);
nand U1128 (N_1128,N_1001,N_1024);
or U1129 (N_1129,N_1046,N_1038);
xnor U1130 (N_1130,N_1032,N_1016);
or U1131 (N_1131,N_1085,N_1067);
xnor U1132 (N_1132,N_1034,N_1062);
nor U1133 (N_1133,N_1011,N_1055);
nor U1134 (N_1134,N_1012,N_1053);
nand U1135 (N_1135,N_1049,N_1058);
and U1136 (N_1136,N_1051,N_1097);
nand U1137 (N_1137,N_1070,N_1044);
nand U1138 (N_1138,N_1056,N_1045);
nand U1139 (N_1139,N_1076,N_1048);
nand U1140 (N_1140,N_1084,N_1063);
nand U1141 (N_1141,N_1010,N_1089);
nand U1142 (N_1142,N_1093,N_1078);
nand U1143 (N_1143,N_1083,N_1021);
nand U1144 (N_1144,N_1020,N_1095);
nand U1145 (N_1145,N_1013,N_1065);
and U1146 (N_1146,N_1079,N_1098);
xor U1147 (N_1147,N_1036,N_1081);
nand U1148 (N_1148,N_1050,N_1004);
or U1149 (N_1149,N_1074,N_1082);
or U1150 (N_1150,N_1042,N_1012);
nor U1151 (N_1151,N_1075,N_1090);
or U1152 (N_1152,N_1089,N_1056);
nor U1153 (N_1153,N_1077,N_1050);
nor U1154 (N_1154,N_1061,N_1032);
and U1155 (N_1155,N_1058,N_1073);
xor U1156 (N_1156,N_1091,N_1078);
or U1157 (N_1157,N_1014,N_1098);
or U1158 (N_1158,N_1073,N_1081);
xnor U1159 (N_1159,N_1067,N_1010);
and U1160 (N_1160,N_1014,N_1082);
and U1161 (N_1161,N_1028,N_1008);
nor U1162 (N_1162,N_1064,N_1063);
nand U1163 (N_1163,N_1015,N_1062);
nand U1164 (N_1164,N_1079,N_1096);
and U1165 (N_1165,N_1007,N_1005);
and U1166 (N_1166,N_1028,N_1020);
or U1167 (N_1167,N_1066,N_1007);
nand U1168 (N_1168,N_1031,N_1043);
nor U1169 (N_1169,N_1063,N_1002);
nand U1170 (N_1170,N_1020,N_1078);
or U1171 (N_1171,N_1064,N_1001);
nor U1172 (N_1172,N_1053,N_1065);
and U1173 (N_1173,N_1091,N_1024);
nand U1174 (N_1174,N_1097,N_1056);
nand U1175 (N_1175,N_1008,N_1092);
nor U1176 (N_1176,N_1018,N_1025);
xor U1177 (N_1177,N_1083,N_1017);
and U1178 (N_1178,N_1052,N_1033);
and U1179 (N_1179,N_1056,N_1077);
xnor U1180 (N_1180,N_1082,N_1040);
nand U1181 (N_1181,N_1016,N_1073);
and U1182 (N_1182,N_1085,N_1046);
nor U1183 (N_1183,N_1023,N_1026);
xor U1184 (N_1184,N_1073,N_1010);
nor U1185 (N_1185,N_1012,N_1050);
nor U1186 (N_1186,N_1069,N_1044);
xnor U1187 (N_1187,N_1088,N_1082);
nor U1188 (N_1188,N_1045,N_1041);
and U1189 (N_1189,N_1053,N_1055);
nor U1190 (N_1190,N_1059,N_1027);
and U1191 (N_1191,N_1037,N_1098);
nor U1192 (N_1192,N_1068,N_1004);
and U1193 (N_1193,N_1036,N_1023);
or U1194 (N_1194,N_1029,N_1017);
and U1195 (N_1195,N_1049,N_1031);
xnor U1196 (N_1196,N_1074,N_1016);
or U1197 (N_1197,N_1020,N_1026);
nor U1198 (N_1198,N_1054,N_1039);
xnor U1199 (N_1199,N_1087,N_1097);
or U1200 (N_1200,N_1193,N_1113);
nor U1201 (N_1201,N_1146,N_1116);
and U1202 (N_1202,N_1103,N_1130);
xor U1203 (N_1203,N_1133,N_1104);
nand U1204 (N_1204,N_1157,N_1166);
nand U1205 (N_1205,N_1100,N_1131);
nand U1206 (N_1206,N_1141,N_1192);
xor U1207 (N_1207,N_1152,N_1196);
nand U1208 (N_1208,N_1136,N_1129);
nand U1209 (N_1209,N_1162,N_1165);
and U1210 (N_1210,N_1160,N_1138);
nor U1211 (N_1211,N_1188,N_1110);
or U1212 (N_1212,N_1198,N_1164);
and U1213 (N_1213,N_1148,N_1153);
and U1214 (N_1214,N_1173,N_1119);
nand U1215 (N_1215,N_1174,N_1191);
nand U1216 (N_1216,N_1183,N_1195);
and U1217 (N_1217,N_1142,N_1144);
and U1218 (N_1218,N_1186,N_1135);
xnor U1219 (N_1219,N_1108,N_1132);
nor U1220 (N_1220,N_1159,N_1125);
xnor U1221 (N_1221,N_1149,N_1163);
or U1222 (N_1222,N_1158,N_1189);
or U1223 (N_1223,N_1126,N_1105);
nand U1224 (N_1224,N_1150,N_1147);
and U1225 (N_1225,N_1155,N_1184);
nor U1226 (N_1226,N_1115,N_1176);
and U1227 (N_1227,N_1154,N_1127);
nand U1228 (N_1228,N_1102,N_1109);
nor U1229 (N_1229,N_1167,N_1194);
nor U1230 (N_1230,N_1134,N_1177);
nand U1231 (N_1231,N_1118,N_1145);
or U1232 (N_1232,N_1107,N_1190);
nor U1233 (N_1233,N_1143,N_1171);
or U1234 (N_1234,N_1197,N_1114);
or U1235 (N_1235,N_1128,N_1178);
and U1236 (N_1236,N_1151,N_1106);
xor U1237 (N_1237,N_1179,N_1101);
or U1238 (N_1238,N_1180,N_1137);
nand U1239 (N_1239,N_1140,N_1161);
and U1240 (N_1240,N_1139,N_1187);
or U1241 (N_1241,N_1123,N_1168);
nor U1242 (N_1242,N_1182,N_1169);
and U1243 (N_1243,N_1175,N_1124);
and U1244 (N_1244,N_1170,N_1181);
nand U1245 (N_1245,N_1120,N_1122);
nor U1246 (N_1246,N_1111,N_1112);
or U1247 (N_1247,N_1172,N_1156);
or U1248 (N_1248,N_1121,N_1185);
nand U1249 (N_1249,N_1117,N_1199);
nor U1250 (N_1250,N_1101,N_1129);
xnor U1251 (N_1251,N_1143,N_1142);
and U1252 (N_1252,N_1199,N_1162);
nor U1253 (N_1253,N_1172,N_1151);
nand U1254 (N_1254,N_1173,N_1185);
or U1255 (N_1255,N_1186,N_1123);
or U1256 (N_1256,N_1117,N_1146);
or U1257 (N_1257,N_1108,N_1106);
xor U1258 (N_1258,N_1176,N_1180);
nor U1259 (N_1259,N_1148,N_1161);
nand U1260 (N_1260,N_1110,N_1163);
and U1261 (N_1261,N_1164,N_1101);
and U1262 (N_1262,N_1185,N_1115);
nand U1263 (N_1263,N_1152,N_1110);
or U1264 (N_1264,N_1189,N_1168);
nand U1265 (N_1265,N_1129,N_1118);
nand U1266 (N_1266,N_1165,N_1179);
or U1267 (N_1267,N_1199,N_1178);
and U1268 (N_1268,N_1124,N_1166);
or U1269 (N_1269,N_1122,N_1170);
xor U1270 (N_1270,N_1195,N_1188);
nand U1271 (N_1271,N_1162,N_1154);
nand U1272 (N_1272,N_1181,N_1128);
and U1273 (N_1273,N_1198,N_1111);
or U1274 (N_1274,N_1108,N_1184);
or U1275 (N_1275,N_1103,N_1148);
nand U1276 (N_1276,N_1187,N_1115);
nor U1277 (N_1277,N_1163,N_1108);
and U1278 (N_1278,N_1102,N_1114);
nand U1279 (N_1279,N_1127,N_1120);
xor U1280 (N_1280,N_1149,N_1196);
and U1281 (N_1281,N_1177,N_1152);
nand U1282 (N_1282,N_1122,N_1160);
and U1283 (N_1283,N_1103,N_1193);
nand U1284 (N_1284,N_1125,N_1165);
xnor U1285 (N_1285,N_1129,N_1134);
nor U1286 (N_1286,N_1186,N_1196);
or U1287 (N_1287,N_1176,N_1161);
and U1288 (N_1288,N_1183,N_1124);
xnor U1289 (N_1289,N_1104,N_1189);
nand U1290 (N_1290,N_1154,N_1116);
nand U1291 (N_1291,N_1108,N_1181);
and U1292 (N_1292,N_1117,N_1197);
nand U1293 (N_1293,N_1197,N_1123);
xor U1294 (N_1294,N_1154,N_1182);
xnor U1295 (N_1295,N_1117,N_1192);
nor U1296 (N_1296,N_1194,N_1153);
and U1297 (N_1297,N_1165,N_1138);
and U1298 (N_1298,N_1190,N_1125);
nand U1299 (N_1299,N_1117,N_1156);
and U1300 (N_1300,N_1231,N_1291);
nor U1301 (N_1301,N_1240,N_1262);
nor U1302 (N_1302,N_1247,N_1290);
nor U1303 (N_1303,N_1203,N_1243);
or U1304 (N_1304,N_1229,N_1285);
and U1305 (N_1305,N_1225,N_1268);
nor U1306 (N_1306,N_1296,N_1213);
nor U1307 (N_1307,N_1219,N_1207);
or U1308 (N_1308,N_1298,N_1275);
and U1309 (N_1309,N_1277,N_1235);
nand U1310 (N_1310,N_1221,N_1270);
and U1311 (N_1311,N_1214,N_1281);
nor U1312 (N_1312,N_1236,N_1256);
and U1313 (N_1313,N_1228,N_1211);
nor U1314 (N_1314,N_1241,N_1254);
or U1315 (N_1315,N_1226,N_1222);
nor U1316 (N_1316,N_1255,N_1295);
or U1317 (N_1317,N_1279,N_1218);
and U1318 (N_1318,N_1234,N_1215);
nand U1319 (N_1319,N_1259,N_1249);
nand U1320 (N_1320,N_1284,N_1257);
nor U1321 (N_1321,N_1239,N_1200);
and U1322 (N_1322,N_1299,N_1250);
and U1323 (N_1323,N_1245,N_1253);
and U1324 (N_1324,N_1283,N_1274);
and U1325 (N_1325,N_1280,N_1244);
and U1326 (N_1326,N_1265,N_1264);
or U1327 (N_1327,N_1209,N_1205);
and U1328 (N_1328,N_1278,N_1204);
or U1329 (N_1329,N_1282,N_1272);
nor U1330 (N_1330,N_1230,N_1217);
and U1331 (N_1331,N_1267,N_1201);
nor U1332 (N_1332,N_1227,N_1206);
nand U1333 (N_1333,N_1276,N_1233);
nand U1334 (N_1334,N_1242,N_1289);
nor U1335 (N_1335,N_1293,N_1224);
nand U1336 (N_1336,N_1288,N_1246);
xor U1337 (N_1337,N_1202,N_1220);
and U1338 (N_1338,N_1212,N_1223);
or U1339 (N_1339,N_1273,N_1261);
and U1340 (N_1340,N_1251,N_1208);
nand U1341 (N_1341,N_1258,N_1269);
xnor U1342 (N_1342,N_1292,N_1297);
and U1343 (N_1343,N_1232,N_1210);
nor U1344 (N_1344,N_1287,N_1294);
or U1345 (N_1345,N_1260,N_1271);
nor U1346 (N_1346,N_1216,N_1252);
nor U1347 (N_1347,N_1238,N_1286);
or U1348 (N_1348,N_1237,N_1248);
or U1349 (N_1349,N_1266,N_1263);
nand U1350 (N_1350,N_1270,N_1287);
or U1351 (N_1351,N_1240,N_1292);
and U1352 (N_1352,N_1264,N_1237);
and U1353 (N_1353,N_1246,N_1268);
nor U1354 (N_1354,N_1257,N_1291);
and U1355 (N_1355,N_1228,N_1296);
nand U1356 (N_1356,N_1227,N_1294);
and U1357 (N_1357,N_1287,N_1256);
nand U1358 (N_1358,N_1222,N_1240);
xnor U1359 (N_1359,N_1231,N_1281);
or U1360 (N_1360,N_1250,N_1253);
xor U1361 (N_1361,N_1278,N_1256);
and U1362 (N_1362,N_1223,N_1280);
or U1363 (N_1363,N_1242,N_1286);
and U1364 (N_1364,N_1216,N_1291);
or U1365 (N_1365,N_1294,N_1299);
or U1366 (N_1366,N_1245,N_1209);
nand U1367 (N_1367,N_1211,N_1235);
nor U1368 (N_1368,N_1254,N_1244);
nor U1369 (N_1369,N_1271,N_1252);
xor U1370 (N_1370,N_1236,N_1258);
nor U1371 (N_1371,N_1236,N_1294);
or U1372 (N_1372,N_1257,N_1212);
or U1373 (N_1373,N_1272,N_1214);
nand U1374 (N_1374,N_1277,N_1222);
nor U1375 (N_1375,N_1219,N_1200);
and U1376 (N_1376,N_1222,N_1272);
and U1377 (N_1377,N_1258,N_1251);
xor U1378 (N_1378,N_1217,N_1299);
xor U1379 (N_1379,N_1273,N_1244);
nor U1380 (N_1380,N_1275,N_1272);
and U1381 (N_1381,N_1274,N_1204);
and U1382 (N_1382,N_1206,N_1273);
or U1383 (N_1383,N_1203,N_1262);
and U1384 (N_1384,N_1289,N_1287);
xnor U1385 (N_1385,N_1275,N_1232);
and U1386 (N_1386,N_1227,N_1261);
or U1387 (N_1387,N_1235,N_1296);
nand U1388 (N_1388,N_1266,N_1293);
nand U1389 (N_1389,N_1260,N_1235);
or U1390 (N_1390,N_1238,N_1201);
or U1391 (N_1391,N_1219,N_1209);
nor U1392 (N_1392,N_1255,N_1251);
or U1393 (N_1393,N_1233,N_1238);
xor U1394 (N_1394,N_1264,N_1292);
nor U1395 (N_1395,N_1228,N_1279);
or U1396 (N_1396,N_1262,N_1269);
nand U1397 (N_1397,N_1224,N_1251);
and U1398 (N_1398,N_1213,N_1240);
or U1399 (N_1399,N_1285,N_1246);
nand U1400 (N_1400,N_1324,N_1305);
nor U1401 (N_1401,N_1376,N_1389);
nand U1402 (N_1402,N_1353,N_1307);
or U1403 (N_1403,N_1335,N_1343);
and U1404 (N_1404,N_1361,N_1345);
nand U1405 (N_1405,N_1312,N_1366);
and U1406 (N_1406,N_1330,N_1338);
nand U1407 (N_1407,N_1357,N_1381);
nand U1408 (N_1408,N_1315,N_1304);
or U1409 (N_1409,N_1308,N_1314);
and U1410 (N_1410,N_1311,N_1367);
nand U1411 (N_1411,N_1309,N_1369);
and U1412 (N_1412,N_1346,N_1347);
and U1413 (N_1413,N_1378,N_1337);
nand U1414 (N_1414,N_1328,N_1374);
or U1415 (N_1415,N_1306,N_1386);
or U1416 (N_1416,N_1331,N_1349);
nor U1417 (N_1417,N_1388,N_1332);
nor U1418 (N_1418,N_1360,N_1380);
nand U1419 (N_1419,N_1375,N_1333);
and U1420 (N_1420,N_1336,N_1363);
or U1421 (N_1421,N_1316,N_1302);
nor U1422 (N_1422,N_1390,N_1303);
xnor U1423 (N_1423,N_1320,N_1364);
and U1424 (N_1424,N_1319,N_1365);
xnor U1425 (N_1425,N_1354,N_1370);
and U1426 (N_1426,N_1323,N_1395);
or U1427 (N_1427,N_1396,N_1377);
nor U1428 (N_1428,N_1313,N_1341);
nand U1429 (N_1429,N_1379,N_1385);
xor U1430 (N_1430,N_1356,N_1384);
xnor U1431 (N_1431,N_1317,N_1326);
or U1432 (N_1432,N_1362,N_1399);
or U1433 (N_1433,N_1321,N_1334);
nor U1434 (N_1434,N_1359,N_1351);
nor U1435 (N_1435,N_1352,N_1325);
nand U1436 (N_1436,N_1329,N_1398);
nand U1437 (N_1437,N_1397,N_1391);
nand U1438 (N_1438,N_1383,N_1371);
and U1439 (N_1439,N_1340,N_1300);
and U1440 (N_1440,N_1382,N_1387);
xnor U1441 (N_1441,N_1327,N_1348);
and U1442 (N_1442,N_1344,N_1372);
and U1443 (N_1443,N_1358,N_1355);
and U1444 (N_1444,N_1339,N_1392);
nand U1445 (N_1445,N_1301,N_1322);
xor U1446 (N_1446,N_1350,N_1393);
xor U1447 (N_1447,N_1310,N_1373);
xnor U1448 (N_1448,N_1318,N_1368);
nand U1449 (N_1449,N_1342,N_1394);
nand U1450 (N_1450,N_1385,N_1315);
nor U1451 (N_1451,N_1344,N_1351);
nor U1452 (N_1452,N_1331,N_1361);
and U1453 (N_1453,N_1301,N_1377);
nor U1454 (N_1454,N_1349,N_1376);
or U1455 (N_1455,N_1375,N_1313);
nand U1456 (N_1456,N_1352,N_1391);
and U1457 (N_1457,N_1318,N_1374);
and U1458 (N_1458,N_1353,N_1345);
and U1459 (N_1459,N_1317,N_1337);
nand U1460 (N_1460,N_1304,N_1394);
and U1461 (N_1461,N_1337,N_1397);
or U1462 (N_1462,N_1311,N_1397);
and U1463 (N_1463,N_1330,N_1321);
nor U1464 (N_1464,N_1364,N_1300);
nor U1465 (N_1465,N_1303,N_1301);
nand U1466 (N_1466,N_1329,N_1381);
or U1467 (N_1467,N_1348,N_1388);
nand U1468 (N_1468,N_1365,N_1324);
and U1469 (N_1469,N_1369,N_1362);
and U1470 (N_1470,N_1379,N_1328);
nand U1471 (N_1471,N_1326,N_1344);
and U1472 (N_1472,N_1391,N_1376);
xnor U1473 (N_1473,N_1322,N_1334);
and U1474 (N_1474,N_1378,N_1367);
and U1475 (N_1475,N_1351,N_1317);
and U1476 (N_1476,N_1319,N_1353);
and U1477 (N_1477,N_1316,N_1308);
xor U1478 (N_1478,N_1316,N_1360);
nor U1479 (N_1479,N_1354,N_1363);
and U1480 (N_1480,N_1369,N_1325);
nor U1481 (N_1481,N_1351,N_1357);
nor U1482 (N_1482,N_1326,N_1371);
xnor U1483 (N_1483,N_1342,N_1329);
nand U1484 (N_1484,N_1382,N_1319);
or U1485 (N_1485,N_1307,N_1319);
and U1486 (N_1486,N_1303,N_1321);
nor U1487 (N_1487,N_1306,N_1350);
nand U1488 (N_1488,N_1379,N_1318);
and U1489 (N_1489,N_1313,N_1348);
or U1490 (N_1490,N_1389,N_1364);
and U1491 (N_1491,N_1312,N_1339);
nand U1492 (N_1492,N_1323,N_1353);
nand U1493 (N_1493,N_1317,N_1373);
nand U1494 (N_1494,N_1338,N_1393);
or U1495 (N_1495,N_1378,N_1374);
nand U1496 (N_1496,N_1393,N_1342);
nor U1497 (N_1497,N_1357,N_1356);
and U1498 (N_1498,N_1300,N_1351);
nand U1499 (N_1499,N_1310,N_1341);
or U1500 (N_1500,N_1441,N_1428);
and U1501 (N_1501,N_1449,N_1487);
nor U1502 (N_1502,N_1413,N_1494);
nor U1503 (N_1503,N_1453,N_1433);
and U1504 (N_1504,N_1430,N_1470);
or U1505 (N_1505,N_1419,N_1451);
and U1506 (N_1506,N_1468,N_1416);
nor U1507 (N_1507,N_1417,N_1415);
xnor U1508 (N_1508,N_1426,N_1401);
nand U1509 (N_1509,N_1469,N_1499);
nand U1510 (N_1510,N_1485,N_1407);
nor U1511 (N_1511,N_1400,N_1475);
or U1512 (N_1512,N_1405,N_1412);
and U1513 (N_1513,N_1489,N_1488);
nand U1514 (N_1514,N_1444,N_1458);
xor U1515 (N_1515,N_1457,N_1491);
xor U1516 (N_1516,N_1402,N_1464);
nor U1517 (N_1517,N_1425,N_1498);
and U1518 (N_1518,N_1493,N_1438);
nand U1519 (N_1519,N_1482,N_1445);
or U1520 (N_1520,N_1462,N_1456);
nor U1521 (N_1521,N_1459,N_1414);
or U1522 (N_1522,N_1474,N_1461);
and U1523 (N_1523,N_1406,N_1479);
nor U1524 (N_1524,N_1421,N_1477);
or U1525 (N_1525,N_1427,N_1447);
or U1526 (N_1526,N_1439,N_1423);
or U1527 (N_1527,N_1431,N_1435);
nor U1528 (N_1528,N_1455,N_1409);
nand U1529 (N_1529,N_1429,N_1496);
nor U1530 (N_1530,N_1448,N_1437);
nor U1531 (N_1531,N_1446,N_1436);
or U1532 (N_1532,N_1484,N_1483);
or U1533 (N_1533,N_1478,N_1418);
nand U1534 (N_1534,N_1410,N_1404);
nand U1535 (N_1535,N_1442,N_1466);
nand U1536 (N_1536,N_1424,N_1473);
or U1537 (N_1537,N_1480,N_1432);
nand U1538 (N_1538,N_1490,N_1408);
nand U1539 (N_1539,N_1497,N_1403);
xor U1540 (N_1540,N_1411,N_1434);
or U1541 (N_1541,N_1495,N_1476);
or U1542 (N_1542,N_1471,N_1472);
and U1543 (N_1543,N_1440,N_1481);
nor U1544 (N_1544,N_1492,N_1460);
or U1545 (N_1545,N_1422,N_1443);
nand U1546 (N_1546,N_1465,N_1486);
nand U1547 (N_1547,N_1454,N_1467);
xor U1548 (N_1548,N_1452,N_1450);
nor U1549 (N_1549,N_1463,N_1420);
nor U1550 (N_1550,N_1473,N_1413);
or U1551 (N_1551,N_1489,N_1433);
nand U1552 (N_1552,N_1436,N_1423);
or U1553 (N_1553,N_1403,N_1492);
nor U1554 (N_1554,N_1451,N_1408);
nor U1555 (N_1555,N_1433,N_1444);
and U1556 (N_1556,N_1464,N_1433);
and U1557 (N_1557,N_1453,N_1428);
and U1558 (N_1558,N_1408,N_1420);
or U1559 (N_1559,N_1452,N_1444);
or U1560 (N_1560,N_1450,N_1481);
or U1561 (N_1561,N_1411,N_1488);
nand U1562 (N_1562,N_1423,N_1401);
nand U1563 (N_1563,N_1411,N_1499);
and U1564 (N_1564,N_1420,N_1431);
nor U1565 (N_1565,N_1452,N_1415);
xor U1566 (N_1566,N_1400,N_1473);
nor U1567 (N_1567,N_1456,N_1428);
or U1568 (N_1568,N_1431,N_1464);
nor U1569 (N_1569,N_1402,N_1455);
or U1570 (N_1570,N_1400,N_1409);
or U1571 (N_1571,N_1406,N_1477);
or U1572 (N_1572,N_1408,N_1464);
nand U1573 (N_1573,N_1487,N_1437);
or U1574 (N_1574,N_1498,N_1434);
nor U1575 (N_1575,N_1466,N_1478);
and U1576 (N_1576,N_1483,N_1499);
or U1577 (N_1577,N_1478,N_1438);
nor U1578 (N_1578,N_1414,N_1438);
and U1579 (N_1579,N_1452,N_1463);
nor U1580 (N_1580,N_1484,N_1492);
or U1581 (N_1581,N_1459,N_1403);
or U1582 (N_1582,N_1437,N_1480);
or U1583 (N_1583,N_1409,N_1467);
nor U1584 (N_1584,N_1490,N_1448);
nand U1585 (N_1585,N_1471,N_1489);
and U1586 (N_1586,N_1475,N_1443);
or U1587 (N_1587,N_1410,N_1492);
and U1588 (N_1588,N_1432,N_1455);
and U1589 (N_1589,N_1421,N_1464);
nor U1590 (N_1590,N_1479,N_1480);
xnor U1591 (N_1591,N_1475,N_1457);
nand U1592 (N_1592,N_1406,N_1443);
nor U1593 (N_1593,N_1430,N_1445);
xnor U1594 (N_1594,N_1484,N_1493);
nor U1595 (N_1595,N_1493,N_1423);
nand U1596 (N_1596,N_1435,N_1481);
nand U1597 (N_1597,N_1446,N_1480);
or U1598 (N_1598,N_1417,N_1425);
xnor U1599 (N_1599,N_1497,N_1488);
and U1600 (N_1600,N_1546,N_1586);
and U1601 (N_1601,N_1547,N_1570);
and U1602 (N_1602,N_1598,N_1560);
nor U1603 (N_1603,N_1561,N_1568);
nor U1604 (N_1604,N_1514,N_1507);
nand U1605 (N_1605,N_1573,N_1524);
nor U1606 (N_1606,N_1530,N_1505);
nand U1607 (N_1607,N_1563,N_1516);
or U1608 (N_1608,N_1535,N_1562);
nor U1609 (N_1609,N_1582,N_1525);
nor U1610 (N_1610,N_1571,N_1567);
nand U1611 (N_1611,N_1528,N_1579);
or U1612 (N_1612,N_1503,N_1520);
and U1613 (N_1613,N_1554,N_1513);
xnor U1614 (N_1614,N_1550,N_1555);
nand U1615 (N_1615,N_1595,N_1572);
and U1616 (N_1616,N_1578,N_1545);
and U1617 (N_1617,N_1588,N_1575);
or U1618 (N_1618,N_1511,N_1536);
and U1619 (N_1619,N_1527,N_1506);
xnor U1620 (N_1620,N_1534,N_1540);
and U1621 (N_1621,N_1591,N_1538);
and U1622 (N_1622,N_1577,N_1504);
nor U1623 (N_1623,N_1502,N_1517);
and U1624 (N_1624,N_1529,N_1576);
xor U1625 (N_1625,N_1549,N_1596);
or U1626 (N_1626,N_1592,N_1539);
nor U1627 (N_1627,N_1597,N_1522);
nand U1628 (N_1628,N_1594,N_1564);
and U1629 (N_1629,N_1510,N_1551);
xor U1630 (N_1630,N_1565,N_1569);
and U1631 (N_1631,N_1593,N_1553);
and U1632 (N_1632,N_1584,N_1501);
or U1633 (N_1633,N_1526,N_1533);
and U1634 (N_1634,N_1581,N_1541);
or U1635 (N_1635,N_1589,N_1580);
or U1636 (N_1636,N_1585,N_1587);
or U1637 (N_1637,N_1552,N_1508);
nand U1638 (N_1638,N_1544,N_1599);
or U1639 (N_1639,N_1512,N_1557);
or U1640 (N_1640,N_1574,N_1518);
or U1641 (N_1641,N_1543,N_1559);
xor U1642 (N_1642,N_1531,N_1521);
nor U1643 (N_1643,N_1583,N_1509);
nand U1644 (N_1644,N_1519,N_1548);
and U1645 (N_1645,N_1500,N_1537);
nor U1646 (N_1646,N_1532,N_1542);
nor U1647 (N_1647,N_1556,N_1523);
nor U1648 (N_1648,N_1515,N_1566);
nor U1649 (N_1649,N_1558,N_1590);
or U1650 (N_1650,N_1543,N_1528);
and U1651 (N_1651,N_1576,N_1502);
nand U1652 (N_1652,N_1561,N_1548);
or U1653 (N_1653,N_1519,N_1588);
or U1654 (N_1654,N_1570,N_1530);
nor U1655 (N_1655,N_1524,N_1561);
nor U1656 (N_1656,N_1536,N_1554);
and U1657 (N_1657,N_1514,N_1515);
or U1658 (N_1658,N_1502,N_1588);
or U1659 (N_1659,N_1526,N_1535);
and U1660 (N_1660,N_1595,N_1570);
nor U1661 (N_1661,N_1567,N_1532);
or U1662 (N_1662,N_1587,N_1532);
and U1663 (N_1663,N_1532,N_1519);
and U1664 (N_1664,N_1502,N_1558);
or U1665 (N_1665,N_1513,N_1588);
nand U1666 (N_1666,N_1546,N_1538);
and U1667 (N_1667,N_1550,N_1531);
and U1668 (N_1668,N_1569,N_1545);
nor U1669 (N_1669,N_1580,N_1544);
or U1670 (N_1670,N_1556,N_1504);
nand U1671 (N_1671,N_1520,N_1587);
xor U1672 (N_1672,N_1536,N_1595);
nand U1673 (N_1673,N_1560,N_1518);
nor U1674 (N_1674,N_1561,N_1500);
nand U1675 (N_1675,N_1562,N_1543);
nor U1676 (N_1676,N_1506,N_1540);
nand U1677 (N_1677,N_1584,N_1598);
or U1678 (N_1678,N_1571,N_1514);
or U1679 (N_1679,N_1561,N_1556);
or U1680 (N_1680,N_1539,N_1570);
or U1681 (N_1681,N_1557,N_1510);
or U1682 (N_1682,N_1534,N_1531);
or U1683 (N_1683,N_1582,N_1572);
and U1684 (N_1684,N_1540,N_1565);
or U1685 (N_1685,N_1568,N_1533);
nand U1686 (N_1686,N_1556,N_1571);
xor U1687 (N_1687,N_1570,N_1525);
nand U1688 (N_1688,N_1555,N_1563);
xnor U1689 (N_1689,N_1517,N_1537);
nand U1690 (N_1690,N_1530,N_1586);
nor U1691 (N_1691,N_1542,N_1525);
and U1692 (N_1692,N_1510,N_1507);
nand U1693 (N_1693,N_1569,N_1573);
nor U1694 (N_1694,N_1508,N_1573);
nor U1695 (N_1695,N_1565,N_1530);
or U1696 (N_1696,N_1529,N_1523);
and U1697 (N_1697,N_1533,N_1547);
xnor U1698 (N_1698,N_1572,N_1593);
nor U1699 (N_1699,N_1514,N_1535);
nor U1700 (N_1700,N_1669,N_1601);
nor U1701 (N_1701,N_1612,N_1618);
and U1702 (N_1702,N_1687,N_1657);
nor U1703 (N_1703,N_1627,N_1609);
nand U1704 (N_1704,N_1625,N_1680);
xnor U1705 (N_1705,N_1651,N_1605);
and U1706 (N_1706,N_1613,N_1673);
nor U1707 (N_1707,N_1654,N_1642);
and U1708 (N_1708,N_1647,N_1626);
xnor U1709 (N_1709,N_1694,N_1659);
nand U1710 (N_1710,N_1636,N_1600);
xor U1711 (N_1711,N_1632,N_1629);
nor U1712 (N_1712,N_1663,N_1630);
and U1713 (N_1713,N_1634,N_1689);
nand U1714 (N_1714,N_1633,N_1695);
or U1715 (N_1715,N_1691,N_1666);
nor U1716 (N_1716,N_1697,N_1648);
xor U1717 (N_1717,N_1660,N_1682);
nand U1718 (N_1718,N_1641,N_1602);
nor U1719 (N_1719,N_1685,N_1635);
and U1720 (N_1720,N_1683,N_1646);
nand U1721 (N_1721,N_1645,N_1640);
nand U1722 (N_1722,N_1628,N_1631);
and U1723 (N_1723,N_1675,N_1606);
and U1724 (N_1724,N_1653,N_1698);
or U1725 (N_1725,N_1637,N_1644);
and U1726 (N_1726,N_1693,N_1655);
nor U1727 (N_1727,N_1686,N_1649);
nor U1728 (N_1728,N_1664,N_1622);
nand U1729 (N_1729,N_1604,N_1615);
nor U1730 (N_1730,N_1677,N_1674);
and U1731 (N_1731,N_1610,N_1603);
or U1732 (N_1732,N_1690,N_1696);
and U1733 (N_1733,N_1671,N_1608);
or U1734 (N_1734,N_1607,N_1624);
nand U1735 (N_1735,N_1678,N_1670);
nand U1736 (N_1736,N_1667,N_1620);
xnor U1737 (N_1737,N_1672,N_1652);
nor U1738 (N_1738,N_1614,N_1623);
nand U1739 (N_1739,N_1656,N_1639);
or U1740 (N_1740,N_1676,N_1658);
or U1741 (N_1741,N_1688,N_1619);
xnor U1742 (N_1742,N_1668,N_1643);
xor U1743 (N_1743,N_1684,N_1617);
nor U1744 (N_1744,N_1661,N_1681);
or U1745 (N_1745,N_1679,N_1692);
and U1746 (N_1746,N_1699,N_1638);
and U1747 (N_1747,N_1611,N_1621);
nand U1748 (N_1748,N_1616,N_1650);
nor U1749 (N_1749,N_1662,N_1665);
and U1750 (N_1750,N_1685,N_1632);
xor U1751 (N_1751,N_1684,N_1652);
and U1752 (N_1752,N_1669,N_1677);
or U1753 (N_1753,N_1691,N_1637);
and U1754 (N_1754,N_1641,N_1616);
and U1755 (N_1755,N_1627,N_1617);
and U1756 (N_1756,N_1695,N_1657);
nand U1757 (N_1757,N_1647,N_1640);
nor U1758 (N_1758,N_1645,N_1683);
or U1759 (N_1759,N_1669,N_1630);
nand U1760 (N_1760,N_1635,N_1696);
nand U1761 (N_1761,N_1681,N_1686);
or U1762 (N_1762,N_1622,N_1631);
and U1763 (N_1763,N_1630,N_1646);
and U1764 (N_1764,N_1644,N_1699);
or U1765 (N_1765,N_1616,N_1648);
and U1766 (N_1766,N_1612,N_1631);
or U1767 (N_1767,N_1620,N_1603);
nand U1768 (N_1768,N_1642,N_1619);
xnor U1769 (N_1769,N_1683,N_1635);
nor U1770 (N_1770,N_1603,N_1682);
nor U1771 (N_1771,N_1684,N_1601);
and U1772 (N_1772,N_1673,N_1681);
nand U1773 (N_1773,N_1620,N_1613);
nor U1774 (N_1774,N_1665,N_1694);
and U1775 (N_1775,N_1641,N_1671);
or U1776 (N_1776,N_1600,N_1625);
nand U1777 (N_1777,N_1648,N_1688);
nor U1778 (N_1778,N_1603,N_1691);
nor U1779 (N_1779,N_1682,N_1696);
nor U1780 (N_1780,N_1643,N_1601);
nor U1781 (N_1781,N_1687,N_1645);
nor U1782 (N_1782,N_1688,N_1678);
xnor U1783 (N_1783,N_1664,N_1663);
nor U1784 (N_1784,N_1676,N_1684);
xor U1785 (N_1785,N_1691,N_1662);
and U1786 (N_1786,N_1637,N_1623);
nor U1787 (N_1787,N_1674,N_1635);
nor U1788 (N_1788,N_1636,N_1622);
nor U1789 (N_1789,N_1648,N_1692);
nor U1790 (N_1790,N_1672,N_1661);
or U1791 (N_1791,N_1639,N_1681);
and U1792 (N_1792,N_1673,N_1675);
nor U1793 (N_1793,N_1698,N_1650);
or U1794 (N_1794,N_1649,N_1624);
nand U1795 (N_1795,N_1683,N_1662);
nand U1796 (N_1796,N_1603,N_1688);
xnor U1797 (N_1797,N_1683,N_1637);
and U1798 (N_1798,N_1633,N_1699);
nand U1799 (N_1799,N_1662,N_1604);
nand U1800 (N_1800,N_1758,N_1713);
nor U1801 (N_1801,N_1738,N_1779);
nor U1802 (N_1802,N_1705,N_1744);
xnor U1803 (N_1803,N_1799,N_1759);
and U1804 (N_1804,N_1726,N_1700);
or U1805 (N_1805,N_1720,N_1767);
and U1806 (N_1806,N_1786,N_1787);
nor U1807 (N_1807,N_1712,N_1798);
nand U1808 (N_1808,N_1765,N_1764);
or U1809 (N_1809,N_1703,N_1714);
nor U1810 (N_1810,N_1701,N_1788);
nor U1811 (N_1811,N_1721,N_1776);
nor U1812 (N_1812,N_1747,N_1741);
and U1813 (N_1813,N_1794,N_1711);
nand U1814 (N_1814,N_1774,N_1746);
or U1815 (N_1815,N_1743,N_1715);
or U1816 (N_1816,N_1732,N_1768);
or U1817 (N_1817,N_1761,N_1754);
and U1818 (N_1818,N_1708,N_1797);
nand U1819 (N_1819,N_1775,N_1763);
and U1820 (N_1820,N_1706,N_1772);
nand U1821 (N_1821,N_1737,N_1792);
or U1822 (N_1822,N_1760,N_1780);
or U1823 (N_1823,N_1756,N_1725);
nor U1824 (N_1824,N_1748,N_1778);
or U1825 (N_1825,N_1752,N_1782);
nand U1826 (N_1826,N_1777,N_1718);
xor U1827 (N_1827,N_1771,N_1745);
nand U1828 (N_1828,N_1722,N_1724);
nor U1829 (N_1829,N_1762,N_1729);
nand U1830 (N_1830,N_1769,N_1728);
nand U1831 (N_1831,N_1753,N_1719);
and U1832 (N_1832,N_1736,N_1734);
nand U1833 (N_1833,N_1727,N_1735);
nor U1834 (N_1834,N_1702,N_1751);
or U1835 (N_1835,N_1795,N_1723);
or U1836 (N_1836,N_1793,N_1757);
or U1837 (N_1837,N_1740,N_1770);
nand U1838 (N_1838,N_1716,N_1789);
xor U1839 (N_1839,N_1704,N_1784);
and U1840 (N_1840,N_1796,N_1766);
or U1841 (N_1841,N_1742,N_1773);
xnor U1842 (N_1842,N_1785,N_1731);
and U1843 (N_1843,N_1739,N_1755);
nand U1844 (N_1844,N_1783,N_1750);
and U1845 (N_1845,N_1710,N_1709);
nor U1846 (N_1846,N_1717,N_1707);
and U1847 (N_1847,N_1749,N_1791);
or U1848 (N_1848,N_1781,N_1733);
nand U1849 (N_1849,N_1730,N_1790);
xnor U1850 (N_1850,N_1704,N_1770);
nand U1851 (N_1851,N_1711,N_1743);
nand U1852 (N_1852,N_1751,N_1704);
or U1853 (N_1853,N_1766,N_1732);
or U1854 (N_1854,N_1751,N_1786);
nor U1855 (N_1855,N_1766,N_1736);
or U1856 (N_1856,N_1729,N_1776);
nand U1857 (N_1857,N_1766,N_1719);
or U1858 (N_1858,N_1729,N_1761);
and U1859 (N_1859,N_1706,N_1738);
and U1860 (N_1860,N_1731,N_1746);
nor U1861 (N_1861,N_1787,N_1723);
nand U1862 (N_1862,N_1733,N_1798);
nor U1863 (N_1863,N_1737,N_1710);
and U1864 (N_1864,N_1771,N_1788);
or U1865 (N_1865,N_1765,N_1768);
nor U1866 (N_1866,N_1712,N_1784);
and U1867 (N_1867,N_1725,N_1720);
nor U1868 (N_1868,N_1754,N_1755);
nand U1869 (N_1869,N_1779,N_1776);
nor U1870 (N_1870,N_1787,N_1725);
and U1871 (N_1871,N_1760,N_1799);
xor U1872 (N_1872,N_1703,N_1787);
and U1873 (N_1873,N_1734,N_1723);
and U1874 (N_1874,N_1704,N_1753);
or U1875 (N_1875,N_1721,N_1748);
nand U1876 (N_1876,N_1777,N_1712);
and U1877 (N_1877,N_1772,N_1725);
or U1878 (N_1878,N_1787,N_1760);
or U1879 (N_1879,N_1705,N_1787);
nor U1880 (N_1880,N_1703,N_1797);
or U1881 (N_1881,N_1773,N_1767);
and U1882 (N_1882,N_1780,N_1764);
nand U1883 (N_1883,N_1798,N_1745);
nand U1884 (N_1884,N_1761,N_1769);
nor U1885 (N_1885,N_1759,N_1793);
nor U1886 (N_1886,N_1754,N_1766);
xor U1887 (N_1887,N_1745,N_1770);
or U1888 (N_1888,N_1738,N_1742);
and U1889 (N_1889,N_1726,N_1740);
xnor U1890 (N_1890,N_1758,N_1701);
nor U1891 (N_1891,N_1756,N_1727);
and U1892 (N_1892,N_1790,N_1745);
and U1893 (N_1893,N_1719,N_1723);
nand U1894 (N_1894,N_1786,N_1718);
or U1895 (N_1895,N_1702,N_1723);
nand U1896 (N_1896,N_1702,N_1736);
nand U1897 (N_1897,N_1708,N_1761);
nor U1898 (N_1898,N_1769,N_1774);
and U1899 (N_1899,N_1747,N_1762);
nand U1900 (N_1900,N_1807,N_1827);
and U1901 (N_1901,N_1882,N_1876);
and U1902 (N_1902,N_1813,N_1852);
or U1903 (N_1903,N_1802,N_1870);
xnor U1904 (N_1904,N_1898,N_1844);
xor U1905 (N_1905,N_1843,N_1808);
xor U1906 (N_1906,N_1848,N_1873);
nand U1907 (N_1907,N_1824,N_1828);
xor U1908 (N_1908,N_1879,N_1834);
and U1909 (N_1909,N_1842,N_1819);
and U1910 (N_1910,N_1845,N_1855);
nor U1911 (N_1911,N_1887,N_1829);
nand U1912 (N_1912,N_1877,N_1854);
xnor U1913 (N_1913,N_1821,N_1899);
or U1914 (N_1914,N_1884,N_1818);
or U1915 (N_1915,N_1892,N_1810);
and U1916 (N_1916,N_1874,N_1889);
nor U1917 (N_1917,N_1841,N_1860);
or U1918 (N_1918,N_1851,N_1835);
xor U1919 (N_1919,N_1896,N_1814);
nand U1920 (N_1920,N_1862,N_1832);
xnor U1921 (N_1921,N_1812,N_1867);
nor U1922 (N_1922,N_1857,N_1811);
or U1923 (N_1923,N_1800,N_1809);
xor U1924 (N_1924,N_1866,N_1839);
xnor U1925 (N_1925,N_1849,N_1806);
or U1926 (N_1926,N_1847,N_1886);
or U1927 (N_1927,N_1850,N_1803);
xnor U1928 (N_1928,N_1893,N_1880);
nor U1929 (N_1929,N_1826,N_1817);
and U1930 (N_1930,N_1859,N_1816);
nor U1931 (N_1931,N_1837,N_1853);
nand U1932 (N_1932,N_1846,N_1840);
or U1933 (N_1933,N_1885,N_1897);
nand U1934 (N_1934,N_1805,N_1864);
nand U1935 (N_1935,N_1830,N_1804);
or U1936 (N_1936,N_1868,N_1878);
nand U1937 (N_1937,N_1863,N_1838);
nor U1938 (N_1938,N_1883,N_1823);
or U1939 (N_1939,N_1858,N_1831);
nand U1940 (N_1940,N_1895,N_1865);
or U1941 (N_1941,N_1856,N_1871);
xnor U1942 (N_1942,N_1801,N_1894);
nand U1943 (N_1943,N_1891,N_1888);
xnor U1944 (N_1944,N_1881,N_1825);
or U1945 (N_1945,N_1872,N_1815);
or U1946 (N_1946,N_1822,N_1890);
or U1947 (N_1947,N_1820,N_1833);
and U1948 (N_1948,N_1869,N_1836);
nand U1949 (N_1949,N_1861,N_1875);
nand U1950 (N_1950,N_1830,N_1891);
nor U1951 (N_1951,N_1821,N_1898);
nor U1952 (N_1952,N_1894,N_1828);
nand U1953 (N_1953,N_1838,N_1854);
or U1954 (N_1954,N_1878,N_1887);
and U1955 (N_1955,N_1850,N_1885);
xor U1956 (N_1956,N_1813,N_1874);
and U1957 (N_1957,N_1809,N_1817);
xor U1958 (N_1958,N_1864,N_1859);
or U1959 (N_1959,N_1882,N_1801);
nor U1960 (N_1960,N_1836,N_1838);
nor U1961 (N_1961,N_1891,N_1814);
xor U1962 (N_1962,N_1800,N_1829);
nand U1963 (N_1963,N_1842,N_1868);
nor U1964 (N_1964,N_1892,N_1811);
and U1965 (N_1965,N_1843,N_1814);
or U1966 (N_1966,N_1867,N_1852);
and U1967 (N_1967,N_1836,N_1863);
nand U1968 (N_1968,N_1819,N_1834);
nand U1969 (N_1969,N_1843,N_1822);
and U1970 (N_1970,N_1875,N_1897);
nand U1971 (N_1971,N_1899,N_1825);
nand U1972 (N_1972,N_1849,N_1848);
nand U1973 (N_1973,N_1877,N_1896);
xor U1974 (N_1974,N_1863,N_1862);
and U1975 (N_1975,N_1825,N_1855);
and U1976 (N_1976,N_1824,N_1860);
nand U1977 (N_1977,N_1815,N_1861);
and U1978 (N_1978,N_1853,N_1869);
nand U1979 (N_1979,N_1899,N_1860);
xnor U1980 (N_1980,N_1857,N_1845);
nor U1981 (N_1981,N_1857,N_1846);
or U1982 (N_1982,N_1887,N_1801);
nand U1983 (N_1983,N_1886,N_1882);
nand U1984 (N_1984,N_1842,N_1884);
nand U1985 (N_1985,N_1879,N_1802);
nor U1986 (N_1986,N_1889,N_1817);
nand U1987 (N_1987,N_1815,N_1834);
nand U1988 (N_1988,N_1888,N_1802);
nand U1989 (N_1989,N_1840,N_1841);
nand U1990 (N_1990,N_1804,N_1835);
nand U1991 (N_1991,N_1846,N_1862);
nand U1992 (N_1992,N_1895,N_1864);
nand U1993 (N_1993,N_1888,N_1813);
or U1994 (N_1994,N_1830,N_1815);
nand U1995 (N_1995,N_1865,N_1803);
or U1996 (N_1996,N_1840,N_1833);
nor U1997 (N_1997,N_1848,N_1819);
nor U1998 (N_1998,N_1834,N_1833);
nand U1999 (N_1999,N_1816,N_1804);
xor U2000 (N_2000,N_1988,N_1905);
nor U2001 (N_2001,N_1969,N_1944);
nand U2002 (N_2002,N_1939,N_1950);
xor U2003 (N_2003,N_1959,N_1966);
or U2004 (N_2004,N_1979,N_1990);
nor U2005 (N_2005,N_1954,N_1921);
or U2006 (N_2006,N_1951,N_1945);
xor U2007 (N_2007,N_1927,N_1903);
nor U2008 (N_2008,N_1948,N_1914);
or U2009 (N_2009,N_1992,N_1996);
and U2010 (N_2010,N_1961,N_1952);
and U2011 (N_2011,N_1955,N_1929);
and U2012 (N_2012,N_1920,N_1922);
and U2013 (N_2013,N_1989,N_1981);
nand U2014 (N_2014,N_1912,N_1975);
nand U2015 (N_2015,N_1940,N_1984);
nor U2016 (N_2016,N_1962,N_1997);
and U2017 (N_2017,N_1946,N_1973);
or U2018 (N_2018,N_1931,N_1924);
nand U2019 (N_2019,N_1917,N_1998);
nor U2020 (N_2020,N_1915,N_1933);
or U2021 (N_2021,N_1980,N_1938);
xnor U2022 (N_2022,N_1908,N_1906);
nand U2023 (N_2023,N_1986,N_1904);
xnor U2024 (N_2024,N_1971,N_1991);
and U2025 (N_2025,N_1918,N_1956);
and U2026 (N_2026,N_1926,N_1923);
nand U2027 (N_2027,N_1993,N_1970);
nor U2028 (N_2028,N_1943,N_1982);
nor U2029 (N_2029,N_1941,N_1974);
nor U2030 (N_2030,N_1947,N_1963);
xnor U2031 (N_2031,N_1983,N_1958);
and U2032 (N_2032,N_1999,N_1911);
nor U2033 (N_2033,N_1978,N_1942);
xnor U2034 (N_2034,N_1901,N_1900);
and U2035 (N_2035,N_1964,N_1953);
nand U2036 (N_2036,N_1965,N_1977);
or U2037 (N_2037,N_1913,N_1930);
or U2038 (N_2038,N_1967,N_1995);
or U2039 (N_2039,N_1968,N_1985);
and U2040 (N_2040,N_1928,N_1976);
nand U2041 (N_2041,N_1919,N_1987);
and U2042 (N_2042,N_1925,N_1932);
nor U2043 (N_2043,N_1949,N_1994);
or U2044 (N_2044,N_1916,N_1935);
and U2045 (N_2045,N_1910,N_1936);
nor U2046 (N_2046,N_1907,N_1972);
and U2047 (N_2047,N_1960,N_1937);
and U2048 (N_2048,N_1934,N_1902);
and U2049 (N_2049,N_1909,N_1957);
or U2050 (N_2050,N_1913,N_1995);
xnor U2051 (N_2051,N_1952,N_1911);
or U2052 (N_2052,N_1950,N_1949);
nand U2053 (N_2053,N_1920,N_1916);
nand U2054 (N_2054,N_1911,N_1941);
or U2055 (N_2055,N_1905,N_1987);
nand U2056 (N_2056,N_1921,N_1909);
or U2057 (N_2057,N_1918,N_1909);
nand U2058 (N_2058,N_1924,N_1921);
and U2059 (N_2059,N_1987,N_1900);
nand U2060 (N_2060,N_1925,N_1917);
nor U2061 (N_2061,N_1916,N_1954);
or U2062 (N_2062,N_1962,N_1939);
nor U2063 (N_2063,N_1948,N_1974);
xor U2064 (N_2064,N_1922,N_1946);
xnor U2065 (N_2065,N_1965,N_1919);
or U2066 (N_2066,N_1924,N_1917);
or U2067 (N_2067,N_1952,N_1936);
nand U2068 (N_2068,N_1910,N_1994);
xnor U2069 (N_2069,N_1971,N_1986);
and U2070 (N_2070,N_1935,N_1994);
nor U2071 (N_2071,N_1976,N_1933);
nand U2072 (N_2072,N_1932,N_1909);
xnor U2073 (N_2073,N_1994,N_1914);
nand U2074 (N_2074,N_1982,N_1935);
and U2075 (N_2075,N_1963,N_1957);
and U2076 (N_2076,N_1963,N_1992);
nand U2077 (N_2077,N_1983,N_1903);
and U2078 (N_2078,N_1944,N_1956);
xor U2079 (N_2079,N_1922,N_1953);
nand U2080 (N_2080,N_1900,N_1935);
nand U2081 (N_2081,N_1915,N_1928);
nor U2082 (N_2082,N_1958,N_1985);
and U2083 (N_2083,N_1979,N_1959);
nand U2084 (N_2084,N_1987,N_1980);
and U2085 (N_2085,N_1905,N_1913);
nand U2086 (N_2086,N_1976,N_1925);
or U2087 (N_2087,N_1923,N_1955);
or U2088 (N_2088,N_1901,N_1993);
xnor U2089 (N_2089,N_1975,N_1905);
and U2090 (N_2090,N_1987,N_1963);
and U2091 (N_2091,N_1958,N_1948);
nand U2092 (N_2092,N_1989,N_1982);
nand U2093 (N_2093,N_1959,N_1935);
nor U2094 (N_2094,N_1947,N_1976);
xor U2095 (N_2095,N_1958,N_1996);
xnor U2096 (N_2096,N_1968,N_1927);
and U2097 (N_2097,N_1961,N_1918);
nand U2098 (N_2098,N_1902,N_1904);
or U2099 (N_2099,N_1959,N_1910);
nor U2100 (N_2100,N_2018,N_2083);
nand U2101 (N_2101,N_2076,N_2050);
or U2102 (N_2102,N_2012,N_2031);
nor U2103 (N_2103,N_2042,N_2023);
and U2104 (N_2104,N_2049,N_2041);
xnor U2105 (N_2105,N_2069,N_2089);
nor U2106 (N_2106,N_2040,N_2030);
nand U2107 (N_2107,N_2066,N_2084);
and U2108 (N_2108,N_2005,N_2071);
xnor U2109 (N_2109,N_2019,N_2096);
or U2110 (N_2110,N_2044,N_2022);
xor U2111 (N_2111,N_2015,N_2059);
nand U2112 (N_2112,N_2046,N_2007);
and U2113 (N_2113,N_2036,N_2025);
nor U2114 (N_2114,N_2016,N_2011);
and U2115 (N_2115,N_2087,N_2056);
and U2116 (N_2116,N_2010,N_2038);
and U2117 (N_2117,N_2091,N_2065);
nand U2118 (N_2118,N_2034,N_2064);
or U2119 (N_2119,N_2004,N_2098);
nand U2120 (N_2120,N_2047,N_2073);
nor U2121 (N_2121,N_2000,N_2099);
and U2122 (N_2122,N_2080,N_2002);
or U2123 (N_2123,N_2020,N_2053);
nor U2124 (N_2124,N_2088,N_2075);
nor U2125 (N_2125,N_2063,N_2039);
and U2126 (N_2126,N_2074,N_2061);
xor U2127 (N_2127,N_2068,N_2057);
or U2128 (N_2128,N_2013,N_2090);
xnor U2129 (N_2129,N_2055,N_2035);
or U2130 (N_2130,N_2093,N_2085);
nand U2131 (N_2131,N_2060,N_2048);
nor U2132 (N_2132,N_2052,N_2009);
or U2133 (N_2133,N_2045,N_2062);
or U2134 (N_2134,N_2021,N_2094);
nor U2135 (N_2135,N_2072,N_2033);
nand U2136 (N_2136,N_2051,N_2095);
and U2137 (N_2137,N_2017,N_2054);
nor U2138 (N_2138,N_2077,N_2014);
or U2139 (N_2139,N_2070,N_2082);
and U2140 (N_2140,N_2086,N_2027);
and U2141 (N_2141,N_2097,N_2078);
nand U2142 (N_2142,N_2001,N_2079);
nand U2143 (N_2143,N_2043,N_2006);
nor U2144 (N_2144,N_2081,N_2037);
and U2145 (N_2145,N_2067,N_2032);
or U2146 (N_2146,N_2003,N_2092);
or U2147 (N_2147,N_2028,N_2024);
nor U2148 (N_2148,N_2026,N_2008);
and U2149 (N_2149,N_2029,N_2058);
and U2150 (N_2150,N_2080,N_2085);
nand U2151 (N_2151,N_2050,N_2088);
and U2152 (N_2152,N_2020,N_2048);
xnor U2153 (N_2153,N_2075,N_2068);
or U2154 (N_2154,N_2014,N_2029);
nand U2155 (N_2155,N_2033,N_2093);
nor U2156 (N_2156,N_2092,N_2051);
xor U2157 (N_2157,N_2088,N_2008);
and U2158 (N_2158,N_2052,N_2081);
or U2159 (N_2159,N_2082,N_2092);
nand U2160 (N_2160,N_2030,N_2036);
and U2161 (N_2161,N_2014,N_2026);
and U2162 (N_2162,N_2066,N_2016);
or U2163 (N_2163,N_2037,N_2057);
nand U2164 (N_2164,N_2004,N_2042);
and U2165 (N_2165,N_2083,N_2017);
and U2166 (N_2166,N_2012,N_2033);
nor U2167 (N_2167,N_2020,N_2035);
nor U2168 (N_2168,N_2076,N_2043);
nor U2169 (N_2169,N_2008,N_2040);
nor U2170 (N_2170,N_2027,N_2025);
nand U2171 (N_2171,N_2028,N_2009);
nand U2172 (N_2172,N_2011,N_2056);
or U2173 (N_2173,N_2089,N_2057);
nor U2174 (N_2174,N_2013,N_2079);
nor U2175 (N_2175,N_2026,N_2001);
nor U2176 (N_2176,N_2092,N_2033);
xnor U2177 (N_2177,N_2090,N_2021);
and U2178 (N_2178,N_2035,N_2010);
nand U2179 (N_2179,N_2036,N_2034);
and U2180 (N_2180,N_2068,N_2084);
and U2181 (N_2181,N_2084,N_2092);
nor U2182 (N_2182,N_2070,N_2092);
nand U2183 (N_2183,N_2069,N_2019);
and U2184 (N_2184,N_2096,N_2008);
nand U2185 (N_2185,N_2014,N_2089);
nand U2186 (N_2186,N_2019,N_2092);
or U2187 (N_2187,N_2035,N_2074);
nor U2188 (N_2188,N_2060,N_2030);
or U2189 (N_2189,N_2046,N_2010);
and U2190 (N_2190,N_2083,N_2001);
and U2191 (N_2191,N_2097,N_2013);
or U2192 (N_2192,N_2060,N_2053);
xor U2193 (N_2193,N_2005,N_2039);
xnor U2194 (N_2194,N_2085,N_2033);
and U2195 (N_2195,N_2003,N_2088);
nor U2196 (N_2196,N_2031,N_2044);
or U2197 (N_2197,N_2049,N_2085);
or U2198 (N_2198,N_2079,N_2029);
or U2199 (N_2199,N_2055,N_2031);
and U2200 (N_2200,N_2123,N_2111);
and U2201 (N_2201,N_2107,N_2175);
and U2202 (N_2202,N_2177,N_2159);
or U2203 (N_2203,N_2134,N_2190);
nor U2204 (N_2204,N_2194,N_2127);
nor U2205 (N_2205,N_2112,N_2145);
nor U2206 (N_2206,N_2152,N_2120);
or U2207 (N_2207,N_2105,N_2121);
nor U2208 (N_2208,N_2176,N_2181);
and U2209 (N_2209,N_2189,N_2114);
nor U2210 (N_2210,N_2163,N_2165);
nor U2211 (N_2211,N_2183,N_2170);
or U2212 (N_2212,N_2137,N_2160);
nor U2213 (N_2213,N_2199,N_2122);
nand U2214 (N_2214,N_2106,N_2125);
nand U2215 (N_2215,N_2180,N_2158);
and U2216 (N_2216,N_2157,N_2128);
nand U2217 (N_2217,N_2119,N_2117);
and U2218 (N_2218,N_2130,N_2168);
and U2219 (N_2219,N_2191,N_2133);
and U2220 (N_2220,N_2193,N_2100);
and U2221 (N_2221,N_2108,N_2167);
and U2222 (N_2222,N_2148,N_2103);
nand U2223 (N_2223,N_2192,N_2118);
and U2224 (N_2224,N_2172,N_2186);
nor U2225 (N_2225,N_2161,N_2169);
and U2226 (N_2226,N_2185,N_2138);
and U2227 (N_2227,N_2173,N_2198);
or U2228 (N_2228,N_2124,N_2101);
nand U2229 (N_2229,N_2151,N_2156);
or U2230 (N_2230,N_2196,N_2116);
xor U2231 (N_2231,N_2142,N_2187);
nor U2232 (N_2232,N_2131,N_2144);
xnor U2233 (N_2233,N_2102,N_2182);
xnor U2234 (N_2234,N_2146,N_2150);
xor U2235 (N_2235,N_2155,N_2162);
nor U2236 (N_2236,N_2115,N_2174);
nand U2237 (N_2237,N_2143,N_2141);
xor U2238 (N_2238,N_2154,N_2110);
and U2239 (N_2239,N_2140,N_2136);
and U2240 (N_2240,N_2184,N_2147);
xnor U2241 (N_2241,N_2164,N_2171);
nand U2242 (N_2242,N_2126,N_2197);
and U2243 (N_2243,N_2149,N_2139);
and U2244 (N_2244,N_2132,N_2109);
nor U2245 (N_2245,N_2129,N_2166);
xnor U2246 (N_2246,N_2113,N_2178);
nor U2247 (N_2247,N_2179,N_2195);
nand U2248 (N_2248,N_2135,N_2188);
nor U2249 (N_2249,N_2153,N_2104);
nor U2250 (N_2250,N_2170,N_2164);
nand U2251 (N_2251,N_2179,N_2162);
nor U2252 (N_2252,N_2199,N_2196);
nor U2253 (N_2253,N_2153,N_2108);
and U2254 (N_2254,N_2188,N_2179);
or U2255 (N_2255,N_2126,N_2102);
nor U2256 (N_2256,N_2136,N_2107);
nor U2257 (N_2257,N_2185,N_2146);
nand U2258 (N_2258,N_2109,N_2196);
nor U2259 (N_2259,N_2146,N_2145);
or U2260 (N_2260,N_2137,N_2146);
nand U2261 (N_2261,N_2193,N_2161);
or U2262 (N_2262,N_2163,N_2193);
nor U2263 (N_2263,N_2151,N_2154);
and U2264 (N_2264,N_2186,N_2109);
nor U2265 (N_2265,N_2186,N_2150);
xor U2266 (N_2266,N_2140,N_2155);
and U2267 (N_2267,N_2169,N_2145);
or U2268 (N_2268,N_2176,N_2137);
or U2269 (N_2269,N_2163,N_2115);
or U2270 (N_2270,N_2104,N_2110);
nand U2271 (N_2271,N_2117,N_2163);
nand U2272 (N_2272,N_2152,N_2142);
or U2273 (N_2273,N_2175,N_2186);
nor U2274 (N_2274,N_2177,N_2156);
nand U2275 (N_2275,N_2174,N_2183);
and U2276 (N_2276,N_2175,N_2137);
or U2277 (N_2277,N_2162,N_2102);
xnor U2278 (N_2278,N_2115,N_2154);
and U2279 (N_2279,N_2143,N_2100);
or U2280 (N_2280,N_2138,N_2168);
nor U2281 (N_2281,N_2135,N_2186);
nand U2282 (N_2282,N_2145,N_2101);
and U2283 (N_2283,N_2172,N_2150);
nor U2284 (N_2284,N_2127,N_2134);
or U2285 (N_2285,N_2125,N_2197);
nand U2286 (N_2286,N_2180,N_2166);
or U2287 (N_2287,N_2131,N_2128);
nand U2288 (N_2288,N_2118,N_2131);
or U2289 (N_2289,N_2103,N_2183);
or U2290 (N_2290,N_2108,N_2165);
nand U2291 (N_2291,N_2100,N_2152);
and U2292 (N_2292,N_2117,N_2127);
nor U2293 (N_2293,N_2118,N_2136);
or U2294 (N_2294,N_2164,N_2153);
nand U2295 (N_2295,N_2146,N_2194);
or U2296 (N_2296,N_2183,N_2191);
or U2297 (N_2297,N_2158,N_2112);
and U2298 (N_2298,N_2116,N_2183);
and U2299 (N_2299,N_2131,N_2107);
or U2300 (N_2300,N_2246,N_2206);
and U2301 (N_2301,N_2245,N_2213);
and U2302 (N_2302,N_2231,N_2235);
nand U2303 (N_2303,N_2211,N_2200);
and U2304 (N_2304,N_2215,N_2227);
and U2305 (N_2305,N_2296,N_2252);
nand U2306 (N_2306,N_2265,N_2266);
xor U2307 (N_2307,N_2278,N_2279);
xor U2308 (N_2308,N_2268,N_2255);
or U2309 (N_2309,N_2277,N_2273);
nor U2310 (N_2310,N_2230,N_2250);
or U2311 (N_2311,N_2299,N_2244);
and U2312 (N_2312,N_2205,N_2261);
nor U2313 (N_2313,N_2292,N_2247);
nand U2314 (N_2314,N_2280,N_2276);
and U2315 (N_2315,N_2254,N_2288);
nor U2316 (N_2316,N_2289,N_2294);
or U2317 (N_2317,N_2241,N_2256);
nor U2318 (N_2318,N_2238,N_2282);
nand U2319 (N_2319,N_2290,N_2228);
and U2320 (N_2320,N_2239,N_2214);
or U2321 (N_2321,N_2269,N_2207);
xnor U2322 (N_2322,N_2201,N_2218);
xor U2323 (N_2323,N_2223,N_2291);
or U2324 (N_2324,N_2234,N_2293);
and U2325 (N_2325,N_2210,N_2226);
nor U2326 (N_2326,N_2233,N_2259);
and U2327 (N_2327,N_2267,N_2283);
nand U2328 (N_2328,N_2253,N_2203);
nor U2329 (N_2329,N_2216,N_2281);
or U2330 (N_2330,N_2204,N_2242);
or U2331 (N_2331,N_2251,N_2224);
or U2332 (N_2332,N_2208,N_2209);
nor U2333 (N_2333,N_2237,N_2260);
xnor U2334 (N_2334,N_2202,N_2270);
and U2335 (N_2335,N_2263,N_2225);
or U2336 (N_2336,N_2220,N_2221);
or U2337 (N_2337,N_2229,N_2212);
and U2338 (N_2338,N_2274,N_2284);
nor U2339 (N_2339,N_2287,N_2286);
nand U2340 (N_2340,N_2236,N_2217);
or U2341 (N_2341,N_2240,N_2232);
nand U2342 (N_2342,N_2285,N_2295);
nor U2343 (N_2343,N_2249,N_2222);
xor U2344 (N_2344,N_2264,N_2297);
nor U2345 (N_2345,N_2258,N_2262);
nor U2346 (N_2346,N_2275,N_2248);
nand U2347 (N_2347,N_2257,N_2298);
nor U2348 (N_2348,N_2272,N_2243);
or U2349 (N_2349,N_2219,N_2271);
xor U2350 (N_2350,N_2219,N_2215);
nand U2351 (N_2351,N_2228,N_2216);
or U2352 (N_2352,N_2268,N_2224);
or U2353 (N_2353,N_2231,N_2207);
nand U2354 (N_2354,N_2293,N_2244);
and U2355 (N_2355,N_2275,N_2249);
and U2356 (N_2356,N_2248,N_2232);
or U2357 (N_2357,N_2294,N_2266);
or U2358 (N_2358,N_2270,N_2217);
nand U2359 (N_2359,N_2235,N_2257);
nand U2360 (N_2360,N_2280,N_2217);
or U2361 (N_2361,N_2227,N_2271);
nand U2362 (N_2362,N_2283,N_2263);
or U2363 (N_2363,N_2244,N_2285);
nand U2364 (N_2364,N_2260,N_2261);
or U2365 (N_2365,N_2254,N_2248);
nand U2366 (N_2366,N_2288,N_2273);
or U2367 (N_2367,N_2261,N_2285);
xor U2368 (N_2368,N_2222,N_2287);
or U2369 (N_2369,N_2251,N_2270);
nor U2370 (N_2370,N_2206,N_2217);
nor U2371 (N_2371,N_2288,N_2201);
or U2372 (N_2372,N_2295,N_2283);
nand U2373 (N_2373,N_2215,N_2269);
and U2374 (N_2374,N_2281,N_2243);
or U2375 (N_2375,N_2224,N_2297);
nand U2376 (N_2376,N_2292,N_2239);
nor U2377 (N_2377,N_2294,N_2224);
nand U2378 (N_2378,N_2258,N_2299);
or U2379 (N_2379,N_2221,N_2273);
nand U2380 (N_2380,N_2261,N_2215);
and U2381 (N_2381,N_2229,N_2289);
or U2382 (N_2382,N_2289,N_2250);
and U2383 (N_2383,N_2210,N_2286);
and U2384 (N_2384,N_2257,N_2238);
nor U2385 (N_2385,N_2231,N_2280);
nor U2386 (N_2386,N_2260,N_2257);
nand U2387 (N_2387,N_2286,N_2250);
or U2388 (N_2388,N_2299,N_2242);
nor U2389 (N_2389,N_2213,N_2252);
or U2390 (N_2390,N_2230,N_2227);
nand U2391 (N_2391,N_2233,N_2265);
nand U2392 (N_2392,N_2268,N_2296);
nor U2393 (N_2393,N_2211,N_2234);
xor U2394 (N_2394,N_2207,N_2220);
xnor U2395 (N_2395,N_2235,N_2252);
or U2396 (N_2396,N_2202,N_2228);
and U2397 (N_2397,N_2253,N_2263);
or U2398 (N_2398,N_2209,N_2200);
and U2399 (N_2399,N_2258,N_2245);
and U2400 (N_2400,N_2319,N_2312);
and U2401 (N_2401,N_2334,N_2385);
xnor U2402 (N_2402,N_2311,N_2373);
xor U2403 (N_2403,N_2304,N_2300);
xnor U2404 (N_2404,N_2364,N_2383);
or U2405 (N_2405,N_2326,N_2344);
xnor U2406 (N_2406,N_2374,N_2320);
nor U2407 (N_2407,N_2305,N_2372);
and U2408 (N_2408,N_2313,N_2356);
nand U2409 (N_2409,N_2331,N_2324);
and U2410 (N_2410,N_2370,N_2395);
nand U2411 (N_2411,N_2302,N_2382);
or U2412 (N_2412,N_2307,N_2361);
xor U2413 (N_2413,N_2301,N_2399);
or U2414 (N_2414,N_2323,N_2368);
and U2415 (N_2415,N_2354,N_2365);
nor U2416 (N_2416,N_2387,N_2343);
and U2417 (N_2417,N_2371,N_2316);
or U2418 (N_2418,N_2315,N_2380);
nor U2419 (N_2419,N_2366,N_2393);
nor U2420 (N_2420,N_2321,N_2329);
or U2421 (N_2421,N_2336,N_2359);
and U2422 (N_2422,N_2322,N_2338);
nand U2423 (N_2423,N_2310,N_2363);
or U2424 (N_2424,N_2394,N_2389);
xor U2425 (N_2425,N_2335,N_2340);
nor U2426 (N_2426,N_2381,N_2391);
or U2427 (N_2427,N_2339,N_2396);
and U2428 (N_2428,N_2328,N_2306);
or U2429 (N_2429,N_2349,N_2347);
or U2430 (N_2430,N_2352,N_2386);
and U2431 (N_2431,N_2346,N_2309);
and U2432 (N_2432,N_2342,N_2350);
and U2433 (N_2433,N_2358,N_2314);
or U2434 (N_2434,N_2303,N_2308);
and U2435 (N_2435,N_2369,N_2397);
nor U2436 (N_2436,N_2379,N_2360);
nor U2437 (N_2437,N_2377,N_2317);
xor U2438 (N_2438,N_2348,N_2330);
nand U2439 (N_2439,N_2392,N_2375);
nand U2440 (N_2440,N_2362,N_2357);
or U2441 (N_2441,N_2376,N_2390);
and U2442 (N_2442,N_2388,N_2353);
or U2443 (N_2443,N_2318,N_2332);
and U2444 (N_2444,N_2333,N_2384);
and U2445 (N_2445,N_2378,N_2327);
nor U2446 (N_2446,N_2398,N_2341);
xor U2447 (N_2447,N_2355,N_2345);
or U2448 (N_2448,N_2337,N_2351);
or U2449 (N_2449,N_2325,N_2367);
or U2450 (N_2450,N_2304,N_2365);
xnor U2451 (N_2451,N_2303,N_2360);
nand U2452 (N_2452,N_2384,N_2368);
nand U2453 (N_2453,N_2356,N_2336);
and U2454 (N_2454,N_2379,N_2384);
nor U2455 (N_2455,N_2318,N_2325);
nor U2456 (N_2456,N_2341,N_2394);
nand U2457 (N_2457,N_2302,N_2333);
and U2458 (N_2458,N_2357,N_2366);
nand U2459 (N_2459,N_2305,N_2307);
nand U2460 (N_2460,N_2340,N_2387);
or U2461 (N_2461,N_2375,N_2313);
nor U2462 (N_2462,N_2311,N_2395);
nand U2463 (N_2463,N_2322,N_2301);
or U2464 (N_2464,N_2389,N_2386);
nand U2465 (N_2465,N_2303,N_2340);
or U2466 (N_2466,N_2338,N_2314);
or U2467 (N_2467,N_2359,N_2387);
xor U2468 (N_2468,N_2371,N_2320);
nand U2469 (N_2469,N_2360,N_2344);
and U2470 (N_2470,N_2349,N_2355);
nor U2471 (N_2471,N_2307,N_2380);
nand U2472 (N_2472,N_2303,N_2382);
or U2473 (N_2473,N_2314,N_2328);
nand U2474 (N_2474,N_2332,N_2354);
and U2475 (N_2475,N_2316,N_2304);
and U2476 (N_2476,N_2346,N_2320);
nand U2477 (N_2477,N_2347,N_2320);
nor U2478 (N_2478,N_2319,N_2384);
and U2479 (N_2479,N_2361,N_2341);
nand U2480 (N_2480,N_2307,N_2331);
nand U2481 (N_2481,N_2320,N_2357);
nor U2482 (N_2482,N_2383,N_2317);
and U2483 (N_2483,N_2312,N_2375);
and U2484 (N_2484,N_2396,N_2380);
and U2485 (N_2485,N_2344,N_2316);
nand U2486 (N_2486,N_2326,N_2397);
and U2487 (N_2487,N_2305,N_2328);
nand U2488 (N_2488,N_2332,N_2373);
and U2489 (N_2489,N_2333,N_2325);
nand U2490 (N_2490,N_2312,N_2353);
nor U2491 (N_2491,N_2323,N_2377);
nor U2492 (N_2492,N_2340,N_2349);
or U2493 (N_2493,N_2325,N_2337);
and U2494 (N_2494,N_2399,N_2345);
and U2495 (N_2495,N_2324,N_2321);
nor U2496 (N_2496,N_2369,N_2348);
and U2497 (N_2497,N_2319,N_2367);
nand U2498 (N_2498,N_2345,N_2327);
nand U2499 (N_2499,N_2342,N_2317);
nand U2500 (N_2500,N_2441,N_2400);
nand U2501 (N_2501,N_2463,N_2469);
or U2502 (N_2502,N_2452,N_2409);
nand U2503 (N_2503,N_2481,N_2450);
nand U2504 (N_2504,N_2487,N_2453);
or U2505 (N_2505,N_2478,N_2454);
or U2506 (N_2506,N_2422,N_2423);
and U2507 (N_2507,N_2421,N_2444);
nand U2508 (N_2508,N_2430,N_2424);
or U2509 (N_2509,N_2451,N_2494);
or U2510 (N_2510,N_2425,N_2483);
and U2511 (N_2511,N_2435,N_2417);
nor U2512 (N_2512,N_2429,N_2490);
nor U2513 (N_2513,N_2499,N_2447);
nand U2514 (N_2514,N_2406,N_2471);
nand U2515 (N_2515,N_2467,N_2436);
nor U2516 (N_2516,N_2489,N_2411);
or U2517 (N_2517,N_2443,N_2464);
nor U2518 (N_2518,N_2412,N_2437);
nand U2519 (N_2519,N_2474,N_2468);
nor U2520 (N_2520,N_2457,N_2488);
nand U2521 (N_2521,N_2479,N_2413);
nor U2522 (N_2522,N_2404,N_2475);
or U2523 (N_2523,N_2456,N_2431);
nand U2524 (N_2524,N_2466,N_2432);
xor U2525 (N_2525,N_2473,N_2458);
nor U2526 (N_2526,N_2416,N_2414);
nor U2527 (N_2527,N_2484,N_2495);
or U2528 (N_2528,N_2497,N_2445);
nand U2529 (N_2529,N_2465,N_2485);
and U2530 (N_2530,N_2407,N_2442);
nand U2531 (N_2531,N_2402,N_2438);
nor U2532 (N_2532,N_2420,N_2428);
and U2533 (N_2533,N_2493,N_2415);
and U2534 (N_2534,N_2403,N_2480);
nor U2535 (N_2535,N_2472,N_2460);
nand U2536 (N_2536,N_2470,N_2440);
and U2537 (N_2537,N_2492,N_2496);
nand U2538 (N_2538,N_2486,N_2434);
xnor U2539 (N_2539,N_2476,N_2439);
nand U2540 (N_2540,N_2401,N_2448);
or U2541 (N_2541,N_2419,N_2477);
nor U2542 (N_2542,N_2446,N_2408);
xor U2543 (N_2543,N_2433,N_2498);
xor U2544 (N_2544,N_2418,N_2459);
and U2545 (N_2545,N_2427,N_2462);
or U2546 (N_2546,N_2426,N_2455);
or U2547 (N_2547,N_2491,N_2449);
xor U2548 (N_2548,N_2482,N_2410);
xor U2549 (N_2549,N_2405,N_2461);
xor U2550 (N_2550,N_2456,N_2441);
nor U2551 (N_2551,N_2429,N_2451);
nor U2552 (N_2552,N_2443,N_2494);
nor U2553 (N_2553,N_2494,N_2460);
or U2554 (N_2554,N_2431,N_2451);
nor U2555 (N_2555,N_2412,N_2459);
or U2556 (N_2556,N_2411,N_2445);
xor U2557 (N_2557,N_2405,N_2485);
or U2558 (N_2558,N_2402,N_2428);
and U2559 (N_2559,N_2448,N_2414);
and U2560 (N_2560,N_2451,N_2476);
nand U2561 (N_2561,N_2497,N_2494);
nor U2562 (N_2562,N_2486,N_2470);
nor U2563 (N_2563,N_2499,N_2466);
and U2564 (N_2564,N_2461,N_2451);
or U2565 (N_2565,N_2429,N_2447);
or U2566 (N_2566,N_2450,N_2451);
nand U2567 (N_2567,N_2462,N_2475);
nor U2568 (N_2568,N_2418,N_2454);
nand U2569 (N_2569,N_2440,N_2463);
nor U2570 (N_2570,N_2412,N_2496);
and U2571 (N_2571,N_2454,N_2461);
xor U2572 (N_2572,N_2423,N_2470);
or U2573 (N_2573,N_2403,N_2482);
and U2574 (N_2574,N_2458,N_2411);
and U2575 (N_2575,N_2474,N_2495);
xor U2576 (N_2576,N_2431,N_2429);
and U2577 (N_2577,N_2444,N_2416);
nand U2578 (N_2578,N_2472,N_2490);
and U2579 (N_2579,N_2485,N_2464);
and U2580 (N_2580,N_2476,N_2412);
nand U2581 (N_2581,N_2492,N_2409);
and U2582 (N_2582,N_2433,N_2447);
nor U2583 (N_2583,N_2478,N_2458);
or U2584 (N_2584,N_2488,N_2458);
or U2585 (N_2585,N_2489,N_2490);
or U2586 (N_2586,N_2439,N_2424);
and U2587 (N_2587,N_2436,N_2448);
or U2588 (N_2588,N_2420,N_2436);
nor U2589 (N_2589,N_2409,N_2429);
or U2590 (N_2590,N_2497,N_2409);
or U2591 (N_2591,N_2422,N_2426);
nor U2592 (N_2592,N_2499,N_2467);
and U2593 (N_2593,N_2430,N_2460);
nand U2594 (N_2594,N_2451,N_2403);
and U2595 (N_2595,N_2476,N_2459);
nor U2596 (N_2596,N_2420,N_2480);
nand U2597 (N_2597,N_2447,N_2424);
nand U2598 (N_2598,N_2440,N_2491);
nand U2599 (N_2599,N_2460,N_2412);
or U2600 (N_2600,N_2553,N_2589);
and U2601 (N_2601,N_2504,N_2544);
nand U2602 (N_2602,N_2575,N_2555);
nor U2603 (N_2603,N_2551,N_2523);
nor U2604 (N_2604,N_2583,N_2581);
nor U2605 (N_2605,N_2570,N_2522);
or U2606 (N_2606,N_2543,N_2516);
xor U2607 (N_2607,N_2509,N_2538);
or U2608 (N_2608,N_2530,N_2500);
xor U2609 (N_2609,N_2556,N_2532);
and U2610 (N_2610,N_2557,N_2592);
nand U2611 (N_2611,N_2528,N_2537);
and U2612 (N_2612,N_2579,N_2565);
and U2613 (N_2613,N_2534,N_2529);
or U2614 (N_2614,N_2513,N_2518);
nand U2615 (N_2615,N_2547,N_2560);
nand U2616 (N_2616,N_2584,N_2587);
nand U2617 (N_2617,N_2514,N_2545);
and U2618 (N_2618,N_2519,N_2503);
and U2619 (N_2619,N_2595,N_2566);
nor U2620 (N_2620,N_2505,N_2586);
nand U2621 (N_2621,N_2520,N_2517);
nand U2622 (N_2622,N_2533,N_2502);
nand U2623 (N_2623,N_2541,N_2552);
nand U2624 (N_2624,N_2550,N_2524);
nor U2625 (N_2625,N_2563,N_2507);
or U2626 (N_2626,N_2588,N_2549);
xnor U2627 (N_2627,N_2527,N_2511);
or U2628 (N_2628,N_2572,N_2510);
and U2629 (N_2629,N_2578,N_2594);
and U2630 (N_2630,N_2546,N_2512);
or U2631 (N_2631,N_2568,N_2508);
or U2632 (N_2632,N_2580,N_2536);
xnor U2633 (N_2633,N_2599,N_2597);
or U2634 (N_2634,N_2559,N_2561);
nand U2635 (N_2635,N_2596,N_2554);
and U2636 (N_2636,N_2535,N_2573);
and U2637 (N_2637,N_2562,N_2593);
and U2638 (N_2638,N_2576,N_2540);
nand U2639 (N_2639,N_2585,N_2539);
nor U2640 (N_2640,N_2569,N_2567);
and U2641 (N_2641,N_2574,N_2582);
nor U2642 (N_2642,N_2577,N_2591);
nand U2643 (N_2643,N_2526,N_2531);
or U2644 (N_2644,N_2506,N_2598);
and U2645 (N_2645,N_2558,N_2521);
xnor U2646 (N_2646,N_2515,N_2542);
xor U2647 (N_2647,N_2548,N_2590);
and U2648 (N_2648,N_2501,N_2564);
nor U2649 (N_2649,N_2571,N_2525);
nor U2650 (N_2650,N_2560,N_2577);
xor U2651 (N_2651,N_2598,N_2582);
nand U2652 (N_2652,N_2561,N_2580);
nor U2653 (N_2653,N_2529,N_2509);
nand U2654 (N_2654,N_2508,N_2530);
or U2655 (N_2655,N_2557,N_2502);
nand U2656 (N_2656,N_2598,N_2555);
nand U2657 (N_2657,N_2577,N_2554);
nor U2658 (N_2658,N_2528,N_2544);
nand U2659 (N_2659,N_2583,N_2594);
or U2660 (N_2660,N_2532,N_2585);
xor U2661 (N_2661,N_2510,N_2533);
nand U2662 (N_2662,N_2546,N_2552);
and U2663 (N_2663,N_2545,N_2527);
or U2664 (N_2664,N_2569,N_2565);
nand U2665 (N_2665,N_2507,N_2558);
or U2666 (N_2666,N_2538,N_2521);
nor U2667 (N_2667,N_2569,N_2502);
and U2668 (N_2668,N_2530,N_2538);
xnor U2669 (N_2669,N_2557,N_2505);
or U2670 (N_2670,N_2572,N_2518);
nor U2671 (N_2671,N_2586,N_2580);
or U2672 (N_2672,N_2546,N_2533);
nor U2673 (N_2673,N_2546,N_2562);
nor U2674 (N_2674,N_2527,N_2531);
nor U2675 (N_2675,N_2521,N_2512);
nor U2676 (N_2676,N_2520,N_2540);
or U2677 (N_2677,N_2549,N_2593);
nand U2678 (N_2678,N_2544,N_2568);
nor U2679 (N_2679,N_2579,N_2500);
nand U2680 (N_2680,N_2531,N_2540);
and U2681 (N_2681,N_2545,N_2561);
nor U2682 (N_2682,N_2510,N_2526);
and U2683 (N_2683,N_2533,N_2544);
nor U2684 (N_2684,N_2530,N_2571);
nand U2685 (N_2685,N_2581,N_2516);
nor U2686 (N_2686,N_2539,N_2587);
nor U2687 (N_2687,N_2562,N_2594);
nor U2688 (N_2688,N_2503,N_2539);
nand U2689 (N_2689,N_2539,N_2591);
nor U2690 (N_2690,N_2557,N_2595);
nor U2691 (N_2691,N_2574,N_2503);
or U2692 (N_2692,N_2576,N_2596);
nor U2693 (N_2693,N_2552,N_2585);
and U2694 (N_2694,N_2567,N_2599);
nor U2695 (N_2695,N_2530,N_2562);
nor U2696 (N_2696,N_2561,N_2527);
and U2697 (N_2697,N_2501,N_2540);
nor U2698 (N_2698,N_2594,N_2596);
or U2699 (N_2699,N_2563,N_2588);
or U2700 (N_2700,N_2648,N_2677);
nand U2701 (N_2701,N_2641,N_2653);
nor U2702 (N_2702,N_2628,N_2682);
and U2703 (N_2703,N_2694,N_2614);
or U2704 (N_2704,N_2674,N_2671);
or U2705 (N_2705,N_2600,N_2611);
nand U2706 (N_2706,N_2607,N_2623);
nor U2707 (N_2707,N_2602,N_2624);
nand U2708 (N_2708,N_2657,N_2620);
and U2709 (N_2709,N_2660,N_2689);
nor U2710 (N_2710,N_2634,N_2696);
xor U2711 (N_2711,N_2687,N_2629);
or U2712 (N_2712,N_2627,N_2678);
nand U2713 (N_2713,N_2681,N_2655);
or U2714 (N_2714,N_2699,N_2659);
nand U2715 (N_2715,N_2669,N_2613);
nand U2716 (N_2716,N_2639,N_2668);
nor U2717 (N_2717,N_2680,N_2665);
and U2718 (N_2718,N_2606,N_2676);
nand U2719 (N_2719,N_2612,N_2632);
or U2720 (N_2720,N_2650,N_2615);
nand U2721 (N_2721,N_2636,N_2652);
or U2722 (N_2722,N_2651,N_2656);
nand U2723 (N_2723,N_2686,N_2630);
or U2724 (N_2724,N_2617,N_2643);
nor U2725 (N_2725,N_2626,N_2667);
or U2726 (N_2726,N_2679,N_2645);
and U2727 (N_2727,N_2610,N_2697);
nand U2728 (N_2728,N_2685,N_2640);
nor U2729 (N_2729,N_2663,N_2601);
xnor U2730 (N_2730,N_2688,N_2608);
nand U2731 (N_2731,N_2642,N_2684);
and U2732 (N_2732,N_2619,N_2662);
nand U2733 (N_2733,N_2654,N_2633);
nand U2734 (N_2734,N_2621,N_2693);
nand U2735 (N_2735,N_2695,N_2649);
nor U2736 (N_2736,N_2618,N_2646);
or U2737 (N_2737,N_2622,N_2664);
or U2738 (N_2738,N_2683,N_2604);
or U2739 (N_2739,N_2661,N_2609);
or U2740 (N_2740,N_2675,N_2638);
and U2741 (N_2741,N_2625,N_2692);
or U2742 (N_2742,N_2666,N_2605);
nand U2743 (N_2743,N_2616,N_2672);
or U2744 (N_2744,N_2670,N_2691);
and U2745 (N_2745,N_2603,N_2658);
and U2746 (N_2746,N_2647,N_2644);
and U2747 (N_2747,N_2637,N_2631);
nor U2748 (N_2748,N_2690,N_2698);
nand U2749 (N_2749,N_2635,N_2673);
or U2750 (N_2750,N_2641,N_2658);
and U2751 (N_2751,N_2648,N_2637);
nor U2752 (N_2752,N_2668,N_2672);
nor U2753 (N_2753,N_2678,N_2605);
nor U2754 (N_2754,N_2679,N_2695);
and U2755 (N_2755,N_2618,N_2637);
and U2756 (N_2756,N_2611,N_2610);
nand U2757 (N_2757,N_2607,N_2626);
xor U2758 (N_2758,N_2653,N_2688);
nor U2759 (N_2759,N_2645,N_2632);
xnor U2760 (N_2760,N_2656,N_2638);
or U2761 (N_2761,N_2658,N_2642);
and U2762 (N_2762,N_2682,N_2699);
or U2763 (N_2763,N_2659,N_2672);
xnor U2764 (N_2764,N_2669,N_2643);
or U2765 (N_2765,N_2650,N_2697);
nor U2766 (N_2766,N_2674,N_2676);
or U2767 (N_2767,N_2694,N_2679);
nor U2768 (N_2768,N_2655,N_2627);
nor U2769 (N_2769,N_2600,N_2610);
and U2770 (N_2770,N_2681,N_2619);
nand U2771 (N_2771,N_2650,N_2618);
or U2772 (N_2772,N_2672,N_2638);
or U2773 (N_2773,N_2670,N_2604);
xnor U2774 (N_2774,N_2615,N_2626);
or U2775 (N_2775,N_2696,N_2690);
or U2776 (N_2776,N_2684,N_2696);
and U2777 (N_2777,N_2680,N_2648);
nand U2778 (N_2778,N_2670,N_2615);
nor U2779 (N_2779,N_2671,N_2638);
xnor U2780 (N_2780,N_2613,N_2654);
nand U2781 (N_2781,N_2611,N_2631);
nor U2782 (N_2782,N_2666,N_2604);
and U2783 (N_2783,N_2674,N_2687);
nand U2784 (N_2784,N_2667,N_2671);
and U2785 (N_2785,N_2670,N_2642);
xor U2786 (N_2786,N_2698,N_2670);
or U2787 (N_2787,N_2668,N_2634);
nand U2788 (N_2788,N_2634,N_2651);
nand U2789 (N_2789,N_2659,N_2635);
nand U2790 (N_2790,N_2630,N_2633);
or U2791 (N_2791,N_2604,N_2653);
and U2792 (N_2792,N_2680,N_2670);
nor U2793 (N_2793,N_2604,N_2615);
xor U2794 (N_2794,N_2638,N_2642);
nand U2795 (N_2795,N_2657,N_2624);
nor U2796 (N_2796,N_2658,N_2650);
nand U2797 (N_2797,N_2692,N_2685);
nor U2798 (N_2798,N_2663,N_2699);
nand U2799 (N_2799,N_2688,N_2619);
nor U2800 (N_2800,N_2704,N_2745);
nor U2801 (N_2801,N_2790,N_2768);
nand U2802 (N_2802,N_2744,N_2736);
or U2803 (N_2803,N_2718,N_2750);
or U2804 (N_2804,N_2735,N_2746);
xnor U2805 (N_2805,N_2751,N_2723);
and U2806 (N_2806,N_2795,N_2726);
nand U2807 (N_2807,N_2743,N_2793);
nor U2808 (N_2808,N_2703,N_2724);
and U2809 (N_2809,N_2774,N_2758);
nor U2810 (N_2810,N_2738,N_2787);
nor U2811 (N_2811,N_2717,N_2709);
and U2812 (N_2812,N_2792,N_2765);
nor U2813 (N_2813,N_2759,N_2728);
and U2814 (N_2814,N_2782,N_2729);
nor U2815 (N_2815,N_2770,N_2741);
nor U2816 (N_2816,N_2720,N_2712);
and U2817 (N_2817,N_2791,N_2776);
and U2818 (N_2818,N_2798,N_2727);
nand U2819 (N_2819,N_2749,N_2702);
and U2820 (N_2820,N_2756,N_2714);
or U2821 (N_2821,N_2761,N_2757);
and U2822 (N_2822,N_2760,N_2732);
nor U2823 (N_2823,N_2769,N_2773);
and U2824 (N_2824,N_2713,N_2762);
nor U2825 (N_2825,N_2734,N_2710);
or U2826 (N_2826,N_2772,N_2715);
or U2827 (N_2827,N_2786,N_2747);
or U2828 (N_2828,N_2767,N_2708);
nand U2829 (N_2829,N_2771,N_2733);
or U2830 (N_2830,N_2785,N_2722);
nor U2831 (N_2831,N_2706,N_2783);
nand U2832 (N_2832,N_2755,N_2766);
nor U2833 (N_2833,N_2777,N_2796);
nand U2834 (N_2834,N_2753,N_2797);
nand U2835 (N_2835,N_2778,N_2799);
nand U2836 (N_2836,N_2737,N_2763);
and U2837 (N_2837,N_2784,N_2731);
nor U2838 (N_2838,N_2779,N_2707);
or U2839 (N_2839,N_2730,N_2719);
or U2840 (N_2840,N_2721,N_2789);
nor U2841 (N_2841,N_2711,N_2794);
nand U2842 (N_2842,N_2781,N_2775);
nor U2843 (N_2843,N_2752,N_2705);
nor U2844 (N_2844,N_2748,N_2754);
or U2845 (N_2845,N_2788,N_2740);
and U2846 (N_2846,N_2716,N_2725);
nand U2847 (N_2847,N_2764,N_2780);
nor U2848 (N_2848,N_2701,N_2742);
nand U2849 (N_2849,N_2700,N_2739);
nand U2850 (N_2850,N_2711,N_2753);
or U2851 (N_2851,N_2768,N_2712);
nor U2852 (N_2852,N_2724,N_2754);
or U2853 (N_2853,N_2788,N_2745);
xor U2854 (N_2854,N_2744,N_2780);
nand U2855 (N_2855,N_2721,N_2706);
and U2856 (N_2856,N_2722,N_2724);
nor U2857 (N_2857,N_2730,N_2785);
nand U2858 (N_2858,N_2719,N_2780);
and U2859 (N_2859,N_2741,N_2788);
and U2860 (N_2860,N_2744,N_2786);
nand U2861 (N_2861,N_2765,N_2762);
and U2862 (N_2862,N_2776,N_2725);
and U2863 (N_2863,N_2763,N_2726);
xnor U2864 (N_2864,N_2711,N_2743);
or U2865 (N_2865,N_2797,N_2732);
and U2866 (N_2866,N_2787,N_2791);
and U2867 (N_2867,N_2762,N_2740);
nand U2868 (N_2868,N_2748,N_2776);
nand U2869 (N_2869,N_2766,N_2738);
or U2870 (N_2870,N_2765,N_2793);
nor U2871 (N_2871,N_2733,N_2784);
and U2872 (N_2872,N_2707,N_2784);
nor U2873 (N_2873,N_2732,N_2757);
and U2874 (N_2874,N_2747,N_2796);
nand U2875 (N_2875,N_2776,N_2710);
xor U2876 (N_2876,N_2723,N_2757);
nand U2877 (N_2877,N_2795,N_2754);
nor U2878 (N_2878,N_2736,N_2729);
xnor U2879 (N_2879,N_2786,N_2731);
xnor U2880 (N_2880,N_2797,N_2750);
nor U2881 (N_2881,N_2758,N_2752);
and U2882 (N_2882,N_2738,N_2772);
nor U2883 (N_2883,N_2702,N_2771);
and U2884 (N_2884,N_2708,N_2794);
nand U2885 (N_2885,N_2767,N_2732);
xor U2886 (N_2886,N_2724,N_2705);
nand U2887 (N_2887,N_2773,N_2713);
or U2888 (N_2888,N_2722,N_2735);
nand U2889 (N_2889,N_2792,N_2752);
nand U2890 (N_2890,N_2714,N_2767);
and U2891 (N_2891,N_2718,N_2702);
nand U2892 (N_2892,N_2789,N_2705);
xor U2893 (N_2893,N_2760,N_2704);
nor U2894 (N_2894,N_2711,N_2723);
xnor U2895 (N_2895,N_2758,N_2785);
and U2896 (N_2896,N_2739,N_2776);
and U2897 (N_2897,N_2752,N_2769);
xor U2898 (N_2898,N_2774,N_2776);
or U2899 (N_2899,N_2743,N_2746);
nand U2900 (N_2900,N_2827,N_2895);
or U2901 (N_2901,N_2828,N_2889);
and U2902 (N_2902,N_2886,N_2812);
nor U2903 (N_2903,N_2804,N_2854);
nand U2904 (N_2904,N_2803,N_2808);
or U2905 (N_2905,N_2851,N_2826);
nand U2906 (N_2906,N_2845,N_2834);
and U2907 (N_2907,N_2818,N_2801);
or U2908 (N_2908,N_2825,N_2894);
nand U2909 (N_2909,N_2867,N_2836);
or U2910 (N_2910,N_2810,N_2800);
nand U2911 (N_2911,N_2870,N_2875);
and U2912 (N_2912,N_2863,N_2860);
or U2913 (N_2913,N_2823,N_2880);
and U2914 (N_2914,N_2855,N_2842);
nand U2915 (N_2915,N_2849,N_2848);
nor U2916 (N_2916,N_2853,N_2824);
nor U2917 (N_2917,N_2840,N_2852);
nor U2918 (N_2918,N_2832,N_2893);
xor U2919 (N_2919,N_2838,N_2887);
nor U2920 (N_2920,N_2865,N_2876);
and U2921 (N_2921,N_2819,N_2897);
or U2922 (N_2922,N_2878,N_2874);
nor U2923 (N_2923,N_2813,N_2806);
nand U2924 (N_2924,N_2861,N_2805);
nand U2925 (N_2925,N_2879,N_2837);
or U2926 (N_2926,N_2869,N_2817);
and U2927 (N_2927,N_2822,N_2857);
and U2928 (N_2928,N_2862,N_2866);
xor U2929 (N_2929,N_2884,N_2816);
or U2930 (N_2930,N_2882,N_2843);
nand U2931 (N_2931,N_2841,N_2871);
or U2932 (N_2932,N_2858,N_2891);
nand U2933 (N_2933,N_2821,N_2868);
nand U2934 (N_2934,N_2864,N_2859);
or U2935 (N_2935,N_2839,N_2830);
and U2936 (N_2936,N_2835,N_2899);
nand U2937 (N_2937,N_2807,N_2890);
nor U2938 (N_2938,N_2829,N_2885);
nand U2939 (N_2939,N_2814,N_2850);
nand U2940 (N_2940,N_2844,N_2802);
nor U2941 (N_2941,N_2809,N_2847);
nor U2942 (N_2942,N_2831,N_2877);
nand U2943 (N_2943,N_2815,N_2883);
nor U2944 (N_2944,N_2896,N_2888);
nor U2945 (N_2945,N_2873,N_2892);
or U2946 (N_2946,N_2820,N_2856);
or U2947 (N_2947,N_2846,N_2811);
xnor U2948 (N_2948,N_2833,N_2898);
xnor U2949 (N_2949,N_2872,N_2881);
or U2950 (N_2950,N_2899,N_2855);
and U2951 (N_2951,N_2843,N_2834);
xnor U2952 (N_2952,N_2844,N_2800);
nand U2953 (N_2953,N_2896,N_2835);
nor U2954 (N_2954,N_2887,N_2860);
and U2955 (N_2955,N_2886,N_2880);
and U2956 (N_2956,N_2828,N_2844);
nand U2957 (N_2957,N_2816,N_2845);
nor U2958 (N_2958,N_2820,N_2872);
nand U2959 (N_2959,N_2835,N_2887);
and U2960 (N_2960,N_2838,N_2872);
nand U2961 (N_2961,N_2891,N_2837);
nor U2962 (N_2962,N_2800,N_2808);
or U2963 (N_2963,N_2804,N_2857);
and U2964 (N_2964,N_2856,N_2882);
nand U2965 (N_2965,N_2829,N_2852);
or U2966 (N_2966,N_2807,N_2878);
nor U2967 (N_2967,N_2869,N_2810);
and U2968 (N_2968,N_2875,N_2846);
nand U2969 (N_2969,N_2876,N_2856);
or U2970 (N_2970,N_2872,N_2888);
nor U2971 (N_2971,N_2816,N_2873);
nand U2972 (N_2972,N_2856,N_2883);
or U2973 (N_2973,N_2824,N_2864);
nand U2974 (N_2974,N_2838,N_2868);
or U2975 (N_2975,N_2898,N_2858);
or U2976 (N_2976,N_2812,N_2815);
nand U2977 (N_2977,N_2874,N_2842);
nand U2978 (N_2978,N_2805,N_2812);
and U2979 (N_2979,N_2838,N_2840);
or U2980 (N_2980,N_2823,N_2841);
nor U2981 (N_2981,N_2850,N_2801);
or U2982 (N_2982,N_2878,N_2833);
nor U2983 (N_2983,N_2805,N_2884);
nor U2984 (N_2984,N_2868,N_2872);
nor U2985 (N_2985,N_2879,N_2832);
and U2986 (N_2986,N_2859,N_2838);
xnor U2987 (N_2987,N_2894,N_2867);
and U2988 (N_2988,N_2822,N_2898);
and U2989 (N_2989,N_2812,N_2844);
and U2990 (N_2990,N_2857,N_2843);
nand U2991 (N_2991,N_2850,N_2891);
nor U2992 (N_2992,N_2853,N_2825);
nand U2993 (N_2993,N_2866,N_2852);
or U2994 (N_2994,N_2848,N_2804);
or U2995 (N_2995,N_2856,N_2840);
nand U2996 (N_2996,N_2835,N_2814);
nor U2997 (N_2997,N_2808,N_2813);
or U2998 (N_2998,N_2822,N_2860);
and U2999 (N_2999,N_2864,N_2885);
nor UO_0 (O_0,N_2929,N_2966);
or UO_1 (O_1,N_2968,N_2926);
or UO_2 (O_2,N_2913,N_2969);
and UO_3 (O_3,N_2943,N_2902);
or UO_4 (O_4,N_2952,N_2935);
nand UO_5 (O_5,N_2936,N_2965);
nor UO_6 (O_6,N_2993,N_2971);
nand UO_7 (O_7,N_2951,N_2995);
and UO_8 (O_8,N_2991,N_2958);
nor UO_9 (O_9,N_2915,N_2973);
or UO_10 (O_10,N_2927,N_2959);
nand UO_11 (O_11,N_2997,N_2950);
and UO_12 (O_12,N_2941,N_2978);
or UO_13 (O_13,N_2904,N_2908);
nand UO_14 (O_14,N_2949,N_2985);
nor UO_15 (O_15,N_2903,N_2901);
or UO_16 (O_16,N_2940,N_2944);
nand UO_17 (O_17,N_2933,N_2994);
nand UO_18 (O_18,N_2911,N_2960);
or UO_19 (O_19,N_2924,N_2980);
and UO_20 (O_20,N_2976,N_2919);
nor UO_21 (O_21,N_2923,N_2999);
and UO_22 (O_22,N_2914,N_2916);
nand UO_23 (O_23,N_2922,N_2931);
nand UO_24 (O_24,N_2975,N_2942);
or UO_25 (O_25,N_2930,N_2945);
and UO_26 (O_26,N_2961,N_2998);
xnor UO_27 (O_27,N_2939,N_2964);
nand UO_28 (O_28,N_2990,N_2909);
nand UO_29 (O_29,N_2928,N_2967);
nor UO_30 (O_30,N_2912,N_2986);
nand UO_31 (O_31,N_2925,N_2948);
and UO_32 (O_32,N_2970,N_2979);
nor UO_33 (O_33,N_2937,N_2918);
or UO_34 (O_34,N_2996,N_2947);
nand UO_35 (O_35,N_2963,N_2988);
nor UO_36 (O_36,N_2955,N_2932);
nor UO_37 (O_37,N_2921,N_2954);
nor UO_38 (O_38,N_2974,N_2920);
or UO_39 (O_39,N_2962,N_2938);
or UO_40 (O_40,N_2905,N_2917);
nand UO_41 (O_41,N_2984,N_2907);
nor UO_42 (O_42,N_2953,N_2946);
or UO_43 (O_43,N_2987,N_2910);
nor UO_44 (O_44,N_2972,N_2982);
or UO_45 (O_45,N_2956,N_2977);
or UO_46 (O_46,N_2957,N_2989);
xnor UO_47 (O_47,N_2934,N_2983);
nand UO_48 (O_48,N_2900,N_2981);
and UO_49 (O_49,N_2906,N_2992);
and UO_50 (O_50,N_2963,N_2987);
xnor UO_51 (O_51,N_2964,N_2928);
nand UO_52 (O_52,N_2999,N_2924);
nand UO_53 (O_53,N_2904,N_2923);
nor UO_54 (O_54,N_2989,N_2907);
or UO_55 (O_55,N_2990,N_2913);
nor UO_56 (O_56,N_2926,N_2937);
and UO_57 (O_57,N_2950,N_2970);
or UO_58 (O_58,N_2922,N_2997);
xor UO_59 (O_59,N_2949,N_2993);
nor UO_60 (O_60,N_2912,N_2907);
or UO_61 (O_61,N_2917,N_2937);
and UO_62 (O_62,N_2942,N_2951);
nand UO_63 (O_63,N_2907,N_2929);
and UO_64 (O_64,N_2947,N_2941);
and UO_65 (O_65,N_2956,N_2960);
nor UO_66 (O_66,N_2981,N_2966);
or UO_67 (O_67,N_2950,N_2930);
nor UO_68 (O_68,N_2903,N_2938);
xor UO_69 (O_69,N_2951,N_2991);
or UO_70 (O_70,N_2910,N_2990);
and UO_71 (O_71,N_2955,N_2945);
nor UO_72 (O_72,N_2905,N_2955);
nand UO_73 (O_73,N_2994,N_2928);
nor UO_74 (O_74,N_2917,N_2900);
nor UO_75 (O_75,N_2920,N_2912);
and UO_76 (O_76,N_2930,N_2979);
nand UO_77 (O_77,N_2986,N_2936);
nand UO_78 (O_78,N_2945,N_2971);
nor UO_79 (O_79,N_2923,N_2968);
nand UO_80 (O_80,N_2902,N_2983);
or UO_81 (O_81,N_2978,N_2997);
nor UO_82 (O_82,N_2910,N_2915);
nand UO_83 (O_83,N_2925,N_2969);
nand UO_84 (O_84,N_2995,N_2904);
nor UO_85 (O_85,N_2972,N_2991);
xor UO_86 (O_86,N_2935,N_2904);
or UO_87 (O_87,N_2972,N_2969);
and UO_88 (O_88,N_2993,N_2931);
nand UO_89 (O_89,N_2976,N_2997);
nor UO_90 (O_90,N_2924,N_2937);
nor UO_91 (O_91,N_2970,N_2985);
nor UO_92 (O_92,N_2954,N_2994);
nand UO_93 (O_93,N_2932,N_2964);
and UO_94 (O_94,N_2954,N_2975);
or UO_95 (O_95,N_2946,N_2902);
nand UO_96 (O_96,N_2979,N_2960);
or UO_97 (O_97,N_2959,N_2965);
nor UO_98 (O_98,N_2913,N_2987);
nor UO_99 (O_99,N_2999,N_2913);
xor UO_100 (O_100,N_2952,N_2922);
or UO_101 (O_101,N_2976,N_2961);
nor UO_102 (O_102,N_2993,N_2950);
nor UO_103 (O_103,N_2971,N_2989);
nand UO_104 (O_104,N_2909,N_2955);
or UO_105 (O_105,N_2926,N_2956);
nor UO_106 (O_106,N_2905,N_2950);
nor UO_107 (O_107,N_2996,N_2992);
nor UO_108 (O_108,N_2931,N_2978);
nor UO_109 (O_109,N_2912,N_2952);
or UO_110 (O_110,N_2954,N_2957);
nand UO_111 (O_111,N_2961,N_2944);
or UO_112 (O_112,N_2926,N_2985);
or UO_113 (O_113,N_2916,N_2970);
nand UO_114 (O_114,N_2954,N_2943);
nand UO_115 (O_115,N_2985,N_2938);
nand UO_116 (O_116,N_2984,N_2991);
and UO_117 (O_117,N_2933,N_2983);
or UO_118 (O_118,N_2941,N_2991);
and UO_119 (O_119,N_2953,N_2915);
nand UO_120 (O_120,N_2975,N_2918);
nand UO_121 (O_121,N_2987,N_2945);
and UO_122 (O_122,N_2966,N_2941);
or UO_123 (O_123,N_2968,N_2982);
and UO_124 (O_124,N_2913,N_2906);
or UO_125 (O_125,N_2906,N_2964);
or UO_126 (O_126,N_2931,N_2962);
and UO_127 (O_127,N_2984,N_2925);
nand UO_128 (O_128,N_2934,N_2917);
and UO_129 (O_129,N_2937,N_2964);
and UO_130 (O_130,N_2964,N_2990);
or UO_131 (O_131,N_2938,N_2934);
nor UO_132 (O_132,N_2900,N_2957);
or UO_133 (O_133,N_2916,N_2996);
nand UO_134 (O_134,N_2949,N_2921);
xnor UO_135 (O_135,N_2940,N_2947);
nor UO_136 (O_136,N_2937,N_2915);
nor UO_137 (O_137,N_2925,N_2964);
and UO_138 (O_138,N_2940,N_2950);
nor UO_139 (O_139,N_2970,N_2940);
nor UO_140 (O_140,N_2949,N_2989);
nor UO_141 (O_141,N_2978,N_2933);
and UO_142 (O_142,N_2902,N_2960);
nor UO_143 (O_143,N_2924,N_2982);
or UO_144 (O_144,N_2930,N_2927);
nand UO_145 (O_145,N_2952,N_2945);
nor UO_146 (O_146,N_2990,N_2945);
or UO_147 (O_147,N_2947,N_2911);
nand UO_148 (O_148,N_2984,N_2966);
and UO_149 (O_149,N_2916,N_2949);
nor UO_150 (O_150,N_2973,N_2974);
or UO_151 (O_151,N_2906,N_2983);
and UO_152 (O_152,N_2918,N_2947);
nand UO_153 (O_153,N_2931,N_2999);
or UO_154 (O_154,N_2958,N_2986);
and UO_155 (O_155,N_2960,N_2953);
nor UO_156 (O_156,N_2988,N_2974);
xnor UO_157 (O_157,N_2906,N_2940);
and UO_158 (O_158,N_2910,N_2992);
nor UO_159 (O_159,N_2918,N_2965);
and UO_160 (O_160,N_2943,N_2908);
nor UO_161 (O_161,N_2948,N_2904);
or UO_162 (O_162,N_2951,N_2997);
nand UO_163 (O_163,N_2951,N_2931);
or UO_164 (O_164,N_2915,N_2987);
or UO_165 (O_165,N_2998,N_2936);
and UO_166 (O_166,N_2931,N_2952);
or UO_167 (O_167,N_2979,N_2912);
and UO_168 (O_168,N_2957,N_2907);
nor UO_169 (O_169,N_2996,N_2981);
and UO_170 (O_170,N_2919,N_2912);
nor UO_171 (O_171,N_2955,N_2938);
or UO_172 (O_172,N_2930,N_2933);
nor UO_173 (O_173,N_2995,N_2964);
and UO_174 (O_174,N_2967,N_2994);
nor UO_175 (O_175,N_2917,N_2976);
or UO_176 (O_176,N_2938,N_2980);
and UO_177 (O_177,N_2959,N_2996);
nor UO_178 (O_178,N_2907,N_2941);
nand UO_179 (O_179,N_2983,N_2909);
nand UO_180 (O_180,N_2976,N_2952);
nand UO_181 (O_181,N_2976,N_2967);
or UO_182 (O_182,N_2910,N_2969);
nor UO_183 (O_183,N_2936,N_2902);
nand UO_184 (O_184,N_2975,N_2916);
nand UO_185 (O_185,N_2954,N_2937);
or UO_186 (O_186,N_2990,N_2950);
nand UO_187 (O_187,N_2936,N_2956);
or UO_188 (O_188,N_2961,N_2907);
or UO_189 (O_189,N_2916,N_2969);
nor UO_190 (O_190,N_2979,N_2995);
nor UO_191 (O_191,N_2978,N_2972);
or UO_192 (O_192,N_2943,N_2912);
xor UO_193 (O_193,N_2922,N_2988);
or UO_194 (O_194,N_2905,N_2999);
nand UO_195 (O_195,N_2906,N_2908);
nand UO_196 (O_196,N_2903,N_2993);
or UO_197 (O_197,N_2918,N_2922);
or UO_198 (O_198,N_2922,N_2901);
nor UO_199 (O_199,N_2999,N_2962);
and UO_200 (O_200,N_2936,N_2922);
nand UO_201 (O_201,N_2916,N_2955);
nor UO_202 (O_202,N_2908,N_2931);
xnor UO_203 (O_203,N_2968,N_2962);
nand UO_204 (O_204,N_2947,N_2912);
xnor UO_205 (O_205,N_2988,N_2909);
and UO_206 (O_206,N_2995,N_2909);
and UO_207 (O_207,N_2956,N_2975);
and UO_208 (O_208,N_2978,N_2990);
or UO_209 (O_209,N_2957,N_2942);
or UO_210 (O_210,N_2959,N_2931);
nand UO_211 (O_211,N_2979,N_2988);
or UO_212 (O_212,N_2967,N_2981);
nor UO_213 (O_213,N_2910,N_2949);
xnor UO_214 (O_214,N_2904,N_2911);
nand UO_215 (O_215,N_2977,N_2953);
or UO_216 (O_216,N_2995,N_2945);
nor UO_217 (O_217,N_2999,N_2992);
or UO_218 (O_218,N_2941,N_2934);
and UO_219 (O_219,N_2967,N_2939);
xnor UO_220 (O_220,N_2970,N_2943);
and UO_221 (O_221,N_2963,N_2911);
nor UO_222 (O_222,N_2914,N_2943);
and UO_223 (O_223,N_2964,N_2904);
nor UO_224 (O_224,N_2966,N_2976);
and UO_225 (O_225,N_2960,N_2978);
or UO_226 (O_226,N_2963,N_2919);
or UO_227 (O_227,N_2961,N_2992);
and UO_228 (O_228,N_2935,N_2940);
nor UO_229 (O_229,N_2968,N_2928);
or UO_230 (O_230,N_2914,N_2989);
nand UO_231 (O_231,N_2934,N_2975);
and UO_232 (O_232,N_2973,N_2991);
or UO_233 (O_233,N_2939,N_2968);
or UO_234 (O_234,N_2911,N_2983);
or UO_235 (O_235,N_2900,N_2979);
nor UO_236 (O_236,N_2990,N_2954);
nor UO_237 (O_237,N_2985,N_2942);
or UO_238 (O_238,N_2953,N_2976);
nand UO_239 (O_239,N_2924,N_2989);
nand UO_240 (O_240,N_2986,N_2940);
nor UO_241 (O_241,N_2914,N_2928);
nand UO_242 (O_242,N_2957,N_2903);
xor UO_243 (O_243,N_2952,N_2977);
xnor UO_244 (O_244,N_2963,N_2991);
nor UO_245 (O_245,N_2959,N_2991);
nor UO_246 (O_246,N_2949,N_2956);
xnor UO_247 (O_247,N_2924,N_2957);
nand UO_248 (O_248,N_2986,N_2920);
and UO_249 (O_249,N_2996,N_2915);
nor UO_250 (O_250,N_2969,N_2912);
nand UO_251 (O_251,N_2948,N_2977);
nand UO_252 (O_252,N_2904,N_2972);
and UO_253 (O_253,N_2980,N_2996);
nand UO_254 (O_254,N_2959,N_2930);
or UO_255 (O_255,N_2984,N_2943);
and UO_256 (O_256,N_2996,N_2973);
and UO_257 (O_257,N_2979,N_2951);
nor UO_258 (O_258,N_2926,N_2987);
and UO_259 (O_259,N_2969,N_2991);
nor UO_260 (O_260,N_2990,N_2936);
or UO_261 (O_261,N_2901,N_2952);
nor UO_262 (O_262,N_2992,N_2977);
nor UO_263 (O_263,N_2981,N_2968);
or UO_264 (O_264,N_2991,N_2927);
and UO_265 (O_265,N_2914,N_2922);
xnor UO_266 (O_266,N_2963,N_2966);
and UO_267 (O_267,N_2999,N_2969);
nand UO_268 (O_268,N_2999,N_2976);
and UO_269 (O_269,N_2973,N_2999);
or UO_270 (O_270,N_2996,N_2934);
nand UO_271 (O_271,N_2939,N_2993);
and UO_272 (O_272,N_2927,N_2990);
nand UO_273 (O_273,N_2900,N_2986);
nor UO_274 (O_274,N_2938,N_2945);
xnor UO_275 (O_275,N_2950,N_2943);
nor UO_276 (O_276,N_2968,N_2970);
and UO_277 (O_277,N_2998,N_2994);
nand UO_278 (O_278,N_2908,N_2990);
or UO_279 (O_279,N_2969,N_2980);
or UO_280 (O_280,N_2905,N_2942);
xnor UO_281 (O_281,N_2957,N_2960);
or UO_282 (O_282,N_2992,N_2989);
or UO_283 (O_283,N_2904,N_2938);
nand UO_284 (O_284,N_2903,N_2933);
nand UO_285 (O_285,N_2920,N_2959);
or UO_286 (O_286,N_2989,N_2970);
nand UO_287 (O_287,N_2989,N_2916);
or UO_288 (O_288,N_2962,N_2911);
and UO_289 (O_289,N_2958,N_2969);
and UO_290 (O_290,N_2926,N_2903);
and UO_291 (O_291,N_2924,N_2904);
nor UO_292 (O_292,N_2904,N_2925);
and UO_293 (O_293,N_2947,N_2973);
xnor UO_294 (O_294,N_2952,N_2998);
and UO_295 (O_295,N_2943,N_2919);
nor UO_296 (O_296,N_2929,N_2914);
nand UO_297 (O_297,N_2924,N_2987);
nand UO_298 (O_298,N_2978,N_2967);
nand UO_299 (O_299,N_2955,N_2985);
nor UO_300 (O_300,N_2990,N_2985);
and UO_301 (O_301,N_2943,N_2994);
nand UO_302 (O_302,N_2971,N_2972);
nor UO_303 (O_303,N_2996,N_2965);
or UO_304 (O_304,N_2961,N_2990);
or UO_305 (O_305,N_2901,N_2908);
nand UO_306 (O_306,N_2995,N_2940);
and UO_307 (O_307,N_2941,N_2953);
nor UO_308 (O_308,N_2923,N_2963);
nor UO_309 (O_309,N_2934,N_2982);
nand UO_310 (O_310,N_2973,N_2905);
and UO_311 (O_311,N_2900,N_2955);
nand UO_312 (O_312,N_2988,N_2991);
or UO_313 (O_313,N_2911,N_2915);
and UO_314 (O_314,N_2917,N_2943);
and UO_315 (O_315,N_2991,N_2926);
and UO_316 (O_316,N_2997,N_2963);
or UO_317 (O_317,N_2966,N_2905);
nor UO_318 (O_318,N_2964,N_2948);
or UO_319 (O_319,N_2946,N_2933);
and UO_320 (O_320,N_2946,N_2980);
or UO_321 (O_321,N_2959,N_2966);
nand UO_322 (O_322,N_2987,N_2949);
or UO_323 (O_323,N_2997,N_2931);
or UO_324 (O_324,N_2934,N_2946);
nor UO_325 (O_325,N_2993,N_2995);
nand UO_326 (O_326,N_2937,N_2910);
nand UO_327 (O_327,N_2976,N_2980);
and UO_328 (O_328,N_2905,N_2951);
nor UO_329 (O_329,N_2984,N_2953);
and UO_330 (O_330,N_2939,N_2991);
nor UO_331 (O_331,N_2954,N_2967);
and UO_332 (O_332,N_2918,N_2928);
and UO_333 (O_333,N_2929,N_2916);
nor UO_334 (O_334,N_2979,N_2925);
and UO_335 (O_335,N_2935,N_2930);
and UO_336 (O_336,N_2998,N_2980);
xnor UO_337 (O_337,N_2926,N_2965);
or UO_338 (O_338,N_2902,N_2918);
and UO_339 (O_339,N_2996,N_2907);
nand UO_340 (O_340,N_2981,N_2969);
nor UO_341 (O_341,N_2958,N_2968);
nor UO_342 (O_342,N_2925,N_2935);
or UO_343 (O_343,N_2970,N_2922);
nand UO_344 (O_344,N_2996,N_2942);
nand UO_345 (O_345,N_2969,N_2982);
nor UO_346 (O_346,N_2944,N_2977);
and UO_347 (O_347,N_2994,N_2957);
nor UO_348 (O_348,N_2954,N_2951);
xor UO_349 (O_349,N_2994,N_2903);
and UO_350 (O_350,N_2961,N_2983);
and UO_351 (O_351,N_2984,N_2988);
nor UO_352 (O_352,N_2901,N_2943);
nor UO_353 (O_353,N_2984,N_2967);
xnor UO_354 (O_354,N_2959,N_2921);
and UO_355 (O_355,N_2905,N_2968);
and UO_356 (O_356,N_2908,N_2989);
nand UO_357 (O_357,N_2973,N_2960);
and UO_358 (O_358,N_2914,N_2973);
xnor UO_359 (O_359,N_2951,N_2966);
or UO_360 (O_360,N_2974,N_2967);
and UO_361 (O_361,N_2973,N_2957);
nor UO_362 (O_362,N_2966,N_2910);
or UO_363 (O_363,N_2972,N_2934);
nor UO_364 (O_364,N_2912,N_2978);
nand UO_365 (O_365,N_2914,N_2921);
or UO_366 (O_366,N_2965,N_2982);
or UO_367 (O_367,N_2950,N_2918);
or UO_368 (O_368,N_2922,N_2905);
or UO_369 (O_369,N_2971,N_2929);
xor UO_370 (O_370,N_2985,N_2921);
nor UO_371 (O_371,N_2983,N_2946);
nand UO_372 (O_372,N_2945,N_2942);
nand UO_373 (O_373,N_2966,N_2940);
or UO_374 (O_374,N_2997,N_2920);
or UO_375 (O_375,N_2944,N_2929);
nor UO_376 (O_376,N_2989,N_2968);
xor UO_377 (O_377,N_2957,N_2970);
nand UO_378 (O_378,N_2970,N_2927);
and UO_379 (O_379,N_2986,N_2929);
nor UO_380 (O_380,N_2999,N_2986);
nor UO_381 (O_381,N_2992,N_2902);
and UO_382 (O_382,N_2929,N_2923);
and UO_383 (O_383,N_2945,N_2985);
or UO_384 (O_384,N_2927,N_2941);
and UO_385 (O_385,N_2969,N_2938);
nand UO_386 (O_386,N_2972,N_2996);
nand UO_387 (O_387,N_2935,N_2957);
or UO_388 (O_388,N_2914,N_2959);
or UO_389 (O_389,N_2930,N_2912);
nor UO_390 (O_390,N_2977,N_2990);
nand UO_391 (O_391,N_2975,N_2914);
xor UO_392 (O_392,N_2944,N_2913);
and UO_393 (O_393,N_2957,N_2963);
and UO_394 (O_394,N_2938,N_2942);
and UO_395 (O_395,N_2914,N_2946);
nand UO_396 (O_396,N_2976,N_2932);
nor UO_397 (O_397,N_2968,N_2977);
or UO_398 (O_398,N_2967,N_2902);
or UO_399 (O_399,N_2915,N_2960);
nor UO_400 (O_400,N_2980,N_2913);
nor UO_401 (O_401,N_2903,N_2995);
or UO_402 (O_402,N_2930,N_2971);
nand UO_403 (O_403,N_2913,N_2967);
nor UO_404 (O_404,N_2952,N_2908);
or UO_405 (O_405,N_2931,N_2902);
and UO_406 (O_406,N_2939,N_2982);
and UO_407 (O_407,N_2913,N_2989);
nand UO_408 (O_408,N_2919,N_2982);
and UO_409 (O_409,N_2932,N_2915);
nor UO_410 (O_410,N_2915,N_2978);
nor UO_411 (O_411,N_2965,N_2902);
nand UO_412 (O_412,N_2942,N_2920);
nand UO_413 (O_413,N_2910,N_2944);
nand UO_414 (O_414,N_2954,N_2953);
nor UO_415 (O_415,N_2997,N_2914);
and UO_416 (O_416,N_2928,N_2936);
or UO_417 (O_417,N_2982,N_2989);
and UO_418 (O_418,N_2972,N_2903);
or UO_419 (O_419,N_2953,N_2963);
nand UO_420 (O_420,N_2961,N_2901);
nand UO_421 (O_421,N_2994,N_2997);
nand UO_422 (O_422,N_2948,N_2933);
nor UO_423 (O_423,N_2976,N_2947);
and UO_424 (O_424,N_2954,N_2956);
and UO_425 (O_425,N_2909,N_2993);
nor UO_426 (O_426,N_2944,N_2916);
or UO_427 (O_427,N_2995,N_2976);
and UO_428 (O_428,N_2993,N_2953);
nor UO_429 (O_429,N_2971,N_2938);
nor UO_430 (O_430,N_2912,N_2939);
and UO_431 (O_431,N_2961,N_2957);
and UO_432 (O_432,N_2935,N_2915);
nor UO_433 (O_433,N_2914,N_2925);
or UO_434 (O_434,N_2928,N_2990);
xnor UO_435 (O_435,N_2974,N_2997);
nand UO_436 (O_436,N_2951,N_2937);
or UO_437 (O_437,N_2983,N_2951);
nand UO_438 (O_438,N_2928,N_2980);
xnor UO_439 (O_439,N_2966,N_2973);
and UO_440 (O_440,N_2904,N_2961);
nor UO_441 (O_441,N_2950,N_2969);
nor UO_442 (O_442,N_2951,N_2986);
or UO_443 (O_443,N_2960,N_2926);
and UO_444 (O_444,N_2981,N_2992);
xor UO_445 (O_445,N_2959,N_2964);
nand UO_446 (O_446,N_2962,N_2997);
nand UO_447 (O_447,N_2912,N_2950);
nand UO_448 (O_448,N_2942,N_2915);
and UO_449 (O_449,N_2997,N_2993);
nand UO_450 (O_450,N_2980,N_2912);
nor UO_451 (O_451,N_2931,N_2976);
nor UO_452 (O_452,N_2959,N_2958);
xnor UO_453 (O_453,N_2963,N_2999);
or UO_454 (O_454,N_2945,N_2989);
nor UO_455 (O_455,N_2908,N_2994);
and UO_456 (O_456,N_2903,N_2999);
xor UO_457 (O_457,N_2987,N_2908);
and UO_458 (O_458,N_2959,N_2995);
nor UO_459 (O_459,N_2980,N_2974);
nor UO_460 (O_460,N_2934,N_2995);
nor UO_461 (O_461,N_2909,N_2967);
and UO_462 (O_462,N_2936,N_2978);
xnor UO_463 (O_463,N_2936,N_2989);
nor UO_464 (O_464,N_2923,N_2997);
nor UO_465 (O_465,N_2984,N_2938);
or UO_466 (O_466,N_2951,N_2920);
nor UO_467 (O_467,N_2941,N_2999);
and UO_468 (O_468,N_2941,N_2948);
nor UO_469 (O_469,N_2917,N_2985);
and UO_470 (O_470,N_2918,N_2911);
and UO_471 (O_471,N_2996,N_2937);
nand UO_472 (O_472,N_2915,N_2958);
nor UO_473 (O_473,N_2981,N_2933);
or UO_474 (O_474,N_2931,N_2929);
xnor UO_475 (O_475,N_2993,N_2990);
xor UO_476 (O_476,N_2994,N_2932);
and UO_477 (O_477,N_2998,N_2940);
nand UO_478 (O_478,N_2969,N_2915);
nor UO_479 (O_479,N_2943,N_2987);
nand UO_480 (O_480,N_2908,N_2950);
and UO_481 (O_481,N_2972,N_2917);
nand UO_482 (O_482,N_2937,N_2907);
and UO_483 (O_483,N_2959,N_2972);
or UO_484 (O_484,N_2979,N_2905);
xor UO_485 (O_485,N_2925,N_2906);
xor UO_486 (O_486,N_2937,N_2919);
xnor UO_487 (O_487,N_2919,N_2964);
and UO_488 (O_488,N_2910,N_2967);
and UO_489 (O_489,N_2952,N_2926);
or UO_490 (O_490,N_2967,N_2972);
or UO_491 (O_491,N_2934,N_2961);
or UO_492 (O_492,N_2959,N_2939);
nand UO_493 (O_493,N_2984,N_2909);
and UO_494 (O_494,N_2962,N_2958);
or UO_495 (O_495,N_2970,N_2946);
and UO_496 (O_496,N_2984,N_2904);
or UO_497 (O_497,N_2936,N_2958);
and UO_498 (O_498,N_2900,N_2949);
and UO_499 (O_499,N_2922,N_2917);
endmodule