module basic_1000_10000_1500_2_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5004,N_5005,N_5006,N_5007,N_5008,N_5011,N_5012,N_5014,N_5015,N_5016,N_5017,N_5019,N_5021,N_5024,N_5025,N_5026,N_5028,N_5029,N_5031,N_5034,N_5035,N_5037,N_5038,N_5039,N_5041,N_5043,N_5044,N_5046,N_5047,N_5049,N_5050,N_5053,N_5058,N_5060,N_5062,N_5063,N_5064,N_5065,N_5066,N_5068,N_5069,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5086,N_5089,N_5090,N_5093,N_5094,N_5097,N_5099,N_5100,N_5101,N_5102,N_5103,N_5105,N_5106,N_5107,N_5108,N_5109,N_5112,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5126,N_5127,N_5129,N_5132,N_5133,N_5134,N_5136,N_5137,N_5140,N_5141,N_5144,N_5145,N_5148,N_5150,N_5151,N_5152,N_5155,N_5157,N_5158,N_5159,N_5163,N_5164,N_5166,N_5167,N_5169,N_5170,N_5171,N_5172,N_5177,N_5180,N_5185,N_5186,N_5187,N_5188,N_5191,N_5192,N_5193,N_5194,N_5197,N_5198,N_5199,N_5200,N_5202,N_5204,N_5205,N_5206,N_5207,N_5209,N_5210,N_5211,N_5212,N_5215,N_5216,N_5217,N_5218,N_5220,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5231,N_5232,N_5238,N_5239,N_5240,N_5241,N_5242,N_5244,N_5245,N_5247,N_5250,N_5251,N_5252,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5273,N_5274,N_5275,N_5278,N_5279,N_5280,N_5281,N_5282,N_5284,N_5286,N_5287,N_5289,N_5292,N_5294,N_5296,N_5298,N_5302,N_5304,N_5305,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5317,N_5318,N_5319,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5334,N_5335,N_5336,N_5338,N_5340,N_5344,N_5345,N_5348,N_5351,N_5352,N_5354,N_5357,N_5358,N_5359,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5373,N_5374,N_5375,N_5377,N_5381,N_5382,N_5385,N_5387,N_5388,N_5389,N_5390,N_5393,N_5394,N_5397,N_5398,N_5399,N_5400,N_5403,N_5404,N_5405,N_5409,N_5410,N_5412,N_5413,N_5415,N_5416,N_5417,N_5418,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5433,N_5434,N_5436,N_5438,N_5441,N_5442,N_5443,N_5447,N_5448,N_5450,N_5452,N_5453,N_5454,N_5456,N_5457,N_5460,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5474,N_5478,N_5481,N_5483,N_5486,N_5487,N_5488,N_5489,N_5490,N_5492,N_5494,N_5495,N_5496,N_5497,N_5498,N_5501,N_5502,N_5503,N_5504,N_5506,N_5512,N_5513,N_5514,N_5517,N_5518,N_5524,N_5526,N_5527,N_5529,N_5530,N_5535,N_5536,N_5537,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5560,N_5561,N_5562,N_5563,N_5564,N_5566,N_5567,N_5568,N_5570,N_5571,N_5572,N_5574,N_5575,N_5577,N_5578,N_5579,N_5580,N_5581,N_5583,N_5584,N_5585,N_5586,N_5588,N_5590,N_5592,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5607,N_5609,N_5611,N_5612,N_5615,N_5618,N_5619,N_5621,N_5622,N_5625,N_5627,N_5628,N_5631,N_5632,N_5635,N_5636,N_5637,N_5640,N_5644,N_5645,N_5647,N_5648,N_5649,N_5651,N_5654,N_5655,N_5657,N_5659,N_5660,N_5662,N_5663,N_5664,N_5665,N_5666,N_5668,N_5669,N_5670,N_5672,N_5675,N_5677,N_5679,N_5680,N_5681,N_5682,N_5684,N_5685,N_5687,N_5688,N_5689,N_5690,N_5693,N_5697,N_5700,N_5701,N_5702,N_5703,N_5707,N_5708,N_5709,N_5710,N_5711,N_5713,N_5714,N_5715,N_5716,N_5718,N_5719,N_5721,N_5723,N_5725,N_5727,N_5729,N_5730,N_5734,N_5736,N_5737,N_5739,N_5742,N_5743,N_5745,N_5746,N_5747,N_5748,N_5750,N_5753,N_5754,N_5756,N_5758,N_5760,N_5762,N_5763,N_5764,N_5765,N_5766,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5776,N_5780,N_5783,N_5786,N_5788,N_5790,N_5791,N_5792,N_5793,N_5796,N_5797,N_5798,N_5801,N_5802,N_5803,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5820,N_5821,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5834,N_5835,N_5836,N_5841,N_5842,N_5845,N_5846,N_5848,N_5852,N_5854,N_5855,N_5856,N_5858,N_5860,N_5862,N_5863,N_5865,N_5866,N_5869,N_5872,N_5873,N_5874,N_5877,N_5879,N_5880,N_5881,N_5883,N_5884,N_5887,N_5892,N_5893,N_5894,N_5896,N_5897,N_5899,N_5901,N_5902,N_5904,N_5905,N_5906,N_5909,N_5910,N_5913,N_5914,N_5915,N_5917,N_5918,N_5920,N_5923,N_5926,N_5928,N_5929,N_5936,N_5939,N_5940,N_5941,N_5943,N_5945,N_5946,N_5947,N_5948,N_5951,N_5952,N_5953,N_5954,N_5956,N_5958,N_5960,N_5961,N_5963,N_5964,N_5965,N_5967,N_5969,N_5970,N_5972,N_5975,N_5977,N_5978,N_5979,N_5982,N_5983,N_5984,N_5986,N_5987,N_5988,N_5989,N_5990,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6005,N_6006,N_6007,N_6009,N_6010,N_6011,N_6013,N_6014,N_6016,N_6018,N_6020,N_6021,N_6022,N_6023,N_6024,N_6026,N_6027,N_6028,N_6030,N_6032,N_6034,N_6036,N_6037,N_6039,N_6040,N_6041,N_6043,N_6047,N_6049,N_6051,N_6052,N_6054,N_6055,N_6057,N_6058,N_6059,N_6060,N_6062,N_6063,N_6065,N_6066,N_6067,N_6068,N_6070,N_6071,N_6074,N_6076,N_6077,N_6078,N_6081,N_6083,N_6084,N_6085,N_6088,N_6089,N_6090,N_6092,N_6093,N_6096,N_6097,N_6098,N_6100,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6119,N_6122,N_6124,N_6125,N_6126,N_6127,N_6128,N_6131,N_6132,N_6133,N_6134,N_6135,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6147,N_6148,N_6149,N_6154,N_6155,N_6157,N_6160,N_6161,N_6162,N_6164,N_6167,N_6170,N_6171,N_6175,N_6176,N_6177,N_6179,N_6180,N_6181,N_6183,N_6185,N_6186,N_6198,N_6201,N_6203,N_6204,N_6205,N_6208,N_6209,N_6212,N_6213,N_6214,N_6215,N_6216,N_6218,N_6219,N_6223,N_6224,N_6225,N_6226,N_6229,N_6230,N_6231,N_6233,N_6234,N_6236,N_6240,N_6241,N_6243,N_6246,N_6247,N_6248,N_6249,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6261,N_6262,N_6266,N_6267,N_6268,N_6269,N_6271,N_6272,N_6274,N_6276,N_6277,N_6278,N_6279,N_6282,N_6284,N_6285,N_6286,N_6287,N_6291,N_6292,N_6293,N_6297,N_6302,N_6305,N_6306,N_6308,N_6309,N_6310,N_6312,N_6314,N_6317,N_6319,N_6322,N_6323,N_6324,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6335,N_6336,N_6337,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6350,N_6352,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6365,N_6366,N_6367,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6378,N_6382,N_6383,N_6384,N_6388,N_6389,N_6390,N_6392,N_6394,N_6395,N_6396,N_6397,N_6399,N_6400,N_6402,N_6403,N_6407,N_6408,N_6409,N_6412,N_6413,N_6415,N_6416,N_6417,N_6419,N_6420,N_6423,N_6424,N_6425,N_6426,N_6428,N_6429,N_6431,N_6434,N_6435,N_6437,N_6439,N_6440,N_6442,N_6443,N_6445,N_6446,N_6447,N_6448,N_6449,N_6451,N_6452,N_6453,N_6454,N_6455,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6468,N_6469,N_6470,N_6471,N_6474,N_6475,N_6479,N_6480,N_6481,N_6482,N_6486,N_6490,N_6491,N_6492,N_6495,N_6497,N_6498,N_6499,N_6502,N_6503,N_6504,N_6505,N_6506,N_6508,N_6509,N_6510,N_6513,N_6515,N_6518,N_6520,N_6521,N_6524,N_6525,N_6529,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6540,N_6543,N_6544,N_6545,N_6547,N_6549,N_6551,N_6555,N_6556,N_6557,N_6560,N_6561,N_6562,N_6563,N_6565,N_6566,N_6567,N_6569,N_6570,N_6572,N_6574,N_6575,N_6576,N_6577,N_6579,N_6581,N_6582,N_6583,N_6585,N_6586,N_6587,N_6588,N_6591,N_6594,N_6596,N_6600,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6610,N_6612,N_6613,N_6617,N_6619,N_6622,N_6623,N_6624,N_6629,N_6630,N_6631,N_6632,N_6633,N_6635,N_6637,N_6638,N_6642,N_6643,N_6645,N_6649,N_6651,N_6653,N_6658,N_6661,N_6662,N_6664,N_6665,N_6666,N_6667,N_6668,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6681,N_6682,N_6684,N_6685,N_6688,N_6690,N_6692,N_6693,N_6694,N_6695,N_6700,N_6701,N_6702,N_6703,N_6706,N_6709,N_6712,N_6713,N_6714,N_6715,N_6719,N_6720,N_6721,N_6722,N_6723,N_6725,N_6726,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6739,N_6740,N_6741,N_6743,N_6744,N_6745,N_6746,N_6749,N_6750,N_6751,N_6753,N_6754,N_6755,N_6756,N_6757,N_6759,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6781,N_6786,N_6788,N_6792,N_6793,N_6798,N_6803,N_6804,N_6805,N_6806,N_6808,N_6814,N_6815,N_6817,N_6818,N_6819,N_6822,N_6825,N_6827,N_6829,N_6830,N_6833,N_6835,N_6837,N_6838,N_6840,N_6842,N_6843,N_6846,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6855,N_6856,N_6857,N_6858,N_6860,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6869,N_6870,N_6871,N_6873,N_6876,N_6877,N_6878,N_6879,N_6880,N_6883,N_6884,N_6885,N_6886,N_6887,N_6889,N_6890,N_6893,N_6894,N_6895,N_6896,N_6899,N_6900,N_6902,N_6903,N_6905,N_6906,N_6907,N_6909,N_6910,N_6911,N_6914,N_6915,N_6916,N_6917,N_6920,N_6921,N_6922,N_6925,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6938,N_6941,N_6942,N_6943,N_6944,N_6945,N_6950,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6963,N_6967,N_6968,N_6970,N_6971,N_6972,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6981,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_7004,N_7005,N_7006,N_7009,N_7011,N_7013,N_7016,N_7020,N_7021,N_7027,N_7028,N_7037,N_7039,N_7040,N_7042,N_7043,N_7045,N_7048,N_7052,N_7053,N_7057,N_7058,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7073,N_7074,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7092,N_7093,N_7094,N_7095,N_7097,N_7099,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7113,N_7114,N_7116,N_7118,N_7119,N_7120,N_7121,N_7124,N_7126,N_7127,N_7129,N_7131,N_7134,N_7136,N_7137,N_7138,N_7139,N_7142,N_7144,N_7146,N_7147,N_7148,N_7149,N_7151,N_7152,N_7153,N_7155,N_7156,N_7157,N_7158,N_7160,N_7161,N_7164,N_7168,N_7169,N_7170,N_7171,N_7172,N_7176,N_7178,N_7182,N_7183,N_7184,N_7185,N_7187,N_7188,N_7190,N_7191,N_7197,N_7198,N_7200,N_7202,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7222,N_7223,N_7226,N_7227,N_7228,N_7232,N_7233,N_7236,N_7237,N_7238,N_7240,N_7242,N_7243,N_7244,N_7246,N_7247,N_7248,N_7249,N_7253,N_7254,N_7256,N_7257,N_7258,N_7259,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7269,N_7270,N_7271,N_7272,N_7273,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7284,N_7287,N_7291,N_7293,N_7294,N_7295,N_7296,N_7298,N_7300,N_7302,N_7305,N_7306,N_7307,N_7309,N_7310,N_7311,N_7313,N_7314,N_7315,N_7316,N_7317,N_7321,N_7323,N_7324,N_7326,N_7327,N_7330,N_7331,N_7332,N_7335,N_7336,N_7337,N_7338,N_7339,N_7341,N_7342,N_7347,N_7348,N_7350,N_7351,N_7352,N_7353,N_7355,N_7356,N_7358,N_7359,N_7360,N_7362,N_7363,N_7366,N_7373,N_7374,N_7376,N_7377,N_7379,N_7381,N_7382,N_7383,N_7386,N_7387,N_7388,N_7389,N_7391,N_7392,N_7395,N_7397,N_7400,N_7401,N_7405,N_7407,N_7408,N_7409,N_7411,N_7412,N_7413,N_7414,N_7416,N_7417,N_7418,N_7421,N_7422,N_7423,N_7425,N_7427,N_7428,N_7429,N_7431,N_7432,N_7433,N_7434,N_7437,N_7438,N_7439,N_7444,N_7447,N_7448,N_7449,N_7452,N_7456,N_7457,N_7458,N_7459,N_7462,N_7464,N_7466,N_7468,N_7469,N_7472,N_7473,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7492,N_7493,N_7495,N_7496,N_7497,N_7498,N_7499,N_7503,N_7508,N_7509,N_7510,N_7511,N_7512,N_7514,N_7515,N_7516,N_7520,N_7521,N_7522,N_7523,N_7524,N_7526,N_7531,N_7532,N_7533,N_7534,N_7536,N_7538,N_7542,N_7543,N_7544,N_7548,N_7549,N_7550,N_7551,N_7553,N_7554,N_7556,N_7557,N_7560,N_7561,N_7563,N_7567,N_7569,N_7570,N_7571,N_7573,N_7574,N_7577,N_7578,N_7580,N_7581,N_7582,N_7584,N_7585,N_7587,N_7590,N_7592,N_7593,N_7594,N_7598,N_7599,N_7603,N_7604,N_7605,N_7606,N_7607,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7618,N_7620,N_7621,N_7623,N_7625,N_7626,N_7627,N_7629,N_7632,N_7633,N_7635,N_7637,N_7642,N_7645,N_7646,N_7648,N_7649,N_7650,N_7651,N_7656,N_7657,N_7658,N_7662,N_7663,N_7664,N_7666,N_7667,N_7668,N_7669,N_7672,N_7673,N_7674,N_7675,N_7676,N_7678,N_7680,N_7681,N_7682,N_7683,N_7684,N_7687,N_7688,N_7691,N_7694,N_7697,N_7699,N_7700,N_7703,N_7705,N_7706,N_7707,N_7710,N_7711,N_7713,N_7714,N_7715,N_7716,N_7718,N_7720,N_7722,N_7723,N_7724,N_7725,N_7727,N_7728,N_7729,N_7730,N_7731,N_7735,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7744,N_7746,N_7747,N_7748,N_7754,N_7759,N_7760,N_7761,N_7762,N_7764,N_7765,N_7766,N_7769,N_7770,N_7771,N_7774,N_7775,N_7777,N_7779,N_7780,N_7781,N_7784,N_7786,N_7787,N_7788,N_7790,N_7792,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7805,N_7806,N_7809,N_7811,N_7812,N_7814,N_7816,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7830,N_7831,N_7832,N_7833,N_7835,N_7836,N_7838,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7851,N_7852,N_7853,N_7854,N_7858,N_7859,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7870,N_7875,N_7876,N_7877,N_7878,N_7880,N_7882,N_7883,N_7884,N_7886,N_7888,N_7891,N_7892,N_7893,N_7895,N_7898,N_7899,N_7900,N_7901,N_7903,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7919,N_7921,N_7923,N_7925,N_7929,N_7930,N_7932,N_7935,N_7936,N_7939,N_7940,N_7943,N_7945,N_7950,N_7954,N_7956,N_7958,N_7959,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7969,N_7970,N_7971,N_7973,N_7975,N_7979,N_7980,N_7983,N_7984,N_7986,N_7991,N_7994,N_7995,N_7996,N_7998,N_7999,N_8000,N_8001,N_8003,N_8004,N_8008,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8017,N_8018,N_8020,N_8022,N_8025,N_8026,N_8027,N_8028,N_8029,N_8033,N_8034,N_8035,N_8037,N_8039,N_8046,N_8048,N_8050,N_8053,N_8054,N_8055,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8074,N_8075,N_8076,N_8077,N_8078,N_8080,N_8082,N_8083,N_8086,N_8088,N_8089,N_8090,N_8092,N_8093,N_8094,N_8096,N_8099,N_8100,N_8104,N_8106,N_8107,N_8109,N_8110,N_8111,N_8112,N_8116,N_8117,N_8118,N_8120,N_8121,N_8122,N_8124,N_8125,N_8126,N_8128,N_8129,N_8131,N_8132,N_8133,N_8134,N_8136,N_8139,N_8143,N_8144,N_8146,N_8147,N_8148,N_8149,N_8151,N_8152,N_8157,N_8158,N_8160,N_8161,N_8162,N_8164,N_8165,N_8166,N_8167,N_8172,N_8174,N_8175,N_8176,N_8177,N_8179,N_8180,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8190,N_8191,N_8192,N_8193,N_8200,N_8202,N_8203,N_8204,N_8206,N_8207,N_8208,N_8211,N_8214,N_8215,N_8216,N_8218,N_8220,N_8221,N_8224,N_8229,N_8230,N_8232,N_8233,N_8234,N_8235,N_8237,N_8239,N_8240,N_8241,N_8243,N_8244,N_8246,N_8252,N_8253,N_8255,N_8257,N_8258,N_8259,N_8260,N_8261,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8271,N_8273,N_8275,N_8276,N_8277,N_8278,N_8279,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8290,N_8291,N_8292,N_8293,N_8294,N_8297,N_8300,N_8301,N_8302,N_8304,N_8306,N_8307,N_8308,N_8312,N_8313,N_8314,N_8316,N_8317,N_8318,N_8323,N_8325,N_8326,N_8331,N_8332,N_8333,N_8334,N_8336,N_8339,N_8340,N_8344,N_8346,N_8347,N_8349,N_8350,N_8351,N_8355,N_8356,N_8359,N_8360,N_8364,N_8368,N_8369,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8380,N_8381,N_8382,N_8383,N_8385,N_8386,N_8389,N_8390,N_8393,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8405,N_8406,N_8407,N_8408,N_8413,N_8415,N_8417,N_8420,N_8421,N_8425,N_8426,N_8429,N_8430,N_8431,N_8438,N_8439,N_8440,N_8441,N_8443,N_8444,N_8445,N_8448,N_8449,N_8450,N_8452,N_8453,N_8454,N_8456,N_8457,N_8460,N_8464,N_8468,N_8471,N_8473,N_8474,N_8475,N_8476,N_8479,N_8481,N_8482,N_8483,N_8486,N_8488,N_8491,N_8493,N_8494,N_8496,N_8499,N_8501,N_8502,N_8503,N_8508,N_8509,N_8510,N_8511,N_8512,N_8516,N_8519,N_8523,N_8528,N_8529,N_8532,N_8533,N_8536,N_8537,N_8538,N_8540,N_8543,N_8545,N_8547,N_8549,N_8551,N_8552,N_8554,N_8555,N_8556,N_8558,N_8559,N_8560,N_8561,N_8565,N_8568,N_8569,N_8572,N_8573,N_8575,N_8578,N_8579,N_8581,N_8582,N_8583,N_8586,N_8587,N_8588,N_8590,N_8591,N_8594,N_8597,N_8599,N_8600,N_8605,N_8607,N_8608,N_8611,N_8615,N_8617,N_8618,N_8620,N_8623,N_8626,N_8627,N_8631,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8643,N_8644,N_8646,N_8648,N_8650,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8660,N_8661,N_8662,N_8663,N_8664,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8675,N_8676,N_8678,N_8679,N_8682,N_8683,N_8684,N_8686,N_8687,N_8688,N_8689,N_8690,N_8696,N_8699,N_8700,N_8701,N_8702,N_8703,N_8705,N_8707,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8716,N_8717,N_8719,N_8721,N_8725,N_8726,N_8727,N_8729,N_8732,N_8733,N_8734,N_8736,N_8739,N_8740,N_8742,N_8743,N_8744,N_8745,N_8748,N_8749,N_8750,N_8751,N_8753,N_8756,N_8758,N_8762,N_8764,N_8766,N_8767,N_8768,N_8769,N_8772,N_8777,N_8780,N_8782,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8794,N_8795,N_8799,N_8800,N_8801,N_8802,N_8803,N_8806,N_8808,N_8809,N_8810,N_8811,N_8817,N_8818,N_8819,N_8820,N_8821,N_8823,N_8824,N_8826,N_8827,N_8828,N_8829,N_8831,N_8834,N_8836,N_8837,N_8838,N_8839,N_8840,N_8844,N_8846,N_8847,N_8849,N_8852,N_8853,N_8855,N_8857,N_8858,N_8859,N_8865,N_8866,N_8867,N_8868,N_8869,N_8871,N_8872,N_8873,N_8874,N_8876,N_8879,N_8880,N_8881,N_8883,N_8886,N_8889,N_8890,N_8892,N_8893,N_8895,N_8896,N_8897,N_8900,N_8901,N_8902,N_8904,N_8905,N_8910,N_8911,N_8913,N_8914,N_8916,N_8917,N_8920,N_8921,N_8922,N_8929,N_8931,N_8933,N_8934,N_8935,N_8936,N_8939,N_8941,N_8942,N_8944,N_8945,N_8947,N_8948,N_8949,N_8950,N_8952,N_8953,N_8955,N_8957,N_8959,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8972,N_8973,N_8975,N_8977,N_8978,N_8979,N_8980,N_8982,N_8983,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8994,N_8996,N_8998,N_9000,N_9001,N_9002,N_9003,N_9005,N_9006,N_9008,N_9010,N_9011,N_9012,N_9014,N_9016,N_9017,N_9018,N_9019,N_9022,N_9023,N_9024,N_9028,N_9031,N_9033,N_9034,N_9036,N_9037,N_9038,N_9039,N_9042,N_9044,N_9046,N_9047,N_9049,N_9051,N_9052,N_9053,N_9055,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9065,N_9066,N_9067,N_9070,N_9072,N_9075,N_9076,N_9077,N_9078,N_9082,N_9084,N_9087,N_9088,N_9089,N_9090,N_9093,N_9096,N_9098,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9114,N_9115,N_9117,N_9118,N_9120,N_9121,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9135,N_9136,N_9138,N_9140,N_9141,N_9142,N_9144,N_9145,N_9148,N_9150,N_9151,N_9153,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9162,N_9163,N_9164,N_9165,N_9166,N_9169,N_9170,N_9171,N_9174,N_9175,N_9179,N_9180,N_9183,N_9186,N_9187,N_9188,N_9189,N_9191,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9206,N_9208,N_9209,N_9211,N_9213,N_9214,N_9215,N_9217,N_9218,N_9220,N_9222,N_9224,N_9229,N_9230,N_9231,N_9233,N_9236,N_9237,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9248,N_9249,N_9250,N_9252,N_9256,N_9257,N_9258,N_9259,N_9261,N_9262,N_9265,N_9267,N_9269,N_9271,N_9272,N_9274,N_9278,N_9281,N_9283,N_9284,N_9286,N_9287,N_9288,N_9290,N_9293,N_9295,N_9296,N_9297,N_9299,N_9301,N_9302,N_9304,N_9306,N_9307,N_9309,N_9311,N_9312,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9323,N_9325,N_9326,N_9327,N_9328,N_9331,N_9332,N_9334,N_9335,N_9338,N_9339,N_9343,N_9345,N_9347,N_9348,N_9352,N_9353,N_9355,N_9356,N_9357,N_9359,N_9360,N_9361,N_9364,N_9365,N_9366,N_9367,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9378,N_9379,N_9381,N_9382,N_9383,N_9385,N_9386,N_9387,N_9389,N_9390,N_9391,N_9392,N_9394,N_9396,N_9397,N_9401,N_9402,N_9403,N_9405,N_9406,N_9407,N_9409,N_9410,N_9411,N_9415,N_9416,N_9419,N_9428,N_9429,N_9432,N_9433,N_9434,N_9435,N_9438,N_9439,N_9441,N_9442,N_9444,N_9447,N_9449,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9459,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9473,N_9474,N_9477,N_9479,N_9480,N_9481,N_9482,N_9483,N_9485,N_9486,N_9488,N_9490,N_9493,N_9495,N_9497,N_9498,N_9501,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9511,N_9512,N_9513,N_9514,N_9516,N_9517,N_9525,N_9527,N_9528,N_9529,N_9530,N_9532,N_9537,N_9538,N_9540,N_9541,N_9545,N_9546,N_9547,N_9550,N_9554,N_9555,N_9556,N_9558,N_9559,N_9560,N_9564,N_9565,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9575,N_9576,N_9577,N_9578,N_9579,N_9583,N_9584,N_9585,N_9586,N_9589,N_9590,N_9591,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9610,N_9612,N_9616,N_9620,N_9622,N_9623,N_9626,N_9627,N_9628,N_9629,N_9632,N_9633,N_9636,N_9637,N_9640,N_9642,N_9643,N_9645,N_9649,N_9652,N_9654,N_9655,N_9657,N_9659,N_9660,N_9661,N_9665,N_9668,N_9669,N_9672,N_9673,N_9676,N_9677,N_9679,N_9680,N_9681,N_9682,N_9684,N_9686,N_9687,N_9688,N_9689,N_9691,N_9692,N_9696,N_9698,N_9700,N_9702,N_9703,N_9704,N_9705,N_9707,N_9708,N_9709,N_9712,N_9713,N_9714,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9729,N_9732,N_9734,N_9735,N_9736,N_9738,N_9740,N_9742,N_9744,N_9745,N_9747,N_9748,N_9750,N_9753,N_9754,N_9755,N_9756,N_9760,N_9761,N_9762,N_9764,N_9765,N_9766,N_9767,N_9774,N_9775,N_9776,N_9777,N_9779,N_9784,N_9785,N_9787,N_9788,N_9790,N_9791,N_9792,N_9793,N_9799,N_9800,N_9802,N_9803,N_9804,N_9805,N_9807,N_9808,N_9809,N_9811,N_9812,N_9813,N_9814,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9825,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9837,N_9838,N_9839,N_9840,N_9843,N_9844,N_9845,N_9846,N_9848,N_9849,N_9850,N_9852,N_9856,N_9857,N_9858,N_9859,N_9861,N_9863,N_9864,N_9865,N_9867,N_9868,N_9869,N_9870,N_9873,N_9874,N_9875,N_9877,N_9878,N_9879,N_9880,N_9882,N_9883,N_9884,N_9885,N_9886,N_9888,N_9889,N_9890,N_9892,N_9893,N_9896,N_9897,N_9899,N_9904,N_9905,N_9908,N_9909,N_9910,N_9911,N_9912,N_9914,N_9916,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9925,N_9926,N_9927,N_9928,N_9929,N_9931,N_9932,N_9933,N_9935,N_9937,N_9939,N_9942,N_9946,N_9948,N_9949,N_9950,N_9954,N_9958,N_9959,N_9962,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9971,N_9973,N_9974,N_9975,N_9976,N_9977,N_9979,N_9980,N_9983,N_9985,N_9986,N_9989,N_9990,N_9993,N_9994,N_9995,N_9996,N_9997,N_9999;
and U0 (N_0,In_945,In_609);
nor U1 (N_1,In_25,In_370);
and U2 (N_2,In_283,In_716);
or U3 (N_3,In_274,In_151);
and U4 (N_4,In_602,In_873);
nand U5 (N_5,In_207,In_613);
or U6 (N_6,In_11,In_931);
and U7 (N_7,In_148,In_682);
and U8 (N_8,In_233,In_941);
and U9 (N_9,In_639,In_728);
and U10 (N_10,In_28,In_14);
nor U11 (N_11,In_778,In_54);
or U12 (N_12,In_40,In_831);
nor U13 (N_13,In_813,In_449);
or U14 (N_14,In_900,In_278);
nor U15 (N_15,In_184,In_896);
nand U16 (N_16,In_255,In_275);
nor U17 (N_17,In_629,In_976);
or U18 (N_18,In_38,In_348);
nor U19 (N_19,In_9,In_322);
or U20 (N_20,In_339,In_628);
nand U21 (N_21,In_756,In_371);
nor U22 (N_22,In_467,In_817);
nand U23 (N_23,In_897,In_500);
nor U24 (N_24,In_169,In_520);
and U25 (N_25,In_21,In_460);
or U26 (N_26,In_83,In_804);
or U27 (N_27,In_487,In_236);
or U28 (N_28,In_329,In_267);
or U29 (N_29,In_443,In_819);
nand U30 (N_30,In_225,In_424);
or U31 (N_31,In_928,In_195);
and U32 (N_32,In_97,In_916);
or U33 (N_33,In_358,In_893);
nor U34 (N_34,In_361,In_212);
or U35 (N_35,In_310,In_986);
nand U36 (N_36,In_781,In_395);
or U37 (N_37,In_431,In_191);
and U38 (N_38,In_159,In_874);
nand U39 (N_39,In_718,In_49);
nand U40 (N_40,In_4,In_347);
or U41 (N_41,In_806,In_394);
or U42 (N_42,In_122,In_930);
or U43 (N_43,In_492,In_3);
nand U44 (N_44,In_702,In_232);
nor U45 (N_45,In_209,In_989);
or U46 (N_46,In_344,In_37);
and U47 (N_47,In_827,In_437);
or U48 (N_48,In_170,In_414);
or U49 (N_49,In_853,In_301);
nor U50 (N_50,In_39,In_509);
nand U51 (N_51,In_338,In_112);
and U52 (N_52,In_803,In_118);
and U53 (N_53,In_636,In_528);
nor U54 (N_54,In_109,In_997);
nand U55 (N_55,In_953,In_904);
or U56 (N_56,In_811,In_768);
nor U57 (N_57,In_889,In_459);
or U58 (N_58,In_511,In_651);
and U59 (N_59,In_674,In_747);
nor U60 (N_60,In_452,In_470);
nand U61 (N_61,In_421,In_825);
and U62 (N_62,In_497,In_248);
or U63 (N_63,In_375,In_563);
or U64 (N_64,In_712,In_480);
nand U65 (N_65,In_489,In_918);
nand U66 (N_66,In_942,In_643);
nor U67 (N_67,In_15,In_554);
and U68 (N_68,In_741,In_998);
nand U69 (N_69,In_504,In_534);
and U70 (N_70,In_955,In_136);
and U71 (N_71,In_245,In_271);
nor U72 (N_72,In_693,In_525);
or U73 (N_73,In_672,In_564);
and U74 (N_74,In_357,In_679);
or U75 (N_75,In_968,In_915);
nand U76 (N_76,In_911,In_273);
nor U77 (N_77,In_216,In_321);
and U78 (N_78,In_192,In_517);
nor U79 (N_79,In_752,In_346);
nor U80 (N_80,In_802,In_201);
or U81 (N_81,In_886,In_164);
nor U82 (N_82,In_972,In_48);
nor U83 (N_83,In_105,In_836);
nand U84 (N_84,In_971,In_320);
or U85 (N_85,In_566,In_24);
and U86 (N_86,In_570,In_65);
xnor U87 (N_87,In_128,In_155);
nand U88 (N_88,In_656,In_202);
and U89 (N_89,In_632,In_457);
nor U90 (N_90,In_389,In_582);
nor U91 (N_91,In_603,In_352);
or U92 (N_92,In_568,In_75);
nand U93 (N_93,In_678,In_964);
nor U94 (N_94,In_765,In_743);
and U95 (N_95,In_469,In_579);
nand U96 (N_96,In_797,In_518);
xnor U97 (N_97,In_992,In_120);
xnor U98 (N_98,In_295,In_466);
or U99 (N_99,In_77,In_982);
nand U100 (N_100,In_513,In_556);
nor U101 (N_101,In_531,In_58);
nand U102 (N_102,In_872,In_841);
or U103 (N_103,In_816,In_277);
nor U104 (N_104,In_445,In_724);
or U105 (N_105,In_117,In_411);
nand U106 (N_106,In_464,In_826);
or U107 (N_107,In_405,In_547);
or U108 (N_108,In_345,In_887);
and U109 (N_109,In_709,In_296);
nor U110 (N_110,In_219,In_843);
and U111 (N_111,In_516,In_689);
nor U112 (N_112,In_397,In_313);
nand U113 (N_113,In_221,In_150);
nor U114 (N_114,In_910,In_95);
or U115 (N_115,In_635,In_734);
and U116 (N_116,In_199,In_454);
nand U117 (N_117,In_108,In_10);
nand U118 (N_118,In_922,In_455);
and U119 (N_119,In_61,In_850);
and U120 (N_120,In_879,In_481);
or U121 (N_121,In_828,In_549);
nor U122 (N_122,In_933,In_145);
and U123 (N_123,In_875,In_400);
nand U124 (N_124,In_533,In_490);
or U125 (N_125,In_735,In_623);
and U126 (N_126,In_576,In_994);
or U127 (N_127,In_965,In_494);
or U128 (N_128,In_434,In_641);
nor U129 (N_129,In_798,In_81);
and U130 (N_130,In_606,In_809);
nand U131 (N_131,In_152,In_305);
nor U132 (N_132,In_263,In_823);
or U133 (N_133,In_272,In_697);
nand U134 (N_134,In_433,In_572);
nand U135 (N_135,In_608,In_349);
nor U136 (N_136,In_589,In_407);
nor U137 (N_137,In_762,In_393);
or U138 (N_138,In_304,In_43);
or U139 (N_139,In_12,In_343);
and U140 (N_140,In_858,In_746);
nor U141 (N_141,In_103,In_124);
nor U142 (N_142,In_574,In_367);
nor U143 (N_143,In_440,In_234);
nand U144 (N_144,In_413,In_404);
or U145 (N_145,In_388,In_140);
nand U146 (N_146,In_591,In_260);
nor U147 (N_147,In_607,In_56);
xnor U148 (N_148,In_204,In_426);
and U149 (N_149,In_259,In_732);
and U150 (N_150,In_753,In_156);
nor U151 (N_151,In_585,In_261);
nand U152 (N_152,In_439,In_314);
or U153 (N_153,In_90,In_829);
nor U154 (N_154,In_451,In_241);
or U155 (N_155,In_175,In_557);
nor U156 (N_156,In_91,In_22);
or U157 (N_157,In_427,In_666);
and U158 (N_158,In_485,In_146);
or U159 (N_159,In_415,In_761);
nand U160 (N_160,In_665,In_754);
xor U161 (N_161,In_316,In_921);
nand U162 (N_162,In_412,In_383);
nand U163 (N_163,In_331,In_929);
nor U164 (N_164,In_93,In_795);
nand U165 (N_165,In_799,In_227);
nand U166 (N_166,In_782,In_26);
or U167 (N_167,In_611,In_392);
or U168 (N_168,In_281,In_612);
nor U169 (N_169,In_884,In_174);
and U170 (N_170,In_950,In_704);
nand U171 (N_171,In_715,In_744);
xnor U172 (N_172,In_581,In_162);
nand U173 (N_173,In_94,In_948);
nand U174 (N_174,In_726,In_142);
and U175 (N_175,In_340,In_23);
nor U176 (N_176,In_569,In_293);
nand U177 (N_177,In_44,In_845);
or U178 (N_178,In_129,In_740);
or U179 (N_179,In_699,In_189);
and U180 (N_180,In_420,In_544);
nand U181 (N_181,In_777,In_963);
nor U182 (N_182,In_220,In_441);
nand U183 (N_183,In_327,In_330);
nand U184 (N_184,In_805,In_332);
or U185 (N_185,In_398,In_88);
or U186 (N_186,In_378,In_890);
and U187 (N_187,In_498,In_961);
nand U188 (N_188,In_840,In_106);
and U189 (N_189,In_832,In_640);
nand U190 (N_190,In_542,In_101);
or U191 (N_191,In_610,In_700);
and U192 (N_192,In_537,In_707);
nor U193 (N_193,In_815,In_903);
or U194 (N_194,In_710,In_962);
or U195 (N_195,In_409,In_917);
nor U196 (N_196,In_265,In_226);
or U197 (N_197,In_33,In_229);
and U198 (N_198,In_299,In_157);
nor U199 (N_199,In_791,In_512);
or U200 (N_200,In_16,In_92);
and U201 (N_201,In_645,In_599);
nand U202 (N_202,In_792,In_503);
and U203 (N_203,In_317,In_954);
nand U204 (N_204,In_901,In_76);
and U205 (N_205,In_308,In_67);
or U206 (N_206,In_359,In_658);
or U207 (N_207,In_369,In_578);
nor U208 (N_208,In_333,In_760);
or U209 (N_209,In_486,In_914);
nand U210 (N_210,In_973,In_7);
xor U211 (N_211,In_84,In_461);
nand U212 (N_212,In_324,In_661);
nand U213 (N_213,In_771,In_113);
or U214 (N_214,In_794,In_130);
or U215 (N_215,In_864,In_834);
nand U216 (N_216,In_690,In_172);
nor U217 (N_217,In_720,In_228);
nor U218 (N_218,In_264,In_750);
and U219 (N_219,In_714,In_319);
nor U220 (N_220,In_692,In_402);
nand U221 (N_221,In_42,In_733);
and U222 (N_222,In_685,In_684);
nand U223 (N_223,In_247,In_515);
and U224 (N_224,In_708,In_934);
nor U225 (N_225,In_68,In_844);
nor U226 (N_226,In_725,In_208);
or U227 (N_227,In_631,In_307);
nor U228 (N_228,In_379,In_671);
nor U229 (N_229,In_507,In_558);
or U230 (N_230,In_303,In_981);
nor U231 (N_231,In_738,In_550);
nor U232 (N_232,In_165,In_362);
xor U233 (N_233,In_462,In_252);
and U234 (N_234,In_865,In_104);
nand U235 (N_235,In_430,In_979);
nor U236 (N_236,In_772,In_885);
nor U237 (N_237,In_892,In_824);
nor U238 (N_238,In_337,In_996);
or U239 (N_239,In_620,In_438);
or U240 (N_240,In_687,In_924);
nor U241 (N_241,In_217,In_131);
nor U242 (N_242,In_800,In_302);
nor U243 (N_243,In_648,In_616);
or U244 (N_244,In_126,In_253);
nor U245 (N_245,In_959,In_851);
or U246 (N_246,In_597,In_2);
and U247 (N_247,In_250,In_479);
xnor U248 (N_248,In_240,In_354);
nor U249 (N_249,In_860,In_980);
and U250 (N_250,In_244,In_399);
nor U251 (N_251,In_650,In_677);
nor U252 (N_252,In_653,In_417);
and U253 (N_253,In_571,In_475);
or U254 (N_254,In_553,In_315);
nand U255 (N_255,In_759,In_231);
nor U256 (N_256,In_6,In_154);
and U257 (N_257,In_766,In_284);
and U258 (N_258,In_842,In_652);
or U259 (N_259,In_213,In_71);
nor U260 (N_260,In_510,In_453);
nand U261 (N_261,In_654,In_655);
xnor U262 (N_262,In_495,In_618);
and U263 (N_263,In_861,In_180);
and U264 (N_264,In_990,In_123);
nand U265 (N_265,In_133,In_871);
nand U266 (N_266,In_908,In_902);
nor U267 (N_267,In_270,In_664);
or U268 (N_268,In_465,In_203);
nor U269 (N_269,In_755,In_416);
and U270 (N_270,In_300,In_138);
nand U271 (N_271,In_541,In_215);
and U272 (N_272,In_211,In_880);
or U273 (N_273,In_560,In_214);
and U274 (N_274,In_974,In_89);
xnor U275 (N_275,In_717,In_907);
or U276 (N_276,In_855,In_977);
nand U277 (N_277,In_121,In_206);
nor U278 (N_278,In_696,In_539);
nand U279 (N_279,In_291,In_775);
and U280 (N_280,In_403,In_983);
nand U281 (N_281,In_630,In_730);
and U282 (N_282,In_626,In_17);
or U283 (N_283,In_246,In_944);
nand U284 (N_284,In_312,In_999);
or U285 (N_285,In_551,In_913);
nand U286 (N_286,In_237,In_188);
nor U287 (N_287,In_482,In_595);
or U288 (N_288,In_177,In_670);
nand U289 (N_289,In_20,In_477);
or U290 (N_290,In_456,In_521);
nand U291 (N_291,In_776,In_736);
nand U292 (N_292,In_698,In_705);
and U293 (N_293,In_135,In_625);
and U294 (N_294,In_269,In_519);
nor U295 (N_295,In_298,In_739);
or U296 (N_296,In_662,In_642);
nand U297 (N_297,In_31,In_287);
nand U298 (N_298,In_562,In_341);
or U299 (N_299,In_601,In_18);
nor U300 (N_300,In_70,In_428);
nand U301 (N_301,In_868,In_767);
nand U302 (N_302,In_205,In_268);
or U303 (N_303,In_182,In_168);
and U304 (N_304,In_238,In_149);
and U305 (N_305,In_178,In_691);
nor U306 (N_306,In_731,In_659);
nor U307 (N_307,In_906,In_545);
nor U308 (N_308,In_53,In_555);
nand U309 (N_309,In_527,In_854);
or U310 (N_310,In_139,In_952);
nor U311 (N_311,In_644,In_115);
or U312 (N_312,In_649,In_970);
xor U313 (N_313,In_450,In_158);
or U314 (N_314,In_160,In_141);
and U315 (N_315,In_143,In_780);
nor U316 (N_316,In_198,In_583);
or U317 (N_317,In_529,In_926);
nand U318 (N_318,In_364,In_619);
or U319 (N_319,In_988,In_96);
nor U320 (N_320,In_496,In_669);
or U321 (N_321,In_505,In_748);
nor U322 (N_322,In_111,In_502);
nand U323 (N_323,In_432,In_51);
nand U324 (N_324,In_862,In_366);
and U325 (N_325,In_723,In_350);
or U326 (N_326,In_969,In_787);
nand U327 (N_327,In_458,In_64);
nor U328 (N_328,In_943,In_688);
and U329 (N_329,In_290,In_763);
or U330 (N_330,In_491,In_668);
nor U331 (N_331,In_373,In_72);
or U332 (N_332,In_894,In_377);
nand U333 (N_333,In_737,In_592);
nand U334 (N_334,In_183,In_186);
or U335 (N_335,In_222,In_757);
nor U336 (N_336,In_835,In_663);
and U337 (N_337,In_821,In_565);
nor U338 (N_338,In_615,In_385);
nand U339 (N_339,In_622,In_919);
or U340 (N_340,In_978,In_559);
and U341 (N_341,In_586,In_99);
or U342 (N_342,In_288,In_790);
or U343 (N_343,In_985,In_584);
nor U344 (N_344,In_325,In_27);
or U345 (N_345,In_881,In_524);
and U346 (N_346,In_634,In_975);
or U347 (N_347,In_171,In_624);
and U348 (N_348,In_719,In_167);
and U349 (N_349,In_444,In_788);
nor U350 (N_350,In_258,In_50);
nand U351 (N_351,In_764,In_257);
and U352 (N_352,In_243,In_137);
nand U353 (N_353,In_870,In_423);
nor U354 (N_354,In_535,In_769);
nor U355 (N_355,In_605,In_617);
or U356 (N_356,In_355,In_386);
nor U357 (N_357,In_883,In_633);
and U358 (N_358,In_848,In_401);
nand U359 (N_359,In_722,In_749);
nand U360 (N_360,In_727,In_957);
nand U361 (N_361,In_446,In_476);
nor U362 (N_362,In_960,In_538);
or U363 (N_363,In_74,In_144);
nand U364 (N_364,In_758,In_822);
nor U365 (N_365,In_254,In_604);
nor U366 (N_366,In_577,In_856);
or U367 (N_367,In_311,In_82);
nand U368 (N_368,In_888,In_849);
and U369 (N_369,In_695,In_334);
and U370 (N_370,In_193,In_590);
or U371 (N_371,In_5,In_125);
and U372 (N_372,In_472,In_703);
nor U373 (N_373,In_543,In_947);
nor U374 (N_374,In_36,In_132);
or U375 (N_375,In_380,In_60);
or U376 (N_376,In_587,In_627);
nor U377 (N_377,In_673,In_242);
or U378 (N_378,In_593,In_368);
nand U379 (N_379,In_161,In_408);
xor U380 (N_380,In_523,In_891);
or U381 (N_381,In_289,In_374);
or U382 (N_382,In_938,In_173);
nand U383 (N_383,In_79,In_418);
nand U384 (N_384,In_176,In_867);
or U385 (N_385,In_41,In_29);
and U386 (N_386,In_898,In_223);
or U387 (N_387,In_116,In_384);
nand U388 (N_388,In_830,In_683);
nor U389 (N_389,In_483,In_779);
nand U390 (N_390,In_478,In_471);
and U391 (N_391,In_909,In_647);
and U392 (N_392,In_69,In_442);
nor U393 (N_393,In_210,In_711);
or U394 (N_394,In_360,In_114);
or U395 (N_395,In_540,In_306);
or U396 (N_396,In_573,In_882);
nor U397 (N_397,In_966,In_701);
nand U398 (N_398,In_808,In_35);
xnor U399 (N_399,In_530,In_80);
and U400 (N_400,In_935,In_770);
or U401 (N_401,In_163,In_958);
nand U402 (N_402,In_102,In_838);
nand U403 (N_403,In_179,In_87);
nor U404 (N_404,In_895,In_190);
nor U405 (N_405,In_680,In_396);
or U406 (N_406,In_694,In_425);
nor U407 (N_407,In_837,In_796);
nand U408 (N_408,In_110,In_575);
nand U409 (N_409,In_66,In_372);
or U410 (N_410,In_390,In_419);
nand U411 (N_411,In_532,In_448);
nand U412 (N_412,In_774,In_925);
and U413 (N_413,In_660,In_127);
nand U414 (N_414,In_46,In_376);
and U415 (N_415,In_807,In_493);
or U416 (N_416,In_993,In_561);
and U417 (N_417,In_499,In_936);
nand U418 (N_418,In_614,In_85);
xnor U419 (N_419,In_422,In_920);
nor U420 (N_420,In_351,In_59);
nor U421 (N_421,In_73,In_596);
nand U422 (N_422,In_967,In_580);
and U423 (N_423,In_107,In_335);
nor U424 (N_424,In_818,In_282);
nand U425 (N_425,In_536,In_847);
nand U426 (N_426,In_857,In_19);
nand U427 (N_427,In_342,In_429);
xnor U428 (N_428,In_62,In_742);
nand U429 (N_429,In_353,In_745);
nor U430 (N_430,In_100,In_729);
or U431 (N_431,In_436,In_323);
nor U432 (N_432,In_1,In_147);
or U433 (N_433,In_899,In_789);
or U434 (N_434,In_912,In_773);
and U435 (N_435,In_514,In_667);
nor U436 (N_436,In_356,In_256);
nor U437 (N_437,In_235,In_166);
or U438 (N_438,In_949,In_546);
and U439 (N_439,In_52,In_279);
or U440 (N_440,In_297,In_859);
or U441 (N_441,In_506,In_318);
or U442 (N_442,In_713,In_638);
and U443 (N_443,In_751,In_34);
and U444 (N_444,In_435,In_363);
nor U445 (N_445,In_280,In_951);
nor U446 (N_446,In_181,In_224);
and U447 (N_447,In_946,In_63);
nand U448 (N_448,In_852,In_447);
or U449 (N_449,In_187,In_681);
nand U450 (N_450,In_686,In_995);
nand U451 (N_451,In_783,In_328);
or U452 (N_452,In_508,In_251);
nor U453 (N_453,In_230,In_839);
or U454 (N_454,In_676,In_32);
nor U455 (N_455,In_47,In_387);
and U456 (N_456,In_294,In_13);
and U457 (N_457,In_78,In_292);
nand U458 (N_458,In_869,In_937);
nand U459 (N_459,In_637,In_336);
and U460 (N_460,In_923,In_391);
and U461 (N_461,In_526,In_382);
and U462 (N_462,In_286,In_468);
nand U463 (N_463,In_249,In_984);
nor U464 (N_464,In_8,In_927);
or U465 (N_465,In_474,In_185);
nand U466 (N_466,In_820,In_785);
and U467 (N_467,In_876,In_721);
or U468 (N_468,In_134,In_197);
and U469 (N_469,In_45,In_877);
nand U470 (N_470,In_98,In_365);
or U471 (N_471,In_932,In_55);
nand U472 (N_472,In_940,In_552);
nor U473 (N_473,In_600,In_987);
nand U474 (N_474,In_0,In_706);
or U475 (N_475,In_309,In_86);
and U476 (N_476,In_956,In_239);
nor U477 (N_477,In_621,In_218);
nor U478 (N_478,In_588,In_793);
nor U479 (N_479,In_866,In_410);
or U480 (N_480,In_833,In_194);
or U481 (N_481,In_810,In_657);
or U482 (N_482,In_488,In_262);
nor U483 (N_483,In_786,In_646);
and U484 (N_484,In_266,In_285);
or U485 (N_485,In_801,In_30);
or U486 (N_486,In_598,In_814);
nor U487 (N_487,In_675,In_119);
nor U488 (N_488,In_276,In_326);
and U489 (N_489,In_548,In_473);
nand U490 (N_490,In_484,In_878);
or U491 (N_491,In_863,In_784);
nor U492 (N_492,In_196,In_991);
and U493 (N_493,In_905,In_463);
xnor U494 (N_494,In_594,In_812);
nand U495 (N_495,In_567,In_501);
or U496 (N_496,In_522,In_381);
or U497 (N_497,In_406,In_200);
and U498 (N_498,In_153,In_846);
nor U499 (N_499,In_939,In_57);
or U500 (N_500,In_834,In_957);
nand U501 (N_501,In_753,In_614);
or U502 (N_502,In_367,In_161);
or U503 (N_503,In_513,In_923);
nor U504 (N_504,In_142,In_470);
nor U505 (N_505,In_824,In_959);
nor U506 (N_506,In_327,In_58);
and U507 (N_507,In_3,In_246);
and U508 (N_508,In_590,In_615);
nand U509 (N_509,In_182,In_156);
and U510 (N_510,In_632,In_44);
and U511 (N_511,In_365,In_766);
and U512 (N_512,In_993,In_797);
or U513 (N_513,In_451,In_911);
nand U514 (N_514,In_951,In_526);
or U515 (N_515,In_791,In_110);
and U516 (N_516,In_688,In_435);
and U517 (N_517,In_921,In_293);
nand U518 (N_518,In_864,In_494);
nand U519 (N_519,In_230,In_748);
and U520 (N_520,In_132,In_969);
nor U521 (N_521,In_824,In_571);
nor U522 (N_522,In_525,In_56);
or U523 (N_523,In_105,In_893);
nor U524 (N_524,In_474,In_193);
and U525 (N_525,In_816,In_794);
nor U526 (N_526,In_253,In_738);
and U527 (N_527,In_226,In_768);
nand U528 (N_528,In_195,In_877);
and U529 (N_529,In_979,In_439);
nand U530 (N_530,In_291,In_527);
nor U531 (N_531,In_135,In_917);
nor U532 (N_532,In_77,In_382);
and U533 (N_533,In_473,In_592);
nand U534 (N_534,In_879,In_964);
nor U535 (N_535,In_496,In_280);
or U536 (N_536,In_169,In_753);
nand U537 (N_537,In_974,In_796);
or U538 (N_538,In_824,In_936);
or U539 (N_539,In_863,In_156);
and U540 (N_540,In_480,In_680);
and U541 (N_541,In_327,In_902);
nor U542 (N_542,In_665,In_410);
nor U543 (N_543,In_155,In_630);
nor U544 (N_544,In_171,In_1);
nor U545 (N_545,In_257,In_136);
nand U546 (N_546,In_578,In_288);
and U547 (N_547,In_253,In_214);
or U548 (N_548,In_734,In_441);
or U549 (N_549,In_363,In_634);
nand U550 (N_550,In_244,In_948);
nor U551 (N_551,In_993,In_386);
or U552 (N_552,In_244,In_766);
nand U553 (N_553,In_543,In_282);
nor U554 (N_554,In_486,In_653);
or U555 (N_555,In_952,In_622);
and U556 (N_556,In_664,In_857);
or U557 (N_557,In_471,In_522);
xor U558 (N_558,In_921,In_808);
and U559 (N_559,In_16,In_846);
and U560 (N_560,In_987,In_806);
or U561 (N_561,In_267,In_558);
and U562 (N_562,In_124,In_826);
nor U563 (N_563,In_336,In_386);
or U564 (N_564,In_276,In_676);
and U565 (N_565,In_553,In_366);
and U566 (N_566,In_611,In_361);
and U567 (N_567,In_341,In_798);
nand U568 (N_568,In_222,In_808);
or U569 (N_569,In_340,In_254);
or U570 (N_570,In_987,In_678);
nand U571 (N_571,In_424,In_927);
nor U572 (N_572,In_119,In_906);
or U573 (N_573,In_967,In_100);
and U574 (N_574,In_692,In_467);
or U575 (N_575,In_620,In_567);
nor U576 (N_576,In_540,In_613);
and U577 (N_577,In_18,In_0);
xnor U578 (N_578,In_257,In_457);
nor U579 (N_579,In_467,In_114);
nand U580 (N_580,In_762,In_553);
nand U581 (N_581,In_135,In_945);
and U582 (N_582,In_41,In_446);
and U583 (N_583,In_246,In_60);
nor U584 (N_584,In_829,In_841);
nor U585 (N_585,In_830,In_317);
or U586 (N_586,In_134,In_584);
nor U587 (N_587,In_38,In_666);
nor U588 (N_588,In_847,In_709);
xnor U589 (N_589,In_923,In_920);
or U590 (N_590,In_166,In_120);
nor U591 (N_591,In_503,In_610);
and U592 (N_592,In_253,In_580);
or U593 (N_593,In_500,In_806);
or U594 (N_594,In_731,In_473);
and U595 (N_595,In_645,In_887);
nand U596 (N_596,In_403,In_735);
or U597 (N_597,In_14,In_319);
nand U598 (N_598,In_465,In_834);
and U599 (N_599,In_831,In_866);
nor U600 (N_600,In_328,In_305);
nand U601 (N_601,In_645,In_719);
nand U602 (N_602,In_879,In_444);
and U603 (N_603,In_908,In_85);
or U604 (N_604,In_407,In_623);
and U605 (N_605,In_837,In_563);
or U606 (N_606,In_113,In_676);
and U607 (N_607,In_558,In_956);
nand U608 (N_608,In_334,In_885);
and U609 (N_609,In_822,In_675);
or U610 (N_610,In_541,In_6);
nor U611 (N_611,In_838,In_849);
nand U612 (N_612,In_273,In_667);
and U613 (N_613,In_358,In_115);
and U614 (N_614,In_64,In_283);
nor U615 (N_615,In_996,In_987);
nor U616 (N_616,In_846,In_712);
nand U617 (N_617,In_795,In_390);
nor U618 (N_618,In_813,In_651);
nand U619 (N_619,In_501,In_155);
nor U620 (N_620,In_377,In_637);
nor U621 (N_621,In_604,In_275);
nand U622 (N_622,In_745,In_661);
xnor U623 (N_623,In_300,In_702);
or U624 (N_624,In_386,In_422);
nor U625 (N_625,In_367,In_357);
and U626 (N_626,In_537,In_172);
nand U627 (N_627,In_14,In_541);
nand U628 (N_628,In_793,In_387);
and U629 (N_629,In_174,In_840);
or U630 (N_630,In_32,In_969);
and U631 (N_631,In_562,In_209);
nor U632 (N_632,In_759,In_785);
xnor U633 (N_633,In_636,In_454);
nand U634 (N_634,In_656,In_433);
nand U635 (N_635,In_89,In_799);
nand U636 (N_636,In_582,In_186);
and U637 (N_637,In_375,In_125);
or U638 (N_638,In_887,In_386);
or U639 (N_639,In_40,In_351);
and U640 (N_640,In_960,In_908);
nand U641 (N_641,In_493,In_851);
and U642 (N_642,In_19,In_59);
nand U643 (N_643,In_671,In_76);
or U644 (N_644,In_530,In_665);
and U645 (N_645,In_301,In_437);
nor U646 (N_646,In_275,In_649);
or U647 (N_647,In_641,In_616);
nor U648 (N_648,In_88,In_820);
and U649 (N_649,In_466,In_790);
or U650 (N_650,In_343,In_358);
and U651 (N_651,In_803,In_894);
nand U652 (N_652,In_379,In_436);
nand U653 (N_653,In_899,In_391);
nor U654 (N_654,In_396,In_126);
nor U655 (N_655,In_488,In_918);
and U656 (N_656,In_94,In_200);
nand U657 (N_657,In_932,In_367);
or U658 (N_658,In_177,In_290);
nand U659 (N_659,In_152,In_231);
or U660 (N_660,In_496,In_303);
or U661 (N_661,In_621,In_681);
or U662 (N_662,In_724,In_318);
or U663 (N_663,In_0,In_989);
or U664 (N_664,In_862,In_447);
nor U665 (N_665,In_979,In_931);
nand U666 (N_666,In_718,In_598);
nor U667 (N_667,In_677,In_839);
and U668 (N_668,In_379,In_777);
or U669 (N_669,In_827,In_293);
and U670 (N_670,In_356,In_451);
or U671 (N_671,In_385,In_311);
and U672 (N_672,In_124,In_134);
nor U673 (N_673,In_354,In_811);
or U674 (N_674,In_571,In_739);
or U675 (N_675,In_407,In_24);
and U676 (N_676,In_261,In_348);
and U677 (N_677,In_455,In_818);
nor U678 (N_678,In_519,In_433);
and U679 (N_679,In_462,In_698);
or U680 (N_680,In_170,In_964);
nand U681 (N_681,In_521,In_713);
and U682 (N_682,In_403,In_810);
nand U683 (N_683,In_593,In_437);
nor U684 (N_684,In_197,In_582);
nor U685 (N_685,In_693,In_65);
or U686 (N_686,In_378,In_619);
nor U687 (N_687,In_235,In_436);
nor U688 (N_688,In_593,In_904);
nor U689 (N_689,In_594,In_983);
or U690 (N_690,In_364,In_839);
nand U691 (N_691,In_612,In_852);
nor U692 (N_692,In_916,In_807);
nor U693 (N_693,In_461,In_191);
nor U694 (N_694,In_559,In_81);
nor U695 (N_695,In_476,In_375);
nand U696 (N_696,In_268,In_451);
nor U697 (N_697,In_626,In_990);
and U698 (N_698,In_896,In_386);
and U699 (N_699,In_491,In_266);
or U700 (N_700,In_97,In_526);
or U701 (N_701,In_298,In_870);
or U702 (N_702,In_925,In_753);
or U703 (N_703,In_608,In_486);
or U704 (N_704,In_692,In_735);
nor U705 (N_705,In_138,In_752);
nor U706 (N_706,In_443,In_785);
or U707 (N_707,In_538,In_270);
or U708 (N_708,In_67,In_389);
nand U709 (N_709,In_81,In_125);
and U710 (N_710,In_862,In_161);
nor U711 (N_711,In_40,In_994);
nor U712 (N_712,In_982,In_590);
nor U713 (N_713,In_806,In_93);
nor U714 (N_714,In_643,In_493);
or U715 (N_715,In_291,In_695);
and U716 (N_716,In_496,In_9);
and U717 (N_717,In_670,In_738);
and U718 (N_718,In_161,In_251);
nor U719 (N_719,In_958,In_183);
or U720 (N_720,In_783,In_697);
nor U721 (N_721,In_779,In_194);
and U722 (N_722,In_837,In_685);
nor U723 (N_723,In_336,In_434);
nand U724 (N_724,In_185,In_351);
nor U725 (N_725,In_8,In_262);
and U726 (N_726,In_779,In_580);
or U727 (N_727,In_736,In_867);
and U728 (N_728,In_53,In_638);
or U729 (N_729,In_991,In_867);
nand U730 (N_730,In_280,In_602);
nand U731 (N_731,In_306,In_816);
and U732 (N_732,In_891,In_730);
or U733 (N_733,In_111,In_418);
nand U734 (N_734,In_467,In_37);
nand U735 (N_735,In_613,In_58);
nor U736 (N_736,In_119,In_8);
nor U737 (N_737,In_753,In_599);
nor U738 (N_738,In_92,In_280);
and U739 (N_739,In_544,In_131);
nor U740 (N_740,In_771,In_21);
or U741 (N_741,In_95,In_665);
and U742 (N_742,In_255,In_624);
nor U743 (N_743,In_395,In_972);
nor U744 (N_744,In_318,In_987);
nor U745 (N_745,In_714,In_715);
nand U746 (N_746,In_612,In_988);
and U747 (N_747,In_968,In_507);
nand U748 (N_748,In_544,In_15);
nand U749 (N_749,In_254,In_389);
or U750 (N_750,In_852,In_187);
nand U751 (N_751,In_494,In_154);
nor U752 (N_752,In_541,In_841);
nor U753 (N_753,In_55,In_287);
and U754 (N_754,In_543,In_410);
and U755 (N_755,In_923,In_379);
nand U756 (N_756,In_610,In_733);
or U757 (N_757,In_702,In_84);
or U758 (N_758,In_377,In_430);
nand U759 (N_759,In_323,In_236);
nor U760 (N_760,In_861,In_938);
and U761 (N_761,In_756,In_47);
or U762 (N_762,In_710,In_396);
nand U763 (N_763,In_125,In_768);
or U764 (N_764,In_880,In_160);
or U765 (N_765,In_865,In_491);
and U766 (N_766,In_298,In_330);
nor U767 (N_767,In_922,In_229);
nand U768 (N_768,In_979,In_951);
and U769 (N_769,In_444,In_461);
and U770 (N_770,In_999,In_163);
and U771 (N_771,In_665,In_438);
nor U772 (N_772,In_431,In_568);
and U773 (N_773,In_230,In_952);
or U774 (N_774,In_827,In_862);
or U775 (N_775,In_635,In_319);
nand U776 (N_776,In_153,In_911);
and U777 (N_777,In_210,In_548);
and U778 (N_778,In_725,In_936);
or U779 (N_779,In_275,In_799);
and U780 (N_780,In_65,In_728);
or U781 (N_781,In_771,In_650);
nor U782 (N_782,In_854,In_491);
or U783 (N_783,In_190,In_879);
nor U784 (N_784,In_678,In_300);
nand U785 (N_785,In_219,In_799);
nor U786 (N_786,In_317,In_91);
nand U787 (N_787,In_454,In_122);
or U788 (N_788,In_298,In_892);
and U789 (N_789,In_343,In_420);
and U790 (N_790,In_968,In_899);
or U791 (N_791,In_627,In_436);
or U792 (N_792,In_515,In_588);
or U793 (N_793,In_58,In_48);
and U794 (N_794,In_444,In_383);
and U795 (N_795,In_176,In_731);
xor U796 (N_796,In_3,In_31);
nand U797 (N_797,In_976,In_163);
and U798 (N_798,In_64,In_575);
nand U799 (N_799,In_136,In_707);
nor U800 (N_800,In_146,In_566);
and U801 (N_801,In_799,In_33);
and U802 (N_802,In_325,In_717);
and U803 (N_803,In_763,In_505);
or U804 (N_804,In_99,In_180);
and U805 (N_805,In_205,In_837);
or U806 (N_806,In_306,In_494);
nor U807 (N_807,In_100,In_179);
nand U808 (N_808,In_143,In_421);
or U809 (N_809,In_456,In_31);
nand U810 (N_810,In_157,In_877);
xnor U811 (N_811,In_175,In_999);
nor U812 (N_812,In_883,In_421);
or U813 (N_813,In_554,In_910);
or U814 (N_814,In_77,In_705);
or U815 (N_815,In_289,In_526);
nor U816 (N_816,In_897,In_753);
nor U817 (N_817,In_328,In_912);
nand U818 (N_818,In_68,In_644);
or U819 (N_819,In_99,In_507);
and U820 (N_820,In_623,In_308);
or U821 (N_821,In_499,In_84);
nor U822 (N_822,In_994,In_75);
or U823 (N_823,In_427,In_354);
and U824 (N_824,In_444,In_791);
or U825 (N_825,In_328,In_88);
or U826 (N_826,In_395,In_686);
nand U827 (N_827,In_338,In_512);
or U828 (N_828,In_590,In_415);
nand U829 (N_829,In_824,In_841);
and U830 (N_830,In_745,In_73);
or U831 (N_831,In_900,In_294);
and U832 (N_832,In_605,In_203);
and U833 (N_833,In_307,In_767);
nand U834 (N_834,In_78,In_306);
nand U835 (N_835,In_720,In_408);
nor U836 (N_836,In_594,In_516);
nand U837 (N_837,In_603,In_63);
nor U838 (N_838,In_290,In_636);
nor U839 (N_839,In_142,In_47);
nor U840 (N_840,In_797,In_521);
nand U841 (N_841,In_651,In_850);
or U842 (N_842,In_599,In_39);
or U843 (N_843,In_578,In_72);
or U844 (N_844,In_554,In_964);
nand U845 (N_845,In_160,In_290);
or U846 (N_846,In_263,In_342);
nor U847 (N_847,In_370,In_266);
or U848 (N_848,In_912,In_842);
and U849 (N_849,In_927,In_70);
nor U850 (N_850,In_621,In_841);
nand U851 (N_851,In_63,In_186);
nand U852 (N_852,In_57,In_560);
xnor U853 (N_853,In_635,In_825);
or U854 (N_854,In_376,In_987);
and U855 (N_855,In_590,In_745);
or U856 (N_856,In_248,In_203);
nor U857 (N_857,In_376,In_804);
or U858 (N_858,In_547,In_531);
and U859 (N_859,In_770,In_820);
nand U860 (N_860,In_227,In_290);
or U861 (N_861,In_743,In_307);
nand U862 (N_862,In_671,In_732);
nor U863 (N_863,In_707,In_168);
or U864 (N_864,In_592,In_778);
nor U865 (N_865,In_802,In_27);
nor U866 (N_866,In_94,In_335);
nor U867 (N_867,In_720,In_71);
and U868 (N_868,In_333,In_245);
xor U869 (N_869,In_572,In_516);
and U870 (N_870,In_384,In_132);
and U871 (N_871,In_418,In_669);
or U872 (N_872,In_238,In_785);
nor U873 (N_873,In_208,In_768);
and U874 (N_874,In_450,In_693);
nand U875 (N_875,In_91,In_808);
nor U876 (N_876,In_441,In_861);
and U877 (N_877,In_917,In_284);
nor U878 (N_878,In_837,In_590);
and U879 (N_879,In_35,In_257);
or U880 (N_880,In_606,In_192);
nand U881 (N_881,In_388,In_261);
nand U882 (N_882,In_157,In_677);
nor U883 (N_883,In_238,In_265);
xnor U884 (N_884,In_85,In_360);
nor U885 (N_885,In_725,In_853);
and U886 (N_886,In_232,In_79);
or U887 (N_887,In_499,In_378);
nand U888 (N_888,In_645,In_846);
nand U889 (N_889,In_836,In_500);
nor U890 (N_890,In_408,In_952);
xnor U891 (N_891,In_795,In_62);
and U892 (N_892,In_69,In_507);
nor U893 (N_893,In_756,In_63);
or U894 (N_894,In_270,In_756);
nor U895 (N_895,In_271,In_144);
and U896 (N_896,In_247,In_197);
nor U897 (N_897,In_817,In_984);
nor U898 (N_898,In_436,In_6);
or U899 (N_899,In_182,In_223);
xor U900 (N_900,In_806,In_617);
nor U901 (N_901,In_719,In_821);
nand U902 (N_902,In_859,In_810);
nand U903 (N_903,In_278,In_201);
and U904 (N_904,In_170,In_294);
and U905 (N_905,In_834,In_258);
and U906 (N_906,In_717,In_735);
nor U907 (N_907,In_352,In_697);
nor U908 (N_908,In_452,In_264);
nor U909 (N_909,In_609,In_379);
nand U910 (N_910,In_10,In_303);
or U911 (N_911,In_677,In_242);
or U912 (N_912,In_405,In_253);
and U913 (N_913,In_375,In_248);
nor U914 (N_914,In_589,In_703);
or U915 (N_915,In_978,In_928);
or U916 (N_916,In_912,In_6);
nand U917 (N_917,In_535,In_198);
nand U918 (N_918,In_515,In_506);
and U919 (N_919,In_525,In_54);
nand U920 (N_920,In_788,In_239);
nand U921 (N_921,In_923,In_845);
nor U922 (N_922,In_834,In_121);
nand U923 (N_923,In_650,In_421);
and U924 (N_924,In_127,In_420);
nor U925 (N_925,In_284,In_986);
nand U926 (N_926,In_987,In_58);
or U927 (N_927,In_712,In_648);
and U928 (N_928,In_626,In_715);
and U929 (N_929,In_154,In_513);
and U930 (N_930,In_856,In_854);
nand U931 (N_931,In_295,In_244);
nand U932 (N_932,In_452,In_56);
nand U933 (N_933,In_432,In_47);
nor U934 (N_934,In_248,In_924);
and U935 (N_935,In_971,In_621);
xor U936 (N_936,In_120,In_849);
nand U937 (N_937,In_48,In_148);
or U938 (N_938,In_978,In_977);
nand U939 (N_939,In_255,In_462);
nand U940 (N_940,In_65,In_596);
and U941 (N_941,In_394,In_28);
and U942 (N_942,In_466,In_705);
or U943 (N_943,In_32,In_112);
nor U944 (N_944,In_200,In_609);
and U945 (N_945,In_552,In_402);
nand U946 (N_946,In_150,In_136);
and U947 (N_947,In_333,In_767);
nand U948 (N_948,In_241,In_93);
and U949 (N_949,In_452,In_946);
nor U950 (N_950,In_729,In_985);
nand U951 (N_951,In_169,In_80);
nor U952 (N_952,In_63,In_626);
xnor U953 (N_953,In_768,In_481);
or U954 (N_954,In_749,In_826);
and U955 (N_955,In_983,In_841);
and U956 (N_956,In_388,In_631);
nor U957 (N_957,In_160,In_999);
xnor U958 (N_958,In_598,In_545);
and U959 (N_959,In_250,In_802);
nor U960 (N_960,In_482,In_276);
and U961 (N_961,In_69,In_47);
and U962 (N_962,In_438,In_367);
or U963 (N_963,In_644,In_948);
nand U964 (N_964,In_248,In_238);
nor U965 (N_965,In_843,In_565);
and U966 (N_966,In_735,In_541);
nand U967 (N_967,In_161,In_306);
or U968 (N_968,In_219,In_680);
nor U969 (N_969,In_419,In_749);
and U970 (N_970,In_701,In_419);
and U971 (N_971,In_580,In_933);
and U972 (N_972,In_494,In_23);
or U973 (N_973,In_578,In_532);
and U974 (N_974,In_730,In_303);
nor U975 (N_975,In_252,In_148);
nand U976 (N_976,In_874,In_990);
nand U977 (N_977,In_48,In_681);
nand U978 (N_978,In_577,In_348);
nand U979 (N_979,In_122,In_894);
and U980 (N_980,In_600,In_279);
nand U981 (N_981,In_427,In_973);
and U982 (N_982,In_416,In_956);
or U983 (N_983,In_488,In_643);
nand U984 (N_984,In_242,In_917);
nand U985 (N_985,In_368,In_569);
nor U986 (N_986,In_4,In_473);
nor U987 (N_987,In_274,In_53);
and U988 (N_988,In_768,In_460);
nand U989 (N_989,In_106,In_225);
nor U990 (N_990,In_340,In_56);
or U991 (N_991,In_381,In_708);
and U992 (N_992,In_32,In_808);
and U993 (N_993,In_327,In_591);
and U994 (N_994,In_601,In_700);
nand U995 (N_995,In_85,In_172);
and U996 (N_996,In_596,In_645);
and U997 (N_997,In_797,In_252);
and U998 (N_998,In_518,In_934);
and U999 (N_999,In_948,In_215);
and U1000 (N_1000,In_937,In_993);
nor U1001 (N_1001,In_194,In_898);
and U1002 (N_1002,In_603,In_462);
nor U1003 (N_1003,In_516,In_713);
or U1004 (N_1004,In_800,In_778);
nor U1005 (N_1005,In_995,In_340);
nand U1006 (N_1006,In_379,In_644);
or U1007 (N_1007,In_23,In_8);
nor U1008 (N_1008,In_319,In_770);
or U1009 (N_1009,In_761,In_497);
and U1010 (N_1010,In_582,In_919);
and U1011 (N_1011,In_562,In_639);
and U1012 (N_1012,In_356,In_794);
nor U1013 (N_1013,In_192,In_586);
or U1014 (N_1014,In_252,In_138);
nand U1015 (N_1015,In_975,In_729);
and U1016 (N_1016,In_934,In_223);
nand U1017 (N_1017,In_722,In_846);
and U1018 (N_1018,In_495,In_804);
or U1019 (N_1019,In_73,In_156);
or U1020 (N_1020,In_240,In_324);
or U1021 (N_1021,In_540,In_5);
and U1022 (N_1022,In_576,In_156);
xnor U1023 (N_1023,In_664,In_584);
nand U1024 (N_1024,In_391,In_942);
or U1025 (N_1025,In_415,In_105);
and U1026 (N_1026,In_371,In_497);
or U1027 (N_1027,In_383,In_713);
and U1028 (N_1028,In_376,In_563);
and U1029 (N_1029,In_613,In_276);
nor U1030 (N_1030,In_964,In_637);
and U1031 (N_1031,In_852,In_46);
or U1032 (N_1032,In_728,In_877);
nor U1033 (N_1033,In_229,In_152);
nand U1034 (N_1034,In_669,In_334);
and U1035 (N_1035,In_781,In_416);
nand U1036 (N_1036,In_258,In_186);
or U1037 (N_1037,In_793,In_151);
xnor U1038 (N_1038,In_696,In_498);
nor U1039 (N_1039,In_933,In_680);
and U1040 (N_1040,In_291,In_216);
or U1041 (N_1041,In_343,In_14);
nand U1042 (N_1042,In_482,In_85);
or U1043 (N_1043,In_437,In_653);
nor U1044 (N_1044,In_607,In_569);
nand U1045 (N_1045,In_986,In_344);
and U1046 (N_1046,In_630,In_211);
and U1047 (N_1047,In_587,In_148);
xnor U1048 (N_1048,In_822,In_309);
nand U1049 (N_1049,In_611,In_994);
nor U1050 (N_1050,In_942,In_171);
or U1051 (N_1051,In_982,In_540);
nor U1052 (N_1052,In_72,In_222);
and U1053 (N_1053,In_9,In_784);
nor U1054 (N_1054,In_939,In_128);
nor U1055 (N_1055,In_281,In_499);
nor U1056 (N_1056,In_836,In_380);
and U1057 (N_1057,In_735,In_118);
nor U1058 (N_1058,In_616,In_83);
nor U1059 (N_1059,In_705,In_825);
nor U1060 (N_1060,In_111,In_899);
and U1061 (N_1061,In_786,In_376);
or U1062 (N_1062,In_645,In_144);
and U1063 (N_1063,In_412,In_653);
nor U1064 (N_1064,In_154,In_471);
nor U1065 (N_1065,In_267,In_911);
and U1066 (N_1066,In_434,In_139);
nor U1067 (N_1067,In_728,In_994);
or U1068 (N_1068,In_519,In_30);
and U1069 (N_1069,In_533,In_559);
or U1070 (N_1070,In_784,In_190);
or U1071 (N_1071,In_827,In_424);
and U1072 (N_1072,In_994,In_762);
and U1073 (N_1073,In_883,In_438);
or U1074 (N_1074,In_743,In_824);
nor U1075 (N_1075,In_960,In_456);
nor U1076 (N_1076,In_697,In_709);
or U1077 (N_1077,In_348,In_919);
nand U1078 (N_1078,In_619,In_415);
nand U1079 (N_1079,In_831,In_345);
nand U1080 (N_1080,In_175,In_144);
or U1081 (N_1081,In_195,In_673);
or U1082 (N_1082,In_369,In_34);
and U1083 (N_1083,In_237,In_216);
or U1084 (N_1084,In_742,In_186);
nor U1085 (N_1085,In_402,In_156);
and U1086 (N_1086,In_186,In_520);
and U1087 (N_1087,In_23,In_92);
xnor U1088 (N_1088,In_453,In_401);
nor U1089 (N_1089,In_653,In_626);
and U1090 (N_1090,In_344,In_229);
nand U1091 (N_1091,In_755,In_751);
or U1092 (N_1092,In_992,In_960);
or U1093 (N_1093,In_143,In_969);
nor U1094 (N_1094,In_175,In_960);
nor U1095 (N_1095,In_925,In_958);
or U1096 (N_1096,In_643,In_793);
nor U1097 (N_1097,In_633,In_33);
nor U1098 (N_1098,In_287,In_644);
nand U1099 (N_1099,In_940,In_320);
nor U1100 (N_1100,In_271,In_468);
nor U1101 (N_1101,In_556,In_467);
or U1102 (N_1102,In_550,In_150);
or U1103 (N_1103,In_757,In_331);
and U1104 (N_1104,In_353,In_617);
nor U1105 (N_1105,In_482,In_8);
nor U1106 (N_1106,In_166,In_545);
xnor U1107 (N_1107,In_218,In_827);
and U1108 (N_1108,In_672,In_719);
xor U1109 (N_1109,In_734,In_60);
nor U1110 (N_1110,In_345,In_261);
nor U1111 (N_1111,In_703,In_858);
or U1112 (N_1112,In_818,In_342);
and U1113 (N_1113,In_583,In_739);
nand U1114 (N_1114,In_778,In_297);
nand U1115 (N_1115,In_436,In_660);
and U1116 (N_1116,In_622,In_225);
and U1117 (N_1117,In_352,In_676);
and U1118 (N_1118,In_9,In_160);
nor U1119 (N_1119,In_210,In_383);
and U1120 (N_1120,In_669,In_207);
nor U1121 (N_1121,In_588,In_168);
nor U1122 (N_1122,In_681,In_591);
or U1123 (N_1123,In_305,In_431);
or U1124 (N_1124,In_443,In_132);
nor U1125 (N_1125,In_627,In_807);
nand U1126 (N_1126,In_571,In_657);
and U1127 (N_1127,In_829,In_270);
nor U1128 (N_1128,In_955,In_794);
or U1129 (N_1129,In_308,In_35);
nor U1130 (N_1130,In_390,In_114);
or U1131 (N_1131,In_427,In_22);
or U1132 (N_1132,In_772,In_105);
or U1133 (N_1133,In_220,In_472);
nor U1134 (N_1134,In_618,In_803);
nand U1135 (N_1135,In_255,In_274);
nand U1136 (N_1136,In_751,In_162);
nor U1137 (N_1137,In_204,In_779);
and U1138 (N_1138,In_730,In_175);
and U1139 (N_1139,In_863,In_489);
and U1140 (N_1140,In_443,In_458);
and U1141 (N_1141,In_794,In_650);
nor U1142 (N_1142,In_89,In_545);
nor U1143 (N_1143,In_79,In_94);
and U1144 (N_1144,In_682,In_112);
or U1145 (N_1145,In_445,In_834);
nor U1146 (N_1146,In_784,In_19);
nor U1147 (N_1147,In_796,In_529);
xor U1148 (N_1148,In_819,In_122);
nand U1149 (N_1149,In_531,In_785);
or U1150 (N_1150,In_186,In_84);
nor U1151 (N_1151,In_481,In_450);
nor U1152 (N_1152,In_704,In_222);
nand U1153 (N_1153,In_676,In_563);
nor U1154 (N_1154,In_158,In_795);
or U1155 (N_1155,In_890,In_105);
nand U1156 (N_1156,In_651,In_117);
or U1157 (N_1157,In_822,In_299);
and U1158 (N_1158,In_588,In_565);
and U1159 (N_1159,In_123,In_457);
nor U1160 (N_1160,In_500,In_124);
or U1161 (N_1161,In_143,In_47);
or U1162 (N_1162,In_568,In_955);
nand U1163 (N_1163,In_838,In_495);
and U1164 (N_1164,In_520,In_480);
nor U1165 (N_1165,In_679,In_48);
nor U1166 (N_1166,In_423,In_926);
and U1167 (N_1167,In_92,In_957);
or U1168 (N_1168,In_970,In_73);
and U1169 (N_1169,In_435,In_746);
and U1170 (N_1170,In_142,In_865);
nor U1171 (N_1171,In_267,In_281);
or U1172 (N_1172,In_988,In_454);
nand U1173 (N_1173,In_773,In_105);
and U1174 (N_1174,In_966,In_252);
or U1175 (N_1175,In_373,In_5);
nand U1176 (N_1176,In_516,In_821);
nand U1177 (N_1177,In_231,In_831);
nand U1178 (N_1178,In_468,In_20);
nand U1179 (N_1179,In_618,In_785);
nand U1180 (N_1180,In_267,In_859);
nand U1181 (N_1181,In_967,In_711);
or U1182 (N_1182,In_666,In_511);
nand U1183 (N_1183,In_634,In_755);
nor U1184 (N_1184,In_554,In_116);
nand U1185 (N_1185,In_233,In_222);
and U1186 (N_1186,In_847,In_910);
and U1187 (N_1187,In_692,In_687);
xor U1188 (N_1188,In_279,In_575);
nor U1189 (N_1189,In_905,In_317);
and U1190 (N_1190,In_883,In_670);
or U1191 (N_1191,In_856,In_414);
or U1192 (N_1192,In_86,In_517);
or U1193 (N_1193,In_286,In_541);
and U1194 (N_1194,In_482,In_869);
nand U1195 (N_1195,In_138,In_444);
and U1196 (N_1196,In_444,In_577);
and U1197 (N_1197,In_708,In_812);
nand U1198 (N_1198,In_131,In_690);
and U1199 (N_1199,In_460,In_762);
or U1200 (N_1200,In_623,In_664);
or U1201 (N_1201,In_953,In_770);
nor U1202 (N_1202,In_914,In_766);
nand U1203 (N_1203,In_21,In_901);
or U1204 (N_1204,In_690,In_501);
nor U1205 (N_1205,In_457,In_693);
nand U1206 (N_1206,In_265,In_922);
or U1207 (N_1207,In_740,In_489);
nor U1208 (N_1208,In_122,In_165);
and U1209 (N_1209,In_86,In_884);
and U1210 (N_1210,In_873,In_624);
or U1211 (N_1211,In_885,In_671);
nor U1212 (N_1212,In_199,In_910);
and U1213 (N_1213,In_807,In_200);
nor U1214 (N_1214,In_139,In_946);
nand U1215 (N_1215,In_452,In_503);
or U1216 (N_1216,In_180,In_737);
or U1217 (N_1217,In_213,In_944);
and U1218 (N_1218,In_844,In_117);
or U1219 (N_1219,In_159,In_110);
nor U1220 (N_1220,In_439,In_63);
nand U1221 (N_1221,In_629,In_922);
nand U1222 (N_1222,In_576,In_177);
nor U1223 (N_1223,In_996,In_378);
and U1224 (N_1224,In_723,In_929);
or U1225 (N_1225,In_688,In_655);
or U1226 (N_1226,In_668,In_304);
nor U1227 (N_1227,In_1,In_21);
or U1228 (N_1228,In_798,In_766);
nor U1229 (N_1229,In_144,In_731);
nand U1230 (N_1230,In_113,In_732);
nand U1231 (N_1231,In_145,In_200);
and U1232 (N_1232,In_545,In_242);
nor U1233 (N_1233,In_82,In_635);
and U1234 (N_1234,In_390,In_58);
and U1235 (N_1235,In_931,In_626);
nor U1236 (N_1236,In_771,In_447);
or U1237 (N_1237,In_383,In_331);
nor U1238 (N_1238,In_960,In_544);
nor U1239 (N_1239,In_990,In_317);
or U1240 (N_1240,In_870,In_740);
xnor U1241 (N_1241,In_851,In_838);
and U1242 (N_1242,In_441,In_134);
and U1243 (N_1243,In_532,In_336);
and U1244 (N_1244,In_276,In_848);
and U1245 (N_1245,In_2,In_935);
nor U1246 (N_1246,In_721,In_849);
and U1247 (N_1247,In_387,In_925);
nand U1248 (N_1248,In_451,In_50);
nand U1249 (N_1249,In_829,In_601);
and U1250 (N_1250,In_310,In_935);
nand U1251 (N_1251,In_729,In_466);
or U1252 (N_1252,In_338,In_94);
or U1253 (N_1253,In_675,In_967);
xnor U1254 (N_1254,In_945,In_713);
and U1255 (N_1255,In_771,In_787);
nand U1256 (N_1256,In_285,In_784);
and U1257 (N_1257,In_439,In_490);
nand U1258 (N_1258,In_394,In_113);
and U1259 (N_1259,In_51,In_177);
nor U1260 (N_1260,In_440,In_615);
nor U1261 (N_1261,In_559,In_608);
nor U1262 (N_1262,In_689,In_493);
nand U1263 (N_1263,In_337,In_950);
and U1264 (N_1264,In_437,In_960);
nor U1265 (N_1265,In_290,In_269);
nand U1266 (N_1266,In_593,In_261);
or U1267 (N_1267,In_24,In_282);
or U1268 (N_1268,In_199,In_805);
nand U1269 (N_1269,In_171,In_286);
nand U1270 (N_1270,In_717,In_109);
or U1271 (N_1271,In_455,In_442);
and U1272 (N_1272,In_959,In_47);
and U1273 (N_1273,In_527,In_320);
nand U1274 (N_1274,In_707,In_566);
and U1275 (N_1275,In_437,In_677);
or U1276 (N_1276,In_498,In_154);
and U1277 (N_1277,In_723,In_83);
xor U1278 (N_1278,In_203,In_201);
or U1279 (N_1279,In_773,In_981);
nand U1280 (N_1280,In_880,In_929);
and U1281 (N_1281,In_539,In_156);
or U1282 (N_1282,In_361,In_554);
or U1283 (N_1283,In_231,In_920);
nand U1284 (N_1284,In_794,In_515);
nor U1285 (N_1285,In_65,In_17);
nor U1286 (N_1286,In_959,In_467);
nand U1287 (N_1287,In_570,In_783);
xor U1288 (N_1288,In_570,In_786);
or U1289 (N_1289,In_763,In_325);
and U1290 (N_1290,In_487,In_625);
xor U1291 (N_1291,In_759,In_699);
nor U1292 (N_1292,In_451,In_139);
nor U1293 (N_1293,In_741,In_965);
nand U1294 (N_1294,In_376,In_921);
and U1295 (N_1295,In_935,In_106);
or U1296 (N_1296,In_977,In_88);
xor U1297 (N_1297,In_409,In_935);
or U1298 (N_1298,In_842,In_846);
and U1299 (N_1299,In_287,In_865);
and U1300 (N_1300,In_415,In_896);
or U1301 (N_1301,In_848,In_800);
nand U1302 (N_1302,In_936,In_127);
and U1303 (N_1303,In_667,In_190);
and U1304 (N_1304,In_972,In_486);
and U1305 (N_1305,In_80,In_468);
nor U1306 (N_1306,In_858,In_219);
nor U1307 (N_1307,In_311,In_895);
nand U1308 (N_1308,In_576,In_454);
nand U1309 (N_1309,In_742,In_430);
and U1310 (N_1310,In_943,In_207);
and U1311 (N_1311,In_778,In_80);
nor U1312 (N_1312,In_585,In_135);
nand U1313 (N_1313,In_408,In_881);
xnor U1314 (N_1314,In_334,In_140);
nand U1315 (N_1315,In_8,In_40);
or U1316 (N_1316,In_611,In_679);
or U1317 (N_1317,In_78,In_71);
and U1318 (N_1318,In_653,In_880);
nor U1319 (N_1319,In_432,In_873);
nor U1320 (N_1320,In_890,In_286);
nand U1321 (N_1321,In_480,In_177);
nand U1322 (N_1322,In_281,In_212);
nor U1323 (N_1323,In_878,In_835);
or U1324 (N_1324,In_138,In_753);
or U1325 (N_1325,In_84,In_492);
nand U1326 (N_1326,In_723,In_40);
nand U1327 (N_1327,In_344,In_709);
or U1328 (N_1328,In_106,In_989);
nor U1329 (N_1329,In_193,In_476);
nand U1330 (N_1330,In_682,In_270);
nor U1331 (N_1331,In_477,In_83);
and U1332 (N_1332,In_627,In_865);
or U1333 (N_1333,In_34,In_549);
nand U1334 (N_1334,In_46,In_300);
or U1335 (N_1335,In_911,In_29);
or U1336 (N_1336,In_288,In_678);
nand U1337 (N_1337,In_523,In_24);
nand U1338 (N_1338,In_754,In_491);
nor U1339 (N_1339,In_638,In_164);
and U1340 (N_1340,In_396,In_299);
nor U1341 (N_1341,In_810,In_517);
nand U1342 (N_1342,In_541,In_138);
nand U1343 (N_1343,In_234,In_759);
or U1344 (N_1344,In_626,In_85);
and U1345 (N_1345,In_648,In_49);
nor U1346 (N_1346,In_508,In_288);
and U1347 (N_1347,In_617,In_604);
nand U1348 (N_1348,In_266,In_24);
and U1349 (N_1349,In_378,In_751);
nor U1350 (N_1350,In_476,In_414);
nor U1351 (N_1351,In_389,In_120);
nor U1352 (N_1352,In_940,In_571);
nand U1353 (N_1353,In_801,In_418);
or U1354 (N_1354,In_839,In_829);
and U1355 (N_1355,In_459,In_413);
xor U1356 (N_1356,In_218,In_776);
nand U1357 (N_1357,In_437,In_121);
nor U1358 (N_1358,In_230,In_111);
and U1359 (N_1359,In_26,In_776);
nand U1360 (N_1360,In_788,In_740);
or U1361 (N_1361,In_173,In_566);
or U1362 (N_1362,In_441,In_552);
nor U1363 (N_1363,In_189,In_564);
nor U1364 (N_1364,In_993,In_67);
nand U1365 (N_1365,In_971,In_474);
or U1366 (N_1366,In_243,In_662);
and U1367 (N_1367,In_524,In_861);
nor U1368 (N_1368,In_987,In_636);
and U1369 (N_1369,In_452,In_74);
and U1370 (N_1370,In_617,In_913);
and U1371 (N_1371,In_34,In_739);
and U1372 (N_1372,In_408,In_467);
and U1373 (N_1373,In_614,In_860);
nor U1374 (N_1374,In_419,In_537);
nand U1375 (N_1375,In_840,In_576);
nand U1376 (N_1376,In_955,In_677);
nand U1377 (N_1377,In_245,In_204);
nand U1378 (N_1378,In_966,In_683);
nand U1379 (N_1379,In_976,In_181);
nor U1380 (N_1380,In_162,In_400);
xnor U1381 (N_1381,In_37,In_107);
nand U1382 (N_1382,In_548,In_602);
or U1383 (N_1383,In_194,In_28);
and U1384 (N_1384,In_795,In_76);
nor U1385 (N_1385,In_469,In_555);
nand U1386 (N_1386,In_727,In_45);
nand U1387 (N_1387,In_616,In_485);
and U1388 (N_1388,In_283,In_520);
and U1389 (N_1389,In_640,In_385);
and U1390 (N_1390,In_991,In_902);
or U1391 (N_1391,In_393,In_114);
nand U1392 (N_1392,In_825,In_509);
and U1393 (N_1393,In_574,In_769);
nand U1394 (N_1394,In_34,In_980);
and U1395 (N_1395,In_968,In_615);
and U1396 (N_1396,In_170,In_211);
or U1397 (N_1397,In_692,In_996);
nor U1398 (N_1398,In_821,In_584);
xor U1399 (N_1399,In_903,In_839);
and U1400 (N_1400,In_5,In_460);
xor U1401 (N_1401,In_943,In_592);
or U1402 (N_1402,In_152,In_359);
nand U1403 (N_1403,In_108,In_516);
nor U1404 (N_1404,In_952,In_856);
nor U1405 (N_1405,In_656,In_748);
or U1406 (N_1406,In_374,In_871);
nand U1407 (N_1407,In_400,In_245);
nor U1408 (N_1408,In_411,In_584);
and U1409 (N_1409,In_683,In_300);
or U1410 (N_1410,In_456,In_169);
nand U1411 (N_1411,In_109,In_126);
nand U1412 (N_1412,In_598,In_311);
nor U1413 (N_1413,In_103,In_850);
nand U1414 (N_1414,In_706,In_732);
and U1415 (N_1415,In_89,In_283);
and U1416 (N_1416,In_841,In_888);
or U1417 (N_1417,In_442,In_113);
or U1418 (N_1418,In_289,In_365);
and U1419 (N_1419,In_292,In_888);
nor U1420 (N_1420,In_571,In_797);
nor U1421 (N_1421,In_345,In_687);
nand U1422 (N_1422,In_81,In_587);
nand U1423 (N_1423,In_9,In_122);
or U1424 (N_1424,In_719,In_153);
or U1425 (N_1425,In_254,In_513);
or U1426 (N_1426,In_985,In_371);
nand U1427 (N_1427,In_737,In_330);
and U1428 (N_1428,In_430,In_483);
nor U1429 (N_1429,In_659,In_31);
or U1430 (N_1430,In_736,In_616);
nand U1431 (N_1431,In_720,In_713);
and U1432 (N_1432,In_215,In_972);
nor U1433 (N_1433,In_788,In_927);
or U1434 (N_1434,In_571,In_516);
and U1435 (N_1435,In_135,In_42);
or U1436 (N_1436,In_163,In_446);
and U1437 (N_1437,In_335,In_419);
or U1438 (N_1438,In_334,In_451);
nand U1439 (N_1439,In_514,In_51);
nand U1440 (N_1440,In_506,In_730);
and U1441 (N_1441,In_36,In_833);
nand U1442 (N_1442,In_262,In_956);
or U1443 (N_1443,In_701,In_44);
nand U1444 (N_1444,In_774,In_889);
or U1445 (N_1445,In_857,In_942);
or U1446 (N_1446,In_394,In_976);
and U1447 (N_1447,In_865,In_763);
nor U1448 (N_1448,In_23,In_391);
nand U1449 (N_1449,In_9,In_583);
xnor U1450 (N_1450,In_301,In_396);
nand U1451 (N_1451,In_855,In_266);
or U1452 (N_1452,In_534,In_467);
nor U1453 (N_1453,In_859,In_326);
and U1454 (N_1454,In_435,In_239);
or U1455 (N_1455,In_29,In_804);
nor U1456 (N_1456,In_616,In_633);
nor U1457 (N_1457,In_68,In_591);
nor U1458 (N_1458,In_930,In_899);
and U1459 (N_1459,In_246,In_672);
nand U1460 (N_1460,In_965,In_419);
nor U1461 (N_1461,In_214,In_650);
or U1462 (N_1462,In_616,In_614);
and U1463 (N_1463,In_42,In_513);
or U1464 (N_1464,In_289,In_624);
nor U1465 (N_1465,In_934,In_584);
nand U1466 (N_1466,In_439,In_791);
nand U1467 (N_1467,In_690,In_868);
or U1468 (N_1468,In_857,In_584);
and U1469 (N_1469,In_791,In_47);
or U1470 (N_1470,In_14,In_525);
nand U1471 (N_1471,In_394,In_914);
or U1472 (N_1472,In_977,In_102);
nand U1473 (N_1473,In_571,In_659);
and U1474 (N_1474,In_248,In_480);
nand U1475 (N_1475,In_484,In_743);
or U1476 (N_1476,In_508,In_958);
nor U1477 (N_1477,In_996,In_321);
or U1478 (N_1478,In_379,In_949);
or U1479 (N_1479,In_492,In_919);
or U1480 (N_1480,In_871,In_168);
nand U1481 (N_1481,In_784,In_820);
and U1482 (N_1482,In_948,In_317);
nand U1483 (N_1483,In_759,In_564);
or U1484 (N_1484,In_700,In_795);
and U1485 (N_1485,In_421,In_685);
nand U1486 (N_1486,In_410,In_681);
and U1487 (N_1487,In_158,In_208);
nand U1488 (N_1488,In_270,In_844);
and U1489 (N_1489,In_137,In_925);
nor U1490 (N_1490,In_104,In_823);
xor U1491 (N_1491,In_281,In_703);
and U1492 (N_1492,In_589,In_740);
nand U1493 (N_1493,In_497,In_22);
and U1494 (N_1494,In_906,In_692);
and U1495 (N_1495,In_277,In_369);
or U1496 (N_1496,In_639,In_679);
or U1497 (N_1497,In_651,In_958);
nand U1498 (N_1498,In_403,In_629);
or U1499 (N_1499,In_96,In_49);
or U1500 (N_1500,In_666,In_638);
and U1501 (N_1501,In_253,In_491);
and U1502 (N_1502,In_461,In_128);
and U1503 (N_1503,In_254,In_888);
nor U1504 (N_1504,In_159,In_499);
nor U1505 (N_1505,In_153,In_518);
and U1506 (N_1506,In_999,In_501);
and U1507 (N_1507,In_634,In_188);
and U1508 (N_1508,In_484,In_740);
and U1509 (N_1509,In_314,In_651);
or U1510 (N_1510,In_159,In_342);
nand U1511 (N_1511,In_244,In_306);
or U1512 (N_1512,In_805,In_423);
and U1513 (N_1513,In_263,In_678);
or U1514 (N_1514,In_4,In_79);
and U1515 (N_1515,In_707,In_459);
nor U1516 (N_1516,In_180,In_826);
or U1517 (N_1517,In_425,In_357);
or U1518 (N_1518,In_519,In_699);
and U1519 (N_1519,In_277,In_425);
nor U1520 (N_1520,In_727,In_740);
nand U1521 (N_1521,In_754,In_277);
nand U1522 (N_1522,In_805,In_927);
nor U1523 (N_1523,In_608,In_142);
and U1524 (N_1524,In_412,In_808);
nor U1525 (N_1525,In_904,In_74);
or U1526 (N_1526,In_905,In_527);
and U1527 (N_1527,In_510,In_329);
nor U1528 (N_1528,In_264,In_147);
nor U1529 (N_1529,In_422,In_244);
nand U1530 (N_1530,In_688,In_564);
or U1531 (N_1531,In_523,In_642);
nor U1532 (N_1532,In_919,In_314);
nor U1533 (N_1533,In_547,In_897);
nand U1534 (N_1534,In_444,In_566);
nor U1535 (N_1535,In_234,In_532);
and U1536 (N_1536,In_12,In_695);
nor U1537 (N_1537,In_13,In_567);
or U1538 (N_1538,In_712,In_401);
nor U1539 (N_1539,In_288,In_709);
nor U1540 (N_1540,In_821,In_827);
xor U1541 (N_1541,In_145,In_462);
and U1542 (N_1542,In_8,In_11);
and U1543 (N_1543,In_522,In_752);
nand U1544 (N_1544,In_202,In_513);
nand U1545 (N_1545,In_958,In_2);
or U1546 (N_1546,In_214,In_718);
or U1547 (N_1547,In_526,In_936);
or U1548 (N_1548,In_677,In_899);
and U1549 (N_1549,In_545,In_540);
or U1550 (N_1550,In_87,In_169);
or U1551 (N_1551,In_894,In_772);
nand U1552 (N_1552,In_566,In_571);
nor U1553 (N_1553,In_375,In_983);
and U1554 (N_1554,In_131,In_565);
nor U1555 (N_1555,In_862,In_582);
nand U1556 (N_1556,In_798,In_657);
nand U1557 (N_1557,In_146,In_791);
nand U1558 (N_1558,In_690,In_975);
nand U1559 (N_1559,In_17,In_884);
or U1560 (N_1560,In_645,In_453);
or U1561 (N_1561,In_530,In_333);
or U1562 (N_1562,In_214,In_570);
nand U1563 (N_1563,In_650,In_234);
xnor U1564 (N_1564,In_792,In_371);
nand U1565 (N_1565,In_184,In_137);
nor U1566 (N_1566,In_562,In_437);
nor U1567 (N_1567,In_812,In_202);
or U1568 (N_1568,In_263,In_18);
nor U1569 (N_1569,In_54,In_586);
nand U1570 (N_1570,In_226,In_897);
or U1571 (N_1571,In_352,In_191);
and U1572 (N_1572,In_732,In_159);
nor U1573 (N_1573,In_652,In_382);
or U1574 (N_1574,In_935,In_204);
or U1575 (N_1575,In_67,In_107);
xor U1576 (N_1576,In_572,In_599);
nand U1577 (N_1577,In_16,In_924);
nand U1578 (N_1578,In_710,In_275);
and U1579 (N_1579,In_196,In_409);
nand U1580 (N_1580,In_882,In_987);
or U1581 (N_1581,In_669,In_769);
nand U1582 (N_1582,In_931,In_634);
nand U1583 (N_1583,In_715,In_770);
nor U1584 (N_1584,In_548,In_704);
nand U1585 (N_1585,In_684,In_196);
nor U1586 (N_1586,In_242,In_751);
nor U1587 (N_1587,In_97,In_738);
and U1588 (N_1588,In_522,In_237);
or U1589 (N_1589,In_225,In_119);
nand U1590 (N_1590,In_416,In_803);
nor U1591 (N_1591,In_234,In_444);
and U1592 (N_1592,In_327,In_600);
xor U1593 (N_1593,In_688,In_991);
nor U1594 (N_1594,In_689,In_76);
nand U1595 (N_1595,In_295,In_652);
or U1596 (N_1596,In_955,In_303);
or U1597 (N_1597,In_665,In_270);
and U1598 (N_1598,In_363,In_685);
nand U1599 (N_1599,In_857,In_92);
or U1600 (N_1600,In_275,In_594);
nand U1601 (N_1601,In_621,In_632);
nand U1602 (N_1602,In_275,In_30);
or U1603 (N_1603,In_494,In_388);
and U1604 (N_1604,In_798,In_928);
nand U1605 (N_1605,In_777,In_751);
nor U1606 (N_1606,In_82,In_200);
xnor U1607 (N_1607,In_979,In_706);
and U1608 (N_1608,In_544,In_880);
and U1609 (N_1609,In_255,In_690);
or U1610 (N_1610,In_716,In_674);
and U1611 (N_1611,In_475,In_687);
nand U1612 (N_1612,In_499,In_36);
and U1613 (N_1613,In_954,In_425);
or U1614 (N_1614,In_438,In_301);
nand U1615 (N_1615,In_110,In_669);
or U1616 (N_1616,In_9,In_870);
and U1617 (N_1617,In_448,In_990);
nor U1618 (N_1618,In_806,In_215);
and U1619 (N_1619,In_361,In_100);
or U1620 (N_1620,In_494,In_493);
nand U1621 (N_1621,In_384,In_423);
and U1622 (N_1622,In_386,In_568);
or U1623 (N_1623,In_815,In_447);
and U1624 (N_1624,In_215,In_868);
nand U1625 (N_1625,In_982,In_781);
and U1626 (N_1626,In_576,In_427);
and U1627 (N_1627,In_755,In_69);
or U1628 (N_1628,In_965,In_341);
or U1629 (N_1629,In_691,In_122);
nand U1630 (N_1630,In_215,In_432);
nor U1631 (N_1631,In_701,In_56);
nor U1632 (N_1632,In_674,In_774);
and U1633 (N_1633,In_94,In_489);
nand U1634 (N_1634,In_900,In_474);
nor U1635 (N_1635,In_300,In_645);
and U1636 (N_1636,In_624,In_66);
and U1637 (N_1637,In_407,In_451);
nand U1638 (N_1638,In_170,In_968);
nand U1639 (N_1639,In_184,In_220);
nand U1640 (N_1640,In_953,In_448);
nand U1641 (N_1641,In_230,In_568);
and U1642 (N_1642,In_589,In_264);
nor U1643 (N_1643,In_330,In_151);
and U1644 (N_1644,In_338,In_452);
or U1645 (N_1645,In_538,In_296);
nor U1646 (N_1646,In_746,In_286);
or U1647 (N_1647,In_144,In_494);
and U1648 (N_1648,In_524,In_235);
xor U1649 (N_1649,In_785,In_975);
or U1650 (N_1650,In_801,In_90);
nor U1651 (N_1651,In_804,In_842);
xor U1652 (N_1652,In_167,In_929);
nor U1653 (N_1653,In_528,In_520);
nor U1654 (N_1654,In_193,In_927);
nand U1655 (N_1655,In_546,In_436);
nand U1656 (N_1656,In_965,In_709);
nor U1657 (N_1657,In_161,In_727);
or U1658 (N_1658,In_784,In_531);
or U1659 (N_1659,In_460,In_401);
nor U1660 (N_1660,In_246,In_609);
nor U1661 (N_1661,In_308,In_926);
and U1662 (N_1662,In_294,In_855);
and U1663 (N_1663,In_329,In_709);
or U1664 (N_1664,In_108,In_189);
nand U1665 (N_1665,In_742,In_265);
or U1666 (N_1666,In_694,In_703);
nor U1667 (N_1667,In_773,In_859);
and U1668 (N_1668,In_543,In_565);
and U1669 (N_1669,In_433,In_814);
and U1670 (N_1670,In_141,In_894);
xor U1671 (N_1671,In_292,In_902);
xor U1672 (N_1672,In_408,In_51);
nor U1673 (N_1673,In_395,In_618);
or U1674 (N_1674,In_719,In_892);
nand U1675 (N_1675,In_671,In_70);
and U1676 (N_1676,In_356,In_447);
or U1677 (N_1677,In_942,In_398);
nand U1678 (N_1678,In_365,In_214);
or U1679 (N_1679,In_653,In_758);
nand U1680 (N_1680,In_487,In_428);
and U1681 (N_1681,In_577,In_472);
or U1682 (N_1682,In_305,In_89);
or U1683 (N_1683,In_503,In_276);
nor U1684 (N_1684,In_45,In_250);
nand U1685 (N_1685,In_58,In_441);
and U1686 (N_1686,In_19,In_832);
nand U1687 (N_1687,In_745,In_367);
and U1688 (N_1688,In_836,In_680);
or U1689 (N_1689,In_311,In_599);
nor U1690 (N_1690,In_969,In_74);
or U1691 (N_1691,In_431,In_764);
nand U1692 (N_1692,In_144,In_921);
nand U1693 (N_1693,In_883,In_959);
nand U1694 (N_1694,In_239,In_290);
nand U1695 (N_1695,In_289,In_963);
nor U1696 (N_1696,In_375,In_589);
nand U1697 (N_1697,In_255,In_502);
and U1698 (N_1698,In_258,In_464);
nand U1699 (N_1699,In_244,In_748);
and U1700 (N_1700,In_962,In_923);
nand U1701 (N_1701,In_378,In_514);
and U1702 (N_1702,In_608,In_338);
and U1703 (N_1703,In_673,In_18);
and U1704 (N_1704,In_873,In_212);
or U1705 (N_1705,In_895,In_584);
nor U1706 (N_1706,In_737,In_733);
nand U1707 (N_1707,In_925,In_527);
xor U1708 (N_1708,In_335,In_495);
and U1709 (N_1709,In_949,In_301);
nand U1710 (N_1710,In_71,In_502);
nor U1711 (N_1711,In_181,In_442);
nand U1712 (N_1712,In_8,In_921);
nor U1713 (N_1713,In_32,In_209);
nor U1714 (N_1714,In_89,In_416);
nand U1715 (N_1715,In_95,In_64);
nor U1716 (N_1716,In_892,In_264);
nor U1717 (N_1717,In_244,In_985);
nand U1718 (N_1718,In_187,In_328);
nor U1719 (N_1719,In_757,In_186);
and U1720 (N_1720,In_160,In_52);
nand U1721 (N_1721,In_587,In_5);
nor U1722 (N_1722,In_253,In_787);
nor U1723 (N_1723,In_669,In_564);
or U1724 (N_1724,In_787,In_108);
and U1725 (N_1725,In_476,In_315);
nand U1726 (N_1726,In_938,In_314);
and U1727 (N_1727,In_552,In_329);
and U1728 (N_1728,In_25,In_722);
nor U1729 (N_1729,In_211,In_203);
nor U1730 (N_1730,In_902,In_786);
or U1731 (N_1731,In_589,In_523);
nand U1732 (N_1732,In_411,In_270);
or U1733 (N_1733,In_908,In_694);
nand U1734 (N_1734,In_583,In_749);
and U1735 (N_1735,In_849,In_59);
nor U1736 (N_1736,In_795,In_144);
nor U1737 (N_1737,In_671,In_716);
and U1738 (N_1738,In_47,In_942);
or U1739 (N_1739,In_944,In_837);
and U1740 (N_1740,In_478,In_994);
nor U1741 (N_1741,In_217,In_756);
nor U1742 (N_1742,In_541,In_136);
or U1743 (N_1743,In_327,In_772);
xnor U1744 (N_1744,In_82,In_714);
or U1745 (N_1745,In_834,In_527);
or U1746 (N_1746,In_582,In_577);
and U1747 (N_1747,In_473,In_24);
nand U1748 (N_1748,In_300,In_80);
or U1749 (N_1749,In_144,In_328);
nand U1750 (N_1750,In_468,In_519);
or U1751 (N_1751,In_104,In_333);
or U1752 (N_1752,In_21,In_667);
and U1753 (N_1753,In_13,In_350);
or U1754 (N_1754,In_829,In_29);
and U1755 (N_1755,In_541,In_41);
or U1756 (N_1756,In_38,In_985);
or U1757 (N_1757,In_656,In_700);
or U1758 (N_1758,In_700,In_56);
xnor U1759 (N_1759,In_482,In_559);
and U1760 (N_1760,In_747,In_225);
and U1761 (N_1761,In_609,In_828);
xnor U1762 (N_1762,In_312,In_118);
or U1763 (N_1763,In_711,In_740);
nand U1764 (N_1764,In_778,In_255);
and U1765 (N_1765,In_952,In_158);
or U1766 (N_1766,In_335,In_606);
nor U1767 (N_1767,In_412,In_52);
nand U1768 (N_1768,In_611,In_176);
and U1769 (N_1769,In_661,In_462);
nor U1770 (N_1770,In_748,In_219);
xnor U1771 (N_1771,In_183,In_723);
nand U1772 (N_1772,In_762,In_62);
xor U1773 (N_1773,In_557,In_4);
nand U1774 (N_1774,In_408,In_716);
and U1775 (N_1775,In_25,In_367);
or U1776 (N_1776,In_597,In_887);
or U1777 (N_1777,In_669,In_585);
and U1778 (N_1778,In_160,In_500);
or U1779 (N_1779,In_626,In_799);
and U1780 (N_1780,In_577,In_458);
or U1781 (N_1781,In_572,In_492);
nand U1782 (N_1782,In_457,In_246);
xor U1783 (N_1783,In_151,In_77);
or U1784 (N_1784,In_89,In_924);
nand U1785 (N_1785,In_306,In_300);
nand U1786 (N_1786,In_590,In_466);
nand U1787 (N_1787,In_547,In_754);
and U1788 (N_1788,In_9,In_468);
nand U1789 (N_1789,In_115,In_817);
nor U1790 (N_1790,In_617,In_993);
and U1791 (N_1791,In_326,In_256);
nor U1792 (N_1792,In_802,In_85);
nand U1793 (N_1793,In_524,In_760);
or U1794 (N_1794,In_301,In_545);
nand U1795 (N_1795,In_725,In_538);
nor U1796 (N_1796,In_594,In_781);
nor U1797 (N_1797,In_677,In_201);
or U1798 (N_1798,In_892,In_947);
or U1799 (N_1799,In_568,In_246);
or U1800 (N_1800,In_730,In_335);
xnor U1801 (N_1801,In_876,In_402);
nand U1802 (N_1802,In_821,In_356);
or U1803 (N_1803,In_133,In_505);
and U1804 (N_1804,In_628,In_800);
or U1805 (N_1805,In_676,In_859);
nand U1806 (N_1806,In_348,In_44);
nand U1807 (N_1807,In_185,In_165);
and U1808 (N_1808,In_922,In_790);
or U1809 (N_1809,In_924,In_828);
nand U1810 (N_1810,In_574,In_595);
or U1811 (N_1811,In_356,In_85);
nor U1812 (N_1812,In_935,In_806);
nor U1813 (N_1813,In_43,In_161);
or U1814 (N_1814,In_415,In_439);
or U1815 (N_1815,In_901,In_407);
or U1816 (N_1816,In_390,In_366);
and U1817 (N_1817,In_910,In_16);
nand U1818 (N_1818,In_294,In_561);
nor U1819 (N_1819,In_100,In_983);
xnor U1820 (N_1820,In_777,In_525);
nand U1821 (N_1821,In_27,In_420);
nor U1822 (N_1822,In_488,In_585);
nor U1823 (N_1823,In_812,In_149);
and U1824 (N_1824,In_322,In_695);
nand U1825 (N_1825,In_552,In_675);
and U1826 (N_1826,In_123,In_630);
nand U1827 (N_1827,In_988,In_588);
or U1828 (N_1828,In_348,In_956);
nor U1829 (N_1829,In_571,In_154);
and U1830 (N_1830,In_677,In_494);
nor U1831 (N_1831,In_508,In_443);
and U1832 (N_1832,In_23,In_419);
nand U1833 (N_1833,In_204,In_682);
and U1834 (N_1834,In_63,In_763);
nand U1835 (N_1835,In_695,In_680);
and U1836 (N_1836,In_234,In_92);
nand U1837 (N_1837,In_771,In_615);
nand U1838 (N_1838,In_703,In_328);
and U1839 (N_1839,In_24,In_98);
and U1840 (N_1840,In_121,In_178);
or U1841 (N_1841,In_715,In_21);
and U1842 (N_1842,In_766,In_937);
and U1843 (N_1843,In_448,In_387);
or U1844 (N_1844,In_465,In_440);
nand U1845 (N_1845,In_574,In_344);
nor U1846 (N_1846,In_580,In_644);
nand U1847 (N_1847,In_420,In_243);
nor U1848 (N_1848,In_945,In_482);
nor U1849 (N_1849,In_515,In_3);
or U1850 (N_1850,In_112,In_782);
and U1851 (N_1851,In_0,In_851);
or U1852 (N_1852,In_591,In_709);
and U1853 (N_1853,In_152,In_481);
and U1854 (N_1854,In_128,In_73);
or U1855 (N_1855,In_498,In_288);
nand U1856 (N_1856,In_388,In_921);
nor U1857 (N_1857,In_741,In_103);
and U1858 (N_1858,In_834,In_646);
nor U1859 (N_1859,In_805,In_125);
nand U1860 (N_1860,In_63,In_361);
nand U1861 (N_1861,In_887,In_311);
nor U1862 (N_1862,In_513,In_555);
or U1863 (N_1863,In_161,In_718);
or U1864 (N_1864,In_385,In_233);
or U1865 (N_1865,In_181,In_852);
nor U1866 (N_1866,In_4,In_281);
nor U1867 (N_1867,In_245,In_519);
and U1868 (N_1868,In_931,In_238);
nor U1869 (N_1869,In_618,In_290);
nor U1870 (N_1870,In_288,In_557);
and U1871 (N_1871,In_576,In_75);
nand U1872 (N_1872,In_419,In_489);
and U1873 (N_1873,In_802,In_956);
nor U1874 (N_1874,In_93,In_383);
nand U1875 (N_1875,In_678,In_456);
and U1876 (N_1876,In_309,In_334);
or U1877 (N_1877,In_145,In_567);
or U1878 (N_1878,In_652,In_3);
and U1879 (N_1879,In_355,In_71);
or U1880 (N_1880,In_996,In_76);
xor U1881 (N_1881,In_905,In_345);
nor U1882 (N_1882,In_215,In_901);
nand U1883 (N_1883,In_33,In_39);
and U1884 (N_1884,In_652,In_891);
or U1885 (N_1885,In_596,In_104);
or U1886 (N_1886,In_531,In_838);
and U1887 (N_1887,In_1,In_503);
nand U1888 (N_1888,In_916,In_245);
nand U1889 (N_1889,In_97,In_594);
and U1890 (N_1890,In_463,In_426);
nand U1891 (N_1891,In_420,In_858);
nand U1892 (N_1892,In_810,In_401);
or U1893 (N_1893,In_154,In_619);
nand U1894 (N_1894,In_7,In_231);
nand U1895 (N_1895,In_723,In_760);
xor U1896 (N_1896,In_220,In_258);
or U1897 (N_1897,In_807,In_504);
or U1898 (N_1898,In_573,In_99);
xor U1899 (N_1899,In_631,In_931);
xnor U1900 (N_1900,In_660,In_446);
or U1901 (N_1901,In_823,In_126);
or U1902 (N_1902,In_395,In_919);
nor U1903 (N_1903,In_49,In_484);
nor U1904 (N_1904,In_924,In_709);
nor U1905 (N_1905,In_598,In_213);
or U1906 (N_1906,In_828,In_221);
nand U1907 (N_1907,In_971,In_206);
xnor U1908 (N_1908,In_550,In_930);
or U1909 (N_1909,In_690,In_681);
and U1910 (N_1910,In_178,In_914);
and U1911 (N_1911,In_400,In_932);
nor U1912 (N_1912,In_74,In_403);
and U1913 (N_1913,In_521,In_430);
or U1914 (N_1914,In_616,In_853);
nor U1915 (N_1915,In_578,In_260);
nand U1916 (N_1916,In_149,In_803);
nor U1917 (N_1917,In_465,In_943);
and U1918 (N_1918,In_794,In_304);
and U1919 (N_1919,In_20,In_429);
nor U1920 (N_1920,In_109,In_946);
and U1921 (N_1921,In_82,In_286);
nand U1922 (N_1922,In_698,In_115);
or U1923 (N_1923,In_976,In_879);
and U1924 (N_1924,In_995,In_607);
and U1925 (N_1925,In_981,In_182);
or U1926 (N_1926,In_461,In_416);
nor U1927 (N_1927,In_291,In_990);
and U1928 (N_1928,In_316,In_675);
nand U1929 (N_1929,In_672,In_553);
and U1930 (N_1930,In_195,In_316);
nor U1931 (N_1931,In_621,In_938);
and U1932 (N_1932,In_538,In_177);
or U1933 (N_1933,In_142,In_473);
nor U1934 (N_1934,In_891,In_635);
and U1935 (N_1935,In_995,In_846);
and U1936 (N_1936,In_310,In_125);
nand U1937 (N_1937,In_586,In_471);
or U1938 (N_1938,In_452,In_801);
xor U1939 (N_1939,In_399,In_865);
nand U1940 (N_1940,In_741,In_301);
or U1941 (N_1941,In_200,In_399);
nand U1942 (N_1942,In_705,In_982);
or U1943 (N_1943,In_324,In_787);
nor U1944 (N_1944,In_272,In_338);
nor U1945 (N_1945,In_776,In_328);
or U1946 (N_1946,In_514,In_739);
and U1947 (N_1947,In_799,In_154);
nand U1948 (N_1948,In_478,In_870);
and U1949 (N_1949,In_443,In_159);
and U1950 (N_1950,In_461,In_88);
xnor U1951 (N_1951,In_544,In_457);
nand U1952 (N_1952,In_407,In_666);
nor U1953 (N_1953,In_116,In_793);
and U1954 (N_1954,In_695,In_757);
nor U1955 (N_1955,In_111,In_659);
nand U1956 (N_1956,In_115,In_221);
and U1957 (N_1957,In_95,In_635);
nor U1958 (N_1958,In_387,In_18);
nand U1959 (N_1959,In_848,In_957);
xnor U1960 (N_1960,In_845,In_473);
nand U1961 (N_1961,In_433,In_523);
nand U1962 (N_1962,In_924,In_321);
nand U1963 (N_1963,In_440,In_183);
nor U1964 (N_1964,In_197,In_199);
or U1965 (N_1965,In_589,In_609);
and U1966 (N_1966,In_332,In_825);
or U1967 (N_1967,In_447,In_498);
nor U1968 (N_1968,In_500,In_594);
or U1969 (N_1969,In_185,In_741);
nand U1970 (N_1970,In_227,In_173);
or U1971 (N_1971,In_789,In_393);
or U1972 (N_1972,In_384,In_886);
and U1973 (N_1973,In_640,In_759);
nand U1974 (N_1974,In_41,In_294);
or U1975 (N_1975,In_254,In_541);
nand U1976 (N_1976,In_941,In_437);
nor U1977 (N_1977,In_3,In_90);
nor U1978 (N_1978,In_724,In_836);
nand U1979 (N_1979,In_53,In_826);
nor U1980 (N_1980,In_669,In_65);
and U1981 (N_1981,In_931,In_312);
nor U1982 (N_1982,In_44,In_875);
or U1983 (N_1983,In_907,In_454);
or U1984 (N_1984,In_745,In_549);
nor U1985 (N_1985,In_734,In_281);
and U1986 (N_1986,In_464,In_487);
and U1987 (N_1987,In_472,In_97);
and U1988 (N_1988,In_151,In_931);
nand U1989 (N_1989,In_192,In_403);
or U1990 (N_1990,In_612,In_599);
nand U1991 (N_1991,In_274,In_647);
nand U1992 (N_1992,In_448,In_250);
nand U1993 (N_1993,In_600,In_10);
nand U1994 (N_1994,In_496,In_740);
and U1995 (N_1995,In_938,In_446);
nand U1996 (N_1996,In_575,In_294);
nand U1997 (N_1997,In_56,In_886);
nor U1998 (N_1998,In_710,In_562);
or U1999 (N_1999,In_399,In_517);
nand U2000 (N_2000,In_888,In_713);
or U2001 (N_2001,In_983,In_425);
or U2002 (N_2002,In_801,In_19);
or U2003 (N_2003,In_504,In_673);
xor U2004 (N_2004,In_404,In_406);
nor U2005 (N_2005,In_960,In_496);
nand U2006 (N_2006,In_697,In_637);
and U2007 (N_2007,In_67,In_293);
xnor U2008 (N_2008,In_687,In_588);
or U2009 (N_2009,In_444,In_723);
and U2010 (N_2010,In_407,In_860);
and U2011 (N_2011,In_633,In_390);
nor U2012 (N_2012,In_497,In_966);
nand U2013 (N_2013,In_951,In_801);
and U2014 (N_2014,In_481,In_803);
or U2015 (N_2015,In_472,In_888);
nor U2016 (N_2016,In_516,In_358);
and U2017 (N_2017,In_176,In_174);
nand U2018 (N_2018,In_677,In_412);
or U2019 (N_2019,In_752,In_592);
and U2020 (N_2020,In_170,In_898);
or U2021 (N_2021,In_476,In_280);
nand U2022 (N_2022,In_914,In_139);
or U2023 (N_2023,In_569,In_535);
nand U2024 (N_2024,In_182,In_463);
and U2025 (N_2025,In_997,In_509);
nand U2026 (N_2026,In_598,In_91);
and U2027 (N_2027,In_69,In_441);
and U2028 (N_2028,In_589,In_591);
or U2029 (N_2029,In_986,In_346);
nor U2030 (N_2030,In_78,In_725);
or U2031 (N_2031,In_665,In_839);
or U2032 (N_2032,In_489,In_119);
nand U2033 (N_2033,In_495,In_179);
and U2034 (N_2034,In_166,In_114);
or U2035 (N_2035,In_108,In_500);
nor U2036 (N_2036,In_58,In_627);
and U2037 (N_2037,In_44,In_144);
or U2038 (N_2038,In_663,In_358);
nand U2039 (N_2039,In_916,In_342);
and U2040 (N_2040,In_718,In_832);
nor U2041 (N_2041,In_522,In_533);
and U2042 (N_2042,In_238,In_188);
or U2043 (N_2043,In_951,In_231);
xor U2044 (N_2044,In_832,In_566);
and U2045 (N_2045,In_61,In_646);
and U2046 (N_2046,In_236,In_862);
nor U2047 (N_2047,In_924,In_609);
xnor U2048 (N_2048,In_4,In_722);
or U2049 (N_2049,In_991,In_508);
nor U2050 (N_2050,In_983,In_62);
nor U2051 (N_2051,In_947,In_351);
and U2052 (N_2052,In_714,In_122);
nand U2053 (N_2053,In_853,In_127);
xor U2054 (N_2054,In_810,In_494);
nor U2055 (N_2055,In_215,In_809);
and U2056 (N_2056,In_866,In_130);
or U2057 (N_2057,In_980,In_402);
and U2058 (N_2058,In_857,In_424);
or U2059 (N_2059,In_60,In_497);
or U2060 (N_2060,In_348,In_634);
and U2061 (N_2061,In_261,In_339);
nand U2062 (N_2062,In_570,In_813);
nor U2063 (N_2063,In_919,In_858);
and U2064 (N_2064,In_289,In_830);
nor U2065 (N_2065,In_946,In_614);
nor U2066 (N_2066,In_64,In_326);
nor U2067 (N_2067,In_2,In_321);
and U2068 (N_2068,In_304,In_286);
nand U2069 (N_2069,In_608,In_363);
nand U2070 (N_2070,In_796,In_423);
or U2071 (N_2071,In_44,In_451);
nor U2072 (N_2072,In_410,In_584);
nor U2073 (N_2073,In_866,In_11);
and U2074 (N_2074,In_630,In_270);
nand U2075 (N_2075,In_473,In_859);
nor U2076 (N_2076,In_938,In_237);
nand U2077 (N_2077,In_648,In_875);
nand U2078 (N_2078,In_377,In_814);
or U2079 (N_2079,In_976,In_622);
and U2080 (N_2080,In_19,In_446);
nor U2081 (N_2081,In_938,In_603);
nand U2082 (N_2082,In_558,In_519);
or U2083 (N_2083,In_849,In_341);
nor U2084 (N_2084,In_100,In_370);
nand U2085 (N_2085,In_437,In_415);
or U2086 (N_2086,In_563,In_244);
nor U2087 (N_2087,In_376,In_747);
or U2088 (N_2088,In_434,In_100);
and U2089 (N_2089,In_22,In_61);
and U2090 (N_2090,In_400,In_382);
or U2091 (N_2091,In_494,In_834);
or U2092 (N_2092,In_746,In_759);
and U2093 (N_2093,In_822,In_357);
and U2094 (N_2094,In_445,In_772);
or U2095 (N_2095,In_175,In_819);
nand U2096 (N_2096,In_202,In_126);
nand U2097 (N_2097,In_936,In_542);
nand U2098 (N_2098,In_457,In_20);
nand U2099 (N_2099,In_371,In_341);
nand U2100 (N_2100,In_216,In_142);
and U2101 (N_2101,In_200,In_217);
or U2102 (N_2102,In_993,In_559);
nand U2103 (N_2103,In_96,In_197);
or U2104 (N_2104,In_783,In_517);
nand U2105 (N_2105,In_843,In_225);
nor U2106 (N_2106,In_570,In_543);
nor U2107 (N_2107,In_729,In_531);
nand U2108 (N_2108,In_911,In_512);
and U2109 (N_2109,In_738,In_631);
or U2110 (N_2110,In_618,In_112);
nand U2111 (N_2111,In_947,In_99);
nand U2112 (N_2112,In_578,In_993);
nor U2113 (N_2113,In_318,In_18);
or U2114 (N_2114,In_870,In_31);
nor U2115 (N_2115,In_74,In_250);
xnor U2116 (N_2116,In_660,In_749);
nor U2117 (N_2117,In_449,In_302);
nor U2118 (N_2118,In_146,In_899);
xnor U2119 (N_2119,In_694,In_928);
nand U2120 (N_2120,In_943,In_604);
and U2121 (N_2121,In_239,In_939);
and U2122 (N_2122,In_105,In_797);
nor U2123 (N_2123,In_767,In_571);
or U2124 (N_2124,In_101,In_881);
or U2125 (N_2125,In_732,In_976);
and U2126 (N_2126,In_298,In_557);
or U2127 (N_2127,In_869,In_127);
or U2128 (N_2128,In_241,In_100);
or U2129 (N_2129,In_877,In_44);
and U2130 (N_2130,In_756,In_158);
and U2131 (N_2131,In_119,In_743);
or U2132 (N_2132,In_969,In_991);
nand U2133 (N_2133,In_877,In_952);
and U2134 (N_2134,In_469,In_118);
nand U2135 (N_2135,In_671,In_446);
and U2136 (N_2136,In_880,In_376);
or U2137 (N_2137,In_0,In_966);
or U2138 (N_2138,In_331,In_404);
nand U2139 (N_2139,In_278,In_823);
nand U2140 (N_2140,In_960,In_537);
and U2141 (N_2141,In_586,In_351);
and U2142 (N_2142,In_854,In_112);
and U2143 (N_2143,In_515,In_402);
xnor U2144 (N_2144,In_132,In_886);
nor U2145 (N_2145,In_841,In_403);
nand U2146 (N_2146,In_583,In_300);
or U2147 (N_2147,In_942,In_948);
nand U2148 (N_2148,In_422,In_795);
nand U2149 (N_2149,In_160,In_21);
nand U2150 (N_2150,In_488,In_812);
and U2151 (N_2151,In_993,In_202);
nand U2152 (N_2152,In_168,In_297);
nand U2153 (N_2153,In_923,In_474);
or U2154 (N_2154,In_872,In_381);
nor U2155 (N_2155,In_290,In_583);
or U2156 (N_2156,In_285,In_898);
nor U2157 (N_2157,In_964,In_377);
xor U2158 (N_2158,In_456,In_391);
nor U2159 (N_2159,In_855,In_632);
or U2160 (N_2160,In_330,In_869);
nor U2161 (N_2161,In_433,In_336);
and U2162 (N_2162,In_379,In_487);
or U2163 (N_2163,In_987,In_610);
and U2164 (N_2164,In_970,In_40);
or U2165 (N_2165,In_616,In_53);
nor U2166 (N_2166,In_960,In_188);
and U2167 (N_2167,In_921,In_945);
or U2168 (N_2168,In_380,In_297);
or U2169 (N_2169,In_192,In_749);
nand U2170 (N_2170,In_245,In_390);
nand U2171 (N_2171,In_575,In_912);
and U2172 (N_2172,In_625,In_233);
nand U2173 (N_2173,In_934,In_249);
nand U2174 (N_2174,In_198,In_987);
nor U2175 (N_2175,In_848,In_587);
xor U2176 (N_2176,In_272,In_96);
xnor U2177 (N_2177,In_569,In_443);
and U2178 (N_2178,In_377,In_247);
and U2179 (N_2179,In_133,In_170);
nor U2180 (N_2180,In_27,In_938);
nor U2181 (N_2181,In_632,In_880);
nand U2182 (N_2182,In_714,In_945);
nor U2183 (N_2183,In_791,In_457);
or U2184 (N_2184,In_569,In_860);
or U2185 (N_2185,In_425,In_707);
nor U2186 (N_2186,In_798,In_623);
nor U2187 (N_2187,In_486,In_765);
nand U2188 (N_2188,In_30,In_15);
nand U2189 (N_2189,In_37,In_251);
nand U2190 (N_2190,In_563,In_50);
and U2191 (N_2191,In_612,In_45);
and U2192 (N_2192,In_304,In_327);
and U2193 (N_2193,In_237,In_555);
nand U2194 (N_2194,In_589,In_513);
nor U2195 (N_2195,In_30,In_100);
and U2196 (N_2196,In_758,In_178);
nor U2197 (N_2197,In_984,In_816);
nand U2198 (N_2198,In_211,In_840);
nor U2199 (N_2199,In_904,In_149);
nand U2200 (N_2200,In_284,In_494);
nor U2201 (N_2201,In_877,In_671);
or U2202 (N_2202,In_453,In_653);
or U2203 (N_2203,In_294,In_0);
nand U2204 (N_2204,In_642,In_770);
nand U2205 (N_2205,In_934,In_925);
and U2206 (N_2206,In_878,In_12);
nand U2207 (N_2207,In_743,In_48);
xnor U2208 (N_2208,In_808,In_24);
or U2209 (N_2209,In_116,In_430);
nor U2210 (N_2210,In_594,In_132);
and U2211 (N_2211,In_899,In_813);
nor U2212 (N_2212,In_42,In_761);
or U2213 (N_2213,In_490,In_554);
or U2214 (N_2214,In_32,In_994);
nor U2215 (N_2215,In_643,In_631);
nand U2216 (N_2216,In_810,In_563);
nand U2217 (N_2217,In_930,In_449);
nor U2218 (N_2218,In_54,In_249);
nor U2219 (N_2219,In_45,In_519);
nand U2220 (N_2220,In_942,In_378);
or U2221 (N_2221,In_584,In_375);
and U2222 (N_2222,In_120,In_392);
nor U2223 (N_2223,In_209,In_833);
nor U2224 (N_2224,In_871,In_752);
nand U2225 (N_2225,In_703,In_892);
or U2226 (N_2226,In_545,In_521);
or U2227 (N_2227,In_477,In_881);
and U2228 (N_2228,In_908,In_353);
or U2229 (N_2229,In_95,In_127);
nand U2230 (N_2230,In_432,In_999);
or U2231 (N_2231,In_891,In_26);
nand U2232 (N_2232,In_503,In_897);
nor U2233 (N_2233,In_532,In_41);
or U2234 (N_2234,In_653,In_621);
nor U2235 (N_2235,In_885,In_912);
nor U2236 (N_2236,In_633,In_395);
or U2237 (N_2237,In_606,In_867);
nand U2238 (N_2238,In_876,In_397);
xnor U2239 (N_2239,In_915,In_559);
and U2240 (N_2240,In_934,In_281);
nor U2241 (N_2241,In_687,In_927);
or U2242 (N_2242,In_621,In_698);
nor U2243 (N_2243,In_432,In_899);
nor U2244 (N_2244,In_864,In_235);
xor U2245 (N_2245,In_410,In_562);
and U2246 (N_2246,In_20,In_746);
nand U2247 (N_2247,In_542,In_546);
and U2248 (N_2248,In_325,In_447);
and U2249 (N_2249,In_452,In_909);
nor U2250 (N_2250,In_567,In_553);
nand U2251 (N_2251,In_147,In_358);
nand U2252 (N_2252,In_692,In_777);
or U2253 (N_2253,In_111,In_450);
nand U2254 (N_2254,In_247,In_998);
and U2255 (N_2255,In_854,In_166);
and U2256 (N_2256,In_492,In_68);
and U2257 (N_2257,In_943,In_359);
nor U2258 (N_2258,In_301,In_923);
nor U2259 (N_2259,In_836,In_440);
nor U2260 (N_2260,In_286,In_325);
nand U2261 (N_2261,In_673,In_972);
nor U2262 (N_2262,In_991,In_839);
nor U2263 (N_2263,In_626,In_38);
nand U2264 (N_2264,In_444,In_356);
nor U2265 (N_2265,In_685,In_110);
nand U2266 (N_2266,In_29,In_824);
nand U2267 (N_2267,In_961,In_999);
or U2268 (N_2268,In_398,In_257);
nor U2269 (N_2269,In_72,In_564);
or U2270 (N_2270,In_377,In_865);
and U2271 (N_2271,In_336,In_838);
nand U2272 (N_2272,In_722,In_389);
nand U2273 (N_2273,In_841,In_889);
nand U2274 (N_2274,In_596,In_728);
nor U2275 (N_2275,In_71,In_388);
and U2276 (N_2276,In_109,In_208);
or U2277 (N_2277,In_379,In_790);
and U2278 (N_2278,In_124,In_23);
nor U2279 (N_2279,In_662,In_108);
or U2280 (N_2280,In_400,In_706);
or U2281 (N_2281,In_920,In_778);
nor U2282 (N_2282,In_57,In_290);
nand U2283 (N_2283,In_507,In_421);
or U2284 (N_2284,In_491,In_86);
or U2285 (N_2285,In_941,In_794);
nand U2286 (N_2286,In_716,In_796);
nor U2287 (N_2287,In_841,In_717);
nand U2288 (N_2288,In_558,In_249);
and U2289 (N_2289,In_920,In_227);
nand U2290 (N_2290,In_49,In_789);
or U2291 (N_2291,In_822,In_998);
nand U2292 (N_2292,In_614,In_30);
and U2293 (N_2293,In_368,In_336);
or U2294 (N_2294,In_420,In_481);
nor U2295 (N_2295,In_120,In_685);
nand U2296 (N_2296,In_865,In_207);
nor U2297 (N_2297,In_186,In_252);
or U2298 (N_2298,In_870,In_114);
nor U2299 (N_2299,In_761,In_16);
nor U2300 (N_2300,In_12,In_420);
nand U2301 (N_2301,In_150,In_118);
and U2302 (N_2302,In_427,In_162);
and U2303 (N_2303,In_636,In_214);
nor U2304 (N_2304,In_735,In_639);
nand U2305 (N_2305,In_490,In_795);
and U2306 (N_2306,In_718,In_635);
nor U2307 (N_2307,In_445,In_915);
and U2308 (N_2308,In_247,In_821);
nand U2309 (N_2309,In_739,In_650);
nand U2310 (N_2310,In_497,In_492);
or U2311 (N_2311,In_82,In_655);
or U2312 (N_2312,In_667,In_748);
or U2313 (N_2313,In_520,In_601);
nor U2314 (N_2314,In_774,In_122);
or U2315 (N_2315,In_682,In_223);
or U2316 (N_2316,In_661,In_280);
nand U2317 (N_2317,In_108,In_626);
and U2318 (N_2318,In_713,In_372);
or U2319 (N_2319,In_82,In_529);
or U2320 (N_2320,In_201,In_647);
xnor U2321 (N_2321,In_755,In_834);
nand U2322 (N_2322,In_559,In_0);
and U2323 (N_2323,In_142,In_538);
nor U2324 (N_2324,In_79,In_377);
and U2325 (N_2325,In_277,In_89);
nand U2326 (N_2326,In_106,In_353);
nor U2327 (N_2327,In_645,In_434);
nand U2328 (N_2328,In_776,In_221);
or U2329 (N_2329,In_868,In_358);
or U2330 (N_2330,In_37,In_790);
nand U2331 (N_2331,In_972,In_443);
and U2332 (N_2332,In_591,In_987);
nand U2333 (N_2333,In_981,In_728);
nor U2334 (N_2334,In_90,In_91);
nor U2335 (N_2335,In_832,In_455);
or U2336 (N_2336,In_596,In_327);
nand U2337 (N_2337,In_680,In_489);
nor U2338 (N_2338,In_766,In_190);
nand U2339 (N_2339,In_667,In_940);
nor U2340 (N_2340,In_22,In_402);
nand U2341 (N_2341,In_606,In_185);
nand U2342 (N_2342,In_590,In_506);
or U2343 (N_2343,In_445,In_653);
or U2344 (N_2344,In_43,In_811);
and U2345 (N_2345,In_600,In_301);
and U2346 (N_2346,In_610,In_766);
nor U2347 (N_2347,In_984,In_558);
or U2348 (N_2348,In_991,In_435);
nor U2349 (N_2349,In_123,In_342);
or U2350 (N_2350,In_803,In_329);
or U2351 (N_2351,In_238,In_886);
nor U2352 (N_2352,In_39,In_264);
or U2353 (N_2353,In_537,In_0);
nor U2354 (N_2354,In_538,In_0);
and U2355 (N_2355,In_495,In_368);
or U2356 (N_2356,In_751,In_23);
and U2357 (N_2357,In_982,In_515);
and U2358 (N_2358,In_349,In_348);
or U2359 (N_2359,In_691,In_100);
nand U2360 (N_2360,In_746,In_369);
nor U2361 (N_2361,In_714,In_754);
xor U2362 (N_2362,In_542,In_308);
nor U2363 (N_2363,In_604,In_627);
or U2364 (N_2364,In_888,In_601);
or U2365 (N_2365,In_429,In_755);
nand U2366 (N_2366,In_859,In_26);
nor U2367 (N_2367,In_389,In_809);
nand U2368 (N_2368,In_258,In_430);
or U2369 (N_2369,In_849,In_666);
or U2370 (N_2370,In_264,In_148);
or U2371 (N_2371,In_928,In_489);
nand U2372 (N_2372,In_22,In_584);
or U2373 (N_2373,In_243,In_887);
and U2374 (N_2374,In_902,In_14);
nand U2375 (N_2375,In_952,In_975);
nor U2376 (N_2376,In_441,In_889);
nor U2377 (N_2377,In_632,In_825);
nor U2378 (N_2378,In_293,In_319);
and U2379 (N_2379,In_498,In_905);
nand U2380 (N_2380,In_958,In_503);
nor U2381 (N_2381,In_1,In_990);
or U2382 (N_2382,In_490,In_144);
and U2383 (N_2383,In_409,In_655);
nor U2384 (N_2384,In_609,In_74);
and U2385 (N_2385,In_339,In_245);
or U2386 (N_2386,In_350,In_524);
nand U2387 (N_2387,In_82,In_980);
and U2388 (N_2388,In_556,In_967);
xor U2389 (N_2389,In_111,In_109);
nor U2390 (N_2390,In_455,In_121);
and U2391 (N_2391,In_65,In_606);
nand U2392 (N_2392,In_441,In_124);
or U2393 (N_2393,In_932,In_235);
nor U2394 (N_2394,In_366,In_707);
nor U2395 (N_2395,In_478,In_522);
nor U2396 (N_2396,In_750,In_403);
or U2397 (N_2397,In_829,In_527);
nor U2398 (N_2398,In_239,In_375);
nand U2399 (N_2399,In_945,In_2);
nand U2400 (N_2400,In_978,In_901);
or U2401 (N_2401,In_565,In_340);
nor U2402 (N_2402,In_851,In_688);
or U2403 (N_2403,In_724,In_885);
and U2404 (N_2404,In_584,In_300);
or U2405 (N_2405,In_131,In_728);
nor U2406 (N_2406,In_781,In_69);
and U2407 (N_2407,In_26,In_744);
nand U2408 (N_2408,In_619,In_360);
nor U2409 (N_2409,In_810,In_209);
nor U2410 (N_2410,In_282,In_36);
nand U2411 (N_2411,In_419,In_421);
and U2412 (N_2412,In_34,In_612);
nor U2413 (N_2413,In_485,In_493);
or U2414 (N_2414,In_247,In_995);
or U2415 (N_2415,In_841,In_208);
nand U2416 (N_2416,In_441,In_738);
nand U2417 (N_2417,In_965,In_557);
nand U2418 (N_2418,In_580,In_216);
nand U2419 (N_2419,In_89,In_792);
or U2420 (N_2420,In_359,In_720);
and U2421 (N_2421,In_611,In_900);
nor U2422 (N_2422,In_383,In_638);
and U2423 (N_2423,In_222,In_82);
or U2424 (N_2424,In_991,In_729);
or U2425 (N_2425,In_704,In_392);
and U2426 (N_2426,In_907,In_58);
nor U2427 (N_2427,In_204,In_786);
and U2428 (N_2428,In_379,In_207);
nand U2429 (N_2429,In_65,In_917);
or U2430 (N_2430,In_509,In_891);
and U2431 (N_2431,In_685,In_627);
nor U2432 (N_2432,In_385,In_927);
and U2433 (N_2433,In_59,In_709);
or U2434 (N_2434,In_610,In_971);
nor U2435 (N_2435,In_548,In_909);
nor U2436 (N_2436,In_119,In_194);
or U2437 (N_2437,In_893,In_693);
or U2438 (N_2438,In_359,In_667);
or U2439 (N_2439,In_349,In_97);
nand U2440 (N_2440,In_805,In_885);
nor U2441 (N_2441,In_131,In_315);
nand U2442 (N_2442,In_522,In_196);
nor U2443 (N_2443,In_290,In_543);
nand U2444 (N_2444,In_981,In_807);
nand U2445 (N_2445,In_908,In_245);
and U2446 (N_2446,In_236,In_987);
nand U2447 (N_2447,In_886,In_374);
xnor U2448 (N_2448,In_656,In_853);
nor U2449 (N_2449,In_885,In_624);
and U2450 (N_2450,In_365,In_302);
and U2451 (N_2451,In_128,In_962);
nor U2452 (N_2452,In_294,In_584);
nand U2453 (N_2453,In_372,In_546);
and U2454 (N_2454,In_897,In_184);
or U2455 (N_2455,In_546,In_213);
nand U2456 (N_2456,In_279,In_832);
or U2457 (N_2457,In_991,In_773);
nand U2458 (N_2458,In_478,In_334);
nand U2459 (N_2459,In_521,In_648);
xnor U2460 (N_2460,In_504,In_372);
nor U2461 (N_2461,In_6,In_786);
nand U2462 (N_2462,In_44,In_353);
and U2463 (N_2463,In_254,In_365);
nor U2464 (N_2464,In_760,In_165);
nand U2465 (N_2465,In_734,In_866);
nor U2466 (N_2466,In_494,In_860);
or U2467 (N_2467,In_214,In_311);
or U2468 (N_2468,In_306,In_481);
and U2469 (N_2469,In_611,In_747);
or U2470 (N_2470,In_504,In_749);
and U2471 (N_2471,In_326,In_485);
and U2472 (N_2472,In_517,In_665);
nor U2473 (N_2473,In_706,In_598);
nor U2474 (N_2474,In_26,In_133);
or U2475 (N_2475,In_24,In_63);
and U2476 (N_2476,In_726,In_674);
nand U2477 (N_2477,In_911,In_1);
nor U2478 (N_2478,In_350,In_434);
nand U2479 (N_2479,In_888,In_415);
nor U2480 (N_2480,In_977,In_158);
nor U2481 (N_2481,In_35,In_440);
nor U2482 (N_2482,In_605,In_506);
and U2483 (N_2483,In_526,In_26);
and U2484 (N_2484,In_122,In_442);
and U2485 (N_2485,In_377,In_215);
nor U2486 (N_2486,In_564,In_756);
nor U2487 (N_2487,In_122,In_396);
or U2488 (N_2488,In_374,In_426);
nor U2489 (N_2489,In_448,In_583);
or U2490 (N_2490,In_684,In_930);
and U2491 (N_2491,In_938,In_574);
and U2492 (N_2492,In_346,In_379);
nand U2493 (N_2493,In_938,In_211);
nor U2494 (N_2494,In_358,In_508);
and U2495 (N_2495,In_147,In_464);
and U2496 (N_2496,In_737,In_30);
or U2497 (N_2497,In_758,In_745);
nand U2498 (N_2498,In_999,In_192);
and U2499 (N_2499,In_829,In_711);
and U2500 (N_2500,In_725,In_379);
xnor U2501 (N_2501,In_285,In_831);
nor U2502 (N_2502,In_735,In_116);
or U2503 (N_2503,In_912,In_938);
or U2504 (N_2504,In_878,In_290);
nand U2505 (N_2505,In_71,In_106);
nor U2506 (N_2506,In_203,In_836);
nor U2507 (N_2507,In_61,In_23);
and U2508 (N_2508,In_665,In_279);
nand U2509 (N_2509,In_229,In_77);
nor U2510 (N_2510,In_212,In_728);
nor U2511 (N_2511,In_851,In_411);
or U2512 (N_2512,In_466,In_154);
nor U2513 (N_2513,In_616,In_525);
or U2514 (N_2514,In_440,In_278);
nand U2515 (N_2515,In_634,In_148);
nand U2516 (N_2516,In_870,In_39);
or U2517 (N_2517,In_436,In_399);
and U2518 (N_2518,In_557,In_499);
nand U2519 (N_2519,In_236,In_275);
nor U2520 (N_2520,In_330,In_930);
and U2521 (N_2521,In_447,In_703);
or U2522 (N_2522,In_894,In_534);
nand U2523 (N_2523,In_357,In_248);
nand U2524 (N_2524,In_154,In_976);
or U2525 (N_2525,In_734,In_372);
and U2526 (N_2526,In_632,In_334);
and U2527 (N_2527,In_715,In_4);
nand U2528 (N_2528,In_3,In_291);
and U2529 (N_2529,In_140,In_186);
and U2530 (N_2530,In_939,In_680);
or U2531 (N_2531,In_504,In_984);
and U2532 (N_2532,In_974,In_790);
nor U2533 (N_2533,In_956,In_684);
nor U2534 (N_2534,In_745,In_739);
or U2535 (N_2535,In_693,In_398);
and U2536 (N_2536,In_33,In_222);
nand U2537 (N_2537,In_206,In_651);
or U2538 (N_2538,In_283,In_933);
nand U2539 (N_2539,In_337,In_960);
or U2540 (N_2540,In_373,In_453);
nand U2541 (N_2541,In_73,In_985);
and U2542 (N_2542,In_792,In_825);
or U2543 (N_2543,In_91,In_662);
nand U2544 (N_2544,In_407,In_795);
nor U2545 (N_2545,In_351,In_384);
nor U2546 (N_2546,In_256,In_366);
nor U2547 (N_2547,In_427,In_444);
nor U2548 (N_2548,In_988,In_407);
nand U2549 (N_2549,In_547,In_916);
nor U2550 (N_2550,In_822,In_162);
and U2551 (N_2551,In_830,In_566);
and U2552 (N_2552,In_722,In_250);
nand U2553 (N_2553,In_793,In_704);
or U2554 (N_2554,In_962,In_116);
or U2555 (N_2555,In_170,In_278);
nor U2556 (N_2556,In_984,In_823);
and U2557 (N_2557,In_877,In_610);
nor U2558 (N_2558,In_981,In_833);
and U2559 (N_2559,In_356,In_43);
and U2560 (N_2560,In_312,In_169);
nand U2561 (N_2561,In_961,In_659);
nand U2562 (N_2562,In_331,In_691);
or U2563 (N_2563,In_531,In_250);
or U2564 (N_2564,In_929,In_146);
or U2565 (N_2565,In_571,In_0);
and U2566 (N_2566,In_412,In_573);
or U2567 (N_2567,In_883,In_372);
nand U2568 (N_2568,In_203,In_62);
nor U2569 (N_2569,In_193,In_775);
nand U2570 (N_2570,In_804,In_388);
nor U2571 (N_2571,In_591,In_12);
nand U2572 (N_2572,In_263,In_693);
and U2573 (N_2573,In_302,In_316);
or U2574 (N_2574,In_567,In_835);
nor U2575 (N_2575,In_624,In_58);
or U2576 (N_2576,In_758,In_674);
nor U2577 (N_2577,In_631,In_891);
and U2578 (N_2578,In_446,In_691);
nand U2579 (N_2579,In_268,In_207);
nor U2580 (N_2580,In_593,In_289);
and U2581 (N_2581,In_531,In_999);
and U2582 (N_2582,In_205,In_136);
nand U2583 (N_2583,In_336,In_114);
or U2584 (N_2584,In_568,In_396);
nor U2585 (N_2585,In_601,In_75);
nand U2586 (N_2586,In_856,In_438);
or U2587 (N_2587,In_881,In_535);
or U2588 (N_2588,In_908,In_764);
and U2589 (N_2589,In_420,In_400);
nor U2590 (N_2590,In_722,In_540);
nor U2591 (N_2591,In_259,In_884);
or U2592 (N_2592,In_126,In_183);
or U2593 (N_2593,In_962,In_594);
or U2594 (N_2594,In_458,In_403);
and U2595 (N_2595,In_96,In_373);
nor U2596 (N_2596,In_937,In_483);
nand U2597 (N_2597,In_463,In_882);
and U2598 (N_2598,In_400,In_512);
nand U2599 (N_2599,In_940,In_588);
and U2600 (N_2600,In_952,In_470);
and U2601 (N_2601,In_712,In_981);
nor U2602 (N_2602,In_962,In_549);
and U2603 (N_2603,In_900,In_864);
nand U2604 (N_2604,In_100,In_430);
nand U2605 (N_2605,In_193,In_894);
nor U2606 (N_2606,In_24,In_555);
nor U2607 (N_2607,In_509,In_387);
nand U2608 (N_2608,In_300,In_384);
and U2609 (N_2609,In_241,In_291);
nor U2610 (N_2610,In_808,In_695);
nand U2611 (N_2611,In_361,In_298);
or U2612 (N_2612,In_911,In_672);
nor U2613 (N_2613,In_248,In_49);
and U2614 (N_2614,In_977,In_869);
nor U2615 (N_2615,In_683,In_878);
xor U2616 (N_2616,In_777,In_232);
nor U2617 (N_2617,In_346,In_228);
nor U2618 (N_2618,In_973,In_679);
or U2619 (N_2619,In_337,In_826);
nor U2620 (N_2620,In_87,In_32);
and U2621 (N_2621,In_751,In_282);
nand U2622 (N_2622,In_403,In_836);
nand U2623 (N_2623,In_184,In_157);
or U2624 (N_2624,In_141,In_335);
and U2625 (N_2625,In_615,In_796);
nand U2626 (N_2626,In_39,In_863);
nor U2627 (N_2627,In_569,In_349);
nand U2628 (N_2628,In_223,In_167);
nor U2629 (N_2629,In_75,In_228);
or U2630 (N_2630,In_658,In_265);
nor U2631 (N_2631,In_558,In_218);
nor U2632 (N_2632,In_653,In_23);
nor U2633 (N_2633,In_575,In_931);
or U2634 (N_2634,In_725,In_172);
nand U2635 (N_2635,In_274,In_47);
nand U2636 (N_2636,In_589,In_308);
and U2637 (N_2637,In_652,In_726);
nand U2638 (N_2638,In_657,In_232);
nor U2639 (N_2639,In_783,In_835);
and U2640 (N_2640,In_330,In_803);
or U2641 (N_2641,In_805,In_407);
and U2642 (N_2642,In_872,In_674);
nand U2643 (N_2643,In_288,In_596);
or U2644 (N_2644,In_746,In_871);
xnor U2645 (N_2645,In_586,In_253);
nor U2646 (N_2646,In_847,In_212);
and U2647 (N_2647,In_813,In_994);
nand U2648 (N_2648,In_229,In_329);
or U2649 (N_2649,In_410,In_921);
and U2650 (N_2650,In_497,In_904);
or U2651 (N_2651,In_348,In_477);
or U2652 (N_2652,In_584,In_874);
or U2653 (N_2653,In_610,In_861);
nand U2654 (N_2654,In_683,In_769);
and U2655 (N_2655,In_362,In_176);
nor U2656 (N_2656,In_139,In_279);
or U2657 (N_2657,In_252,In_760);
nor U2658 (N_2658,In_582,In_868);
and U2659 (N_2659,In_547,In_691);
nand U2660 (N_2660,In_699,In_807);
nor U2661 (N_2661,In_549,In_983);
and U2662 (N_2662,In_990,In_691);
nor U2663 (N_2663,In_454,In_144);
xor U2664 (N_2664,In_573,In_79);
and U2665 (N_2665,In_617,In_802);
and U2666 (N_2666,In_531,In_852);
and U2667 (N_2667,In_36,In_365);
and U2668 (N_2668,In_301,In_139);
nand U2669 (N_2669,In_68,In_339);
or U2670 (N_2670,In_123,In_90);
nor U2671 (N_2671,In_190,In_156);
nor U2672 (N_2672,In_271,In_430);
nand U2673 (N_2673,In_169,In_496);
and U2674 (N_2674,In_336,In_612);
and U2675 (N_2675,In_348,In_902);
nor U2676 (N_2676,In_38,In_69);
and U2677 (N_2677,In_400,In_540);
nand U2678 (N_2678,In_274,In_239);
nand U2679 (N_2679,In_183,In_627);
or U2680 (N_2680,In_221,In_640);
nand U2681 (N_2681,In_260,In_143);
nand U2682 (N_2682,In_203,In_498);
and U2683 (N_2683,In_514,In_553);
and U2684 (N_2684,In_315,In_781);
nand U2685 (N_2685,In_484,In_727);
and U2686 (N_2686,In_559,In_653);
or U2687 (N_2687,In_541,In_659);
nor U2688 (N_2688,In_416,In_936);
nand U2689 (N_2689,In_713,In_60);
or U2690 (N_2690,In_999,In_45);
and U2691 (N_2691,In_862,In_267);
xnor U2692 (N_2692,In_135,In_71);
nor U2693 (N_2693,In_228,In_696);
nor U2694 (N_2694,In_871,In_621);
and U2695 (N_2695,In_285,In_559);
nor U2696 (N_2696,In_150,In_881);
or U2697 (N_2697,In_48,In_760);
and U2698 (N_2698,In_303,In_961);
or U2699 (N_2699,In_27,In_285);
and U2700 (N_2700,In_586,In_792);
nor U2701 (N_2701,In_486,In_188);
or U2702 (N_2702,In_295,In_628);
and U2703 (N_2703,In_2,In_474);
or U2704 (N_2704,In_841,In_730);
nand U2705 (N_2705,In_460,In_702);
nand U2706 (N_2706,In_614,In_414);
or U2707 (N_2707,In_280,In_909);
or U2708 (N_2708,In_557,In_729);
or U2709 (N_2709,In_158,In_520);
and U2710 (N_2710,In_919,In_964);
nor U2711 (N_2711,In_950,In_67);
or U2712 (N_2712,In_69,In_124);
or U2713 (N_2713,In_340,In_521);
nor U2714 (N_2714,In_495,In_199);
or U2715 (N_2715,In_57,In_680);
and U2716 (N_2716,In_197,In_761);
and U2717 (N_2717,In_845,In_774);
nor U2718 (N_2718,In_947,In_151);
or U2719 (N_2719,In_479,In_965);
or U2720 (N_2720,In_444,In_231);
or U2721 (N_2721,In_207,In_322);
nand U2722 (N_2722,In_507,In_700);
or U2723 (N_2723,In_902,In_798);
or U2724 (N_2724,In_697,In_147);
or U2725 (N_2725,In_49,In_953);
and U2726 (N_2726,In_858,In_758);
and U2727 (N_2727,In_269,In_360);
and U2728 (N_2728,In_541,In_228);
nor U2729 (N_2729,In_784,In_73);
and U2730 (N_2730,In_370,In_179);
nor U2731 (N_2731,In_795,In_227);
or U2732 (N_2732,In_502,In_819);
nand U2733 (N_2733,In_451,In_67);
nor U2734 (N_2734,In_292,In_900);
or U2735 (N_2735,In_167,In_668);
nor U2736 (N_2736,In_709,In_101);
or U2737 (N_2737,In_239,In_588);
nor U2738 (N_2738,In_682,In_392);
and U2739 (N_2739,In_449,In_340);
nor U2740 (N_2740,In_862,In_369);
nor U2741 (N_2741,In_887,In_501);
and U2742 (N_2742,In_127,In_576);
and U2743 (N_2743,In_769,In_236);
nor U2744 (N_2744,In_652,In_475);
nand U2745 (N_2745,In_851,In_161);
nor U2746 (N_2746,In_960,In_773);
and U2747 (N_2747,In_134,In_826);
nand U2748 (N_2748,In_165,In_480);
and U2749 (N_2749,In_238,In_667);
nand U2750 (N_2750,In_926,In_46);
nor U2751 (N_2751,In_140,In_543);
or U2752 (N_2752,In_566,In_320);
xnor U2753 (N_2753,In_855,In_826);
nor U2754 (N_2754,In_220,In_341);
or U2755 (N_2755,In_395,In_307);
or U2756 (N_2756,In_838,In_274);
nor U2757 (N_2757,In_284,In_604);
nor U2758 (N_2758,In_884,In_798);
and U2759 (N_2759,In_320,In_34);
or U2760 (N_2760,In_906,In_109);
nor U2761 (N_2761,In_152,In_251);
nand U2762 (N_2762,In_842,In_541);
nor U2763 (N_2763,In_689,In_654);
or U2764 (N_2764,In_437,In_269);
nand U2765 (N_2765,In_856,In_304);
nor U2766 (N_2766,In_349,In_928);
xnor U2767 (N_2767,In_36,In_41);
nor U2768 (N_2768,In_823,In_359);
or U2769 (N_2769,In_134,In_932);
and U2770 (N_2770,In_950,In_43);
or U2771 (N_2771,In_649,In_880);
nor U2772 (N_2772,In_583,In_946);
and U2773 (N_2773,In_854,In_870);
or U2774 (N_2774,In_692,In_889);
nor U2775 (N_2775,In_827,In_534);
nand U2776 (N_2776,In_953,In_920);
nor U2777 (N_2777,In_415,In_116);
xor U2778 (N_2778,In_594,In_867);
and U2779 (N_2779,In_767,In_903);
and U2780 (N_2780,In_90,In_959);
nor U2781 (N_2781,In_234,In_614);
or U2782 (N_2782,In_745,In_679);
and U2783 (N_2783,In_407,In_728);
nor U2784 (N_2784,In_674,In_518);
or U2785 (N_2785,In_331,In_307);
or U2786 (N_2786,In_210,In_302);
nand U2787 (N_2787,In_775,In_774);
or U2788 (N_2788,In_796,In_536);
nor U2789 (N_2789,In_505,In_684);
nand U2790 (N_2790,In_496,In_980);
or U2791 (N_2791,In_343,In_745);
or U2792 (N_2792,In_642,In_400);
nand U2793 (N_2793,In_328,In_395);
and U2794 (N_2794,In_865,In_880);
and U2795 (N_2795,In_735,In_570);
or U2796 (N_2796,In_410,In_927);
nor U2797 (N_2797,In_807,In_889);
or U2798 (N_2798,In_59,In_453);
nor U2799 (N_2799,In_467,In_885);
and U2800 (N_2800,In_822,In_770);
nand U2801 (N_2801,In_141,In_869);
or U2802 (N_2802,In_606,In_214);
and U2803 (N_2803,In_44,In_558);
nor U2804 (N_2804,In_19,In_234);
nand U2805 (N_2805,In_969,In_355);
nor U2806 (N_2806,In_266,In_444);
and U2807 (N_2807,In_679,In_165);
or U2808 (N_2808,In_684,In_356);
or U2809 (N_2809,In_815,In_111);
nor U2810 (N_2810,In_307,In_979);
nor U2811 (N_2811,In_38,In_660);
or U2812 (N_2812,In_880,In_740);
and U2813 (N_2813,In_354,In_97);
nand U2814 (N_2814,In_505,In_492);
nand U2815 (N_2815,In_867,In_157);
nand U2816 (N_2816,In_231,In_620);
or U2817 (N_2817,In_467,In_296);
nor U2818 (N_2818,In_652,In_246);
or U2819 (N_2819,In_458,In_926);
nor U2820 (N_2820,In_11,In_843);
nor U2821 (N_2821,In_845,In_430);
and U2822 (N_2822,In_78,In_450);
or U2823 (N_2823,In_698,In_827);
or U2824 (N_2824,In_452,In_3);
and U2825 (N_2825,In_1,In_554);
or U2826 (N_2826,In_549,In_919);
nand U2827 (N_2827,In_445,In_988);
nor U2828 (N_2828,In_576,In_387);
and U2829 (N_2829,In_961,In_563);
nor U2830 (N_2830,In_744,In_164);
nand U2831 (N_2831,In_958,In_110);
nor U2832 (N_2832,In_887,In_44);
and U2833 (N_2833,In_880,In_566);
and U2834 (N_2834,In_128,In_728);
and U2835 (N_2835,In_357,In_602);
nand U2836 (N_2836,In_429,In_213);
and U2837 (N_2837,In_660,In_861);
and U2838 (N_2838,In_440,In_26);
and U2839 (N_2839,In_225,In_416);
or U2840 (N_2840,In_404,In_164);
and U2841 (N_2841,In_363,In_956);
nor U2842 (N_2842,In_875,In_461);
or U2843 (N_2843,In_885,In_768);
and U2844 (N_2844,In_428,In_41);
nor U2845 (N_2845,In_917,In_143);
or U2846 (N_2846,In_308,In_187);
nand U2847 (N_2847,In_147,In_875);
or U2848 (N_2848,In_350,In_501);
and U2849 (N_2849,In_187,In_117);
and U2850 (N_2850,In_380,In_923);
nor U2851 (N_2851,In_772,In_289);
nand U2852 (N_2852,In_163,In_573);
nand U2853 (N_2853,In_959,In_431);
nor U2854 (N_2854,In_33,In_827);
and U2855 (N_2855,In_716,In_566);
or U2856 (N_2856,In_342,In_524);
nand U2857 (N_2857,In_439,In_589);
or U2858 (N_2858,In_923,In_855);
or U2859 (N_2859,In_545,In_990);
nand U2860 (N_2860,In_546,In_52);
nor U2861 (N_2861,In_925,In_322);
nand U2862 (N_2862,In_859,In_517);
or U2863 (N_2863,In_157,In_623);
nor U2864 (N_2864,In_585,In_27);
nand U2865 (N_2865,In_480,In_35);
nand U2866 (N_2866,In_308,In_304);
nand U2867 (N_2867,In_260,In_33);
nor U2868 (N_2868,In_131,In_938);
and U2869 (N_2869,In_945,In_84);
or U2870 (N_2870,In_782,In_723);
nand U2871 (N_2871,In_491,In_268);
nand U2872 (N_2872,In_319,In_514);
nor U2873 (N_2873,In_419,In_759);
or U2874 (N_2874,In_940,In_500);
nor U2875 (N_2875,In_598,In_22);
and U2876 (N_2876,In_766,In_640);
and U2877 (N_2877,In_612,In_619);
nor U2878 (N_2878,In_399,In_246);
and U2879 (N_2879,In_158,In_750);
and U2880 (N_2880,In_365,In_510);
or U2881 (N_2881,In_705,In_452);
nor U2882 (N_2882,In_328,In_607);
and U2883 (N_2883,In_772,In_6);
nor U2884 (N_2884,In_651,In_668);
or U2885 (N_2885,In_570,In_659);
and U2886 (N_2886,In_504,In_876);
or U2887 (N_2887,In_478,In_859);
nand U2888 (N_2888,In_782,In_500);
or U2889 (N_2889,In_953,In_776);
or U2890 (N_2890,In_410,In_762);
and U2891 (N_2891,In_101,In_626);
or U2892 (N_2892,In_436,In_619);
and U2893 (N_2893,In_605,In_453);
and U2894 (N_2894,In_688,In_980);
or U2895 (N_2895,In_551,In_216);
nand U2896 (N_2896,In_753,In_935);
or U2897 (N_2897,In_607,In_605);
nand U2898 (N_2898,In_504,In_897);
and U2899 (N_2899,In_863,In_467);
nand U2900 (N_2900,In_944,In_301);
or U2901 (N_2901,In_213,In_292);
or U2902 (N_2902,In_969,In_164);
nand U2903 (N_2903,In_560,In_383);
and U2904 (N_2904,In_722,In_534);
nor U2905 (N_2905,In_666,In_936);
or U2906 (N_2906,In_606,In_379);
nor U2907 (N_2907,In_57,In_331);
nor U2908 (N_2908,In_981,In_759);
or U2909 (N_2909,In_579,In_206);
or U2910 (N_2910,In_344,In_27);
nor U2911 (N_2911,In_236,In_651);
nor U2912 (N_2912,In_54,In_958);
nand U2913 (N_2913,In_468,In_369);
or U2914 (N_2914,In_961,In_985);
or U2915 (N_2915,In_331,In_213);
nand U2916 (N_2916,In_207,In_70);
nand U2917 (N_2917,In_164,In_413);
and U2918 (N_2918,In_985,In_789);
or U2919 (N_2919,In_674,In_680);
or U2920 (N_2920,In_88,In_891);
and U2921 (N_2921,In_699,In_969);
nor U2922 (N_2922,In_981,In_314);
nor U2923 (N_2923,In_364,In_109);
and U2924 (N_2924,In_847,In_557);
nor U2925 (N_2925,In_458,In_234);
nand U2926 (N_2926,In_104,In_103);
and U2927 (N_2927,In_877,In_113);
or U2928 (N_2928,In_387,In_875);
or U2929 (N_2929,In_822,In_24);
nor U2930 (N_2930,In_549,In_856);
nand U2931 (N_2931,In_22,In_396);
xor U2932 (N_2932,In_515,In_962);
nor U2933 (N_2933,In_647,In_308);
or U2934 (N_2934,In_626,In_742);
or U2935 (N_2935,In_449,In_96);
and U2936 (N_2936,In_195,In_581);
or U2937 (N_2937,In_816,In_652);
nor U2938 (N_2938,In_551,In_379);
nand U2939 (N_2939,In_785,In_768);
nor U2940 (N_2940,In_766,In_418);
or U2941 (N_2941,In_305,In_911);
or U2942 (N_2942,In_3,In_746);
nand U2943 (N_2943,In_51,In_296);
nor U2944 (N_2944,In_730,In_913);
and U2945 (N_2945,In_80,In_78);
nand U2946 (N_2946,In_39,In_834);
and U2947 (N_2947,In_662,In_561);
nor U2948 (N_2948,In_940,In_430);
nor U2949 (N_2949,In_387,In_751);
and U2950 (N_2950,In_954,In_674);
nand U2951 (N_2951,In_287,In_617);
and U2952 (N_2952,In_219,In_926);
nor U2953 (N_2953,In_949,In_103);
nand U2954 (N_2954,In_56,In_497);
nor U2955 (N_2955,In_143,In_794);
nor U2956 (N_2956,In_940,In_980);
or U2957 (N_2957,In_96,In_848);
nand U2958 (N_2958,In_529,In_338);
or U2959 (N_2959,In_183,In_168);
nand U2960 (N_2960,In_611,In_23);
nor U2961 (N_2961,In_877,In_178);
nor U2962 (N_2962,In_284,In_439);
nor U2963 (N_2963,In_728,In_16);
nor U2964 (N_2964,In_447,In_788);
and U2965 (N_2965,In_25,In_352);
nor U2966 (N_2966,In_158,In_206);
or U2967 (N_2967,In_531,In_920);
nor U2968 (N_2968,In_90,In_162);
or U2969 (N_2969,In_760,In_228);
and U2970 (N_2970,In_338,In_206);
nor U2971 (N_2971,In_281,In_803);
nand U2972 (N_2972,In_949,In_131);
or U2973 (N_2973,In_711,In_800);
nand U2974 (N_2974,In_376,In_101);
and U2975 (N_2975,In_89,In_368);
nor U2976 (N_2976,In_577,In_802);
or U2977 (N_2977,In_480,In_32);
nand U2978 (N_2978,In_677,In_233);
and U2979 (N_2979,In_55,In_669);
nand U2980 (N_2980,In_363,In_39);
and U2981 (N_2981,In_98,In_628);
xor U2982 (N_2982,In_7,In_841);
nand U2983 (N_2983,In_613,In_774);
nor U2984 (N_2984,In_527,In_746);
nor U2985 (N_2985,In_150,In_756);
or U2986 (N_2986,In_301,In_585);
nor U2987 (N_2987,In_555,In_772);
and U2988 (N_2988,In_22,In_155);
and U2989 (N_2989,In_0,In_308);
nand U2990 (N_2990,In_572,In_406);
or U2991 (N_2991,In_76,In_124);
nand U2992 (N_2992,In_219,In_32);
and U2993 (N_2993,In_45,In_677);
nor U2994 (N_2994,In_413,In_475);
or U2995 (N_2995,In_485,In_59);
and U2996 (N_2996,In_702,In_67);
or U2997 (N_2997,In_44,In_91);
nor U2998 (N_2998,In_375,In_529);
nand U2999 (N_2999,In_208,In_745);
or U3000 (N_3000,In_124,In_960);
or U3001 (N_3001,In_507,In_630);
and U3002 (N_3002,In_250,In_204);
nand U3003 (N_3003,In_805,In_253);
and U3004 (N_3004,In_950,In_560);
nor U3005 (N_3005,In_704,In_466);
nor U3006 (N_3006,In_160,In_841);
nor U3007 (N_3007,In_336,In_989);
nand U3008 (N_3008,In_73,In_40);
or U3009 (N_3009,In_145,In_233);
or U3010 (N_3010,In_59,In_822);
and U3011 (N_3011,In_770,In_638);
nand U3012 (N_3012,In_820,In_399);
nor U3013 (N_3013,In_151,In_897);
nand U3014 (N_3014,In_365,In_134);
nor U3015 (N_3015,In_861,In_669);
nand U3016 (N_3016,In_842,In_779);
nand U3017 (N_3017,In_31,In_122);
nand U3018 (N_3018,In_504,In_612);
or U3019 (N_3019,In_8,In_629);
nand U3020 (N_3020,In_553,In_749);
and U3021 (N_3021,In_651,In_127);
nor U3022 (N_3022,In_867,In_851);
nor U3023 (N_3023,In_12,In_392);
nor U3024 (N_3024,In_394,In_252);
nor U3025 (N_3025,In_9,In_551);
nand U3026 (N_3026,In_652,In_486);
and U3027 (N_3027,In_89,In_357);
nand U3028 (N_3028,In_505,In_314);
nor U3029 (N_3029,In_745,In_507);
or U3030 (N_3030,In_710,In_674);
nand U3031 (N_3031,In_332,In_57);
nand U3032 (N_3032,In_829,In_525);
and U3033 (N_3033,In_345,In_600);
or U3034 (N_3034,In_837,In_159);
and U3035 (N_3035,In_505,In_738);
nand U3036 (N_3036,In_116,In_624);
and U3037 (N_3037,In_151,In_915);
or U3038 (N_3038,In_92,In_989);
nand U3039 (N_3039,In_535,In_537);
or U3040 (N_3040,In_313,In_907);
and U3041 (N_3041,In_165,In_896);
nor U3042 (N_3042,In_400,In_90);
nor U3043 (N_3043,In_556,In_158);
nor U3044 (N_3044,In_14,In_591);
nor U3045 (N_3045,In_220,In_246);
nor U3046 (N_3046,In_247,In_381);
nand U3047 (N_3047,In_997,In_79);
nor U3048 (N_3048,In_563,In_213);
and U3049 (N_3049,In_477,In_833);
nand U3050 (N_3050,In_883,In_977);
nor U3051 (N_3051,In_552,In_524);
xor U3052 (N_3052,In_543,In_118);
nor U3053 (N_3053,In_576,In_253);
xnor U3054 (N_3054,In_590,In_186);
or U3055 (N_3055,In_821,In_861);
nand U3056 (N_3056,In_773,In_141);
nand U3057 (N_3057,In_350,In_237);
and U3058 (N_3058,In_395,In_256);
or U3059 (N_3059,In_612,In_567);
nand U3060 (N_3060,In_517,In_210);
nand U3061 (N_3061,In_223,In_98);
and U3062 (N_3062,In_95,In_317);
nor U3063 (N_3063,In_274,In_462);
and U3064 (N_3064,In_562,In_809);
nor U3065 (N_3065,In_653,In_536);
or U3066 (N_3066,In_801,In_361);
nand U3067 (N_3067,In_848,In_713);
or U3068 (N_3068,In_811,In_358);
nand U3069 (N_3069,In_847,In_722);
nor U3070 (N_3070,In_878,In_450);
nand U3071 (N_3071,In_368,In_636);
or U3072 (N_3072,In_236,In_4);
nand U3073 (N_3073,In_939,In_480);
nand U3074 (N_3074,In_243,In_585);
nor U3075 (N_3075,In_782,In_708);
nor U3076 (N_3076,In_624,In_895);
or U3077 (N_3077,In_506,In_627);
nand U3078 (N_3078,In_474,In_209);
nand U3079 (N_3079,In_872,In_97);
nand U3080 (N_3080,In_228,In_230);
xor U3081 (N_3081,In_268,In_23);
or U3082 (N_3082,In_19,In_878);
and U3083 (N_3083,In_609,In_21);
or U3084 (N_3084,In_994,In_503);
nor U3085 (N_3085,In_261,In_483);
or U3086 (N_3086,In_50,In_173);
and U3087 (N_3087,In_689,In_99);
nor U3088 (N_3088,In_852,In_366);
nand U3089 (N_3089,In_562,In_814);
and U3090 (N_3090,In_455,In_298);
nor U3091 (N_3091,In_824,In_209);
and U3092 (N_3092,In_480,In_906);
or U3093 (N_3093,In_46,In_432);
and U3094 (N_3094,In_925,In_984);
nand U3095 (N_3095,In_147,In_468);
nor U3096 (N_3096,In_403,In_37);
or U3097 (N_3097,In_40,In_438);
or U3098 (N_3098,In_905,In_914);
nor U3099 (N_3099,In_686,In_827);
nor U3100 (N_3100,In_762,In_471);
nand U3101 (N_3101,In_774,In_55);
or U3102 (N_3102,In_519,In_430);
and U3103 (N_3103,In_551,In_186);
nand U3104 (N_3104,In_484,In_941);
or U3105 (N_3105,In_184,In_374);
nand U3106 (N_3106,In_699,In_636);
nand U3107 (N_3107,In_999,In_43);
and U3108 (N_3108,In_438,In_890);
nor U3109 (N_3109,In_684,In_927);
or U3110 (N_3110,In_9,In_526);
and U3111 (N_3111,In_604,In_969);
nor U3112 (N_3112,In_741,In_492);
or U3113 (N_3113,In_343,In_550);
or U3114 (N_3114,In_640,In_945);
nand U3115 (N_3115,In_510,In_774);
or U3116 (N_3116,In_617,In_197);
and U3117 (N_3117,In_799,In_68);
nand U3118 (N_3118,In_347,In_79);
or U3119 (N_3119,In_956,In_779);
nand U3120 (N_3120,In_947,In_556);
and U3121 (N_3121,In_519,In_4);
nor U3122 (N_3122,In_168,In_465);
or U3123 (N_3123,In_618,In_541);
xor U3124 (N_3124,In_369,In_633);
and U3125 (N_3125,In_820,In_465);
or U3126 (N_3126,In_582,In_415);
and U3127 (N_3127,In_9,In_762);
or U3128 (N_3128,In_330,In_10);
or U3129 (N_3129,In_945,In_639);
nor U3130 (N_3130,In_526,In_867);
nor U3131 (N_3131,In_842,In_101);
nand U3132 (N_3132,In_387,In_462);
or U3133 (N_3133,In_332,In_166);
nor U3134 (N_3134,In_536,In_697);
and U3135 (N_3135,In_99,In_552);
or U3136 (N_3136,In_185,In_388);
nand U3137 (N_3137,In_545,In_860);
or U3138 (N_3138,In_462,In_628);
or U3139 (N_3139,In_419,In_491);
nand U3140 (N_3140,In_858,In_203);
nand U3141 (N_3141,In_276,In_404);
and U3142 (N_3142,In_880,In_710);
and U3143 (N_3143,In_282,In_705);
nand U3144 (N_3144,In_584,In_457);
nor U3145 (N_3145,In_939,In_793);
and U3146 (N_3146,In_193,In_151);
nand U3147 (N_3147,In_426,In_301);
xor U3148 (N_3148,In_64,In_69);
nor U3149 (N_3149,In_497,In_509);
or U3150 (N_3150,In_657,In_56);
nand U3151 (N_3151,In_396,In_18);
nand U3152 (N_3152,In_372,In_91);
or U3153 (N_3153,In_894,In_362);
or U3154 (N_3154,In_872,In_815);
or U3155 (N_3155,In_953,In_539);
nand U3156 (N_3156,In_631,In_67);
and U3157 (N_3157,In_235,In_565);
or U3158 (N_3158,In_942,In_609);
and U3159 (N_3159,In_526,In_974);
nor U3160 (N_3160,In_395,In_551);
or U3161 (N_3161,In_976,In_428);
nor U3162 (N_3162,In_468,In_447);
nor U3163 (N_3163,In_269,In_356);
or U3164 (N_3164,In_311,In_472);
nand U3165 (N_3165,In_485,In_628);
nand U3166 (N_3166,In_389,In_996);
nor U3167 (N_3167,In_818,In_310);
nor U3168 (N_3168,In_155,In_573);
nor U3169 (N_3169,In_359,In_975);
nor U3170 (N_3170,In_714,In_834);
nor U3171 (N_3171,In_147,In_884);
nor U3172 (N_3172,In_176,In_487);
and U3173 (N_3173,In_366,In_418);
or U3174 (N_3174,In_437,In_274);
or U3175 (N_3175,In_333,In_707);
nor U3176 (N_3176,In_415,In_330);
nor U3177 (N_3177,In_386,In_888);
or U3178 (N_3178,In_590,In_802);
xor U3179 (N_3179,In_656,In_273);
or U3180 (N_3180,In_168,In_55);
nand U3181 (N_3181,In_765,In_403);
nand U3182 (N_3182,In_455,In_990);
xor U3183 (N_3183,In_813,In_609);
or U3184 (N_3184,In_733,In_213);
nand U3185 (N_3185,In_183,In_56);
and U3186 (N_3186,In_315,In_820);
nand U3187 (N_3187,In_668,In_459);
nand U3188 (N_3188,In_543,In_187);
or U3189 (N_3189,In_741,In_753);
nand U3190 (N_3190,In_54,In_766);
or U3191 (N_3191,In_904,In_479);
or U3192 (N_3192,In_237,In_474);
and U3193 (N_3193,In_172,In_327);
or U3194 (N_3194,In_316,In_286);
xor U3195 (N_3195,In_545,In_707);
or U3196 (N_3196,In_477,In_570);
or U3197 (N_3197,In_843,In_483);
and U3198 (N_3198,In_914,In_807);
nor U3199 (N_3199,In_483,In_394);
xnor U3200 (N_3200,In_294,In_463);
xnor U3201 (N_3201,In_928,In_270);
nand U3202 (N_3202,In_896,In_252);
nor U3203 (N_3203,In_196,In_357);
or U3204 (N_3204,In_81,In_638);
or U3205 (N_3205,In_604,In_470);
and U3206 (N_3206,In_44,In_953);
and U3207 (N_3207,In_960,In_236);
or U3208 (N_3208,In_83,In_101);
or U3209 (N_3209,In_573,In_276);
nor U3210 (N_3210,In_792,In_456);
or U3211 (N_3211,In_242,In_928);
or U3212 (N_3212,In_112,In_427);
or U3213 (N_3213,In_639,In_149);
or U3214 (N_3214,In_484,In_581);
and U3215 (N_3215,In_207,In_412);
nand U3216 (N_3216,In_451,In_190);
nor U3217 (N_3217,In_157,In_133);
and U3218 (N_3218,In_626,In_874);
nand U3219 (N_3219,In_569,In_493);
xor U3220 (N_3220,In_2,In_690);
nor U3221 (N_3221,In_49,In_425);
nand U3222 (N_3222,In_971,In_818);
and U3223 (N_3223,In_193,In_938);
nor U3224 (N_3224,In_303,In_465);
and U3225 (N_3225,In_538,In_990);
and U3226 (N_3226,In_782,In_678);
and U3227 (N_3227,In_121,In_829);
and U3228 (N_3228,In_503,In_596);
or U3229 (N_3229,In_276,In_310);
or U3230 (N_3230,In_631,In_615);
and U3231 (N_3231,In_176,In_692);
and U3232 (N_3232,In_141,In_284);
and U3233 (N_3233,In_15,In_433);
nor U3234 (N_3234,In_327,In_217);
or U3235 (N_3235,In_779,In_186);
and U3236 (N_3236,In_553,In_274);
nor U3237 (N_3237,In_568,In_667);
and U3238 (N_3238,In_397,In_457);
or U3239 (N_3239,In_147,In_776);
or U3240 (N_3240,In_242,In_737);
nand U3241 (N_3241,In_596,In_583);
and U3242 (N_3242,In_880,In_490);
and U3243 (N_3243,In_425,In_191);
nor U3244 (N_3244,In_773,In_575);
nand U3245 (N_3245,In_672,In_872);
nand U3246 (N_3246,In_458,In_619);
nand U3247 (N_3247,In_756,In_212);
nor U3248 (N_3248,In_768,In_253);
nor U3249 (N_3249,In_816,In_838);
nor U3250 (N_3250,In_171,In_256);
nor U3251 (N_3251,In_510,In_555);
and U3252 (N_3252,In_8,In_582);
and U3253 (N_3253,In_679,In_80);
nor U3254 (N_3254,In_568,In_577);
and U3255 (N_3255,In_96,In_720);
and U3256 (N_3256,In_90,In_543);
nor U3257 (N_3257,In_926,In_755);
or U3258 (N_3258,In_60,In_27);
nand U3259 (N_3259,In_629,In_241);
or U3260 (N_3260,In_297,In_812);
nor U3261 (N_3261,In_295,In_241);
or U3262 (N_3262,In_799,In_109);
or U3263 (N_3263,In_116,In_170);
nor U3264 (N_3264,In_220,In_550);
or U3265 (N_3265,In_26,In_44);
or U3266 (N_3266,In_30,In_579);
and U3267 (N_3267,In_414,In_38);
and U3268 (N_3268,In_194,In_689);
nor U3269 (N_3269,In_504,In_584);
nor U3270 (N_3270,In_304,In_294);
or U3271 (N_3271,In_306,In_41);
nor U3272 (N_3272,In_161,In_920);
nand U3273 (N_3273,In_606,In_868);
or U3274 (N_3274,In_997,In_759);
or U3275 (N_3275,In_249,In_334);
nand U3276 (N_3276,In_583,In_304);
nand U3277 (N_3277,In_203,In_177);
nor U3278 (N_3278,In_418,In_437);
or U3279 (N_3279,In_900,In_498);
nor U3280 (N_3280,In_58,In_708);
xnor U3281 (N_3281,In_697,In_68);
and U3282 (N_3282,In_342,In_449);
and U3283 (N_3283,In_158,In_854);
nand U3284 (N_3284,In_609,In_694);
or U3285 (N_3285,In_192,In_763);
or U3286 (N_3286,In_761,In_801);
and U3287 (N_3287,In_648,In_775);
or U3288 (N_3288,In_974,In_682);
nand U3289 (N_3289,In_914,In_935);
nor U3290 (N_3290,In_726,In_379);
nor U3291 (N_3291,In_307,In_323);
nor U3292 (N_3292,In_384,In_96);
or U3293 (N_3293,In_507,In_612);
nand U3294 (N_3294,In_817,In_775);
nand U3295 (N_3295,In_644,In_208);
and U3296 (N_3296,In_688,In_250);
nand U3297 (N_3297,In_700,In_3);
xor U3298 (N_3298,In_72,In_274);
and U3299 (N_3299,In_29,In_553);
nand U3300 (N_3300,In_776,In_368);
nor U3301 (N_3301,In_513,In_456);
nand U3302 (N_3302,In_730,In_857);
nor U3303 (N_3303,In_792,In_341);
and U3304 (N_3304,In_95,In_51);
and U3305 (N_3305,In_965,In_236);
nor U3306 (N_3306,In_984,In_898);
or U3307 (N_3307,In_760,In_681);
xnor U3308 (N_3308,In_972,In_456);
nand U3309 (N_3309,In_433,In_992);
nor U3310 (N_3310,In_307,In_128);
nand U3311 (N_3311,In_966,In_279);
and U3312 (N_3312,In_380,In_750);
or U3313 (N_3313,In_542,In_140);
xor U3314 (N_3314,In_38,In_598);
nor U3315 (N_3315,In_81,In_844);
or U3316 (N_3316,In_285,In_617);
nor U3317 (N_3317,In_76,In_415);
and U3318 (N_3318,In_82,In_49);
nor U3319 (N_3319,In_950,In_398);
or U3320 (N_3320,In_651,In_195);
and U3321 (N_3321,In_133,In_981);
and U3322 (N_3322,In_364,In_412);
nor U3323 (N_3323,In_619,In_911);
and U3324 (N_3324,In_440,In_774);
or U3325 (N_3325,In_52,In_720);
or U3326 (N_3326,In_704,In_871);
or U3327 (N_3327,In_694,In_68);
or U3328 (N_3328,In_880,In_434);
nand U3329 (N_3329,In_740,In_237);
and U3330 (N_3330,In_587,In_217);
nand U3331 (N_3331,In_816,In_877);
nand U3332 (N_3332,In_275,In_923);
and U3333 (N_3333,In_430,In_270);
and U3334 (N_3334,In_275,In_614);
or U3335 (N_3335,In_333,In_363);
nor U3336 (N_3336,In_657,In_409);
nand U3337 (N_3337,In_141,In_586);
and U3338 (N_3338,In_41,In_747);
nand U3339 (N_3339,In_277,In_578);
nor U3340 (N_3340,In_6,In_259);
or U3341 (N_3341,In_817,In_755);
or U3342 (N_3342,In_502,In_569);
or U3343 (N_3343,In_180,In_897);
nor U3344 (N_3344,In_355,In_854);
nor U3345 (N_3345,In_863,In_860);
nor U3346 (N_3346,In_912,In_273);
nand U3347 (N_3347,In_819,In_864);
or U3348 (N_3348,In_680,In_971);
or U3349 (N_3349,In_601,In_793);
nand U3350 (N_3350,In_287,In_954);
or U3351 (N_3351,In_254,In_113);
and U3352 (N_3352,In_726,In_316);
or U3353 (N_3353,In_445,In_103);
or U3354 (N_3354,In_973,In_330);
and U3355 (N_3355,In_434,In_366);
and U3356 (N_3356,In_163,In_390);
nor U3357 (N_3357,In_878,In_442);
nor U3358 (N_3358,In_903,In_467);
nor U3359 (N_3359,In_348,In_482);
nor U3360 (N_3360,In_907,In_434);
nor U3361 (N_3361,In_413,In_30);
or U3362 (N_3362,In_777,In_849);
nor U3363 (N_3363,In_274,In_668);
and U3364 (N_3364,In_942,In_514);
and U3365 (N_3365,In_305,In_532);
or U3366 (N_3366,In_882,In_947);
and U3367 (N_3367,In_473,In_878);
or U3368 (N_3368,In_627,In_360);
and U3369 (N_3369,In_354,In_188);
nor U3370 (N_3370,In_282,In_60);
or U3371 (N_3371,In_521,In_453);
nand U3372 (N_3372,In_359,In_226);
and U3373 (N_3373,In_763,In_375);
xnor U3374 (N_3374,In_152,In_833);
nand U3375 (N_3375,In_893,In_337);
or U3376 (N_3376,In_868,In_711);
nor U3377 (N_3377,In_568,In_65);
nand U3378 (N_3378,In_584,In_677);
nor U3379 (N_3379,In_616,In_643);
nand U3380 (N_3380,In_553,In_877);
nand U3381 (N_3381,In_587,In_452);
nand U3382 (N_3382,In_838,In_286);
nor U3383 (N_3383,In_241,In_111);
or U3384 (N_3384,In_823,In_945);
nand U3385 (N_3385,In_134,In_934);
nor U3386 (N_3386,In_119,In_479);
nor U3387 (N_3387,In_276,In_325);
and U3388 (N_3388,In_743,In_462);
or U3389 (N_3389,In_657,In_509);
and U3390 (N_3390,In_892,In_621);
and U3391 (N_3391,In_369,In_606);
nor U3392 (N_3392,In_750,In_720);
nand U3393 (N_3393,In_397,In_635);
nand U3394 (N_3394,In_260,In_107);
and U3395 (N_3395,In_993,In_225);
nor U3396 (N_3396,In_590,In_805);
and U3397 (N_3397,In_396,In_374);
nor U3398 (N_3398,In_153,In_104);
and U3399 (N_3399,In_710,In_233);
or U3400 (N_3400,In_431,In_116);
and U3401 (N_3401,In_37,In_277);
nand U3402 (N_3402,In_787,In_813);
and U3403 (N_3403,In_881,In_185);
nor U3404 (N_3404,In_130,In_890);
nor U3405 (N_3405,In_664,In_966);
or U3406 (N_3406,In_35,In_230);
and U3407 (N_3407,In_633,In_753);
and U3408 (N_3408,In_918,In_221);
and U3409 (N_3409,In_140,In_640);
and U3410 (N_3410,In_934,In_360);
or U3411 (N_3411,In_904,In_777);
nand U3412 (N_3412,In_543,In_399);
nor U3413 (N_3413,In_935,In_633);
nand U3414 (N_3414,In_967,In_17);
and U3415 (N_3415,In_162,In_102);
nand U3416 (N_3416,In_819,In_21);
nor U3417 (N_3417,In_485,In_645);
and U3418 (N_3418,In_844,In_376);
or U3419 (N_3419,In_921,In_196);
and U3420 (N_3420,In_330,In_225);
nand U3421 (N_3421,In_714,In_982);
and U3422 (N_3422,In_968,In_762);
nand U3423 (N_3423,In_920,In_237);
nor U3424 (N_3424,In_937,In_931);
and U3425 (N_3425,In_23,In_27);
nor U3426 (N_3426,In_244,In_743);
nor U3427 (N_3427,In_103,In_533);
nand U3428 (N_3428,In_473,In_84);
nor U3429 (N_3429,In_304,In_611);
or U3430 (N_3430,In_144,In_407);
or U3431 (N_3431,In_198,In_976);
or U3432 (N_3432,In_652,In_934);
nand U3433 (N_3433,In_596,In_924);
nand U3434 (N_3434,In_642,In_370);
nor U3435 (N_3435,In_322,In_139);
and U3436 (N_3436,In_388,In_335);
nand U3437 (N_3437,In_764,In_92);
nand U3438 (N_3438,In_610,In_750);
and U3439 (N_3439,In_353,In_943);
nor U3440 (N_3440,In_472,In_292);
nand U3441 (N_3441,In_572,In_20);
nor U3442 (N_3442,In_684,In_824);
nand U3443 (N_3443,In_331,In_174);
or U3444 (N_3444,In_537,In_831);
and U3445 (N_3445,In_140,In_141);
and U3446 (N_3446,In_547,In_517);
or U3447 (N_3447,In_926,In_82);
or U3448 (N_3448,In_931,In_948);
and U3449 (N_3449,In_466,In_17);
nor U3450 (N_3450,In_969,In_382);
or U3451 (N_3451,In_476,In_4);
nand U3452 (N_3452,In_888,In_305);
nor U3453 (N_3453,In_307,In_713);
nor U3454 (N_3454,In_159,In_418);
nor U3455 (N_3455,In_23,In_438);
or U3456 (N_3456,In_438,In_495);
nor U3457 (N_3457,In_854,In_982);
nor U3458 (N_3458,In_90,In_338);
nand U3459 (N_3459,In_675,In_609);
and U3460 (N_3460,In_945,In_478);
and U3461 (N_3461,In_994,In_83);
nor U3462 (N_3462,In_9,In_10);
and U3463 (N_3463,In_701,In_217);
and U3464 (N_3464,In_404,In_610);
nand U3465 (N_3465,In_371,In_387);
or U3466 (N_3466,In_329,In_138);
or U3467 (N_3467,In_851,In_383);
xor U3468 (N_3468,In_111,In_646);
xor U3469 (N_3469,In_769,In_840);
nor U3470 (N_3470,In_734,In_4);
xor U3471 (N_3471,In_730,In_600);
nand U3472 (N_3472,In_154,In_788);
and U3473 (N_3473,In_897,In_832);
xnor U3474 (N_3474,In_78,In_615);
or U3475 (N_3475,In_439,In_756);
or U3476 (N_3476,In_547,In_38);
or U3477 (N_3477,In_633,In_902);
or U3478 (N_3478,In_56,In_526);
and U3479 (N_3479,In_314,In_90);
nand U3480 (N_3480,In_41,In_243);
and U3481 (N_3481,In_226,In_9);
or U3482 (N_3482,In_697,In_371);
and U3483 (N_3483,In_105,In_98);
nand U3484 (N_3484,In_878,In_59);
nand U3485 (N_3485,In_893,In_573);
and U3486 (N_3486,In_395,In_520);
or U3487 (N_3487,In_664,In_900);
nor U3488 (N_3488,In_32,In_323);
and U3489 (N_3489,In_412,In_897);
or U3490 (N_3490,In_139,In_925);
nor U3491 (N_3491,In_331,In_970);
nand U3492 (N_3492,In_338,In_173);
or U3493 (N_3493,In_648,In_272);
nand U3494 (N_3494,In_366,In_868);
xnor U3495 (N_3495,In_568,In_422);
or U3496 (N_3496,In_371,In_340);
or U3497 (N_3497,In_734,In_217);
nand U3498 (N_3498,In_934,In_705);
and U3499 (N_3499,In_362,In_803);
and U3500 (N_3500,In_450,In_630);
xnor U3501 (N_3501,In_318,In_454);
and U3502 (N_3502,In_189,In_54);
nor U3503 (N_3503,In_235,In_72);
or U3504 (N_3504,In_211,In_166);
and U3505 (N_3505,In_623,In_453);
nor U3506 (N_3506,In_876,In_925);
nor U3507 (N_3507,In_23,In_592);
nand U3508 (N_3508,In_112,In_925);
or U3509 (N_3509,In_106,In_543);
nor U3510 (N_3510,In_767,In_70);
or U3511 (N_3511,In_852,In_543);
or U3512 (N_3512,In_883,In_303);
or U3513 (N_3513,In_982,In_847);
xor U3514 (N_3514,In_12,In_457);
or U3515 (N_3515,In_822,In_813);
or U3516 (N_3516,In_97,In_815);
or U3517 (N_3517,In_154,In_542);
or U3518 (N_3518,In_317,In_150);
or U3519 (N_3519,In_480,In_360);
nor U3520 (N_3520,In_595,In_497);
nand U3521 (N_3521,In_647,In_144);
nor U3522 (N_3522,In_117,In_86);
nor U3523 (N_3523,In_548,In_705);
or U3524 (N_3524,In_974,In_170);
and U3525 (N_3525,In_274,In_277);
nand U3526 (N_3526,In_349,In_541);
and U3527 (N_3527,In_138,In_747);
and U3528 (N_3528,In_901,In_563);
or U3529 (N_3529,In_532,In_732);
and U3530 (N_3530,In_283,In_592);
and U3531 (N_3531,In_295,In_740);
and U3532 (N_3532,In_795,In_447);
xnor U3533 (N_3533,In_307,In_394);
nor U3534 (N_3534,In_798,In_245);
nor U3535 (N_3535,In_461,In_718);
or U3536 (N_3536,In_314,In_219);
nand U3537 (N_3537,In_55,In_161);
nand U3538 (N_3538,In_888,In_921);
or U3539 (N_3539,In_185,In_861);
nand U3540 (N_3540,In_939,In_732);
nand U3541 (N_3541,In_405,In_504);
and U3542 (N_3542,In_107,In_956);
nand U3543 (N_3543,In_895,In_105);
nor U3544 (N_3544,In_204,In_715);
and U3545 (N_3545,In_107,In_909);
nor U3546 (N_3546,In_828,In_7);
and U3547 (N_3547,In_436,In_51);
xnor U3548 (N_3548,In_894,In_170);
and U3549 (N_3549,In_698,In_14);
nand U3550 (N_3550,In_254,In_402);
nand U3551 (N_3551,In_154,In_239);
and U3552 (N_3552,In_116,In_135);
or U3553 (N_3553,In_882,In_337);
nor U3554 (N_3554,In_966,In_461);
nand U3555 (N_3555,In_421,In_776);
nor U3556 (N_3556,In_146,In_563);
nand U3557 (N_3557,In_466,In_43);
nor U3558 (N_3558,In_751,In_907);
and U3559 (N_3559,In_2,In_297);
and U3560 (N_3560,In_887,In_98);
and U3561 (N_3561,In_784,In_651);
nor U3562 (N_3562,In_810,In_801);
nor U3563 (N_3563,In_587,In_951);
and U3564 (N_3564,In_829,In_489);
or U3565 (N_3565,In_943,In_727);
nand U3566 (N_3566,In_9,In_138);
nand U3567 (N_3567,In_34,In_947);
and U3568 (N_3568,In_350,In_828);
or U3569 (N_3569,In_21,In_658);
or U3570 (N_3570,In_684,In_217);
nor U3571 (N_3571,In_611,In_132);
and U3572 (N_3572,In_975,In_657);
or U3573 (N_3573,In_423,In_659);
nand U3574 (N_3574,In_336,In_39);
and U3575 (N_3575,In_954,In_160);
and U3576 (N_3576,In_39,In_457);
nand U3577 (N_3577,In_25,In_609);
or U3578 (N_3578,In_487,In_444);
nor U3579 (N_3579,In_637,In_25);
xnor U3580 (N_3580,In_646,In_985);
nor U3581 (N_3581,In_673,In_306);
nand U3582 (N_3582,In_791,In_126);
or U3583 (N_3583,In_635,In_791);
nand U3584 (N_3584,In_504,In_952);
nand U3585 (N_3585,In_303,In_925);
or U3586 (N_3586,In_36,In_227);
nand U3587 (N_3587,In_715,In_509);
nand U3588 (N_3588,In_890,In_52);
nand U3589 (N_3589,In_328,In_494);
and U3590 (N_3590,In_818,In_413);
or U3591 (N_3591,In_879,In_994);
nand U3592 (N_3592,In_210,In_515);
or U3593 (N_3593,In_685,In_125);
nand U3594 (N_3594,In_756,In_279);
nor U3595 (N_3595,In_616,In_873);
or U3596 (N_3596,In_324,In_239);
or U3597 (N_3597,In_679,In_696);
or U3598 (N_3598,In_44,In_483);
nand U3599 (N_3599,In_595,In_512);
nor U3600 (N_3600,In_218,In_632);
nand U3601 (N_3601,In_888,In_945);
and U3602 (N_3602,In_747,In_26);
nand U3603 (N_3603,In_352,In_203);
nor U3604 (N_3604,In_60,In_132);
nor U3605 (N_3605,In_130,In_518);
or U3606 (N_3606,In_17,In_932);
or U3607 (N_3607,In_452,In_179);
nor U3608 (N_3608,In_782,In_27);
or U3609 (N_3609,In_863,In_567);
nor U3610 (N_3610,In_773,In_757);
or U3611 (N_3611,In_80,In_945);
and U3612 (N_3612,In_133,In_688);
and U3613 (N_3613,In_63,In_240);
nor U3614 (N_3614,In_954,In_46);
nor U3615 (N_3615,In_121,In_374);
and U3616 (N_3616,In_658,In_665);
nand U3617 (N_3617,In_801,In_482);
nand U3618 (N_3618,In_876,In_696);
and U3619 (N_3619,In_210,In_990);
nand U3620 (N_3620,In_180,In_307);
nand U3621 (N_3621,In_314,In_187);
and U3622 (N_3622,In_413,In_274);
nand U3623 (N_3623,In_980,In_421);
nand U3624 (N_3624,In_756,In_851);
or U3625 (N_3625,In_929,In_788);
and U3626 (N_3626,In_334,In_479);
and U3627 (N_3627,In_506,In_429);
xor U3628 (N_3628,In_760,In_408);
nor U3629 (N_3629,In_514,In_239);
or U3630 (N_3630,In_642,In_611);
or U3631 (N_3631,In_653,In_481);
nor U3632 (N_3632,In_877,In_893);
and U3633 (N_3633,In_370,In_282);
and U3634 (N_3634,In_546,In_793);
nand U3635 (N_3635,In_376,In_968);
nand U3636 (N_3636,In_264,In_342);
nand U3637 (N_3637,In_936,In_640);
and U3638 (N_3638,In_896,In_4);
or U3639 (N_3639,In_22,In_636);
and U3640 (N_3640,In_898,In_335);
or U3641 (N_3641,In_197,In_615);
nor U3642 (N_3642,In_358,In_764);
or U3643 (N_3643,In_869,In_495);
nor U3644 (N_3644,In_479,In_259);
or U3645 (N_3645,In_761,In_790);
nand U3646 (N_3646,In_550,In_681);
and U3647 (N_3647,In_256,In_873);
nand U3648 (N_3648,In_966,In_416);
nor U3649 (N_3649,In_466,In_585);
nand U3650 (N_3650,In_403,In_830);
and U3651 (N_3651,In_914,In_171);
or U3652 (N_3652,In_263,In_238);
and U3653 (N_3653,In_37,In_158);
and U3654 (N_3654,In_134,In_526);
xor U3655 (N_3655,In_248,In_802);
or U3656 (N_3656,In_602,In_273);
nand U3657 (N_3657,In_249,In_509);
or U3658 (N_3658,In_964,In_471);
or U3659 (N_3659,In_628,In_391);
nand U3660 (N_3660,In_485,In_61);
nand U3661 (N_3661,In_172,In_288);
nor U3662 (N_3662,In_300,In_948);
nor U3663 (N_3663,In_143,In_901);
and U3664 (N_3664,In_738,In_22);
nand U3665 (N_3665,In_902,In_290);
nor U3666 (N_3666,In_501,In_250);
nor U3667 (N_3667,In_776,In_850);
nand U3668 (N_3668,In_803,In_154);
nor U3669 (N_3669,In_693,In_827);
or U3670 (N_3670,In_521,In_592);
nor U3671 (N_3671,In_654,In_255);
nand U3672 (N_3672,In_255,In_273);
or U3673 (N_3673,In_418,In_276);
or U3674 (N_3674,In_925,In_72);
or U3675 (N_3675,In_693,In_492);
or U3676 (N_3676,In_866,In_267);
or U3677 (N_3677,In_298,In_825);
xnor U3678 (N_3678,In_156,In_89);
nor U3679 (N_3679,In_645,In_539);
and U3680 (N_3680,In_155,In_918);
or U3681 (N_3681,In_307,In_940);
nand U3682 (N_3682,In_962,In_74);
or U3683 (N_3683,In_658,In_224);
nor U3684 (N_3684,In_908,In_220);
nor U3685 (N_3685,In_702,In_83);
or U3686 (N_3686,In_679,In_722);
or U3687 (N_3687,In_192,In_550);
nand U3688 (N_3688,In_631,In_970);
or U3689 (N_3689,In_356,In_478);
and U3690 (N_3690,In_764,In_634);
nor U3691 (N_3691,In_676,In_552);
xor U3692 (N_3692,In_105,In_384);
or U3693 (N_3693,In_58,In_365);
and U3694 (N_3694,In_352,In_595);
nand U3695 (N_3695,In_489,In_962);
nand U3696 (N_3696,In_210,In_547);
and U3697 (N_3697,In_514,In_241);
or U3698 (N_3698,In_527,In_556);
and U3699 (N_3699,In_777,In_301);
nor U3700 (N_3700,In_271,In_912);
nor U3701 (N_3701,In_401,In_646);
and U3702 (N_3702,In_316,In_149);
or U3703 (N_3703,In_52,In_725);
nand U3704 (N_3704,In_125,In_409);
and U3705 (N_3705,In_612,In_62);
and U3706 (N_3706,In_447,In_63);
nor U3707 (N_3707,In_928,In_516);
and U3708 (N_3708,In_66,In_734);
or U3709 (N_3709,In_359,In_229);
or U3710 (N_3710,In_620,In_228);
nand U3711 (N_3711,In_511,In_869);
or U3712 (N_3712,In_591,In_933);
xnor U3713 (N_3713,In_292,In_390);
and U3714 (N_3714,In_345,In_951);
nor U3715 (N_3715,In_970,In_519);
nor U3716 (N_3716,In_448,In_12);
and U3717 (N_3717,In_383,In_3);
and U3718 (N_3718,In_337,In_654);
nand U3719 (N_3719,In_443,In_479);
nand U3720 (N_3720,In_282,In_329);
xnor U3721 (N_3721,In_199,In_442);
nand U3722 (N_3722,In_824,In_786);
nand U3723 (N_3723,In_197,In_101);
or U3724 (N_3724,In_598,In_680);
nor U3725 (N_3725,In_338,In_174);
nand U3726 (N_3726,In_813,In_603);
or U3727 (N_3727,In_444,In_9);
nand U3728 (N_3728,In_834,In_651);
or U3729 (N_3729,In_789,In_55);
nor U3730 (N_3730,In_145,In_503);
nand U3731 (N_3731,In_494,In_230);
and U3732 (N_3732,In_44,In_695);
or U3733 (N_3733,In_901,In_584);
or U3734 (N_3734,In_254,In_476);
or U3735 (N_3735,In_351,In_952);
or U3736 (N_3736,In_380,In_640);
nor U3737 (N_3737,In_562,In_93);
nor U3738 (N_3738,In_240,In_79);
nand U3739 (N_3739,In_312,In_508);
or U3740 (N_3740,In_21,In_47);
or U3741 (N_3741,In_283,In_422);
nor U3742 (N_3742,In_772,In_233);
and U3743 (N_3743,In_424,In_941);
nand U3744 (N_3744,In_62,In_447);
and U3745 (N_3745,In_754,In_20);
nand U3746 (N_3746,In_366,In_355);
nand U3747 (N_3747,In_935,In_495);
or U3748 (N_3748,In_230,In_817);
or U3749 (N_3749,In_780,In_759);
and U3750 (N_3750,In_118,In_402);
or U3751 (N_3751,In_87,In_707);
and U3752 (N_3752,In_954,In_831);
nand U3753 (N_3753,In_950,In_714);
or U3754 (N_3754,In_761,In_218);
nor U3755 (N_3755,In_237,In_389);
and U3756 (N_3756,In_293,In_764);
and U3757 (N_3757,In_527,In_967);
nand U3758 (N_3758,In_222,In_330);
or U3759 (N_3759,In_826,In_614);
or U3760 (N_3760,In_223,In_173);
and U3761 (N_3761,In_389,In_970);
nor U3762 (N_3762,In_463,In_401);
nor U3763 (N_3763,In_485,In_43);
nor U3764 (N_3764,In_766,In_756);
or U3765 (N_3765,In_121,In_109);
and U3766 (N_3766,In_937,In_363);
and U3767 (N_3767,In_261,In_53);
and U3768 (N_3768,In_486,In_25);
or U3769 (N_3769,In_432,In_177);
xor U3770 (N_3770,In_555,In_518);
nand U3771 (N_3771,In_348,In_182);
nor U3772 (N_3772,In_197,In_263);
nor U3773 (N_3773,In_214,In_720);
and U3774 (N_3774,In_630,In_509);
nor U3775 (N_3775,In_442,In_966);
nand U3776 (N_3776,In_777,In_363);
nor U3777 (N_3777,In_894,In_880);
and U3778 (N_3778,In_225,In_190);
nor U3779 (N_3779,In_387,In_588);
nand U3780 (N_3780,In_525,In_502);
nor U3781 (N_3781,In_475,In_922);
and U3782 (N_3782,In_741,In_293);
and U3783 (N_3783,In_296,In_517);
xnor U3784 (N_3784,In_347,In_27);
or U3785 (N_3785,In_764,In_920);
or U3786 (N_3786,In_199,In_812);
or U3787 (N_3787,In_288,In_853);
and U3788 (N_3788,In_978,In_265);
nor U3789 (N_3789,In_29,In_163);
nand U3790 (N_3790,In_791,In_847);
nor U3791 (N_3791,In_949,In_377);
and U3792 (N_3792,In_478,In_790);
nor U3793 (N_3793,In_978,In_584);
or U3794 (N_3794,In_879,In_186);
or U3795 (N_3795,In_74,In_857);
or U3796 (N_3796,In_938,In_433);
and U3797 (N_3797,In_353,In_906);
nand U3798 (N_3798,In_248,In_889);
or U3799 (N_3799,In_996,In_657);
and U3800 (N_3800,In_113,In_670);
and U3801 (N_3801,In_750,In_725);
and U3802 (N_3802,In_945,In_205);
or U3803 (N_3803,In_699,In_870);
and U3804 (N_3804,In_845,In_8);
and U3805 (N_3805,In_564,In_396);
and U3806 (N_3806,In_586,In_334);
nor U3807 (N_3807,In_368,In_860);
or U3808 (N_3808,In_318,In_988);
nor U3809 (N_3809,In_900,In_43);
nand U3810 (N_3810,In_684,In_7);
and U3811 (N_3811,In_874,In_92);
or U3812 (N_3812,In_106,In_275);
or U3813 (N_3813,In_885,In_157);
or U3814 (N_3814,In_1,In_776);
or U3815 (N_3815,In_291,In_89);
nand U3816 (N_3816,In_918,In_26);
xor U3817 (N_3817,In_106,In_704);
and U3818 (N_3818,In_580,In_887);
xor U3819 (N_3819,In_260,In_994);
and U3820 (N_3820,In_443,In_675);
and U3821 (N_3821,In_384,In_34);
nor U3822 (N_3822,In_911,In_862);
and U3823 (N_3823,In_384,In_354);
and U3824 (N_3824,In_473,In_751);
and U3825 (N_3825,In_345,In_436);
xnor U3826 (N_3826,In_243,In_196);
or U3827 (N_3827,In_951,In_524);
nor U3828 (N_3828,In_590,In_31);
or U3829 (N_3829,In_439,In_719);
or U3830 (N_3830,In_627,In_99);
and U3831 (N_3831,In_391,In_512);
nand U3832 (N_3832,In_553,In_612);
or U3833 (N_3833,In_493,In_660);
nand U3834 (N_3834,In_404,In_98);
nand U3835 (N_3835,In_395,In_611);
nor U3836 (N_3836,In_275,In_975);
nand U3837 (N_3837,In_631,In_922);
nand U3838 (N_3838,In_873,In_147);
nand U3839 (N_3839,In_475,In_110);
nand U3840 (N_3840,In_670,In_117);
and U3841 (N_3841,In_107,In_104);
nor U3842 (N_3842,In_450,In_556);
nor U3843 (N_3843,In_924,In_565);
and U3844 (N_3844,In_714,In_875);
nor U3845 (N_3845,In_505,In_341);
and U3846 (N_3846,In_799,In_101);
nand U3847 (N_3847,In_849,In_817);
and U3848 (N_3848,In_136,In_498);
or U3849 (N_3849,In_472,In_715);
or U3850 (N_3850,In_149,In_723);
or U3851 (N_3851,In_844,In_414);
nor U3852 (N_3852,In_140,In_824);
nand U3853 (N_3853,In_751,In_911);
nor U3854 (N_3854,In_527,In_565);
nand U3855 (N_3855,In_132,In_635);
or U3856 (N_3856,In_590,In_51);
nor U3857 (N_3857,In_916,In_932);
nand U3858 (N_3858,In_689,In_819);
nor U3859 (N_3859,In_661,In_786);
or U3860 (N_3860,In_200,In_603);
nor U3861 (N_3861,In_244,In_612);
or U3862 (N_3862,In_396,In_335);
nand U3863 (N_3863,In_692,In_328);
or U3864 (N_3864,In_548,In_865);
and U3865 (N_3865,In_103,In_248);
nor U3866 (N_3866,In_98,In_508);
and U3867 (N_3867,In_923,In_984);
nand U3868 (N_3868,In_0,In_667);
nand U3869 (N_3869,In_80,In_260);
nand U3870 (N_3870,In_774,In_59);
nor U3871 (N_3871,In_369,In_558);
or U3872 (N_3872,In_212,In_392);
and U3873 (N_3873,In_422,In_773);
nand U3874 (N_3874,In_751,In_443);
nor U3875 (N_3875,In_535,In_303);
and U3876 (N_3876,In_789,In_136);
or U3877 (N_3877,In_798,In_455);
and U3878 (N_3878,In_716,In_736);
or U3879 (N_3879,In_2,In_640);
nand U3880 (N_3880,In_311,In_278);
nand U3881 (N_3881,In_1,In_471);
nand U3882 (N_3882,In_863,In_433);
and U3883 (N_3883,In_498,In_281);
nor U3884 (N_3884,In_133,In_763);
or U3885 (N_3885,In_268,In_48);
or U3886 (N_3886,In_457,In_202);
nor U3887 (N_3887,In_914,In_872);
or U3888 (N_3888,In_764,In_277);
or U3889 (N_3889,In_97,In_473);
and U3890 (N_3890,In_414,In_343);
and U3891 (N_3891,In_563,In_878);
or U3892 (N_3892,In_218,In_869);
nor U3893 (N_3893,In_846,In_857);
or U3894 (N_3894,In_125,In_895);
or U3895 (N_3895,In_73,In_297);
nand U3896 (N_3896,In_210,In_70);
nor U3897 (N_3897,In_866,In_151);
and U3898 (N_3898,In_433,In_118);
nand U3899 (N_3899,In_744,In_587);
or U3900 (N_3900,In_365,In_486);
nor U3901 (N_3901,In_671,In_685);
or U3902 (N_3902,In_254,In_67);
and U3903 (N_3903,In_970,In_307);
nand U3904 (N_3904,In_304,In_235);
nand U3905 (N_3905,In_274,In_76);
or U3906 (N_3906,In_296,In_749);
and U3907 (N_3907,In_424,In_152);
nand U3908 (N_3908,In_439,In_172);
or U3909 (N_3909,In_971,In_781);
and U3910 (N_3910,In_340,In_365);
nand U3911 (N_3911,In_545,In_887);
nand U3912 (N_3912,In_778,In_569);
or U3913 (N_3913,In_299,In_768);
nor U3914 (N_3914,In_998,In_662);
and U3915 (N_3915,In_609,In_163);
and U3916 (N_3916,In_900,In_782);
and U3917 (N_3917,In_876,In_916);
or U3918 (N_3918,In_560,In_379);
or U3919 (N_3919,In_662,In_887);
nor U3920 (N_3920,In_650,In_55);
nor U3921 (N_3921,In_818,In_387);
and U3922 (N_3922,In_524,In_99);
nand U3923 (N_3923,In_387,In_693);
nor U3924 (N_3924,In_683,In_406);
and U3925 (N_3925,In_138,In_20);
or U3926 (N_3926,In_571,In_983);
or U3927 (N_3927,In_607,In_705);
nand U3928 (N_3928,In_313,In_653);
nand U3929 (N_3929,In_55,In_992);
nor U3930 (N_3930,In_129,In_346);
and U3931 (N_3931,In_482,In_251);
nor U3932 (N_3932,In_105,In_16);
nor U3933 (N_3933,In_651,In_24);
nand U3934 (N_3934,In_380,In_185);
nand U3935 (N_3935,In_201,In_387);
nor U3936 (N_3936,In_357,In_390);
or U3937 (N_3937,In_965,In_90);
nand U3938 (N_3938,In_985,In_643);
nand U3939 (N_3939,In_850,In_961);
nand U3940 (N_3940,In_409,In_415);
nor U3941 (N_3941,In_728,In_817);
nor U3942 (N_3942,In_335,In_743);
nor U3943 (N_3943,In_572,In_946);
nand U3944 (N_3944,In_893,In_873);
nor U3945 (N_3945,In_48,In_774);
nand U3946 (N_3946,In_78,In_740);
or U3947 (N_3947,In_576,In_963);
or U3948 (N_3948,In_545,In_967);
nand U3949 (N_3949,In_315,In_678);
or U3950 (N_3950,In_646,In_954);
nand U3951 (N_3951,In_510,In_501);
nor U3952 (N_3952,In_379,In_960);
or U3953 (N_3953,In_401,In_567);
nor U3954 (N_3954,In_682,In_110);
and U3955 (N_3955,In_194,In_57);
nor U3956 (N_3956,In_831,In_180);
or U3957 (N_3957,In_181,In_550);
nand U3958 (N_3958,In_408,In_454);
and U3959 (N_3959,In_335,In_909);
nor U3960 (N_3960,In_962,In_841);
nor U3961 (N_3961,In_951,In_510);
nor U3962 (N_3962,In_763,In_94);
or U3963 (N_3963,In_9,In_193);
nand U3964 (N_3964,In_68,In_172);
and U3965 (N_3965,In_896,In_846);
or U3966 (N_3966,In_446,In_167);
and U3967 (N_3967,In_154,In_588);
xor U3968 (N_3968,In_745,In_72);
nand U3969 (N_3969,In_590,In_951);
nand U3970 (N_3970,In_509,In_856);
nand U3971 (N_3971,In_683,In_54);
nand U3972 (N_3972,In_168,In_908);
or U3973 (N_3973,In_401,In_794);
nor U3974 (N_3974,In_819,In_941);
or U3975 (N_3975,In_596,In_204);
and U3976 (N_3976,In_643,In_234);
or U3977 (N_3977,In_349,In_201);
or U3978 (N_3978,In_764,In_474);
and U3979 (N_3979,In_194,In_739);
nor U3980 (N_3980,In_786,In_915);
or U3981 (N_3981,In_814,In_661);
or U3982 (N_3982,In_882,In_316);
or U3983 (N_3983,In_402,In_323);
or U3984 (N_3984,In_500,In_39);
or U3985 (N_3985,In_841,In_918);
and U3986 (N_3986,In_441,In_673);
nor U3987 (N_3987,In_157,In_543);
xnor U3988 (N_3988,In_993,In_758);
nor U3989 (N_3989,In_35,In_779);
nor U3990 (N_3990,In_757,In_170);
and U3991 (N_3991,In_234,In_855);
nand U3992 (N_3992,In_38,In_140);
nand U3993 (N_3993,In_936,In_460);
and U3994 (N_3994,In_513,In_761);
and U3995 (N_3995,In_64,In_112);
nor U3996 (N_3996,In_39,In_160);
nand U3997 (N_3997,In_361,In_671);
nand U3998 (N_3998,In_518,In_73);
or U3999 (N_3999,In_87,In_613);
and U4000 (N_4000,In_819,In_960);
nor U4001 (N_4001,In_566,In_373);
nand U4002 (N_4002,In_69,In_278);
and U4003 (N_4003,In_450,In_69);
nor U4004 (N_4004,In_507,In_189);
nand U4005 (N_4005,In_949,In_933);
or U4006 (N_4006,In_288,In_328);
nor U4007 (N_4007,In_30,In_891);
and U4008 (N_4008,In_430,In_514);
and U4009 (N_4009,In_236,In_106);
and U4010 (N_4010,In_483,In_877);
or U4011 (N_4011,In_74,In_258);
nor U4012 (N_4012,In_340,In_847);
nand U4013 (N_4013,In_370,In_182);
and U4014 (N_4014,In_167,In_497);
nor U4015 (N_4015,In_171,In_586);
or U4016 (N_4016,In_500,In_245);
nand U4017 (N_4017,In_224,In_11);
and U4018 (N_4018,In_883,In_337);
or U4019 (N_4019,In_975,In_742);
xnor U4020 (N_4020,In_585,In_907);
or U4021 (N_4021,In_870,In_649);
and U4022 (N_4022,In_622,In_241);
nand U4023 (N_4023,In_829,In_265);
and U4024 (N_4024,In_251,In_392);
and U4025 (N_4025,In_372,In_880);
and U4026 (N_4026,In_966,In_34);
and U4027 (N_4027,In_130,In_746);
or U4028 (N_4028,In_146,In_110);
or U4029 (N_4029,In_574,In_935);
or U4030 (N_4030,In_367,In_683);
xor U4031 (N_4031,In_479,In_372);
and U4032 (N_4032,In_382,In_495);
or U4033 (N_4033,In_131,In_332);
nand U4034 (N_4034,In_142,In_221);
nor U4035 (N_4035,In_773,In_494);
and U4036 (N_4036,In_310,In_316);
nor U4037 (N_4037,In_870,In_977);
and U4038 (N_4038,In_438,In_434);
or U4039 (N_4039,In_725,In_594);
nand U4040 (N_4040,In_57,In_132);
and U4041 (N_4041,In_492,In_488);
nand U4042 (N_4042,In_155,In_153);
nand U4043 (N_4043,In_31,In_448);
or U4044 (N_4044,In_188,In_756);
nor U4045 (N_4045,In_571,In_883);
nor U4046 (N_4046,In_519,In_867);
nand U4047 (N_4047,In_641,In_614);
nor U4048 (N_4048,In_894,In_221);
nor U4049 (N_4049,In_412,In_914);
nor U4050 (N_4050,In_59,In_109);
nor U4051 (N_4051,In_391,In_702);
xor U4052 (N_4052,In_870,In_206);
nor U4053 (N_4053,In_758,In_285);
nor U4054 (N_4054,In_130,In_36);
nand U4055 (N_4055,In_222,In_186);
or U4056 (N_4056,In_697,In_494);
and U4057 (N_4057,In_425,In_218);
nor U4058 (N_4058,In_440,In_604);
and U4059 (N_4059,In_339,In_750);
nand U4060 (N_4060,In_815,In_720);
nand U4061 (N_4061,In_159,In_947);
and U4062 (N_4062,In_862,In_18);
nand U4063 (N_4063,In_126,In_422);
nor U4064 (N_4064,In_335,In_269);
nand U4065 (N_4065,In_537,In_165);
or U4066 (N_4066,In_697,In_350);
and U4067 (N_4067,In_243,In_215);
nand U4068 (N_4068,In_243,In_248);
or U4069 (N_4069,In_642,In_688);
nand U4070 (N_4070,In_863,In_33);
nand U4071 (N_4071,In_44,In_654);
and U4072 (N_4072,In_434,In_288);
and U4073 (N_4073,In_378,In_236);
nor U4074 (N_4074,In_543,In_950);
and U4075 (N_4075,In_935,In_832);
or U4076 (N_4076,In_220,In_329);
and U4077 (N_4077,In_508,In_138);
nor U4078 (N_4078,In_720,In_873);
nor U4079 (N_4079,In_801,In_699);
or U4080 (N_4080,In_56,In_182);
or U4081 (N_4081,In_229,In_296);
nand U4082 (N_4082,In_926,In_906);
and U4083 (N_4083,In_672,In_709);
or U4084 (N_4084,In_980,In_865);
nor U4085 (N_4085,In_24,In_290);
and U4086 (N_4086,In_913,In_702);
nor U4087 (N_4087,In_400,In_560);
nand U4088 (N_4088,In_987,In_732);
nor U4089 (N_4089,In_789,In_81);
xor U4090 (N_4090,In_392,In_727);
or U4091 (N_4091,In_695,In_972);
nand U4092 (N_4092,In_409,In_516);
nand U4093 (N_4093,In_326,In_370);
and U4094 (N_4094,In_969,In_341);
nand U4095 (N_4095,In_998,In_22);
nor U4096 (N_4096,In_229,In_14);
and U4097 (N_4097,In_399,In_566);
nor U4098 (N_4098,In_367,In_339);
nand U4099 (N_4099,In_466,In_684);
and U4100 (N_4100,In_834,In_163);
nor U4101 (N_4101,In_910,In_325);
nand U4102 (N_4102,In_141,In_631);
nand U4103 (N_4103,In_218,In_437);
nand U4104 (N_4104,In_541,In_977);
or U4105 (N_4105,In_402,In_822);
and U4106 (N_4106,In_21,In_491);
or U4107 (N_4107,In_418,In_774);
and U4108 (N_4108,In_122,In_635);
and U4109 (N_4109,In_141,In_138);
nor U4110 (N_4110,In_427,In_726);
nand U4111 (N_4111,In_100,In_574);
xor U4112 (N_4112,In_930,In_822);
and U4113 (N_4113,In_887,In_328);
nand U4114 (N_4114,In_161,In_159);
and U4115 (N_4115,In_767,In_827);
nand U4116 (N_4116,In_77,In_26);
nor U4117 (N_4117,In_479,In_485);
nor U4118 (N_4118,In_743,In_552);
nand U4119 (N_4119,In_159,In_37);
nand U4120 (N_4120,In_733,In_984);
nand U4121 (N_4121,In_695,In_439);
or U4122 (N_4122,In_906,In_73);
nand U4123 (N_4123,In_30,In_825);
and U4124 (N_4124,In_68,In_540);
and U4125 (N_4125,In_41,In_988);
and U4126 (N_4126,In_499,In_758);
xor U4127 (N_4127,In_911,In_748);
or U4128 (N_4128,In_419,In_476);
or U4129 (N_4129,In_981,In_58);
or U4130 (N_4130,In_682,In_398);
nand U4131 (N_4131,In_970,In_857);
nand U4132 (N_4132,In_88,In_779);
nor U4133 (N_4133,In_358,In_455);
nor U4134 (N_4134,In_906,In_947);
or U4135 (N_4135,In_541,In_43);
or U4136 (N_4136,In_72,In_171);
and U4137 (N_4137,In_610,In_830);
nand U4138 (N_4138,In_579,In_719);
nand U4139 (N_4139,In_833,In_296);
or U4140 (N_4140,In_874,In_117);
or U4141 (N_4141,In_864,In_803);
xnor U4142 (N_4142,In_208,In_12);
xnor U4143 (N_4143,In_64,In_875);
nand U4144 (N_4144,In_937,In_532);
nand U4145 (N_4145,In_103,In_395);
or U4146 (N_4146,In_127,In_303);
nand U4147 (N_4147,In_312,In_349);
nor U4148 (N_4148,In_175,In_651);
or U4149 (N_4149,In_764,In_111);
nor U4150 (N_4150,In_317,In_252);
or U4151 (N_4151,In_445,In_342);
xnor U4152 (N_4152,In_453,In_624);
nand U4153 (N_4153,In_229,In_46);
or U4154 (N_4154,In_549,In_710);
and U4155 (N_4155,In_799,In_263);
nand U4156 (N_4156,In_836,In_22);
nor U4157 (N_4157,In_462,In_983);
nand U4158 (N_4158,In_87,In_289);
nor U4159 (N_4159,In_927,In_154);
and U4160 (N_4160,In_31,In_222);
and U4161 (N_4161,In_514,In_670);
or U4162 (N_4162,In_570,In_463);
nand U4163 (N_4163,In_240,In_200);
or U4164 (N_4164,In_462,In_449);
and U4165 (N_4165,In_401,In_489);
nand U4166 (N_4166,In_646,In_979);
and U4167 (N_4167,In_274,In_286);
nor U4168 (N_4168,In_672,In_389);
xor U4169 (N_4169,In_701,In_583);
nand U4170 (N_4170,In_191,In_310);
or U4171 (N_4171,In_994,In_779);
nor U4172 (N_4172,In_143,In_720);
nand U4173 (N_4173,In_123,In_61);
or U4174 (N_4174,In_750,In_413);
or U4175 (N_4175,In_895,In_455);
or U4176 (N_4176,In_36,In_857);
nor U4177 (N_4177,In_227,In_202);
nor U4178 (N_4178,In_89,In_889);
nor U4179 (N_4179,In_644,In_366);
nor U4180 (N_4180,In_245,In_936);
nor U4181 (N_4181,In_953,In_642);
nand U4182 (N_4182,In_870,In_326);
and U4183 (N_4183,In_187,In_158);
and U4184 (N_4184,In_773,In_800);
and U4185 (N_4185,In_944,In_186);
nand U4186 (N_4186,In_920,In_837);
or U4187 (N_4187,In_989,In_330);
or U4188 (N_4188,In_464,In_597);
nand U4189 (N_4189,In_942,In_487);
nand U4190 (N_4190,In_725,In_580);
nand U4191 (N_4191,In_128,In_929);
nand U4192 (N_4192,In_14,In_139);
and U4193 (N_4193,In_99,In_945);
nand U4194 (N_4194,In_655,In_239);
nor U4195 (N_4195,In_598,In_88);
nor U4196 (N_4196,In_452,In_563);
or U4197 (N_4197,In_32,In_35);
xor U4198 (N_4198,In_519,In_567);
nand U4199 (N_4199,In_871,In_667);
nor U4200 (N_4200,In_927,In_379);
or U4201 (N_4201,In_565,In_530);
nor U4202 (N_4202,In_231,In_847);
or U4203 (N_4203,In_410,In_778);
nand U4204 (N_4204,In_921,In_358);
nor U4205 (N_4205,In_399,In_372);
and U4206 (N_4206,In_324,In_754);
and U4207 (N_4207,In_26,In_522);
nand U4208 (N_4208,In_631,In_374);
nand U4209 (N_4209,In_404,In_71);
and U4210 (N_4210,In_890,In_272);
or U4211 (N_4211,In_128,In_367);
or U4212 (N_4212,In_13,In_99);
nand U4213 (N_4213,In_299,In_617);
nor U4214 (N_4214,In_364,In_862);
nand U4215 (N_4215,In_22,In_677);
and U4216 (N_4216,In_647,In_89);
nand U4217 (N_4217,In_687,In_945);
and U4218 (N_4218,In_612,In_187);
or U4219 (N_4219,In_246,In_910);
and U4220 (N_4220,In_760,In_712);
and U4221 (N_4221,In_813,In_524);
nor U4222 (N_4222,In_469,In_183);
nor U4223 (N_4223,In_392,In_395);
nand U4224 (N_4224,In_319,In_976);
nand U4225 (N_4225,In_515,In_728);
nor U4226 (N_4226,In_291,In_612);
and U4227 (N_4227,In_625,In_230);
and U4228 (N_4228,In_349,In_698);
and U4229 (N_4229,In_191,In_762);
nor U4230 (N_4230,In_133,In_58);
or U4231 (N_4231,In_839,In_992);
nand U4232 (N_4232,In_679,In_762);
nand U4233 (N_4233,In_615,In_533);
or U4234 (N_4234,In_226,In_949);
and U4235 (N_4235,In_669,In_324);
nand U4236 (N_4236,In_201,In_989);
or U4237 (N_4237,In_249,In_582);
nand U4238 (N_4238,In_550,In_451);
nor U4239 (N_4239,In_19,In_486);
and U4240 (N_4240,In_262,In_287);
and U4241 (N_4241,In_118,In_66);
nand U4242 (N_4242,In_387,In_609);
and U4243 (N_4243,In_71,In_79);
or U4244 (N_4244,In_941,In_304);
or U4245 (N_4245,In_492,In_383);
nand U4246 (N_4246,In_89,In_595);
nand U4247 (N_4247,In_179,In_544);
or U4248 (N_4248,In_203,In_782);
nor U4249 (N_4249,In_251,In_761);
nor U4250 (N_4250,In_379,In_976);
and U4251 (N_4251,In_110,In_224);
and U4252 (N_4252,In_109,In_320);
nor U4253 (N_4253,In_631,In_860);
nand U4254 (N_4254,In_761,In_469);
or U4255 (N_4255,In_681,In_534);
or U4256 (N_4256,In_456,In_333);
and U4257 (N_4257,In_264,In_940);
nor U4258 (N_4258,In_526,In_18);
and U4259 (N_4259,In_160,In_484);
and U4260 (N_4260,In_757,In_990);
nor U4261 (N_4261,In_100,In_760);
or U4262 (N_4262,In_652,In_43);
nand U4263 (N_4263,In_33,In_271);
and U4264 (N_4264,In_659,In_376);
nor U4265 (N_4265,In_102,In_902);
or U4266 (N_4266,In_257,In_893);
nand U4267 (N_4267,In_685,In_882);
or U4268 (N_4268,In_50,In_552);
and U4269 (N_4269,In_261,In_954);
and U4270 (N_4270,In_385,In_375);
nor U4271 (N_4271,In_849,In_29);
or U4272 (N_4272,In_484,In_550);
nor U4273 (N_4273,In_586,In_489);
nor U4274 (N_4274,In_352,In_592);
nand U4275 (N_4275,In_888,In_990);
or U4276 (N_4276,In_279,In_919);
or U4277 (N_4277,In_407,In_155);
nand U4278 (N_4278,In_204,In_997);
and U4279 (N_4279,In_948,In_963);
nand U4280 (N_4280,In_357,In_641);
nand U4281 (N_4281,In_446,In_31);
nand U4282 (N_4282,In_644,In_203);
nand U4283 (N_4283,In_77,In_658);
and U4284 (N_4284,In_986,In_579);
xnor U4285 (N_4285,In_682,In_591);
or U4286 (N_4286,In_371,In_728);
nand U4287 (N_4287,In_113,In_91);
nor U4288 (N_4288,In_877,In_802);
or U4289 (N_4289,In_423,In_341);
or U4290 (N_4290,In_142,In_358);
nor U4291 (N_4291,In_237,In_113);
or U4292 (N_4292,In_925,In_56);
and U4293 (N_4293,In_429,In_566);
or U4294 (N_4294,In_836,In_783);
or U4295 (N_4295,In_249,In_657);
nor U4296 (N_4296,In_855,In_916);
and U4297 (N_4297,In_633,In_994);
nor U4298 (N_4298,In_567,In_497);
nand U4299 (N_4299,In_365,In_956);
or U4300 (N_4300,In_113,In_716);
nand U4301 (N_4301,In_240,In_685);
and U4302 (N_4302,In_22,In_565);
nor U4303 (N_4303,In_568,In_991);
nand U4304 (N_4304,In_416,In_492);
nand U4305 (N_4305,In_570,In_537);
or U4306 (N_4306,In_659,In_632);
nand U4307 (N_4307,In_78,In_28);
nand U4308 (N_4308,In_63,In_540);
nand U4309 (N_4309,In_206,In_73);
nor U4310 (N_4310,In_836,In_880);
xnor U4311 (N_4311,In_405,In_610);
or U4312 (N_4312,In_171,In_929);
nand U4313 (N_4313,In_698,In_948);
nor U4314 (N_4314,In_241,In_42);
nor U4315 (N_4315,In_432,In_807);
nor U4316 (N_4316,In_633,In_958);
and U4317 (N_4317,In_410,In_307);
nand U4318 (N_4318,In_204,In_760);
nor U4319 (N_4319,In_589,In_792);
nor U4320 (N_4320,In_526,In_544);
nand U4321 (N_4321,In_670,In_513);
and U4322 (N_4322,In_80,In_794);
or U4323 (N_4323,In_365,In_451);
nand U4324 (N_4324,In_661,In_482);
or U4325 (N_4325,In_107,In_375);
and U4326 (N_4326,In_781,In_579);
and U4327 (N_4327,In_323,In_335);
nand U4328 (N_4328,In_182,In_469);
and U4329 (N_4329,In_940,In_484);
and U4330 (N_4330,In_688,In_913);
nand U4331 (N_4331,In_150,In_308);
nor U4332 (N_4332,In_589,In_748);
nand U4333 (N_4333,In_903,In_241);
and U4334 (N_4334,In_285,In_62);
nand U4335 (N_4335,In_16,In_812);
and U4336 (N_4336,In_484,In_249);
nor U4337 (N_4337,In_184,In_620);
nor U4338 (N_4338,In_427,In_1);
nor U4339 (N_4339,In_484,In_189);
xor U4340 (N_4340,In_78,In_284);
nor U4341 (N_4341,In_412,In_300);
nand U4342 (N_4342,In_957,In_533);
nor U4343 (N_4343,In_698,In_242);
or U4344 (N_4344,In_523,In_756);
nor U4345 (N_4345,In_426,In_258);
or U4346 (N_4346,In_332,In_349);
and U4347 (N_4347,In_645,In_579);
nand U4348 (N_4348,In_704,In_196);
nand U4349 (N_4349,In_766,In_534);
xnor U4350 (N_4350,In_276,In_265);
nand U4351 (N_4351,In_259,In_254);
nor U4352 (N_4352,In_524,In_822);
nand U4353 (N_4353,In_297,In_322);
nor U4354 (N_4354,In_961,In_956);
or U4355 (N_4355,In_426,In_123);
nor U4356 (N_4356,In_310,In_422);
nand U4357 (N_4357,In_287,In_0);
nand U4358 (N_4358,In_68,In_464);
nor U4359 (N_4359,In_570,In_646);
or U4360 (N_4360,In_384,In_630);
and U4361 (N_4361,In_977,In_519);
nor U4362 (N_4362,In_799,In_983);
or U4363 (N_4363,In_829,In_286);
nor U4364 (N_4364,In_302,In_686);
xnor U4365 (N_4365,In_502,In_43);
xor U4366 (N_4366,In_348,In_597);
nor U4367 (N_4367,In_956,In_975);
and U4368 (N_4368,In_687,In_278);
or U4369 (N_4369,In_93,In_552);
nand U4370 (N_4370,In_469,In_584);
nor U4371 (N_4371,In_945,In_593);
or U4372 (N_4372,In_855,In_586);
nor U4373 (N_4373,In_965,In_40);
and U4374 (N_4374,In_617,In_183);
nor U4375 (N_4375,In_232,In_810);
xnor U4376 (N_4376,In_180,In_544);
and U4377 (N_4377,In_563,In_351);
or U4378 (N_4378,In_590,In_85);
nor U4379 (N_4379,In_62,In_189);
nand U4380 (N_4380,In_10,In_459);
nor U4381 (N_4381,In_981,In_168);
nor U4382 (N_4382,In_775,In_276);
nor U4383 (N_4383,In_487,In_312);
and U4384 (N_4384,In_636,In_60);
or U4385 (N_4385,In_919,In_538);
or U4386 (N_4386,In_735,In_293);
or U4387 (N_4387,In_256,In_677);
nand U4388 (N_4388,In_236,In_788);
and U4389 (N_4389,In_79,In_309);
nor U4390 (N_4390,In_294,In_227);
or U4391 (N_4391,In_478,In_101);
nand U4392 (N_4392,In_684,In_555);
nor U4393 (N_4393,In_874,In_951);
nor U4394 (N_4394,In_250,In_64);
or U4395 (N_4395,In_368,In_361);
nand U4396 (N_4396,In_751,In_565);
nor U4397 (N_4397,In_251,In_832);
and U4398 (N_4398,In_932,In_275);
nand U4399 (N_4399,In_511,In_451);
and U4400 (N_4400,In_143,In_88);
nor U4401 (N_4401,In_730,In_958);
or U4402 (N_4402,In_34,In_265);
and U4403 (N_4403,In_327,In_0);
or U4404 (N_4404,In_109,In_509);
and U4405 (N_4405,In_681,In_486);
nand U4406 (N_4406,In_957,In_913);
and U4407 (N_4407,In_48,In_883);
nor U4408 (N_4408,In_844,In_261);
nor U4409 (N_4409,In_456,In_596);
nor U4410 (N_4410,In_727,In_428);
and U4411 (N_4411,In_742,In_47);
nand U4412 (N_4412,In_118,In_84);
nand U4413 (N_4413,In_236,In_755);
and U4414 (N_4414,In_849,In_58);
and U4415 (N_4415,In_499,In_307);
and U4416 (N_4416,In_34,In_24);
nor U4417 (N_4417,In_650,In_852);
nand U4418 (N_4418,In_753,In_409);
or U4419 (N_4419,In_519,In_639);
nand U4420 (N_4420,In_232,In_23);
or U4421 (N_4421,In_417,In_207);
or U4422 (N_4422,In_155,In_686);
and U4423 (N_4423,In_751,In_596);
or U4424 (N_4424,In_353,In_867);
or U4425 (N_4425,In_742,In_805);
or U4426 (N_4426,In_773,In_820);
nand U4427 (N_4427,In_299,In_787);
nor U4428 (N_4428,In_346,In_166);
nand U4429 (N_4429,In_459,In_268);
nand U4430 (N_4430,In_703,In_97);
or U4431 (N_4431,In_730,In_213);
or U4432 (N_4432,In_99,In_181);
nor U4433 (N_4433,In_277,In_51);
nor U4434 (N_4434,In_123,In_728);
and U4435 (N_4435,In_833,In_248);
and U4436 (N_4436,In_925,In_639);
and U4437 (N_4437,In_531,In_836);
and U4438 (N_4438,In_826,In_924);
nor U4439 (N_4439,In_813,In_548);
and U4440 (N_4440,In_535,In_88);
nor U4441 (N_4441,In_376,In_477);
nand U4442 (N_4442,In_131,In_883);
and U4443 (N_4443,In_731,In_807);
nand U4444 (N_4444,In_90,In_395);
nand U4445 (N_4445,In_891,In_180);
nand U4446 (N_4446,In_643,In_895);
nor U4447 (N_4447,In_852,In_333);
and U4448 (N_4448,In_270,In_353);
nand U4449 (N_4449,In_799,In_746);
or U4450 (N_4450,In_789,In_792);
nand U4451 (N_4451,In_484,In_892);
nor U4452 (N_4452,In_366,In_505);
or U4453 (N_4453,In_588,In_176);
and U4454 (N_4454,In_439,In_780);
nor U4455 (N_4455,In_183,In_798);
and U4456 (N_4456,In_850,In_754);
nor U4457 (N_4457,In_129,In_800);
nand U4458 (N_4458,In_706,In_881);
nor U4459 (N_4459,In_373,In_578);
nand U4460 (N_4460,In_71,In_319);
xor U4461 (N_4461,In_34,In_281);
xor U4462 (N_4462,In_802,In_73);
or U4463 (N_4463,In_45,In_453);
nor U4464 (N_4464,In_314,In_428);
and U4465 (N_4465,In_412,In_784);
xnor U4466 (N_4466,In_617,In_510);
and U4467 (N_4467,In_259,In_991);
and U4468 (N_4468,In_661,In_125);
or U4469 (N_4469,In_329,In_894);
or U4470 (N_4470,In_138,In_34);
and U4471 (N_4471,In_81,In_293);
nand U4472 (N_4472,In_374,In_435);
nor U4473 (N_4473,In_332,In_949);
or U4474 (N_4474,In_264,In_3);
xor U4475 (N_4475,In_369,In_639);
and U4476 (N_4476,In_189,In_115);
nand U4477 (N_4477,In_67,In_289);
nor U4478 (N_4478,In_410,In_310);
or U4479 (N_4479,In_6,In_208);
nor U4480 (N_4480,In_54,In_378);
nand U4481 (N_4481,In_744,In_867);
nor U4482 (N_4482,In_729,In_713);
nor U4483 (N_4483,In_416,In_750);
or U4484 (N_4484,In_948,In_879);
xnor U4485 (N_4485,In_875,In_840);
nand U4486 (N_4486,In_882,In_236);
and U4487 (N_4487,In_749,In_595);
nor U4488 (N_4488,In_546,In_238);
nand U4489 (N_4489,In_347,In_391);
and U4490 (N_4490,In_670,In_110);
and U4491 (N_4491,In_841,In_816);
or U4492 (N_4492,In_890,In_967);
nor U4493 (N_4493,In_760,In_827);
or U4494 (N_4494,In_283,In_931);
nand U4495 (N_4495,In_127,In_178);
or U4496 (N_4496,In_495,In_209);
and U4497 (N_4497,In_225,In_115);
nand U4498 (N_4498,In_953,In_995);
or U4499 (N_4499,In_864,In_565);
and U4500 (N_4500,In_102,In_822);
or U4501 (N_4501,In_447,In_54);
nor U4502 (N_4502,In_703,In_105);
nand U4503 (N_4503,In_62,In_282);
and U4504 (N_4504,In_900,In_895);
nand U4505 (N_4505,In_394,In_646);
nor U4506 (N_4506,In_968,In_984);
and U4507 (N_4507,In_309,In_363);
or U4508 (N_4508,In_438,In_387);
xnor U4509 (N_4509,In_680,In_707);
nor U4510 (N_4510,In_693,In_363);
or U4511 (N_4511,In_359,In_934);
and U4512 (N_4512,In_539,In_294);
and U4513 (N_4513,In_847,In_201);
and U4514 (N_4514,In_357,In_670);
nor U4515 (N_4515,In_801,In_310);
or U4516 (N_4516,In_135,In_714);
nor U4517 (N_4517,In_265,In_709);
nand U4518 (N_4518,In_889,In_961);
or U4519 (N_4519,In_958,In_116);
nand U4520 (N_4520,In_110,In_691);
nor U4521 (N_4521,In_40,In_231);
and U4522 (N_4522,In_903,In_991);
or U4523 (N_4523,In_110,In_893);
and U4524 (N_4524,In_590,In_978);
nand U4525 (N_4525,In_538,In_694);
nor U4526 (N_4526,In_764,In_499);
nand U4527 (N_4527,In_579,In_723);
or U4528 (N_4528,In_96,In_29);
nor U4529 (N_4529,In_450,In_470);
and U4530 (N_4530,In_978,In_951);
or U4531 (N_4531,In_35,In_798);
nand U4532 (N_4532,In_547,In_767);
or U4533 (N_4533,In_347,In_862);
and U4534 (N_4534,In_811,In_515);
nor U4535 (N_4535,In_109,In_827);
or U4536 (N_4536,In_12,In_724);
nand U4537 (N_4537,In_444,In_939);
or U4538 (N_4538,In_351,In_866);
nor U4539 (N_4539,In_303,In_293);
nand U4540 (N_4540,In_761,In_383);
nand U4541 (N_4541,In_758,In_617);
nor U4542 (N_4542,In_300,In_950);
or U4543 (N_4543,In_130,In_696);
and U4544 (N_4544,In_578,In_902);
nand U4545 (N_4545,In_235,In_701);
nand U4546 (N_4546,In_675,In_781);
nand U4547 (N_4547,In_595,In_693);
and U4548 (N_4548,In_492,In_431);
nor U4549 (N_4549,In_156,In_229);
or U4550 (N_4550,In_953,In_801);
xor U4551 (N_4551,In_361,In_709);
nand U4552 (N_4552,In_208,In_581);
nand U4553 (N_4553,In_211,In_456);
nor U4554 (N_4554,In_830,In_822);
nor U4555 (N_4555,In_612,In_375);
or U4556 (N_4556,In_789,In_838);
nand U4557 (N_4557,In_462,In_152);
or U4558 (N_4558,In_301,In_931);
nor U4559 (N_4559,In_867,In_903);
and U4560 (N_4560,In_509,In_48);
and U4561 (N_4561,In_948,In_913);
xor U4562 (N_4562,In_879,In_289);
nor U4563 (N_4563,In_75,In_967);
nor U4564 (N_4564,In_516,In_824);
nor U4565 (N_4565,In_363,In_532);
or U4566 (N_4566,In_807,In_464);
nor U4567 (N_4567,In_366,In_715);
and U4568 (N_4568,In_535,In_906);
and U4569 (N_4569,In_752,In_785);
or U4570 (N_4570,In_964,In_34);
or U4571 (N_4571,In_320,In_187);
nand U4572 (N_4572,In_832,In_736);
nand U4573 (N_4573,In_256,In_425);
or U4574 (N_4574,In_392,In_133);
and U4575 (N_4575,In_677,In_553);
nand U4576 (N_4576,In_174,In_320);
and U4577 (N_4577,In_99,In_409);
and U4578 (N_4578,In_997,In_117);
or U4579 (N_4579,In_865,In_384);
or U4580 (N_4580,In_807,In_697);
or U4581 (N_4581,In_216,In_87);
nor U4582 (N_4582,In_589,In_344);
and U4583 (N_4583,In_868,In_220);
and U4584 (N_4584,In_585,In_663);
nand U4585 (N_4585,In_111,In_257);
and U4586 (N_4586,In_310,In_961);
or U4587 (N_4587,In_308,In_454);
or U4588 (N_4588,In_165,In_310);
or U4589 (N_4589,In_501,In_624);
and U4590 (N_4590,In_766,In_398);
nor U4591 (N_4591,In_738,In_653);
and U4592 (N_4592,In_750,In_476);
nand U4593 (N_4593,In_478,In_916);
and U4594 (N_4594,In_848,In_204);
and U4595 (N_4595,In_299,In_771);
nor U4596 (N_4596,In_688,In_413);
and U4597 (N_4597,In_477,In_793);
or U4598 (N_4598,In_980,In_870);
and U4599 (N_4599,In_988,In_420);
and U4600 (N_4600,In_533,In_191);
nand U4601 (N_4601,In_427,In_296);
or U4602 (N_4602,In_603,In_440);
nor U4603 (N_4603,In_125,In_194);
nand U4604 (N_4604,In_169,In_653);
nor U4605 (N_4605,In_43,In_680);
nand U4606 (N_4606,In_260,In_864);
xor U4607 (N_4607,In_197,In_875);
xnor U4608 (N_4608,In_778,In_528);
nor U4609 (N_4609,In_353,In_768);
or U4610 (N_4610,In_395,In_836);
or U4611 (N_4611,In_897,In_325);
nand U4612 (N_4612,In_624,In_550);
nand U4613 (N_4613,In_263,In_154);
and U4614 (N_4614,In_944,In_749);
nand U4615 (N_4615,In_425,In_956);
nor U4616 (N_4616,In_714,In_159);
nand U4617 (N_4617,In_309,In_236);
and U4618 (N_4618,In_136,In_682);
nor U4619 (N_4619,In_562,In_696);
or U4620 (N_4620,In_970,In_410);
nand U4621 (N_4621,In_571,In_131);
nand U4622 (N_4622,In_697,In_425);
nand U4623 (N_4623,In_902,In_261);
or U4624 (N_4624,In_13,In_836);
nor U4625 (N_4625,In_633,In_383);
and U4626 (N_4626,In_474,In_320);
and U4627 (N_4627,In_925,In_49);
and U4628 (N_4628,In_25,In_63);
and U4629 (N_4629,In_402,In_96);
nand U4630 (N_4630,In_713,In_862);
and U4631 (N_4631,In_896,In_245);
nand U4632 (N_4632,In_970,In_552);
and U4633 (N_4633,In_493,In_881);
and U4634 (N_4634,In_297,In_35);
or U4635 (N_4635,In_550,In_740);
and U4636 (N_4636,In_560,In_576);
nor U4637 (N_4637,In_897,In_671);
nor U4638 (N_4638,In_20,In_820);
or U4639 (N_4639,In_645,In_14);
nor U4640 (N_4640,In_757,In_317);
nand U4641 (N_4641,In_681,In_611);
nand U4642 (N_4642,In_774,In_661);
nor U4643 (N_4643,In_405,In_453);
and U4644 (N_4644,In_942,In_637);
nand U4645 (N_4645,In_978,In_132);
or U4646 (N_4646,In_329,In_734);
nor U4647 (N_4647,In_337,In_46);
or U4648 (N_4648,In_735,In_628);
and U4649 (N_4649,In_899,In_671);
nor U4650 (N_4650,In_559,In_470);
nor U4651 (N_4651,In_485,In_75);
nand U4652 (N_4652,In_61,In_721);
nand U4653 (N_4653,In_666,In_314);
nand U4654 (N_4654,In_834,In_837);
nor U4655 (N_4655,In_123,In_270);
and U4656 (N_4656,In_329,In_972);
and U4657 (N_4657,In_853,In_416);
or U4658 (N_4658,In_878,In_898);
or U4659 (N_4659,In_648,In_672);
or U4660 (N_4660,In_175,In_830);
or U4661 (N_4661,In_168,In_48);
nor U4662 (N_4662,In_112,In_349);
or U4663 (N_4663,In_863,In_521);
nand U4664 (N_4664,In_691,In_606);
and U4665 (N_4665,In_518,In_425);
or U4666 (N_4666,In_953,In_952);
and U4667 (N_4667,In_343,In_216);
nand U4668 (N_4668,In_97,In_417);
or U4669 (N_4669,In_858,In_869);
nand U4670 (N_4670,In_408,In_359);
nor U4671 (N_4671,In_890,In_947);
or U4672 (N_4672,In_585,In_701);
nand U4673 (N_4673,In_85,In_668);
nand U4674 (N_4674,In_701,In_905);
and U4675 (N_4675,In_581,In_341);
nand U4676 (N_4676,In_748,In_379);
and U4677 (N_4677,In_524,In_704);
and U4678 (N_4678,In_99,In_928);
nor U4679 (N_4679,In_0,In_950);
or U4680 (N_4680,In_288,In_710);
nand U4681 (N_4681,In_718,In_489);
nor U4682 (N_4682,In_935,In_593);
or U4683 (N_4683,In_189,In_154);
nand U4684 (N_4684,In_430,In_182);
and U4685 (N_4685,In_692,In_10);
and U4686 (N_4686,In_246,In_374);
nor U4687 (N_4687,In_226,In_217);
and U4688 (N_4688,In_336,In_901);
and U4689 (N_4689,In_686,In_945);
nand U4690 (N_4690,In_580,In_256);
and U4691 (N_4691,In_632,In_504);
or U4692 (N_4692,In_395,In_123);
or U4693 (N_4693,In_451,In_430);
nor U4694 (N_4694,In_559,In_292);
nand U4695 (N_4695,In_807,In_69);
and U4696 (N_4696,In_521,In_828);
nor U4697 (N_4697,In_706,In_585);
nand U4698 (N_4698,In_983,In_817);
and U4699 (N_4699,In_934,In_907);
and U4700 (N_4700,In_668,In_197);
nand U4701 (N_4701,In_941,In_400);
nand U4702 (N_4702,In_719,In_93);
nor U4703 (N_4703,In_744,In_889);
nand U4704 (N_4704,In_951,In_66);
nor U4705 (N_4705,In_217,In_801);
or U4706 (N_4706,In_257,In_828);
and U4707 (N_4707,In_809,In_197);
or U4708 (N_4708,In_952,In_756);
xnor U4709 (N_4709,In_472,In_806);
and U4710 (N_4710,In_985,In_663);
or U4711 (N_4711,In_832,In_695);
or U4712 (N_4712,In_476,In_990);
and U4713 (N_4713,In_2,In_611);
nand U4714 (N_4714,In_29,In_836);
nor U4715 (N_4715,In_911,In_250);
nand U4716 (N_4716,In_664,In_212);
and U4717 (N_4717,In_726,In_515);
or U4718 (N_4718,In_520,In_562);
or U4719 (N_4719,In_676,In_967);
nand U4720 (N_4720,In_782,In_562);
nand U4721 (N_4721,In_968,In_986);
or U4722 (N_4722,In_248,In_401);
nand U4723 (N_4723,In_655,In_825);
nor U4724 (N_4724,In_929,In_191);
nand U4725 (N_4725,In_862,In_595);
and U4726 (N_4726,In_99,In_464);
or U4727 (N_4727,In_694,In_409);
xnor U4728 (N_4728,In_558,In_121);
nand U4729 (N_4729,In_992,In_884);
nand U4730 (N_4730,In_247,In_769);
nand U4731 (N_4731,In_390,In_61);
or U4732 (N_4732,In_317,In_494);
nor U4733 (N_4733,In_168,In_502);
nor U4734 (N_4734,In_64,In_0);
and U4735 (N_4735,In_4,In_483);
nor U4736 (N_4736,In_320,In_759);
nor U4737 (N_4737,In_207,In_611);
xor U4738 (N_4738,In_141,In_294);
nand U4739 (N_4739,In_50,In_298);
and U4740 (N_4740,In_80,In_701);
or U4741 (N_4741,In_51,In_504);
and U4742 (N_4742,In_94,In_84);
nor U4743 (N_4743,In_2,In_53);
and U4744 (N_4744,In_691,In_563);
or U4745 (N_4745,In_938,In_641);
or U4746 (N_4746,In_957,In_266);
nand U4747 (N_4747,In_50,In_446);
nor U4748 (N_4748,In_359,In_491);
or U4749 (N_4749,In_483,In_782);
nor U4750 (N_4750,In_148,In_580);
or U4751 (N_4751,In_124,In_160);
and U4752 (N_4752,In_241,In_978);
and U4753 (N_4753,In_909,In_887);
and U4754 (N_4754,In_852,In_976);
nand U4755 (N_4755,In_788,In_225);
nor U4756 (N_4756,In_485,In_153);
nand U4757 (N_4757,In_516,In_867);
and U4758 (N_4758,In_439,In_893);
nand U4759 (N_4759,In_973,In_138);
nand U4760 (N_4760,In_208,In_99);
xor U4761 (N_4761,In_902,In_426);
and U4762 (N_4762,In_192,In_847);
or U4763 (N_4763,In_470,In_616);
nand U4764 (N_4764,In_810,In_108);
and U4765 (N_4765,In_349,In_994);
or U4766 (N_4766,In_849,In_714);
nor U4767 (N_4767,In_232,In_481);
nand U4768 (N_4768,In_578,In_18);
xnor U4769 (N_4769,In_326,In_856);
and U4770 (N_4770,In_469,In_204);
or U4771 (N_4771,In_574,In_421);
nand U4772 (N_4772,In_558,In_830);
nor U4773 (N_4773,In_96,In_283);
nand U4774 (N_4774,In_647,In_411);
nand U4775 (N_4775,In_319,In_954);
nand U4776 (N_4776,In_673,In_185);
nor U4777 (N_4777,In_427,In_80);
or U4778 (N_4778,In_659,In_654);
nor U4779 (N_4779,In_948,In_828);
and U4780 (N_4780,In_963,In_697);
or U4781 (N_4781,In_890,In_572);
nor U4782 (N_4782,In_937,In_809);
nand U4783 (N_4783,In_328,In_663);
or U4784 (N_4784,In_928,In_217);
nand U4785 (N_4785,In_796,In_881);
nor U4786 (N_4786,In_732,In_815);
and U4787 (N_4787,In_345,In_955);
nor U4788 (N_4788,In_564,In_690);
and U4789 (N_4789,In_591,In_225);
nand U4790 (N_4790,In_396,In_186);
and U4791 (N_4791,In_845,In_741);
nand U4792 (N_4792,In_738,In_985);
nor U4793 (N_4793,In_530,In_140);
and U4794 (N_4794,In_416,In_438);
and U4795 (N_4795,In_957,In_70);
or U4796 (N_4796,In_384,In_443);
nor U4797 (N_4797,In_739,In_919);
nand U4798 (N_4798,In_297,In_409);
and U4799 (N_4799,In_45,In_324);
xor U4800 (N_4800,In_292,In_793);
or U4801 (N_4801,In_605,In_525);
and U4802 (N_4802,In_918,In_220);
nor U4803 (N_4803,In_661,In_534);
and U4804 (N_4804,In_101,In_473);
or U4805 (N_4805,In_392,In_853);
xnor U4806 (N_4806,In_995,In_117);
or U4807 (N_4807,In_193,In_680);
nand U4808 (N_4808,In_787,In_744);
or U4809 (N_4809,In_518,In_885);
and U4810 (N_4810,In_446,In_566);
or U4811 (N_4811,In_595,In_855);
nor U4812 (N_4812,In_446,In_265);
and U4813 (N_4813,In_454,In_971);
or U4814 (N_4814,In_357,In_788);
or U4815 (N_4815,In_399,In_324);
nand U4816 (N_4816,In_791,In_433);
or U4817 (N_4817,In_87,In_215);
nor U4818 (N_4818,In_474,In_382);
or U4819 (N_4819,In_252,In_180);
xnor U4820 (N_4820,In_910,In_852);
nor U4821 (N_4821,In_71,In_91);
or U4822 (N_4822,In_563,In_756);
and U4823 (N_4823,In_783,In_588);
and U4824 (N_4824,In_595,In_946);
or U4825 (N_4825,In_59,In_985);
and U4826 (N_4826,In_158,In_704);
or U4827 (N_4827,In_751,In_664);
nor U4828 (N_4828,In_909,In_658);
nor U4829 (N_4829,In_369,In_422);
nand U4830 (N_4830,In_342,In_283);
nand U4831 (N_4831,In_643,In_930);
nor U4832 (N_4832,In_107,In_314);
or U4833 (N_4833,In_999,In_539);
nor U4834 (N_4834,In_504,In_316);
or U4835 (N_4835,In_589,In_112);
or U4836 (N_4836,In_133,In_440);
or U4837 (N_4837,In_564,In_339);
and U4838 (N_4838,In_867,In_334);
or U4839 (N_4839,In_673,In_131);
and U4840 (N_4840,In_431,In_928);
nand U4841 (N_4841,In_229,In_380);
nand U4842 (N_4842,In_930,In_693);
or U4843 (N_4843,In_702,In_13);
xor U4844 (N_4844,In_129,In_284);
nand U4845 (N_4845,In_143,In_532);
or U4846 (N_4846,In_75,In_962);
and U4847 (N_4847,In_19,In_658);
or U4848 (N_4848,In_245,In_494);
or U4849 (N_4849,In_386,In_853);
or U4850 (N_4850,In_624,In_386);
or U4851 (N_4851,In_36,In_318);
and U4852 (N_4852,In_389,In_677);
and U4853 (N_4853,In_888,In_47);
nor U4854 (N_4854,In_271,In_16);
nor U4855 (N_4855,In_305,In_106);
or U4856 (N_4856,In_584,In_231);
or U4857 (N_4857,In_83,In_289);
xnor U4858 (N_4858,In_794,In_817);
or U4859 (N_4859,In_777,In_767);
xor U4860 (N_4860,In_981,In_429);
or U4861 (N_4861,In_925,In_672);
nor U4862 (N_4862,In_753,In_807);
and U4863 (N_4863,In_166,In_827);
nor U4864 (N_4864,In_822,In_888);
nor U4865 (N_4865,In_300,In_847);
or U4866 (N_4866,In_420,In_349);
nand U4867 (N_4867,In_637,In_649);
nand U4868 (N_4868,In_514,In_227);
nor U4869 (N_4869,In_932,In_578);
and U4870 (N_4870,In_149,In_404);
and U4871 (N_4871,In_69,In_361);
nor U4872 (N_4872,In_205,In_60);
or U4873 (N_4873,In_411,In_415);
nand U4874 (N_4874,In_108,In_583);
or U4875 (N_4875,In_39,In_654);
nand U4876 (N_4876,In_87,In_952);
nor U4877 (N_4877,In_9,In_179);
nor U4878 (N_4878,In_138,In_598);
nand U4879 (N_4879,In_20,In_252);
and U4880 (N_4880,In_338,In_332);
or U4881 (N_4881,In_611,In_248);
nor U4882 (N_4882,In_597,In_866);
or U4883 (N_4883,In_297,In_38);
and U4884 (N_4884,In_330,In_854);
nand U4885 (N_4885,In_7,In_642);
or U4886 (N_4886,In_774,In_422);
and U4887 (N_4887,In_166,In_720);
nor U4888 (N_4888,In_667,In_542);
and U4889 (N_4889,In_774,In_979);
xnor U4890 (N_4890,In_432,In_567);
and U4891 (N_4891,In_79,In_215);
and U4892 (N_4892,In_266,In_859);
or U4893 (N_4893,In_109,In_463);
nor U4894 (N_4894,In_756,In_105);
nor U4895 (N_4895,In_519,In_481);
nand U4896 (N_4896,In_909,In_362);
nor U4897 (N_4897,In_293,In_50);
nand U4898 (N_4898,In_97,In_83);
and U4899 (N_4899,In_662,In_574);
nor U4900 (N_4900,In_291,In_264);
or U4901 (N_4901,In_970,In_604);
nor U4902 (N_4902,In_764,In_143);
nand U4903 (N_4903,In_226,In_927);
and U4904 (N_4904,In_288,In_573);
nor U4905 (N_4905,In_752,In_98);
nor U4906 (N_4906,In_894,In_364);
nor U4907 (N_4907,In_12,In_594);
nor U4908 (N_4908,In_701,In_74);
and U4909 (N_4909,In_698,In_31);
nor U4910 (N_4910,In_280,In_391);
or U4911 (N_4911,In_157,In_825);
or U4912 (N_4912,In_172,In_286);
and U4913 (N_4913,In_714,In_260);
nand U4914 (N_4914,In_92,In_244);
nor U4915 (N_4915,In_719,In_118);
or U4916 (N_4916,In_579,In_201);
nand U4917 (N_4917,In_399,In_948);
nand U4918 (N_4918,In_259,In_170);
nand U4919 (N_4919,In_170,In_468);
nor U4920 (N_4920,In_428,In_23);
or U4921 (N_4921,In_60,In_415);
and U4922 (N_4922,In_474,In_861);
or U4923 (N_4923,In_677,In_206);
or U4924 (N_4924,In_917,In_568);
or U4925 (N_4925,In_281,In_127);
xnor U4926 (N_4926,In_849,In_306);
and U4927 (N_4927,In_929,In_985);
and U4928 (N_4928,In_755,In_921);
or U4929 (N_4929,In_195,In_994);
and U4930 (N_4930,In_932,In_756);
nor U4931 (N_4931,In_753,In_689);
xor U4932 (N_4932,In_42,In_859);
nand U4933 (N_4933,In_164,In_551);
or U4934 (N_4934,In_272,In_866);
nor U4935 (N_4935,In_638,In_965);
and U4936 (N_4936,In_131,In_400);
or U4937 (N_4937,In_826,In_543);
nor U4938 (N_4938,In_393,In_852);
xnor U4939 (N_4939,In_143,In_212);
nand U4940 (N_4940,In_228,In_33);
and U4941 (N_4941,In_748,In_241);
nor U4942 (N_4942,In_528,In_954);
or U4943 (N_4943,In_493,In_205);
or U4944 (N_4944,In_606,In_922);
nand U4945 (N_4945,In_94,In_233);
and U4946 (N_4946,In_879,In_346);
nor U4947 (N_4947,In_587,In_193);
nor U4948 (N_4948,In_727,In_842);
nor U4949 (N_4949,In_736,In_38);
and U4950 (N_4950,In_347,In_177);
nand U4951 (N_4951,In_409,In_132);
or U4952 (N_4952,In_792,In_302);
nand U4953 (N_4953,In_485,In_607);
and U4954 (N_4954,In_767,In_941);
or U4955 (N_4955,In_515,In_85);
and U4956 (N_4956,In_581,In_101);
nor U4957 (N_4957,In_505,In_578);
and U4958 (N_4958,In_780,In_483);
and U4959 (N_4959,In_248,In_862);
or U4960 (N_4960,In_266,In_273);
nor U4961 (N_4961,In_54,In_37);
nand U4962 (N_4962,In_216,In_498);
nand U4963 (N_4963,In_905,In_326);
or U4964 (N_4964,In_530,In_586);
and U4965 (N_4965,In_776,In_3);
and U4966 (N_4966,In_488,In_343);
or U4967 (N_4967,In_368,In_30);
or U4968 (N_4968,In_159,In_269);
or U4969 (N_4969,In_595,In_348);
nor U4970 (N_4970,In_848,In_600);
and U4971 (N_4971,In_990,In_258);
and U4972 (N_4972,In_673,In_588);
and U4973 (N_4973,In_87,In_120);
or U4974 (N_4974,In_117,In_250);
or U4975 (N_4975,In_836,In_178);
nand U4976 (N_4976,In_977,In_626);
or U4977 (N_4977,In_537,In_329);
nor U4978 (N_4978,In_643,In_722);
and U4979 (N_4979,In_375,In_552);
nor U4980 (N_4980,In_956,In_74);
or U4981 (N_4981,In_116,In_971);
or U4982 (N_4982,In_439,In_367);
nor U4983 (N_4983,In_225,In_957);
and U4984 (N_4984,In_103,In_675);
nand U4985 (N_4985,In_6,In_60);
nand U4986 (N_4986,In_270,In_862);
and U4987 (N_4987,In_784,In_282);
or U4988 (N_4988,In_810,In_622);
nor U4989 (N_4989,In_665,In_406);
or U4990 (N_4990,In_792,In_602);
and U4991 (N_4991,In_829,In_369);
or U4992 (N_4992,In_499,In_52);
nor U4993 (N_4993,In_788,In_194);
nand U4994 (N_4994,In_961,In_119);
nand U4995 (N_4995,In_482,In_944);
nand U4996 (N_4996,In_700,In_698);
nand U4997 (N_4997,In_683,In_365);
nand U4998 (N_4998,In_88,In_742);
or U4999 (N_4999,In_243,In_625);
nor U5000 (N_5000,N_1310,N_2989);
nand U5001 (N_5001,N_3964,N_4678);
nor U5002 (N_5002,N_4673,N_51);
nor U5003 (N_5003,N_2536,N_3573);
nor U5004 (N_5004,N_907,N_1304);
and U5005 (N_5005,N_3762,N_2062);
or U5006 (N_5006,N_4768,N_3831);
nand U5007 (N_5007,N_2142,N_3871);
nor U5008 (N_5008,N_4272,N_3424);
nand U5009 (N_5009,N_3583,N_1130);
or U5010 (N_5010,N_2171,N_969);
nand U5011 (N_5011,N_3621,N_835);
and U5012 (N_5012,N_2321,N_3225);
nor U5013 (N_5013,N_1690,N_1461);
and U5014 (N_5014,N_4130,N_1290);
or U5015 (N_5015,N_478,N_4201);
and U5016 (N_5016,N_961,N_742);
nand U5017 (N_5017,N_2364,N_4065);
and U5018 (N_5018,N_3833,N_2825);
and U5019 (N_5019,N_3343,N_1893);
and U5020 (N_5020,N_1256,N_343);
xor U5021 (N_5021,N_2465,N_3847);
nand U5022 (N_5022,N_2766,N_3646);
nor U5023 (N_5023,N_4661,N_934);
nor U5024 (N_5024,N_3035,N_3332);
and U5025 (N_5025,N_4615,N_4927);
nor U5026 (N_5026,N_4829,N_121);
nor U5027 (N_5027,N_931,N_2813);
nor U5028 (N_5028,N_3023,N_1020);
or U5029 (N_5029,N_4077,N_167);
nand U5030 (N_5030,N_4142,N_4102);
xor U5031 (N_5031,N_4915,N_194);
nand U5032 (N_5032,N_3290,N_295);
nand U5033 (N_5033,N_999,N_1727);
and U5034 (N_5034,N_4220,N_1540);
or U5035 (N_5035,N_1433,N_373);
and U5036 (N_5036,N_1875,N_1435);
xnor U5037 (N_5037,N_159,N_4838);
nand U5038 (N_5038,N_834,N_1505);
nand U5039 (N_5039,N_3369,N_3641);
nand U5040 (N_5040,N_530,N_1728);
and U5041 (N_5041,N_1264,N_738);
and U5042 (N_5042,N_1914,N_1792);
or U5043 (N_5043,N_4252,N_2925);
or U5044 (N_5044,N_599,N_3920);
nand U5045 (N_5045,N_2937,N_2230);
nor U5046 (N_5046,N_1923,N_1880);
nor U5047 (N_5047,N_3510,N_3466);
and U5048 (N_5048,N_4264,N_2201);
and U5049 (N_5049,N_4479,N_785);
and U5050 (N_5050,N_862,N_2840);
nand U5051 (N_5051,N_3313,N_1267);
nor U5052 (N_5052,N_891,N_118);
nor U5053 (N_5053,N_2674,N_828);
or U5054 (N_5054,N_2819,N_3031);
or U5055 (N_5055,N_4742,N_1819);
or U5056 (N_5056,N_780,N_2558);
or U5057 (N_5057,N_1037,N_4056);
or U5058 (N_5058,N_4262,N_4613);
xnor U5059 (N_5059,N_1682,N_2810);
nor U5060 (N_5060,N_2186,N_3653);
nor U5061 (N_5061,N_3101,N_1558);
nand U5062 (N_5062,N_4800,N_4402);
nor U5063 (N_5063,N_60,N_3296);
or U5064 (N_5064,N_4752,N_3073);
nor U5065 (N_5065,N_4563,N_2385);
and U5066 (N_5066,N_2426,N_4680);
or U5067 (N_5067,N_4235,N_1824);
nor U5068 (N_5068,N_2758,N_1467);
nor U5069 (N_5069,N_213,N_1543);
xor U5070 (N_5070,N_2804,N_3188);
nand U5071 (N_5071,N_157,N_2777);
and U5072 (N_5072,N_2362,N_4633);
or U5073 (N_5073,N_3973,N_1634);
nor U5074 (N_5074,N_864,N_611);
and U5075 (N_5075,N_921,N_4277);
nand U5076 (N_5076,N_318,N_1647);
or U5077 (N_5077,N_2635,N_1254);
nand U5078 (N_5078,N_4575,N_116);
and U5079 (N_5079,N_4675,N_1485);
nor U5080 (N_5080,N_3544,N_3324);
or U5081 (N_5081,N_2651,N_4648);
nor U5082 (N_5082,N_2018,N_4331);
and U5083 (N_5083,N_1090,N_2311);
nand U5084 (N_5084,N_1599,N_3231);
nand U5085 (N_5085,N_1570,N_3375);
and U5086 (N_5086,N_4592,N_4221);
and U5087 (N_5087,N_2907,N_4336);
nor U5088 (N_5088,N_3816,N_3988);
nand U5089 (N_5089,N_4516,N_4093);
and U5090 (N_5090,N_3880,N_1076);
nor U5091 (N_5091,N_1409,N_1906);
nor U5092 (N_5092,N_4072,N_3044);
nand U5093 (N_5093,N_384,N_1743);
and U5094 (N_5094,N_4112,N_655);
and U5095 (N_5095,N_2908,N_4285);
and U5096 (N_5096,N_811,N_1896);
and U5097 (N_5097,N_2210,N_2286);
nand U5098 (N_5098,N_3608,N_1741);
or U5099 (N_5099,N_4907,N_620);
nor U5100 (N_5100,N_2643,N_2007);
or U5101 (N_5101,N_1432,N_1444);
and U5102 (N_5102,N_3901,N_2931);
and U5103 (N_5103,N_2887,N_3);
and U5104 (N_5104,N_3148,N_4750);
and U5105 (N_5105,N_2541,N_2435);
and U5106 (N_5106,N_4154,N_3948);
or U5107 (N_5107,N_518,N_2271);
or U5108 (N_5108,N_4952,N_3215);
or U5109 (N_5109,N_2607,N_1989);
and U5110 (N_5110,N_1268,N_2519);
and U5111 (N_5111,N_3700,N_494);
nand U5112 (N_5112,N_1152,N_3884);
nor U5113 (N_5113,N_733,N_1036);
nor U5114 (N_5114,N_512,N_4769);
nand U5115 (N_5115,N_3087,N_3971);
or U5116 (N_5116,N_557,N_382);
xor U5117 (N_5117,N_1587,N_2064);
nor U5118 (N_5118,N_2670,N_1063);
and U5119 (N_5119,N_714,N_2055);
xnor U5120 (N_5120,N_4208,N_4271);
nor U5121 (N_5121,N_3584,N_3434);
nand U5122 (N_5122,N_4055,N_2707);
nor U5123 (N_5123,N_3407,N_4215);
and U5124 (N_5124,N_2748,N_4367);
and U5125 (N_5125,N_686,N_1207);
or U5126 (N_5126,N_4568,N_3850);
nand U5127 (N_5127,N_1289,N_2730);
nand U5128 (N_5128,N_1422,N_764);
and U5129 (N_5129,N_1248,N_2097);
nand U5130 (N_5130,N_3160,N_161);
or U5131 (N_5131,N_560,N_2653);
or U5132 (N_5132,N_4760,N_2481);
and U5133 (N_5133,N_207,N_3076);
xor U5134 (N_5134,N_3502,N_508);
and U5135 (N_5135,N_2543,N_452);
and U5136 (N_5136,N_1426,N_3553);
nor U5137 (N_5137,N_4260,N_3380);
nand U5138 (N_5138,N_1837,N_301);
nor U5139 (N_5139,N_3534,N_2951);
or U5140 (N_5140,N_4749,N_4978);
nor U5141 (N_5141,N_643,N_3356);
nor U5142 (N_5142,N_4969,N_2767);
or U5143 (N_5143,N_2875,N_4033);
nand U5144 (N_5144,N_3515,N_1628);
or U5145 (N_5145,N_4510,N_438);
and U5146 (N_5146,N_2837,N_1338);
nand U5147 (N_5147,N_3066,N_1892);
nor U5148 (N_5148,N_4804,N_4273);
nand U5149 (N_5149,N_323,N_3269);
and U5150 (N_5150,N_2127,N_1501);
or U5151 (N_5151,N_2559,N_3654);
and U5152 (N_5152,N_713,N_4270);
nand U5153 (N_5153,N_408,N_4945);
nor U5154 (N_5154,N_898,N_2282);
and U5155 (N_5155,N_1815,N_805);
and U5156 (N_5156,N_4544,N_2665);
nand U5157 (N_5157,N_2520,N_3385);
and U5158 (N_5158,N_2374,N_3648);
and U5159 (N_5159,N_289,N_3602);
nand U5160 (N_5160,N_1303,N_715);
or U5161 (N_5161,N_3048,N_3582);
nand U5162 (N_5162,N_2329,N_757);
and U5163 (N_5163,N_2068,N_196);
nor U5164 (N_5164,N_1738,N_3259);
nor U5165 (N_5165,N_423,N_2721);
or U5166 (N_5166,N_1613,N_2704);
and U5167 (N_5167,N_2081,N_3720);
xor U5168 (N_5168,N_4667,N_4013);
nand U5169 (N_5169,N_3824,N_726);
or U5170 (N_5170,N_303,N_4160);
nor U5171 (N_5171,N_2043,N_3123);
or U5172 (N_5172,N_2262,N_519);
nand U5173 (N_5173,N_888,N_4627);
nand U5174 (N_5174,N_625,N_4481);
nor U5175 (N_5175,N_1410,N_4288);
or U5176 (N_5176,N_4015,N_4038);
and U5177 (N_5177,N_1689,N_4526);
and U5178 (N_5178,N_2560,N_4135);
nor U5179 (N_5179,N_1523,N_4036);
and U5180 (N_5180,N_3368,N_3491);
nor U5181 (N_5181,N_1598,N_76);
nand U5182 (N_5182,N_340,N_4014);
or U5183 (N_5183,N_4407,N_2410);
or U5184 (N_5184,N_2727,N_3861);
and U5185 (N_5185,N_1292,N_1360);
and U5186 (N_5186,N_38,N_3704);
nand U5187 (N_5187,N_216,N_3374);
and U5188 (N_5188,N_3522,N_4751);
nand U5189 (N_5189,N_903,N_3206);
and U5190 (N_5190,N_3435,N_1380);
and U5191 (N_5191,N_1226,N_1873);
nand U5192 (N_5192,N_3624,N_265);
nand U5193 (N_5193,N_2178,N_3392);
or U5194 (N_5194,N_4095,N_2679);
or U5195 (N_5195,N_3308,N_1677);
nand U5196 (N_5196,N_503,N_1631);
nand U5197 (N_5197,N_1674,N_618);
or U5198 (N_5198,N_4736,N_278);
nor U5199 (N_5199,N_2854,N_4898);
nand U5200 (N_5200,N_4097,N_4929);
and U5201 (N_5201,N_2188,N_2156);
nand U5202 (N_5202,N_4576,N_4618);
and U5203 (N_5203,N_4641,N_4798);
or U5204 (N_5204,N_2216,N_2408);
and U5205 (N_5205,N_2921,N_3154);
and U5206 (N_5206,N_4146,N_4194);
nor U5207 (N_5207,N_1367,N_1552);
and U5208 (N_5208,N_4373,N_1032);
xor U5209 (N_5209,N_4333,N_2391);
or U5210 (N_5210,N_3316,N_3086);
and U5211 (N_5211,N_3433,N_150);
and U5212 (N_5212,N_952,N_4424);
nor U5213 (N_5213,N_2054,N_2888);
and U5214 (N_5214,N_4746,N_3490);
and U5215 (N_5215,N_3963,N_4230);
and U5216 (N_5216,N_3543,N_1196);
nor U5217 (N_5217,N_2846,N_4832);
or U5218 (N_5218,N_803,N_4256);
and U5219 (N_5219,N_3987,N_1252);
xor U5220 (N_5220,N_2561,N_2177);
or U5221 (N_5221,N_4921,N_306);
and U5222 (N_5222,N_4983,N_275);
xor U5223 (N_5223,N_4027,N_689);
or U5224 (N_5224,N_3352,N_4885);
nand U5225 (N_5225,N_4420,N_4595);
nand U5226 (N_5226,N_2586,N_460);
or U5227 (N_5227,N_3415,N_3479);
nor U5228 (N_5228,N_3775,N_1178);
or U5229 (N_5229,N_3656,N_2390);
and U5230 (N_5230,N_4995,N_4989);
nor U5231 (N_5231,N_2749,N_1487);
or U5232 (N_5232,N_1723,N_3881);
nor U5233 (N_5233,N_942,N_963);
nor U5234 (N_5234,N_2169,N_4933);
and U5235 (N_5235,N_30,N_2631);
or U5236 (N_5236,N_3939,N_54);
or U5237 (N_5237,N_1155,N_1403);
nor U5238 (N_5238,N_4939,N_2445);
nand U5239 (N_5239,N_4843,N_995);
and U5240 (N_5240,N_2428,N_668);
nor U5241 (N_5241,N_3328,N_2012);
or U5242 (N_5242,N_1132,N_1049);
nor U5243 (N_5243,N_966,N_2089);
and U5244 (N_5244,N_1503,N_4069);
nor U5245 (N_5245,N_3671,N_539);
and U5246 (N_5246,N_2366,N_4934);
or U5247 (N_5247,N_2982,N_3567);
xnor U5248 (N_5248,N_3790,N_3454);
and U5249 (N_5249,N_2056,N_1314);
and U5250 (N_5250,N_4779,N_1162);
nand U5251 (N_5251,N_2058,N_2165);
and U5252 (N_5252,N_3617,N_3683);
or U5253 (N_5253,N_2473,N_1545);
nand U5254 (N_5254,N_1332,N_3756);
or U5255 (N_5255,N_2108,N_1640);
or U5256 (N_5256,N_2330,N_2332);
nand U5257 (N_5257,N_1497,N_1740);
or U5258 (N_5258,N_3868,N_139);
or U5259 (N_5259,N_3451,N_1220);
and U5260 (N_5260,N_2038,N_1583);
or U5261 (N_5261,N_2630,N_4868);
or U5262 (N_5262,N_2745,N_1167);
nor U5263 (N_5263,N_3969,N_3983);
and U5264 (N_5264,N_3933,N_2847);
nand U5265 (N_5265,N_3032,N_1074);
nor U5266 (N_5266,N_2192,N_2673);
or U5267 (N_5267,N_3929,N_964);
or U5268 (N_5268,N_3942,N_3834);
nand U5269 (N_5269,N_145,N_923);
nor U5270 (N_5270,N_4418,N_449);
or U5271 (N_5271,N_4283,N_3242);
and U5272 (N_5272,N_2351,N_2022);
or U5273 (N_5273,N_2028,N_292);
nor U5274 (N_5274,N_2008,N_3972);
nor U5275 (N_5275,N_4651,N_2677);
or U5276 (N_5276,N_4930,N_1786);
or U5277 (N_5277,N_2413,N_3612);
nand U5278 (N_5278,N_506,N_4266);
nand U5279 (N_5279,N_4844,N_4248);
nand U5280 (N_5280,N_1548,N_1542);
and U5281 (N_5281,N_763,N_4274);
and U5282 (N_5282,N_1626,N_2615);
nand U5283 (N_5283,N_1034,N_2961);
or U5284 (N_5284,N_1514,N_3517);
or U5285 (N_5285,N_3472,N_5);
nand U5286 (N_5286,N_511,N_3974);
and U5287 (N_5287,N_481,N_4527);
nand U5288 (N_5288,N_131,N_2689);
or U5289 (N_5289,N_3223,N_2109);
nor U5290 (N_5290,N_4758,N_4801);
nand U5291 (N_5291,N_4532,N_4192);
or U5292 (N_5292,N_917,N_378);
nand U5293 (N_5293,N_1278,N_4891);
nor U5294 (N_5294,N_4708,N_82);
nor U5295 (N_5295,N_3586,N_4845);
and U5296 (N_5296,N_3554,N_3266);
or U5297 (N_5297,N_3114,N_4118);
nand U5298 (N_5298,N_23,N_4179);
nand U5299 (N_5299,N_2452,N_2485);
and U5300 (N_5300,N_4805,N_747);
nor U5301 (N_5301,N_4491,N_4696);
nand U5302 (N_5302,N_4968,N_3357);
or U5303 (N_5303,N_317,N_4133);
or U5304 (N_5304,N_3765,N_826);
or U5305 (N_5305,N_2221,N_420);
xnor U5306 (N_5306,N_3449,N_313);
nand U5307 (N_5307,N_471,N_3864);
nand U5308 (N_5308,N_2244,N_960);
or U5309 (N_5309,N_1428,N_2274);
and U5310 (N_5310,N_4582,N_1646);
nor U5311 (N_5311,N_4383,N_4403);
and U5312 (N_5312,N_1042,N_2952);
nand U5313 (N_5313,N_1495,N_1962);
nor U5314 (N_5314,N_2167,N_2832);
or U5315 (N_5315,N_1698,N_1838);
or U5316 (N_5316,N_3842,N_1616);
nor U5317 (N_5317,N_484,N_1954);
and U5318 (N_5318,N_4190,N_2660);
nor U5319 (N_5319,N_1055,N_3161);
or U5320 (N_5320,N_4021,N_3823);
or U5321 (N_5321,N_205,N_1151);
or U5322 (N_5322,N_4761,N_2479);
nand U5323 (N_5323,N_3755,N_3278);
nor U5324 (N_5324,N_1431,N_3173);
or U5325 (N_5325,N_1714,N_3692);
or U5326 (N_5326,N_2917,N_456);
nand U5327 (N_5327,N_1774,N_2650);
or U5328 (N_5328,N_922,N_4637);
nor U5329 (N_5329,N_2988,N_671);
nand U5330 (N_5330,N_1054,N_1601);
nor U5331 (N_5331,N_4173,N_4175);
and U5332 (N_5332,N_3258,N_526);
xnor U5333 (N_5333,N_2879,N_1607);
nand U5334 (N_5334,N_1011,N_4067);
nor U5335 (N_5335,N_2429,N_2256);
nor U5336 (N_5336,N_2870,N_899);
or U5337 (N_5337,N_1771,N_142);
nor U5338 (N_5338,N_1105,N_1483);
nand U5339 (N_5339,N_1676,N_1203);
and U5340 (N_5340,N_2250,N_2360);
or U5341 (N_5341,N_796,N_4344);
nor U5342 (N_5342,N_3955,N_489);
nor U5343 (N_5343,N_4267,N_439);
and U5344 (N_5344,N_2489,N_4059);
xnor U5345 (N_5345,N_3777,N_2496);
nor U5346 (N_5346,N_1357,N_4622);
nor U5347 (N_5347,N_3229,N_4882);
nor U5348 (N_5348,N_2316,N_3688);
and U5349 (N_5349,N_2335,N_4387);
and U5350 (N_5350,N_462,N_1166);
nand U5351 (N_5351,N_154,N_2269);
nor U5352 (N_5352,N_2593,N_4366);
nand U5353 (N_5353,N_1418,N_1911);
or U5354 (N_5354,N_2273,N_2654);
and U5355 (N_5355,N_3975,N_3622);
and U5356 (N_5356,N_2884,N_4520);
and U5357 (N_5357,N_1293,N_3200);
nor U5358 (N_5358,N_2471,N_4653);
xor U5359 (N_5359,N_4773,N_2310);
and U5360 (N_5360,N_3507,N_972);
and U5361 (N_5361,N_3379,N_4570);
nand U5362 (N_5362,N_2202,N_269);
or U5363 (N_5363,N_4075,N_2579);
and U5364 (N_5364,N_4860,N_2786);
nand U5365 (N_5365,N_381,N_2838);
or U5366 (N_5366,N_1748,N_3458);
or U5367 (N_5367,N_3088,N_1014);
nor U5368 (N_5368,N_1161,N_4376);
nand U5369 (N_5369,N_2499,N_865);
or U5370 (N_5370,N_2009,N_4497);
nand U5371 (N_5371,N_536,N_1029);
and U5372 (N_5372,N_900,N_3321);
nor U5373 (N_5373,N_3124,N_2814);
nor U5374 (N_5374,N_2328,N_3480);
nor U5375 (N_5375,N_2912,N_2432);
nor U5376 (N_5376,N_1135,N_426);
nor U5377 (N_5377,N_848,N_753);
nor U5378 (N_5378,N_756,N_2755);
nor U5379 (N_5379,N_2005,N_3666);
nor U5380 (N_5380,N_2088,N_892);
or U5381 (N_5381,N_957,N_2728);
and U5382 (N_5382,N_4011,N_3572);
xor U5383 (N_5383,N_2708,N_4878);
nand U5384 (N_5384,N_1478,N_1809);
or U5385 (N_5385,N_3542,N_3156);
and U5386 (N_5386,N_4312,N_4370);
nor U5387 (N_5387,N_4743,N_1961);
nor U5388 (N_5388,N_1804,N_2085);
nand U5389 (N_5389,N_3947,N_2011);
and U5390 (N_5390,N_4553,N_3630);
nand U5391 (N_5391,N_2798,N_434);
nor U5392 (N_5392,N_2947,N_1956);
and U5393 (N_5393,N_3960,N_3403);
and U5394 (N_5394,N_2260,N_1159);
nand U5395 (N_5395,N_203,N_1412);
and U5396 (N_5396,N_3506,N_108);
nand U5397 (N_5397,N_1806,N_2079);
nor U5398 (N_5398,N_2304,N_364);
nand U5399 (N_5399,N_3325,N_4797);
and U5400 (N_5400,N_3503,N_745);
or U5401 (N_5401,N_2238,N_1294);
or U5402 (N_5402,N_2641,N_3168);
and U5403 (N_5403,N_2678,N_1863);
and U5404 (N_5404,N_706,N_2845);
and U5405 (N_5405,N_4782,N_2853);
nand U5406 (N_5406,N_701,N_1572);
and U5407 (N_5407,N_947,N_3748);
nand U5408 (N_5408,N_4920,N_59);
or U5409 (N_5409,N_3956,N_3391);
nand U5410 (N_5410,N_1898,N_4433);
nor U5411 (N_5411,N_4956,N_1527);
and U5412 (N_5412,N_4901,N_2388);
and U5413 (N_5413,N_4811,N_570);
nand U5414 (N_5414,N_3725,N_2437);
and U5415 (N_5415,N_4035,N_941);
nand U5416 (N_5416,N_1789,N_1720);
nor U5417 (N_5417,N_3408,N_4524);
or U5418 (N_5418,N_1713,N_3440);
or U5419 (N_5419,N_3873,N_3844);
and U5420 (N_5420,N_2603,N_1088);
nand U5421 (N_5421,N_951,N_4963);
and U5422 (N_5422,N_1145,N_124);
nor U5423 (N_5423,N_1950,N_1885);
and U5424 (N_5424,N_4478,N_1300);
nand U5425 (N_5425,N_3026,N_965);
nor U5426 (N_5426,N_3595,N_2048);
nand U5427 (N_5427,N_4870,N_3991);
nor U5428 (N_5428,N_398,N_1793);
nor U5429 (N_5429,N_52,N_3800);
and U5430 (N_5430,N_1944,N_1079);
nor U5431 (N_5431,N_1107,N_4167);
xnor U5432 (N_5432,N_629,N_1562);
nand U5433 (N_5433,N_4296,N_1747);
or U5434 (N_5434,N_2544,N_1705);
or U5435 (N_5435,N_1903,N_1343);
or U5436 (N_5436,N_2322,N_3793);
or U5437 (N_5437,N_3798,N_3931);
xor U5438 (N_5438,N_2037,N_3989);
and U5439 (N_5439,N_2556,N_2583);
or U5440 (N_5440,N_2633,N_331);
and U5441 (N_5441,N_2072,N_3845);
and U5442 (N_5442,N_2792,N_3717);
nand U5443 (N_5443,N_493,N_1566);
nor U5444 (N_5444,N_470,N_677);
or U5445 (N_5445,N_3548,N_741);
or U5446 (N_5446,N_649,N_406);
or U5447 (N_5447,N_4786,N_1296);
and U5448 (N_5448,N_435,N_2829);
and U5449 (N_5449,N_2243,N_1271);
or U5450 (N_5450,N_4139,N_949);
or U5451 (N_5451,N_72,N_4207);
nor U5452 (N_5452,N_4425,N_147);
nor U5453 (N_5453,N_3074,N_3607);
and U5454 (N_5454,N_1651,N_514);
nor U5455 (N_5455,N_874,N_2203);
or U5456 (N_5456,N_4084,N_1320);
nor U5457 (N_5457,N_4006,N_619);
or U5458 (N_5458,N_3298,N_3981);
and U5459 (N_5459,N_3749,N_2996);
xor U5460 (N_5460,N_2956,N_2151);
nand U5461 (N_5461,N_792,N_3294);
nand U5462 (N_5462,N_2817,N_2433);
nor U5463 (N_5463,N_1812,N_4827);
nand U5464 (N_5464,N_126,N_2275);
nand U5465 (N_5465,N_1553,N_4634);
nand U5466 (N_5466,N_1216,N_3806);
nor U5467 (N_5467,N_1319,N_1184);
or U5468 (N_5468,N_2913,N_3552);
and U5469 (N_5469,N_1766,N_918);
or U5470 (N_5470,N_1986,N_4440);
and U5471 (N_5471,N_215,N_4783);
nor U5472 (N_5472,N_4645,N_1773);
nor U5473 (N_5473,N_4658,N_2240);
and U5474 (N_5474,N_1661,N_3518);
and U5475 (N_5475,N_474,N_1669);
nand U5476 (N_5476,N_405,N_4295);
xor U5477 (N_5477,N_43,N_606);
or U5478 (N_5478,N_553,N_4831);
nand U5479 (N_5479,N_1150,N_4477);
nand U5480 (N_5480,N_2163,N_3675);
or U5481 (N_5481,N_409,N_421);
nor U5482 (N_5482,N_4321,N_705);
nor U5483 (N_5483,N_3922,N_1883);
nor U5484 (N_5484,N_2239,N_590);
nand U5485 (N_5485,N_4541,N_4444);
nand U5486 (N_5486,N_2591,N_3219);
and U5487 (N_5487,N_4287,N_3444);
or U5488 (N_5488,N_4625,N_1362);
nand U5489 (N_5489,N_1737,N_1610);
and U5490 (N_5490,N_4345,N_4755);
nor U5491 (N_5491,N_3670,N_600);
nand U5492 (N_5492,N_1139,N_4078);
or U5493 (N_5493,N_1614,N_4614);
or U5494 (N_5494,N_2716,N_958);
xor U5495 (N_5495,N_940,N_390);
nand U5496 (N_5496,N_2460,N_836);
and U5497 (N_5497,N_4971,N_1504);
nand U5498 (N_5498,N_3333,N_2623);
nor U5499 (N_5499,N_4030,N_3930);
nor U5500 (N_5500,N_3005,N_3889);
nor U5501 (N_5501,N_3853,N_3661);
and U5502 (N_5502,N_754,N_4772);
or U5503 (N_5503,N_2461,N_1958);
and U5504 (N_5504,N_1882,N_1494);
xor U5505 (N_5505,N_4620,N_672);
nand U5506 (N_5506,N_109,N_4498);
nand U5507 (N_5507,N_3926,N_3075);
nand U5508 (N_5508,N_2480,N_3878);
nand U5509 (N_5509,N_1655,N_887);
nor U5510 (N_5510,N_25,N_1106);
nand U5511 (N_5511,N_2312,N_1935);
and U5512 (N_5512,N_2207,N_1317);
xor U5513 (N_5513,N_4662,N_3689);
nor U5514 (N_5514,N_1930,N_4600);
or U5515 (N_5515,N_1810,N_3516);
and U5516 (N_5516,N_3059,N_339);
or U5517 (N_5517,N_304,N_1460);
nor U5518 (N_5518,N_3276,N_222);
or U5519 (N_5519,N_4787,N_2107);
nor U5520 (N_5520,N_1718,N_2448);
nand U5521 (N_5521,N_1627,N_3815);
and U5522 (N_5522,N_3134,N_3773);
or U5523 (N_5523,N_3460,N_664);
or U5524 (N_5524,N_520,N_1000);
or U5525 (N_5525,N_638,N_998);
or U5526 (N_5526,N_476,N_3338);
or U5527 (N_5527,N_4753,N_4812);
nor U5528 (N_5528,N_407,N_114);
or U5529 (N_5529,N_1850,N_3663);
or U5530 (N_5530,N_3175,N_4247);
and U5531 (N_5531,N_1442,N_363);
or U5532 (N_5532,N_4429,N_4825);
or U5533 (N_5533,N_4778,N_1811);
and U5534 (N_5534,N_4664,N_4919);
and U5535 (N_5535,N_1295,N_1595);
or U5536 (N_5536,N_4813,N_4581);
or U5537 (N_5537,N_1799,N_4297);
and U5538 (N_5538,N_3138,N_1828);
and U5539 (N_5539,N_3851,N_1694);
or U5540 (N_5540,N_1604,N_2978);
xnor U5541 (N_5541,N_1568,N_2100);
nand U5542 (N_5542,N_1437,N_1174);
or U5543 (N_5543,N_3751,N_4341);
nand U5544 (N_5544,N_218,N_3091);
nand U5545 (N_5545,N_254,N_1381);
and U5546 (N_5546,N_2865,N_2923);
nor U5547 (N_5547,N_354,N_2434);
nand U5548 (N_5548,N_4339,N_3182);
nand U5549 (N_5549,N_801,N_1933);
nand U5550 (N_5550,N_622,N_4531);
nor U5551 (N_5551,N_392,N_2006);
nor U5552 (N_5552,N_3797,N_1556);
nor U5553 (N_5553,N_3260,N_2930);
nor U5554 (N_5554,N_348,N_986);
nor U5555 (N_5555,N_4301,N_3710);
or U5556 (N_5556,N_3303,N_2742);
nor U5557 (N_5557,N_4087,N_4849);
nand U5558 (N_5558,N_3337,N_2587);
or U5559 (N_5559,N_4739,N_4803);
and U5560 (N_5560,N_4213,N_1817);
nor U5561 (N_5561,N_3825,N_74);
nor U5562 (N_5562,N_3537,N_44);
and U5563 (N_5563,N_1998,N_4051);
and U5564 (N_5564,N_3908,N_4676);
and U5565 (N_5565,N_90,N_2509);
or U5566 (N_5566,N_1038,N_2938);
nand U5567 (N_5567,N_485,N_3257);
nand U5568 (N_5568,N_3082,N_103);
or U5569 (N_5569,N_7,N_3619);
nor U5570 (N_5570,N_4872,N_2719);
nand U5571 (N_5571,N_1010,N_1801);
nand U5572 (N_5572,N_528,N_4763);
nand U5573 (N_5573,N_3898,N_177);
nor U5574 (N_5574,N_2449,N_914);
or U5575 (N_5575,N_2359,N_2622);
nor U5576 (N_5576,N_4090,N_4902);
and U5577 (N_5577,N_3151,N_4143);
and U5578 (N_5578,N_3928,N_2959);
nand U5579 (N_5579,N_580,N_595);
and U5580 (N_5580,N_2675,N_110);
nand U5581 (N_5581,N_3669,N_3876);
and U5582 (N_5582,N_4454,N_2114);
nand U5583 (N_5583,N_4347,N_4437);
nor U5584 (N_5584,N_4350,N_3915);
nand U5585 (N_5585,N_4317,N_63);
and U5586 (N_5586,N_743,N_3166);
or U5587 (N_5587,N_95,N_3514);
or U5588 (N_5588,N_4391,N_1330);
nand U5589 (N_5589,N_2189,N_3406);
nand U5590 (N_5590,N_2096,N_1546);
or U5591 (N_5591,N_574,N_4226);
and U5592 (N_5592,N_1206,N_497);
and U5593 (N_5593,N_3202,N_1425);
xnor U5594 (N_5594,N_1041,N_2928);
nand U5595 (N_5595,N_1411,N_1102);
nand U5596 (N_5596,N_3940,N_3843);
or U5597 (N_5597,N_584,N_854);
and U5598 (N_5598,N_2739,N_4233);
or U5599 (N_5599,N_4840,N_1449);
nand U5600 (N_5600,N_913,N_4399);
nor U5601 (N_5601,N_1739,N_4494);
nand U5602 (N_5602,N_4228,N_4748);
or U5603 (N_5603,N_2293,N_3982);
nor U5604 (N_5604,N_2033,N_3107);
or U5605 (N_5605,N_3270,N_608);
and U5606 (N_5606,N_2743,N_3304);
nor U5607 (N_5607,N_3330,N_1867);
nor U5608 (N_5608,N_1975,N_2363);
nor U5609 (N_5609,N_2276,N_830);
and U5610 (N_5610,N_3137,N_3994);
nor U5611 (N_5611,N_2789,N_1305);
nor U5612 (N_5612,N_337,N_4774);
and U5613 (N_5613,N_1498,N_1565);
and U5614 (N_5614,N_1522,N_123);
or U5615 (N_5615,N_3350,N_994);
or U5616 (N_5616,N_3596,N_4874);
xnor U5617 (N_5617,N_4180,N_1990);
nand U5618 (N_5618,N_1650,N_1922);
and U5619 (N_5619,N_4422,N_1755);
or U5620 (N_5620,N_1829,N_956);
nand U5621 (N_5621,N_2268,N_174);
or U5622 (N_5622,N_2365,N_652);
and U5623 (N_5623,N_3183,N_4623);
or U5624 (N_5624,N_3527,N_451);
or U5625 (N_5625,N_1180,N_4385);
and U5626 (N_5626,N_2944,N_1458);
nand U5627 (N_5627,N_765,N_3830);
and U5628 (N_5628,N_1301,N_2051);
or U5629 (N_5629,N_1325,N_1350);
nand U5630 (N_5630,N_2289,N_1476);
and U5631 (N_5631,N_4062,N_1322);
nand U5632 (N_5632,N_4091,N_616);
nor U5633 (N_5633,N_2219,N_4924);
and U5634 (N_5634,N_1642,N_3209);
or U5635 (N_5635,N_3381,N_2147);
and U5636 (N_5636,N_3037,N_3760);
nor U5637 (N_5637,N_821,N_280);
and U5638 (N_5638,N_2876,N_1608);
nor U5639 (N_5639,N_1653,N_4147);
nor U5640 (N_5640,N_1355,N_4630);
and U5641 (N_5641,N_2979,N_2512);
and U5642 (N_5642,N_783,N_344);
or U5643 (N_5643,N_2850,N_117);
nand U5644 (N_5644,N_2569,N_2726);
or U5645 (N_5645,N_1110,N_422);
or U5646 (N_5646,N_3421,N_262);
xor U5647 (N_5647,N_1230,N_875);
nand U5648 (N_5648,N_1561,N_2827);
xnor U5649 (N_5649,N_1752,N_2182);
nand U5650 (N_5650,N_2032,N_2842);
and U5651 (N_5651,N_1632,N_4409);
nand U5652 (N_5652,N_163,N_3702);
and U5653 (N_5653,N_2574,N_4116);
or U5654 (N_5654,N_720,N_2);
and U5655 (N_5655,N_3759,N_3769);
or U5656 (N_5656,N_1544,N_1851);
xor U5657 (N_5657,N_2416,N_577);
nor U5658 (N_5658,N_3359,N_1615);
xor U5659 (N_5659,N_4324,N_1529);
nand U5660 (N_5660,N_2815,N_55);
or U5661 (N_5661,N_3606,N_1820);
nand U5662 (N_5662,N_1517,N_3241);
or U5663 (N_5663,N_989,N_680);
or U5664 (N_5664,N_450,N_3519);
and U5665 (N_5665,N_2999,N_4597);
and U5666 (N_5666,N_4258,N_3985);
nand U5667 (N_5667,N_1949,N_807);
and U5668 (N_5668,N_3895,N_4903);
or U5669 (N_5669,N_3620,N_4298);
and U5670 (N_5670,N_53,N_1179);
and U5671 (N_5671,N_3113,N_2656);
and U5672 (N_5672,N_2098,N_933);
and U5673 (N_5673,N_2892,N_4218);
and U5674 (N_5674,N_4219,N_1973);
and U5675 (N_5675,N_740,N_365);
or U5676 (N_5676,N_3470,N_4854);
nor U5677 (N_5677,N_4940,N_2336);
nor U5678 (N_5678,N_2524,N_825);
nor U5679 (N_5679,N_3581,N_3651);
and U5680 (N_5680,N_2769,N_1441);
nor U5681 (N_5681,N_1589,N_324);
nor U5682 (N_5682,N_697,N_4504);
nor U5683 (N_5683,N_3724,N_2023);
nor U5684 (N_5684,N_2376,N_83);
or U5685 (N_5685,N_2206,N_224);
xnor U5686 (N_5686,N_561,N_256);
nor U5687 (N_5687,N_1692,N_4307);
nor U5688 (N_5688,N_3286,N_3251);
or U5689 (N_5689,N_700,N_263);
nor U5690 (N_5690,N_3508,N_943);
nor U5691 (N_5691,N_2939,N_1104);
nand U5692 (N_5692,N_2972,N_873);
and U5693 (N_5693,N_3351,N_3540);
nand U5694 (N_5694,N_4950,N_1416);
nand U5695 (N_5695,N_3912,N_704);
nor U5696 (N_5696,N_1716,N_2920);
nand U5697 (N_5697,N_1193,N_1537);
or U5698 (N_5698,N_4231,N_1266);
and U5699 (N_5699,N_3309,N_1237);
nor U5700 (N_5700,N_3423,N_28);
or U5701 (N_5701,N_4163,N_4290);
nor U5702 (N_5702,N_2320,N_2833);
or U5703 (N_5703,N_4727,N_2862);
or U5704 (N_5704,N_3664,N_2124);
nand U5705 (N_5705,N_4377,N_4359);
nor U5706 (N_5706,N_3050,N_4253);
or U5707 (N_5707,N_1822,N_1378);
nand U5708 (N_5708,N_2800,N_2709);
or U5709 (N_5709,N_3789,N_3264);
nand U5710 (N_5710,N_2478,N_4996);
nand U5711 (N_5711,N_4871,N_2317);
nand U5712 (N_5712,N_1477,N_3329);
and U5713 (N_5713,N_4652,N_1005);
or U5714 (N_5714,N_2115,N_2458);
nand U5715 (N_5715,N_4607,N_3852);
nor U5716 (N_5716,N_1847,N_2375);
and U5717 (N_5717,N_3525,N_4202);
xnor U5718 (N_5718,N_2076,N_1168);
or U5719 (N_5719,N_3549,N_2502);
nor U5720 (N_5720,N_3904,N_3807);
and U5721 (N_5721,N_400,N_746);
and U5722 (N_5722,N_1085,N_1280);
and U5723 (N_5723,N_3126,N_2657);
and U5724 (N_5724,N_34,N_3185);
and U5725 (N_5725,N_492,N_1345);
or U5726 (N_5726,N_77,N_552);
and U5727 (N_5727,N_4560,N_4837);
nand U5728 (N_5728,N_2441,N_4354);
or U5729 (N_5729,N_3078,N_3623);
nand U5730 (N_5730,N_488,N_3860);
nor U5731 (N_5731,N_1126,N_3627);
or U5732 (N_5732,N_3935,N_3966);
or U5733 (N_5733,N_2205,N_3089);
nor U5734 (N_5734,N_4559,N_401);
and U5735 (N_5735,N_587,N_1900);
nor U5736 (N_5736,N_279,N_766);
or U5737 (N_5737,N_314,N_2746);
and U5738 (N_5738,N_2849,N_1341);
and U5739 (N_5739,N_4389,N_1093);
and U5740 (N_5740,N_3672,N_1836);
and U5741 (N_5741,N_2688,N_4954);
and U5742 (N_5742,N_2162,N_4161);
or U5743 (N_5743,N_3283,N_2609);
nand U5744 (N_5744,N_1508,N_653);
or U5745 (N_5745,N_500,N_1349);
or U5746 (N_5746,N_1735,N_4263);
and U5747 (N_5747,N_4292,N_1291);
nand U5748 (N_5748,N_179,N_48);
or U5749 (N_5749,N_3681,N_1192);
nor U5750 (N_5750,N_2612,N_1756);
nand U5751 (N_5751,N_3020,N_4378);
nor U5752 (N_5752,N_1056,N_4502);
and U5753 (N_5753,N_3932,N_1987);
nand U5754 (N_5754,N_281,N_2797);
nand U5755 (N_5755,N_1018,N_1326);
nand U5756 (N_5756,N_3632,N_4732);
nand U5757 (N_5757,N_173,N_437);
and U5758 (N_5758,N_1427,N_735);
nand U5759 (N_5759,N_4925,N_1299);
nor U5760 (N_5760,N_3027,N_1131);
nand U5761 (N_5761,N_1996,N_2265);
or U5762 (N_5762,N_2785,N_4775);
and U5763 (N_5763,N_4964,N_4507);
nor U5764 (N_5764,N_1879,N_1327);
nor U5765 (N_5765,N_1834,N_361);
and U5766 (N_5766,N_1154,N_4632);
nor U5767 (N_5767,N_627,N_2300);
and U5768 (N_5768,N_791,N_498);
nand U5769 (N_5769,N_3300,N_3443);
or U5770 (N_5770,N_3839,N_4474);
and U5771 (N_5771,N_11,N_1157);
nand U5772 (N_5772,N_2601,N_4795);
nor U5773 (N_5773,N_4522,N_2632);
and U5774 (N_5774,N_3575,N_4303);
or U5775 (N_5775,N_1160,N_2974);
nor U5776 (N_5776,N_2872,N_1573);
and U5777 (N_5777,N_1843,N_3237);
xnor U5778 (N_5778,N_4716,N_2916);
and U5779 (N_5779,N_4895,N_882);
xor U5780 (N_5780,N_257,N_4125);
nand U5781 (N_5781,N_832,N_1645);
nand U5782 (N_5782,N_128,N_1685);
and U5783 (N_5783,N_3053,N_3158);
nor U5784 (N_5784,N_4269,N_911);
nor U5785 (N_5785,N_1369,N_3945);
nor U5786 (N_5786,N_2213,N_3835);
and U5787 (N_5787,N_3721,N_85);
or U5788 (N_5788,N_4137,N_4711);
nand U5789 (N_5789,N_3341,N_4709);
nand U5790 (N_5790,N_4476,N_242);
and U5791 (N_5791,N_149,N_1204);
nand U5792 (N_5792,N_1955,N_2883);
nand U5793 (N_5793,N_2987,N_4611);
or U5794 (N_5794,N_879,N_845);
nand U5795 (N_5795,N_2522,N_2751);
or U5796 (N_5796,N_2647,N_402);
nand U5797 (N_5797,N_2929,N_239);
and U5798 (N_5798,N_2602,N_4565);
nand U5799 (N_5799,N_1044,N_1340);
nor U5800 (N_5800,N_2638,N_2700);
nor U5801 (N_5801,N_2457,N_4353);
nor U5802 (N_5802,N_4111,N_1648);
or U5803 (N_5803,N_3402,N_62);
and U5804 (N_5804,N_1001,N_115);
nor U5805 (N_5805,N_4103,N_1424);
or U5806 (N_5806,N_1050,N_3943);
nor U5807 (N_5807,N_1993,N_1352);
or U5808 (N_5808,N_4603,N_3235);
and U5809 (N_5809,N_3867,N_2152);
nor U5810 (N_5810,N_1652,N_1078);
nand U5811 (N_5811,N_1901,N_843);
nand U5812 (N_5812,N_1940,N_2034);
or U5813 (N_5813,N_4236,N_4529);
or U5814 (N_5814,N_4856,N_3979);
or U5815 (N_5815,N_3605,N_2475);
xor U5816 (N_5816,N_1096,N_3442);
and U5817 (N_5817,N_1721,N_14);
or U5818 (N_5818,N_4470,N_2693);
or U5819 (N_5819,N_4428,N_1969);
and U5820 (N_5820,N_777,N_12);
nor U5821 (N_5821,N_2090,N_2629);
nor U5822 (N_5822,N_3457,N_1112);
nor U5823 (N_5823,N_3397,N_3757);
nand U5824 (N_5824,N_169,N_4311);
xor U5825 (N_5825,N_3636,N_3492);
and U5826 (N_5826,N_2936,N_837);
xor U5827 (N_5827,N_2752,N_4717);
xnor U5828 (N_5828,N_1782,N_80);
or U5829 (N_5829,N_4496,N_3531);
nand U5830 (N_5830,N_1238,N_991);
and U5831 (N_5831,N_2788,N_443);
nand U5832 (N_5832,N_4958,N_3695);
nand U5833 (N_5833,N_3745,N_3794);
nor U5834 (N_5834,N_2232,N_3108);
nand U5835 (N_5835,N_4548,N_1062);
or U5836 (N_5836,N_4697,N_1957);
and U5837 (N_5837,N_555,N_4737);
nand U5838 (N_5838,N_2042,N_4240);
and U5839 (N_5839,N_2381,N_2950);
nand U5840 (N_5840,N_3163,N_2659);
and U5841 (N_5841,N_1354,N_21);
nand U5842 (N_5842,N_2699,N_4047);
or U5843 (N_5843,N_928,N_4280);
and U5844 (N_5844,N_477,N_2809);
or U5845 (N_5845,N_2744,N_839);
or U5846 (N_5846,N_4257,N_1198);
nand U5847 (N_5847,N_1968,N_136);
or U5848 (N_5848,N_4032,N_1995);
nand U5849 (N_5849,N_3520,N_1331);
nor U5850 (N_5850,N_2222,N_2309);
and U5851 (N_5851,N_3079,N_3455);
and U5852 (N_5852,N_2447,N_708);
or U5853 (N_5853,N_1312,N_1569);
or U5854 (N_5854,N_630,N_4199);
and U5855 (N_5855,N_824,N_3657);
nor U5856 (N_5856,N_2183,N_3859);
nor U5857 (N_5857,N_1447,N_3293);
and U5858 (N_5858,N_345,N_3535);
or U5859 (N_5859,N_4557,N_2970);
nor U5860 (N_5860,N_1623,N_2223);
and U5861 (N_5861,N_1639,N_572);
and U5862 (N_5862,N_2249,N_1874);
nor U5863 (N_5863,N_3291,N_3150);
nand U5864 (N_5864,N_1022,N_1194);
nand U5865 (N_5865,N_1732,N_380);
and U5866 (N_5866,N_1686,N_4883);
nor U5867 (N_5867,N_4583,N_3996);
nor U5868 (N_5868,N_1313,N_285);
nand U5869 (N_5869,N_1328,N_4314);
nor U5870 (N_5870,N_2308,N_4371);
nand U5871 (N_5871,N_58,N_2450);
nand U5872 (N_5872,N_234,N_3903);
nand U5873 (N_5873,N_3854,N_4699);
nand U5874 (N_5874,N_1757,N_245);
and U5875 (N_5875,N_863,N_2573);
and U5876 (N_5876,N_1684,N_3214);
and U5877 (N_5877,N_3279,N_1489);
or U5878 (N_5878,N_125,N_3204);
or U5879 (N_5879,N_2155,N_1284);
and U5880 (N_5880,N_3401,N_930);
or U5881 (N_5881,N_1511,N_1579);
nor U5882 (N_5882,N_3363,N_6);
nor U5883 (N_5883,N_3658,N_3068);
nor U5884 (N_5884,N_465,N_1656);
and U5885 (N_5885,N_480,N_4426);
and U5886 (N_5886,N_4917,N_1082);
nor U5887 (N_5887,N_4537,N_1399);
nor U5888 (N_5888,N_527,N_1963);
nor U5889 (N_5889,N_1202,N_2294);
nor U5890 (N_5890,N_692,N_4701);
nand U5891 (N_5891,N_4140,N_3744);
xor U5892 (N_5892,N_3927,N_42);
and U5893 (N_5893,N_1858,N_290);
nand U5894 (N_5894,N_75,N_3767);
xor U5895 (N_5895,N_1187,N_1668);
nor U5896 (N_5896,N_3348,N_4109);
or U5897 (N_5897,N_298,N_1436);
and U5898 (N_5898,N_1229,N_4265);
and U5899 (N_5899,N_3849,N_1137);
and U5900 (N_5900,N_1274,N_2398);
nor U5901 (N_5901,N_3342,N_4413);
or U5902 (N_5902,N_1143,N_4887);
or U5903 (N_5903,N_789,N_3288);
nand U5904 (N_5904,N_2771,N_2757);
or U5905 (N_5905,N_2666,N_1943);
or U5906 (N_5906,N_3232,N_2095);
and U5907 (N_5907,N_4605,N_3780);
or U5908 (N_5908,N_4519,N_1842);
nor U5909 (N_5909,N_495,N_182);
nor U5910 (N_5910,N_4394,N_3735);
or U5911 (N_5911,N_272,N_3469);
and U5912 (N_5912,N_4332,N_1469);
nor U5913 (N_5913,N_2501,N_3957);
xor U5914 (N_5914,N_1833,N_3819);
and U5915 (N_5915,N_3804,N_3616);
or U5916 (N_5916,N_1976,N_3587);
nor U5917 (N_5917,N_4355,N_3285);
or U5918 (N_5918,N_683,N_2776);
nor U5919 (N_5919,N_782,N_4037);
nor U5920 (N_5920,N_2873,N_626);
and U5921 (N_5921,N_2077,N_383);
nand U5922 (N_5922,N_4083,N_3894);
nor U5923 (N_5923,N_1577,N_4936);
or U5924 (N_5924,N_601,N_3473);
or U5925 (N_5925,N_3883,N_2723);
and U5926 (N_5926,N_4119,N_781);
or U5927 (N_5927,N_2953,N_571);
and U5928 (N_5928,N_2957,N_4540);
and U5929 (N_5929,N_4928,N_130);
nor U5930 (N_5930,N_3419,N_870);
and U5931 (N_5931,N_642,N_4666);
nor U5932 (N_5932,N_2490,N_3733);
xnor U5933 (N_5933,N_1120,N_1832);
nand U5934 (N_5934,N_2225,N_3112);
or U5935 (N_5935,N_3224,N_311);
nor U5936 (N_5936,N_3153,N_2242);
or U5937 (N_5937,N_4943,N_816);
or U5938 (N_5938,N_4735,N_3533);
nor U5939 (N_5939,N_2564,N_1007);
nor U5940 (N_5940,N_3233,N_327);
nor U5941 (N_5941,N_2732,N_1719);
or U5942 (N_5942,N_1115,N_639);
nand U5943 (N_5943,N_2039,N_4712);
nand U5944 (N_5944,N_2765,N_4134);
or U5945 (N_5945,N_2333,N_104);
and U5946 (N_5946,N_3358,N_2231);
and U5947 (N_5947,N_3667,N_3128);
nor U5948 (N_5948,N_138,N_2281);
nand U5949 (N_5949,N_3320,N_2910);
nor U5950 (N_5950,N_4822,N_94);
nand U5951 (N_5951,N_3716,N_1835);
nor U5952 (N_5952,N_1097,N_4959);
or U5953 (N_5953,N_4922,N_3105);
nor U5954 (N_5954,N_2986,N_3696);
or U5955 (N_5955,N_1803,N_2417);
nor U5956 (N_5956,N_4585,N_4517);
nand U5957 (N_5957,N_3737,N_1);
or U5958 (N_5958,N_2245,N_1515);
and U5959 (N_5959,N_2024,N_424);
and U5960 (N_5960,N_2291,N_3077);
and U5961 (N_5961,N_475,N_3164);
and U5962 (N_5962,N_3498,N_4973);
or U5963 (N_5963,N_2634,N_1777);
and U5964 (N_5964,N_3340,N_1069);
nand U5965 (N_5965,N_4198,N_4485);
or U5966 (N_5966,N_684,N_4001);
xnor U5967 (N_5967,N_181,N_3591);
nand U5968 (N_5968,N_950,N_3811);
nor U5969 (N_5969,N_3326,N_3039);
or U5970 (N_5970,N_4025,N_1047);
nand U5971 (N_5971,N_4348,N_3677);
or U5972 (N_5972,N_4944,N_675);
or U5973 (N_5973,N_1117,N_3384);
or U5974 (N_5974,N_734,N_3618);
and U5975 (N_5975,N_4523,N_3732);
or U5976 (N_5976,N_2774,N_2992);
nand U5977 (N_5977,N_4738,N_1999);
nor U5978 (N_5978,N_3684,N_4828);
nor U5979 (N_5979,N_3255,N_2995);
xnor U5980 (N_5980,N_1855,N_1492);
nor U5981 (N_5981,N_4506,N_2078);
nand U5982 (N_5982,N_4911,N_925);
or U5983 (N_5983,N_538,N_4687);
and U5984 (N_5984,N_4584,N_2172);
or U5985 (N_5985,N_1733,N_948);
or U5986 (N_5986,N_3147,N_2355);
nand U5987 (N_5987,N_1865,N_3768);
nor U5988 (N_5988,N_1026,N_1480);
or U5989 (N_5989,N_650,N_3803);
and U5990 (N_5990,N_4923,N_3060);
and U5991 (N_5991,N_3146,N_1525);
or U5992 (N_5992,N_4484,N_3256);
and U5993 (N_5993,N_4579,N_3093);
nor U5994 (N_5994,N_160,N_1887);
nor U5995 (N_5995,N_1215,N_4423);
nor U5996 (N_5996,N_2148,N_2802);
nor U5997 (N_5997,N_4626,N_3836);
and U5998 (N_5998,N_1816,N_2044);
nand U5999 (N_5999,N_4227,N_1574);
or U6000 (N_6000,N_3610,N_1073);
and U6001 (N_6001,N_4665,N_1890);
nor U6002 (N_6002,N_4796,N_3404);
and U6003 (N_6003,N_4182,N_4534);
and U6004 (N_6004,N_1413,N_809);
nand U6005 (N_6005,N_3121,N_628);
nor U6006 (N_6006,N_583,N_1907);
nand U6007 (N_6007,N_4416,N_607);
or U6008 (N_6008,N_2857,N_2046);
and U6009 (N_6009,N_2267,N_387);
and U6010 (N_6010,N_4279,N_3495);
or U6011 (N_6011,N_1212,N_4547);
nand U6012 (N_6012,N_4511,N_632);
nand U6013 (N_6013,N_3801,N_134);
or U6014 (N_6014,N_3923,N_2881);
and U6015 (N_6015,N_534,N_2821);
nand U6016 (N_6016,N_3267,N_1173);
nor U6017 (N_6017,N_3383,N_3588);
or U6018 (N_6018,N_4456,N_338);
nor U6019 (N_6019,N_1926,N_504);
xnor U6020 (N_6020,N_153,N_4636);
and U6021 (N_6021,N_3295,N_1337);
or U6022 (N_6022,N_3709,N_3715);
or U6023 (N_6023,N_3085,N_1586);
and U6024 (N_6024,N_3355,N_4589);
or U6025 (N_6025,N_1902,N_3428);
nand U6026 (N_6026,N_3754,N_237);
nand U6027 (N_6027,N_1538,N_3585);
or U6028 (N_6028,N_353,N_973);
nor U6029 (N_6029,N_190,N_4744);
nor U6030 (N_6030,N_4723,N_1470);
or U6031 (N_6031,N_1019,N_4362);
or U6032 (N_6032,N_2834,N_229);
or U6033 (N_6033,N_3254,N_2555);
and U6034 (N_6034,N_4587,N_3788);
nor U6035 (N_6035,N_4692,N_3529);
nand U6036 (N_6036,N_3070,N_1533);
nor U6037 (N_6037,N_3055,N_1499);
xor U6038 (N_6038,N_4049,N_1783);
nand U6039 (N_6039,N_3727,N_3437);
nand U6040 (N_6040,N_4346,N_4642);
or U6041 (N_6041,N_1941,N_3367);
nor U6042 (N_6042,N_641,N_4320);
and U6043 (N_6043,N_4865,N_3208);
or U6044 (N_6044,N_226,N_1625);
and U6045 (N_6045,N_2101,N_1960);
nor U6046 (N_6046,N_562,N_1323);
and U6047 (N_6047,N_3145,N_1396);
nand U6048 (N_6048,N_249,N_1321);
and U6049 (N_6049,N_2590,N_2571);
xor U6050 (N_6050,N_3949,N_979);
nand U6051 (N_6051,N_2442,N_4515);
and U6052 (N_6052,N_1228,N_4703);
or U6053 (N_6053,N_1778,N_3040);
nor U6054 (N_6054,N_3129,N_2720);
or U6055 (N_6055,N_2306,N_180);
and U6056 (N_6056,N_3281,N_739);
nor U6057 (N_6057,N_1951,N_2472);
and U6058 (N_6058,N_1700,N_4105);
and U6059 (N_6059,N_1393,N_838);
and U6060 (N_6060,N_3886,N_1849);
and U6061 (N_6061,N_4619,N_4170);
or U6062 (N_6062,N_4777,N_2060);
and U6063 (N_6063,N_937,N_3282);
and U6064 (N_6064,N_3353,N_924);
and U6065 (N_6065,N_3863,N_2053);
nor U6066 (N_6066,N_1365,N_3305);
or U6067 (N_6067,N_3345,N_1671);
and U6068 (N_6068,N_1391,N_3746);
nor U6069 (N_6069,N_4206,N_788);
and U6070 (N_6070,N_1479,N_4185);
or U6071 (N_6071,N_464,N_4186);
or U6072 (N_6072,N_2266,N_3738);
nand U6073 (N_6073,N_3875,N_419);
or U6074 (N_6074,N_1214,N_2637);
xnor U6075 (N_6075,N_3081,N_648);
nand U6076 (N_6076,N_3579,N_1776);
nand U6077 (N_6077,N_1823,N_158);
nor U6078 (N_6078,N_3592,N_4432);
nand U6079 (N_6079,N_3980,N_4993);
or U6080 (N_6080,N_3420,N_3371);
nor U6081 (N_6081,N_4718,N_2577);
xnor U6082 (N_6082,N_2117,N_4117);
and U6083 (N_6083,N_3888,N_1015);
and U6084 (N_6084,N_1927,N_1965);
nand U6085 (N_6085,N_731,N_1169);
nor U6086 (N_6086,N_3373,N_976);
or U6087 (N_6087,N_984,N_3905);
nand U6088 (N_6088,N_2504,N_4360);
or U6089 (N_6089,N_3708,N_2902);
and U6090 (N_6090,N_2030,N_1500);
nor U6091 (N_6091,N_3967,N_762);
xnor U6092 (N_6092,N_168,N_3758);
xor U6093 (N_6093,N_3680,N_129);
and U6094 (N_6094,N_2958,N_4070);
xor U6095 (N_6095,N_3174,N_4410);
and U6096 (N_6096,N_2173,N_1466);
or U6097 (N_6097,N_1709,N_2542);
xnor U6098 (N_6098,N_1484,N_1356);
or U6099 (N_6099,N_4889,N_3007);
nor U6100 (N_6100,N_4156,N_2229);
and U6101 (N_6101,N_4115,N_3140);
nor U6102 (N_6102,N_1118,N_981);
nand U6103 (N_6103,N_3659,N_369);
or U6104 (N_6104,N_2639,N_744);
nor U6105 (N_6105,N_1860,N_3047);
xnor U6106 (N_6106,N_2474,N_255);
or U6107 (N_6107,N_336,N_4340);
and U6108 (N_6108,N_1218,N_1039);
nor U6109 (N_6109,N_350,N_186);
nor U6110 (N_6110,N_3877,N_3740);
nor U6111 (N_6111,N_3558,N_3196);
or U6112 (N_6112,N_3781,N_4380);
nand U6113 (N_6113,N_1236,N_1895);
and U6114 (N_6114,N_3436,N_10);
or U6115 (N_6115,N_3099,N_2980);
nand U6116 (N_6116,N_2780,N_4593);
and U6117 (N_6117,N_1100,N_3475);
or U6118 (N_6118,N_2357,N_990);
nor U6119 (N_6119,N_3509,N_2604);
nor U6120 (N_6120,N_274,N_4881);
xor U6121 (N_6121,N_2277,N_847);
or U6122 (N_6122,N_4483,N_342);
and U6123 (N_6123,N_1932,N_2015);
nand U6124 (N_6124,N_2343,N_3812);
nand U6125 (N_6125,N_4171,N_3190);
and U6126 (N_6126,N_926,N_2505);
or U6127 (N_6127,N_3921,N_2476);
nor U6128 (N_6128,N_2710,N_533);
nand U6129 (N_6129,N_1602,N_1455);
or U6130 (N_6130,N_1846,N_1695);
nor U6131 (N_6131,N_1519,N_3327);
and U6132 (N_6132,N_2683,N_3389);
and U6133 (N_6133,N_2782,N_4855);
or U6134 (N_6134,N_2288,N_4897);
and U6135 (N_6135,N_1931,N_291);
xor U6136 (N_6136,N_2280,N_800);
and U6137 (N_6137,N_3778,N_4282);
and U6138 (N_6138,N_1952,N_4794);
and U6139 (N_6139,N_3808,N_1258);
nand U6140 (N_6140,N_3826,N_1638);
or U6141 (N_6141,N_1845,N_1612);
nor U6142 (N_6142,N_4168,N_4574);
or U6143 (N_6143,N_889,N_3486);
nor U6144 (N_6144,N_367,N_1045);
or U6145 (N_6145,N_1767,N_240);
and U6146 (N_6146,N_1269,N_4747);
and U6147 (N_6147,N_2302,N_978);
and U6148 (N_6148,N_4644,N_2506);
and U6149 (N_6149,N_4688,N_3559);
nor U6150 (N_6150,N_3818,N_3022);
or U6151 (N_6151,N_1798,N_2527);
or U6152 (N_6152,N_3564,N_3012);
or U6153 (N_6153,N_662,N_851);
nor U6154 (N_6154,N_267,N_457);
nor U6155 (N_6155,N_2123,N_1905);
nand U6156 (N_6156,N_758,N_712);
or U6157 (N_6157,N_2627,N_4053);
nor U6158 (N_6158,N_1734,N_39);
or U6159 (N_6159,N_4144,N_3919);
nor U6160 (N_6160,N_1977,N_3951);
and U6161 (N_6161,N_1394,N_2869);
or U6162 (N_6162,N_1770,N_1840);
nor U6163 (N_6163,N_4464,N_2001);
nor U6164 (N_6164,N_208,N_4318);
or U6165 (N_6165,N_2866,N_4395);
nor U6166 (N_6166,N_3297,N_4040);
or U6167 (N_6167,N_4162,N_2218);
nand U6168 (N_6168,N_375,N_200);
and U6169 (N_6169,N_3576,N_3541);
and U6170 (N_6170,N_521,N_4094);
and U6171 (N_6171,N_3438,N_31);
or U6172 (N_6172,N_1886,N_3234);
and U6173 (N_6173,N_1439,N_4217);
nand U6174 (N_6174,N_4834,N_2010);
or U6175 (N_6175,N_2258,N_2084);
or U6176 (N_6176,N_3307,N_3743);
and U6177 (N_6177,N_2488,N_4976);
nand U6178 (N_6178,N_1912,N_2334);
and U6179 (N_6179,N_3783,N_2942);
or U6180 (N_6180,N_4276,N_2352);
nor U6181 (N_6181,N_1273,N_2597);
xor U6182 (N_6182,N_4184,N_107);
nor U6183 (N_6183,N_2801,N_4088);
nand U6184 (N_6184,N_4724,N_4690);
and U6185 (N_6185,N_2065,N_1496);
nor U6186 (N_6186,N_417,N_4064);
or U6187 (N_6187,N_728,N_4445);
nor U6188 (N_6188,N_3615,N_3043);
nor U6189 (N_6189,N_852,N_2111);
xor U6190 (N_6190,N_4241,N_2701);
and U6191 (N_6191,N_305,N_2791);
or U6192 (N_6192,N_2157,N_586);
or U6193 (N_6193,N_1619,N_3067);
and U6194 (N_6194,N_4859,N_3869);
and U6195 (N_6195,N_4980,N_4571);
or U6196 (N_6196,N_2234,N_877);
nand U6197 (N_6197,N_2969,N_2420);
nor U6198 (N_6198,N_2099,N_1377);
and U6199 (N_6199,N_4128,N_2158);
nor U6200 (N_6200,N_3187,N_4988);
and U6201 (N_6201,N_2796,N_1920);
and U6202 (N_6202,N_4200,N_2523);
or U6203 (N_6203,N_241,N_2761);
or U6204 (N_6204,N_4098,N_3944);
nor U6205 (N_6205,N_1402,N_4598);
nand U6206 (N_6206,N_696,N_3563);
or U6207 (N_6207,N_3019,N_4017);
nor U6208 (N_6208,N_4602,N_4224);
xor U6209 (N_6209,N_3386,N_2685);
and U6210 (N_6210,N_2844,N_366);
and U6211 (N_6211,N_4259,N_3292);
nor U6212 (N_6212,N_2759,N_334);
and U6213 (N_6213,N_351,N_1894);
nor U6214 (N_6214,N_3155,N_2477);
nor U6215 (N_6215,N_4164,N_4042);
nand U6216 (N_6216,N_945,N_46);
nor U6217 (N_6217,N_3698,N_1233);
nor U6218 (N_6218,N_2915,N_4145);
or U6219 (N_6219,N_4024,N_68);
or U6220 (N_6220,N_4079,N_483);
or U6221 (N_6221,N_4610,N_2984);
nand U6222 (N_6222,N_3827,N_1551);
and U6223 (N_6223,N_2383,N_3924);
nand U6224 (N_6224,N_47,N_4858);
nor U6225 (N_6225,N_3016,N_4862);
and U6226 (N_6226,N_2818,N_1600);
or U6227 (N_6227,N_3998,N_231);
nand U6228 (N_6228,N_2725,N_248);
nand U6229 (N_6229,N_3049,N_4508);
nand U6230 (N_6230,N_3565,N_4214);
or U6231 (N_6231,N_602,N_2392);
or U6232 (N_6232,N_4309,N_1560);
nor U6233 (N_6233,N_2295,N_1649);
nand U6234 (N_6234,N_4734,N_3238);
xor U6235 (N_6235,N_3360,N_1023);
nand U6236 (N_6236,N_1929,N_3753);
or U6237 (N_6237,N_3496,N_2074);
nand U6238 (N_6238,N_2790,N_3649);
or U6239 (N_6239,N_993,N_2971);
nor U6240 (N_6240,N_2965,N_878);
xor U6241 (N_6241,N_4159,N_2411);
nand U6242 (N_6242,N_2135,N_4513);
xnor U6243 (N_6243,N_2236,N_165);
nand U6244 (N_6244,N_2768,N_4876);
nor U6245 (N_6245,N_4698,N_1916);
xnor U6246 (N_6246,N_711,N_487);
nor U6247 (N_6247,N_1438,N_1818);
xor U6248 (N_6248,N_2525,N_2314);
and U6249 (N_6249,N_3062,N_4628);
nand U6250 (N_6250,N_771,N_690);
and U6251 (N_6251,N_4204,N_2284);
nand U6252 (N_6252,N_3463,N_4677);
and U6253 (N_6253,N_2052,N_1768);
or U6254 (N_6254,N_2733,N_1617);
nand U6255 (N_6255,N_3418,N_4023);
and U6256 (N_6256,N_4471,N_2104);
nor U6257 (N_6257,N_812,N_2526);
or U6258 (N_6258,N_3643,N_4216);
or U6259 (N_6259,N_770,N_1430);
nand U6260 (N_6260,N_4654,N_3252);
or U6261 (N_6261,N_4438,N_718);
nand U6262 (N_6262,N_2462,N_3445);
and U6263 (N_6263,N_3766,N_3879);
and U6264 (N_6264,N_1909,N_2949);
or U6265 (N_6265,N_1101,N_1149);
nor U6266 (N_6266,N_2575,N_1122);
nand U6267 (N_6267,N_2283,N_49);
nand U6268 (N_6268,N_3747,N_388);
and U6269 (N_6269,N_2134,N_3858);
nand U6270 (N_6270,N_3100,N_3315);
and U6271 (N_6271,N_1231,N_3993);
and U6272 (N_6272,N_3705,N_872);
nor U6273 (N_6273,N_3977,N_1443);
and U6274 (N_6274,N_1526,N_1318);
and U6275 (N_6275,N_4918,N_2567);
nor U6276 (N_6276,N_4694,N_2344);
and U6277 (N_6277,N_2900,N_540);
nand U6278 (N_6278,N_1928,N_2611);
or U6279 (N_6279,N_2919,N_3538);
nor U6280 (N_6280,N_3779,N_1384);
xnor U6281 (N_6281,N_2453,N_2402);
and U6282 (N_6282,N_4806,N_3395);
nor U6283 (N_6283,N_1924,N_4669);
nor U6284 (N_6284,N_1934,N_3430);
nor U6285 (N_6285,N_4946,N_2595);
nor U6286 (N_6286,N_3130,N_1660);
nand U6287 (N_6287,N_1222,N_4390);
and U6288 (N_6288,N_3122,N_1790);
and U6289 (N_6289,N_2270,N_4588);
nand U6290 (N_6290,N_1133,N_3729);
or U6291 (N_6291,N_4417,N_4364);
nand U6292 (N_6292,N_2494,N_4728);
nand U6293 (N_6293,N_455,N_946);
xor U6294 (N_6294,N_211,N_2071);
and U6295 (N_6295,N_24,N_1547);
nor U6296 (N_6296,N_2874,N_4671);
nor U6297 (N_6297,N_4685,N_1510);
and U6298 (N_6298,N_386,N_4535);
and U6299 (N_6299,N_3431,N_4899);
and U6300 (N_6300,N_220,N_775);
or U6301 (N_6301,N_853,N_4990);
or U6302 (N_6302,N_621,N_2718);
nand U6303 (N_6303,N_4104,N_3965);
nor U6304 (N_6304,N_20,N_4984);
nor U6305 (N_6305,N_695,N_3603);
nor U6306 (N_6306,N_2891,N_2412);
nor U6307 (N_6307,N_4970,N_4335);
nor U6308 (N_6308,N_2444,N_3772);
and U6309 (N_6309,N_3561,N_235);
and U6310 (N_6310,N_1448,N_2263);
and U6311 (N_6311,N_228,N_2026);
xor U6312 (N_6312,N_4101,N_326);
xnor U6313 (N_6313,N_333,N_2347);
or U6314 (N_6314,N_1277,N_2760);
and U6315 (N_6315,N_3387,N_1270);
nor U6316 (N_6316,N_2324,N_3095);
nand U6317 (N_6317,N_4686,N_4906);
nand U6318 (N_6318,N_2105,N_663);
nand U6319 (N_6319,N_3220,N_1250);
and U6320 (N_6320,N_4448,N_3306);
nand U6321 (N_6321,N_1308,N_1520);
or U6322 (N_6322,N_3205,N_221);
or U6323 (N_6323,N_1942,N_3247);
and U6324 (N_6324,N_4029,N_4401);
and U6325 (N_6325,N_432,N_448);
nor U6326 (N_6326,N_4998,N_436);
and U6327 (N_6327,N_3312,N_2349);
or U6328 (N_6328,N_1375,N_549);
nand U6329 (N_6329,N_4244,N_2464);
nand U6330 (N_6330,N_2805,N_3083);
or U6331 (N_6331,N_2624,N_4375);
and U6332 (N_6332,N_2662,N_156);
or U6333 (N_6333,N_4873,N_2517);
and U6334 (N_6334,N_4586,N_3056);
nor U6335 (N_6335,N_804,N_3513);
and U6336 (N_6336,N_4799,N_352);
and U6337 (N_6337,N_92,N_4647);
xnor U6338 (N_6338,N_433,N_3719);
nor U6339 (N_6339,N_868,N_4008);
and U6340 (N_6340,N_1065,N_4542);
or U6341 (N_6341,N_859,N_112);
or U6342 (N_6342,N_3536,N_4791);
nor U6343 (N_6343,N_4974,N_1103);
nand U6344 (N_6344,N_2722,N_132);
nand U6345 (N_6345,N_1852,N_1813);
nand U6346 (N_6346,N_2532,N_4606);
or U6347 (N_6347,N_1978,N_1040);
and U6348 (N_6348,N_1725,N_2977);
nor U6349 (N_6349,N_4999,N_246);
nor U6350 (N_6350,N_4890,N_1171);
nand U6351 (N_6351,N_1938,N_3562);
nor U6352 (N_6352,N_840,N_4558);
nand U6353 (N_6353,N_1596,N_3464);
nor U6354 (N_6354,N_4085,N_4205);
and U6355 (N_6355,N_143,N_1591);
or U6356 (N_6356,N_1657,N_4835);
or U6357 (N_6357,N_148,N_3841);
and U6358 (N_6358,N_776,N_3786);
nor U6359 (N_6359,N_4846,N_2975);
or U6360 (N_6360,N_3501,N_1590);
nor U6361 (N_6361,N_2803,N_2816);
or U6362 (N_6362,N_3176,N_2264);
nand U6363 (N_6363,N_2695,N_69);
and U6364 (N_6364,N_1017,N_4655);
or U6365 (N_6365,N_26,N_490);
and U6366 (N_6366,N_4002,N_636);
nand U6367 (N_6367,N_1633,N_3626);
nor U6368 (N_6368,N_886,N_1287);
nor U6369 (N_6369,N_3426,N_795);
or U6370 (N_6370,N_3809,N_4222);
nor U6371 (N_6371,N_2762,N_1831);
xnor U6372 (N_6372,N_1307,N_1946);
xor U6373 (N_6373,N_3165,N_593);
or U6374 (N_6374,N_1201,N_2620);
nor U6375 (N_6375,N_1794,N_3865);
or U6376 (N_6376,N_896,N_974);
and U6377 (N_6377,N_1245,N_4172);
and U6378 (N_6378,N_2086,N_3580);
nand U6379 (N_6379,N_4382,N_2861);
nand U6380 (N_6380,N_445,N_1658);
nand U6381 (N_6381,N_3410,N_970);
nand U6382 (N_6382,N_3322,N_2013);
nor U6383 (N_6383,N_1787,N_2535);
nor U6384 (N_6384,N_4461,N_2712);
nor U6385 (N_6385,N_2823,N_1306);
or U6386 (N_6386,N_1795,N_1780);
nand U6387 (N_6387,N_1138,N_2557);
and U6388 (N_6388,N_2698,N_890);
or U6389 (N_6389,N_3914,N_4082);
or U6390 (N_6390,N_141,N_1800);
xnor U6391 (N_6391,N_3601,N_396);
nand U6392 (N_6392,N_3685,N_357);
nor U6393 (N_6393,N_1678,N_1051);
and U6394 (N_6394,N_2208,N_2418);
nand U6395 (N_6395,N_2669,N_1870);
nand U6396 (N_6396,N_4657,N_1098);
nand U6397 (N_6397,N_4501,N_3221);
nand U6398 (N_6398,N_3065,N_2414);
or U6399 (N_6399,N_802,N_4809);
nor U6400 (N_6400,N_403,N_2764);
nor U6401 (N_6401,N_1680,N_4705);
or U6402 (N_6402,N_3025,N_4343);
nor U6403 (N_6403,N_732,N_2563);
nor U6404 (N_6404,N_78,N_170);
nor U6405 (N_6405,N_415,N_4459);
and U6406 (N_6406,N_1234,N_2423);
nand U6407 (N_6407,N_3180,N_1918);
or U6408 (N_6408,N_669,N_3718);
nand U6409 (N_6409,N_270,N_1753);
nor U6410 (N_6410,N_2153,N_3393);
nand U6411 (N_6411,N_2836,N_2598);
and U6412 (N_6412,N_2787,N_3530);
or U6413 (N_6413,N_1061,N_1261);
and U6414 (N_6414,N_4766,N_2692);
and U6415 (N_6415,N_1434,N_603);
xnor U6416 (N_6416,N_308,N_905);
nor U6417 (N_6417,N_3484,N_820);
nand U6418 (N_6418,N_996,N_3950);
or U6419 (N_6419,N_4590,N_87);
and U6420 (N_6420,N_2852,N_3429);
nand U6421 (N_6421,N_191,N_1333);
nand U6422 (N_6422,N_4189,N_370);
or U6423 (N_6423,N_1462,N_105);
nand U6424 (N_6424,N_3172,N_3170);
and U6425 (N_6425,N_3693,N_1471);
nor U6426 (N_6426,N_772,N_858);
nor U6427 (N_6427,N_592,N_2668);
nor U6428 (N_6428,N_1013,N_1701);
and U6429 (N_6429,N_3682,N_1688);
nand U6430 (N_6430,N_679,N_3897);
nor U6431 (N_6431,N_2279,N_573);
nand U6432 (N_6432,N_230,N_2824);
nor U6433 (N_6433,N_4771,N_197);
and U6434 (N_6434,N_3551,N_4368);
nand U6435 (N_6435,N_4278,N_385);
nor U6436 (N_6436,N_4446,N_1401);
nand U6437 (N_6437,N_2040,N_4713);
or U6438 (N_6438,N_2550,N_1009);
and U6439 (N_6439,N_2946,N_4238);
nor U6440 (N_6440,N_3934,N_3396);
or U6441 (N_6441,N_2893,N_3024);
nor U6442 (N_6442,N_4762,N_1121);
or U6443 (N_6443,N_881,N_1336);
nand U6444 (N_6444,N_4022,N_3739);
and U6445 (N_6445,N_968,N_2617);
or U6446 (N_6446,N_575,N_1606);
xor U6447 (N_6447,N_2092,N_2175);
nor U6448 (N_6448,N_4337,N_1239);
or U6449 (N_6449,N_3478,N_4460);
or U6450 (N_6450,N_2652,N_1243);
nand U6451 (N_6451,N_2397,N_1057);
nor U6452 (N_6452,N_1407,N_4909);
and U6453 (N_6453,N_1841,N_1908);
nand U6454 (N_6454,N_2589,N_247);
or U6455 (N_6455,N_2903,N_1125);
or U6456 (N_6456,N_3961,N_564);
and U6457 (N_6457,N_418,N_1983);
and U6458 (N_6458,N_2935,N_2036);
nor U6459 (N_6459,N_1707,N_1939);
nand U6460 (N_6460,N_3015,N_2087);
nand U6461 (N_6461,N_2934,N_4472);
nor U6462 (N_6462,N_4966,N_3311);
or U6463 (N_6463,N_4546,N_532);
or U6464 (N_6464,N_2736,N_2741);
and U6465 (N_6465,N_1397,N_1664);
and U6466 (N_6466,N_287,N_1282);
nor U6467 (N_6467,N_3556,N_962);
and U6468 (N_6468,N_4674,N_3524);
nor U6469 (N_6469,N_2486,N_4961);
nor U6470 (N_6470,N_1311,N_1984);
and U6471 (N_6471,N_4621,N_988);
or U6472 (N_6472,N_2687,N_767);
nand U6473 (N_6473,N_3936,N_1213);
or U6474 (N_6474,N_4068,N_1861);
nor U6475 (N_6475,N_4792,N_1181);
or U6476 (N_6476,N_2940,N_581);
and U6477 (N_6477,N_4110,N_3952);
nand U6478 (N_6478,N_3763,N_349);
or U6479 (N_6479,N_3633,N_359);
or U6480 (N_6480,N_4681,N_29);
and U6481 (N_6481,N_286,N_2325);
nand U6482 (N_6482,N_3701,N_4152);
nand U6483 (N_6483,N_3791,N_4942);
nand U6484 (N_6484,N_1967,N_2190);
nand U6485 (N_6485,N_3009,N_703);
nor U6486 (N_6486,N_2181,N_2470);
nand U6487 (N_6487,N_1711,N_893);
nand U6488 (N_6488,N_3485,N_779);
nor U6489 (N_6489,N_2533,N_2345);
nand U6490 (N_6490,N_1693,N_40);
or U6491 (N_6491,N_4044,N_4916);
or U6492 (N_6492,N_1872,N_3645);
nand U6493 (N_6493,N_4289,N_3730);
nor U6494 (N_6494,N_2793,N_3802);
or U6495 (N_6495,N_4784,N_1609);
or U6496 (N_6496,N_4495,N_1025);
or U6497 (N_6497,N_360,N_515);
nor U6498 (N_6498,N_86,N_3157);
nor U6499 (N_6499,N_2116,N_987);
nand U6500 (N_6500,N_855,N_1750);
and U6501 (N_6501,N_3593,N_4660);
nand U6502 (N_6502,N_2440,N_260);
nor U6503 (N_6503,N_1637,N_2436);
and U6504 (N_6504,N_4505,N_1364);
nand U6505 (N_6505,N_1490,N_32);
and U6506 (N_6506,N_568,N_909);
and U6507 (N_6507,N_4323,N_2372);
and U6508 (N_6508,N_635,N_3103);
nor U6509 (N_6509,N_3691,N_2545);
nor U6510 (N_6510,N_3069,N_98);
or U6511 (N_6511,N_414,N_2973);
nand U6512 (N_6512,N_1502,N_1889);
and U6513 (N_6513,N_4120,N_806);
nor U6514 (N_6514,N_698,N_1374);
or U6515 (N_6515,N_591,N_2122);
or U6516 (N_6516,N_1754,N_2469);
nor U6517 (N_6517,N_787,N_4638);
nor U6518 (N_6518,N_3731,N_1265);
or U6519 (N_6519,N_3736,N_2409);
or U6520 (N_6520,N_2799,N_187);
and U6521 (N_6521,N_243,N_2400);
xnor U6522 (N_6522,N_4043,N_2297);
or U6523 (N_6523,N_212,N_3557);
or U6524 (N_6524,N_4415,N_4759);
or U6525 (N_6525,N_3560,N_4599);
nor U6526 (N_6526,N_1785,N_3071);
or U6527 (N_6527,N_2753,N_2327);
nor U6528 (N_6528,N_1094,N_1964);
nor U6529 (N_6529,N_4957,N_1531);
nand U6530 (N_6530,N_1176,N_1376);
and U6531 (N_6531,N_4815,N_1059);
or U6532 (N_6532,N_2511,N_1696);
nor U6533 (N_6533,N_3038,N_2356);
nor U6534 (N_6534,N_774,N_597);
nand U6535 (N_6535,N_1315,N_688);
and U6536 (N_6536,N_2326,N_1235);
nand U6537 (N_6537,N_3319,N_1575);
nand U6538 (N_6538,N_15,N_2337);
and U6539 (N_6539,N_861,N_232);
and U6540 (N_6540,N_1982,N_4250);
and U6541 (N_6541,N_4754,N_2588);
nor U6542 (N_6542,N_3499,N_1876);
nand U6543 (N_6543,N_4411,N_1624);
nand U6544 (N_6544,N_4099,N_18);
nand U6545 (N_6545,N_3388,N_70);
or U6546 (N_6546,N_1083,N_2361);
and U6547 (N_6547,N_3051,N_4689);
xnor U6548 (N_6548,N_3589,N_1557);
and U6549 (N_6549,N_1128,N_312);
nand U6550 (N_6550,N_3250,N_2967);
or U6551 (N_6551,N_1456,N_2551);
xnor U6552 (N_6552,N_563,N_1588);
nand U6553 (N_6553,N_517,N_3003);
and U6554 (N_6554,N_1452,N_2880);
nor U6555 (N_6555,N_2091,N_1744);
nor U6556 (N_6556,N_3992,N_1417);
nor U6557 (N_6557,N_4245,N_674);
nand U6558 (N_6558,N_1673,N_3193);
nand U6559 (N_6559,N_184,N_4322);
nor U6560 (N_6560,N_3362,N_1891);
nor U6561 (N_6561,N_2808,N_486);
and U6562 (N_6562,N_4316,N_3002);
and U6563 (N_6563,N_1210,N_3042);
and U6564 (N_6564,N_654,N_2537);
and U6565 (N_6565,N_4879,N_4315);
nand U6566 (N_6566,N_4994,N_3244);
and U6567 (N_6567,N_2848,N_3668);
nand U6568 (N_6568,N_4695,N_1997);
nand U6569 (N_6569,N_4369,N_2981);
nand U6570 (N_6570,N_4237,N_3432);
nor U6571 (N_6571,N_3274,N_4334);
or U6572 (N_6572,N_4617,N_4566);
nand U6573 (N_6573,N_4356,N_3013);
nor U6574 (N_6574,N_722,N_164);
nand U6575 (N_6575,N_3857,N_472);
and U6576 (N_6576,N_4126,N_4294);
nor U6577 (N_6577,N_2226,N_2610);
and U6578 (N_6578,N_1559,N_1854);
nand U6579 (N_6579,N_3872,N_3021);
nand U6580 (N_6580,N_2779,N_355);
nand U6581 (N_6581,N_4114,N_4325);
or U6582 (N_6582,N_4129,N_454);
nor U6583 (N_6583,N_140,N_4393);
or U6584 (N_6584,N_111,N_4521);
nor U6585 (N_6585,N_1971,N_469);
or U6586 (N_6586,N_1124,N_1405);
and U6587 (N_6587,N_2422,N_310);
or U6588 (N_6588,N_1075,N_2049);
nor U6589 (N_6589,N_2212,N_716);
and U6590 (N_6590,N_657,N_3799);
nor U6591 (N_6591,N_330,N_3655);
or U6592 (N_6592,N_3450,N_3917);
and U6593 (N_6593,N_1802,N_3029);
nand U6594 (N_6594,N_1746,N_516);
xnor U6595 (N_6595,N_3179,N_1263);
nor U6596 (N_6596,N_3446,N_4169);
or U6597 (N_6597,N_545,N_4884);
and U6598 (N_6598,N_1334,N_1199);
or U6599 (N_6599,N_4361,N_908);
and U6600 (N_6600,N_4196,N_3785);
nand U6601 (N_6601,N_1862,N_1012);
xor U6602 (N_6602,N_2393,N_3678);
nor U6603 (N_6603,N_3838,N_1188);
nand U6604 (N_6604,N_189,N_2906);
or U6605 (N_6605,N_2396,N_440);
and U6606 (N_6606,N_1454,N_2425);
nor U6607 (N_6607,N_4405,N_1383);
xor U6608 (N_6608,N_610,N_2515);
or U6609 (N_6609,N_1915,N_670);
nor U6610 (N_6610,N_1972,N_992);
nand U6611 (N_6611,N_2705,N_1031);
xor U6612 (N_6612,N_2783,N_1981);
nor U6613 (N_6613,N_4482,N_3080);
or U6614 (N_6614,N_3159,N_3207);
or U6615 (N_6615,N_1389,N_2619);
nor U6616 (N_6616,N_2706,N_135);
or U6617 (N_6617,N_3909,N_13);
nand U6618 (N_6618,N_3954,N_1183);
nand U6619 (N_6619,N_883,N_2690);
or U6620 (N_6620,N_4300,N_137);
or U6621 (N_6621,N_1344,N_2063);
and U6622 (N_6622,N_615,N_4572);
nor U6623 (N_6623,N_3199,N_3117);
or U6624 (N_6624,N_2606,N_1227);
nand U6625 (N_6625,N_2482,N_3115);
nand U6626 (N_6626,N_2830,N_4608);
nand U6627 (N_6627,N_2497,N_223);
and U6628 (N_6628,N_2513,N_529);
nand U6629 (N_6629,N_4953,N_1468);
or U6630 (N_6630,N_1072,N_2484);
nand U6631 (N_6631,N_1420,N_1342);
nor U6632 (N_6632,N_3317,N_2136);
and U6633 (N_6633,N_939,N_1379);
nand U6634 (N_6634,N_1400,N_2443);
and U6635 (N_6635,N_91,N_4596);
and U6636 (N_6636,N_3277,N_3913);
or U6637 (N_6637,N_316,N_3239);
and U6638 (N_6638,N_127,N_2209);
and U6639 (N_6639,N_691,N_1272);
and U6640 (N_6640,N_681,N_1217);
nand U6641 (N_6641,N_1464,N_1316);
nor U6642 (N_6642,N_4396,N_3090);
nand U6643 (N_6643,N_1781,N_1146);
nand U6644 (N_6644,N_2164,N_2976);
nor U6645 (N_6645,N_2964,N_4329);
nand U6646 (N_6646,N_4538,N_2247);
and U6647 (N_6647,N_4839,N_2658);
and U6648 (N_6648,N_4275,N_3650);
nor U6649 (N_6649,N_3452,N_727);
nor U6650 (N_6650,N_2918,N_2628);
or U6651 (N_6651,N_857,N_2616);
and U6652 (N_6652,N_554,N_3694);
and U6653 (N_6653,N_391,N_3959);
nand U6654 (N_6654,N_2794,N_1482);
nand U6655 (N_6655,N_1826,N_2518);
and U6656 (N_6656,N_505,N_833);
nor U6657 (N_6657,N_1002,N_1936);
and U6658 (N_6658,N_2174,N_4041);
nor U6659 (N_6659,N_3346,N_2645);
and U6660 (N_6660,N_4451,N_1156);
or U6661 (N_6661,N_2795,N_1745);
nor U6662 (N_6662,N_2125,N_499);
and U6663 (N_6663,N_3376,N_3246);
nand U6664 (N_6664,N_1724,N_2735);
nor U6665 (N_6665,N_1141,N_578);
nor U6666 (N_6666,N_2184,N_151);
and U6667 (N_6667,N_4210,N_3004);
nor U6668 (N_6668,N_120,N_2682);
or U6669 (N_6669,N_3459,N_1567);
nand U6670 (N_6670,N_4731,N_2599);
or U6671 (N_6671,N_3526,N_1177);
nand U6672 (N_6672,N_3722,N_172);
or U6673 (N_6673,N_661,N_2663);
or U6674 (N_6674,N_2851,N_3637);
nand U6675 (N_6675,N_379,N_3910);
and U6676 (N_6676,N_1622,N_453);
nand U6677 (N_6677,N_4528,N_496);
nor U6678 (N_6678,N_2407,N_4121);
nand U6679 (N_6679,N_2547,N_2261);
or U6680 (N_6680,N_320,N_4977);
and U6681 (N_6681,N_3488,N_3568);
and U6682 (N_6682,N_3770,N_2191);
and U6683 (N_6683,N_3862,N_2341);
and U6684 (N_6684,N_3893,N_3686);
nand U6685 (N_6685,N_841,N_1092);
and U6686 (N_6686,N_4209,N_4514);
nor U6687 (N_6687,N_3690,N_4010);
nor U6688 (N_6688,N_4352,N_4948);
or U6689 (N_6689,N_2770,N_3855);
nor U6690 (N_6690,N_2415,N_3171);
and U6691 (N_6691,N_2578,N_2287);
and U6692 (N_6692,N_2031,N_3970);
or U6693 (N_6693,N_631,N_1119);
nand U6694 (N_6694,N_637,N_3644);
or U6695 (N_6695,N_299,N_3707);
nand U6696 (N_6696,N_2737,N_1670);
nand U6697 (N_6697,N_2676,N_3323);
or U6698 (N_6698,N_67,N_1643);
nand U6699 (N_6699,N_4048,N_4725);
or U6700 (N_6700,N_2340,N_2594);
nand U6701 (N_6701,N_1260,N_2894);
and U6702 (N_6702,N_4733,N_319);
and U6703 (N_6703,N_3354,N_2514);
and U6704 (N_6704,N_3228,N_1446);
or U6705 (N_6705,N_3837,N_871);
or U6706 (N_6706,N_2553,N_2843);
and U6707 (N_6707,N_3030,N_867);
nor U6708 (N_6708,N_3774,N_1324);
or U6709 (N_6709,N_2858,N_4914);
and U6710 (N_6710,N_4123,N_3474);
and U6711 (N_6711,N_4908,N_271);
and U6712 (N_6712,N_4639,N_3262);
nor U6713 (N_6713,N_2456,N_1387);
and U6714 (N_6714,N_2740,N_1512);
nand U6715 (N_6715,N_4430,N_4398);
nand U6716 (N_6716,N_1406,N_2636);
nand U6717 (N_6717,N_1945,N_3810);
or U6718 (N_6718,N_4894,N_4672);
nor U6719 (N_6719,N_3962,N_3416);
nand U6720 (N_6720,N_2066,N_447);
nand U6721 (N_6721,N_4308,N_4306);
and U6722 (N_6722,N_2738,N_3634);
nand U6723 (N_6723,N_106,N_3167);
and U6724 (N_6724,N_4489,N_4926);
and U6725 (N_6725,N_3144,N_328);
or U6726 (N_6726,N_1064,N_84);
and U6727 (N_6727,N_550,N_4549);
and U6728 (N_6728,N_1715,N_2027);
and U6729 (N_6729,N_1077,N_1888);
nand U6730 (N_6730,N_444,N_3203);
and U6731 (N_6731,N_1491,N_3275);
nor U6732 (N_6732,N_4358,N_3566);
and U6733 (N_6733,N_1249,N_3628);
nor U6734 (N_6734,N_1474,N_1288);
nand U6735 (N_6735,N_4165,N_3461);
or U6736 (N_6736,N_3483,N_3336);
or U6737 (N_6737,N_3477,N_3006);
and U6738 (N_6738,N_1571,N_3261);
nor U6739 (N_6739,N_2353,N_2251);
and U6740 (N_6740,N_1225,N_277);
nand U6741 (N_6741,N_3776,N_102);
nand U6742 (N_6742,N_935,N_2642);
nand U6743 (N_6743,N_1386,N_4338);
nand U6744 (N_6744,N_1108,N_4328);
and U6745 (N_6745,N_4005,N_4710);
and U6746 (N_6746,N_2093,N_2831);
and U6747 (N_6747,N_4028,N_524);
nor U6748 (N_6748,N_1662,N_2323);
or U6749 (N_6749,N_4819,N_9);
nor U6750 (N_6750,N_2911,N_3057);
or U6751 (N_6751,N_1158,N_1373);
nor U6752 (N_6752,N_2315,N_850);
nand U6753 (N_6753,N_1111,N_3639);
nand U6754 (N_6754,N_3273,N_2983);
nor U6755 (N_6755,N_4050,N_1925);
nor U6756 (N_6756,N_2233,N_1582);
xor U6757 (N_6757,N_725,N_2835);
nor U6758 (N_6758,N_4938,N_1507);
nor U6759 (N_6759,N_4452,N_3482);
nor U6760 (N_6760,N_3569,N_4704);
or U6761 (N_6761,N_3425,N_569);
or U6762 (N_6762,N_1257,N_4458);
or U6763 (N_6763,N_4158,N_2899);
or U6764 (N_6764,N_1848,N_2528);
and U6765 (N_6765,N_1208,N_3046);
xor U6766 (N_6766,N_605,N_2954);
and U6767 (N_6767,N_1550,N_4979);
nor U6768 (N_6768,N_2014,N_558);
nor U6769 (N_6769,N_3210,N_2047);
nand U6770 (N_6770,N_4981,N_4327);
and U6771 (N_6771,N_1904,N_214);
nor U6772 (N_6772,N_2778,N_3625);
or U6773 (N_6773,N_1970,N_4441);
and U6774 (N_6774,N_3813,N_2901);
and U6775 (N_6775,N_1788,N_4012);
xnor U6776 (N_6776,N_1028,N_1241);
nand U6777 (N_6777,N_920,N_1170);
nand U6778 (N_6778,N_1910,N_547);
nor U6779 (N_6779,N_3611,N_2035);
nand U6780 (N_6780,N_2215,N_1683);
or U6781 (N_6781,N_4561,N_377);
nor U6782 (N_6782,N_3181,N_217);
xnor U6783 (N_6783,N_459,N_4551);
or U6784 (N_6784,N_4195,N_2554);
or U6785 (N_6785,N_2070,N_2145);
nor U6786 (N_6786,N_2339,N_1247);
or U6787 (N_6787,N_3687,N_2446);
nor U6788 (N_6788,N_936,N_1066);
nor U6789 (N_6789,N_2161,N_1346);
and U6790 (N_6790,N_752,N_2889);
or U6791 (N_6791,N_3453,N_1421);
and U6792 (N_6792,N_376,N_3302);
nand U6793 (N_6793,N_1953,N_2367);
nor U6794 (N_6794,N_793,N_446);
or U6795 (N_6795,N_3248,N_856);
nand U6796 (N_6796,N_4905,N_3906);
xnor U6797 (N_6797,N_2069,N_1363);
and U6798 (N_6798,N_3036,N_3364);
and U6799 (N_6799,N_702,N_2806);
or U6800 (N_6800,N_1992,N_3784);
and U6801 (N_6801,N_3400,N_4286);
nand U6802 (N_6802,N_2029,N_4039);
nand U6803 (N_6803,N_4061,N_4388);
nand U6804 (N_6804,N_2045,N_2170);
nand U6805 (N_6805,N_1224,N_4178);
nand U6806 (N_6806,N_4229,N_1524);
and U6807 (N_6807,N_1440,N_2103);
or U6808 (N_6808,N_4122,N_183);
nor U6809 (N_6809,N_3033,N_1223);
nor U6810 (N_6810,N_3310,N_3821);
nor U6811 (N_6811,N_678,N_3211);
and U6812 (N_6812,N_3084,N_3197);
nand U6813 (N_6813,N_4243,N_463);
or U6814 (N_6814,N_724,N_2194);
and U6815 (N_6815,N_2997,N_1388);
nand U6816 (N_6816,N_1279,N_206);
nor U6817 (N_6817,N_315,N_193);
and U6818 (N_6818,N_4379,N_3712);
or U6819 (N_6819,N_238,N_2681);
nor U6820 (N_6820,N_2784,N_2299);
nand U6821 (N_6821,N_458,N_1534);
or U6822 (N_6822,N_3571,N_399);
nor U6823 (N_6823,N_88,N_4475);
or U6824 (N_6824,N_4567,N_3111);
or U6825 (N_6825,N_1114,N_2885);
and U6826 (N_6826,N_1382,N_1775);
and U6827 (N_6827,N_2565,N_4153);
and U6828 (N_6828,N_2926,N_1024);
or U6829 (N_6829,N_544,N_2235);
nand U6830 (N_6830,N_751,N_3828);
nor U6831 (N_6831,N_4503,N_831);
and U6832 (N_6832,N_1281,N_2828);
xor U6833 (N_6833,N_3139,N_3119);
nor U6834 (N_6834,N_1175,N_261);
nor U6835 (N_6835,N_4108,N_4670);
nor U6836 (N_6836,N_3253,N_2562);
or U6837 (N_6837,N_2540,N_4076);
or U6838 (N_6838,N_1988,N_3178);
or U6839 (N_6839,N_2121,N_2204);
and U6840 (N_6840,N_3599,N_1004);
nand U6841 (N_6841,N_2369,N_2455);
nor U6842 (N_6842,N_2924,N_1749);
or U6843 (N_6843,N_667,N_4781);
nand U6844 (N_6844,N_1576,N_4);
and U6845 (N_6845,N_4406,N_1555);
nand U6846 (N_6846,N_4536,N_36);
and U6847 (N_6847,N_4486,N_1140);
nor U6848 (N_6848,N_4991,N_4612);
or U6849 (N_6849,N_4412,N_687);
and U6850 (N_6850,N_430,N_1742);
or U6851 (N_6851,N_3064,N_4616);
xnor U6852 (N_6852,N_3856,N_4730);
nand U6853 (N_6853,N_959,N_3752);
and U6854 (N_6854,N_4960,N_441);
nand U6855 (N_6855,N_3118,N_4026);
or U6856 (N_6856,N_2566,N_2807);
or U6857 (N_6857,N_1532,N_4518);
nor U6858 (N_6858,N_3481,N_3796);
nor U6859 (N_6859,N_2401,N_3699);
nand U6860 (N_6860,N_1414,N_1003);
or U6861 (N_6861,N_1182,N_155);
nor U6862 (N_6862,N_1869,N_4741);
and U6863 (N_6863,N_1611,N_542);
or U6864 (N_6864,N_613,N_468);
nor U6865 (N_6865,N_594,N_3008);
or U6866 (N_6866,N_3726,N_1726);
and U6867 (N_6867,N_178,N_1398);
nor U6868 (N_6868,N_1099,N_2301);
nor U6869 (N_6869,N_294,N_3660);
or U6870 (N_6870,N_1298,N_2050);
nand U6871 (N_6871,N_4729,N_4629);
and U6872 (N_6872,N_1761,N_1351);
or U6873 (N_6873,N_4850,N_717);
and U6874 (N_6874,N_4530,N_4249);
and U6875 (N_6875,N_3184,N_332);
or U6876 (N_6876,N_3462,N_2811);
nor U6877 (N_6877,N_4702,N_4714);
and U6878 (N_6878,N_264,N_4261);
and U6879 (N_6879,N_2773,N_1712);
or U6880 (N_6880,N_4400,N_3399);
or U6881 (N_6881,N_3546,N_201);
nor U6882 (N_6882,N_3577,N_2495);
nor U6883 (N_6883,N_3805,N_522);
nor U6884 (N_6884,N_4246,N_565);
nand U6885 (N_6885,N_491,N_2747);
nand U6886 (N_6886,N_634,N_3230);
and U6887 (N_6887,N_3465,N_1191);
nand U6888 (N_6888,N_1335,N_2259);
or U6889 (N_6889,N_523,N_3911);
nor U6890 (N_6890,N_3240,N_737);
or U6891 (N_6891,N_866,N_3217);
nor U6892 (N_6892,N_4554,N_1697);
nand U6893 (N_6893,N_4058,N_2419);
and U6894 (N_6894,N_3014,N_3706);
and U6895 (N_6895,N_944,N_2867);
and U6896 (N_6896,N_3674,N_2386);
or U6897 (N_6897,N_1459,N_4469);
nor U6898 (N_6898,N_1884,N_1251);
nor U6899 (N_6899,N_3891,N_3594);
nand U6900 (N_6900,N_4089,N_3471);
nand U6901 (N_6901,N_4211,N_2878);
nand U6902 (N_6902,N_4888,N_4183);
or U6903 (N_6903,N_233,N_2467);
or U6904 (N_6904,N_2195,N_682);
nor U6905 (N_6905,N_2640,N_4404);
or U6906 (N_6906,N_273,N_4284);
nand U6907 (N_6907,N_2451,N_3011);
or U6908 (N_6908,N_2404,N_3640);
nand U6909 (N_6909,N_4525,N_3997);
nand U6910 (N_6910,N_707,N_4239);
or U6911 (N_6911,N_2021,N_3476);
nor U6912 (N_6912,N_3555,N_4408);
nand U6913 (N_6913,N_1068,N_967);
nand U6914 (N_6914,N_393,N_2487);
and U6915 (N_6915,N_531,N_2549);
nor U6916 (N_6916,N_860,N_3984);
or U6917 (N_6917,N_3723,N_582);
xnor U6918 (N_6918,N_258,N_1636);
and U6919 (N_6919,N_3195,N_2348);
nor U6920 (N_6920,N_1580,N_4493);
or U6921 (N_6921,N_2516,N_3339);
nand U6922 (N_6922,N_4092,N_1730);
nor U6923 (N_6923,N_730,N_2399);
and U6924 (N_6924,N_300,N_1046);
or U6925 (N_6925,N_2019,N_1937);
nand U6926 (N_6926,N_4656,N_829);
nor U6927 (N_6927,N_4789,N_646);
nand U6928 (N_6928,N_4935,N_2492);
or U6929 (N_6929,N_1620,N_3422);
and U6930 (N_6930,N_2781,N_3045);
nand U6931 (N_6931,N_4683,N_61);
or U6932 (N_6932,N_3265,N_4562);
nand U6933 (N_6933,N_2128,N_4057);
or U6934 (N_6934,N_4937,N_2896);
or U6935 (N_6935,N_885,N_1853);
or U6936 (N_6936,N_2198,N_81);
nor U6937 (N_6937,N_467,N_3226);
or U6938 (N_6938,N_2004,N_1109);
nand U6939 (N_6939,N_624,N_2378);
or U6940 (N_6940,N_1871,N_144);
and U6941 (N_6941,N_2016,N_566);
nor U6942 (N_6942,N_2149,N_4071);
or U6943 (N_6943,N_4254,N_1086);
nor U6944 (N_6944,N_1535,N_4682);
or U6945 (N_6945,N_2439,N_1917);
nor U6946 (N_6946,N_794,N_2139);
nand U6947 (N_6947,N_283,N_4141);
or U6948 (N_6948,N_322,N_2667);
nor U6949 (N_6949,N_2570,N_1016);
nor U6950 (N_6950,N_510,N_4349);
nand U6951 (N_6951,N_4465,N_4468);
and U6952 (N_6952,N_1148,N_4004);
or U6953 (N_6953,N_2129,N_2529);
nor U6954 (N_6954,N_2350,N_1878);
and U6955 (N_6955,N_329,N_3887);
nand U6956 (N_6956,N_660,N_101);
or U6957 (N_6957,N_4609,N_4631);
and U6958 (N_6958,N_2278,N_3052);
and U6959 (N_6959,N_2897,N_4985);
and U6960 (N_6960,N_3600,N_609);
nand U6961 (N_6961,N_2826,N_3814);
nor U6962 (N_6962,N_3532,N_1021);
nand U6963 (N_6963,N_1283,N_1691);
or U6964 (N_6964,N_2990,N_1518);
or U6965 (N_6965,N_1592,N_1844);
nor U6966 (N_6966,N_3866,N_122);
nor U6967 (N_6967,N_2075,N_842);
or U6968 (N_6968,N_2252,N_4824);
nor U6969 (N_6969,N_3314,N_814);
or U6970 (N_6970,N_3116,N_3347);
nand U6971 (N_6971,N_2717,N_709);
and U6972 (N_6972,N_3280,N_659);
nor U6973 (N_6973,N_507,N_4310);
and U6974 (N_6974,N_3131,N_2150);
or U6975 (N_6975,N_4900,N_2083);
or U6976 (N_6976,N_4449,N_3054);
nor U6977 (N_6977,N_1603,N_4268);
nor U6978 (N_6978,N_2584,N_3331);
or U6979 (N_6979,N_2421,N_1839);
or U6980 (N_6980,N_3468,N_1758);
and U6981 (N_6981,N_3665,N_4203);
nor U6982 (N_6982,N_3822,N_2572);
or U6983 (N_6983,N_2290,N_1991);
and U6984 (N_6984,N_596,N_3938);
nand U6985 (N_6985,N_2955,N_876);
and U6986 (N_6986,N_3177,N_1493);
nor U6987 (N_6987,N_1060,N_693);
nor U6988 (N_6988,N_1702,N_35);
nand U6989 (N_6989,N_368,N_1665);
and U6990 (N_6990,N_3713,N_198);
nand U6991 (N_6991,N_2424,N_3098);
and U6992 (N_6992,N_4931,N_1445);
nor U6993 (N_6993,N_2211,N_2694);
nor U6994 (N_6994,N_3102,N_3829);
nand U6995 (N_6995,N_1667,N_2179);
or U6996 (N_6996,N_4764,N_2126);
or U6997 (N_6997,N_769,N_953);
or U6998 (N_6998,N_210,N_4234);
or U6999 (N_6999,N_4635,N_296);
and U7000 (N_7000,N_4363,N_2812);
nand U7001 (N_7001,N_1679,N_2285);
nor U7002 (N_7002,N_3133,N_56);
or U7003 (N_7003,N_37,N_895);
nand U7004 (N_7004,N_1276,N_1663);
nor U7005 (N_7005,N_4578,N_3487);
and U7006 (N_7006,N_3299,N_589);
or U7007 (N_7007,N_3135,N_2600);
or U7008 (N_7008,N_2895,N_3750);
nand U7009 (N_7009,N_3771,N_576);
nand U7010 (N_7010,N_473,N_1205);
nand U7011 (N_7011,N_1089,N_3136);
xnor U7012 (N_7012,N_2890,N_537);
and U7013 (N_7013,N_4780,N_4841);
or U7014 (N_7014,N_2898,N_4419);
nand U7015 (N_7015,N_1859,N_4896);
nand U7016 (N_7016,N_4949,N_647);
nand U7017 (N_7017,N_4003,N_162);
nor U7018 (N_7018,N_1246,N_4965);
or U7019 (N_7019,N_2296,N_3110);
nor U7020 (N_7020,N_710,N_4127);
and U7021 (N_7021,N_3271,N_2775);
nor U7022 (N_7022,N_4293,N_2904);
and U7023 (N_7023,N_699,N_2154);
nor U7024 (N_7024,N_658,N_2648);
and U7025 (N_7025,N_3545,N_3817);
nor U7026 (N_7026,N_1262,N_750);
and U7027 (N_7027,N_2257,N_2168);
nand U7028 (N_7028,N_4893,N_253);
and U7029 (N_7029,N_815,N_823);
and U7030 (N_7030,N_3941,N_869);
or U7031 (N_7031,N_3377,N_4790);
and U7032 (N_7032,N_2468,N_4912);
nand U7033 (N_7033,N_604,N_3017);
and U7034 (N_7034,N_1390,N_3918);
or U7035 (N_7035,N_656,N_2463);
nand U7036 (N_7036,N_4193,N_73);
nand U7037 (N_7037,N_4374,N_1681);
or U7038 (N_7038,N_1371,N_4073);
nand U7039 (N_7039,N_2697,N_356);
or U7040 (N_7040,N_2057,N_1821);
nand U7041 (N_7041,N_2227,N_2176);
or U7042 (N_7042,N_2871,N_428);
or U7043 (N_7043,N_4000,N_4955);
nor U7044 (N_7044,N_1706,N_4132);
or U7045 (N_7045,N_4421,N_2933);
nor U7046 (N_7046,N_2371,N_2166);
nor U7047 (N_7047,N_982,N_4299);
or U7048 (N_7048,N_2493,N_723);
nand U7049 (N_7049,N_1339,N_1451);
or U7050 (N_7050,N_3590,N_1759);
and U7051 (N_7051,N_4693,N_1549);
and U7052 (N_7052,N_3272,N_4564);
or U7053 (N_7053,N_4543,N_2430);
xnor U7054 (N_7054,N_2531,N_2373);
and U7055 (N_7055,N_4700,N_1581);
xor U7056 (N_7056,N_3642,N_3142);
nor U7057 (N_7057,N_4392,N_4802);
nor U7058 (N_7058,N_4555,N_3874);
or U7059 (N_7059,N_4054,N_1419);
nor U7060 (N_7060,N_3679,N_4962);
nand U7061 (N_7061,N_1539,N_4913);
xnor U7062 (N_7062,N_4601,N_827);
and U7063 (N_7063,N_2927,N_1593);
and U7064 (N_7064,N_4975,N_288);
nand U7065 (N_7065,N_1370,N_4500);
nand U7066 (N_7066,N_1536,N_4987);
or U7067 (N_7067,N_2143,N_3001);
or U7068 (N_7068,N_4823,N_4080);
and U7069 (N_7069,N_543,N_748);
nand U7070 (N_7070,N_3334,N_2394);
or U7071 (N_7071,N_176,N_2945);
nand U7072 (N_7072,N_3638,N_897);
or U7073 (N_7073,N_4776,N_502);
or U7074 (N_7074,N_2241,N_3946);
or U7075 (N_7075,N_3840,N_3216);
or U7076 (N_7076,N_4569,N_2120);
nor U7077 (N_7077,N_1353,N_19);
and U7078 (N_7078,N_3058,N_293);
or U7079 (N_7079,N_4223,N_3848);
xnor U7080 (N_7080,N_2255,N_1450);
nand U7081 (N_7081,N_3907,N_1033);
or U7082 (N_7082,N_4149,N_1134);
nor U7083 (N_7083,N_676,N_2384);
nor U7084 (N_7084,N_1784,N_3198);
xnor U7085 (N_7085,N_3448,N_1605);
or U7086 (N_7086,N_4046,N_276);
xnor U7087 (N_7087,N_3097,N_880);
and U7088 (N_7088,N_1129,N_225);
nor U7089 (N_7089,N_2197,N_4138);
and U7090 (N_7090,N_2237,N_2319);
and U7091 (N_7091,N_4745,N_3598);
and U7092 (N_7092,N_4031,N_2141);
and U7093 (N_7093,N_4177,N_1361);
or U7094 (N_7094,N_321,N_4381);
or U7095 (N_7095,N_4487,N_2772);
xor U7096 (N_7096,N_1144,N_4074);
nand U7097 (N_7097,N_2859,N_3900);
and U7098 (N_7098,N_1067,N_980);
nor U7099 (N_7099,N_2621,N_2909);
nor U7100 (N_7100,N_2082,N_307);
or U7101 (N_7101,N_2608,N_3467);
and U7102 (N_7102,N_3999,N_4242);
or U7103 (N_7103,N_3574,N_4857);
or U7104 (N_7104,N_3968,N_3318);
and U7105 (N_7105,N_347,N_4351);
nor U7106 (N_7106,N_2305,N_2199);
nor U7107 (N_7107,N_1372,N_79);
and U7108 (N_7108,N_4869,N_1329);
and U7109 (N_7109,N_975,N_1197);
nor U7110 (N_7110,N_1232,N_2380);
nand U7111 (N_7111,N_2248,N_4932);
nor U7112 (N_7112,N_4545,N_3344);
nor U7113 (N_7113,N_1242,N_2731);
or U7114 (N_7114,N_3764,N_2538);
or U7115 (N_7115,N_202,N_3795);
and U7116 (N_7116,N_65,N_2993);
nand U7117 (N_7117,N_3034,N_3578);
nand U7118 (N_7118,N_1751,N_1081);
nor U7119 (N_7119,N_1048,N_509);
and U7120 (N_7120,N_297,N_1881);
nand U7121 (N_7121,N_466,N_4197);
or U7122 (N_7122,N_3882,N_2131);
or U7123 (N_7123,N_4721,N_1530);
nand U7124 (N_7124,N_3263,N_4463);
nand U7125 (N_7125,N_2132,N_721);
nor U7126 (N_7126,N_4691,N_394);
nor U7127 (N_7127,N_4107,N_244);
or U7128 (N_7128,N_17,N_3604);
and U7129 (N_7129,N_3500,N_3703);
or U7130 (N_7130,N_3287,N_645);
or U7131 (N_7131,N_1913,N_1058);
nand U7132 (N_7132,N_4251,N_2754);
nor U7133 (N_7133,N_3629,N_1297);
nand U7134 (N_7134,N_3417,N_45);
or U7135 (N_7135,N_2466,N_3409);
or U7136 (N_7136,N_27,N_3000);
xnor U7137 (N_7137,N_4770,N_4434);
and U7138 (N_7138,N_3189,N_3149);
nand U7139 (N_7139,N_1516,N_2822);
nor U7140 (N_7140,N_3249,N_2750);
and U7141 (N_7141,N_397,N_3104);
nor U7142 (N_7142,N_2644,N_2948);
and U7143 (N_7143,N_3041,N_259);
and U7144 (N_7144,N_4007,N_4591);
nand U7145 (N_7145,N_3365,N_3390);
nand U7146 (N_7146,N_3218,N_2841);
or U7147 (N_7147,N_4719,N_97);
and U7148 (N_7148,N_175,N_1994);
nor U7149 (N_7149,N_1142,N_4052);
nor U7150 (N_7150,N_3405,N_1219);
nor U7151 (N_7151,N_2059,N_559);
nor U7152 (N_7152,N_2585,N_2672);
nor U7153 (N_7153,N_1030,N_1255);
nand U7154 (N_7154,N_3631,N_209);
nor U7155 (N_7155,N_2724,N_614);
and U7156 (N_7156,N_4255,N_100);
and U7157 (N_7157,N_3236,N_8);
nor U7158 (N_7158,N_759,N_1644);
and U7159 (N_7159,N_4473,N_2106);
nor U7160 (N_7160,N_4892,N_3127);
and U7161 (N_7161,N_3711,N_3976);
nor U7162 (N_7162,N_2220,N_2626);
or U7163 (N_7163,N_673,N_1666);
or U7164 (N_7164,N_1513,N_4722);
and U7165 (N_7165,N_3061,N_2298);
and U7166 (N_7166,N_4086,N_1762);
or U7167 (N_7167,N_362,N_2020);
nand U7168 (N_7168,N_3647,N_4814);
nor U7169 (N_7169,N_1123,N_1486);
or U7170 (N_7170,N_1814,N_1165);
nor U7171 (N_7171,N_3162,N_2377);
or U7172 (N_7172,N_4490,N_1722);
nor U7173 (N_7173,N_2855,N_915);
nand U7174 (N_7174,N_1731,N_2539);
or U7175 (N_7175,N_1710,N_3366);
nor U7176 (N_7176,N_2661,N_2498);
nor U7177 (N_7177,N_3412,N_3978);
or U7178 (N_7178,N_1153,N_2200);
xor U7179 (N_7179,N_96,N_3243);
and U7180 (N_7180,N_3870,N_4715);
or U7181 (N_7181,N_4967,N_4982);
or U7182 (N_7182,N_1465,N_4594);
or U7183 (N_7183,N_4155,N_1488);
or U7184 (N_7184,N_3635,N_1985);
nand U7185 (N_7185,N_3662,N_1070);
nand U7186 (N_7186,N_3132,N_2686);
or U7187 (N_7187,N_4150,N_3892);
nand U7188 (N_7188,N_309,N_1597);
and U7189 (N_7189,N_1899,N_617);
nand U7190 (N_7190,N_1209,N_41);
and U7191 (N_7191,N_1717,N_1415);
xnor U7192 (N_7192,N_4131,N_4342);
or U7193 (N_7193,N_1043,N_2729);
nand U7194 (N_7194,N_1027,N_1052);
nand U7195 (N_7195,N_4826,N_778);
or U7196 (N_7196,N_3609,N_4767);
nand U7197 (N_7197,N_2863,N_1830);
and U7198 (N_7198,N_1095,N_1008);
nor U7199 (N_7199,N_4679,N_410);
xor U7200 (N_7200,N_2763,N_1392);
or U7201 (N_7201,N_4100,N_4992);
nor U7202 (N_7202,N_1947,N_4556);
and U7203 (N_7203,N_2354,N_3335);
and U7204 (N_7204,N_2985,N_760);
nand U7205 (N_7205,N_2882,N_2582);
or U7206 (N_7206,N_4414,N_1868);
and U7207 (N_7207,N_4533,N_3398);
and U7208 (N_7208,N_2405,N_4096);
and U7209 (N_7209,N_1703,N_4848);
or U7210 (N_7210,N_3761,N_4016);
nor U7211 (N_7211,N_219,N_1618);
nand U7212 (N_7212,N_784,N_4580);
nand U7213 (N_7213,N_4807,N_3570);
or U7214 (N_7214,N_66,N_1584);
and U7215 (N_7215,N_4467,N_919);
xnor U7216 (N_7216,N_4847,N_1948);
nand U7217 (N_7217,N_4863,N_849);
xor U7218 (N_7218,N_3523,N_644);
nand U7219 (N_7219,N_4875,N_2715);
or U7220 (N_7220,N_612,N_251);
or U7221 (N_7221,N_146,N_4492);
nor U7222 (N_7222,N_1080,N_358);
xnor U7223 (N_7223,N_1473,N_1736);
nand U7224 (N_7224,N_1675,N_3792);
nor U7225 (N_7225,N_1195,N_1457);
or U7226 (N_7226,N_2703,N_2994);
nor U7227 (N_7227,N_4853,N_3953);
and U7228 (N_7228,N_372,N_1368);
or U7229 (N_7229,N_2454,N_2960);
nor U7230 (N_7230,N_906,N_325);
nor U7231 (N_7231,N_4972,N_1087);
or U7232 (N_7232,N_3109,N_1791);
nand U7233 (N_7233,N_2507,N_4431);
xnor U7234 (N_7234,N_3370,N_4668);
xnor U7235 (N_7235,N_2521,N_3284);
and U7236 (N_7236,N_2968,N_431);
and U7237 (N_7237,N_567,N_902);
and U7238 (N_7238,N_1286,N_3141);
or U7239 (N_7239,N_2119,N_425);
nor U7240 (N_7240,N_3916,N_2922);
nor U7241 (N_7241,N_4372,N_799);
or U7242 (N_7242,N_2886,N_4818);
nand U7243 (N_7243,N_2146,N_2596);
nand U7244 (N_7244,N_1827,N_3547);
and U7245 (N_7245,N_411,N_1921);
or U7246 (N_7246,N_1866,N_2991);
or U7247 (N_7247,N_4706,N_2110);
or U7248 (N_7248,N_4232,N_822);
or U7249 (N_7249,N_2017,N_3201);
nor U7250 (N_7250,N_2180,N_3885);
or U7251 (N_7251,N_1053,N_4646);
and U7252 (N_7252,N_1528,N_3192);
or U7253 (N_7253,N_719,N_284);
or U7254 (N_7254,N_268,N_2254);
nand U7255 (N_7255,N_2196,N_4357);
nor U7256 (N_7256,N_3120,N_1404);
nor U7257 (N_7257,N_3143,N_736);
nand U7258 (N_7258,N_4457,N_1408);
and U7259 (N_7259,N_3995,N_579);
nand U7260 (N_7260,N_3832,N_2137);
or U7261 (N_7261,N_3539,N_427);
nand U7262 (N_7262,N_501,N_694);
nand U7263 (N_7263,N_2614,N_1808);
nor U7264 (N_7264,N_4384,N_1385);
nor U7265 (N_7265,N_954,N_4810);
nand U7266 (N_7266,N_3896,N_685);
xnor U7267 (N_7267,N_2368,N_797);
or U7268 (N_7268,N_927,N_904);
nand U7269 (N_7269,N_4319,N_884);
and U7270 (N_7270,N_808,N_1704);
or U7271 (N_7271,N_2605,N_1672);
nand U7272 (N_7272,N_1563,N_2133);
nor U7273 (N_7273,N_4365,N_2358);
or U7274 (N_7274,N_4176,N_4009);
nor U7275 (N_7275,N_4864,N_1190);
nor U7276 (N_7276,N_2646,N_2592);
nand U7277 (N_7277,N_3441,N_651);
and U7278 (N_7278,N_4539,N_1857);
nor U7279 (N_7279,N_3439,N_985);
nand U7280 (N_7280,N_2067,N_416);
or U7281 (N_7281,N_2144,N_1630);
and U7282 (N_7282,N_546,N_2680);
and U7283 (N_7283,N_4305,N_3846);
nand U7284 (N_7284,N_252,N_1147);
nor U7285 (N_7285,N_3741,N_3106);
and U7286 (N_7286,N_4861,N_3494);
nor U7287 (N_7287,N_4034,N_1760);
and U7288 (N_7288,N_57,N_2113);
nor U7289 (N_7289,N_3614,N_2272);
nand U7290 (N_7290,N_4439,N_2080);
and U7291 (N_7291,N_1366,N_3301);
nand U7292 (N_7292,N_4124,N_1453);
nand U7293 (N_7293,N_4330,N_4817);
or U7294 (N_7294,N_932,N_1463);
or U7295 (N_7295,N_535,N_2618);
nor U7296 (N_7296,N_929,N_2438);
nand U7297 (N_7297,N_818,N_4455);
nand U7298 (N_7298,N_1285,N_4550);
and U7299 (N_7299,N_1629,N_585);
and U7300 (N_7300,N_548,N_4302);
nand U7301 (N_7301,N_666,N_983);
or U7302 (N_7302,N_2002,N_819);
or U7303 (N_7303,N_4867,N_185);
nor U7304 (N_7304,N_4225,N_1585);
and U7305 (N_7305,N_1091,N_2820);
nand U7306 (N_7306,N_2130,N_4166);
nor U7307 (N_7307,N_482,N_2998);
nor U7308 (N_7308,N_71,N_846);
xnor U7309 (N_7309,N_1979,N_2503);
nand U7310 (N_7310,N_3096,N_166);
and U7311 (N_7311,N_1240,N_2387);
nor U7312 (N_7312,N_1309,N_1423);
or U7313 (N_7313,N_4466,N_4442);
nor U7314 (N_7314,N_2962,N_773);
and U7315 (N_7315,N_1765,N_977);
or U7316 (N_7316,N_729,N_2346);
nand U7317 (N_7317,N_2649,N_1797);
or U7318 (N_7318,N_4151,N_2003);
and U7319 (N_7319,N_99,N_4886);
and U7320 (N_7320,N_798,N_93);
and U7321 (N_7321,N_4788,N_346);
or U7322 (N_7322,N_1429,N_4986);
and U7323 (N_7323,N_3125,N_4281);
and U7324 (N_7324,N_1211,N_3063);
nor U7325 (N_7325,N_3550,N_2963);
or U7326 (N_7326,N_2185,N_3268);
and U7327 (N_7327,N_2691,N_4941);
nand U7328 (N_7328,N_2102,N_3010);
nor U7329 (N_7329,N_4066,N_4450);
nand U7330 (N_7330,N_204,N_2713);
nand U7331 (N_7331,N_2655,N_4304);
nor U7332 (N_7332,N_3372,N_236);
nand U7333 (N_7333,N_1172,N_541);
and U7334 (N_7334,N_2839,N_4436);
xnor U7335 (N_7335,N_2966,N_2061);
and U7336 (N_7336,N_2159,N_1769);
nor U7337 (N_7337,N_1856,N_4018);
or U7338 (N_7338,N_266,N_282);
nor U7339 (N_7339,N_588,N_3245);
nor U7340 (N_7340,N_2868,N_1035);
and U7341 (N_7341,N_2342,N_1654);
nor U7342 (N_7342,N_4435,N_2217);
xor U7343 (N_7343,N_4757,N_2403);
nand U7344 (N_7344,N_810,N_1472);
or U7345 (N_7345,N_4947,N_3528);
or U7346 (N_7346,N_374,N_461);
or U7347 (N_7347,N_3378,N_4397);
nand U7348 (N_7348,N_22,N_1347);
and U7349 (N_7349,N_1071,N_2864);
and U7350 (N_7350,N_1687,N_188);
nand U7351 (N_7351,N_4624,N_89);
and U7352 (N_7352,N_3152,N_1621);
and U7353 (N_7353,N_1275,N_1136);
or U7354 (N_7354,N_1578,N_1772);
and U7355 (N_7355,N_4726,N_3489);
or U7356 (N_7356,N_4756,N_2379);
nand U7357 (N_7357,N_2427,N_1521);
and U7358 (N_7358,N_4851,N_4640);
and U7359 (N_7359,N_3958,N_2318);
nand U7360 (N_7360,N_404,N_1974);
and U7361 (N_7361,N_3902,N_4512);
nand U7362 (N_7362,N_3787,N_3512);
or U7363 (N_7363,N_2459,N_2671);
and U7364 (N_7364,N_3613,N_633);
nor U7365 (N_7365,N_2548,N_2860);
and U7366 (N_7366,N_817,N_1825);
and U7367 (N_7367,N_2581,N_1200);
nor U7368 (N_7368,N_2856,N_2160);
nand U7369 (N_7369,N_4060,N_3782);
or U7370 (N_7370,N_4136,N_3394);
or U7371 (N_7371,N_4852,N_4212);
nand U7372 (N_7372,N_3493,N_1006);
or U7373 (N_7373,N_4386,N_3925);
and U7374 (N_7374,N_113,N_910);
or U7375 (N_7375,N_3213,N_3194);
and U7376 (N_7376,N_2303,N_4174);
or U7377 (N_7377,N_2576,N_479);
and U7378 (N_7378,N_3504,N_3714);
and U7379 (N_7379,N_4552,N_901);
nor U7380 (N_7380,N_2073,N_250);
or U7381 (N_7381,N_1302,N_2932);
or U7382 (N_7382,N_4643,N_2292);
nor U7383 (N_7383,N_4808,N_749);
or U7384 (N_7384,N_389,N_2041);
and U7385 (N_7385,N_199,N_1779);
or U7386 (N_7386,N_3414,N_4488);
xnor U7387 (N_7387,N_2530,N_2483);
and U7388 (N_7388,N_4842,N_3413);
nand U7389 (N_7389,N_412,N_2534);
nand U7390 (N_7390,N_1163,N_4326);
and U7391 (N_7391,N_2395,N_442);
or U7392 (N_7392,N_335,N_4765);
nand U7393 (N_7393,N_4910,N_2568);
nand U7394 (N_7394,N_2877,N_4188);
and U7395 (N_7395,N_0,N_2406);
or U7396 (N_7396,N_1659,N_4447);
nand U7397 (N_7397,N_152,N_133);
or U7398 (N_7398,N_3361,N_2508);
or U7399 (N_7399,N_3169,N_2625);
nor U7400 (N_7400,N_1897,N_3597);
nor U7401 (N_7401,N_2431,N_813);
nand U7402 (N_7402,N_1564,N_4453);
and U7403 (N_7403,N_1509,N_894);
nor U7404 (N_7404,N_1641,N_2914);
or U7405 (N_7405,N_4820,N_4020);
nand U7406 (N_7406,N_1358,N_2331);
nand U7407 (N_7407,N_3890,N_912);
and U7408 (N_7408,N_513,N_2246);
nand U7409 (N_7409,N_4816,N_3092);
nor U7410 (N_7410,N_3521,N_3191);
and U7411 (N_7411,N_1244,N_2943);
and U7412 (N_7412,N_1807,N_3497);
nor U7413 (N_7413,N_4187,N_1877);
or U7414 (N_7414,N_4106,N_2138);
or U7415 (N_7415,N_3094,N_4081);
nand U7416 (N_7416,N_1506,N_955);
and U7417 (N_7417,N_3511,N_1959);
nand U7418 (N_7418,N_341,N_1796);
nand U7419 (N_7419,N_1763,N_2307);
nor U7420 (N_7420,N_4443,N_2756);
nand U7421 (N_7421,N_844,N_2000);
and U7422 (N_7422,N_2094,N_1708);
xnor U7423 (N_7423,N_1395,N_1189);
nor U7424 (N_7424,N_3673,N_938);
or U7425 (N_7425,N_1127,N_3447);
and U7426 (N_7426,N_302,N_2696);
and U7427 (N_7427,N_1348,N_3411);
or U7428 (N_7428,N_3990,N_2684);
and U7429 (N_7429,N_429,N_2193);
or U7430 (N_7430,N_3072,N_195);
and U7431 (N_7431,N_4509,N_16);
and U7432 (N_7432,N_1221,N_2214);
and U7433 (N_7433,N_4113,N_4148);
nor U7434 (N_7434,N_4740,N_3427);
and U7435 (N_7435,N_4291,N_556);
or U7436 (N_7436,N_4019,N_1541);
nor U7437 (N_7437,N_3652,N_4499);
or U7438 (N_7438,N_4659,N_1185);
and U7439 (N_7439,N_1113,N_768);
nand U7440 (N_7440,N_4427,N_4649);
and U7441 (N_7441,N_665,N_4577);
nand U7442 (N_7442,N_2313,N_2382);
or U7443 (N_7443,N_1481,N_4836);
nand U7444 (N_7444,N_2140,N_3227);
or U7445 (N_7445,N_3349,N_525);
or U7446 (N_7446,N_1635,N_119);
nor U7447 (N_7447,N_4045,N_1116);
or U7448 (N_7448,N_598,N_4157);
nand U7449 (N_7449,N_1805,N_3676);
or U7450 (N_7450,N_1919,N_640);
nand U7451 (N_7451,N_2389,N_1966);
and U7452 (N_7452,N_4951,N_2025);
nand U7453 (N_7453,N_2711,N_4880);
and U7454 (N_7454,N_3728,N_3986);
nand U7455 (N_7455,N_2187,N_3456);
or U7456 (N_7456,N_371,N_1554);
nand U7457 (N_7457,N_1164,N_3222);
or U7458 (N_7458,N_4063,N_4480);
nand U7459 (N_7459,N_790,N_33);
nand U7460 (N_7460,N_4313,N_623);
nor U7461 (N_7461,N_395,N_2552);
and U7462 (N_7462,N_3212,N_2905);
nor U7463 (N_7463,N_2224,N_1864);
or U7464 (N_7464,N_3937,N_916);
or U7465 (N_7465,N_2338,N_4821);
or U7466 (N_7466,N_3742,N_2546);
nand U7467 (N_7467,N_3697,N_3018);
and U7468 (N_7468,N_2664,N_1084);
and U7469 (N_7469,N_1259,N_2580);
nand U7470 (N_7470,N_4191,N_997);
nand U7471 (N_7471,N_1359,N_3186);
nand U7472 (N_7472,N_2228,N_1186);
nand U7473 (N_7473,N_413,N_4604);
or U7474 (N_7474,N_3505,N_2112);
or U7475 (N_7475,N_2714,N_192);
nor U7476 (N_7476,N_1475,N_3289);
and U7477 (N_7477,N_761,N_2702);
nor U7478 (N_7478,N_1594,N_4650);
and U7479 (N_7479,N_3028,N_2510);
or U7480 (N_7480,N_1980,N_4720);
and U7481 (N_7481,N_755,N_4877);
nor U7482 (N_7482,N_3734,N_3899);
or U7483 (N_7483,N_2491,N_4707);
nor U7484 (N_7484,N_4181,N_4830);
and U7485 (N_7485,N_4785,N_1764);
and U7486 (N_7486,N_2253,N_1699);
or U7487 (N_7487,N_3820,N_2941);
nand U7488 (N_7488,N_64,N_971);
nor U7489 (N_7489,N_171,N_2500);
and U7490 (N_7490,N_1253,N_4462);
nand U7491 (N_7491,N_4663,N_551);
nor U7492 (N_7492,N_786,N_2118);
nand U7493 (N_7493,N_3382,N_4904);
and U7494 (N_7494,N_2613,N_4684);
or U7495 (N_7495,N_50,N_2734);
and U7496 (N_7496,N_4793,N_227);
and U7497 (N_7497,N_4573,N_4833);
and U7498 (N_7498,N_4997,N_2370);
nor U7499 (N_7499,N_4866,N_1729);
nor U7500 (N_7500,N_1299,N_1925);
or U7501 (N_7501,N_1945,N_2363);
or U7502 (N_7502,N_1831,N_4980);
and U7503 (N_7503,N_2632,N_3652);
and U7504 (N_7504,N_306,N_1524);
nor U7505 (N_7505,N_928,N_2747);
nor U7506 (N_7506,N_192,N_4161);
nor U7507 (N_7507,N_3153,N_1572);
and U7508 (N_7508,N_1191,N_4218);
nor U7509 (N_7509,N_3479,N_4824);
nand U7510 (N_7510,N_4225,N_1540);
and U7511 (N_7511,N_4685,N_1585);
and U7512 (N_7512,N_3882,N_326);
and U7513 (N_7513,N_556,N_4849);
nor U7514 (N_7514,N_3214,N_2013);
nor U7515 (N_7515,N_2323,N_4861);
or U7516 (N_7516,N_2638,N_2560);
and U7517 (N_7517,N_2993,N_4740);
xnor U7518 (N_7518,N_1648,N_2701);
or U7519 (N_7519,N_1471,N_2299);
nand U7520 (N_7520,N_1301,N_2585);
and U7521 (N_7521,N_1818,N_2791);
or U7522 (N_7522,N_4687,N_1914);
or U7523 (N_7523,N_442,N_2839);
nor U7524 (N_7524,N_1619,N_4622);
nor U7525 (N_7525,N_740,N_1182);
and U7526 (N_7526,N_3919,N_3862);
or U7527 (N_7527,N_124,N_2120);
or U7528 (N_7528,N_1575,N_3391);
or U7529 (N_7529,N_2641,N_2727);
xor U7530 (N_7530,N_4658,N_4833);
nor U7531 (N_7531,N_1939,N_1191);
nor U7532 (N_7532,N_4964,N_2696);
and U7533 (N_7533,N_4548,N_4307);
or U7534 (N_7534,N_1349,N_119);
and U7535 (N_7535,N_4005,N_4711);
nand U7536 (N_7536,N_1905,N_4827);
and U7537 (N_7537,N_2867,N_3433);
and U7538 (N_7538,N_193,N_2138);
nor U7539 (N_7539,N_1770,N_699);
nor U7540 (N_7540,N_3403,N_3901);
nor U7541 (N_7541,N_3773,N_4026);
nor U7542 (N_7542,N_2446,N_3603);
nor U7543 (N_7543,N_804,N_1580);
or U7544 (N_7544,N_162,N_4820);
and U7545 (N_7545,N_4713,N_2670);
nor U7546 (N_7546,N_2275,N_2836);
or U7547 (N_7547,N_2348,N_2799);
nand U7548 (N_7548,N_2325,N_1284);
nor U7549 (N_7549,N_1726,N_4805);
or U7550 (N_7550,N_2015,N_1907);
nand U7551 (N_7551,N_68,N_2932);
nor U7552 (N_7552,N_1783,N_1201);
and U7553 (N_7553,N_1499,N_2563);
xor U7554 (N_7554,N_2024,N_2780);
or U7555 (N_7555,N_535,N_2842);
nand U7556 (N_7556,N_4353,N_839);
or U7557 (N_7557,N_2599,N_3499);
nand U7558 (N_7558,N_4255,N_3125);
nor U7559 (N_7559,N_1576,N_3458);
nand U7560 (N_7560,N_370,N_277);
nor U7561 (N_7561,N_2822,N_4352);
nand U7562 (N_7562,N_2420,N_1829);
nand U7563 (N_7563,N_1646,N_2900);
nand U7564 (N_7564,N_1316,N_2279);
nand U7565 (N_7565,N_2938,N_1534);
and U7566 (N_7566,N_4804,N_4347);
or U7567 (N_7567,N_3230,N_2031);
nor U7568 (N_7568,N_2147,N_2380);
and U7569 (N_7569,N_3900,N_4849);
nor U7570 (N_7570,N_3393,N_1467);
nor U7571 (N_7571,N_3224,N_2375);
and U7572 (N_7572,N_1356,N_1378);
nor U7573 (N_7573,N_2912,N_1071);
or U7574 (N_7574,N_1714,N_4984);
or U7575 (N_7575,N_4508,N_1165);
nand U7576 (N_7576,N_4363,N_4021);
nand U7577 (N_7577,N_883,N_766);
xor U7578 (N_7578,N_4314,N_4196);
and U7579 (N_7579,N_3466,N_2329);
nand U7580 (N_7580,N_1783,N_3769);
or U7581 (N_7581,N_2575,N_1278);
xnor U7582 (N_7582,N_1926,N_259);
nor U7583 (N_7583,N_3089,N_1663);
nand U7584 (N_7584,N_3604,N_535);
and U7585 (N_7585,N_4635,N_1877);
nand U7586 (N_7586,N_2511,N_1961);
nand U7587 (N_7587,N_2261,N_2468);
or U7588 (N_7588,N_4010,N_2214);
nor U7589 (N_7589,N_4668,N_2850);
nor U7590 (N_7590,N_4180,N_669);
nand U7591 (N_7591,N_4923,N_4728);
and U7592 (N_7592,N_1903,N_4656);
or U7593 (N_7593,N_3496,N_4752);
xor U7594 (N_7594,N_4225,N_3749);
nand U7595 (N_7595,N_347,N_433);
nor U7596 (N_7596,N_2890,N_1348);
nand U7597 (N_7597,N_41,N_630);
nand U7598 (N_7598,N_4157,N_2464);
nor U7599 (N_7599,N_3469,N_4509);
or U7600 (N_7600,N_3808,N_2987);
and U7601 (N_7601,N_2080,N_2926);
nor U7602 (N_7602,N_2015,N_1638);
or U7603 (N_7603,N_3096,N_704);
and U7604 (N_7604,N_3062,N_4471);
or U7605 (N_7605,N_1177,N_1314);
nand U7606 (N_7606,N_1206,N_3387);
and U7607 (N_7607,N_3286,N_3511);
nand U7608 (N_7608,N_2171,N_3094);
nand U7609 (N_7609,N_377,N_819);
and U7610 (N_7610,N_2527,N_1630);
and U7611 (N_7611,N_4750,N_193);
nor U7612 (N_7612,N_3338,N_970);
nand U7613 (N_7613,N_452,N_3086);
nor U7614 (N_7614,N_743,N_2692);
nor U7615 (N_7615,N_2646,N_300);
or U7616 (N_7616,N_3258,N_3308);
and U7617 (N_7617,N_4821,N_4316);
or U7618 (N_7618,N_1100,N_276);
nand U7619 (N_7619,N_1462,N_4970);
nor U7620 (N_7620,N_698,N_263);
and U7621 (N_7621,N_3491,N_3171);
and U7622 (N_7622,N_14,N_434);
nor U7623 (N_7623,N_233,N_3857);
or U7624 (N_7624,N_3179,N_3549);
nand U7625 (N_7625,N_3045,N_2230);
nand U7626 (N_7626,N_60,N_1525);
nand U7627 (N_7627,N_215,N_3753);
nand U7628 (N_7628,N_1337,N_4659);
nand U7629 (N_7629,N_4994,N_4086);
nor U7630 (N_7630,N_4646,N_4338);
nand U7631 (N_7631,N_4294,N_3719);
and U7632 (N_7632,N_3869,N_866);
nor U7633 (N_7633,N_4230,N_4511);
nand U7634 (N_7634,N_4870,N_694);
and U7635 (N_7635,N_4764,N_3599);
nand U7636 (N_7636,N_904,N_1377);
nor U7637 (N_7637,N_4366,N_3078);
nor U7638 (N_7638,N_3312,N_3871);
and U7639 (N_7639,N_4361,N_2041);
nor U7640 (N_7640,N_4832,N_696);
nand U7641 (N_7641,N_3246,N_2854);
nor U7642 (N_7642,N_2545,N_3444);
nand U7643 (N_7643,N_831,N_1412);
or U7644 (N_7644,N_1115,N_2465);
and U7645 (N_7645,N_2671,N_2654);
and U7646 (N_7646,N_3612,N_1842);
nor U7647 (N_7647,N_3892,N_537);
or U7648 (N_7648,N_1472,N_3077);
or U7649 (N_7649,N_524,N_2548);
nand U7650 (N_7650,N_1967,N_2510);
and U7651 (N_7651,N_2999,N_265);
nand U7652 (N_7652,N_2598,N_1294);
nor U7653 (N_7653,N_2063,N_4489);
nand U7654 (N_7654,N_1079,N_901);
and U7655 (N_7655,N_553,N_1546);
nor U7656 (N_7656,N_2236,N_4914);
nor U7657 (N_7657,N_875,N_2514);
nand U7658 (N_7658,N_2541,N_4882);
nor U7659 (N_7659,N_2646,N_1711);
and U7660 (N_7660,N_2861,N_871);
nor U7661 (N_7661,N_2282,N_1576);
nor U7662 (N_7662,N_4496,N_404);
nor U7663 (N_7663,N_480,N_1726);
nand U7664 (N_7664,N_4041,N_37);
and U7665 (N_7665,N_597,N_277);
and U7666 (N_7666,N_2372,N_1561);
nor U7667 (N_7667,N_350,N_1670);
nand U7668 (N_7668,N_3002,N_3918);
nand U7669 (N_7669,N_253,N_3271);
nand U7670 (N_7670,N_4611,N_2456);
and U7671 (N_7671,N_3953,N_3371);
nor U7672 (N_7672,N_753,N_849);
and U7673 (N_7673,N_3607,N_24);
nand U7674 (N_7674,N_3324,N_1263);
and U7675 (N_7675,N_4976,N_1074);
and U7676 (N_7676,N_967,N_670);
and U7677 (N_7677,N_2012,N_4303);
nor U7678 (N_7678,N_1016,N_1997);
nor U7679 (N_7679,N_578,N_4727);
and U7680 (N_7680,N_1034,N_2969);
or U7681 (N_7681,N_1489,N_2982);
nor U7682 (N_7682,N_51,N_1420);
and U7683 (N_7683,N_2067,N_3435);
or U7684 (N_7684,N_2639,N_1740);
nor U7685 (N_7685,N_4842,N_2062);
and U7686 (N_7686,N_1494,N_2350);
nor U7687 (N_7687,N_932,N_1476);
nand U7688 (N_7688,N_4938,N_2391);
or U7689 (N_7689,N_2116,N_103);
nor U7690 (N_7690,N_3716,N_3123);
xnor U7691 (N_7691,N_1261,N_3737);
nor U7692 (N_7692,N_693,N_2347);
and U7693 (N_7693,N_3370,N_2047);
or U7694 (N_7694,N_3305,N_4138);
nor U7695 (N_7695,N_3716,N_2883);
nand U7696 (N_7696,N_4187,N_4597);
and U7697 (N_7697,N_4461,N_465);
or U7698 (N_7698,N_2692,N_1643);
and U7699 (N_7699,N_3362,N_1822);
nor U7700 (N_7700,N_4348,N_4032);
nor U7701 (N_7701,N_4050,N_2);
xnor U7702 (N_7702,N_1859,N_2055);
nor U7703 (N_7703,N_4334,N_3388);
nor U7704 (N_7704,N_2916,N_377);
and U7705 (N_7705,N_1766,N_1908);
and U7706 (N_7706,N_1761,N_334);
xnor U7707 (N_7707,N_1271,N_1807);
nor U7708 (N_7708,N_989,N_1340);
and U7709 (N_7709,N_4697,N_2187);
and U7710 (N_7710,N_1751,N_45);
or U7711 (N_7711,N_2827,N_187);
xor U7712 (N_7712,N_2193,N_3610);
nand U7713 (N_7713,N_944,N_4227);
nor U7714 (N_7714,N_927,N_2403);
and U7715 (N_7715,N_1440,N_1596);
or U7716 (N_7716,N_1673,N_2087);
nand U7717 (N_7717,N_2815,N_2570);
nand U7718 (N_7718,N_213,N_4866);
or U7719 (N_7719,N_376,N_3270);
nor U7720 (N_7720,N_3049,N_1920);
or U7721 (N_7721,N_728,N_2103);
nand U7722 (N_7722,N_1962,N_2788);
and U7723 (N_7723,N_3626,N_198);
nor U7724 (N_7724,N_1989,N_4278);
or U7725 (N_7725,N_291,N_2458);
nor U7726 (N_7726,N_2955,N_2573);
or U7727 (N_7727,N_3034,N_3757);
or U7728 (N_7728,N_4184,N_1847);
nand U7729 (N_7729,N_881,N_4386);
or U7730 (N_7730,N_1592,N_1085);
nor U7731 (N_7731,N_2010,N_2165);
nand U7732 (N_7732,N_2187,N_3409);
or U7733 (N_7733,N_3538,N_4093);
and U7734 (N_7734,N_3062,N_4582);
and U7735 (N_7735,N_685,N_1949);
nand U7736 (N_7736,N_4095,N_1413);
nor U7737 (N_7737,N_4604,N_168);
nor U7738 (N_7738,N_822,N_4274);
or U7739 (N_7739,N_2703,N_106);
nor U7740 (N_7740,N_978,N_2286);
or U7741 (N_7741,N_2032,N_4354);
nand U7742 (N_7742,N_495,N_1221);
or U7743 (N_7743,N_4854,N_2047);
and U7744 (N_7744,N_2736,N_210);
nor U7745 (N_7745,N_3989,N_4237);
or U7746 (N_7746,N_2678,N_4438);
and U7747 (N_7747,N_1159,N_4071);
nand U7748 (N_7748,N_2325,N_255);
xor U7749 (N_7749,N_535,N_2251);
nor U7750 (N_7750,N_4685,N_4296);
and U7751 (N_7751,N_1119,N_379);
nand U7752 (N_7752,N_4668,N_1924);
nor U7753 (N_7753,N_3828,N_4766);
nor U7754 (N_7754,N_2821,N_3036);
nor U7755 (N_7755,N_4493,N_2382);
and U7756 (N_7756,N_3378,N_2559);
and U7757 (N_7757,N_3234,N_4328);
or U7758 (N_7758,N_3392,N_358);
and U7759 (N_7759,N_2477,N_2);
and U7760 (N_7760,N_3601,N_1515);
nor U7761 (N_7761,N_3421,N_3543);
nand U7762 (N_7762,N_2672,N_2318);
nand U7763 (N_7763,N_926,N_1711);
and U7764 (N_7764,N_99,N_778);
or U7765 (N_7765,N_1758,N_2910);
or U7766 (N_7766,N_2822,N_4469);
nor U7767 (N_7767,N_4638,N_3312);
nand U7768 (N_7768,N_3759,N_1949);
nand U7769 (N_7769,N_2410,N_3311);
nor U7770 (N_7770,N_4876,N_2198);
or U7771 (N_7771,N_1647,N_1557);
and U7772 (N_7772,N_3414,N_4402);
and U7773 (N_7773,N_2048,N_1748);
and U7774 (N_7774,N_2988,N_3366);
nor U7775 (N_7775,N_4060,N_4759);
nor U7776 (N_7776,N_1766,N_787);
nand U7777 (N_7777,N_3662,N_3584);
or U7778 (N_7778,N_4510,N_396);
nor U7779 (N_7779,N_4935,N_1061);
or U7780 (N_7780,N_4732,N_2780);
nor U7781 (N_7781,N_659,N_2801);
nand U7782 (N_7782,N_2833,N_4246);
nor U7783 (N_7783,N_1830,N_592);
or U7784 (N_7784,N_1234,N_4239);
and U7785 (N_7785,N_853,N_664);
nand U7786 (N_7786,N_2004,N_4974);
nor U7787 (N_7787,N_787,N_4725);
and U7788 (N_7788,N_4036,N_1907);
or U7789 (N_7789,N_1668,N_26);
and U7790 (N_7790,N_4564,N_1031);
xnor U7791 (N_7791,N_294,N_925);
nand U7792 (N_7792,N_3180,N_2614);
or U7793 (N_7793,N_4877,N_4475);
nand U7794 (N_7794,N_3399,N_3308);
or U7795 (N_7795,N_4814,N_2166);
or U7796 (N_7796,N_4821,N_919);
or U7797 (N_7797,N_2986,N_3651);
nor U7798 (N_7798,N_2987,N_3535);
nor U7799 (N_7799,N_1616,N_1879);
nand U7800 (N_7800,N_1327,N_2779);
nand U7801 (N_7801,N_1037,N_1266);
or U7802 (N_7802,N_4768,N_1630);
xnor U7803 (N_7803,N_4774,N_1033);
and U7804 (N_7804,N_4257,N_2050);
nor U7805 (N_7805,N_463,N_941);
or U7806 (N_7806,N_3064,N_1234);
or U7807 (N_7807,N_3475,N_1022);
and U7808 (N_7808,N_2535,N_4014);
nand U7809 (N_7809,N_1385,N_1985);
nand U7810 (N_7810,N_1926,N_534);
and U7811 (N_7811,N_3479,N_1219);
nor U7812 (N_7812,N_1521,N_359);
nand U7813 (N_7813,N_710,N_161);
nand U7814 (N_7814,N_1347,N_1633);
nor U7815 (N_7815,N_4713,N_4442);
or U7816 (N_7816,N_4144,N_3321);
or U7817 (N_7817,N_1577,N_4432);
and U7818 (N_7818,N_4549,N_2068);
or U7819 (N_7819,N_3893,N_3271);
or U7820 (N_7820,N_2514,N_4880);
or U7821 (N_7821,N_311,N_832);
nor U7822 (N_7822,N_1167,N_3634);
or U7823 (N_7823,N_2527,N_3852);
and U7824 (N_7824,N_4348,N_4803);
nand U7825 (N_7825,N_1681,N_1492);
nand U7826 (N_7826,N_1073,N_2137);
nand U7827 (N_7827,N_4311,N_667);
nor U7828 (N_7828,N_3799,N_3754);
and U7829 (N_7829,N_2159,N_4165);
nor U7830 (N_7830,N_4265,N_2033);
or U7831 (N_7831,N_1363,N_1561);
or U7832 (N_7832,N_2781,N_3639);
nand U7833 (N_7833,N_1398,N_4846);
and U7834 (N_7834,N_3891,N_668);
or U7835 (N_7835,N_1091,N_4117);
and U7836 (N_7836,N_2369,N_3127);
and U7837 (N_7837,N_4184,N_3984);
nand U7838 (N_7838,N_3128,N_3808);
and U7839 (N_7839,N_325,N_3319);
and U7840 (N_7840,N_1972,N_201);
and U7841 (N_7841,N_1966,N_1801);
nor U7842 (N_7842,N_293,N_2678);
nor U7843 (N_7843,N_684,N_2263);
or U7844 (N_7844,N_2127,N_4058);
or U7845 (N_7845,N_431,N_4180);
or U7846 (N_7846,N_173,N_4002);
xnor U7847 (N_7847,N_1040,N_2123);
or U7848 (N_7848,N_2263,N_821);
and U7849 (N_7849,N_2413,N_4883);
and U7850 (N_7850,N_422,N_3208);
nand U7851 (N_7851,N_4142,N_636);
nor U7852 (N_7852,N_2570,N_2338);
and U7853 (N_7853,N_2043,N_4842);
nor U7854 (N_7854,N_2814,N_2336);
nor U7855 (N_7855,N_4991,N_3958);
nand U7856 (N_7856,N_2024,N_2253);
and U7857 (N_7857,N_974,N_2501);
or U7858 (N_7858,N_1141,N_3311);
or U7859 (N_7859,N_3307,N_740);
nor U7860 (N_7860,N_4104,N_2494);
and U7861 (N_7861,N_4906,N_4355);
and U7862 (N_7862,N_3898,N_3631);
and U7863 (N_7863,N_3981,N_2028);
and U7864 (N_7864,N_4285,N_3753);
and U7865 (N_7865,N_1801,N_4775);
and U7866 (N_7866,N_4837,N_446);
and U7867 (N_7867,N_395,N_2828);
nand U7868 (N_7868,N_3011,N_4610);
or U7869 (N_7869,N_4056,N_2181);
nand U7870 (N_7870,N_2218,N_1974);
and U7871 (N_7871,N_2477,N_4540);
or U7872 (N_7872,N_1882,N_3892);
and U7873 (N_7873,N_4824,N_3431);
nand U7874 (N_7874,N_2084,N_3532);
nand U7875 (N_7875,N_3298,N_2583);
or U7876 (N_7876,N_3124,N_1378);
xnor U7877 (N_7877,N_1687,N_3732);
nor U7878 (N_7878,N_3894,N_2783);
nor U7879 (N_7879,N_1346,N_3706);
or U7880 (N_7880,N_296,N_3417);
and U7881 (N_7881,N_3163,N_1165);
nand U7882 (N_7882,N_218,N_1141);
and U7883 (N_7883,N_2551,N_4492);
nor U7884 (N_7884,N_1184,N_3192);
nor U7885 (N_7885,N_2444,N_1806);
nand U7886 (N_7886,N_2158,N_529);
and U7887 (N_7887,N_4096,N_2715);
nand U7888 (N_7888,N_4354,N_3809);
nand U7889 (N_7889,N_3409,N_903);
nand U7890 (N_7890,N_4225,N_3079);
nand U7891 (N_7891,N_1223,N_1620);
nand U7892 (N_7892,N_1619,N_2038);
nand U7893 (N_7893,N_4229,N_1299);
or U7894 (N_7894,N_1599,N_1338);
nor U7895 (N_7895,N_2262,N_454);
nor U7896 (N_7896,N_2869,N_2254);
nor U7897 (N_7897,N_2059,N_694);
nor U7898 (N_7898,N_4381,N_2405);
or U7899 (N_7899,N_584,N_521);
or U7900 (N_7900,N_853,N_195);
and U7901 (N_7901,N_2920,N_1960);
or U7902 (N_7902,N_4430,N_245);
nor U7903 (N_7903,N_2825,N_3585);
nand U7904 (N_7904,N_282,N_4873);
nor U7905 (N_7905,N_3702,N_915);
and U7906 (N_7906,N_1575,N_1809);
and U7907 (N_7907,N_2947,N_1397);
and U7908 (N_7908,N_3190,N_4763);
or U7909 (N_7909,N_4774,N_2613);
or U7910 (N_7910,N_4145,N_1525);
or U7911 (N_7911,N_1500,N_3089);
and U7912 (N_7912,N_2336,N_1180);
or U7913 (N_7913,N_1590,N_2578);
nor U7914 (N_7914,N_2440,N_1290);
nor U7915 (N_7915,N_3971,N_1468);
and U7916 (N_7916,N_437,N_52);
nand U7917 (N_7917,N_396,N_545);
nor U7918 (N_7918,N_1078,N_1100);
or U7919 (N_7919,N_592,N_2740);
nor U7920 (N_7920,N_643,N_2332);
nand U7921 (N_7921,N_1462,N_2764);
nand U7922 (N_7922,N_2481,N_4284);
or U7923 (N_7923,N_347,N_4157);
or U7924 (N_7924,N_2303,N_4207);
nand U7925 (N_7925,N_606,N_4998);
or U7926 (N_7926,N_1493,N_4601);
nand U7927 (N_7927,N_1605,N_1735);
and U7928 (N_7928,N_1552,N_3435);
nor U7929 (N_7929,N_4370,N_2274);
nand U7930 (N_7930,N_4874,N_3370);
or U7931 (N_7931,N_1828,N_1973);
nor U7932 (N_7932,N_1136,N_2920);
nand U7933 (N_7933,N_4345,N_1714);
or U7934 (N_7934,N_2905,N_285);
and U7935 (N_7935,N_4375,N_4514);
nor U7936 (N_7936,N_4080,N_915);
or U7937 (N_7937,N_3314,N_4605);
nor U7938 (N_7938,N_2860,N_2298);
and U7939 (N_7939,N_2703,N_436);
nand U7940 (N_7940,N_3501,N_3201);
or U7941 (N_7941,N_1389,N_3127);
and U7942 (N_7942,N_3352,N_3937);
nand U7943 (N_7943,N_724,N_4041);
or U7944 (N_7944,N_3500,N_992);
nand U7945 (N_7945,N_2407,N_3420);
nor U7946 (N_7946,N_113,N_4401);
and U7947 (N_7947,N_316,N_3682);
nand U7948 (N_7948,N_1384,N_882);
and U7949 (N_7949,N_3132,N_1085);
nand U7950 (N_7950,N_4364,N_3222);
nand U7951 (N_7951,N_1686,N_4087);
and U7952 (N_7952,N_1179,N_439);
nand U7953 (N_7953,N_4753,N_3536);
xnor U7954 (N_7954,N_1141,N_1573);
nand U7955 (N_7955,N_1798,N_2292);
nand U7956 (N_7956,N_2064,N_4615);
nor U7957 (N_7957,N_141,N_3681);
xor U7958 (N_7958,N_4338,N_2681);
and U7959 (N_7959,N_4281,N_2560);
or U7960 (N_7960,N_3339,N_2285);
nand U7961 (N_7961,N_1121,N_3280);
and U7962 (N_7962,N_1397,N_2817);
and U7963 (N_7963,N_1051,N_4677);
or U7964 (N_7964,N_2418,N_4891);
nor U7965 (N_7965,N_3901,N_3731);
or U7966 (N_7966,N_3707,N_3330);
or U7967 (N_7967,N_2627,N_165);
nor U7968 (N_7968,N_3579,N_4276);
or U7969 (N_7969,N_2001,N_2903);
or U7970 (N_7970,N_2485,N_2336);
nand U7971 (N_7971,N_857,N_911);
and U7972 (N_7972,N_2404,N_1898);
and U7973 (N_7973,N_1985,N_3367);
xor U7974 (N_7974,N_3514,N_478);
nand U7975 (N_7975,N_1401,N_2166);
nand U7976 (N_7976,N_653,N_1434);
nor U7977 (N_7977,N_2353,N_3998);
nor U7978 (N_7978,N_3133,N_2162);
nand U7979 (N_7979,N_3392,N_3686);
or U7980 (N_7980,N_1122,N_2307);
or U7981 (N_7981,N_3238,N_3344);
xor U7982 (N_7982,N_2160,N_551);
and U7983 (N_7983,N_1433,N_3816);
nor U7984 (N_7984,N_4584,N_3421);
nand U7985 (N_7985,N_2985,N_2842);
and U7986 (N_7986,N_487,N_4665);
nor U7987 (N_7987,N_4711,N_3553);
nor U7988 (N_7988,N_4032,N_1035);
nand U7989 (N_7989,N_2082,N_3490);
nor U7990 (N_7990,N_682,N_1643);
nor U7991 (N_7991,N_1472,N_2519);
or U7992 (N_7992,N_356,N_2201);
or U7993 (N_7993,N_564,N_4478);
nor U7994 (N_7994,N_2877,N_4584);
xnor U7995 (N_7995,N_3278,N_2308);
nand U7996 (N_7996,N_4364,N_743);
or U7997 (N_7997,N_1170,N_246);
and U7998 (N_7998,N_3697,N_4752);
nor U7999 (N_7999,N_3885,N_3300);
nor U8000 (N_8000,N_695,N_339);
nand U8001 (N_8001,N_1140,N_2914);
and U8002 (N_8002,N_2436,N_3517);
and U8003 (N_8003,N_676,N_4582);
nor U8004 (N_8004,N_1145,N_3178);
nand U8005 (N_8005,N_4158,N_3524);
nor U8006 (N_8006,N_4380,N_3533);
nand U8007 (N_8007,N_485,N_3939);
and U8008 (N_8008,N_2160,N_202);
nand U8009 (N_8009,N_4808,N_4751);
nand U8010 (N_8010,N_4600,N_4251);
xnor U8011 (N_8011,N_2147,N_2058);
or U8012 (N_8012,N_1012,N_1196);
nand U8013 (N_8013,N_1905,N_2952);
and U8014 (N_8014,N_0,N_3774);
and U8015 (N_8015,N_1871,N_911);
xor U8016 (N_8016,N_4981,N_4322);
nor U8017 (N_8017,N_3848,N_1535);
nor U8018 (N_8018,N_4854,N_4991);
nand U8019 (N_8019,N_3105,N_443);
nand U8020 (N_8020,N_764,N_3418);
nand U8021 (N_8021,N_1084,N_1288);
nor U8022 (N_8022,N_4106,N_2079);
nand U8023 (N_8023,N_3425,N_4807);
and U8024 (N_8024,N_210,N_3412);
nor U8025 (N_8025,N_1466,N_4554);
or U8026 (N_8026,N_4109,N_1036);
nor U8027 (N_8027,N_4155,N_12);
or U8028 (N_8028,N_2855,N_3276);
and U8029 (N_8029,N_2596,N_3549);
nand U8030 (N_8030,N_4496,N_3132);
nor U8031 (N_8031,N_1449,N_2051);
and U8032 (N_8032,N_2122,N_3558);
nor U8033 (N_8033,N_1898,N_300);
or U8034 (N_8034,N_4942,N_4324);
and U8035 (N_8035,N_3606,N_3239);
or U8036 (N_8036,N_4120,N_275);
or U8037 (N_8037,N_3070,N_3437);
and U8038 (N_8038,N_1929,N_4079);
nand U8039 (N_8039,N_3114,N_892);
nor U8040 (N_8040,N_1702,N_1417);
nor U8041 (N_8041,N_4859,N_1355);
or U8042 (N_8042,N_4416,N_1338);
or U8043 (N_8043,N_1196,N_2381);
nor U8044 (N_8044,N_4297,N_2102);
and U8045 (N_8045,N_35,N_1208);
nand U8046 (N_8046,N_4715,N_4030);
nand U8047 (N_8047,N_2244,N_4182);
or U8048 (N_8048,N_3380,N_2191);
and U8049 (N_8049,N_2622,N_2483);
or U8050 (N_8050,N_3526,N_3698);
nor U8051 (N_8051,N_3792,N_2712);
nor U8052 (N_8052,N_1434,N_4630);
or U8053 (N_8053,N_326,N_698);
nor U8054 (N_8054,N_3788,N_1312);
and U8055 (N_8055,N_2440,N_4457);
or U8056 (N_8056,N_3732,N_1069);
nor U8057 (N_8057,N_3332,N_3453);
or U8058 (N_8058,N_1240,N_2389);
xor U8059 (N_8059,N_4814,N_1282);
nand U8060 (N_8060,N_1281,N_780);
nand U8061 (N_8061,N_837,N_3075);
and U8062 (N_8062,N_3194,N_2585);
nand U8063 (N_8063,N_883,N_2994);
and U8064 (N_8064,N_2734,N_1443);
or U8065 (N_8065,N_368,N_3964);
and U8066 (N_8066,N_1748,N_4670);
or U8067 (N_8067,N_3099,N_3831);
and U8068 (N_8068,N_1218,N_1053);
nor U8069 (N_8069,N_2879,N_1916);
or U8070 (N_8070,N_1984,N_2593);
or U8071 (N_8071,N_4657,N_937);
xnor U8072 (N_8072,N_4238,N_1411);
or U8073 (N_8073,N_3264,N_1574);
or U8074 (N_8074,N_527,N_4870);
nor U8075 (N_8075,N_4980,N_1056);
nand U8076 (N_8076,N_1741,N_3583);
nor U8077 (N_8077,N_889,N_4271);
and U8078 (N_8078,N_16,N_4066);
or U8079 (N_8079,N_1127,N_769);
and U8080 (N_8080,N_211,N_1906);
nor U8081 (N_8081,N_4696,N_4125);
and U8082 (N_8082,N_3306,N_3525);
and U8083 (N_8083,N_2535,N_3882);
nor U8084 (N_8084,N_314,N_2854);
nor U8085 (N_8085,N_4331,N_2699);
nand U8086 (N_8086,N_3528,N_3913);
nand U8087 (N_8087,N_3150,N_3821);
nor U8088 (N_8088,N_2199,N_4711);
and U8089 (N_8089,N_4870,N_4259);
nand U8090 (N_8090,N_1535,N_749);
and U8091 (N_8091,N_1707,N_4782);
and U8092 (N_8092,N_1452,N_4876);
nand U8093 (N_8093,N_4401,N_504);
and U8094 (N_8094,N_2697,N_1771);
or U8095 (N_8095,N_2413,N_3527);
nand U8096 (N_8096,N_3518,N_3053);
and U8097 (N_8097,N_367,N_823);
and U8098 (N_8098,N_1038,N_4159);
and U8099 (N_8099,N_2790,N_2813);
or U8100 (N_8100,N_2804,N_4297);
and U8101 (N_8101,N_1601,N_4560);
nand U8102 (N_8102,N_334,N_1777);
nand U8103 (N_8103,N_3187,N_481);
nor U8104 (N_8104,N_1695,N_873);
or U8105 (N_8105,N_1811,N_1713);
nor U8106 (N_8106,N_2074,N_3122);
nand U8107 (N_8107,N_70,N_3743);
nor U8108 (N_8108,N_3244,N_4570);
nor U8109 (N_8109,N_3619,N_4810);
nand U8110 (N_8110,N_4343,N_147);
or U8111 (N_8111,N_4008,N_2152);
and U8112 (N_8112,N_600,N_4096);
or U8113 (N_8113,N_4682,N_2317);
nand U8114 (N_8114,N_1446,N_2175);
nor U8115 (N_8115,N_1549,N_548);
xor U8116 (N_8116,N_878,N_1013);
nor U8117 (N_8117,N_3481,N_3618);
and U8118 (N_8118,N_3611,N_1356);
nand U8119 (N_8119,N_2130,N_64);
nand U8120 (N_8120,N_795,N_2092);
nand U8121 (N_8121,N_2493,N_2428);
and U8122 (N_8122,N_3317,N_2612);
and U8123 (N_8123,N_4537,N_1790);
nor U8124 (N_8124,N_3332,N_2895);
nor U8125 (N_8125,N_3441,N_2020);
or U8126 (N_8126,N_1478,N_4151);
or U8127 (N_8127,N_330,N_4187);
and U8128 (N_8128,N_3779,N_3758);
nor U8129 (N_8129,N_563,N_792);
nand U8130 (N_8130,N_1462,N_2413);
or U8131 (N_8131,N_3771,N_4651);
and U8132 (N_8132,N_269,N_4531);
and U8133 (N_8133,N_3819,N_3146);
or U8134 (N_8134,N_1311,N_2787);
nor U8135 (N_8135,N_3083,N_464);
or U8136 (N_8136,N_360,N_3205);
or U8137 (N_8137,N_1389,N_769);
xor U8138 (N_8138,N_4328,N_1275);
or U8139 (N_8139,N_4809,N_3031);
nor U8140 (N_8140,N_1649,N_4939);
nor U8141 (N_8141,N_3671,N_1547);
or U8142 (N_8142,N_4074,N_1255);
and U8143 (N_8143,N_831,N_2464);
xor U8144 (N_8144,N_1126,N_4529);
nor U8145 (N_8145,N_319,N_308);
or U8146 (N_8146,N_1062,N_4007);
nor U8147 (N_8147,N_2122,N_3352);
or U8148 (N_8148,N_3877,N_4853);
and U8149 (N_8149,N_3684,N_1539);
and U8150 (N_8150,N_3683,N_4003);
and U8151 (N_8151,N_3055,N_2173);
xor U8152 (N_8152,N_1181,N_4428);
or U8153 (N_8153,N_2423,N_4524);
nand U8154 (N_8154,N_3450,N_3376);
and U8155 (N_8155,N_4856,N_726);
or U8156 (N_8156,N_1127,N_887);
nand U8157 (N_8157,N_4002,N_2046);
nand U8158 (N_8158,N_1925,N_355);
nor U8159 (N_8159,N_3575,N_2515);
nand U8160 (N_8160,N_3025,N_462);
and U8161 (N_8161,N_3282,N_1333);
or U8162 (N_8162,N_1469,N_2645);
and U8163 (N_8163,N_115,N_3880);
nor U8164 (N_8164,N_2858,N_2344);
or U8165 (N_8165,N_2464,N_4850);
nor U8166 (N_8166,N_1020,N_4480);
or U8167 (N_8167,N_3821,N_1677);
nand U8168 (N_8168,N_4000,N_4546);
or U8169 (N_8169,N_1962,N_4487);
and U8170 (N_8170,N_2794,N_2787);
nand U8171 (N_8171,N_615,N_3105);
nor U8172 (N_8172,N_4292,N_162);
and U8173 (N_8173,N_4424,N_4354);
and U8174 (N_8174,N_2246,N_1905);
or U8175 (N_8175,N_1315,N_900);
and U8176 (N_8176,N_4711,N_3512);
nor U8177 (N_8177,N_2615,N_4916);
or U8178 (N_8178,N_1931,N_3839);
nand U8179 (N_8179,N_2246,N_1856);
nand U8180 (N_8180,N_575,N_2954);
or U8181 (N_8181,N_195,N_1994);
or U8182 (N_8182,N_3,N_2468);
nand U8183 (N_8183,N_3060,N_3052);
and U8184 (N_8184,N_4679,N_1036);
nand U8185 (N_8185,N_1104,N_1390);
nor U8186 (N_8186,N_3882,N_3231);
nand U8187 (N_8187,N_1559,N_18);
or U8188 (N_8188,N_465,N_4093);
nor U8189 (N_8189,N_1476,N_501);
nand U8190 (N_8190,N_3311,N_4404);
nand U8191 (N_8191,N_2495,N_2907);
and U8192 (N_8192,N_4346,N_4373);
nor U8193 (N_8193,N_4920,N_472);
or U8194 (N_8194,N_3411,N_1964);
or U8195 (N_8195,N_3538,N_1614);
nand U8196 (N_8196,N_4094,N_3249);
and U8197 (N_8197,N_1569,N_3582);
nor U8198 (N_8198,N_4471,N_3466);
or U8199 (N_8199,N_1668,N_1298);
and U8200 (N_8200,N_3879,N_3970);
nor U8201 (N_8201,N_1070,N_1187);
and U8202 (N_8202,N_697,N_1289);
nor U8203 (N_8203,N_3564,N_471);
nand U8204 (N_8204,N_3280,N_4245);
nand U8205 (N_8205,N_1003,N_3285);
nand U8206 (N_8206,N_1494,N_2424);
nand U8207 (N_8207,N_640,N_1174);
and U8208 (N_8208,N_3507,N_153);
and U8209 (N_8209,N_1893,N_1571);
nand U8210 (N_8210,N_1283,N_4823);
and U8211 (N_8211,N_700,N_2998);
or U8212 (N_8212,N_1879,N_3241);
nor U8213 (N_8213,N_183,N_3340);
nor U8214 (N_8214,N_3427,N_921);
nor U8215 (N_8215,N_3415,N_4226);
nand U8216 (N_8216,N_2163,N_2468);
nor U8217 (N_8217,N_2728,N_1001);
or U8218 (N_8218,N_31,N_2977);
and U8219 (N_8219,N_4530,N_4132);
and U8220 (N_8220,N_4149,N_2777);
and U8221 (N_8221,N_3224,N_4199);
nor U8222 (N_8222,N_2124,N_1409);
nand U8223 (N_8223,N_1107,N_2592);
nand U8224 (N_8224,N_1733,N_3169);
or U8225 (N_8225,N_1156,N_3679);
and U8226 (N_8226,N_3513,N_975);
or U8227 (N_8227,N_53,N_3611);
nand U8228 (N_8228,N_1187,N_4948);
and U8229 (N_8229,N_4427,N_2884);
or U8230 (N_8230,N_4203,N_2011);
nand U8231 (N_8231,N_4563,N_2694);
or U8232 (N_8232,N_807,N_3195);
xor U8233 (N_8233,N_4560,N_4432);
nor U8234 (N_8234,N_660,N_3212);
and U8235 (N_8235,N_3494,N_3999);
nand U8236 (N_8236,N_2635,N_1014);
or U8237 (N_8237,N_2557,N_2658);
nand U8238 (N_8238,N_4111,N_2764);
nand U8239 (N_8239,N_729,N_4404);
and U8240 (N_8240,N_4240,N_4059);
nand U8241 (N_8241,N_1719,N_2098);
and U8242 (N_8242,N_1074,N_1917);
and U8243 (N_8243,N_4592,N_3421);
and U8244 (N_8244,N_3770,N_4372);
nand U8245 (N_8245,N_623,N_3507);
and U8246 (N_8246,N_2589,N_3165);
and U8247 (N_8247,N_221,N_3915);
nor U8248 (N_8248,N_2154,N_2623);
nand U8249 (N_8249,N_4096,N_4937);
and U8250 (N_8250,N_4984,N_3094);
and U8251 (N_8251,N_487,N_3462);
nand U8252 (N_8252,N_2153,N_4199);
or U8253 (N_8253,N_2446,N_934);
nor U8254 (N_8254,N_46,N_2340);
nor U8255 (N_8255,N_937,N_3608);
or U8256 (N_8256,N_1066,N_121);
and U8257 (N_8257,N_154,N_2542);
nor U8258 (N_8258,N_1487,N_1447);
nand U8259 (N_8259,N_735,N_2462);
or U8260 (N_8260,N_3077,N_2458);
nand U8261 (N_8261,N_3045,N_4650);
and U8262 (N_8262,N_4800,N_611);
and U8263 (N_8263,N_2760,N_840);
or U8264 (N_8264,N_819,N_3302);
nor U8265 (N_8265,N_1346,N_3461);
or U8266 (N_8266,N_894,N_145);
or U8267 (N_8267,N_2977,N_4709);
nor U8268 (N_8268,N_3430,N_1218);
or U8269 (N_8269,N_664,N_4504);
or U8270 (N_8270,N_997,N_19);
nand U8271 (N_8271,N_4897,N_3419);
or U8272 (N_8272,N_285,N_2237);
nand U8273 (N_8273,N_1940,N_404);
or U8274 (N_8274,N_330,N_4097);
and U8275 (N_8275,N_1608,N_1150);
or U8276 (N_8276,N_2756,N_1451);
nor U8277 (N_8277,N_4314,N_2484);
and U8278 (N_8278,N_4897,N_227);
and U8279 (N_8279,N_1573,N_12);
nand U8280 (N_8280,N_164,N_3176);
and U8281 (N_8281,N_1341,N_1588);
xor U8282 (N_8282,N_10,N_4024);
or U8283 (N_8283,N_3012,N_4816);
nor U8284 (N_8284,N_1465,N_2066);
and U8285 (N_8285,N_4642,N_1208);
or U8286 (N_8286,N_2705,N_2802);
and U8287 (N_8287,N_4506,N_2313);
nand U8288 (N_8288,N_1926,N_1326);
nor U8289 (N_8289,N_2326,N_4477);
and U8290 (N_8290,N_2234,N_2513);
nor U8291 (N_8291,N_1421,N_1781);
nand U8292 (N_8292,N_34,N_1060);
xor U8293 (N_8293,N_3009,N_3766);
nand U8294 (N_8294,N_3889,N_2006);
and U8295 (N_8295,N_577,N_4406);
nand U8296 (N_8296,N_1973,N_2940);
nand U8297 (N_8297,N_1337,N_4665);
nor U8298 (N_8298,N_892,N_2505);
and U8299 (N_8299,N_4699,N_1552);
nor U8300 (N_8300,N_2045,N_4396);
and U8301 (N_8301,N_184,N_4662);
or U8302 (N_8302,N_4555,N_4933);
and U8303 (N_8303,N_3824,N_2943);
and U8304 (N_8304,N_599,N_1236);
and U8305 (N_8305,N_4945,N_4522);
nand U8306 (N_8306,N_2261,N_2588);
or U8307 (N_8307,N_1317,N_294);
and U8308 (N_8308,N_4897,N_1157);
and U8309 (N_8309,N_2232,N_99);
and U8310 (N_8310,N_3767,N_1599);
nand U8311 (N_8311,N_3421,N_794);
and U8312 (N_8312,N_4007,N_3061);
nand U8313 (N_8313,N_4882,N_3096);
nand U8314 (N_8314,N_3232,N_4715);
nor U8315 (N_8315,N_2820,N_2345);
or U8316 (N_8316,N_2271,N_2775);
xnor U8317 (N_8317,N_3403,N_1139);
and U8318 (N_8318,N_4897,N_1622);
xor U8319 (N_8319,N_3083,N_4150);
and U8320 (N_8320,N_4295,N_145);
and U8321 (N_8321,N_2306,N_3464);
or U8322 (N_8322,N_1194,N_1698);
and U8323 (N_8323,N_3511,N_2816);
nand U8324 (N_8324,N_1282,N_4034);
or U8325 (N_8325,N_2204,N_2994);
and U8326 (N_8326,N_4137,N_3808);
nor U8327 (N_8327,N_943,N_4330);
nor U8328 (N_8328,N_2981,N_400);
nand U8329 (N_8329,N_1923,N_4538);
nand U8330 (N_8330,N_3481,N_460);
nand U8331 (N_8331,N_2886,N_2090);
or U8332 (N_8332,N_4859,N_1434);
or U8333 (N_8333,N_2508,N_1762);
or U8334 (N_8334,N_486,N_4126);
nor U8335 (N_8335,N_3610,N_3318);
and U8336 (N_8336,N_3660,N_107);
or U8337 (N_8337,N_1668,N_4113);
and U8338 (N_8338,N_4912,N_886);
or U8339 (N_8339,N_2259,N_3974);
and U8340 (N_8340,N_4403,N_117);
or U8341 (N_8341,N_3482,N_687);
or U8342 (N_8342,N_1793,N_4244);
nor U8343 (N_8343,N_2915,N_1025);
or U8344 (N_8344,N_4835,N_307);
or U8345 (N_8345,N_4441,N_4957);
nand U8346 (N_8346,N_2467,N_4875);
nor U8347 (N_8347,N_919,N_15);
xnor U8348 (N_8348,N_41,N_2937);
nand U8349 (N_8349,N_4930,N_4411);
nand U8350 (N_8350,N_2887,N_4837);
nor U8351 (N_8351,N_4127,N_2844);
or U8352 (N_8352,N_3005,N_1171);
nand U8353 (N_8353,N_319,N_4139);
nor U8354 (N_8354,N_4921,N_3506);
nand U8355 (N_8355,N_4439,N_859);
or U8356 (N_8356,N_1499,N_3162);
nor U8357 (N_8357,N_3192,N_2267);
or U8358 (N_8358,N_2159,N_1403);
nand U8359 (N_8359,N_2734,N_2729);
nand U8360 (N_8360,N_695,N_3669);
and U8361 (N_8361,N_3616,N_2632);
xnor U8362 (N_8362,N_3134,N_3604);
nor U8363 (N_8363,N_3559,N_4858);
and U8364 (N_8364,N_2208,N_4020);
nand U8365 (N_8365,N_3115,N_166);
or U8366 (N_8366,N_124,N_3058);
nor U8367 (N_8367,N_399,N_2285);
and U8368 (N_8368,N_2674,N_3793);
and U8369 (N_8369,N_1507,N_401);
nand U8370 (N_8370,N_1941,N_1083);
nand U8371 (N_8371,N_610,N_1672);
nand U8372 (N_8372,N_4528,N_4074);
nor U8373 (N_8373,N_890,N_175);
xor U8374 (N_8374,N_2782,N_2526);
or U8375 (N_8375,N_2086,N_2846);
nand U8376 (N_8376,N_735,N_2547);
nand U8377 (N_8377,N_3897,N_4350);
nand U8378 (N_8378,N_801,N_4243);
and U8379 (N_8379,N_4198,N_2029);
or U8380 (N_8380,N_2725,N_4317);
and U8381 (N_8381,N_3755,N_855);
or U8382 (N_8382,N_2914,N_3352);
nand U8383 (N_8383,N_2853,N_1005);
or U8384 (N_8384,N_2094,N_2418);
and U8385 (N_8385,N_329,N_580);
nand U8386 (N_8386,N_3059,N_3964);
nor U8387 (N_8387,N_4442,N_3371);
or U8388 (N_8388,N_1584,N_1175);
and U8389 (N_8389,N_2309,N_2730);
nor U8390 (N_8390,N_44,N_2408);
or U8391 (N_8391,N_4939,N_2128);
or U8392 (N_8392,N_4082,N_3129);
nand U8393 (N_8393,N_66,N_2742);
nor U8394 (N_8394,N_2399,N_1946);
nor U8395 (N_8395,N_1877,N_4177);
and U8396 (N_8396,N_3385,N_686);
and U8397 (N_8397,N_121,N_2642);
nand U8398 (N_8398,N_1098,N_3625);
nor U8399 (N_8399,N_2367,N_304);
and U8400 (N_8400,N_4942,N_3477);
or U8401 (N_8401,N_2563,N_4694);
nor U8402 (N_8402,N_285,N_1798);
nor U8403 (N_8403,N_3001,N_239);
or U8404 (N_8404,N_1205,N_2627);
nand U8405 (N_8405,N_3875,N_4722);
or U8406 (N_8406,N_3753,N_1597);
or U8407 (N_8407,N_165,N_3008);
nand U8408 (N_8408,N_4278,N_2086);
nand U8409 (N_8409,N_4669,N_3621);
xor U8410 (N_8410,N_3735,N_181);
or U8411 (N_8411,N_4817,N_4918);
and U8412 (N_8412,N_2345,N_4881);
or U8413 (N_8413,N_2981,N_4643);
nor U8414 (N_8414,N_1252,N_4237);
nand U8415 (N_8415,N_907,N_3773);
or U8416 (N_8416,N_3546,N_3122);
nor U8417 (N_8417,N_4423,N_1586);
and U8418 (N_8418,N_2904,N_2157);
nand U8419 (N_8419,N_1548,N_2684);
nand U8420 (N_8420,N_4767,N_3506);
and U8421 (N_8421,N_4241,N_1652);
nand U8422 (N_8422,N_170,N_2866);
or U8423 (N_8423,N_1937,N_4897);
and U8424 (N_8424,N_4416,N_1075);
or U8425 (N_8425,N_3225,N_3245);
or U8426 (N_8426,N_1641,N_1943);
nand U8427 (N_8427,N_2626,N_3800);
and U8428 (N_8428,N_2511,N_1507);
or U8429 (N_8429,N_2555,N_1762);
nand U8430 (N_8430,N_4190,N_3937);
and U8431 (N_8431,N_2350,N_131);
nor U8432 (N_8432,N_1273,N_516);
or U8433 (N_8433,N_1598,N_3651);
nand U8434 (N_8434,N_2915,N_3734);
nor U8435 (N_8435,N_4679,N_1513);
nand U8436 (N_8436,N_2874,N_889);
or U8437 (N_8437,N_1184,N_774);
nand U8438 (N_8438,N_3942,N_3266);
nand U8439 (N_8439,N_2742,N_443);
or U8440 (N_8440,N_778,N_4131);
nor U8441 (N_8441,N_2138,N_1468);
nand U8442 (N_8442,N_1208,N_4801);
or U8443 (N_8443,N_3497,N_4389);
or U8444 (N_8444,N_1339,N_3443);
nand U8445 (N_8445,N_764,N_3769);
or U8446 (N_8446,N_2762,N_1051);
nand U8447 (N_8447,N_256,N_1000);
nand U8448 (N_8448,N_773,N_2435);
or U8449 (N_8449,N_679,N_2740);
nand U8450 (N_8450,N_327,N_1707);
nand U8451 (N_8451,N_2342,N_1642);
and U8452 (N_8452,N_544,N_541);
nand U8453 (N_8453,N_2068,N_2122);
nor U8454 (N_8454,N_2322,N_3406);
nand U8455 (N_8455,N_4419,N_2265);
and U8456 (N_8456,N_1199,N_2188);
nor U8457 (N_8457,N_1396,N_224);
or U8458 (N_8458,N_2665,N_520);
and U8459 (N_8459,N_1506,N_718);
nand U8460 (N_8460,N_2327,N_1674);
nand U8461 (N_8461,N_1270,N_2062);
and U8462 (N_8462,N_3576,N_2487);
nand U8463 (N_8463,N_2522,N_35);
or U8464 (N_8464,N_3928,N_1907);
nand U8465 (N_8465,N_3603,N_703);
or U8466 (N_8466,N_3510,N_1549);
nand U8467 (N_8467,N_2706,N_3938);
nor U8468 (N_8468,N_3748,N_321);
nor U8469 (N_8469,N_3011,N_758);
and U8470 (N_8470,N_3057,N_3526);
and U8471 (N_8471,N_2853,N_1101);
nand U8472 (N_8472,N_27,N_714);
or U8473 (N_8473,N_3705,N_974);
and U8474 (N_8474,N_3099,N_2293);
nand U8475 (N_8475,N_3135,N_2502);
xor U8476 (N_8476,N_2062,N_2367);
nor U8477 (N_8477,N_1252,N_2725);
and U8478 (N_8478,N_3042,N_3638);
nand U8479 (N_8479,N_2321,N_3383);
nand U8480 (N_8480,N_2168,N_1442);
nand U8481 (N_8481,N_1424,N_4097);
nor U8482 (N_8482,N_820,N_2968);
nand U8483 (N_8483,N_101,N_609);
and U8484 (N_8484,N_1583,N_4371);
nand U8485 (N_8485,N_1728,N_960);
or U8486 (N_8486,N_2215,N_4599);
nand U8487 (N_8487,N_3482,N_3275);
and U8488 (N_8488,N_4766,N_4959);
nor U8489 (N_8489,N_2826,N_1698);
nand U8490 (N_8490,N_3922,N_3252);
and U8491 (N_8491,N_4097,N_4593);
xnor U8492 (N_8492,N_2024,N_909);
or U8493 (N_8493,N_4101,N_116);
and U8494 (N_8494,N_4109,N_1394);
nor U8495 (N_8495,N_625,N_49);
and U8496 (N_8496,N_140,N_3823);
nor U8497 (N_8497,N_2530,N_624);
or U8498 (N_8498,N_3090,N_1575);
nand U8499 (N_8499,N_3821,N_2072);
nor U8500 (N_8500,N_4630,N_4967);
nor U8501 (N_8501,N_3551,N_4347);
nor U8502 (N_8502,N_4256,N_4741);
or U8503 (N_8503,N_1785,N_3174);
or U8504 (N_8504,N_2118,N_2086);
nand U8505 (N_8505,N_687,N_1221);
nand U8506 (N_8506,N_4778,N_975);
nand U8507 (N_8507,N_574,N_3080);
nor U8508 (N_8508,N_2271,N_2083);
and U8509 (N_8509,N_840,N_2786);
nor U8510 (N_8510,N_404,N_4166);
or U8511 (N_8511,N_4429,N_2065);
and U8512 (N_8512,N_67,N_3641);
nand U8513 (N_8513,N_2868,N_386);
xor U8514 (N_8514,N_1687,N_652);
or U8515 (N_8515,N_2562,N_3102);
or U8516 (N_8516,N_1392,N_839);
nor U8517 (N_8517,N_3936,N_912);
nand U8518 (N_8518,N_2286,N_3594);
xor U8519 (N_8519,N_4779,N_1638);
nand U8520 (N_8520,N_3921,N_333);
and U8521 (N_8521,N_3401,N_21);
nand U8522 (N_8522,N_1494,N_367);
or U8523 (N_8523,N_1662,N_3643);
or U8524 (N_8524,N_3137,N_2620);
nor U8525 (N_8525,N_4435,N_731);
and U8526 (N_8526,N_1255,N_4749);
and U8527 (N_8527,N_42,N_1292);
and U8528 (N_8528,N_3508,N_2103);
and U8529 (N_8529,N_578,N_4314);
nor U8530 (N_8530,N_316,N_3790);
nor U8531 (N_8531,N_506,N_549);
nor U8532 (N_8532,N_1492,N_3142);
nand U8533 (N_8533,N_4295,N_1006);
and U8534 (N_8534,N_49,N_2459);
and U8535 (N_8535,N_417,N_2769);
nor U8536 (N_8536,N_799,N_2621);
or U8537 (N_8537,N_4526,N_4415);
nand U8538 (N_8538,N_2631,N_1198);
or U8539 (N_8539,N_563,N_4918);
and U8540 (N_8540,N_1414,N_3026);
or U8541 (N_8541,N_1783,N_4912);
nor U8542 (N_8542,N_2682,N_1547);
or U8543 (N_8543,N_2550,N_931);
nor U8544 (N_8544,N_3244,N_2791);
or U8545 (N_8545,N_759,N_3493);
xnor U8546 (N_8546,N_2174,N_2731);
nor U8547 (N_8547,N_3208,N_1705);
nor U8548 (N_8548,N_751,N_1312);
nand U8549 (N_8549,N_3504,N_4201);
nand U8550 (N_8550,N_1778,N_2966);
nor U8551 (N_8551,N_765,N_2822);
or U8552 (N_8552,N_258,N_3997);
and U8553 (N_8553,N_1961,N_777);
nor U8554 (N_8554,N_4878,N_2413);
or U8555 (N_8555,N_3843,N_3163);
and U8556 (N_8556,N_2106,N_2565);
nand U8557 (N_8557,N_2923,N_3069);
nor U8558 (N_8558,N_317,N_2627);
nand U8559 (N_8559,N_397,N_2470);
nand U8560 (N_8560,N_4043,N_1104);
nor U8561 (N_8561,N_2675,N_1198);
nor U8562 (N_8562,N_2701,N_2743);
nand U8563 (N_8563,N_4511,N_1056);
nor U8564 (N_8564,N_178,N_2222);
nor U8565 (N_8565,N_3360,N_343);
nor U8566 (N_8566,N_3226,N_3685);
or U8567 (N_8567,N_4410,N_2064);
nor U8568 (N_8568,N_1863,N_3545);
and U8569 (N_8569,N_2475,N_879);
or U8570 (N_8570,N_1987,N_1502);
nor U8571 (N_8571,N_4191,N_3540);
nand U8572 (N_8572,N_2682,N_1695);
nor U8573 (N_8573,N_2653,N_2577);
nor U8574 (N_8574,N_2591,N_3135);
or U8575 (N_8575,N_2252,N_4723);
and U8576 (N_8576,N_1782,N_2812);
nand U8577 (N_8577,N_3704,N_1340);
nor U8578 (N_8578,N_3986,N_2645);
nand U8579 (N_8579,N_2591,N_4128);
nor U8580 (N_8580,N_2026,N_4747);
or U8581 (N_8581,N_609,N_1444);
nand U8582 (N_8582,N_225,N_296);
nand U8583 (N_8583,N_4014,N_1320);
nand U8584 (N_8584,N_1426,N_2426);
or U8585 (N_8585,N_3721,N_4271);
nand U8586 (N_8586,N_2350,N_1827);
or U8587 (N_8587,N_4595,N_4494);
and U8588 (N_8588,N_653,N_708);
xnor U8589 (N_8589,N_1757,N_2705);
nand U8590 (N_8590,N_192,N_1751);
and U8591 (N_8591,N_1754,N_4701);
nor U8592 (N_8592,N_2966,N_3026);
or U8593 (N_8593,N_2647,N_991);
nand U8594 (N_8594,N_4473,N_2648);
and U8595 (N_8595,N_4268,N_1226);
nand U8596 (N_8596,N_311,N_1213);
nand U8597 (N_8597,N_1925,N_429);
or U8598 (N_8598,N_3290,N_3244);
nor U8599 (N_8599,N_1819,N_3684);
and U8600 (N_8600,N_3981,N_2035);
and U8601 (N_8601,N_558,N_1772);
nand U8602 (N_8602,N_2244,N_3333);
or U8603 (N_8603,N_2562,N_1365);
nor U8604 (N_8604,N_3691,N_427);
or U8605 (N_8605,N_2364,N_3687);
nor U8606 (N_8606,N_1335,N_4076);
nand U8607 (N_8607,N_2297,N_2683);
nor U8608 (N_8608,N_247,N_3114);
or U8609 (N_8609,N_3876,N_3785);
nor U8610 (N_8610,N_2082,N_1844);
nand U8611 (N_8611,N_2215,N_1510);
nor U8612 (N_8612,N_670,N_1013);
and U8613 (N_8613,N_2619,N_1778);
nor U8614 (N_8614,N_1047,N_2137);
or U8615 (N_8615,N_1493,N_3512);
and U8616 (N_8616,N_1053,N_318);
nor U8617 (N_8617,N_3967,N_4445);
and U8618 (N_8618,N_2354,N_2260);
or U8619 (N_8619,N_3626,N_1265);
nand U8620 (N_8620,N_3997,N_3073);
and U8621 (N_8621,N_3186,N_333);
nand U8622 (N_8622,N_2906,N_679);
nor U8623 (N_8623,N_4364,N_2427);
nor U8624 (N_8624,N_734,N_4929);
and U8625 (N_8625,N_3701,N_1520);
nor U8626 (N_8626,N_2869,N_1436);
nor U8627 (N_8627,N_4229,N_2197);
xnor U8628 (N_8628,N_4441,N_4525);
nor U8629 (N_8629,N_4633,N_923);
or U8630 (N_8630,N_573,N_350);
nand U8631 (N_8631,N_3922,N_2058);
and U8632 (N_8632,N_3006,N_4931);
and U8633 (N_8633,N_857,N_240);
or U8634 (N_8634,N_4508,N_3958);
and U8635 (N_8635,N_3858,N_3675);
or U8636 (N_8636,N_4335,N_1230);
nor U8637 (N_8637,N_710,N_4722);
nand U8638 (N_8638,N_2199,N_4003);
and U8639 (N_8639,N_4381,N_3713);
or U8640 (N_8640,N_3422,N_1678);
and U8641 (N_8641,N_3190,N_458);
and U8642 (N_8642,N_4743,N_3607);
and U8643 (N_8643,N_2923,N_1490);
or U8644 (N_8644,N_3627,N_4452);
or U8645 (N_8645,N_3140,N_4751);
nand U8646 (N_8646,N_2750,N_3600);
nand U8647 (N_8647,N_4239,N_1976);
and U8648 (N_8648,N_1844,N_1931);
and U8649 (N_8649,N_4838,N_4994);
nor U8650 (N_8650,N_4987,N_29);
nand U8651 (N_8651,N_135,N_506);
nand U8652 (N_8652,N_2141,N_3275);
nand U8653 (N_8653,N_887,N_3966);
or U8654 (N_8654,N_4318,N_2781);
or U8655 (N_8655,N_2221,N_1176);
nand U8656 (N_8656,N_954,N_354);
and U8657 (N_8657,N_2214,N_4059);
nand U8658 (N_8658,N_2210,N_4120);
or U8659 (N_8659,N_3490,N_1222);
and U8660 (N_8660,N_553,N_3410);
and U8661 (N_8661,N_3671,N_481);
and U8662 (N_8662,N_3986,N_3649);
and U8663 (N_8663,N_4806,N_2614);
and U8664 (N_8664,N_3854,N_4222);
and U8665 (N_8665,N_812,N_2593);
nand U8666 (N_8666,N_1450,N_1938);
nand U8667 (N_8667,N_3411,N_3226);
nor U8668 (N_8668,N_1446,N_70);
nor U8669 (N_8669,N_4739,N_3966);
or U8670 (N_8670,N_4622,N_2515);
nor U8671 (N_8671,N_1507,N_2573);
and U8672 (N_8672,N_2072,N_2345);
and U8673 (N_8673,N_307,N_2332);
nand U8674 (N_8674,N_3702,N_560);
nor U8675 (N_8675,N_4796,N_3399);
nor U8676 (N_8676,N_3494,N_3580);
nor U8677 (N_8677,N_3313,N_1884);
or U8678 (N_8678,N_1136,N_3361);
nor U8679 (N_8679,N_4836,N_3628);
nand U8680 (N_8680,N_3378,N_2446);
or U8681 (N_8681,N_4400,N_4225);
nand U8682 (N_8682,N_4314,N_4951);
and U8683 (N_8683,N_3365,N_2865);
or U8684 (N_8684,N_1916,N_1370);
and U8685 (N_8685,N_890,N_3996);
nand U8686 (N_8686,N_4271,N_4752);
nand U8687 (N_8687,N_2070,N_2125);
nor U8688 (N_8688,N_4487,N_1254);
nor U8689 (N_8689,N_4290,N_4400);
nand U8690 (N_8690,N_607,N_2373);
and U8691 (N_8691,N_3684,N_1063);
or U8692 (N_8692,N_4597,N_3850);
and U8693 (N_8693,N_2015,N_1201);
and U8694 (N_8694,N_312,N_2310);
and U8695 (N_8695,N_161,N_2625);
or U8696 (N_8696,N_3408,N_2152);
and U8697 (N_8697,N_3626,N_3387);
and U8698 (N_8698,N_4317,N_1098);
or U8699 (N_8699,N_3473,N_4402);
and U8700 (N_8700,N_1984,N_528);
and U8701 (N_8701,N_4107,N_2955);
nand U8702 (N_8702,N_3364,N_1647);
nor U8703 (N_8703,N_3797,N_745);
and U8704 (N_8704,N_1922,N_4712);
or U8705 (N_8705,N_2606,N_2798);
nor U8706 (N_8706,N_3142,N_239);
and U8707 (N_8707,N_2786,N_1240);
and U8708 (N_8708,N_356,N_798);
xnor U8709 (N_8709,N_4576,N_1674);
or U8710 (N_8710,N_93,N_1882);
and U8711 (N_8711,N_230,N_1124);
and U8712 (N_8712,N_4336,N_2774);
nor U8713 (N_8713,N_2442,N_1892);
nor U8714 (N_8714,N_3939,N_1532);
or U8715 (N_8715,N_988,N_606);
or U8716 (N_8716,N_1921,N_2393);
and U8717 (N_8717,N_4408,N_1877);
and U8718 (N_8718,N_2372,N_4339);
nand U8719 (N_8719,N_4940,N_1920);
nor U8720 (N_8720,N_2464,N_4721);
nand U8721 (N_8721,N_330,N_4895);
nor U8722 (N_8722,N_4734,N_324);
nand U8723 (N_8723,N_4544,N_1238);
and U8724 (N_8724,N_2536,N_3907);
or U8725 (N_8725,N_159,N_2388);
nand U8726 (N_8726,N_4909,N_4057);
nor U8727 (N_8727,N_2585,N_2002);
and U8728 (N_8728,N_4797,N_1915);
nor U8729 (N_8729,N_1734,N_749);
nand U8730 (N_8730,N_4356,N_3283);
nor U8731 (N_8731,N_1165,N_1870);
nor U8732 (N_8732,N_3551,N_1235);
nand U8733 (N_8733,N_2650,N_2876);
or U8734 (N_8734,N_56,N_1092);
nand U8735 (N_8735,N_1422,N_368);
and U8736 (N_8736,N_4270,N_1491);
nand U8737 (N_8737,N_1679,N_3162);
or U8738 (N_8738,N_3952,N_3711);
and U8739 (N_8739,N_3114,N_4315);
and U8740 (N_8740,N_2609,N_3010);
or U8741 (N_8741,N_3098,N_3664);
nand U8742 (N_8742,N_1238,N_1335);
nor U8743 (N_8743,N_3851,N_1837);
and U8744 (N_8744,N_4546,N_49);
or U8745 (N_8745,N_2334,N_2676);
nand U8746 (N_8746,N_1738,N_1232);
nor U8747 (N_8747,N_4928,N_3354);
or U8748 (N_8748,N_951,N_3830);
and U8749 (N_8749,N_3600,N_1482);
and U8750 (N_8750,N_3697,N_3573);
nor U8751 (N_8751,N_3063,N_3033);
or U8752 (N_8752,N_1414,N_2440);
or U8753 (N_8753,N_2070,N_4883);
nor U8754 (N_8754,N_1626,N_624);
nor U8755 (N_8755,N_4734,N_4589);
and U8756 (N_8756,N_3344,N_4246);
nor U8757 (N_8757,N_3205,N_371);
nor U8758 (N_8758,N_1422,N_1386);
nand U8759 (N_8759,N_4696,N_1972);
nor U8760 (N_8760,N_1595,N_1953);
or U8761 (N_8761,N_1068,N_4732);
or U8762 (N_8762,N_1286,N_1987);
nor U8763 (N_8763,N_4528,N_4213);
and U8764 (N_8764,N_3732,N_4620);
and U8765 (N_8765,N_1280,N_4738);
nand U8766 (N_8766,N_2874,N_1701);
or U8767 (N_8767,N_4453,N_2742);
and U8768 (N_8768,N_1781,N_587);
and U8769 (N_8769,N_4866,N_3624);
nand U8770 (N_8770,N_2130,N_4552);
or U8771 (N_8771,N_4164,N_3551);
nor U8772 (N_8772,N_2221,N_542);
or U8773 (N_8773,N_124,N_1251);
nand U8774 (N_8774,N_270,N_3392);
nand U8775 (N_8775,N_1796,N_2209);
xor U8776 (N_8776,N_1848,N_1452);
and U8777 (N_8777,N_3329,N_4448);
nor U8778 (N_8778,N_1444,N_4808);
nand U8779 (N_8779,N_2055,N_3854);
nor U8780 (N_8780,N_3990,N_4460);
and U8781 (N_8781,N_3858,N_569);
nand U8782 (N_8782,N_4798,N_4426);
nor U8783 (N_8783,N_2215,N_2685);
and U8784 (N_8784,N_371,N_141);
xnor U8785 (N_8785,N_717,N_571);
nand U8786 (N_8786,N_419,N_637);
nand U8787 (N_8787,N_1699,N_4372);
xnor U8788 (N_8788,N_3760,N_3665);
nand U8789 (N_8789,N_4694,N_2057);
nand U8790 (N_8790,N_582,N_2946);
and U8791 (N_8791,N_47,N_402);
nor U8792 (N_8792,N_2305,N_422);
and U8793 (N_8793,N_467,N_2189);
and U8794 (N_8794,N_907,N_3027);
or U8795 (N_8795,N_3075,N_4944);
or U8796 (N_8796,N_531,N_792);
nand U8797 (N_8797,N_3481,N_3523);
or U8798 (N_8798,N_272,N_506);
nand U8799 (N_8799,N_2914,N_1933);
nand U8800 (N_8800,N_152,N_1374);
nand U8801 (N_8801,N_59,N_633);
and U8802 (N_8802,N_17,N_3916);
nor U8803 (N_8803,N_4298,N_410);
or U8804 (N_8804,N_4052,N_1910);
xor U8805 (N_8805,N_1166,N_620);
nor U8806 (N_8806,N_4868,N_1408);
nor U8807 (N_8807,N_51,N_4771);
and U8808 (N_8808,N_1946,N_3482);
and U8809 (N_8809,N_1690,N_1021);
or U8810 (N_8810,N_3756,N_3738);
nor U8811 (N_8811,N_1225,N_2702);
or U8812 (N_8812,N_828,N_1290);
and U8813 (N_8813,N_1810,N_4173);
and U8814 (N_8814,N_3633,N_1336);
and U8815 (N_8815,N_245,N_3189);
nand U8816 (N_8816,N_3002,N_2604);
and U8817 (N_8817,N_2979,N_4238);
nor U8818 (N_8818,N_2403,N_4093);
nand U8819 (N_8819,N_4410,N_4231);
and U8820 (N_8820,N_4857,N_1648);
or U8821 (N_8821,N_1332,N_1878);
nand U8822 (N_8822,N_203,N_1031);
nor U8823 (N_8823,N_139,N_1638);
nor U8824 (N_8824,N_3078,N_468);
or U8825 (N_8825,N_2641,N_3768);
or U8826 (N_8826,N_3039,N_839);
nor U8827 (N_8827,N_2605,N_1255);
and U8828 (N_8828,N_7,N_19);
or U8829 (N_8829,N_1136,N_932);
nand U8830 (N_8830,N_705,N_25);
nand U8831 (N_8831,N_1061,N_4514);
and U8832 (N_8832,N_1276,N_3405);
nand U8833 (N_8833,N_1879,N_4216);
nor U8834 (N_8834,N_3509,N_1185);
and U8835 (N_8835,N_1417,N_4295);
nor U8836 (N_8836,N_2367,N_4975);
nor U8837 (N_8837,N_2069,N_4654);
and U8838 (N_8838,N_2493,N_4878);
or U8839 (N_8839,N_3022,N_4427);
nand U8840 (N_8840,N_4302,N_4026);
nor U8841 (N_8841,N_3830,N_1153);
or U8842 (N_8842,N_4045,N_1431);
or U8843 (N_8843,N_2703,N_1353);
and U8844 (N_8844,N_3855,N_4742);
or U8845 (N_8845,N_3427,N_3793);
and U8846 (N_8846,N_3597,N_3854);
and U8847 (N_8847,N_888,N_2543);
nor U8848 (N_8848,N_4796,N_3340);
or U8849 (N_8849,N_1263,N_500);
or U8850 (N_8850,N_570,N_4869);
nand U8851 (N_8851,N_2092,N_309);
or U8852 (N_8852,N_67,N_3171);
xnor U8853 (N_8853,N_2998,N_1920);
and U8854 (N_8854,N_341,N_1087);
nand U8855 (N_8855,N_4593,N_3612);
or U8856 (N_8856,N_381,N_2106);
nand U8857 (N_8857,N_2203,N_4766);
or U8858 (N_8858,N_1732,N_2888);
and U8859 (N_8859,N_2216,N_1356);
nor U8860 (N_8860,N_2840,N_636);
nand U8861 (N_8861,N_4396,N_367);
or U8862 (N_8862,N_1820,N_2414);
and U8863 (N_8863,N_2,N_4229);
nor U8864 (N_8864,N_3890,N_4238);
nand U8865 (N_8865,N_4858,N_3498);
nand U8866 (N_8866,N_4581,N_1817);
nand U8867 (N_8867,N_1120,N_1876);
nor U8868 (N_8868,N_4638,N_715);
nand U8869 (N_8869,N_2396,N_632);
and U8870 (N_8870,N_968,N_3417);
or U8871 (N_8871,N_2225,N_2937);
nand U8872 (N_8872,N_2549,N_3185);
nor U8873 (N_8873,N_2256,N_1728);
nand U8874 (N_8874,N_821,N_1036);
or U8875 (N_8875,N_1984,N_742);
nand U8876 (N_8876,N_2783,N_2764);
or U8877 (N_8877,N_4419,N_2481);
nand U8878 (N_8878,N_3793,N_175);
nor U8879 (N_8879,N_2596,N_4141);
nand U8880 (N_8880,N_4738,N_2628);
nor U8881 (N_8881,N_952,N_3236);
or U8882 (N_8882,N_1619,N_1906);
nor U8883 (N_8883,N_3895,N_1803);
nand U8884 (N_8884,N_4797,N_1896);
or U8885 (N_8885,N_3616,N_2611);
nor U8886 (N_8886,N_3831,N_4272);
nand U8887 (N_8887,N_471,N_3626);
or U8888 (N_8888,N_585,N_3208);
nand U8889 (N_8889,N_588,N_1329);
and U8890 (N_8890,N_3971,N_1530);
and U8891 (N_8891,N_2199,N_3134);
and U8892 (N_8892,N_956,N_4101);
and U8893 (N_8893,N_2737,N_4590);
and U8894 (N_8894,N_2337,N_696);
nor U8895 (N_8895,N_3508,N_2918);
nor U8896 (N_8896,N_1819,N_71);
nand U8897 (N_8897,N_4218,N_1359);
nor U8898 (N_8898,N_3454,N_1255);
nor U8899 (N_8899,N_779,N_3208);
and U8900 (N_8900,N_1339,N_2377);
nor U8901 (N_8901,N_899,N_1408);
and U8902 (N_8902,N_4861,N_2904);
nor U8903 (N_8903,N_3050,N_795);
and U8904 (N_8904,N_376,N_4189);
nor U8905 (N_8905,N_1151,N_1092);
nor U8906 (N_8906,N_2391,N_782);
nand U8907 (N_8907,N_3789,N_292);
nor U8908 (N_8908,N_524,N_1123);
or U8909 (N_8909,N_539,N_681);
nor U8910 (N_8910,N_2757,N_4170);
or U8911 (N_8911,N_2679,N_1688);
and U8912 (N_8912,N_4576,N_539);
or U8913 (N_8913,N_1238,N_1791);
nor U8914 (N_8914,N_1878,N_4982);
nor U8915 (N_8915,N_1537,N_306);
xnor U8916 (N_8916,N_2296,N_2339);
nand U8917 (N_8917,N_1205,N_2195);
xnor U8918 (N_8918,N_3327,N_338);
and U8919 (N_8919,N_4459,N_2371);
and U8920 (N_8920,N_462,N_3323);
or U8921 (N_8921,N_327,N_328);
nand U8922 (N_8922,N_4452,N_318);
nor U8923 (N_8923,N_1912,N_1244);
nor U8924 (N_8924,N_3634,N_4495);
and U8925 (N_8925,N_4954,N_4834);
nand U8926 (N_8926,N_1376,N_4582);
or U8927 (N_8927,N_1795,N_4451);
xor U8928 (N_8928,N_1195,N_125);
or U8929 (N_8929,N_4993,N_118);
or U8930 (N_8930,N_2716,N_1503);
nor U8931 (N_8931,N_1795,N_3955);
nand U8932 (N_8932,N_1266,N_1132);
nand U8933 (N_8933,N_3930,N_1263);
nand U8934 (N_8934,N_1056,N_1088);
nand U8935 (N_8935,N_1983,N_3058);
nor U8936 (N_8936,N_1765,N_2422);
nand U8937 (N_8937,N_3940,N_4224);
nand U8938 (N_8938,N_4326,N_1576);
or U8939 (N_8939,N_1936,N_2702);
nor U8940 (N_8940,N_1802,N_1567);
nor U8941 (N_8941,N_2194,N_3871);
nor U8942 (N_8942,N_3549,N_683);
and U8943 (N_8943,N_3342,N_3368);
or U8944 (N_8944,N_2885,N_4436);
and U8945 (N_8945,N_836,N_4334);
and U8946 (N_8946,N_2931,N_308);
or U8947 (N_8947,N_4543,N_3992);
nand U8948 (N_8948,N_2240,N_4144);
nand U8949 (N_8949,N_3254,N_4868);
nor U8950 (N_8950,N_2709,N_3362);
nor U8951 (N_8951,N_644,N_805);
nor U8952 (N_8952,N_4106,N_568);
and U8953 (N_8953,N_2569,N_4533);
and U8954 (N_8954,N_315,N_1716);
or U8955 (N_8955,N_4700,N_3312);
and U8956 (N_8956,N_4734,N_2952);
or U8957 (N_8957,N_2792,N_4552);
and U8958 (N_8958,N_1425,N_1682);
nand U8959 (N_8959,N_4695,N_1963);
and U8960 (N_8960,N_499,N_2185);
nand U8961 (N_8961,N_2610,N_534);
nor U8962 (N_8962,N_1910,N_525);
nand U8963 (N_8963,N_1393,N_1923);
nand U8964 (N_8964,N_1571,N_4871);
or U8965 (N_8965,N_407,N_4221);
nand U8966 (N_8966,N_4722,N_565);
or U8967 (N_8967,N_1279,N_915);
nand U8968 (N_8968,N_1312,N_1449);
nand U8969 (N_8969,N_4827,N_4811);
nor U8970 (N_8970,N_3555,N_2310);
nor U8971 (N_8971,N_341,N_2588);
and U8972 (N_8972,N_1670,N_1275);
nor U8973 (N_8973,N_3176,N_4163);
nand U8974 (N_8974,N_3700,N_2800);
and U8975 (N_8975,N_2710,N_1463);
nand U8976 (N_8976,N_877,N_4926);
and U8977 (N_8977,N_2919,N_431);
and U8978 (N_8978,N_2512,N_2164);
nor U8979 (N_8979,N_1869,N_465);
and U8980 (N_8980,N_2501,N_4549);
nand U8981 (N_8981,N_4787,N_441);
and U8982 (N_8982,N_2234,N_299);
nor U8983 (N_8983,N_3723,N_4257);
or U8984 (N_8984,N_1371,N_4108);
or U8985 (N_8985,N_1143,N_1678);
and U8986 (N_8986,N_4803,N_1669);
or U8987 (N_8987,N_4268,N_3792);
and U8988 (N_8988,N_1499,N_1988);
and U8989 (N_8989,N_2419,N_4117);
and U8990 (N_8990,N_4907,N_2931);
nor U8991 (N_8991,N_191,N_2160);
nor U8992 (N_8992,N_4725,N_951);
or U8993 (N_8993,N_829,N_966);
nand U8994 (N_8994,N_3298,N_3997);
nor U8995 (N_8995,N_4617,N_3187);
or U8996 (N_8996,N_3753,N_1665);
nor U8997 (N_8997,N_241,N_1454);
nor U8998 (N_8998,N_4214,N_3012);
xor U8999 (N_8999,N_2433,N_3217);
nor U9000 (N_9000,N_4967,N_2695);
or U9001 (N_9001,N_1196,N_2426);
nand U9002 (N_9002,N_4060,N_2418);
nand U9003 (N_9003,N_2264,N_2513);
xnor U9004 (N_9004,N_3843,N_2488);
or U9005 (N_9005,N_3655,N_1743);
nand U9006 (N_9006,N_4069,N_2801);
and U9007 (N_9007,N_2706,N_1042);
and U9008 (N_9008,N_3866,N_4119);
and U9009 (N_9009,N_898,N_404);
and U9010 (N_9010,N_2058,N_863);
and U9011 (N_9011,N_1510,N_3594);
nand U9012 (N_9012,N_4555,N_1725);
and U9013 (N_9013,N_262,N_4751);
nor U9014 (N_9014,N_1859,N_3716);
nand U9015 (N_9015,N_832,N_393);
nor U9016 (N_9016,N_2329,N_4701);
and U9017 (N_9017,N_2475,N_136);
or U9018 (N_9018,N_2487,N_3936);
nand U9019 (N_9019,N_335,N_3388);
nor U9020 (N_9020,N_1961,N_3763);
or U9021 (N_9021,N_440,N_3016);
or U9022 (N_9022,N_2652,N_707);
nand U9023 (N_9023,N_4872,N_2905);
nor U9024 (N_9024,N_1518,N_516);
and U9025 (N_9025,N_1459,N_1476);
nor U9026 (N_9026,N_511,N_2797);
and U9027 (N_9027,N_1958,N_2880);
nor U9028 (N_9028,N_1906,N_4334);
nand U9029 (N_9029,N_4867,N_2091);
nand U9030 (N_9030,N_279,N_4384);
nand U9031 (N_9031,N_1973,N_2433);
nor U9032 (N_9032,N_3405,N_493);
or U9033 (N_9033,N_1011,N_4962);
nor U9034 (N_9034,N_4012,N_3687);
and U9035 (N_9035,N_4852,N_2612);
or U9036 (N_9036,N_3854,N_4800);
or U9037 (N_9037,N_4051,N_923);
or U9038 (N_9038,N_4853,N_266);
nand U9039 (N_9039,N_1949,N_2197);
and U9040 (N_9040,N_2291,N_3295);
or U9041 (N_9041,N_3839,N_2003);
or U9042 (N_9042,N_4649,N_4165);
and U9043 (N_9043,N_4435,N_59);
nor U9044 (N_9044,N_3341,N_3553);
xor U9045 (N_9045,N_2046,N_126);
nand U9046 (N_9046,N_658,N_2951);
nand U9047 (N_9047,N_3048,N_4236);
nand U9048 (N_9048,N_3623,N_2739);
and U9049 (N_9049,N_2335,N_2437);
and U9050 (N_9050,N_1801,N_4618);
or U9051 (N_9051,N_4481,N_555);
and U9052 (N_9052,N_4350,N_4271);
nor U9053 (N_9053,N_2200,N_3816);
nand U9054 (N_9054,N_675,N_4914);
xor U9055 (N_9055,N_16,N_2824);
nand U9056 (N_9056,N_3850,N_3729);
and U9057 (N_9057,N_1410,N_3459);
nand U9058 (N_9058,N_951,N_4996);
and U9059 (N_9059,N_2945,N_1020);
nor U9060 (N_9060,N_2247,N_1597);
nor U9061 (N_9061,N_2950,N_1694);
and U9062 (N_9062,N_977,N_3046);
nor U9063 (N_9063,N_3032,N_3156);
nand U9064 (N_9064,N_3060,N_1231);
nor U9065 (N_9065,N_3148,N_510);
and U9066 (N_9066,N_4345,N_2394);
nor U9067 (N_9067,N_3256,N_3419);
or U9068 (N_9068,N_2799,N_232);
nor U9069 (N_9069,N_929,N_612);
nand U9070 (N_9070,N_179,N_2456);
or U9071 (N_9071,N_4631,N_3961);
xnor U9072 (N_9072,N_513,N_1879);
and U9073 (N_9073,N_737,N_4537);
and U9074 (N_9074,N_3729,N_2841);
nor U9075 (N_9075,N_4708,N_4380);
nor U9076 (N_9076,N_2261,N_1508);
and U9077 (N_9077,N_427,N_3885);
or U9078 (N_9078,N_4144,N_2749);
nor U9079 (N_9079,N_2558,N_2679);
and U9080 (N_9080,N_2620,N_281);
or U9081 (N_9081,N_3089,N_4126);
or U9082 (N_9082,N_3684,N_3775);
and U9083 (N_9083,N_3806,N_3571);
or U9084 (N_9084,N_1575,N_4531);
or U9085 (N_9085,N_4569,N_1627);
and U9086 (N_9086,N_1589,N_1006);
nand U9087 (N_9087,N_2974,N_2070);
or U9088 (N_9088,N_3518,N_2019);
and U9089 (N_9089,N_3994,N_961);
or U9090 (N_9090,N_2670,N_2999);
or U9091 (N_9091,N_4672,N_1006);
or U9092 (N_9092,N_374,N_2062);
xor U9093 (N_9093,N_4726,N_2330);
xor U9094 (N_9094,N_1663,N_1222);
and U9095 (N_9095,N_1236,N_3521);
xor U9096 (N_9096,N_2441,N_1999);
or U9097 (N_9097,N_2179,N_4210);
nor U9098 (N_9098,N_1844,N_2011);
nand U9099 (N_9099,N_1952,N_1979);
or U9100 (N_9100,N_1791,N_4681);
nand U9101 (N_9101,N_1820,N_3006);
and U9102 (N_9102,N_3437,N_1);
nor U9103 (N_9103,N_515,N_1778);
and U9104 (N_9104,N_4510,N_4899);
or U9105 (N_9105,N_141,N_2558);
nand U9106 (N_9106,N_490,N_115);
nor U9107 (N_9107,N_4754,N_4749);
or U9108 (N_9108,N_12,N_4296);
or U9109 (N_9109,N_1827,N_57);
nor U9110 (N_9110,N_3485,N_662);
nand U9111 (N_9111,N_4676,N_1982);
and U9112 (N_9112,N_1447,N_737);
nand U9113 (N_9113,N_3314,N_4846);
nor U9114 (N_9114,N_3644,N_3234);
nand U9115 (N_9115,N_367,N_3961);
or U9116 (N_9116,N_2493,N_970);
and U9117 (N_9117,N_1440,N_4137);
and U9118 (N_9118,N_4331,N_4050);
and U9119 (N_9119,N_2142,N_1439);
and U9120 (N_9120,N_2672,N_2867);
nand U9121 (N_9121,N_4738,N_3101);
nand U9122 (N_9122,N_2243,N_937);
or U9123 (N_9123,N_3907,N_437);
or U9124 (N_9124,N_142,N_2037);
nand U9125 (N_9125,N_3451,N_3813);
nand U9126 (N_9126,N_609,N_3486);
nand U9127 (N_9127,N_1400,N_3932);
or U9128 (N_9128,N_1905,N_360);
and U9129 (N_9129,N_263,N_4130);
and U9130 (N_9130,N_2693,N_1031);
nand U9131 (N_9131,N_4789,N_1539);
and U9132 (N_9132,N_1567,N_1559);
nand U9133 (N_9133,N_3086,N_1742);
or U9134 (N_9134,N_3577,N_2220);
or U9135 (N_9135,N_1158,N_338);
and U9136 (N_9136,N_2366,N_2603);
nand U9137 (N_9137,N_3312,N_1055);
nand U9138 (N_9138,N_626,N_587);
nand U9139 (N_9139,N_3164,N_4244);
nand U9140 (N_9140,N_1737,N_1235);
or U9141 (N_9141,N_3353,N_4815);
nor U9142 (N_9142,N_2321,N_3038);
and U9143 (N_9143,N_4445,N_165);
and U9144 (N_9144,N_3119,N_4724);
or U9145 (N_9145,N_4987,N_2965);
nand U9146 (N_9146,N_1170,N_4862);
nor U9147 (N_9147,N_4112,N_4351);
nand U9148 (N_9148,N_744,N_1952);
nand U9149 (N_9149,N_2065,N_1865);
and U9150 (N_9150,N_3987,N_1383);
and U9151 (N_9151,N_1205,N_4761);
nand U9152 (N_9152,N_2757,N_3134);
or U9153 (N_9153,N_1305,N_4789);
nor U9154 (N_9154,N_207,N_4002);
xnor U9155 (N_9155,N_1624,N_874);
nand U9156 (N_9156,N_1964,N_3208);
or U9157 (N_9157,N_3558,N_2910);
nor U9158 (N_9158,N_2928,N_1060);
nor U9159 (N_9159,N_87,N_1401);
xnor U9160 (N_9160,N_4633,N_841);
and U9161 (N_9161,N_2353,N_821);
and U9162 (N_9162,N_4698,N_209);
nand U9163 (N_9163,N_4366,N_447);
and U9164 (N_9164,N_3194,N_3062);
and U9165 (N_9165,N_1457,N_4531);
and U9166 (N_9166,N_2795,N_4061);
and U9167 (N_9167,N_1177,N_3);
or U9168 (N_9168,N_4529,N_151);
or U9169 (N_9169,N_4512,N_1198);
and U9170 (N_9170,N_4441,N_2473);
or U9171 (N_9171,N_3342,N_1797);
xnor U9172 (N_9172,N_942,N_3858);
nand U9173 (N_9173,N_2217,N_4588);
nand U9174 (N_9174,N_9,N_4864);
or U9175 (N_9175,N_3305,N_4713);
and U9176 (N_9176,N_1503,N_1510);
or U9177 (N_9177,N_4550,N_57);
nand U9178 (N_9178,N_4777,N_3816);
or U9179 (N_9179,N_4632,N_1674);
nand U9180 (N_9180,N_368,N_782);
and U9181 (N_9181,N_1909,N_4619);
or U9182 (N_9182,N_2370,N_2048);
nor U9183 (N_9183,N_4044,N_4473);
nor U9184 (N_9184,N_4276,N_1336);
and U9185 (N_9185,N_4421,N_666);
nand U9186 (N_9186,N_863,N_2070);
nand U9187 (N_9187,N_2289,N_4317);
or U9188 (N_9188,N_4620,N_1586);
nor U9189 (N_9189,N_2865,N_4628);
nor U9190 (N_9190,N_4500,N_4957);
nand U9191 (N_9191,N_4439,N_12);
and U9192 (N_9192,N_995,N_3646);
and U9193 (N_9193,N_1688,N_2857);
and U9194 (N_9194,N_1284,N_2378);
and U9195 (N_9195,N_2662,N_141);
nand U9196 (N_9196,N_832,N_4472);
nor U9197 (N_9197,N_2170,N_529);
xnor U9198 (N_9198,N_3450,N_1759);
nand U9199 (N_9199,N_1063,N_1496);
or U9200 (N_9200,N_716,N_57);
nand U9201 (N_9201,N_1069,N_4352);
nor U9202 (N_9202,N_1304,N_3790);
nor U9203 (N_9203,N_1745,N_4216);
nand U9204 (N_9204,N_4010,N_4085);
nand U9205 (N_9205,N_4108,N_4196);
and U9206 (N_9206,N_2835,N_4606);
and U9207 (N_9207,N_3355,N_224);
nand U9208 (N_9208,N_3526,N_3870);
and U9209 (N_9209,N_1644,N_4064);
nor U9210 (N_9210,N_3870,N_368);
nor U9211 (N_9211,N_2830,N_1377);
nor U9212 (N_9212,N_1109,N_4741);
and U9213 (N_9213,N_3592,N_1288);
and U9214 (N_9214,N_4491,N_2796);
or U9215 (N_9215,N_2113,N_2105);
and U9216 (N_9216,N_4986,N_3313);
or U9217 (N_9217,N_219,N_2891);
nand U9218 (N_9218,N_4326,N_524);
and U9219 (N_9219,N_1245,N_3950);
and U9220 (N_9220,N_4157,N_3008);
and U9221 (N_9221,N_3575,N_501);
nand U9222 (N_9222,N_3899,N_4577);
nand U9223 (N_9223,N_4719,N_4615);
or U9224 (N_9224,N_1488,N_2015);
nand U9225 (N_9225,N_4606,N_1767);
or U9226 (N_9226,N_305,N_4187);
nand U9227 (N_9227,N_664,N_1969);
or U9228 (N_9228,N_1568,N_649);
xor U9229 (N_9229,N_2469,N_2334);
nand U9230 (N_9230,N_297,N_2777);
nor U9231 (N_9231,N_3364,N_699);
xnor U9232 (N_9232,N_71,N_2945);
nand U9233 (N_9233,N_2961,N_2739);
nand U9234 (N_9234,N_2000,N_2903);
or U9235 (N_9235,N_2138,N_3275);
or U9236 (N_9236,N_620,N_2997);
nor U9237 (N_9237,N_3608,N_777);
or U9238 (N_9238,N_431,N_4418);
nand U9239 (N_9239,N_1042,N_3858);
and U9240 (N_9240,N_4980,N_2186);
nor U9241 (N_9241,N_1682,N_314);
or U9242 (N_9242,N_1868,N_1063);
nand U9243 (N_9243,N_2819,N_4328);
or U9244 (N_9244,N_2652,N_3016);
nand U9245 (N_9245,N_4583,N_1664);
nand U9246 (N_9246,N_789,N_206);
and U9247 (N_9247,N_3882,N_592);
and U9248 (N_9248,N_569,N_49);
and U9249 (N_9249,N_174,N_4222);
nor U9250 (N_9250,N_1636,N_4619);
and U9251 (N_9251,N_4456,N_3733);
nand U9252 (N_9252,N_1806,N_3325);
nor U9253 (N_9253,N_4221,N_3623);
or U9254 (N_9254,N_3812,N_3758);
and U9255 (N_9255,N_3588,N_4076);
and U9256 (N_9256,N_4431,N_3592);
and U9257 (N_9257,N_2502,N_1685);
or U9258 (N_9258,N_3107,N_822);
and U9259 (N_9259,N_2882,N_4733);
and U9260 (N_9260,N_1833,N_3074);
nor U9261 (N_9261,N_4103,N_4613);
nand U9262 (N_9262,N_4392,N_2258);
or U9263 (N_9263,N_4130,N_2931);
or U9264 (N_9264,N_4730,N_2428);
nor U9265 (N_9265,N_2221,N_242);
nor U9266 (N_9266,N_3534,N_1372);
or U9267 (N_9267,N_4603,N_3029);
and U9268 (N_9268,N_891,N_4037);
or U9269 (N_9269,N_2181,N_1380);
nor U9270 (N_9270,N_1329,N_2114);
nor U9271 (N_9271,N_2761,N_1407);
nand U9272 (N_9272,N_2034,N_3990);
or U9273 (N_9273,N_1237,N_700);
nand U9274 (N_9274,N_1259,N_1581);
or U9275 (N_9275,N_3870,N_3336);
nor U9276 (N_9276,N_891,N_3940);
and U9277 (N_9277,N_2777,N_2017);
nand U9278 (N_9278,N_4116,N_4223);
nor U9279 (N_9279,N_2019,N_4450);
nand U9280 (N_9280,N_2093,N_1472);
and U9281 (N_9281,N_4898,N_1099);
or U9282 (N_9282,N_3291,N_4040);
and U9283 (N_9283,N_4615,N_4383);
nor U9284 (N_9284,N_1049,N_2569);
and U9285 (N_9285,N_3864,N_94);
xor U9286 (N_9286,N_1294,N_4030);
and U9287 (N_9287,N_4593,N_1704);
nor U9288 (N_9288,N_1077,N_3910);
and U9289 (N_9289,N_2222,N_3125);
or U9290 (N_9290,N_288,N_1806);
nand U9291 (N_9291,N_4890,N_2410);
or U9292 (N_9292,N_2336,N_1519);
nor U9293 (N_9293,N_611,N_4189);
nor U9294 (N_9294,N_3270,N_3029);
nor U9295 (N_9295,N_3590,N_3741);
or U9296 (N_9296,N_535,N_835);
or U9297 (N_9297,N_4860,N_3994);
and U9298 (N_9298,N_149,N_1146);
or U9299 (N_9299,N_3307,N_3741);
or U9300 (N_9300,N_191,N_4014);
nor U9301 (N_9301,N_3843,N_1091);
xnor U9302 (N_9302,N_479,N_1921);
nand U9303 (N_9303,N_1496,N_4124);
or U9304 (N_9304,N_2206,N_1437);
nor U9305 (N_9305,N_3005,N_3360);
nand U9306 (N_9306,N_856,N_2429);
nand U9307 (N_9307,N_2516,N_2603);
nor U9308 (N_9308,N_4835,N_32);
or U9309 (N_9309,N_4100,N_123);
nand U9310 (N_9310,N_4029,N_3664);
and U9311 (N_9311,N_1077,N_1308);
nor U9312 (N_9312,N_3390,N_563);
or U9313 (N_9313,N_4705,N_3871);
or U9314 (N_9314,N_1355,N_3099);
and U9315 (N_9315,N_1229,N_4505);
and U9316 (N_9316,N_4632,N_1070);
nand U9317 (N_9317,N_1390,N_329);
or U9318 (N_9318,N_2446,N_2471);
nand U9319 (N_9319,N_3249,N_2262);
and U9320 (N_9320,N_550,N_3310);
or U9321 (N_9321,N_1850,N_3180);
nor U9322 (N_9322,N_2123,N_4239);
nand U9323 (N_9323,N_4247,N_550);
xor U9324 (N_9324,N_2661,N_3713);
nor U9325 (N_9325,N_4107,N_430);
and U9326 (N_9326,N_3682,N_204);
nand U9327 (N_9327,N_2417,N_3559);
and U9328 (N_9328,N_2742,N_1273);
nor U9329 (N_9329,N_2780,N_4383);
nand U9330 (N_9330,N_3168,N_27);
nor U9331 (N_9331,N_4954,N_1882);
nor U9332 (N_9332,N_4410,N_4868);
nor U9333 (N_9333,N_80,N_225);
and U9334 (N_9334,N_2099,N_612);
nor U9335 (N_9335,N_4303,N_4753);
or U9336 (N_9336,N_2612,N_2441);
nor U9337 (N_9337,N_3113,N_2212);
and U9338 (N_9338,N_2476,N_904);
xnor U9339 (N_9339,N_3362,N_912);
nor U9340 (N_9340,N_1104,N_4159);
or U9341 (N_9341,N_3453,N_1429);
and U9342 (N_9342,N_2271,N_4157);
xnor U9343 (N_9343,N_3935,N_1519);
nand U9344 (N_9344,N_4603,N_4130);
nor U9345 (N_9345,N_2561,N_2445);
and U9346 (N_9346,N_4045,N_4270);
and U9347 (N_9347,N_188,N_3871);
or U9348 (N_9348,N_670,N_3826);
nor U9349 (N_9349,N_3704,N_863);
xnor U9350 (N_9350,N_408,N_2249);
and U9351 (N_9351,N_2730,N_966);
xnor U9352 (N_9352,N_1249,N_4133);
and U9353 (N_9353,N_4727,N_4171);
nor U9354 (N_9354,N_3571,N_866);
or U9355 (N_9355,N_321,N_2806);
and U9356 (N_9356,N_3444,N_4239);
or U9357 (N_9357,N_4159,N_125);
and U9358 (N_9358,N_2272,N_4578);
and U9359 (N_9359,N_2366,N_3260);
and U9360 (N_9360,N_466,N_3849);
and U9361 (N_9361,N_3432,N_2589);
nor U9362 (N_9362,N_874,N_1354);
nand U9363 (N_9363,N_2151,N_1397);
and U9364 (N_9364,N_2473,N_3369);
or U9365 (N_9365,N_1386,N_694);
nor U9366 (N_9366,N_3586,N_1773);
xor U9367 (N_9367,N_1138,N_1480);
nand U9368 (N_9368,N_955,N_550);
nor U9369 (N_9369,N_1328,N_4231);
nand U9370 (N_9370,N_1041,N_829);
nand U9371 (N_9371,N_4536,N_2788);
nand U9372 (N_9372,N_191,N_1368);
and U9373 (N_9373,N_1584,N_4637);
or U9374 (N_9374,N_3899,N_2495);
and U9375 (N_9375,N_1857,N_4715);
and U9376 (N_9376,N_873,N_1493);
nor U9377 (N_9377,N_1206,N_4083);
nor U9378 (N_9378,N_1969,N_4145);
and U9379 (N_9379,N_4989,N_1497);
nor U9380 (N_9380,N_2450,N_719);
nand U9381 (N_9381,N_3913,N_4983);
and U9382 (N_9382,N_1873,N_3795);
nor U9383 (N_9383,N_869,N_2347);
nor U9384 (N_9384,N_1225,N_4424);
nor U9385 (N_9385,N_1611,N_2610);
nor U9386 (N_9386,N_2764,N_2924);
or U9387 (N_9387,N_2535,N_116);
and U9388 (N_9388,N_781,N_2339);
or U9389 (N_9389,N_838,N_2712);
nand U9390 (N_9390,N_2403,N_1427);
and U9391 (N_9391,N_1774,N_2931);
nor U9392 (N_9392,N_2832,N_4906);
and U9393 (N_9393,N_936,N_3309);
nand U9394 (N_9394,N_4891,N_3739);
nor U9395 (N_9395,N_4553,N_2189);
xor U9396 (N_9396,N_1498,N_171);
nand U9397 (N_9397,N_3704,N_2497);
nand U9398 (N_9398,N_249,N_3969);
nor U9399 (N_9399,N_3036,N_678);
and U9400 (N_9400,N_1172,N_2903);
nor U9401 (N_9401,N_3686,N_3572);
nor U9402 (N_9402,N_4962,N_603);
nand U9403 (N_9403,N_1337,N_2331);
and U9404 (N_9404,N_1800,N_3550);
and U9405 (N_9405,N_2418,N_4304);
nor U9406 (N_9406,N_164,N_304);
or U9407 (N_9407,N_3647,N_2148);
and U9408 (N_9408,N_1471,N_3339);
or U9409 (N_9409,N_3799,N_367);
and U9410 (N_9410,N_2895,N_666);
nand U9411 (N_9411,N_3647,N_988);
and U9412 (N_9412,N_3409,N_4478);
and U9413 (N_9413,N_3544,N_609);
nand U9414 (N_9414,N_2261,N_1749);
and U9415 (N_9415,N_2424,N_1712);
nor U9416 (N_9416,N_4756,N_298);
and U9417 (N_9417,N_379,N_3544);
or U9418 (N_9418,N_2731,N_368);
nor U9419 (N_9419,N_4125,N_386);
or U9420 (N_9420,N_3760,N_3086);
nor U9421 (N_9421,N_2086,N_3393);
and U9422 (N_9422,N_4682,N_4321);
or U9423 (N_9423,N_1203,N_2299);
nor U9424 (N_9424,N_4689,N_3471);
or U9425 (N_9425,N_2774,N_1807);
nor U9426 (N_9426,N_1526,N_4308);
or U9427 (N_9427,N_1442,N_1086);
nand U9428 (N_9428,N_612,N_4869);
and U9429 (N_9429,N_2876,N_4721);
nor U9430 (N_9430,N_136,N_279);
and U9431 (N_9431,N_473,N_3830);
nand U9432 (N_9432,N_2705,N_3008);
nor U9433 (N_9433,N_4415,N_3153);
or U9434 (N_9434,N_2553,N_2179);
nand U9435 (N_9435,N_569,N_19);
or U9436 (N_9436,N_542,N_3934);
and U9437 (N_9437,N_702,N_2245);
nand U9438 (N_9438,N_2133,N_2722);
or U9439 (N_9439,N_2733,N_4106);
xnor U9440 (N_9440,N_2767,N_1194);
nor U9441 (N_9441,N_1636,N_2112);
and U9442 (N_9442,N_716,N_4725);
nor U9443 (N_9443,N_427,N_3771);
nand U9444 (N_9444,N_4822,N_4106);
nor U9445 (N_9445,N_880,N_2868);
nor U9446 (N_9446,N_1558,N_788);
or U9447 (N_9447,N_618,N_4260);
and U9448 (N_9448,N_2713,N_3948);
nand U9449 (N_9449,N_3831,N_2623);
nor U9450 (N_9450,N_2255,N_2069);
xor U9451 (N_9451,N_4382,N_1342);
or U9452 (N_9452,N_538,N_2975);
xnor U9453 (N_9453,N_704,N_2085);
or U9454 (N_9454,N_299,N_3303);
nand U9455 (N_9455,N_106,N_4450);
nand U9456 (N_9456,N_1883,N_3872);
nand U9457 (N_9457,N_3623,N_2010);
nor U9458 (N_9458,N_4650,N_4822);
xnor U9459 (N_9459,N_875,N_1203);
nor U9460 (N_9460,N_2140,N_1097);
nor U9461 (N_9461,N_1300,N_3602);
and U9462 (N_9462,N_1122,N_2091);
nor U9463 (N_9463,N_4044,N_4007);
or U9464 (N_9464,N_207,N_699);
nor U9465 (N_9465,N_441,N_239);
xnor U9466 (N_9466,N_522,N_206);
nand U9467 (N_9467,N_1992,N_1701);
nand U9468 (N_9468,N_1582,N_2595);
nor U9469 (N_9469,N_2190,N_268);
nand U9470 (N_9470,N_4194,N_4292);
and U9471 (N_9471,N_375,N_3174);
nor U9472 (N_9472,N_209,N_1895);
and U9473 (N_9473,N_1400,N_4988);
nor U9474 (N_9474,N_847,N_3106);
and U9475 (N_9475,N_2502,N_3882);
and U9476 (N_9476,N_333,N_682);
or U9477 (N_9477,N_2766,N_78);
nand U9478 (N_9478,N_4720,N_4670);
nand U9479 (N_9479,N_3313,N_3121);
and U9480 (N_9480,N_660,N_1124);
or U9481 (N_9481,N_1400,N_3101);
nand U9482 (N_9482,N_748,N_1917);
nand U9483 (N_9483,N_914,N_1528);
and U9484 (N_9484,N_3016,N_873);
nor U9485 (N_9485,N_4121,N_4515);
nor U9486 (N_9486,N_502,N_4443);
or U9487 (N_9487,N_2340,N_3147);
nand U9488 (N_9488,N_4673,N_1559);
or U9489 (N_9489,N_4737,N_2623);
nand U9490 (N_9490,N_364,N_1333);
nand U9491 (N_9491,N_3887,N_2248);
and U9492 (N_9492,N_4956,N_2801);
nor U9493 (N_9493,N_3912,N_4454);
nor U9494 (N_9494,N_982,N_3793);
nor U9495 (N_9495,N_327,N_1613);
or U9496 (N_9496,N_3985,N_4967);
or U9497 (N_9497,N_689,N_4880);
nor U9498 (N_9498,N_4797,N_1964);
nor U9499 (N_9499,N_1956,N_2829);
nor U9500 (N_9500,N_457,N_4798);
or U9501 (N_9501,N_4626,N_1931);
xor U9502 (N_9502,N_4634,N_1463);
nand U9503 (N_9503,N_2165,N_2753);
nor U9504 (N_9504,N_2065,N_4786);
nand U9505 (N_9505,N_3798,N_246);
and U9506 (N_9506,N_3350,N_2926);
or U9507 (N_9507,N_122,N_2717);
or U9508 (N_9508,N_3093,N_3921);
or U9509 (N_9509,N_4484,N_3308);
nor U9510 (N_9510,N_2274,N_2314);
nor U9511 (N_9511,N_399,N_3622);
nor U9512 (N_9512,N_4619,N_2834);
or U9513 (N_9513,N_562,N_1819);
and U9514 (N_9514,N_2174,N_2099);
and U9515 (N_9515,N_3820,N_1190);
and U9516 (N_9516,N_3977,N_1109);
and U9517 (N_9517,N_4731,N_116);
or U9518 (N_9518,N_404,N_2679);
nor U9519 (N_9519,N_1615,N_3824);
nand U9520 (N_9520,N_4788,N_4688);
or U9521 (N_9521,N_2655,N_1973);
nand U9522 (N_9522,N_2386,N_1047);
nor U9523 (N_9523,N_4968,N_3308);
nor U9524 (N_9524,N_277,N_441);
and U9525 (N_9525,N_2167,N_119);
and U9526 (N_9526,N_3833,N_203);
and U9527 (N_9527,N_588,N_2360);
or U9528 (N_9528,N_3844,N_2878);
or U9529 (N_9529,N_4059,N_2525);
and U9530 (N_9530,N_600,N_886);
or U9531 (N_9531,N_2380,N_1381);
nand U9532 (N_9532,N_1837,N_1909);
nand U9533 (N_9533,N_541,N_2667);
or U9534 (N_9534,N_40,N_4745);
or U9535 (N_9535,N_3343,N_4929);
nand U9536 (N_9536,N_2396,N_2042);
or U9537 (N_9537,N_3702,N_2621);
or U9538 (N_9538,N_3092,N_2339);
or U9539 (N_9539,N_767,N_2671);
or U9540 (N_9540,N_3740,N_1337);
nor U9541 (N_9541,N_3046,N_3252);
nand U9542 (N_9542,N_3572,N_3621);
and U9543 (N_9543,N_4855,N_2422);
or U9544 (N_9544,N_3499,N_4717);
or U9545 (N_9545,N_1945,N_2994);
nor U9546 (N_9546,N_670,N_2381);
nand U9547 (N_9547,N_1692,N_4189);
nand U9548 (N_9548,N_4172,N_2426);
and U9549 (N_9549,N_2051,N_1214);
or U9550 (N_9550,N_3710,N_1638);
or U9551 (N_9551,N_1998,N_1646);
nor U9552 (N_9552,N_2081,N_339);
and U9553 (N_9553,N_4492,N_2176);
and U9554 (N_9554,N_2532,N_1257);
and U9555 (N_9555,N_2013,N_1110);
nor U9556 (N_9556,N_2826,N_1817);
and U9557 (N_9557,N_3396,N_3158);
xnor U9558 (N_9558,N_709,N_3875);
nand U9559 (N_9559,N_3801,N_1385);
and U9560 (N_9560,N_1360,N_813);
and U9561 (N_9561,N_3376,N_1890);
nor U9562 (N_9562,N_489,N_285);
nor U9563 (N_9563,N_624,N_4804);
and U9564 (N_9564,N_1569,N_2300);
or U9565 (N_9565,N_1411,N_2886);
or U9566 (N_9566,N_2469,N_214);
nor U9567 (N_9567,N_2277,N_1939);
or U9568 (N_9568,N_2266,N_4136);
and U9569 (N_9569,N_1791,N_1006);
and U9570 (N_9570,N_1724,N_3465);
nor U9571 (N_9571,N_3511,N_2644);
nor U9572 (N_9572,N_4658,N_4564);
or U9573 (N_9573,N_3726,N_3919);
nor U9574 (N_9574,N_3388,N_2466);
and U9575 (N_9575,N_1051,N_3007);
or U9576 (N_9576,N_4386,N_1490);
and U9577 (N_9577,N_1513,N_4783);
nor U9578 (N_9578,N_2351,N_3169);
nand U9579 (N_9579,N_285,N_1179);
and U9580 (N_9580,N_3100,N_4270);
or U9581 (N_9581,N_3553,N_2891);
nand U9582 (N_9582,N_2897,N_3489);
xor U9583 (N_9583,N_469,N_2448);
and U9584 (N_9584,N_331,N_2571);
nor U9585 (N_9585,N_4117,N_1916);
nand U9586 (N_9586,N_4773,N_2707);
or U9587 (N_9587,N_4700,N_4286);
or U9588 (N_9588,N_2926,N_3787);
or U9589 (N_9589,N_427,N_2624);
xor U9590 (N_9590,N_2449,N_1784);
or U9591 (N_9591,N_3316,N_1151);
nand U9592 (N_9592,N_2084,N_3592);
and U9593 (N_9593,N_1301,N_1190);
or U9594 (N_9594,N_4477,N_2928);
nor U9595 (N_9595,N_3587,N_3444);
and U9596 (N_9596,N_741,N_2485);
nand U9597 (N_9597,N_883,N_3886);
and U9598 (N_9598,N_2271,N_1999);
nand U9599 (N_9599,N_1608,N_3886);
and U9600 (N_9600,N_635,N_749);
nand U9601 (N_9601,N_1829,N_4296);
nor U9602 (N_9602,N_1100,N_3918);
and U9603 (N_9603,N_1092,N_3776);
or U9604 (N_9604,N_536,N_3439);
or U9605 (N_9605,N_508,N_4312);
and U9606 (N_9606,N_64,N_3456);
xor U9607 (N_9607,N_251,N_1932);
and U9608 (N_9608,N_800,N_4757);
and U9609 (N_9609,N_3318,N_3435);
nand U9610 (N_9610,N_1283,N_1619);
nor U9611 (N_9611,N_3492,N_3488);
or U9612 (N_9612,N_2774,N_1691);
and U9613 (N_9613,N_804,N_2761);
nand U9614 (N_9614,N_1849,N_1265);
or U9615 (N_9615,N_4763,N_2881);
nand U9616 (N_9616,N_1758,N_906);
and U9617 (N_9617,N_2751,N_2794);
nor U9618 (N_9618,N_879,N_346);
nor U9619 (N_9619,N_3355,N_2448);
or U9620 (N_9620,N_2103,N_3949);
and U9621 (N_9621,N_4423,N_3941);
or U9622 (N_9622,N_460,N_2157);
nand U9623 (N_9623,N_2618,N_2050);
nor U9624 (N_9624,N_1634,N_4175);
and U9625 (N_9625,N_3549,N_1750);
and U9626 (N_9626,N_2691,N_4150);
nand U9627 (N_9627,N_2753,N_2177);
or U9628 (N_9628,N_2790,N_4549);
or U9629 (N_9629,N_512,N_1871);
nand U9630 (N_9630,N_4013,N_4524);
nor U9631 (N_9631,N_2281,N_2796);
nand U9632 (N_9632,N_3179,N_152);
nand U9633 (N_9633,N_2563,N_1445);
nor U9634 (N_9634,N_4656,N_1189);
and U9635 (N_9635,N_4326,N_1663);
or U9636 (N_9636,N_3321,N_2594);
or U9637 (N_9637,N_1075,N_1307);
and U9638 (N_9638,N_673,N_1646);
xnor U9639 (N_9639,N_2720,N_3554);
nor U9640 (N_9640,N_4750,N_4769);
nor U9641 (N_9641,N_2492,N_3538);
or U9642 (N_9642,N_4349,N_375);
nor U9643 (N_9643,N_4122,N_334);
and U9644 (N_9644,N_905,N_3148);
nor U9645 (N_9645,N_1102,N_1974);
nand U9646 (N_9646,N_2627,N_1585);
nor U9647 (N_9647,N_2403,N_4005);
or U9648 (N_9648,N_2607,N_4411);
nand U9649 (N_9649,N_1558,N_3481);
and U9650 (N_9650,N_2784,N_2837);
nor U9651 (N_9651,N_3872,N_4641);
nand U9652 (N_9652,N_3326,N_3670);
xnor U9653 (N_9653,N_1430,N_4192);
and U9654 (N_9654,N_696,N_4327);
or U9655 (N_9655,N_3831,N_2068);
nand U9656 (N_9656,N_2141,N_1958);
or U9657 (N_9657,N_275,N_1672);
nand U9658 (N_9658,N_3625,N_1477);
nor U9659 (N_9659,N_3334,N_1391);
xor U9660 (N_9660,N_1621,N_463);
nand U9661 (N_9661,N_3887,N_3729);
and U9662 (N_9662,N_3185,N_2104);
or U9663 (N_9663,N_575,N_3841);
nor U9664 (N_9664,N_4881,N_59);
nand U9665 (N_9665,N_2530,N_3212);
nand U9666 (N_9666,N_3439,N_2043);
or U9667 (N_9667,N_3792,N_3168);
nor U9668 (N_9668,N_4864,N_755);
nor U9669 (N_9669,N_330,N_1594);
and U9670 (N_9670,N_4274,N_1988);
nor U9671 (N_9671,N_1449,N_2577);
and U9672 (N_9672,N_4129,N_3423);
or U9673 (N_9673,N_2907,N_2421);
nand U9674 (N_9674,N_2514,N_2492);
nor U9675 (N_9675,N_2706,N_746);
nor U9676 (N_9676,N_2648,N_1174);
nand U9677 (N_9677,N_1636,N_2970);
nor U9678 (N_9678,N_1636,N_4822);
and U9679 (N_9679,N_1173,N_4039);
nand U9680 (N_9680,N_2225,N_1071);
and U9681 (N_9681,N_814,N_4081);
nor U9682 (N_9682,N_3951,N_3256);
nand U9683 (N_9683,N_3440,N_4200);
xnor U9684 (N_9684,N_3192,N_1397);
nand U9685 (N_9685,N_1691,N_3843);
and U9686 (N_9686,N_1945,N_1925);
nor U9687 (N_9687,N_3152,N_4005);
nand U9688 (N_9688,N_1863,N_4896);
and U9689 (N_9689,N_3583,N_4790);
or U9690 (N_9690,N_4872,N_1201);
or U9691 (N_9691,N_3523,N_4754);
and U9692 (N_9692,N_3313,N_2455);
nand U9693 (N_9693,N_2952,N_4605);
or U9694 (N_9694,N_4224,N_669);
nor U9695 (N_9695,N_21,N_3117);
or U9696 (N_9696,N_1106,N_2193);
or U9697 (N_9697,N_1353,N_3957);
nand U9698 (N_9698,N_3021,N_2388);
nor U9699 (N_9699,N_3149,N_1762);
nor U9700 (N_9700,N_2224,N_2201);
xnor U9701 (N_9701,N_361,N_2430);
or U9702 (N_9702,N_564,N_4811);
and U9703 (N_9703,N_4469,N_3570);
and U9704 (N_9704,N_3951,N_4835);
or U9705 (N_9705,N_2763,N_4941);
and U9706 (N_9706,N_3386,N_4198);
and U9707 (N_9707,N_2153,N_4592);
nor U9708 (N_9708,N_493,N_481);
and U9709 (N_9709,N_1662,N_3115);
or U9710 (N_9710,N_4801,N_2566);
or U9711 (N_9711,N_1194,N_1300);
and U9712 (N_9712,N_3960,N_607);
nand U9713 (N_9713,N_3762,N_3281);
or U9714 (N_9714,N_1904,N_2958);
nor U9715 (N_9715,N_3567,N_3993);
nand U9716 (N_9716,N_2393,N_3266);
and U9717 (N_9717,N_4046,N_1198);
xnor U9718 (N_9718,N_1550,N_4439);
xor U9719 (N_9719,N_715,N_1317);
nor U9720 (N_9720,N_2804,N_4049);
nor U9721 (N_9721,N_3758,N_270);
and U9722 (N_9722,N_3434,N_1002);
and U9723 (N_9723,N_964,N_1471);
nor U9724 (N_9724,N_3453,N_3520);
nand U9725 (N_9725,N_4488,N_2833);
nor U9726 (N_9726,N_2005,N_2354);
and U9727 (N_9727,N_3275,N_1604);
and U9728 (N_9728,N_1002,N_4108);
nand U9729 (N_9729,N_3551,N_2098);
nand U9730 (N_9730,N_2737,N_1925);
nand U9731 (N_9731,N_4524,N_702);
or U9732 (N_9732,N_591,N_3244);
nand U9733 (N_9733,N_1743,N_553);
nand U9734 (N_9734,N_1062,N_2335);
or U9735 (N_9735,N_3107,N_2388);
and U9736 (N_9736,N_1470,N_3894);
nand U9737 (N_9737,N_536,N_1411);
nand U9738 (N_9738,N_4153,N_25);
xnor U9739 (N_9739,N_196,N_1867);
or U9740 (N_9740,N_3175,N_3627);
or U9741 (N_9741,N_4042,N_942);
and U9742 (N_9742,N_1032,N_3164);
or U9743 (N_9743,N_3156,N_1375);
xor U9744 (N_9744,N_1328,N_193);
and U9745 (N_9745,N_1985,N_672);
and U9746 (N_9746,N_652,N_4809);
or U9747 (N_9747,N_1585,N_1555);
nor U9748 (N_9748,N_2107,N_1618);
nor U9749 (N_9749,N_4164,N_3657);
nor U9750 (N_9750,N_3936,N_2568);
and U9751 (N_9751,N_3173,N_164);
and U9752 (N_9752,N_470,N_4668);
and U9753 (N_9753,N_2993,N_2777);
or U9754 (N_9754,N_1777,N_3932);
nor U9755 (N_9755,N_398,N_2587);
and U9756 (N_9756,N_1160,N_1534);
or U9757 (N_9757,N_47,N_3737);
nor U9758 (N_9758,N_1102,N_4407);
and U9759 (N_9759,N_3875,N_170);
or U9760 (N_9760,N_1956,N_4653);
and U9761 (N_9761,N_297,N_3643);
and U9762 (N_9762,N_3405,N_2148);
nand U9763 (N_9763,N_1683,N_3107);
nor U9764 (N_9764,N_4660,N_1309);
nand U9765 (N_9765,N_3112,N_1983);
nor U9766 (N_9766,N_1318,N_3842);
nor U9767 (N_9767,N_4024,N_1949);
nor U9768 (N_9768,N_1968,N_2788);
and U9769 (N_9769,N_275,N_1262);
nor U9770 (N_9770,N_4551,N_456);
nor U9771 (N_9771,N_3755,N_3270);
and U9772 (N_9772,N_3925,N_2944);
nand U9773 (N_9773,N_525,N_215);
nand U9774 (N_9774,N_3557,N_3923);
nand U9775 (N_9775,N_3293,N_825);
nor U9776 (N_9776,N_2014,N_2200);
or U9777 (N_9777,N_4499,N_3572);
or U9778 (N_9778,N_427,N_4678);
and U9779 (N_9779,N_516,N_4696);
and U9780 (N_9780,N_194,N_4122);
nand U9781 (N_9781,N_2565,N_3712);
nor U9782 (N_9782,N_3086,N_2716);
nor U9783 (N_9783,N_3761,N_2532);
or U9784 (N_9784,N_2652,N_4857);
nand U9785 (N_9785,N_3617,N_4356);
nor U9786 (N_9786,N_288,N_2122);
nand U9787 (N_9787,N_18,N_2703);
nor U9788 (N_9788,N_3117,N_2947);
or U9789 (N_9789,N_3298,N_2369);
and U9790 (N_9790,N_4134,N_3263);
or U9791 (N_9791,N_2709,N_3042);
nor U9792 (N_9792,N_549,N_1687);
nand U9793 (N_9793,N_3814,N_3743);
and U9794 (N_9794,N_3099,N_2850);
nand U9795 (N_9795,N_2149,N_993);
and U9796 (N_9796,N_912,N_4247);
nor U9797 (N_9797,N_83,N_4729);
nor U9798 (N_9798,N_2922,N_3278);
xnor U9799 (N_9799,N_818,N_1646);
nand U9800 (N_9800,N_2410,N_208);
or U9801 (N_9801,N_1352,N_1760);
nand U9802 (N_9802,N_3339,N_2533);
and U9803 (N_9803,N_38,N_1463);
nor U9804 (N_9804,N_2623,N_425);
nor U9805 (N_9805,N_4173,N_1911);
nand U9806 (N_9806,N_4062,N_1395);
nand U9807 (N_9807,N_2377,N_1);
or U9808 (N_9808,N_161,N_2717);
nand U9809 (N_9809,N_1794,N_4821);
nand U9810 (N_9810,N_1491,N_1706);
nor U9811 (N_9811,N_3386,N_437);
nand U9812 (N_9812,N_3692,N_1644);
nor U9813 (N_9813,N_3447,N_618);
and U9814 (N_9814,N_3650,N_1496);
nor U9815 (N_9815,N_2259,N_1275);
xor U9816 (N_9816,N_1074,N_4270);
xor U9817 (N_9817,N_4755,N_366);
or U9818 (N_9818,N_60,N_1396);
and U9819 (N_9819,N_1356,N_3670);
and U9820 (N_9820,N_2015,N_2179);
or U9821 (N_9821,N_4058,N_414);
nand U9822 (N_9822,N_2546,N_3523);
nor U9823 (N_9823,N_3208,N_4940);
nor U9824 (N_9824,N_2224,N_2461);
or U9825 (N_9825,N_1184,N_3392);
or U9826 (N_9826,N_1416,N_2385);
nor U9827 (N_9827,N_4839,N_4949);
nand U9828 (N_9828,N_4994,N_2262);
nand U9829 (N_9829,N_2510,N_878);
and U9830 (N_9830,N_4083,N_2848);
and U9831 (N_9831,N_2411,N_2285);
nand U9832 (N_9832,N_1506,N_3497);
and U9833 (N_9833,N_4667,N_2984);
or U9834 (N_9834,N_3638,N_3597);
or U9835 (N_9835,N_889,N_263);
nand U9836 (N_9836,N_2563,N_4956);
nand U9837 (N_9837,N_1641,N_3939);
or U9838 (N_9838,N_4734,N_2076);
and U9839 (N_9839,N_3928,N_1798);
or U9840 (N_9840,N_1209,N_1831);
nor U9841 (N_9841,N_571,N_2928);
nor U9842 (N_9842,N_1109,N_3353);
nor U9843 (N_9843,N_2492,N_242);
and U9844 (N_9844,N_1205,N_3600);
or U9845 (N_9845,N_3844,N_2698);
nand U9846 (N_9846,N_3312,N_3027);
or U9847 (N_9847,N_1369,N_1141);
nor U9848 (N_9848,N_453,N_2498);
xor U9849 (N_9849,N_4836,N_2885);
xnor U9850 (N_9850,N_1791,N_1414);
nor U9851 (N_9851,N_1948,N_2414);
or U9852 (N_9852,N_3341,N_3792);
and U9853 (N_9853,N_3848,N_4601);
nand U9854 (N_9854,N_1216,N_832);
or U9855 (N_9855,N_1933,N_1071);
nor U9856 (N_9856,N_3306,N_2664);
or U9857 (N_9857,N_1252,N_2887);
nand U9858 (N_9858,N_1629,N_2765);
and U9859 (N_9859,N_2861,N_2532);
nor U9860 (N_9860,N_4149,N_1306);
nand U9861 (N_9861,N_8,N_1454);
and U9862 (N_9862,N_4843,N_3402);
and U9863 (N_9863,N_1379,N_1644);
nor U9864 (N_9864,N_128,N_1626);
or U9865 (N_9865,N_3140,N_2108);
and U9866 (N_9866,N_3864,N_1210);
nand U9867 (N_9867,N_1616,N_4869);
nor U9868 (N_9868,N_799,N_3905);
and U9869 (N_9869,N_3324,N_2993);
and U9870 (N_9870,N_3605,N_3736);
or U9871 (N_9871,N_2903,N_3816);
nand U9872 (N_9872,N_4184,N_4202);
and U9873 (N_9873,N_1896,N_2691);
nor U9874 (N_9874,N_2928,N_4921);
nand U9875 (N_9875,N_96,N_2849);
nor U9876 (N_9876,N_1387,N_1428);
and U9877 (N_9877,N_1999,N_1574);
nand U9878 (N_9878,N_3380,N_2836);
nand U9879 (N_9879,N_3788,N_1002);
and U9880 (N_9880,N_1639,N_2655);
nand U9881 (N_9881,N_3487,N_4786);
nor U9882 (N_9882,N_4357,N_2163);
nor U9883 (N_9883,N_760,N_2241);
nand U9884 (N_9884,N_3742,N_2965);
and U9885 (N_9885,N_1891,N_3396);
nand U9886 (N_9886,N_305,N_4831);
nor U9887 (N_9887,N_2683,N_131);
nand U9888 (N_9888,N_1169,N_4532);
and U9889 (N_9889,N_2581,N_1623);
or U9890 (N_9890,N_3284,N_1615);
nor U9891 (N_9891,N_3495,N_1614);
or U9892 (N_9892,N_946,N_2605);
or U9893 (N_9893,N_2354,N_3648);
or U9894 (N_9894,N_635,N_450);
nand U9895 (N_9895,N_4033,N_1273);
nor U9896 (N_9896,N_4495,N_1327);
and U9897 (N_9897,N_1901,N_2174);
xnor U9898 (N_9898,N_1067,N_1373);
nand U9899 (N_9899,N_3566,N_3488);
nor U9900 (N_9900,N_196,N_1075);
nand U9901 (N_9901,N_4607,N_4433);
nand U9902 (N_9902,N_3940,N_2184);
xor U9903 (N_9903,N_375,N_4448);
nor U9904 (N_9904,N_2130,N_1960);
nand U9905 (N_9905,N_4704,N_2839);
nor U9906 (N_9906,N_180,N_4436);
nor U9907 (N_9907,N_1794,N_2095);
and U9908 (N_9908,N_4286,N_3341);
nand U9909 (N_9909,N_1622,N_2618);
xor U9910 (N_9910,N_673,N_3850);
nor U9911 (N_9911,N_4785,N_3768);
and U9912 (N_9912,N_4284,N_2304);
nor U9913 (N_9913,N_2472,N_442);
or U9914 (N_9914,N_2807,N_1268);
or U9915 (N_9915,N_3861,N_54);
or U9916 (N_9916,N_1537,N_723);
or U9917 (N_9917,N_1482,N_4007);
or U9918 (N_9918,N_1055,N_190);
and U9919 (N_9919,N_4268,N_258);
xnor U9920 (N_9920,N_1191,N_2508);
nor U9921 (N_9921,N_4160,N_1219);
nand U9922 (N_9922,N_4150,N_1614);
nand U9923 (N_9923,N_2557,N_878);
nor U9924 (N_9924,N_2572,N_2036);
or U9925 (N_9925,N_2268,N_1074);
nand U9926 (N_9926,N_2242,N_4846);
or U9927 (N_9927,N_399,N_2327);
or U9928 (N_9928,N_1918,N_3440);
nand U9929 (N_9929,N_3562,N_1462);
nand U9930 (N_9930,N_3869,N_4690);
nor U9931 (N_9931,N_14,N_711);
nor U9932 (N_9932,N_4527,N_2447);
nor U9933 (N_9933,N_3275,N_3088);
or U9934 (N_9934,N_2545,N_3168);
and U9935 (N_9935,N_100,N_536);
nor U9936 (N_9936,N_4652,N_3219);
nor U9937 (N_9937,N_2740,N_2765);
nand U9938 (N_9938,N_2628,N_3316);
or U9939 (N_9939,N_2466,N_313);
nor U9940 (N_9940,N_3628,N_4450);
and U9941 (N_9941,N_1541,N_3471);
xor U9942 (N_9942,N_2588,N_2626);
nand U9943 (N_9943,N_376,N_2160);
nor U9944 (N_9944,N_2600,N_793);
xor U9945 (N_9945,N_1085,N_2973);
and U9946 (N_9946,N_4443,N_3162);
nor U9947 (N_9947,N_1052,N_1826);
nand U9948 (N_9948,N_148,N_2510);
nand U9949 (N_9949,N_2133,N_338);
and U9950 (N_9950,N_3822,N_2369);
and U9951 (N_9951,N_3969,N_2712);
nor U9952 (N_9952,N_4698,N_1939);
nor U9953 (N_9953,N_3313,N_1236);
nor U9954 (N_9954,N_2210,N_2702);
or U9955 (N_9955,N_157,N_822);
nor U9956 (N_9956,N_2984,N_3053);
and U9957 (N_9957,N_2303,N_3230);
and U9958 (N_9958,N_4385,N_2348);
nor U9959 (N_9959,N_2102,N_1833);
or U9960 (N_9960,N_1837,N_1612);
nand U9961 (N_9961,N_1427,N_1603);
nor U9962 (N_9962,N_2043,N_4671);
nor U9963 (N_9963,N_2835,N_3921);
nand U9964 (N_9964,N_2187,N_2939);
and U9965 (N_9965,N_1644,N_3090);
and U9966 (N_9966,N_3937,N_1486);
and U9967 (N_9967,N_4503,N_3589);
and U9968 (N_9968,N_790,N_810);
nor U9969 (N_9969,N_2013,N_3756);
or U9970 (N_9970,N_2727,N_1858);
nand U9971 (N_9971,N_4110,N_4364);
nand U9972 (N_9972,N_612,N_4405);
nand U9973 (N_9973,N_1419,N_1554);
nand U9974 (N_9974,N_2,N_4707);
nand U9975 (N_9975,N_4778,N_1134);
xor U9976 (N_9976,N_927,N_3929);
nand U9977 (N_9977,N_3344,N_172);
nand U9978 (N_9978,N_2618,N_1820);
nor U9979 (N_9979,N_3953,N_4366);
and U9980 (N_9980,N_468,N_2604);
nor U9981 (N_9981,N_1130,N_3361);
nor U9982 (N_9982,N_972,N_2057);
or U9983 (N_9983,N_4928,N_2445);
nand U9984 (N_9984,N_3082,N_890);
nand U9985 (N_9985,N_3403,N_207);
or U9986 (N_9986,N_3825,N_2560);
nand U9987 (N_9987,N_1870,N_2592);
and U9988 (N_9988,N_259,N_3813);
nor U9989 (N_9989,N_157,N_3457);
nor U9990 (N_9990,N_2972,N_2109);
nor U9991 (N_9991,N_586,N_3961);
and U9992 (N_9992,N_2765,N_2253);
and U9993 (N_9993,N_1681,N_419);
or U9994 (N_9994,N_2503,N_4571);
or U9995 (N_9995,N_747,N_4740);
or U9996 (N_9996,N_1110,N_2896);
and U9997 (N_9997,N_341,N_2397);
or U9998 (N_9998,N_3937,N_4044);
nor U9999 (N_9999,N_2882,N_3321);
and UO_0 (O_0,N_9231,N_9373);
nor UO_1 (O_1,N_9939,N_8308);
or UO_2 (O_2,N_9256,N_7226);
and UO_3 (O_3,N_7016,N_5998);
nor UO_4 (O_4,N_7642,N_8020);
or UO_5 (O_5,N_7585,N_5050);
or UO_6 (O_6,N_9055,N_8772);
nand UO_7 (O_7,N_5649,N_6959);
nand UO_8 (O_8,N_6837,N_5526);
nor UO_9 (O_9,N_6089,N_9983);
and UO_10 (O_10,N_7336,N_9765);
or UO_11 (O_11,N_6630,N_7105);
nor UO_12 (O_12,N_6543,N_6413);
nor UO_13 (O_13,N_8849,N_8545);
nand UO_14 (O_14,N_7350,N_6319);
and UO_15 (O_15,N_8294,N_7302);
nor UO_16 (O_16,N_9652,N_5747);
nor UO_17 (O_17,N_5524,N_8941);
or UO_18 (O_18,N_9051,N_9556);
nand UO_19 (O_19,N_6161,N_9724);
nor UO_20 (O_20,N_5118,N_6871);
nor UO_21 (O_21,N_9213,N_5140);
and UO_22 (O_22,N_5664,N_5764);
nand UO_23 (O_23,N_9968,N_5654);
nand UO_24 (O_24,N_8588,N_7317);
or UO_25 (O_25,N_5684,N_5963);
nor UO_26 (O_26,N_7323,N_5312);
nand UO_27 (O_27,N_9833,N_7912);
nand UO_28 (O_28,N_9109,N_9875);
nor UO_29 (O_29,N_7612,N_8669);
nor UO_30 (O_30,N_8266,N_7294);
nand UO_31 (O_31,N_5117,N_5148);
xor UO_32 (O_32,N_7499,N_8429);
nand UO_33 (O_33,N_7273,N_7271);
nand UO_34 (O_34,N_6520,N_6822);
nor UO_35 (O_35,N_7039,N_8218);
nand UO_36 (O_36,N_7730,N_7261);
or UO_37 (O_37,N_6027,N_6956);
nand UO_38 (O_38,N_6340,N_8979);
nand UO_39 (O_39,N_5081,N_5335);
nand UO_40 (O_40,N_9555,N_9104);
nand UO_41 (O_41,N_7353,N_9527);
nor UO_42 (O_42,N_7625,N_6439);
nor UO_43 (O_43,N_7218,N_8965);
or UO_44 (O_44,N_6577,N_7794);
nand UO_45 (O_45,N_7915,N_9560);
nor UO_46 (O_46,N_9732,N_8284);
nand UO_47 (O_47,N_9281,N_8847);
and UO_48 (O_48,N_9241,N_8831);
xor UO_49 (O_49,N_8393,N_7971);
nand UO_50 (O_50,N_7919,N_7784);
or UO_51 (O_51,N_8828,N_6278);
nor UO_52 (O_52,N_8301,N_7284);
nor UO_53 (O_53,N_7037,N_9850);
and UO_54 (O_54,N_8177,N_8161);
nand UO_55 (O_55,N_7724,N_6470);
or UO_56 (O_56,N_5460,N_5468);
and UO_57 (O_57,N_9338,N_9209);
nor UO_58 (O_58,N_7656,N_8634);
or UO_59 (O_59,N_8838,N_9353);
xor UO_60 (O_60,N_7621,N_6781);
or UO_61 (O_61,N_9477,N_5245);
nand UO_62 (O_62,N_8782,N_9060);
or UO_63 (O_63,N_7215,N_6805);
or UO_64 (O_64,N_8237,N_9788);
or UO_65 (O_65,N_9719,N_9369);
nand UO_66 (O_66,N_5137,N_8586);
nor UO_67 (O_67,N_9401,N_6549);
xor UO_68 (O_68,N_5262,N_9879);
nand UO_69 (O_69,N_9976,N_6111);
and UO_70 (O_70,N_5456,N_5177);
xor UO_71 (O_71,N_9517,N_7916);
nand UO_72 (O_72,N_6722,N_7254);
nor UO_73 (O_73,N_5969,N_8376);
nand UO_74 (O_74,N_6049,N_9249);
nand UO_75 (O_75,N_8431,N_7867);
nand UO_76 (O_76,N_9909,N_8857);
nand UO_77 (O_77,N_5017,N_7901);
and UO_78 (O_78,N_6726,N_5123);
nor UO_79 (O_79,N_6662,N_5188);
nand UO_80 (O_80,N_9965,N_5163);
and UO_81 (O_81,N_5186,N_5552);
and UO_82 (O_82,N_5330,N_8726);
or UO_83 (O_83,N_6804,N_5987);
nand UO_84 (O_84,N_8809,N_7958);
or UO_85 (O_85,N_6203,N_7520);
nor UO_86 (O_86,N_7663,N_9405);
nand UO_87 (O_87,N_8332,N_7004);
and UO_88 (O_88,N_7408,N_9197);
nor UO_89 (O_89,N_9799,N_9237);
and UO_90 (O_90,N_6332,N_7151);
nand UO_91 (O_91,N_6563,N_9920);
and UO_92 (O_92,N_5305,N_5247);
and UO_93 (O_93,N_9997,N_7208);
and UO_94 (O_94,N_9200,N_5746);
nor UO_95 (O_95,N_8678,N_8707);
nand UO_96 (O_96,N_9822,N_7754);
and UO_97 (O_97,N_8070,N_9364);
and UO_98 (O_98,N_6682,N_9870);
nor UO_99 (O_99,N_6204,N_5913);
nor UO_100 (O_100,N_7618,N_9166);
or UO_101 (O_101,N_9087,N_8221);
and UO_102 (O_102,N_5065,N_8607);
xnor UO_103 (O_103,N_9378,N_6013);
nand UO_104 (O_104,N_5478,N_7080);
nor UO_105 (O_105,N_7316,N_8955);
or UO_106 (O_106,N_8078,N_8880);
or UO_107 (O_107,N_8068,N_9271);
nand UO_108 (O_108,N_9689,N_8687);
or UO_109 (O_109,N_6583,N_5187);
and UO_110 (O_110,N_5702,N_7814);
nand UO_111 (O_111,N_5369,N_7326);
nand UO_112 (O_112,N_6339,N_9688);
nor UO_113 (O_113,N_6243,N_5791);
nand UO_114 (O_114,N_6383,N_8207);
or UO_115 (O_115,N_5498,N_8969);
and UO_116 (O_116,N_5910,N_8012);
nor UO_117 (O_117,N_7095,N_5202);
nor UO_118 (O_118,N_5584,N_5266);
nand UO_119 (O_119,N_7213,N_8216);
nor UO_120 (O_120,N_8881,N_8818);
or UO_121 (O_121,N_9809,N_6975);
nor UO_122 (O_122,N_6715,N_6219);
nand UO_123 (O_123,N_9932,N_6133);
and UO_124 (O_124,N_7592,N_9904);
nand UO_125 (O_125,N_9512,N_6988);
and UO_126 (O_126,N_5628,N_8668);
nor UO_127 (O_127,N_7232,N_8283);
nand UO_128 (O_128,N_5770,N_9942);
nand UO_129 (O_129,N_9462,N_7998);
or UO_130 (O_130,N_5024,N_5792);
and UO_131 (O_131,N_8093,N_6255);
nor UO_132 (O_132,N_7139,N_6224);
nor UO_133 (O_133,N_5834,N_9389);
or UO_134 (O_134,N_5308,N_7739);
nand UO_135 (O_135,N_9818,N_7085);
and UO_136 (O_136,N_9003,N_9402);
or UO_137 (O_137,N_8180,N_6460);
nand UO_138 (O_138,N_9215,N_9873);
or UO_139 (O_139,N_9878,N_8648);
nor UO_140 (O_140,N_9734,N_6028);
nand UO_141 (O_141,N_5596,N_9691);
nand UO_142 (O_142,N_6128,N_8758);
nand UO_143 (O_143,N_7205,N_7412);
nor UO_144 (O_144,N_5014,N_7118);
and UO_145 (O_145,N_9454,N_9861);
or UO_146 (O_146,N_8558,N_8866);
and UO_147 (O_147,N_8936,N_5813);
and UO_148 (O_148,N_7005,N_5842);
and UO_149 (O_149,N_6746,N_6116);
or UO_150 (O_150,N_6612,N_8533);
and UO_151 (O_151,N_9449,N_8132);
nor UO_152 (O_152,N_8122,N_5748);
and UO_153 (O_153,N_5599,N_5721);
or UO_154 (O_154,N_9727,N_9453);
nor UO_155 (O_155,N_8879,N_9886);
nor UO_156 (O_156,N_6588,N_8756);
nand UO_157 (O_157,N_9573,N_7508);
nand UO_158 (O_158,N_6575,N_9919);
and UO_159 (O_159,N_9735,N_8110);
nor UO_160 (O_160,N_8426,N_9272);
nor UO_161 (O_161,N_9242,N_6314);
or UO_162 (O_162,N_5920,N_5992);
nand UO_163 (O_163,N_7149,N_9802);
nand UO_164 (O_164,N_6463,N_8627);
nand UO_165 (O_165,N_8998,N_9250);
nor UO_166 (O_166,N_8839,N_7362);
or UO_167 (O_167,N_5655,N_8871);
nand UO_168 (O_168,N_8022,N_7458);
nand UO_169 (O_169,N_6345,N_5563);
or UO_170 (O_170,N_9295,N_5627);
and UO_171 (O_171,N_6570,N_8532);
nor UO_172 (O_172,N_9036,N_8834);
or UO_173 (O_173,N_6674,N_7021);
and UO_174 (O_174,N_9622,N_8561);
and UO_175 (O_175,N_9923,N_7077);
nand UO_176 (O_176,N_9082,N_9996);
or UO_177 (O_177,N_7835,N_5625);
xor UO_178 (O_178,N_6743,N_6574);
nand UO_179 (O_179,N_5000,N_5958);
and UO_180 (O_180,N_7830,N_9595);
and UO_181 (O_181,N_5417,N_7069);
or UO_182 (O_182,N_7780,N_6555);
nor UO_183 (O_183,N_7983,N_8727);
nand UO_184 (O_184,N_9224,N_5688);
or UO_185 (O_185,N_6468,N_7356);
or UO_186 (O_186,N_5488,N_5737);
xnor UO_187 (O_187,N_5586,N_9451);
nand UO_188 (O_188,N_6497,N_7877);
nor UO_189 (O_189,N_6703,N_9865);
nor UO_190 (O_190,N_8716,N_5282);
or UO_191 (O_191,N_9607,N_8396);
nor UO_192 (O_192,N_5815,N_5494);
and UO_193 (O_193,N_8762,N_9973);
and UO_194 (O_194,N_9383,N_6026);
nand UO_195 (O_195,N_9914,N_5577);
nor UO_196 (O_196,N_6714,N_8193);
nor UO_197 (O_197,N_5470,N_8292);
or UO_198 (O_198,N_6756,N_7553);
nor UO_199 (O_199,N_7052,N_6229);
nand UO_200 (O_200,N_5896,N_6928);
nand UO_201 (O_201,N_5058,N_9304);
or UO_202 (O_202,N_9698,N_6731);
or UO_203 (O_203,N_9274,N_5428);
or UO_204 (O_204,N_7078,N_6474);
and UO_205 (O_205,N_5108,N_6631);
and UO_206 (O_206,N_6768,N_9946);
nor UO_207 (O_207,N_5917,N_7158);
and UO_208 (O_208,N_6915,N_9950);
or UO_209 (O_209,N_5124,N_6132);
xnor UO_210 (O_210,N_9053,N_8660);
nor UO_211 (O_211,N_9977,N_6177);
and UO_212 (O_212,N_6596,N_5585);
nand UO_213 (O_213,N_8751,N_5334);
nor UO_214 (O_214,N_5600,N_6399);
nor UO_215 (O_215,N_6274,N_9111);
nand UO_216 (O_216,N_8339,N_7764);
nor UO_217 (O_217,N_5267,N_8360);
nor UO_218 (O_218,N_9098,N_8453);
nand UO_219 (O_219,N_5855,N_7613);
and UO_220 (O_220,N_7711,N_7347);
nand UO_221 (O_221,N_9600,N_6223);
or UO_222 (O_222,N_6327,N_7898);
and UO_223 (O_223,N_8626,N_8615);
and UO_224 (O_224,N_9432,N_7293);
nand UO_225 (O_225,N_8058,N_5979);
or UO_226 (O_226,N_9511,N_7120);
and UO_227 (O_227,N_8992,N_7533);
or UO_228 (O_228,N_7861,N_6825);
and UO_229 (O_229,N_7060,N_5845);
nor UO_230 (O_230,N_5622,N_6665);
or UO_231 (O_231,N_7358,N_5873);
and UO_232 (O_232,N_6688,N_6600);
nand UO_233 (O_233,N_7991,N_9203);
or UO_234 (O_234,N_5218,N_8146);
or UO_235 (O_235,N_7582,N_6499);
and UO_236 (O_236,N_9929,N_5101);
nor UO_237 (O_237,N_9321,N_6702);
or UO_238 (O_238,N_5323,N_9754);
or UO_239 (O_239,N_7355,N_5029);
nand UO_240 (O_240,N_9993,N_7598);
and UO_241 (O_241,N_9160,N_8508);
and UO_242 (O_242,N_9971,N_9760);
nand UO_243 (O_243,N_7735,N_8116);
and UO_244 (O_244,N_9880,N_5038);
xnor UO_245 (O_245,N_6560,N_9037);
and UO_246 (O_246,N_9564,N_6761);
nor UO_247 (O_247,N_8739,N_8821);
nand UO_248 (O_248,N_5387,N_5571);
nor UO_249 (O_249,N_7561,N_8636);
nor UO_250 (O_250,N_6569,N_7806);
and UO_251 (O_251,N_5086,N_6732);
xor UO_252 (O_252,N_8421,N_7238);
or UO_253 (O_253,N_8597,N_9877);
and UO_254 (O_254,N_7067,N_8767);
or UO_255 (O_255,N_7511,N_8973);
and UO_256 (O_256,N_6788,N_8120);
nand UO_257 (O_257,N_7190,N_8224);
nor UO_258 (O_258,N_5598,N_8107);
nor UO_259 (O_259,N_8873,N_7962);
or UO_260 (O_260,N_7061,N_5793);
nand UO_261 (O_261,N_9108,N_5317);
and UO_262 (O_262,N_8441,N_9736);
nor UO_263 (O_263,N_5899,N_5447);
or UO_264 (O_264,N_5605,N_6415);
or UO_265 (O_265,N_7551,N_9062);
or UO_266 (O_266,N_5047,N_7485);
and UO_267 (O_267,N_5506,N_9761);
and UO_268 (O_268,N_5631,N_5185);
or UO_269 (O_269,N_5258,N_6890);
or UO_270 (O_270,N_9370,N_8060);
nor UO_271 (O_271,N_8511,N_6124);
or UO_272 (O_272,N_5427,N_7854);
nor UO_273 (O_273,N_9016,N_7658);
or UO_274 (O_274,N_5464,N_8963);
nor UO_275 (O_275,N_9110,N_5463);
nor UO_276 (O_276,N_7853,N_6624);
and UO_277 (O_277,N_5818,N_5274);
and UO_278 (O_278,N_6902,N_9657);
and UO_279 (O_279,N_8920,N_8034);
and UO_280 (O_280,N_5773,N_7790);
and UO_281 (O_281,N_6706,N_9012);
xnor UO_282 (O_282,N_9374,N_7429);
nand UO_283 (O_283,N_9248,N_5727);
nand UO_284 (O_284,N_7341,N_9386);
nand UO_285 (O_285,N_5357,N_8000);
nor UO_286 (O_286,N_5443,N_8001);
nand UO_287 (O_287,N_9516,N_6792);
nand UO_288 (O_288,N_9429,N_6344);
nand UO_289 (O_289,N_5619,N_9144);
nand UO_290 (O_290,N_5742,N_7907);
nand UO_291 (O_291,N_7282,N_6424);
and UO_292 (O_292,N_8323,N_7740);
or UO_293 (O_293,N_8559,N_8836);
or UO_294 (O_294,N_8620,N_7892);
nor UO_295 (O_295,N_8111,N_7479);
or UO_296 (O_296,N_9269,N_8824);
nand UO_297 (O_297,N_8208,N_7703);
nor UO_298 (O_298,N_9785,N_6842);
or UO_299 (O_299,N_8444,N_9356);
nor UO_300 (O_300,N_7503,N_7497);
or UO_301 (O_301,N_5662,N_5967);
or UO_302 (O_302,N_9885,N_9813);
nand UO_303 (O_303,N_9057,N_5858);
nor UO_304 (O_304,N_9332,N_9714);
or UO_305 (O_305,N_6443,N_9550);
nand UO_306 (O_306,N_6941,N_6607);
or UO_307 (O_307,N_7481,N_6992);
nor UO_308 (O_308,N_9777,N_9704);
nand UO_309 (O_309,N_6272,N_6505);
nand UO_310 (O_310,N_8203,N_7964);
or UO_311 (O_311,N_6105,N_9434);
nor UO_312 (O_312,N_6562,N_6305);
nand UO_313 (O_313,N_7738,N_9187);
and UO_314 (O_314,N_5570,N_8260);
nand UO_315 (O_315,N_7240,N_8753);
or UO_316 (O_316,N_9834,N_7102);
nand UO_317 (O_317,N_8664,N_6241);
nor UO_318 (O_318,N_6449,N_9455);
nor UO_319 (O_319,N_8980,N_5228);
nand UO_320 (O_320,N_9599,N_9725);
nor UO_321 (O_321,N_8151,N_5501);
nor UO_322 (O_322,N_9962,N_6849);
or UO_323 (O_323,N_5612,N_9867);
and UO_324 (O_324,N_8013,N_6392);
or UO_325 (O_325,N_6214,N_6764);
xnor UO_326 (O_326,N_8646,N_6005);
nand UO_327 (O_327,N_6994,N_7270);
nor UO_328 (O_328,N_7699,N_8271);
nand UO_329 (O_329,N_8897,N_5197);
and UO_330 (O_330,N_9583,N_5194);
nand UO_331 (O_331,N_6637,N_5424);
and UO_332 (O_332,N_9090,N_7444);
nor UO_333 (O_333,N_6331,N_5039);
nor UO_334 (O_334,N_7374,N_5729);
and UO_335 (O_335,N_6503,N_7107);
or UO_336 (O_336,N_8276,N_9687);
xnor UO_337 (O_337,N_8949,N_5659);
and UO_338 (O_338,N_6018,N_9612);
and UO_339 (O_339,N_6107,N_9832);
nand UO_340 (O_340,N_8935,N_8672);
or UO_341 (O_341,N_8892,N_5144);
nor UO_342 (O_342,N_7571,N_7605);
or UO_343 (O_343,N_6952,N_7106);
and UO_344 (O_344,N_7498,N_6006);
nand UO_345 (O_345,N_9791,N_7209);
nand UO_346 (O_346,N_9598,N_8077);
nor UO_347 (O_347,N_8768,N_8608);
nand UO_348 (O_348,N_9163,N_9568);
nor UO_349 (O_349,N_6337,N_8858);
and UO_350 (O_350,N_5530,N_7650);
or UO_351 (O_351,N_6661,N_5465);
and UO_352 (O_352,N_7405,N_8046);
nand UO_353 (O_353,N_5615,N_7865);
nand UO_354 (O_354,N_9457,N_6929);
and UO_355 (O_355,N_8232,N_9493);
and UO_356 (O_356,N_9465,N_8713);
xor UO_357 (O_357,N_7495,N_7161);
and UO_358 (O_358,N_6440,N_9403);
and UO_359 (O_359,N_6977,N_9334);
and UO_360 (O_360,N_6106,N_8543);
or UO_361 (O_361,N_5416,N_6461);
or UO_362 (O_362,N_7683,N_5367);
or UO_363 (O_363,N_8386,N_6603);
and UO_364 (O_364,N_7995,N_5982);
nor UO_365 (O_365,N_8380,N_5103);
and UO_366 (O_366,N_8631,N_6734);
and UO_367 (O_367,N_6856,N_9385);
nor UO_368 (O_368,N_9222,N_5296);
nand UO_369 (O_369,N_7262,N_8869);
xor UO_370 (O_370,N_7536,N_9967);
or UO_371 (O_371,N_9665,N_6772);
nand UO_372 (O_372,N_9703,N_9153);
nand UO_373 (O_373,N_5841,N_6870);
nand UO_374 (O_374,N_7383,N_6215);
nand UO_375 (O_375,N_7425,N_6934);
nand UO_376 (O_376,N_6459,N_5239);
or UO_377 (O_377,N_6063,N_5310);
nor UO_378 (O_378,N_8675,N_7434);
or UO_379 (O_379,N_6695,N_8560);
or UO_380 (O_380,N_8711,N_6071);
nand UO_381 (O_381,N_5254,N_9584);
and UO_382 (O_382,N_6098,N_7798);
or UO_383 (O_383,N_5546,N_6198);
or UO_384 (O_384,N_9776,N_7523);
nand UO_385 (O_385,N_5816,N_5504);
and UO_386 (O_386,N_6533,N_8382);
nand UO_387 (O_387,N_7411,N_6447);
nand UO_388 (O_388,N_5166,N_8889);
or UO_389 (O_389,N_5232,N_8371);
or UO_390 (O_390,N_6148,N_6843);
nor UO_391 (O_391,N_5647,N_6435);
and UO_392 (O_392,N_6055,N_7090);
nand UO_393 (O_393,N_5448,N_8094);
or UO_394 (O_394,N_8509,N_9246);
or UO_395 (O_395,N_9921,N_6878);
nand UO_396 (O_396,N_6846,N_5972);
nor UO_397 (O_397,N_9892,N_7880);
nor UO_398 (O_398,N_6610,N_5309);
or UO_399 (O_399,N_5145,N_5329);
nand UO_400 (O_400,N_9410,N_7930);
nor UO_401 (O_401,N_5994,N_8089);
and UO_402 (O_402,N_7395,N_7560);
nor UO_403 (O_403,N_8377,N_6041);
nor UO_404 (O_404,N_9480,N_8373);
and UO_405 (O_405,N_9843,N_8978);
or UO_406 (O_406,N_8895,N_9156);
nor UO_407 (O_407,N_6201,N_8896);
and UO_408 (O_408,N_7138,N_5810);
nand UO_409 (O_409,N_8590,N_8494);
nand UO_410 (O_410,N_6149,N_7979);
nor UO_411 (O_411,N_8921,N_8067);
nand UO_412 (O_412,N_9245,N_8473);
nand UO_413 (O_413,N_6341,N_7629);
nor UO_414 (O_414,N_5948,N_8644);
and UO_415 (O_415,N_7191,N_9159);
nand UO_416 (O_416,N_6388,N_8599);
nand UO_417 (O_417,N_8143,N_7134);
or UO_418 (O_418,N_8449,N_5025);
nand UO_419 (O_419,N_9753,N_7127);
and UO_420 (O_420,N_7604,N_8326);
nand UO_421 (O_421,N_8202,N_7538);
and UO_422 (O_422,N_9357,N_9508);
nand UO_423 (O_423,N_6378,N_6419);
or UO_424 (O_424,N_7144,N_7486);
nor UO_425 (O_425,N_6147,N_8801);
and UO_426 (O_426,N_7762,N_5259);
nand UO_427 (O_427,N_6452,N_7895);
nor UO_428 (O_428,N_8239,N_7765);
nand UO_429 (O_429,N_5564,N_5289);
and UO_430 (O_430,N_9001,N_6545);
and UO_431 (O_431,N_9323,N_6693);
nor UO_432 (O_432,N_8968,N_8286);
and UO_433 (O_433,N_6426,N_8398);
and UO_434 (O_434,N_5753,N_5026);
nor UO_435 (O_435,N_9435,N_8594);
or UO_436 (O_436,N_8910,N_7421);
nand UO_437 (O_437,N_6658,N_9975);
nand UO_438 (O_438,N_9893,N_7731);
nand UO_439 (O_439,N_8475,N_5730);
nor UO_440 (O_440,N_7999,N_8826);
xor UO_441 (O_441,N_9995,N_6774);
or UO_442 (O_442,N_7462,N_8650);
nor UO_443 (O_443,N_7812,N_7787);
nor UO_444 (O_444,N_7407,N_5327);
nor UO_445 (O_445,N_9537,N_9579);
nand UO_446 (O_446,N_7833,N_9838);
nor UO_447 (O_447,N_8430,N_6894);
or UO_448 (O_448,N_9506,N_6068);
nand UO_449 (O_449,N_8440,N_5766);
nand UO_450 (O_450,N_8491,N_7581);
nand UO_451 (O_451,N_7427,N_9067);
nor UO_452 (O_452,N_9318,N_6030);
and UO_453 (O_453,N_7242,N_7456);
nand UO_454 (O_454,N_5951,N_7148);
nand UO_455 (O_455,N_5543,N_8160);
and UO_456 (O_456,N_6137,N_9726);
nor UO_457 (O_457,N_6932,N_8347);
and UO_458 (O_458,N_9233,N_7563);
nand UO_459 (O_459,N_6358,N_8657);
xor UO_460 (O_460,N_8374,N_9339);
nor UO_461 (O_461,N_9990,N_7649);
nand UO_462 (O_462,N_5518,N_9118);
or UO_463 (O_463,N_7611,N_6943);
and UO_464 (O_464,N_7911,N_6382);
or UO_465 (O_465,N_6403,N_9243);
or UO_466 (O_466,N_7801,N_5364);
nand UO_467 (O_467,N_7009,N_5204);
or UO_468 (O_468,N_8987,N_8827);
or UO_469 (O_469,N_5954,N_6247);
nor UO_470 (O_470,N_5099,N_6267);
xor UO_471 (O_471,N_7759,N_6357);
or UO_472 (O_472,N_7514,N_6375);
or UO_473 (O_473,N_5298,N_9325);
and UO_474 (O_474,N_9381,N_7363);
and UO_475 (O_475,N_9590,N_6521);
nor UO_476 (O_476,N_8503,N_6266);
nand UO_477 (O_477,N_6093,N_5946);
or UO_478 (O_478,N_9382,N_6815);
xnor UO_479 (O_479,N_7573,N_5558);
or UO_480 (O_480,N_6464,N_5648);
nor UO_481 (O_481,N_6078,N_6957);
nand UO_482 (O_482,N_8368,N_8257);
xor UO_483 (O_483,N_6806,N_8670);
xor UO_484 (O_484,N_9863,N_6225);
or UO_485 (O_485,N_8736,N_7452);
nand UO_486 (O_486,N_8931,N_5555);
nand UO_487 (O_487,N_5750,N_9162);
and UO_488 (O_488,N_6987,N_5708);
or UO_489 (O_489,N_7883,N_7672);
nor UO_490 (O_490,N_9668,N_9283);
nand UO_491 (O_491,N_9823,N_5275);
or UO_492 (O_492,N_7433,N_6437);
nor UO_493 (O_493,N_6971,N_9845);
nand UO_494 (O_494,N_6277,N_7335);
nand UO_495 (O_495,N_5561,N_9572);
and UO_496 (O_496,N_9578,N_6594);
nor UO_497 (O_497,N_7101,N_8872);
or UO_498 (O_498,N_6062,N_6996);
nand UO_499 (O_499,N_6867,N_9908);
nor UO_500 (O_500,N_9367,N_7217);
or UO_501 (O_501,N_6310,N_8287);
or UO_502 (O_502,N_5668,N_8942);
nor UO_503 (O_503,N_6402,N_7332);
or UO_504 (O_504,N_5808,N_6619);
nand UO_505 (O_505,N_7836,N_8808);
or UO_506 (O_506,N_9121,N_8460);
nand UO_507 (O_507,N_9469,N_9387);
xor UO_508 (O_508,N_5877,N_7851);
or UO_509 (O_509,N_5798,N_8359);
and UO_510 (O_510,N_7805,N_9066);
and UO_511 (O_511,N_5670,N_7515);
or UO_512 (O_512,N_8983,N_9888);
or UO_513 (O_513,N_9206,N_6504);
or UO_514 (O_514,N_8187,N_7914);
nand UO_515 (O_515,N_9218,N_8096);
or UO_516 (O_516,N_6291,N_7183);
or UO_517 (O_517,N_5557,N_7220);
nand UO_518 (O_518,N_8643,N_6776);
or UO_519 (O_519,N_5109,N_8076);
or UO_520 (O_520,N_7760,N_6668);
and UO_521 (O_521,N_9911,N_5210);
or UO_522 (O_522,N_8390,N_8190);
nand UO_523 (O_523,N_7669,N_6763);
nor UO_524 (O_524,N_6700,N_7966);
and UO_525 (O_525,N_5579,N_5572);
or UO_526 (O_526,N_8917,N_9869);
and UO_527 (O_527,N_6576,N_6074);
nor UO_528 (O_528,N_6818,N_8112);
nand UO_529 (O_529,N_7155,N_7388);
and UO_530 (O_530,N_7973,N_5385);
and UO_531 (O_531,N_9278,N_8452);
and UO_532 (O_532,N_6446,N_9745);
and UO_533 (O_533,N_9135,N_8701);
and UO_534 (O_534,N_5251,N_5560);
and UO_535 (O_535,N_6428,N_6370);
nor UO_536 (O_536,N_5550,N_8977);
or UO_537 (O_537,N_9825,N_6524);
nor UO_538 (O_538,N_6127,N_5497);
or UO_539 (O_539,N_6481,N_5945);
and UO_540 (O_540,N_7386,N_9084);
nor UO_541 (O_541,N_8125,N_7651);
or UO_542 (O_542,N_5939,N_7744);
and UO_543 (O_543,N_5390,N_6181);
nand UO_544 (O_544,N_8064,N_7969);
nor UO_545 (O_545,N_7113,N_8516);
nor UO_546 (O_546,N_8714,N_6877);
and UO_547 (O_547,N_8640,N_7843);
or UO_548 (O_548,N_5393,N_6664);
or UO_549 (O_549,N_6034,N_5848);
or UO_550 (O_550,N_9896,N_9750);
and UO_551 (O_551,N_9756,N_8063);
or UO_552 (O_552,N_5836,N_9299);
or UO_553 (O_553,N_7258,N_7994);
and UO_554 (O_554,N_8635,N_6342);
nand UO_555 (O_555,N_7397,N_6684);
nor UO_556 (O_556,N_7381,N_9044);
xor UO_557 (O_557,N_7680,N_8117);
xnor UO_558 (O_558,N_8540,N_7792);
or UO_559 (O_559,N_5495,N_6605);
or UO_560 (O_560,N_9577,N_8246);
nand UO_561 (O_561,N_7376,N_8088);
nor UO_562 (O_562,N_7584,N_5796);
and UO_563 (O_563,N_5869,N_6635);
nor UO_564 (O_564,N_8240,N_6840);
nor UO_565 (O_565,N_9010,N_6565);
and UO_566 (O_566,N_8211,N_5075);
nor UO_567 (O_567,N_5562,N_5107);
nand UO_568 (O_568,N_8134,N_8666);
or UO_569 (O_569,N_6336,N_6070);
and UO_570 (O_570,N_8749,N_5603);
nor UO_571 (O_571,N_7800,N_6741);
xnor UO_572 (O_572,N_5823,N_7779);
or UO_573 (O_573,N_9589,N_9047);
and UO_574 (O_574,N_5231,N_5807);
nand UO_575 (O_575,N_6376,N_8243);
nand UO_576 (O_576,N_5199,N_8536);
nor UO_577 (O_577,N_8705,N_5012);
or UO_578 (O_578,N_5157,N_5292);
nand UO_579 (O_579,N_5066,N_6479);
or UO_580 (O_580,N_6103,N_6907);
or UO_581 (O_581,N_9150,N_6978);
and UO_582 (O_582,N_5136,N_8721);
and UO_583 (O_583,N_8732,N_9585);
or UO_584 (O_584,N_5351,N_5034);
nand UO_585 (O_585,N_5198,N_5090);
nand UO_586 (O_586,N_7264,N_7714);
nor UO_587 (O_587,N_5682,N_9204);
nand UO_588 (O_588,N_8014,N_8297);
or UO_589 (O_589,N_7959,N_5122);
nor UO_590 (O_590,N_6230,N_5535);
and UO_591 (O_591,N_9916,N_8684);
or UO_592 (O_592,N_8913,N_5651);
nor UO_593 (O_593,N_9864,N_9126);
nand UO_594 (O_594,N_9468,N_9463);
nor UO_595 (O_595,N_9157,N_9889);
or UO_596 (O_596,N_5031,N_6417);
or UO_597 (O_597,N_5373,N_7761);
or UO_598 (O_598,N_6860,N_5588);
nor UO_599 (O_599,N_8846,N_8916);
or UO_600 (O_600,N_6096,N_8638);
xor UO_601 (O_601,N_9189,N_6257);
and UO_602 (O_602,N_7063,N_8493);
nand UO_603 (O_603,N_9170,N_6967);
or UO_604 (O_604,N_8496,N_6852);
xor UO_605 (O_605,N_5011,N_6016);
nor UO_606 (O_606,N_9949,N_9191);
and UO_607 (O_607,N_7899,N_7954);
nand UO_608 (O_608,N_5693,N_7389);
or UO_609 (O_609,N_7099,N_7903);
nand UO_610 (O_610,N_6736,N_9702);
or UO_611 (O_611,N_7214,N_5502);
or UO_612 (O_612,N_8512,N_8136);
nor UO_613 (O_613,N_9202,N_6749);
and UO_614 (O_614,N_5169,N_8803);
nand UO_615 (O_615,N_8029,N_8128);
and UO_616 (O_616,N_8244,N_7309);
and UO_617 (O_617,N_7081,N_6733);
or UO_618 (O_618,N_9406,N_5474);
nor UO_619 (O_619,N_7723,N_9722);
or UO_620 (O_620,N_6955,N_9265);
nor UO_621 (O_621,N_9692,N_7725);
or UO_622 (O_622,N_8810,N_9905);
or UO_623 (O_623,N_6007,N_5805);
nand UO_624 (O_624,N_5601,N_5273);
and UO_625 (O_625,N_6945,N_5265);
nand UO_626 (O_626,N_5229,N_6808);
nor UO_627 (O_627,N_7864,N_9989);
or UO_628 (O_628,N_8991,N_9257);
or UO_629 (O_629,N_5053,N_9174);
nor UO_630 (O_630,N_9479,N_6361);
xnor UO_631 (O_631,N_8676,N_9319);
nand UO_632 (O_632,N_8099,N_6876);
nand UO_633 (O_633,N_6323,N_7437);
nand UO_634 (O_634,N_7799,N_9849);
nor UO_635 (O_635,N_6350,N_9199);
nor UO_636 (O_636,N_8389,N_8402);
and UO_637 (O_637,N_5001,N_7657);
or UO_638 (O_638,N_6143,N_8914);
nand UO_639 (O_639,N_8806,N_5046);
and UO_640 (O_640,N_9474,N_5548);
nand UO_641 (O_641,N_5904,N_7720);
or UO_642 (O_642,N_9490,N_6020);
or UO_643 (O_643,N_5071,N_6258);
nor UO_644 (O_644,N_5513,N_5450);
nand UO_645 (O_645,N_8852,N_6397);
and UO_646 (O_646,N_7603,N_8039);
nand UO_647 (O_647,N_6606,N_7070);
and UO_648 (O_648,N_9142,N_7280);
and UO_649 (O_649,N_9784,N_6442);
and UO_650 (O_650,N_8065,N_5632);
or UO_651 (O_651,N_8174,N_6113);
nand UO_652 (O_652,N_9559,N_8334);
nand UO_653 (O_653,N_7574,N_6076);
nor UO_654 (O_654,N_7848,N_6160);
nor UO_655 (O_655,N_9169,N_5690);
nand UO_656 (O_656,N_9937,N_5019);
nand UO_657 (O_657,N_9681,N_8403);
nand UO_658 (O_658,N_5457,N_6848);
nand UO_659 (O_659,N_5466,N_7265);
and UO_660 (O_660,N_6814,N_5786);
nand UO_661 (O_661,N_6448,N_5536);
nor UO_662 (O_662,N_5527,N_6282);
and UO_663 (O_663,N_7945,N_8600);
nand UO_664 (O_664,N_6054,N_8186);
or UO_665 (O_665,N_7449,N_6125);
and UO_666 (O_666,N_9486,N_7272);
nand UO_667 (O_667,N_6154,N_5923);
nor UO_668 (O_668,N_6367,N_8121);
nand UO_669 (O_669,N_5964,N_5936);
or UO_670 (O_670,N_7492,N_7279);
and UO_671 (O_671,N_8344,N_7900);
or UO_672 (O_672,N_7580,N_5286);
nor UO_673 (O_673,N_5261,N_9024);
or UO_674 (O_674,N_8148,N_7464);
nand UO_675 (O_675,N_8939,N_5783);
nand UO_676 (O_676,N_6985,N_8683);
and UO_677 (O_677,N_9974,N_6909);
and UO_678 (O_678,N_7011,N_7673);
and UO_679 (O_679,N_9723,N_8083);
nand UO_680 (O_680,N_9000,N_7827);
nand UO_681 (O_681,N_8661,N_5797);
or UO_682 (O_682,N_9096,N_7844);
xor UO_683 (O_683,N_9814,N_7674);
or UO_684 (O_684,N_6963,N_6950);
and UO_685 (O_685,N_9201,N_6537);
and UO_686 (O_686,N_7417,N_9352);
nand UO_687 (O_687,N_7366,N_7849);
and UO_688 (O_688,N_9669,N_8192);
nor UO_689 (O_689,N_8318,N_8304);
and UO_690 (O_690,N_5763,N_5325);
and UO_691 (O_691,N_6119,N_7057);
nor UO_692 (O_692,N_7233,N_5037);
or UO_693 (O_693,N_5679,N_9327);
nand UO_694 (O_694,N_9999,N_9019);
nand UO_695 (O_695,N_8124,N_7965);
xor UO_696 (O_696,N_9076,N_8066);
or UO_697 (O_697,N_9926,N_8652);
or UO_698 (O_698,N_7310,N_6083);
nand UO_699 (O_699,N_5941,N_7614);
nand UO_700 (O_700,N_5529,N_7484);
or UO_701 (O_701,N_9171,N_6974);
xor UO_702 (O_702,N_6425,N_5743);
nor UO_703 (O_703,N_7307,N_9293);
nand UO_704 (O_704,N_7594,N_6269);
or UO_705 (O_705,N_9093,N_6835);
nand UO_706 (O_706,N_6236,N_5788);
and UO_707 (O_707,N_7311,N_5879);
and UO_708 (O_708,N_9601,N_7542);
xnor UO_709 (O_709,N_8399,N_6713);
nand UO_710 (O_710,N_7121,N_5928);
or UO_711 (O_711,N_7961,N_7198);
nand UO_712 (O_712,N_7042,N_6084);
nand UO_713 (O_713,N_9452,N_7219);
and UO_714 (O_714,N_8554,N_8255);
nand UO_715 (O_715,N_8750,N_5567);
or UO_716 (O_716,N_5965,N_5041);
and UO_717 (O_717,N_7532,N_8637);
nor UO_718 (O_718,N_5280,N_5909);
or UO_719 (O_719,N_5713,N_6240);
nand UO_720 (O_720,N_8109,N_8302);
nand UO_721 (O_721,N_8573,N_8696);
nand UO_722 (O_722,N_9039,N_9183);
and UO_723 (O_723,N_6276,N_6989);
and UO_724 (O_724,N_7377,N_5866);
nand UO_725 (O_725,N_5441,N_9220);
nor UO_726 (O_726,N_9980,N_6216);
nand UO_727 (O_727,N_8004,N_8529);
nand UO_728 (O_728,N_9628,N_9538);
nand UO_729 (O_729,N_7774,N_6604);
or UO_730 (O_730,N_5578,N_7870);
and UO_731 (O_731,N_8547,N_6900);
and UO_732 (O_732,N_7103,N_9284);
and UO_733 (O_733,N_6047,N_5035);
nor UO_734 (O_734,N_9858,N_6434);
or UO_735 (O_735,N_8719,N_8902);
nand UO_736 (O_736,N_9830,N_7775);
or UO_737 (O_737,N_8967,N_5220);
or UO_738 (O_738,N_8710,N_6366);
nor UO_739 (O_739,N_5970,N_5361);
and UO_740 (O_740,N_7847,N_7116);
nor UO_741 (O_741,N_6097,N_8454);
and UO_742 (O_742,N_8510,N_9466);
and UO_743 (O_743,N_9755,N_9046);
or UO_744 (O_744,N_7468,N_5999);
nand UO_745 (O_745,N_5263,N_5718);
nand UO_746 (O_746,N_5069,N_8378);
or UO_747 (O_747,N_7137,N_7210);
nor UO_748 (O_748,N_7392,N_8438);
or UO_749 (O_749,N_8966,N_8080);
or UO_750 (O_750,N_5089,N_9120);
or UO_751 (O_751,N_5410,N_8568);
and UO_752 (O_752,N_9034,N_5802);
and UO_753 (O_753,N_6666,N_7645);
and UO_754 (O_754,N_7852,N_7109);
nor UO_755 (O_755,N_7339,N_7975);
nand UO_756 (O_756,N_5167,N_7306);
and UO_757 (O_757,N_7064,N_9985);
or UO_758 (O_758,N_8959,N_7092);
and UO_759 (O_759,N_5193,N_6899);
or UO_760 (O_760,N_7074,N_8611);
and UO_761 (O_761,N_5043,N_8406);
nor UO_762 (O_762,N_9637,N_9165);
and UO_763 (O_763,N_9366,N_5672);
nand UO_764 (O_764,N_5880,N_8618);
nor UO_765 (O_765,N_6066,N_9643);
nand UO_766 (O_766,N_7795,N_7746);
nand UO_767 (O_767,N_8290,N_6492);
or UO_768 (O_768,N_6617,N_6384);
nand UO_769 (O_769,N_5412,N_6209);
or UO_770 (O_770,N_5697,N_9812);
nand UO_771 (O_771,N_6613,N_7970);
nand UO_772 (O_772,N_9767,N_5105);
nor UO_773 (O_773,N_6218,N_5754);
or UO_774 (O_774,N_7811,N_6547);
nand UO_775 (O_775,N_7676,N_5212);
nand UO_776 (O_776,N_8425,N_7838);
nor UO_777 (O_777,N_8090,N_6360);
nand UO_778 (O_778,N_9343,N_6972);
or UO_779 (O_779,N_9633,N_5224);
and UO_780 (O_780,N_9317,N_6322);
nor UO_781 (O_781,N_8952,N_8215);
or UO_782 (O_782,N_9459,N_7263);
nand UO_783 (O_783,N_8253,N_6863);
nor UO_784 (O_784,N_6471,N_5215);
nand UO_785 (O_785,N_8689,N_5120);
and UO_786 (O_786,N_6532,N_9391);
and UO_787 (O_787,N_9033,N_9411);
nor UO_788 (O_788,N_8356,N_9856);
nand UO_789 (O_789,N_9890,N_6719);
nand UO_790 (O_790,N_5635,N_6372);
nand UO_791 (O_791,N_8395,N_8229);
nor UO_792 (O_792,N_5211,N_8233);
nor UO_793 (O_793,N_6043,N_6534);
nor UO_794 (O_794,N_9312,N_6286);
or UO_795 (O_795,N_9547,N_7627);
or UO_796 (O_796,N_7606,N_6884);
or UO_797 (O_797,N_9672,N_6183);
nor UO_798 (O_798,N_6911,N_8789);
or UO_799 (O_799,N_6009,N_7781);
or UO_800 (O_800,N_5943,N_7777);
nor UO_801 (O_801,N_6317,N_5222);
or UO_802 (O_802,N_7256,N_8413);
or UO_803 (O_803,N_9464,N_5278);
nor UO_804 (O_804,N_9514,N_5068);
nand UO_805 (O_805,N_7666,N_5687);
or UO_806 (O_806,N_5082,N_9230);
and UO_807 (O_807,N_8769,N_9748);
and UO_808 (O_808,N_6970,N_9787);
or UO_809 (O_809,N_9884,N_7448);
nand UO_810 (O_810,N_5436,N_6023);
nor UO_811 (O_811,N_6179,N_8149);
nor UO_812 (O_812,N_7068,N_8682);
and UO_813 (O_813,N_5126,N_8026);
and UO_814 (O_814,N_6677,N_5846);
nor UO_815 (O_815,N_8025,N_9959);
and UO_816 (O_816,N_8350,N_5541);
nand UO_817 (O_817,N_5637,N_5362);
or UO_818 (O_818,N_7253,N_8263);
nor UO_819 (O_819,N_7129,N_6374);
and UO_820 (O_820,N_9433,N_8035);
nor UO_821 (O_821,N_6889,N_8900);
nand UO_822 (O_822,N_5723,N_8989);
and UO_823 (O_823,N_8565,N_9857);
nand UO_824 (O_824,N_5956,N_6052);
and UO_825 (O_825,N_6186,N_7043);
or UO_826 (O_826,N_6858,N_6979);
and UO_827 (O_827,N_9345,N_6445);
nand UO_828 (O_828,N_7414,N_6510);
or UO_829 (O_829,N_9023,N_8439);
nor UO_830 (O_830,N_7488,N_9361);
nand UO_831 (O_831,N_9258,N_7315);
or UO_832 (O_832,N_8420,N_5978);
nand UO_833 (O_833,N_8375,N_6253);
nand UO_834 (O_834,N_8859,N_9528);
xnor UO_835 (O_835,N_7013,N_9591);
nor UO_836 (O_836,N_7875,N_5926);
and UO_837 (O_837,N_9684,N_5079);
nand UO_838 (O_838,N_9659,N_6914);
nand UO_839 (O_839,N_8415,N_6833);
and UO_840 (O_840,N_9416,N_8712);
and UO_841 (O_841,N_8011,N_7472);
nand UO_842 (O_842,N_7664,N_5675);
or UO_843 (O_843,N_6608,N_6423);
nor UO_844 (O_844,N_8157,N_8372);
or UO_845 (O_845,N_7176,N_5863);
nand UO_846 (O_846,N_9503,N_5902);
nand UO_847 (O_847,N_8538,N_6058);
nor UO_848 (O_848,N_7766,N_5326);
or UO_849 (O_849,N_6879,N_6279);
nand UO_850 (O_850,N_7082,N_9127);
or UO_851 (O_851,N_6246,N_8764);
nor UO_852 (O_852,N_5328,N_5405);
nand UO_853 (O_853,N_9558,N_7295);
nor UO_854 (O_854,N_8537,N_5892);
and UO_855 (O_855,N_8018,N_8742);
and UO_856 (O_856,N_5324,N_5381);
and UO_857 (O_857,N_5359,N_7909);
nand UO_858 (O_858,N_5400,N_9859);
nor UO_859 (O_859,N_9115,N_6256);
nand UO_860 (O_860,N_7257,N_5580);
and UO_861 (O_861,N_5270,N_7184);
nand UO_862 (O_862,N_5354,N_7373);
xor UO_863 (O_863,N_9504,N_8853);
nor UO_864 (O_864,N_8104,N_6077);
and UO_865 (O_865,N_9394,N_8369);
xnor UO_866 (O_866,N_9575,N_7593);
nor UO_867 (O_867,N_7862,N_5883);
and UO_868 (O_868,N_7020,N_9979);
and UO_869 (O_869,N_5547,N_8948);
and UO_870 (O_870,N_8069,N_7187);
nand UO_871 (O_871,N_5790,N_5825);
and UO_872 (O_872,N_9371,N_6176);
nor UO_873 (O_873,N_5645,N_5106);
nor UO_874 (O_874,N_5820,N_8300);
and UO_875 (O_875,N_9925,N_8316);
nand UO_876 (O_876,N_5279,N_6362);
or UO_877 (O_877,N_5454,N_9447);
nor UO_878 (O_878,N_5119,N_5171);
and UO_879 (O_879,N_6933,N_5517);
or UO_880 (O_880,N_8990,N_7040);
nand UO_881 (O_881,N_6930,N_5340);
and UO_882 (O_882,N_8106,N_8639);
nor UO_883 (O_883,N_7543,N_6869);
nor UO_884 (O_884,N_6755,N_8745);
or UO_885 (O_885,N_8893,N_5854);
or UO_886 (O_886,N_6261,N_7986);
or UO_887 (O_887,N_7249,N_8464);
nand UO_888 (O_888,N_7243,N_8486);
and UO_889 (O_889,N_8075,N_7917);
or UO_890 (O_890,N_7521,N_9125);
nand UO_891 (O_891,N_5990,N_8277);
and UO_892 (O_892,N_7244,N_9179);
nand UO_893 (O_893,N_7331,N_9632);
nand UO_894 (O_894,N_9390,N_6725);
and UO_895 (O_895,N_9713,N_6102);
and UO_896 (O_896,N_5060,N_6036);
and UO_897 (O_897,N_9117,N_9586);
or UO_898 (O_898,N_9676,N_7876);
nor UO_899 (O_899,N_7826,N_9790);
and UO_900 (O_900,N_5028,N_8795);
nand UO_901 (O_901,N_7422,N_8688);
or UO_902 (O_902,N_8314,N_6495);
and UO_903 (O_903,N_6544,N_8820);
and UO_904 (O_904,N_6721,N_6162);
nand UO_905 (O_905,N_7868,N_8126);
or UO_906 (O_906,N_5134,N_9679);
and UO_907 (O_907,N_7544,N_7482);
nand UO_908 (O_908,N_8468,N_5881);
and UO_909 (O_909,N_5709,N_5319);
or UO_910 (O_910,N_7313,N_6226);
or UO_911 (O_911,N_7048,N_8325);
or UO_912 (O_912,N_8922,N_6645);
and UO_913 (O_913,N_6067,N_5602);
or UO_914 (O_914,N_5537,N_9744);
or UO_915 (O_915,N_7200,N_7324);
nor UO_916 (O_916,N_6997,N_9570);
and UO_917 (O_917,N_6297,N_6819);
nor UO_918 (O_918,N_7124,N_5238);
nor UO_919 (O_919,N_5568,N_7770);
or UO_920 (O_920,N_6995,N_7086);
nor UO_921 (O_921,N_6540,N_7114);
nand UO_922 (O_922,N_9365,N_6556);
and UO_923 (O_923,N_8780,N_6529);
nor UO_924 (O_924,N_8092,N_5403);
nor UO_925 (O_925,N_6469,N_6513);
nor UO_926 (O_926,N_8336,N_8053);
nor UO_927 (O_927,N_9498,N_5915);
or UO_928 (O_928,N_8293,N_7222);
nor UO_929 (O_929,N_6925,N_8206);
nor UO_930 (O_930,N_6506,N_9262);
nand UO_931 (O_931,N_7382,N_8988);
or UO_932 (O_932,N_8934,N_9927);
and UO_933 (O_933,N_8267,N_6773);
nand UO_934 (O_934,N_7202,N_7493);
nand UO_935 (O_935,N_8471,N_5665);
or UO_936 (O_936,N_8033,N_8313);
nor UO_937 (O_937,N_9883,N_8868);
or UO_938 (O_938,N_5893,N_6508);
and UO_939 (O_939,N_7182,N_7108);
or UO_940 (O_940,N_9485,N_5993);
xnor UO_941 (O_941,N_7884,N_9705);
nand UO_942 (O_942,N_5442,N_5225);
or UO_943 (O_943,N_7607,N_7635);
nand UO_944 (O_944,N_6762,N_5336);
nor UO_945 (O_945,N_9075,N_6352);
or UO_946 (O_946,N_6778,N_9407);
nor UO_947 (O_947,N_5116,N_6998);
or UO_948 (O_948,N_5669,N_9602);
nor UO_949 (O_949,N_5551,N_6866);
and UO_950 (O_950,N_5438,N_9718);
and UO_951 (O_951,N_5472,N_7769);
or UO_952 (O_952,N_6390,N_6551);
and UO_953 (O_953,N_6885,N_9158);
and UO_954 (O_954,N_6335,N_9820);
or UO_955 (O_955,N_6326,N_5077);
and UO_956 (O_956,N_9106,N_5918);
nand UO_957 (O_957,N_7687,N_7246);
or UO_958 (O_958,N_5287,N_5064);
and UO_959 (O_959,N_5100,N_6851);
or UO_960 (O_960,N_8278,N_9438);
nor UO_961 (O_961,N_7891,N_7400);
or UO_962 (O_962,N_6141,N_6359);
nand UO_963 (O_963,N_5409,N_6525);
or UO_964 (O_964,N_6633,N_6396);
and UO_965 (O_965,N_5302,N_8185);
and UO_966 (O_966,N_8874,N_5226);
nor UO_967 (O_967,N_7940,N_5811);
nor UO_968 (O_968,N_7146,N_8823);
nor UO_969 (O_969,N_6429,N_8383);
nand UO_970 (O_970,N_6205,N_6024);
and UO_971 (O_971,N_8183,N_6117);
nor UO_972 (O_972,N_6122,N_7259);
nand UO_973 (O_973,N_7236,N_8552);
and UO_974 (O_974,N_7599,N_9259);
nor UO_975 (O_975,N_6486,N_5986);
nor UO_976 (O_976,N_9419,N_7247);
and UO_977 (O_977,N_7729,N_6535);
or UO_978 (O_978,N_8944,N_9738);
nor UO_979 (O_979,N_9214,N_5268);
nor UO_980 (O_980,N_6653,N_7590);
nor UO_981 (O_981,N_8055,N_8867);
nand UO_982 (O_982,N_9151,N_6786);
nand UO_983 (O_983,N_8528,N_8733);
nand UO_984 (O_984,N_7439,N_8017);
nand UO_985 (O_985,N_8671,N_6651);
and UO_986 (O_986,N_6753,N_9355);
or UO_987 (O_987,N_5015,N_5252);
nand UO_988 (O_988,N_8855,N_5824);
nand UO_989 (O_989,N_6057,N_9061);
and UO_990 (O_990,N_9792,N_8167);
nor UO_991 (O_991,N_8179,N_9835);
nand UO_992 (O_992,N_5281,N_7845);
nor UO_993 (O_993,N_9700,N_9821);
and UO_994 (O_994,N_8483,N_8962);
and UO_995 (O_995,N_5433,N_5707);
or UO_996 (O_996,N_5725,N_6767);
nand UO_997 (O_997,N_7337,N_5514);
or UO_998 (O_998,N_8037,N_5657);
or UO_999 (O_999,N_9296,N_7079);
nor UO_1000 (O_1000,N_9018,N_7688);
xnor UO_1001 (O_1001,N_9155,N_7718);
and UO_1002 (O_1002,N_9473,N_5073);
and UO_1003 (O_1003,N_5914,N_5556);
nor UO_1004 (O_1004,N_6779,N_6180);
nand UO_1005 (O_1005,N_5489,N_5780);
nand UO_1006 (O_1006,N_8744,N_8549);
and UO_1007 (O_1007,N_8953,N_9128);
nand UO_1008 (O_1008,N_5566,N_9868);
xnor UO_1009 (O_1009,N_6100,N_7906);
nor UO_1010 (O_1010,N_6642,N_8028);
nor UO_1011 (O_1011,N_6212,N_9610);
nor UO_1012 (O_1012,N_7447,N_9442);
or UO_1013 (O_1013,N_5852,N_9604);
or UO_1014 (O_1014,N_7626,N_5180);
or UO_1015 (O_1015,N_6138,N_5756);
or UO_1016 (O_1016,N_5542,N_5313);
xor UO_1017 (O_1017,N_6690,N_5680);
nor UO_1018 (O_1018,N_8890,N_6944);
nand UO_1019 (O_1019,N_5768,N_9229);
nor UO_1020 (O_1020,N_5486,N_7570);
xor UO_1021 (O_1021,N_8147,N_8556);
and UO_1022 (O_1022,N_5471,N_9441);
or UO_1023 (O_1023,N_9002,N_5076);
nand UO_1024 (O_1024,N_6931,N_7842);
and UO_1025 (O_1025,N_6011,N_6451);
nand UO_1026 (O_1026,N_6602,N_8901);
and UO_1027 (O_1027,N_7126,N_5311);
nor UO_1028 (O_1028,N_9654,N_6164);
or UO_1029 (O_1029,N_6830,N_6981);
nor UO_1030 (O_1030,N_8794,N_5806);
xnor UO_1031 (O_1031,N_6829,N_8957);
xnor UO_1032 (O_1032,N_8003,N_9805);
nor UO_1033 (O_1033,N_6886,N_6916);
nand UO_1034 (O_1034,N_9078,N_5255);
or UO_1035 (O_1035,N_7281,N_6675);
or UO_1036 (O_1036,N_7615,N_5801);
nor UO_1037 (O_1037,N_6328,N_7788);
nor UO_1038 (O_1038,N_8985,N_9964);
nor UO_1039 (O_1039,N_6185,N_5425);
nand UO_1040 (O_1040,N_5294,N_9261);
nor UO_1041 (O_1041,N_9569,N_5352);
nand UO_1042 (O_1042,N_8162,N_9819);
and UO_1043 (O_1043,N_6040,N_9742);
or UO_1044 (O_1044,N_6457,N_9328);
nor UO_1045 (O_1045,N_8443,N_5835);
nor UO_1046 (O_1046,N_5681,N_8474);
or UO_1047 (O_1047,N_9124,N_5609);
and UO_1048 (O_1048,N_7416,N_9372);
and UO_1049 (O_1049,N_9059,N_9540);
nor UO_1050 (O_1050,N_7932,N_7188);
nor UO_1051 (O_1051,N_7423,N_5677);
nor UO_1052 (O_1052,N_5997,N_7136);
nand UO_1053 (O_1053,N_9645,N_6953);
and UO_1054 (O_1054,N_8176,N_5701);
and UO_1055 (O_1055,N_6917,N_6954);
or UO_1056 (O_1056,N_7457,N_9565);
nor UO_1057 (O_1057,N_8587,N_6827);
nor UO_1058 (O_1058,N_9673,N_6896);
or UO_1059 (O_1059,N_8501,N_9686);
nand UO_1060 (O_1060,N_5739,N_6343);
nand UO_1061 (O_1061,N_6104,N_9011);
nor UO_1062 (O_1062,N_6416,N_6649);
and UO_1063 (O_1063,N_8986,N_9852);
and UO_1064 (O_1064,N_9931,N_8667);
nand UO_1065 (O_1065,N_9846,N_7715);
or UO_1066 (O_1066,N_5097,N_5344);
or UO_1067 (O_1067,N_9505,N_6622);
or UO_1068 (O_1068,N_5947,N_7878);
or UO_1069 (O_1069,N_7266,N_7935);
nand UO_1070 (O_1070,N_7094,N_8481);
nand UO_1071 (O_1071,N_6462,N_6968);
nand UO_1072 (O_1072,N_5512,N_5200);
nor UO_1073 (O_1073,N_5080,N_5640);
and UO_1074 (O_1074,N_9488,N_8663);
and UO_1075 (O_1075,N_9682,N_9288);
and UO_1076 (O_1076,N_7956,N_8653);
nor UO_1077 (O_1077,N_8364,N_5581);
nor UO_1078 (O_1078,N_8264,N_8972);
or UO_1079 (O_1079,N_5257,N_7071);
nand UO_1080 (O_1080,N_6735,N_9897);
or UO_1081 (O_1081,N_7888,N_5575);
nand UO_1082 (O_1082,N_8456,N_5207);
or UO_1083 (O_1083,N_8699,N_7510);
nor UO_1084 (O_1084,N_5894,N_8583);
nor UO_1085 (O_1085,N_9729,N_9236);
and UO_1086 (O_1086,N_6329,N_7223);
or UO_1087 (O_1087,N_5002,N_6302);
and UO_1088 (O_1088,N_9072,N_7300);
or UO_1089 (O_1089,N_6538,N_7803);
nand UO_1090 (O_1090,N_6014,N_5132);
nand UO_1091 (O_1091,N_8131,N_9541);
or UO_1092 (O_1092,N_6887,N_6059);
and UO_1093 (O_1093,N_9359,N_5828);
and UO_1094 (O_1094,N_7298,N_9070);
or UO_1095 (O_1095,N_8703,N_5242);
or UO_1096 (O_1096,N_9014,N_6249);
or UO_1097 (O_1097,N_5192,N_8008);
nand UO_1098 (O_1098,N_5860,N_5318);
or UO_1099 (O_1099,N_8658,N_9217);
nor UO_1100 (O_1100,N_7360,N_5503);
and UO_1101 (O_1101,N_5803,N_8662);
and UO_1102 (O_1102,N_9089,N_5719);
nor UO_1103 (O_1103,N_9623,N_5961);
nand UO_1104 (O_1104,N_8656,N_9576);
or UO_1105 (O_1105,N_8175,N_8654);
or UO_1106 (O_1106,N_9175,N_7984);
nor UO_1107 (O_1107,N_6986,N_7065);
or UO_1108 (O_1108,N_6231,N_6873);
and UO_1109 (O_1109,N_6475,N_5415);
nor UO_1110 (O_1110,N_7062,N_6170);
and UO_1111 (O_1111,N_8844,N_5996);
nand UO_1112 (O_1112,N_8582,N_8191);
or UO_1113 (O_1113,N_9188,N_9636);
xor UO_1114 (O_1114,N_7637,N_9123);
nand UO_1115 (O_1115,N_8010,N_6581);
or UO_1116 (O_1116,N_7119,N_5714);
or UO_1117 (O_1117,N_9397,N_8164);
or UO_1118 (O_1118,N_5205,N_5884);
nand UO_1119 (O_1119,N_7278,N_5636);
or UO_1120 (O_1120,N_9335,N_9311);
and UO_1121 (O_1121,N_9720,N_7348);
nor UO_1122 (O_1122,N_7929,N_6862);
or UO_1123 (O_1123,N_8519,N_9211);
nor UO_1124 (O_1124,N_8381,N_8268);
or UO_1125 (O_1125,N_5621,N_7045);
and UO_1126 (O_1126,N_9301,N_9306);
nor UO_1127 (O_1127,N_8252,N_9392);
nor UO_1128 (O_1128,N_9456,N_8082);
or UO_1129 (O_1129,N_8702,N_8118);
nand UO_1130 (O_1130,N_8261,N_7678);
nand UO_1131 (O_1131,N_5772,N_5960);
nand UO_1132 (O_1132,N_8355,N_6671);
or UO_1133 (O_1133,N_7516,N_5995);
and UO_1134 (O_1134,N_9022,N_7697);
xnor UO_1135 (O_1135,N_7893,N_7084);
or UO_1136 (O_1136,N_9546,N_5453);
nand UO_1137 (O_1137,N_6502,N_5856);
and UO_1138 (O_1138,N_9148,N_5901);
nor UO_1139 (O_1139,N_9107,N_5906);
nor UO_1140 (O_1140,N_7567,N_8448);
nor UO_1141 (O_1141,N_7466,N_7147);
or UO_1142 (O_1142,N_6983,N_7110);
or UO_1143 (O_1143,N_6131,N_7863);
nor UO_1144 (O_1144,N_6701,N_5016);
nand UO_1145 (O_1145,N_5062,N_8700);
nor UO_1146 (O_1146,N_5769,N_5374);
nor UO_1147 (O_1147,N_9164,N_9105);
nand UO_1148 (O_1148,N_7248,N_5241);
nand UO_1149 (O_1149,N_5989,N_5004);
and UO_1150 (O_1150,N_9808,N_5377);
and UO_1151 (O_1151,N_5358,N_5975);
nand UO_1152 (O_1152,N_6306,N_7524);
and UO_1153 (O_1153,N_8317,N_7291);
and UO_1154 (O_1154,N_8165,N_9928);
and UO_1155 (O_1155,N_9140,N_7925);
or UO_1156 (O_1156,N_8786,N_8785);
nor UO_1157 (O_1157,N_7314,N_5260);
and UO_1158 (O_1158,N_5382,N_7633);
and UO_1159 (O_1159,N_7980,N_5826);
and UO_1160 (O_1160,N_6993,N_7913);
or UO_1161 (O_1161,N_9707,N_7428);
nand UO_1162 (O_1162,N_8970,N_5094);
or UO_1163 (O_1163,N_5170,N_6400);
nor UO_1164 (O_1164,N_8679,N_5553);
nor UO_1165 (O_1165,N_6284,N_8790);
nor UO_1166 (O_1166,N_6010,N_9696);
and UO_1167 (O_1167,N_9290,N_9803);
and UO_1168 (O_1168,N_6910,N_7786);
xor UO_1169 (O_1169,N_6572,N_9597);
or UO_1170 (O_1170,N_6115,N_6676);
or UO_1171 (O_1171,N_6850,N_6480);
nand UO_1172 (O_1172,N_5496,N_6730);
and UO_1173 (O_1173,N_5434,N_5715);
and UO_1174 (O_1174,N_5862,N_8230);
or UO_1175 (O_1175,N_6853,N_9136);
nor UO_1176 (O_1176,N_5206,N_5545);
nand UO_1177 (O_1177,N_8883,N_7093);
nand UO_1178 (O_1178,N_8172,N_9428);
or UO_1179 (O_1179,N_5983,N_8581);
nand UO_1180 (O_1180,N_7351,N_5952);
and UO_1181 (O_1181,N_9626,N_7227);
and UO_1182 (O_1182,N_5365,N_6880);
nor UO_1183 (O_1183,N_8351,N_6754);
xnor UO_1184 (O_1184,N_6817,N_5776);
and UO_1185 (O_1185,N_5760,N_8234);
or UO_1186 (O_1186,N_8204,N_8133);
and UO_1187 (O_1187,N_9571,N_7359);
or UO_1188 (O_1188,N_7822,N_5083);
nand UO_1189 (O_1189,N_5874,N_8214);
and UO_1190 (O_1190,N_5607,N_9307);
or UO_1191 (O_1191,N_9839,N_9958);
nand UO_1192 (O_1192,N_5592,N_6893);
and UO_1193 (O_1193,N_8265,N_5021);
nor UO_1194 (O_1194,N_7910,N_8450);
xor UO_1195 (O_1195,N_6740,N_9501);
or UO_1196 (O_1196,N_8050,N_7675);
nor UO_1197 (O_1197,N_6090,N_6373);
and UO_1198 (O_1198,N_8476,N_6561);
xor UO_1199 (O_1199,N_5256,N_8623);
or UO_1200 (O_1200,N_8062,N_6395);
nand UO_1201 (O_1201,N_7216,N_9409);
and UO_1202 (O_1202,N_5827,N_6838);
nand UO_1203 (O_1203,N_9005,N_9347);
nor UO_1204 (O_1204,N_9196,N_7713);
nor UO_1205 (O_1205,N_7846,N_5487);
and UO_1206 (O_1206,N_8865,N_7409);
xor UO_1207 (O_1207,N_8445,N_8074);
or UO_1208 (O_1208,N_6333,N_5397);
or UO_1209 (O_1209,N_7741,N_5007);
and UO_1210 (O_1210,N_7858,N_6694);
or UO_1211 (O_1211,N_6309,N_9077);
nor UO_1212 (O_1212,N_6254,N_5398);
or UO_1213 (O_1213,N_9481,N_5072);
nand UO_1214 (O_1214,N_5159,N_5644);
and UO_1215 (O_1215,N_8285,N_7169);
nor UO_1216 (O_1216,N_6051,N_5217);
or UO_1217 (O_1217,N_9497,N_7662);
nor UO_1218 (O_1218,N_7170,N_7185);
or UO_1219 (O_1219,N_6454,N_6750);
nor UO_1220 (O_1220,N_8945,N_7809);
nor UO_1221 (O_1221,N_9986,N_8933);
and UO_1222 (O_1222,N_8400,N_8569);
or UO_1223 (O_1223,N_7352,N_6389);
nor UO_1224 (O_1224,N_6458,N_7859);
or UO_1225 (O_1225,N_7228,N_6420);
nand UO_1226 (O_1226,N_8905,N_9640);
nor UO_1227 (O_1227,N_6498,N_8982);
or UO_1228 (O_1228,N_5762,N_6453);
or UO_1229 (O_1229,N_6407,N_6883);
or UO_1230 (O_1230,N_8690,N_5736);
nor UO_1231 (O_1231,N_7401,N_9379);
and UO_1232 (O_1232,N_7578,N_6021);
nand UO_1233 (O_1233,N_9740,N_7557);
nor UO_1234 (O_1234,N_5112,N_9811);
nor UO_1235 (O_1235,N_7742,N_5150);
or UO_1236 (O_1236,N_6490,N_9567);
xnor UO_1237 (O_1237,N_6766,N_7550);
and UO_1238 (O_1238,N_8555,N_5865);
nor UO_1239 (O_1239,N_5141,N_9198);
and UO_1240 (O_1240,N_9017,N_7823);
xor UO_1241 (O_1241,N_6678,N_7667);
or UO_1242 (O_1242,N_6536,N_7489);
nor UO_1243 (O_1243,N_6293,N_7700);
or UO_1244 (O_1244,N_9507,N_8385);
nor UO_1245 (O_1245,N_8235,N_5685);
or UO_1246 (O_1246,N_5821,N_8964);
or UO_1247 (O_1247,N_9840,N_8994);
nand UO_1248 (O_1248,N_6060,N_8929);
nand UO_1249 (O_1249,N_8975,N_6394);
nor UO_1250 (O_1250,N_7681,N_7939);
nand UO_1251 (O_1251,N_9966,N_6938);
nand UO_1252 (O_1252,N_7164,N_7197);
and UO_1253 (O_1253,N_6409,N_6673);
nor UO_1254 (O_1254,N_8184,N_9800);
and UO_1255 (O_1255,N_5953,N_9529);
nand UO_1256 (O_1256,N_6857,N_9244);
and UO_1257 (O_1257,N_7710,N_6864);
or UO_1258 (O_1258,N_8479,N_6032);
nand UO_1259 (O_1259,N_5703,N_7321);
and UO_1260 (O_1260,N_6709,N_6065);
and UO_1261 (O_1261,N_5469,N_8259);
nand UO_1262 (O_1262,N_5008,N_7469);
nor UO_1263 (O_1263,N_6112,N_7142);
and UO_1264 (O_1264,N_8061,N_9145);
nand UO_1265 (O_1265,N_5492,N_7620);
nor UO_1266 (O_1266,N_5544,N_6157);
or UO_1267 (O_1267,N_5734,N_8349);
or UO_1268 (O_1268,N_6287,N_7512);
nor UO_1269 (O_1269,N_7816,N_6765);
nand UO_1270 (O_1270,N_7391,N_6759);
nand UO_1271 (O_1271,N_7066,N_7908);
nand UO_1272 (O_1272,N_7269,N_6775);
nor UO_1273 (O_1273,N_6356,N_6903);
nand UO_1274 (O_1274,N_8787,N_6793);
nor UO_1275 (O_1275,N_9360,N_6412);
nand UO_1276 (O_1276,N_6092,N_9774);
nor UO_1277 (O_1277,N_8331,N_5078);
nor UO_1278 (O_1278,N_5716,N_9302);
and UO_1279 (O_1279,N_6586,N_5423);
or UO_1280 (O_1280,N_5689,N_6672);
nor UO_1281 (O_1281,N_9028,N_8523);
nor UO_1282 (O_1282,N_5905,N_7705);
and UO_1283 (O_1283,N_8788,N_5164);
and UO_1284 (O_1284,N_8800,N_7296);
nor UO_1285 (O_1285,N_8572,N_7963);
and UO_1286 (O_1286,N_9655,N_9058);
nand UO_1287 (O_1287,N_6667,N_7153);
nor UO_1288 (O_1288,N_7886,N_8819);
or UO_1289 (O_1289,N_7207,N_8488);
nor UO_1290 (O_1290,N_7832,N_9649);
nand UO_1291 (O_1291,N_7287,N_6855);
or UO_1292 (O_1292,N_9793,N_5711);
or UO_1293 (O_1293,N_6037,N_9112);
nand UO_1294 (O_1294,N_5191,N_6175);
nand UO_1295 (O_1295,N_8482,N_9680);
or UO_1296 (O_1296,N_8802,N_7330);
and UO_1297 (O_1297,N_9807,N_8059);
and UO_1298 (O_1298,N_8071,N_8617);
nor UO_1299 (O_1299,N_6022,N_8166);
or UO_1300 (O_1300,N_6369,N_9186);
xor UO_1301 (O_1301,N_5209,N_8144);
or UO_1302 (O_1302,N_7073,N_5977);
nor UO_1303 (O_1303,N_9766,N_8408);
and UO_1304 (O_1304,N_7728,N_7824);
nor UO_1305 (O_1305,N_9603,N_5467);
or UO_1306 (O_1306,N_7616,N_5240);
nand UO_1307 (O_1307,N_7083,N_7006);
or UO_1308 (O_1308,N_8188,N_9141);
nand UO_1309 (O_1309,N_7088,N_7172);
nor UO_1310 (O_1310,N_9467,N_5663);
or UO_1311 (O_1311,N_8876,N_5331);
nor UO_1312 (O_1312,N_8086,N_8740);
and UO_1313 (O_1313,N_8734,N_6984);
nand UO_1314 (O_1314,N_9286,N_9708);
or UO_1315 (O_1315,N_6745,N_7748);
nand UO_1316 (O_1316,N_5115,N_7418);
nor UO_1317 (O_1317,N_8578,N_9779);
nor UO_1318 (O_1318,N_9804,N_8100);
or UO_1319 (O_1319,N_5590,N_9764);
nor UO_1320 (O_1320,N_6895,N_5554);
nand UO_1321 (O_1321,N_9316,N_8291);
nand UO_1322 (O_1322,N_9954,N_6142);
xnor UO_1323 (O_1323,N_7796,N_5618);
or UO_1324 (O_1324,N_8743,N_9831);
nand UO_1325 (O_1325,N_5250,N_8725);
and UO_1326 (O_1326,N_7413,N_6135);
and UO_1327 (O_1327,N_9252,N_6167);
or UO_1328 (O_1328,N_7771,N_9129);
or UO_1329 (O_1329,N_5006,N_7327);
nand UO_1330 (O_1330,N_7802,N_5483);
and UO_1331 (O_1331,N_5389,N_9629);
or UO_1332 (O_1332,N_6324,N_8139);
nand UO_1333 (O_1333,N_9348,N_8048);
nand UO_1334 (O_1334,N_9006,N_9882);
nor UO_1335 (O_1335,N_7168,N_9320);
and UO_1336 (O_1336,N_9910,N_6585);
nand UO_1337 (O_1337,N_8748,N_5597);
and UO_1338 (O_1338,N_6248,N_9762);
nand UO_1339 (O_1339,N_5074,N_9837);
and UO_1340 (O_1340,N_7569,N_6330);
nor UO_1341 (O_1341,N_7156,N_8709);
nor UO_1342 (O_1342,N_5129,N_9439);
nor UO_1343 (O_1343,N_8766,N_7237);
and UO_1344 (O_1344,N_6312,N_7936);
nor UO_1345 (O_1345,N_5133,N_9331);
and UO_1346 (O_1346,N_5413,N_8717);
or UO_1347 (O_1347,N_5745,N_9712);
and UO_1348 (O_1348,N_6976,N_8729);
nand UO_1349 (O_1349,N_5172,N_7825);
nor UO_1350 (O_1350,N_7338,N_8015);
or UO_1351 (O_1351,N_5583,N_7646);
nand UO_1352 (O_1352,N_7459,N_9114);
or UO_1353 (O_1353,N_9969,N_5988);
and UO_1354 (O_1354,N_7157,N_8457);
nor UO_1355 (O_1355,N_6681,N_5375);
nand UO_1356 (O_1356,N_8312,N_8158);
or UO_1357 (O_1357,N_6408,N_7831);
nor UO_1358 (O_1358,N_7089,N_8072);
or UO_1359 (O_1359,N_5388,N_5872);
nor UO_1360 (O_1360,N_6757,N_6431);
nor UO_1361 (O_1361,N_6371,N_8947);
nor UO_1362 (O_1362,N_7996,N_6712);
and UO_1363 (O_1363,N_7549,N_6643);
and UO_1364 (O_1364,N_5368,N_9052);
and UO_1365 (O_1365,N_7548,N_8575);
nand UO_1366 (O_1366,N_8220,N_7526);
xor UO_1367 (O_1367,N_5604,N_9525);
or UO_1368 (O_1368,N_8655,N_7706);
and UO_1369 (O_1369,N_7387,N_8686);
nor UO_1370 (O_1370,N_8840,N_9049);
xor UO_1371 (O_1371,N_6906,N_7722);
and UO_1372 (O_1372,N_5155,N_7556);
nand UO_1373 (O_1373,N_6308,N_7432);
and UO_1374 (O_1374,N_5771,N_9297);
or UO_1375 (O_1375,N_8129,N_6234);
or UO_1376 (O_1376,N_6567,N_5887);
or UO_1377 (O_1377,N_9918,N_7131);
and UO_1378 (O_1378,N_5929,N_8340);
and UO_1379 (O_1379,N_8307,N_7480);
and UO_1380 (O_1380,N_8273,N_9042);
nand UO_1381 (O_1381,N_9038,N_5216);
nor UO_1382 (O_1382,N_8837,N_6213);
and UO_1383 (O_1383,N_7554,N_5940);
or UO_1384 (O_1384,N_7882,N_9545);
xor UO_1385 (O_1385,N_8502,N_5611);
nand UO_1386 (O_1386,N_7668,N_5394);
or UO_1387 (O_1387,N_7097,N_5809);
or UO_1388 (O_1388,N_5452,N_7522);
or UO_1389 (O_1389,N_6346,N_9444);
or UO_1390 (O_1390,N_8950,N_6685);
or UO_1391 (O_1391,N_6134,N_9912);
or UO_1392 (O_1392,N_8152,N_9326);
and UO_1393 (O_1393,N_6509,N_8275);
or UO_1394 (O_1394,N_9530,N_5244);
nor UO_1395 (O_1395,N_9994,N_5363);
nor UO_1396 (O_1396,N_8417,N_9948);
nor UO_1397 (O_1397,N_8405,N_7950);
and UO_1398 (O_1398,N_6723,N_6455);
and UO_1399 (O_1399,N_6739,N_8401);
and UO_1400 (O_1400,N_5399,N_7058);
or UO_1401 (O_1401,N_9660,N_5660);
and UO_1402 (O_1402,N_6491,N_6591);
and UO_1403 (O_1403,N_6285,N_9642);
and UO_1404 (O_1404,N_7747,N_7623);
nand UO_1405 (O_1405,N_7160,N_8777);
nor UO_1406 (O_1406,N_5151,N_5223);
nand UO_1407 (O_1407,N_5005,N_6638);
or UO_1408 (O_1408,N_7577,N_5812);
and UO_1409 (O_1409,N_5338,N_8054);
or UO_1410 (O_1410,N_5348,N_8288);
nand UO_1411 (O_1411,N_8346,N_7305);
nand UO_1412 (O_1412,N_8258,N_5345);
nand UO_1413 (O_1413,N_8200,N_6515);
nand UO_1414 (O_1414,N_9677,N_9661);
or UO_1415 (O_1415,N_9208,N_6751);
nor UO_1416 (O_1416,N_7727,N_9721);
xnor UO_1417 (O_1417,N_8057,N_9482);
nand UO_1418 (O_1418,N_9287,N_8886);
nand UO_1419 (O_1419,N_6139,N_5897);
or UO_1420 (O_1420,N_7206,N_7087);
nor UO_1421 (O_1421,N_8911,N_6088);
or UO_1422 (O_1422,N_9922,N_5758);
nand UO_1423 (O_1423,N_7152,N_5063);
or UO_1424 (O_1424,N_5102,N_5700);
nand UO_1425 (O_1425,N_8027,N_6798);
nor UO_1426 (O_1426,N_9747,N_9532);
xnor UO_1427 (O_1427,N_6262,N_6271);
nand UO_1428 (O_1428,N_8591,N_5710);
or UO_1429 (O_1429,N_7277,N_7509);
nand UO_1430 (O_1430,N_9620,N_7531);
or UO_1431 (O_1431,N_5574,N_7716);
and UO_1432 (O_1432,N_9267,N_6171);
nand UO_1433 (O_1433,N_7587,N_8904);
and UO_1434 (O_1434,N_7028,N_6126);
nor UO_1435 (O_1435,N_9874,N_9138);
or UO_1436 (O_1436,N_6579,N_9309);
and UO_1437 (O_1437,N_9396,N_7483);
nand UO_1438 (O_1438,N_7178,N_6518);
nor UO_1439 (O_1439,N_7342,N_6557);
and UO_1440 (O_1440,N_5121,N_5127);
and UO_1441 (O_1441,N_5490,N_5774);
and UO_1442 (O_1442,N_6587,N_7691);
nand UO_1443 (O_1443,N_7104,N_7534);
xor UO_1444 (O_1444,N_9008,N_5093);
or UO_1445 (O_1445,N_5817,N_6039);
nand UO_1446 (O_1446,N_7487,N_7496);
and UO_1447 (O_1447,N_9415,N_9180);
nor UO_1448 (O_1448,N_5304,N_6140);
nand UO_1449 (O_1449,N_9899,N_5269);
xor UO_1450 (O_1450,N_8605,N_5158);
or UO_1451 (O_1451,N_6744,N_6208);
xor UO_1452 (O_1452,N_6920,N_5044);
nor UO_1453 (O_1453,N_6958,N_9031);
nor UO_1454 (O_1454,N_9483,N_8811);
and UO_1455 (O_1455,N_7276,N_5666);
or UO_1456 (O_1456,N_8499,N_6632);
xnor UO_1457 (O_1457,N_7905,N_6990);
nand UO_1458 (O_1458,N_9605,N_7171);
nor UO_1459 (O_1459,N_7921,N_6085);
and UO_1460 (O_1460,N_5049,N_5284);
nor UO_1461 (O_1461,N_6623,N_6905);
and UO_1462 (O_1462,N_7923,N_7473);
nand UO_1463 (O_1463,N_6155,N_9088);
nor UO_1464 (O_1464,N_8407,N_7478);
nor UO_1465 (O_1465,N_6803,N_6720);
nor UO_1466 (O_1466,N_9065,N_5227);
or UO_1467 (O_1467,N_5426,N_7431);
nor UO_1468 (O_1468,N_8817,N_9513);
xnor UO_1469 (O_1469,N_6692,N_9627);
nand UO_1470 (O_1470,N_5984,N_6865);
nor UO_1471 (O_1471,N_6268,N_6233);
or UO_1472 (O_1472,N_9616,N_6292);
and UO_1473 (O_1473,N_8279,N_5814);
or UO_1474 (O_1474,N_5418,N_6922);
and UO_1475 (O_1475,N_8996,N_6942);
nor UO_1476 (O_1476,N_9709,N_7632);
nand UO_1477 (O_1477,N_9554,N_6114);
nor UO_1478 (O_1478,N_5404,N_8241);
nand UO_1479 (O_1479,N_6365,N_8551);
and UO_1480 (O_1480,N_7682,N_6777);
nand UO_1481 (O_1481,N_8579,N_6921);
or UO_1482 (O_1482,N_7866,N_7684);
nor UO_1483 (O_1483,N_9935,N_8306);
or UO_1484 (O_1484,N_7648,N_6629);
nand UO_1485 (O_1485,N_9495,N_9596);
and UO_1486 (O_1486,N_7379,N_7737);
and UO_1487 (O_1487,N_6000,N_5765);
or UO_1488 (O_1488,N_5152,N_9844);
nor UO_1489 (O_1489,N_7943,N_6582);
nand UO_1490 (O_1490,N_8799,N_5366);
and UO_1491 (O_1491,N_8397,N_6081);
and UO_1492 (O_1492,N_5481,N_7707);
and UO_1493 (O_1493,N_7027,N_9933);
nor UO_1494 (O_1494,N_7053,N_7694);
or UO_1495 (O_1495,N_9606,N_6566);
nand UO_1496 (O_1496,N_7438,N_8829);
xor UO_1497 (O_1497,N_6482,N_7797);
or UO_1498 (O_1498,N_9775,N_7212);
nor UO_1499 (O_1499,N_8333,N_9848);
endmodule