module basic_1500_15000_2000_30_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_1287,In_51);
and U1 (N_1,In_1470,In_740);
and U2 (N_2,In_1085,In_441);
or U3 (N_3,In_1091,In_1102);
and U4 (N_4,In_1194,In_1113);
nor U5 (N_5,In_1486,In_775);
xor U6 (N_6,In_144,In_449);
or U7 (N_7,In_721,In_40);
and U8 (N_8,In_1433,In_102);
or U9 (N_9,In_1259,In_1483);
xnor U10 (N_10,In_141,In_1369);
nand U11 (N_11,In_1067,In_1362);
or U12 (N_12,In_1344,In_112);
nor U13 (N_13,In_750,In_717);
nor U14 (N_14,In_1318,In_1214);
nand U15 (N_15,In_1295,In_382);
nor U16 (N_16,In_611,In_123);
nor U17 (N_17,In_1336,In_938);
nor U18 (N_18,In_781,In_1345);
and U19 (N_19,In_1276,In_972);
and U20 (N_20,In_1078,In_1041);
nand U21 (N_21,In_981,In_1261);
or U22 (N_22,In_1268,In_1203);
nor U23 (N_23,In_1210,In_347);
nand U24 (N_24,In_1456,In_764);
nor U25 (N_25,In_1332,In_193);
nand U26 (N_26,In_660,In_281);
and U27 (N_27,In_1071,In_1328);
or U28 (N_28,In_591,In_617);
and U29 (N_29,In_706,In_957);
xnor U30 (N_30,In_1263,In_1052);
nor U31 (N_31,In_709,In_1152);
nand U32 (N_32,In_110,In_979);
and U33 (N_33,In_215,In_970);
or U34 (N_34,In_213,In_44);
or U35 (N_35,In_854,In_1428);
or U36 (N_36,In_1015,In_465);
nor U37 (N_37,In_707,In_731);
nor U38 (N_38,In_331,In_900);
nor U39 (N_39,In_204,In_759);
and U40 (N_40,In_700,In_958);
or U41 (N_41,In_104,In_401);
nand U42 (N_42,In_229,In_198);
and U43 (N_43,In_910,In_1283);
nor U44 (N_44,In_101,In_1384);
and U45 (N_45,In_870,In_120);
nor U46 (N_46,In_127,In_969);
and U47 (N_47,In_1448,In_306);
nor U48 (N_48,In_724,In_35);
nor U49 (N_49,In_1151,In_962);
nand U50 (N_50,In_1192,In_921);
nand U51 (N_51,In_472,In_289);
nor U52 (N_52,In_641,In_129);
or U53 (N_53,In_809,In_584);
or U54 (N_54,In_409,In_948);
and U55 (N_55,In_837,In_564);
or U56 (N_56,In_657,In_742);
nand U57 (N_57,In_462,In_1434);
xor U58 (N_58,In_173,In_250);
and U59 (N_59,In_615,In_178);
xor U60 (N_60,In_1045,In_1414);
nand U61 (N_61,In_1218,In_1378);
or U62 (N_62,In_538,In_304);
or U63 (N_63,In_366,In_1451);
nor U64 (N_64,In_1491,In_1458);
and U65 (N_65,In_1084,In_315);
nor U66 (N_66,In_1230,In_240);
and U67 (N_67,In_819,In_1300);
nor U68 (N_68,In_161,In_1278);
nand U69 (N_69,In_165,In_589);
xnor U70 (N_70,In_1440,In_406);
xor U71 (N_71,In_961,In_1396);
xnor U72 (N_72,In_222,In_671);
nor U73 (N_73,In_1316,In_1247);
nand U74 (N_74,In_761,In_29);
nand U75 (N_75,In_41,In_397);
nand U76 (N_76,In_982,In_206);
nand U77 (N_77,In_1020,In_359);
xnor U78 (N_78,In_174,In_540);
nor U79 (N_79,In_189,In_15);
nor U80 (N_80,In_1213,In_105);
nand U81 (N_81,In_664,In_587);
nand U82 (N_82,In_1235,In_708);
nand U83 (N_83,In_182,In_1099);
nor U84 (N_84,In_183,In_220);
nand U85 (N_85,In_224,In_282);
and U86 (N_86,In_603,In_1000);
or U87 (N_87,In_755,In_1055);
or U88 (N_88,In_1157,In_468);
or U89 (N_89,In_1399,In_687);
or U90 (N_90,In_385,In_872);
and U91 (N_91,In_896,In_9);
nor U92 (N_92,In_1307,In_945);
nor U93 (N_93,In_115,In_158);
nor U94 (N_94,In_318,In_484);
or U95 (N_95,In_210,In_1205);
nor U96 (N_96,In_694,In_489);
or U97 (N_97,In_799,In_196);
and U98 (N_98,In_705,In_551);
nand U99 (N_99,In_1086,In_455);
nor U100 (N_100,In_97,In_175);
or U101 (N_101,In_787,In_762);
nand U102 (N_102,In_856,In_776);
nand U103 (N_103,In_1212,In_454);
nor U104 (N_104,In_784,In_121);
nand U105 (N_105,In_581,In_1266);
nor U106 (N_106,In_1221,In_574);
nor U107 (N_107,In_453,In_1273);
or U108 (N_108,In_1348,In_990);
nor U109 (N_109,In_770,In_1056);
or U110 (N_110,In_1473,In_283);
nor U111 (N_111,In_782,In_107);
and U112 (N_112,In_502,In_446);
nor U113 (N_113,In_1068,In_1076);
or U114 (N_114,In_1206,In_667);
nand U115 (N_115,In_866,In_813);
or U116 (N_116,In_6,In_871);
and U117 (N_117,In_350,In_1027);
and U118 (N_118,In_602,In_1393);
nor U119 (N_119,In_1016,In_783);
nand U120 (N_120,In_1379,In_555);
and U121 (N_121,In_874,In_1431);
or U122 (N_122,In_275,In_216);
nand U123 (N_123,In_1341,In_968);
or U124 (N_124,In_648,In_1453);
or U125 (N_125,In_113,In_909);
or U126 (N_126,In_954,In_485);
xnor U127 (N_127,In_1038,In_1329);
xnor U128 (N_128,In_767,In_225);
nand U129 (N_129,In_915,In_1357);
and U130 (N_130,In_1166,In_195);
or U131 (N_131,In_342,In_133);
or U132 (N_132,In_356,In_1251);
nand U133 (N_133,In_839,In_636);
and U134 (N_134,In_821,In_1331);
nand U135 (N_135,In_980,In_207);
nor U136 (N_136,In_199,In_1153);
and U137 (N_137,In_337,In_605);
xnor U138 (N_138,In_1498,In_522);
and U139 (N_139,In_1360,In_1043);
and U140 (N_140,In_124,In_728);
and U141 (N_141,In_596,In_375);
nand U142 (N_142,In_1255,In_1190);
nand U143 (N_143,In_24,In_678);
or U144 (N_144,In_1388,In_1444);
nand U145 (N_145,In_52,In_333);
nand U146 (N_146,In_528,In_1479);
and U147 (N_147,In_310,In_53);
and U148 (N_148,In_801,In_162);
nand U149 (N_149,In_1065,In_467);
or U150 (N_150,In_1439,In_1062);
nand U151 (N_151,In_341,In_883);
and U152 (N_152,In_773,In_736);
nand U153 (N_153,In_274,In_533);
nand U154 (N_154,In_1219,In_1415);
and U155 (N_155,In_499,In_1304);
nor U156 (N_156,In_438,In_1105);
xor U157 (N_157,In_459,In_765);
and U158 (N_158,In_1243,In_1495);
nand U159 (N_159,In_280,In_1058);
xnor U160 (N_160,In_261,In_332);
xor U161 (N_161,In_1004,In_245);
xnor U162 (N_162,In_1216,In_862);
nor U163 (N_163,In_246,In_1042);
and U164 (N_164,In_547,In_1367);
and U165 (N_165,In_685,In_640);
xnor U166 (N_166,In_1392,In_91);
and U167 (N_167,In_748,In_497);
xor U168 (N_168,In_699,In_228);
nor U169 (N_169,In_190,In_418);
and U170 (N_170,In_532,In_1013);
and U171 (N_171,In_975,In_1007);
xor U172 (N_172,In_932,In_1237);
or U173 (N_173,In_188,In_1233);
or U174 (N_174,In_13,In_955);
nor U175 (N_175,In_1461,In_384);
and U176 (N_176,In_1211,In_797);
and U177 (N_177,In_264,In_1073);
nor U178 (N_178,In_435,In_570);
nor U179 (N_179,In_343,In_481);
and U180 (N_180,In_417,In_396);
and U181 (N_181,In_1236,In_427);
nand U182 (N_182,In_208,In_1409);
or U183 (N_183,In_328,In_634);
and U184 (N_184,In_130,In_1454);
nor U185 (N_185,In_1140,In_70);
nor U186 (N_186,In_1093,In_1269);
and U187 (N_187,In_17,In_828);
nand U188 (N_188,In_747,In_1437);
nor U189 (N_189,In_415,In_746);
nand U190 (N_190,In_1292,In_279);
or U191 (N_191,In_30,In_233);
xor U192 (N_192,In_1034,In_1108);
or U193 (N_193,In_1189,In_953);
and U194 (N_194,In_307,In_639);
or U195 (N_195,In_913,In_345);
nor U196 (N_196,In_1466,In_692);
or U197 (N_197,In_774,In_718);
or U198 (N_198,In_623,In_824);
and U199 (N_199,In_749,In_1156);
nand U200 (N_200,In_544,In_231);
nor U201 (N_201,In_22,In_769);
or U202 (N_202,In_847,In_1005);
or U203 (N_203,In_924,In_381);
nor U204 (N_204,In_1204,In_536);
nand U205 (N_205,In_296,In_100);
nor U206 (N_206,In_1137,In_1480);
and U207 (N_207,In_256,In_11);
nand U208 (N_208,In_440,In_569);
nand U209 (N_209,In_807,In_1423);
xnor U210 (N_210,In_1089,In_1303);
nor U211 (N_211,In_1312,In_727);
nand U212 (N_212,In_393,In_1449);
nor U213 (N_213,In_391,In_10);
nand U214 (N_214,In_1010,In_443);
and U215 (N_215,In_1198,In_1242);
or U216 (N_216,In_34,In_83);
xnor U217 (N_217,In_644,In_94);
nand U218 (N_218,In_1253,In_633);
or U219 (N_219,In_157,In_716);
nand U220 (N_220,In_822,In_21);
nor U221 (N_221,In_1310,In_357);
or U222 (N_222,In_1353,In_730);
or U223 (N_223,In_670,In_223);
or U224 (N_224,In_1298,In_802);
or U225 (N_225,In_88,In_1179);
nand U226 (N_226,In_812,In_1280);
and U227 (N_227,In_1185,In_1375);
or U228 (N_228,In_428,In_579);
xnor U229 (N_229,In_803,In_1144);
nand U230 (N_230,In_491,In_624);
nor U231 (N_231,In_1200,In_1047);
or U232 (N_232,In_542,In_493);
xor U233 (N_233,In_646,In_608);
and U234 (N_234,In_1446,In_928);
nor U235 (N_235,In_1199,In_416);
nor U236 (N_236,In_1313,In_136);
or U237 (N_237,In_790,In_726);
or U238 (N_238,In_666,In_563);
or U239 (N_239,In_853,In_202);
or U240 (N_240,In_875,In_1069);
nor U241 (N_241,In_1305,In_1122);
xor U242 (N_242,In_956,In_404);
and U243 (N_243,In_218,In_1469);
nand U244 (N_244,In_876,In_777);
nor U245 (N_245,In_1290,In_934);
xor U246 (N_246,In_595,In_1141);
nor U247 (N_247,In_1077,In_425);
and U248 (N_248,In_805,In_93);
nor U249 (N_249,In_1459,In_926);
and U250 (N_250,In_169,In_612);
nand U251 (N_251,In_1408,In_126);
and U252 (N_252,In_475,In_1035);
nand U253 (N_253,In_663,In_1462);
xor U254 (N_254,In_508,In_65);
nor U255 (N_255,In_92,In_56);
nand U256 (N_256,In_1254,In_1249);
and U257 (N_257,In_1308,In_1285);
nand U258 (N_258,In_498,In_792);
and U259 (N_259,In_861,In_495);
nand U260 (N_260,In_545,In_1334);
and U261 (N_261,In_1180,In_78);
nand U262 (N_262,In_1402,In_673);
and U263 (N_263,In_241,In_576);
and U264 (N_264,In_1394,In_1382);
xor U265 (N_265,In_1342,In_374);
nor U266 (N_266,In_850,In_482);
and U267 (N_267,In_548,In_851);
and U268 (N_268,In_899,In_490);
nor U269 (N_269,In_539,In_890);
nand U270 (N_270,In_60,In_621);
nand U271 (N_271,In_808,In_1244);
nor U272 (N_272,In_451,In_118);
nand U273 (N_273,In_1164,In_1315);
xor U274 (N_274,In_998,In_598);
and U275 (N_275,In_373,In_303);
or U276 (N_276,In_1471,In_146);
nand U277 (N_277,In_1499,In_1172);
nor U278 (N_278,In_630,In_983);
or U279 (N_279,In_1049,In_1054);
xnor U280 (N_280,In_1355,In_1258);
xnor U281 (N_281,In_1340,In_1381);
xor U282 (N_282,In_1317,In_448);
and U283 (N_283,In_849,In_186);
and U284 (N_284,In_58,In_450);
nand U285 (N_285,In_886,In_479);
nor U286 (N_286,In_785,In_679);
nor U287 (N_287,In_1059,In_511);
or U288 (N_288,In_321,In_680);
or U289 (N_289,In_1188,In_902);
and U290 (N_290,In_1358,In_1051);
nor U291 (N_291,In_949,In_713);
or U292 (N_292,In_159,In_487);
nor U293 (N_293,In_71,In_607);
nor U294 (N_294,In_738,In_1492);
nand U295 (N_295,In_818,In_500);
and U296 (N_296,In_372,In_1149);
or U297 (N_297,In_629,In_69);
and U298 (N_298,In_325,In_554);
nor U299 (N_299,In_437,In_1125);
nor U300 (N_300,In_846,In_59);
and U301 (N_301,In_923,In_606);
and U302 (N_302,In_952,In_863);
and U303 (N_303,In_1238,In_230);
nor U304 (N_304,In_838,In_73);
nand U305 (N_305,In_388,In_297);
nand U306 (N_306,In_741,In_269);
and U307 (N_307,In_1174,In_151);
or U308 (N_308,In_831,In_1006);
nor U309 (N_309,In_284,In_1159);
xor U310 (N_310,In_804,In_867);
and U311 (N_311,In_662,In_585);
nand U312 (N_312,In_1252,In_334);
and U313 (N_313,In_766,In_571);
or U314 (N_314,In_1335,In_1240);
nor U315 (N_315,In_816,In_649);
or U316 (N_316,In_160,In_676);
nor U317 (N_317,In_1496,In_757);
and U318 (N_318,In_527,In_798);
or U319 (N_319,In_1264,In_558);
and U320 (N_320,In_413,In_843);
and U321 (N_321,In_888,In_1012);
nand U322 (N_322,In_939,In_211);
nor U323 (N_323,In_55,In_918);
nand U324 (N_324,In_23,In_1484);
nand U325 (N_325,In_908,In_1142);
nand U326 (N_326,In_1103,In_1028);
or U327 (N_327,In_780,In_677);
and U328 (N_328,In_895,In_743);
nor U329 (N_329,In_1031,In_753);
nand U330 (N_330,In_442,In_674);
xnor U331 (N_331,In_826,In_423);
nor U332 (N_332,In_457,In_978);
xor U333 (N_333,In_286,In_627);
nand U334 (N_334,In_609,In_299);
nor U335 (N_335,In_1025,In_496);
or U336 (N_336,In_1468,In_1146);
nor U337 (N_337,In_1272,In_1082);
and U338 (N_338,In_267,In_655);
nand U339 (N_339,In_559,In_535);
or U340 (N_340,In_894,In_255);
or U341 (N_341,In_1044,In_922);
or U342 (N_342,In_349,In_1048);
nand U343 (N_343,In_72,In_31);
or U344 (N_344,In_252,In_1323);
xor U345 (N_345,In_1350,In_1410);
nor U346 (N_346,In_1148,In_1380);
nand U347 (N_347,In_710,In_265);
xor U348 (N_348,In_568,In_594);
xnor U349 (N_349,In_877,In_150);
nand U350 (N_350,In_905,In_32);
nor U351 (N_351,In_562,In_752);
nor U352 (N_352,In_1270,In_278);
or U353 (N_353,In_1139,In_197);
and U354 (N_354,In_1135,In_232);
nor U355 (N_355,In_238,In_1118);
and U356 (N_356,In_26,In_897);
nor U357 (N_357,In_313,In_1222);
and U358 (N_358,In_293,In_965);
nor U359 (N_359,In_1452,In_567);
xor U360 (N_360,In_1248,In_789);
nor U361 (N_361,In_469,In_37);
and U362 (N_362,In_825,In_1101);
or U363 (N_363,In_1296,In_645);
nor U364 (N_364,In_263,In_48);
nor U365 (N_365,In_504,In_301);
xnor U366 (N_366,In_49,In_1387);
nor U367 (N_367,In_669,In_1134);
and U368 (N_368,In_57,In_1224);
nand U369 (N_369,In_758,In_546);
nor U370 (N_370,In_109,In_191);
nor U371 (N_371,In_458,In_378);
nor U372 (N_372,In_362,In_1079);
nor U373 (N_373,In_1053,In_290);
nor U374 (N_374,In_842,In_27);
nor U375 (N_375,In_268,In_419);
or U376 (N_376,In_103,In_407);
nand U377 (N_377,In_1106,In_1225);
nor U378 (N_378,In_702,In_737);
and U379 (N_379,In_1162,In_788);
and U380 (N_380,In_712,In_541);
xnor U381 (N_381,In_778,In_1168);
nor U382 (N_382,In_722,In_181);
nand U383 (N_383,In_1386,In_1314);
xnor U384 (N_384,In_1309,In_1021);
nor U385 (N_385,In_1330,In_1002);
and U386 (N_386,In_1397,In_1165);
and U387 (N_387,In_898,In_474);
or U388 (N_388,In_90,In_1060);
or U389 (N_389,In_486,In_725);
nand U390 (N_390,In_1075,In_1464);
or U391 (N_391,In_148,In_128);
xnor U392 (N_392,In_360,In_620);
nor U393 (N_393,In_1293,In_324);
nand U394 (N_394,In_1363,In_1435);
nor U395 (N_395,In_1232,In_106);
nand U396 (N_396,In_1032,In_1297);
xor U397 (N_397,In_668,In_889);
nand U398 (N_398,In_477,In_1193);
and U399 (N_399,In_1327,In_947);
xor U400 (N_400,In_1081,In_887);
and U401 (N_401,In_33,In_260);
nor U402 (N_402,In_833,In_517);
and U403 (N_403,In_935,In_1361);
nor U404 (N_404,In_1119,In_583);
nor U405 (N_405,In_1346,In_763);
and U406 (N_406,In_1337,In_434);
or U407 (N_407,In_1390,In_857);
xnor U408 (N_408,In_116,In_410);
nand U409 (N_409,In_1282,In_933);
nor U410 (N_410,In_85,In_560);
nand U411 (N_411,In_1147,In_348);
and U412 (N_412,In_96,In_7);
nor U413 (N_413,In_1123,In_445);
xnor U414 (N_414,In_352,In_643);
nor U415 (N_415,In_566,In_844);
nand U416 (N_416,In_995,In_221);
and U417 (N_417,In_672,In_859);
nor U418 (N_418,In_1288,In_248);
xor U419 (N_419,In_39,In_1333);
and U420 (N_420,In_1133,In_1419);
or U421 (N_421,In_512,In_1195);
nand U422 (N_422,In_519,In_860);
or U423 (N_423,In_75,In_411);
xor U424 (N_424,In_944,In_1197);
nand U425 (N_425,In_628,In_1250);
xnor U426 (N_426,In_1245,In_389);
nand U427 (N_427,In_1374,In_156);
nand U428 (N_428,In_1275,In_1405);
nand U429 (N_429,In_214,In_550);
nand U430 (N_430,In_1124,In_1398);
nand U431 (N_431,In_693,In_84);
nand U432 (N_432,In_698,In_914);
and U433 (N_433,In_1087,In_38);
and U434 (N_434,In_1121,In_1181);
and U435 (N_435,In_501,In_994);
and U436 (N_436,In_122,In_1116);
or U437 (N_437,In_1003,In_80);
nand U438 (N_438,In_171,In_1110);
and U439 (N_439,In_1389,In_316);
nor U440 (N_440,In_323,In_1022);
nor U441 (N_441,In_63,In_125);
nor U442 (N_442,In_1354,In_552);
and U443 (N_443,In_1129,In_1370);
and U444 (N_444,In_1325,In_1040);
xor U445 (N_445,In_253,In_892);
or U446 (N_446,In_42,In_1019);
nand U447 (N_447,In_597,In_50);
or U448 (N_448,In_61,In_930);
nand U449 (N_449,In_308,In_631);
or U450 (N_450,In_999,In_919);
or U451 (N_451,In_19,In_739);
and U452 (N_452,In_28,In_1226);
and U453 (N_453,In_1155,In_298);
xnor U454 (N_454,In_656,In_439);
or U455 (N_455,In_1228,In_1072);
nand U456 (N_456,In_920,In_452);
and U457 (N_457,In_212,In_1426);
or U458 (N_458,In_119,In_1406);
or U459 (N_459,In_1112,In_960);
or U460 (N_460,In_937,In_4);
nand U461 (N_461,In_99,In_1161);
nor U462 (N_462,In_1239,In_1395);
nand U463 (N_463,In_976,In_841);
and U464 (N_464,In_1143,In_1063);
xnor U465 (N_465,In_379,In_1030);
nand U466 (N_466,In_665,In_1050);
nor U467 (N_467,In_74,In_247);
or U468 (N_468,In_651,In_1130);
or U469 (N_469,In_1364,In_1256);
or U470 (N_470,In_421,In_371);
xor U471 (N_471,In_1191,In_696);
and U472 (N_472,In_1109,In_989);
or U473 (N_473,In_473,In_794);
nand U474 (N_474,In_340,In_1383);
xor U475 (N_475,In_1088,In_363);
nand U476 (N_476,In_622,In_1115);
xnor U477 (N_477,In_1169,In_537);
xnor U478 (N_478,In_1493,In_1324);
or U479 (N_479,In_735,In_1202);
or U480 (N_480,In_686,In_394);
nor U481 (N_481,In_1445,In_1347);
and U482 (N_482,In_338,In_1138);
nor U483 (N_483,In_365,In_1014);
nand U484 (N_484,In_0,In_412);
nand U485 (N_485,In_134,In_1234);
nor U486 (N_486,In_368,In_1064);
nor U487 (N_487,In_444,In_654);
nor U488 (N_488,In_152,In_262);
nor U489 (N_489,In_695,In_239);
and U490 (N_490,In_588,In_272);
or U491 (N_491,In_236,In_951);
nor U492 (N_492,In_1176,In_1223);
or U493 (N_493,In_276,In_364);
nand U494 (N_494,In_916,In_203);
nand U495 (N_495,In_723,In_79);
nand U496 (N_496,In_1100,In_1472);
nor U497 (N_497,In_1368,In_1131);
nand U498 (N_498,In_1066,In_613);
or U499 (N_499,In_154,In_1279);
xnor U500 (N_500,N_429,In_1404);
or U501 (N_501,N_273,In_483);
or U502 (N_502,In_1167,N_356);
or U503 (N_503,N_239,In_242);
xnor U504 (N_504,N_92,N_486);
or U505 (N_505,In_12,In_399);
nand U506 (N_506,N_150,In_163);
or U507 (N_507,N_418,N_343);
or U508 (N_508,N_334,N_90);
nor U509 (N_509,In_616,N_59);
and U510 (N_510,In_1023,N_473);
or U511 (N_511,N_374,N_307);
xnor U512 (N_512,N_215,N_81);
nor U513 (N_513,N_220,N_258);
and U514 (N_514,In_36,In_771);
or U515 (N_515,N_120,N_478);
nand U516 (N_516,In_1175,N_450);
nand U517 (N_517,In_370,N_240);
nor U518 (N_518,N_362,N_177);
and U519 (N_519,In_466,In_1427);
or U520 (N_520,In_729,In_330);
or U521 (N_521,N_34,In_353);
and U522 (N_522,In_848,In_820);
nor U523 (N_523,In_509,N_119);
and U524 (N_524,N_95,In_1262);
nor U525 (N_525,In_355,N_65);
nor U526 (N_526,In_1485,N_88);
and U527 (N_527,N_189,N_246);
nand U528 (N_528,N_45,N_25);
nor U529 (N_529,In_302,N_139);
and U530 (N_530,N_336,N_134);
nand U531 (N_531,N_387,In_879);
xor U532 (N_532,N_234,In_907);
nor U533 (N_533,N_376,In_82);
or U534 (N_534,N_82,N_216);
nor U535 (N_535,In_494,N_251);
or U536 (N_536,In_185,N_64);
or U537 (N_537,In_1209,In_991);
nand U538 (N_538,In_553,N_12);
and U539 (N_539,In_1417,N_285);
or U540 (N_540,In_912,N_312);
nor U541 (N_541,N_48,In_531);
xnor U542 (N_542,N_70,In_1215);
or U543 (N_543,N_115,N_71);
nand U544 (N_544,N_411,N_147);
nor U545 (N_545,N_200,N_231);
and U546 (N_546,In_732,In_619);
nor U547 (N_547,In_882,N_194);
nand U548 (N_548,N_289,In_243);
nand U549 (N_549,In_285,N_266);
and U550 (N_550,In_1097,In_429);
nor U551 (N_551,In_1432,In_873);
or U552 (N_552,In_386,In_424);
nand U553 (N_553,N_271,N_102);
nand U554 (N_554,In_358,In_209);
nor U555 (N_555,In_369,In_1373);
nor U556 (N_556,In_149,N_152);
xor U557 (N_557,In_526,In_506);
nand U558 (N_558,N_32,N_109);
nor U559 (N_559,In_795,In_806);
and U560 (N_560,N_367,N_17);
nor U561 (N_561,In_632,N_30);
nand U562 (N_562,N_329,In_1154);
nand U563 (N_563,N_181,In_492);
nand U564 (N_564,In_1017,In_426);
or U565 (N_565,N_328,In_1430);
nor U566 (N_566,N_121,In_514);
or U567 (N_567,N_184,In_931);
nand U568 (N_568,In_361,In_320);
and U569 (N_569,N_116,In_719);
and U570 (N_570,N_402,In_1260);
and U571 (N_571,In_1265,N_208);
nor U572 (N_572,N_230,N_153);
nor U573 (N_573,In_614,N_16);
and U574 (N_574,N_388,In_940);
nor U575 (N_575,In_549,N_406);
nand U576 (N_576,In_392,N_209);
nand U577 (N_577,In_436,In_1024);
nor U578 (N_578,N_224,In_1281);
and U579 (N_579,In_1001,N_244);
nand U580 (N_580,In_43,In_1008);
or U581 (N_581,N_203,In_292);
or U582 (N_582,N_104,N_204);
nand U583 (N_583,N_408,In_642);
nor U584 (N_584,N_22,N_213);
nand U585 (N_585,N_435,In_1061);
nor U586 (N_586,N_364,N_471);
or U587 (N_587,N_454,In_1343);
and U588 (N_588,In_1160,In_1246);
or U589 (N_589,In_988,In_420);
xor U590 (N_590,In_433,N_40);
nor U591 (N_591,N_19,In_16);
and U592 (N_592,In_108,In_177);
or U593 (N_593,In_869,N_170);
xor U594 (N_594,In_403,N_103);
nand U595 (N_595,In_1474,In_513);
or U596 (N_596,In_592,In_855);
nand U597 (N_597,In_884,In_987);
or U598 (N_598,In_1450,In_329);
nand U599 (N_599,In_925,N_359);
nor U600 (N_600,N_495,N_449);
nor U601 (N_601,In_1033,N_171);
nand U602 (N_602,In_1196,N_69);
nor U603 (N_603,In_800,N_320);
nand U604 (N_604,In_1420,In_1271);
nor U605 (N_605,In_760,In_963);
or U606 (N_606,N_324,In_87);
and U607 (N_607,In_1029,N_53);
nand U608 (N_608,N_124,In_1460);
xor U609 (N_609,N_396,N_434);
nand U610 (N_610,N_110,N_113);
or U611 (N_611,N_243,In_996);
and U612 (N_612,In_701,N_86);
nor U613 (N_613,N_341,N_155);
and U614 (N_614,In_711,N_197);
nor U615 (N_615,N_142,N_460);
and U616 (N_616,In_557,In_402);
or U617 (N_617,In_1289,N_316);
nor U618 (N_618,In_422,In_964);
or U619 (N_619,In_543,In_529);
xor U620 (N_620,In_76,In_1301);
and U621 (N_621,N_99,In_200);
nor U622 (N_622,N_314,N_118);
and U623 (N_623,N_61,In_682);
nand U624 (N_624,N_299,In_835);
or U625 (N_625,In_131,N_145);
nor U626 (N_626,In_647,N_403);
or U627 (N_627,In_503,In_1201);
nand U628 (N_628,In_959,N_96);
nand U629 (N_629,N_442,N_229);
nand U630 (N_630,N_133,N_232);
nand U631 (N_631,N_13,N_106);
nand U632 (N_632,N_175,N_1);
nor U633 (N_633,In_179,N_474);
and U634 (N_634,In_1411,N_420);
nor U635 (N_635,N_438,N_303);
and U636 (N_636,In_1321,In_1463);
and U637 (N_637,N_487,N_15);
nand U638 (N_638,In_1377,In_1421);
or U639 (N_639,In_1274,In_840);
nand U640 (N_640,N_37,N_368);
nand U641 (N_641,N_399,N_138);
and U642 (N_642,N_39,N_268);
nand U643 (N_643,N_419,In_1424);
or U644 (N_644,N_38,In_135);
xor U645 (N_645,In_187,N_226);
nor U646 (N_646,In_768,N_295);
xor U647 (N_647,N_163,N_262);
or U648 (N_648,In_377,N_249);
nand U649 (N_649,N_340,In_1177);
xor U650 (N_650,In_142,In_561);
or U651 (N_651,In_1482,N_443);
nand U652 (N_652,In_5,In_530);
and U653 (N_653,N_94,In_1092);
and U654 (N_654,N_462,In_1349);
or U655 (N_655,N_457,N_188);
nand U656 (N_656,In_1442,In_64);
nand U657 (N_657,N_43,N_21);
and U658 (N_658,N_24,N_369);
and U659 (N_659,In_1080,In_1220);
nor U660 (N_660,N_379,N_355);
nand U661 (N_661,In_704,In_1046);
nand U662 (N_662,In_1467,In_941);
or U663 (N_663,In_986,N_275);
nand U664 (N_664,In_1366,In_1457);
xor U665 (N_665,In_565,N_57);
and U666 (N_666,In_1497,In_153);
or U667 (N_667,N_100,N_338);
or U668 (N_668,N_265,In_659);
or U669 (N_669,N_186,N_385);
and U670 (N_670,In_367,N_89);
or U671 (N_671,N_453,In_703);
nand U672 (N_672,N_83,In_604);
xor U673 (N_673,In_865,In_1438);
or U674 (N_674,N_440,In_1403);
nor U675 (N_675,N_360,In_77);
and U676 (N_676,In_164,N_72);
nor U677 (N_677,In_405,N_6);
nor U678 (N_678,N_405,In_1422);
nand U679 (N_679,In_1227,N_36);
or U680 (N_680,N_325,In_845);
or U681 (N_681,In_1074,N_330);
nor U682 (N_682,N_270,N_91);
and U683 (N_683,In_1478,In_1476);
and U684 (N_684,N_196,In_47);
nor U685 (N_685,N_395,In_168);
xnor U686 (N_686,In_1186,In_257);
nand U687 (N_687,In_147,In_266);
nor U688 (N_688,In_1401,In_176);
xor U689 (N_689,N_375,N_242);
xnor U690 (N_690,N_143,In_691);
and U691 (N_691,In_893,N_427);
nor U692 (N_692,In_273,In_650);
or U693 (N_693,N_63,In_351);
nor U694 (N_694,N_302,N_452);
nand U695 (N_695,N_66,N_2);
nor U696 (N_696,N_476,N_212);
nor U697 (N_697,In_836,In_1407);
nand U698 (N_698,In_456,In_1322);
nor U699 (N_699,In_1365,In_997);
xor U700 (N_700,In_66,N_237);
and U701 (N_701,N_371,N_353);
nor U702 (N_702,N_27,N_391);
xor U703 (N_703,N_317,N_176);
xnor U704 (N_704,In_45,In_322);
and U705 (N_705,In_1267,In_507);
nor U706 (N_706,In_580,In_319);
or U707 (N_707,In_25,In_201);
or U708 (N_708,N_3,In_138);
or U709 (N_709,N_404,In_317);
xor U710 (N_710,In_1026,In_518);
or U711 (N_711,N_74,N_458);
nand U712 (N_712,In_515,N_437);
xor U713 (N_713,N_112,N_497);
nor U714 (N_714,In_1311,N_107);
and U715 (N_715,In_1494,N_245);
nand U716 (N_716,In_180,N_472);
and U717 (N_717,In_1447,N_187);
xor U718 (N_718,N_217,In_1372);
xor U719 (N_719,In_516,In_992);
and U720 (N_720,N_342,N_221);
nand U721 (N_721,N_5,N_358);
xor U722 (N_722,N_447,N_386);
nor U723 (N_723,In_67,N_219);
nand U724 (N_724,In_971,N_430);
or U725 (N_725,N_9,N_18);
nor U726 (N_726,In_390,In_1217);
xor U727 (N_727,N_46,In_733);
and U728 (N_728,In_1371,N_499);
or U729 (N_729,N_101,In_1351);
xor U730 (N_730,In_827,In_346);
or U731 (N_731,N_370,In_1339);
nand U732 (N_732,In_1241,In_684);
and U733 (N_733,N_425,N_52);
nor U734 (N_734,N_125,N_301);
or U735 (N_735,N_417,N_305);
xor U736 (N_736,In_237,In_878);
or U737 (N_737,In_81,N_47);
xor U738 (N_738,N_267,N_248);
and U739 (N_739,In_1178,N_85);
nor U740 (N_740,In_1443,N_410);
nor U741 (N_741,In_1391,In_398);
xor U742 (N_742,In_1320,N_190);
and U743 (N_743,In_744,In_305);
or U744 (N_744,In_98,N_313);
or U745 (N_745,N_54,N_68);
or U746 (N_746,N_128,In_578);
nor U747 (N_747,N_484,N_286);
nand U748 (N_748,N_205,In_1291);
and U749 (N_749,N_377,In_586);
nor U750 (N_750,N_493,In_745);
nand U751 (N_751,In_635,N_254);
nor U752 (N_752,N_482,N_23);
or U753 (N_753,In_1489,N_252);
nor U754 (N_754,N_214,N_298);
nand U755 (N_755,In_1183,N_127);
and U756 (N_756,N_361,N_297);
nor U757 (N_757,N_227,N_284);
xnor U758 (N_758,N_461,N_8);
or U759 (N_759,N_277,N_401);
or U760 (N_760,N_479,In_510);
nor U761 (N_761,In_823,In_1418);
nand U762 (N_762,In_1098,In_259);
nor U763 (N_763,N_261,In_258);
nor U764 (N_764,N_309,N_287);
nor U765 (N_765,N_201,In_697);
or U766 (N_766,N_78,In_943);
nand U767 (N_767,N_350,N_424);
and U768 (N_768,N_272,N_415);
nand U769 (N_769,N_491,In_505);
nor U770 (N_770,In_1400,In_786);
and U771 (N_771,In_834,N_422);
or U772 (N_772,N_218,In_395);
and U773 (N_773,N_296,In_1208);
nor U774 (N_774,In_1114,In_946);
and U775 (N_775,N_233,In_1257);
or U776 (N_776,In_430,In_327);
or U777 (N_777,In_1136,N_211);
nand U778 (N_778,In_8,N_394);
or U779 (N_779,In_815,In_376);
or U780 (N_780,In_652,N_349);
and U781 (N_781,In_625,In_1018);
nor U782 (N_782,In_291,N_306);
nand U783 (N_783,N_141,In_852);
nand U784 (N_784,In_1011,N_269);
and U785 (N_785,N_346,N_97);
and U786 (N_786,In_1455,In_754);
and U787 (N_787,N_93,N_206);
nor U788 (N_788,N_14,In_681);
and U789 (N_789,N_247,In_885);
or U790 (N_790,N_496,N_381);
xor U791 (N_791,In_170,N_383);
or U792 (N_792,N_77,N_129);
and U793 (N_793,N_409,N_73);
nand U794 (N_794,N_393,In_447);
and U795 (N_795,N_160,N_444);
nor U796 (N_796,N_111,In_217);
and U797 (N_797,In_167,N_455);
xnor U798 (N_798,In_582,In_432);
or U799 (N_799,N_198,In_675);
nand U800 (N_800,In_1120,N_144);
and U801 (N_801,N_477,In_62);
and U802 (N_802,In_1441,N_291);
and U803 (N_803,In_380,In_54);
nor U804 (N_804,In_1488,N_351);
or U805 (N_805,N_31,N_207);
and U806 (N_806,In_1319,In_791);
or U807 (N_807,In_166,In_244);
nand U808 (N_808,N_260,N_498);
or U809 (N_809,N_426,In_194);
or U810 (N_810,In_1352,In_1039);
and U811 (N_811,N_263,In_1376);
and U812 (N_812,In_46,In_1127);
or U813 (N_813,In_140,In_829);
nor U814 (N_814,In_661,N_253);
nor U815 (N_815,N_42,In_1096);
and U816 (N_816,In_927,N_80);
and U817 (N_817,N_41,N_448);
nand U818 (N_818,N_300,In_117);
nor U819 (N_819,N_238,In_295);
and U820 (N_820,In_637,N_439);
xnor U821 (N_821,N_304,In_471);
nand U822 (N_822,N_290,In_300);
or U823 (N_823,In_463,N_35);
nor U824 (N_824,In_1083,In_145);
nor U825 (N_825,N_132,In_720);
or U826 (N_826,N_384,N_58);
nand U827 (N_827,In_525,N_167);
and U828 (N_828,In_575,N_397);
xor U829 (N_829,In_1187,In_756);
nor U830 (N_830,In_1416,In_1338);
and U831 (N_831,N_412,N_149);
or U832 (N_832,In_18,N_459);
xnor U833 (N_833,N_292,In_470);
or U834 (N_834,In_864,N_33);
and U835 (N_835,N_202,N_60);
and U836 (N_836,In_1104,N_492);
nor U837 (N_837,N_446,N_126);
nor U838 (N_838,N_228,N_428);
and U839 (N_839,In_779,In_461);
or U840 (N_840,N_468,In_793);
xnor U841 (N_841,N_421,N_117);
nor U842 (N_842,N_105,In_2);
or U843 (N_843,N_348,N_365);
and U844 (N_844,In_814,N_432);
nand U845 (N_845,In_335,In_1385);
or U846 (N_846,N_282,N_172);
or U847 (N_847,N_413,N_168);
nand U848 (N_848,N_310,N_183);
xnor U849 (N_849,N_293,N_366);
nand U850 (N_850,In_734,N_29);
xnor U851 (N_851,In_1184,N_319);
nand U852 (N_852,In_1132,In_1070);
xnor U853 (N_853,In_520,N_288);
nand U854 (N_854,In_387,In_431);
or U855 (N_855,In_227,In_132);
nand U856 (N_856,In_1229,N_0);
nand U857 (N_857,In_521,In_1107);
or U858 (N_858,N_192,In_1286);
nor U859 (N_859,In_618,N_164);
or U860 (N_860,In_234,In_1490);
nor U861 (N_861,N_475,N_154);
xor U862 (N_862,In_219,In_1299);
or U863 (N_863,In_400,N_256);
and U864 (N_864,In_599,In_626);
nor U865 (N_865,In_942,N_62);
xor U866 (N_866,N_323,N_294);
nand U867 (N_867,In_906,N_140);
nand U868 (N_868,N_223,N_87);
and U869 (N_869,N_122,N_67);
or U870 (N_870,N_169,N_151);
nand U871 (N_871,In_993,In_600);
and U872 (N_872,In_577,In_858);
nand U873 (N_873,In_830,In_184);
nand U874 (N_874,N_463,N_315);
and U875 (N_875,In_1413,In_288);
nor U876 (N_876,N_257,In_714);
and U877 (N_877,In_523,N_55);
nand U878 (N_878,N_264,N_281);
nor U879 (N_879,N_390,In_772);
nand U880 (N_880,N_280,In_1294);
and U881 (N_881,In_880,N_433);
and U882 (N_882,In_235,In_464);
nand U883 (N_883,In_967,In_1150);
nand U884 (N_884,N_7,In_977);
nor U885 (N_885,In_414,N_236);
and U886 (N_886,N_489,N_210);
nand U887 (N_887,In_1429,N_481);
nand U888 (N_888,N_321,N_466);
nand U889 (N_889,In_1036,In_601);
xnor U890 (N_890,N_191,N_274);
xor U891 (N_891,In_610,In_688);
and U892 (N_892,In_326,N_136);
or U893 (N_893,In_1037,N_123);
and U894 (N_894,N_193,N_337);
and U895 (N_895,In_137,N_114);
nor U896 (N_896,In_881,N_276);
nor U897 (N_897,In_339,In_817);
xnor U898 (N_898,In_556,In_478);
nand U899 (N_899,In_1425,N_84);
or U900 (N_900,N_173,N_161);
nor U901 (N_901,N_56,N_326);
and U902 (N_902,N_494,In_155);
nor U903 (N_903,In_832,In_1173);
nor U904 (N_904,In_1475,N_327);
nor U905 (N_905,N_222,In_811);
nand U906 (N_906,N_347,In_344);
or U907 (N_907,In_476,N_180);
and U908 (N_908,In_1465,In_1057);
and U909 (N_909,N_11,In_1207);
nand U910 (N_910,In_488,In_1117);
or U911 (N_911,N_423,In_1128);
nor U912 (N_912,In_251,N_241);
or U913 (N_913,N_311,In_1171);
nor U914 (N_914,N_159,In_1126);
and U915 (N_915,N_345,N_195);
nand U916 (N_916,In_1094,In_1326);
or U917 (N_917,In_1170,In_973);
or U918 (N_918,N_28,N_135);
and U919 (N_919,N_255,N_485);
nand U920 (N_920,N_400,N_398);
or U921 (N_921,N_464,In_715);
or U922 (N_922,N_373,In_3);
and U923 (N_923,In_1487,In_593);
xor U924 (N_924,In_287,In_408);
or U925 (N_925,In_911,In_312);
or U926 (N_926,In_985,In_590);
and U927 (N_927,In_1231,In_1095);
or U928 (N_928,In_480,In_1182);
nand U929 (N_929,N_357,In_294);
and U930 (N_930,N_157,N_382);
or U931 (N_931,In_966,In_336);
and U932 (N_932,N_76,N_322);
or U933 (N_933,In_95,In_277);
nor U934 (N_934,In_1,N_146);
xnor U935 (N_935,N_162,N_354);
and U936 (N_936,In_1111,N_441);
nand U937 (N_937,N_185,N_51);
nor U938 (N_938,N_283,N_50);
and U939 (N_939,In_1306,N_372);
or U940 (N_940,N_10,N_165);
nor U941 (N_941,N_174,In_572);
nand U942 (N_942,In_901,In_460);
or U943 (N_943,N_131,In_89);
nor U944 (N_944,In_205,In_868);
and U945 (N_945,In_891,N_26);
nand U946 (N_946,In_658,N_331);
nand U947 (N_947,N_414,In_1477);
xnor U948 (N_948,N_235,N_416);
nor U949 (N_949,In_314,N_431);
and U950 (N_950,N_156,In_1284);
nand U951 (N_951,In_354,In_270);
nor U952 (N_952,N_137,In_751);
and U953 (N_953,N_44,N_392);
xor U954 (N_954,N_178,N_278);
or U955 (N_955,N_166,N_380);
nand U956 (N_956,In_1163,In_1436);
xnor U957 (N_957,N_445,N_456);
nand U958 (N_958,In_903,N_378);
or U959 (N_959,N_469,In_249);
or U960 (N_960,N_108,In_1302);
nand U961 (N_961,N_407,N_179);
or U962 (N_962,In_524,In_172);
or U963 (N_963,In_254,In_271);
or U964 (N_964,N_225,In_139);
and U965 (N_965,In_936,N_490);
and U966 (N_966,In_1481,In_111);
nor U967 (N_967,N_75,N_389);
nor U968 (N_968,In_20,N_279);
nor U969 (N_969,In_226,In_689);
nand U970 (N_970,In_1277,In_984);
nand U971 (N_971,In_1090,N_199);
nor U972 (N_972,N_352,In_1359);
and U973 (N_973,N_182,In_309);
nor U974 (N_974,In_917,N_470);
and U975 (N_975,N_49,In_143);
nor U976 (N_976,In_14,N_308);
nand U977 (N_977,In_810,In_638);
or U978 (N_978,N_339,N_451);
and U979 (N_979,In_974,N_148);
and U980 (N_980,In_683,In_534);
and U981 (N_981,In_1145,In_1158);
nor U982 (N_982,N_98,In_796);
and U983 (N_983,N_467,N_480);
and U984 (N_984,N_20,N_363);
or U985 (N_985,In_950,In_690);
nor U986 (N_986,In_86,N_130);
and U987 (N_987,N_488,In_311);
nand U988 (N_988,In_573,In_1412);
and U989 (N_989,In_653,N_483);
nor U990 (N_990,N_158,N_250);
nor U991 (N_991,N_335,N_436);
nand U992 (N_992,In_114,In_68);
or U993 (N_993,N_318,N_333);
and U994 (N_994,N_79,N_465);
or U995 (N_995,N_259,N_4);
nand U996 (N_996,In_929,In_1356);
nor U997 (N_997,In_383,In_1009);
or U998 (N_998,In_904,In_192);
and U999 (N_999,N_344,N_332);
or U1000 (N_1000,N_835,N_673);
nor U1001 (N_1001,N_920,N_570);
nand U1002 (N_1002,N_867,N_915);
nand U1003 (N_1003,N_983,N_707);
nor U1004 (N_1004,N_781,N_783);
xor U1005 (N_1005,N_515,N_618);
and U1006 (N_1006,N_885,N_774);
nand U1007 (N_1007,N_569,N_685);
nor U1008 (N_1008,N_821,N_880);
nand U1009 (N_1009,N_695,N_706);
xor U1010 (N_1010,N_993,N_896);
and U1011 (N_1011,N_542,N_757);
nor U1012 (N_1012,N_971,N_933);
xnor U1013 (N_1013,N_625,N_909);
or U1014 (N_1014,N_710,N_646);
nor U1015 (N_1015,N_639,N_592);
or U1016 (N_1016,N_862,N_791);
nand U1017 (N_1017,N_760,N_561);
and U1018 (N_1018,N_982,N_577);
nand U1019 (N_1019,N_770,N_892);
or U1020 (N_1020,N_705,N_614);
and U1021 (N_1021,N_801,N_711);
nand U1022 (N_1022,N_755,N_683);
or U1023 (N_1023,N_923,N_552);
nand U1024 (N_1024,N_884,N_582);
nor U1025 (N_1025,N_881,N_556);
nand U1026 (N_1026,N_979,N_763);
xor U1027 (N_1027,N_930,N_658);
and U1028 (N_1028,N_598,N_860);
and U1029 (N_1029,N_722,N_861);
and U1030 (N_1030,N_546,N_959);
nor U1031 (N_1031,N_626,N_693);
or U1032 (N_1032,N_788,N_822);
nand U1033 (N_1033,N_652,N_708);
nand U1034 (N_1034,N_532,N_654);
nor U1035 (N_1035,N_585,N_777);
and U1036 (N_1036,N_751,N_846);
and U1037 (N_1037,N_962,N_864);
or U1038 (N_1038,N_858,N_938);
xnor U1039 (N_1039,N_634,N_667);
or U1040 (N_1040,N_808,N_502);
or U1041 (N_1041,N_914,N_550);
and U1042 (N_1042,N_537,N_974);
nor U1043 (N_1043,N_629,N_954);
and U1044 (N_1044,N_796,N_630);
or U1045 (N_1045,N_599,N_610);
and U1046 (N_1046,N_507,N_588);
nor U1047 (N_1047,N_919,N_544);
nor U1048 (N_1048,N_735,N_680);
nand U1049 (N_1049,N_698,N_633);
nand U1050 (N_1050,N_522,N_733);
or U1051 (N_1051,N_514,N_622);
nor U1052 (N_1052,N_703,N_752);
nor U1053 (N_1053,N_719,N_779);
xor U1054 (N_1054,N_782,N_603);
and U1055 (N_1055,N_812,N_843);
xor U1056 (N_1056,N_631,N_747);
nand U1057 (N_1057,N_677,N_557);
or U1058 (N_1058,N_593,N_728);
and U1059 (N_1059,N_955,N_551);
or U1060 (N_1060,N_859,N_917);
nor U1061 (N_1061,N_912,N_510);
nand U1062 (N_1062,N_769,N_623);
nor U1063 (N_1063,N_910,N_668);
xor U1064 (N_1064,N_850,N_837);
nand U1065 (N_1065,N_978,N_764);
nand U1066 (N_1066,N_656,N_748);
or U1067 (N_1067,N_823,N_688);
nor U1068 (N_1068,N_824,N_987);
or U1069 (N_1069,N_647,N_718);
nor U1070 (N_1070,N_968,N_619);
or U1071 (N_1071,N_712,N_597);
xnor U1072 (N_1072,N_526,N_804);
and U1073 (N_1073,N_571,N_661);
xnor U1074 (N_1074,N_724,N_977);
xor U1075 (N_1075,N_819,N_513);
nor U1076 (N_1076,N_741,N_746);
or U1077 (N_1077,N_876,N_818);
nand U1078 (N_1078,N_702,N_508);
or U1079 (N_1079,N_538,N_762);
nor U1080 (N_1080,N_809,N_980);
and U1081 (N_1081,N_640,N_701);
xor U1082 (N_1082,N_990,N_607);
and U1083 (N_1083,N_805,N_992);
and U1084 (N_1084,N_574,N_644);
nand U1085 (N_1085,N_612,N_726);
and U1086 (N_1086,N_643,N_567);
nor U1087 (N_1087,N_736,N_744);
or U1088 (N_1088,N_972,N_901);
nor U1089 (N_1089,N_842,N_998);
xor U1090 (N_1090,N_841,N_931);
nor U1091 (N_1091,N_672,N_872);
nand U1092 (N_1092,N_581,N_768);
and U1093 (N_1093,N_676,N_681);
or U1094 (N_1094,N_554,N_628);
and U1095 (N_1095,N_519,N_694);
nor U1096 (N_1096,N_689,N_516);
and U1097 (N_1097,N_590,N_523);
nor U1098 (N_1098,N_601,N_583);
xnor U1099 (N_1099,N_848,N_638);
nor U1100 (N_1100,N_738,N_536);
nand U1101 (N_1101,N_943,N_797);
nand U1102 (N_1102,N_579,N_802);
nor U1103 (N_1103,N_727,N_976);
nand U1104 (N_1104,N_813,N_854);
nand U1105 (N_1105,N_709,N_773);
nor U1106 (N_1106,N_731,N_521);
nand U1107 (N_1107,N_776,N_500);
and U1108 (N_1108,N_820,N_832);
and U1109 (N_1109,N_855,N_602);
or U1110 (N_1110,N_794,N_922);
and U1111 (N_1111,N_965,N_729);
xnor U1112 (N_1112,N_863,N_960);
nand U1113 (N_1113,N_684,N_621);
xor U1114 (N_1114,N_595,N_866);
nand U1115 (N_1115,N_714,N_657);
nor U1116 (N_1116,N_799,N_816);
and U1117 (N_1117,N_947,N_939);
nor U1118 (N_1118,N_834,N_997);
nor U1119 (N_1119,N_995,N_950);
and U1120 (N_1120,N_771,N_525);
or U1121 (N_1121,N_810,N_697);
nor U1122 (N_1122,N_999,N_874);
or U1123 (N_1123,N_991,N_806);
or U1124 (N_1124,N_961,N_682);
xnor U1125 (N_1125,N_568,N_784);
or U1126 (N_1126,N_994,N_753);
nand U1127 (N_1127,N_775,N_948);
nor U1128 (N_1128,N_989,N_749);
nor U1129 (N_1129,N_573,N_509);
and U1130 (N_1130,N_932,N_674);
and U1131 (N_1131,N_678,N_754);
nor U1132 (N_1132,N_615,N_660);
nand U1133 (N_1133,N_966,N_534);
and U1134 (N_1134,N_944,N_870);
nor U1135 (N_1135,N_543,N_566);
nor U1136 (N_1136,N_767,N_565);
or U1137 (N_1137,N_596,N_833);
or U1138 (N_1138,N_845,N_815);
xnor U1139 (N_1139,N_985,N_897);
nor U1140 (N_1140,N_547,N_851);
and U1141 (N_1141,N_576,N_838);
nor U1142 (N_1142,N_575,N_953);
or U1143 (N_1143,N_559,N_716);
xnor U1144 (N_1144,N_975,N_811);
and U1145 (N_1145,N_967,N_642);
nand U1146 (N_1146,N_904,N_969);
nand U1147 (N_1147,N_873,N_758);
or U1148 (N_1148,N_902,N_518);
nor U1149 (N_1149,N_878,N_789);
and U1150 (N_1150,N_928,N_879);
or U1151 (N_1151,N_963,N_996);
nand U1152 (N_1152,N_512,N_605);
nand U1153 (N_1153,N_964,N_692);
nand U1154 (N_1154,N_541,N_888);
or U1155 (N_1155,N_609,N_679);
or U1156 (N_1156,N_732,N_893);
xnor U1157 (N_1157,N_700,N_800);
xnor U1158 (N_1158,N_529,N_555);
and U1159 (N_1159,N_535,N_882);
and U1160 (N_1160,N_869,N_825);
nand U1161 (N_1161,N_949,N_857);
xnor U1162 (N_1162,N_737,N_687);
nor U1163 (N_1163,N_696,N_785);
nand U1164 (N_1164,N_578,N_540);
and U1165 (N_1165,N_600,N_586);
nor U1166 (N_1166,N_887,N_594);
nand U1167 (N_1167,N_986,N_942);
nand U1168 (N_1168,N_505,N_742);
nor U1169 (N_1169,N_827,N_662);
or U1170 (N_1170,N_666,N_759);
xnor U1171 (N_1171,N_911,N_717);
and U1172 (N_1172,N_655,N_756);
nor U1173 (N_1173,N_894,N_527);
or U1174 (N_1174,N_852,N_899);
nor U1175 (N_1175,N_956,N_871);
or U1176 (N_1176,N_958,N_957);
or U1177 (N_1177,N_675,N_814);
nand U1178 (N_1178,N_787,N_608);
nor U1179 (N_1179,N_921,N_686);
and U1180 (N_1180,N_780,N_839);
xnor U1181 (N_1181,N_765,N_511);
or U1182 (N_1182,N_828,N_918);
xnor U1183 (N_1183,N_988,N_831);
or U1184 (N_1184,N_792,N_699);
and U1185 (N_1185,N_984,N_925);
and U1186 (N_1186,N_611,N_793);
or U1187 (N_1187,N_946,N_691);
xor U1188 (N_1188,N_836,N_613);
or U1189 (N_1189,N_665,N_604);
nand U1190 (N_1190,N_637,N_591);
nand U1191 (N_1191,N_635,N_790);
nor U1192 (N_1192,N_890,N_501);
or U1193 (N_1193,N_504,N_648);
or U1194 (N_1194,N_730,N_530);
and U1195 (N_1195,N_506,N_981);
or U1196 (N_1196,N_720,N_934);
or U1197 (N_1197,N_617,N_929);
nand U1198 (N_1198,N_669,N_817);
and U1199 (N_1199,N_589,N_826);
or U1200 (N_1200,N_883,N_649);
and U1201 (N_1201,N_937,N_853);
nor U1202 (N_1202,N_916,N_739);
nor U1203 (N_1203,N_889,N_713);
or U1204 (N_1204,N_723,N_553);
nor U1205 (N_1205,N_690,N_562);
nand U1206 (N_1206,N_645,N_533);
and U1207 (N_1207,N_548,N_905);
and U1208 (N_1208,N_973,N_663);
or U1209 (N_1209,N_725,N_970);
nor U1210 (N_1210,N_903,N_772);
and U1211 (N_1211,N_898,N_524);
xnor U1212 (N_1212,N_795,N_951);
nand U1213 (N_1213,N_952,N_653);
xnor U1214 (N_1214,N_875,N_503);
or U1215 (N_1215,N_520,N_616);
nor U1216 (N_1216,N_913,N_829);
or U1217 (N_1217,N_664,N_580);
or U1218 (N_1218,N_830,N_906);
and U1219 (N_1219,N_778,N_670);
and U1220 (N_1220,N_807,N_908);
nand U1221 (N_1221,N_627,N_844);
or U1222 (N_1222,N_715,N_868);
nor U1223 (N_1223,N_940,N_895);
or U1224 (N_1224,N_935,N_886);
nand U1225 (N_1225,N_606,N_927);
and U1226 (N_1226,N_734,N_704);
nand U1227 (N_1227,N_517,N_651);
nand U1228 (N_1228,N_877,N_761);
nand U1229 (N_1229,N_659,N_624);
nor U1230 (N_1230,N_560,N_766);
nand U1231 (N_1231,N_549,N_721);
or U1232 (N_1232,N_558,N_803);
and U1233 (N_1233,N_650,N_856);
or U1234 (N_1234,N_564,N_926);
and U1235 (N_1235,N_865,N_849);
xor U1236 (N_1236,N_641,N_907);
nor U1237 (N_1237,N_945,N_786);
nor U1238 (N_1238,N_539,N_840);
and U1239 (N_1239,N_545,N_620);
xor U1240 (N_1240,N_900,N_636);
nand U1241 (N_1241,N_743,N_528);
nand U1242 (N_1242,N_632,N_750);
nand U1243 (N_1243,N_572,N_563);
or U1244 (N_1244,N_671,N_936);
nand U1245 (N_1245,N_847,N_531);
nand U1246 (N_1246,N_740,N_891);
or U1247 (N_1247,N_941,N_584);
nor U1248 (N_1248,N_587,N_798);
and U1249 (N_1249,N_924,N_745);
and U1250 (N_1250,N_750,N_557);
nand U1251 (N_1251,N_537,N_751);
nand U1252 (N_1252,N_945,N_961);
nor U1253 (N_1253,N_865,N_963);
or U1254 (N_1254,N_956,N_961);
nand U1255 (N_1255,N_602,N_671);
nor U1256 (N_1256,N_730,N_700);
xnor U1257 (N_1257,N_766,N_996);
nand U1258 (N_1258,N_718,N_512);
and U1259 (N_1259,N_959,N_913);
and U1260 (N_1260,N_799,N_911);
and U1261 (N_1261,N_633,N_746);
and U1262 (N_1262,N_625,N_847);
or U1263 (N_1263,N_851,N_601);
nor U1264 (N_1264,N_967,N_700);
or U1265 (N_1265,N_734,N_858);
xnor U1266 (N_1266,N_578,N_817);
nor U1267 (N_1267,N_825,N_804);
nand U1268 (N_1268,N_820,N_750);
xnor U1269 (N_1269,N_997,N_548);
xor U1270 (N_1270,N_991,N_596);
and U1271 (N_1271,N_793,N_792);
and U1272 (N_1272,N_534,N_677);
or U1273 (N_1273,N_583,N_733);
xnor U1274 (N_1274,N_708,N_820);
and U1275 (N_1275,N_731,N_930);
nand U1276 (N_1276,N_861,N_698);
or U1277 (N_1277,N_607,N_605);
and U1278 (N_1278,N_676,N_758);
xnor U1279 (N_1279,N_794,N_737);
and U1280 (N_1280,N_715,N_583);
or U1281 (N_1281,N_825,N_802);
or U1282 (N_1282,N_623,N_621);
nand U1283 (N_1283,N_826,N_733);
or U1284 (N_1284,N_914,N_840);
nand U1285 (N_1285,N_501,N_815);
xnor U1286 (N_1286,N_988,N_663);
and U1287 (N_1287,N_686,N_933);
and U1288 (N_1288,N_790,N_567);
nand U1289 (N_1289,N_762,N_993);
nor U1290 (N_1290,N_745,N_552);
and U1291 (N_1291,N_686,N_679);
or U1292 (N_1292,N_501,N_939);
nand U1293 (N_1293,N_650,N_658);
nand U1294 (N_1294,N_729,N_792);
and U1295 (N_1295,N_776,N_679);
nand U1296 (N_1296,N_554,N_702);
nand U1297 (N_1297,N_587,N_567);
nand U1298 (N_1298,N_616,N_611);
nor U1299 (N_1299,N_792,N_620);
and U1300 (N_1300,N_847,N_692);
and U1301 (N_1301,N_769,N_886);
nor U1302 (N_1302,N_892,N_729);
or U1303 (N_1303,N_744,N_937);
and U1304 (N_1304,N_876,N_863);
nand U1305 (N_1305,N_887,N_502);
nor U1306 (N_1306,N_927,N_842);
nand U1307 (N_1307,N_663,N_840);
nand U1308 (N_1308,N_579,N_699);
nor U1309 (N_1309,N_985,N_988);
nor U1310 (N_1310,N_503,N_721);
and U1311 (N_1311,N_956,N_720);
nand U1312 (N_1312,N_855,N_797);
and U1313 (N_1313,N_836,N_778);
or U1314 (N_1314,N_528,N_684);
or U1315 (N_1315,N_888,N_957);
nor U1316 (N_1316,N_950,N_988);
nor U1317 (N_1317,N_839,N_875);
nor U1318 (N_1318,N_565,N_831);
nor U1319 (N_1319,N_855,N_868);
nor U1320 (N_1320,N_887,N_552);
xor U1321 (N_1321,N_583,N_656);
nand U1322 (N_1322,N_818,N_755);
nor U1323 (N_1323,N_872,N_809);
nor U1324 (N_1324,N_754,N_511);
and U1325 (N_1325,N_797,N_756);
nor U1326 (N_1326,N_834,N_905);
nand U1327 (N_1327,N_529,N_727);
nor U1328 (N_1328,N_838,N_740);
xor U1329 (N_1329,N_961,N_564);
nor U1330 (N_1330,N_585,N_916);
and U1331 (N_1331,N_765,N_644);
or U1332 (N_1332,N_993,N_819);
and U1333 (N_1333,N_560,N_738);
nand U1334 (N_1334,N_641,N_547);
nor U1335 (N_1335,N_637,N_651);
and U1336 (N_1336,N_861,N_857);
xor U1337 (N_1337,N_655,N_608);
and U1338 (N_1338,N_722,N_977);
nor U1339 (N_1339,N_748,N_818);
nand U1340 (N_1340,N_562,N_788);
and U1341 (N_1341,N_697,N_756);
nand U1342 (N_1342,N_780,N_729);
xor U1343 (N_1343,N_573,N_939);
nor U1344 (N_1344,N_510,N_840);
and U1345 (N_1345,N_873,N_525);
nor U1346 (N_1346,N_912,N_565);
xnor U1347 (N_1347,N_767,N_507);
nand U1348 (N_1348,N_560,N_991);
nand U1349 (N_1349,N_941,N_835);
and U1350 (N_1350,N_638,N_760);
nor U1351 (N_1351,N_865,N_725);
xor U1352 (N_1352,N_910,N_846);
or U1353 (N_1353,N_690,N_875);
nor U1354 (N_1354,N_603,N_597);
xnor U1355 (N_1355,N_904,N_671);
and U1356 (N_1356,N_904,N_573);
nand U1357 (N_1357,N_995,N_915);
nand U1358 (N_1358,N_507,N_746);
nand U1359 (N_1359,N_744,N_703);
and U1360 (N_1360,N_774,N_973);
and U1361 (N_1361,N_551,N_790);
xor U1362 (N_1362,N_630,N_876);
nand U1363 (N_1363,N_702,N_663);
nor U1364 (N_1364,N_893,N_951);
or U1365 (N_1365,N_806,N_718);
nor U1366 (N_1366,N_916,N_551);
and U1367 (N_1367,N_663,N_835);
nor U1368 (N_1368,N_933,N_584);
or U1369 (N_1369,N_778,N_709);
nand U1370 (N_1370,N_856,N_848);
or U1371 (N_1371,N_973,N_532);
nand U1372 (N_1372,N_693,N_531);
nand U1373 (N_1373,N_733,N_624);
nor U1374 (N_1374,N_699,N_937);
or U1375 (N_1375,N_812,N_929);
or U1376 (N_1376,N_629,N_623);
nand U1377 (N_1377,N_991,N_899);
xor U1378 (N_1378,N_603,N_920);
or U1379 (N_1379,N_898,N_587);
and U1380 (N_1380,N_880,N_810);
and U1381 (N_1381,N_986,N_748);
nand U1382 (N_1382,N_774,N_840);
or U1383 (N_1383,N_705,N_858);
nand U1384 (N_1384,N_935,N_700);
or U1385 (N_1385,N_607,N_982);
nor U1386 (N_1386,N_686,N_820);
nor U1387 (N_1387,N_931,N_620);
nand U1388 (N_1388,N_833,N_916);
xnor U1389 (N_1389,N_662,N_915);
and U1390 (N_1390,N_625,N_606);
nand U1391 (N_1391,N_852,N_724);
nand U1392 (N_1392,N_694,N_744);
nor U1393 (N_1393,N_955,N_948);
nor U1394 (N_1394,N_832,N_635);
and U1395 (N_1395,N_936,N_523);
nand U1396 (N_1396,N_639,N_989);
nand U1397 (N_1397,N_615,N_762);
xnor U1398 (N_1398,N_630,N_865);
nand U1399 (N_1399,N_721,N_674);
and U1400 (N_1400,N_540,N_551);
and U1401 (N_1401,N_855,N_753);
nor U1402 (N_1402,N_808,N_939);
or U1403 (N_1403,N_930,N_817);
or U1404 (N_1404,N_563,N_981);
nand U1405 (N_1405,N_912,N_868);
or U1406 (N_1406,N_610,N_851);
and U1407 (N_1407,N_715,N_777);
and U1408 (N_1408,N_724,N_996);
and U1409 (N_1409,N_727,N_782);
nand U1410 (N_1410,N_738,N_797);
or U1411 (N_1411,N_510,N_518);
or U1412 (N_1412,N_957,N_679);
xnor U1413 (N_1413,N_572,N_805);
nor U1414 (N_1414,N_964,N_987);
nand U1415 (N_1415,N_508,N_807);
or U1416 (N_1416,N_686,N_659);
nor U1417 (N_1417,N_762,N_722);
xor U1418 (N_1418,N_829,N_851);
or U1419 (N_1419,N_536,N_715);
nor U1420 (N_1420,N_653,N_861);
nand U1421 (N_1421,N_980,N_726);
nand U1422 (N_1422,N_800,N_706);
nor U1423 (N_1423,N_786,N_872);
nor U1424 (N_1424,N_950,N_517);
nand U1425 (N_1425,N_707,N_974);
or U1426 (N_1426,N_928,N_988);
or U1427 (N_1427,N_952,N_979);
and U1428 (N_1428,N_577,N_766);
or U1429 (N_1429,N_647,N_608);
or U1430 (N_1430,N_867,N_579);
or U1431 (N_1431,N_752,N_571);
or U1432 (N_1432,N_822,N_850);
xor U1433 (N_1433,N_500,N_545);
or U1434 (N_1434,N_526,N_556);
nor U1435 (N_1435,N_868,N_807);
or U1436 (N_1436,N_713,N_887);
nor U1437 (N_1437,N_527,N_721);
or U1438 (N_1438,N_527,N_608);
and U1439 (N_1439,N_959,N_995);
or U1440 (N_1440,N_943,N_791);
nor U1441 (N_1441,N_583,N_887);
or U1442 (N_1442,N_609,N_706);
xnor U1443 (N_1443,N_741,N_770);
nor U1444 (N_1444,N_590,N_545);
or U1445 (N_1445,N_643,N_550);
nor U1446 (N_1446,N_677,N_560);
and U1447 (N_1447,N_853,N_909);
and U1448 (N_1448,N_540,N_929);
xor U1449 (N_1449,N_849,N_765);
nor U1450 (N_1450,N_732,N_566);
or U1451 (N_1451,N_511,N_638);
nand U1452 (N_1452,N_937,N_507);
nand U1453 (N_1453,N_702,N_876);
and U1454 (N_1454,N_569,N_538);
or U1455 (N_1455,N_974,N_543);
xor U1456 (N_1456,N_584,N_553);
xnor U1457 (N_1457,N_749,N_729);
nor U1458 (N_1458,N_839,N_778);
nand U1459 (N_1459,N_996,N_847);
or U1460 (N_1460,N_932,N_849);
and U1461 (N_1461,N_754,N_570);
xor U1462 (N_1462,N_797,N_996);
nor U1463 (N_1463,N_785,N_991);
and U1464 (N_1464,N_513,N_946);
and U1465 (N_1465,N_793,N_631);
nand U1466 (N_1466,N_726,N_630);
or U1467 (N_1467,N_598,N_943);
or U1468 (N_1468,N_642,N_501);
nand U1469 (N_1469,N_557,N_854);
or U1470 (N_1470,N_584,N_965);
nand U1471 (N_1471,N_967,N_577);
or U1472 (N_1472,N_850,N_688);
nand U1473 (N_1473,N_503,N_789);
or U1474 (N_1474,N_545,N_887);
or U1475 (N_1475,N_772,N_760);
nand U1476 (N_1476,N_930,N_829);
and U1477 (N_1477,N_574,N_691);
xnor U1478 (N_1478,N_992,N_537);
nand U1479 (N_1479,N_930,N_563);
or U1480 (N_1480,N_819,N_509);
nor U1481 (N_1481,N_508,N_659);
nand U1482 (N_1482,N_565,N_634);
and U1483 (N_1483,N_952,N_704);
nand U1484 (N_1484,N_998,N_728);
or U1485 (N_1485,N_807,N_901);
nor U1486 (N_1486,N_890,N_654);
nor U1487 (N_1487,N_765,N_931);
nand U1488 (N_1488,N_962,N_924);
nand U1489 (N_1489,N_706,N_647);
and U1490 (N_1490,N_841,N_753);
nor U1491 (N_1491,N_716,N_572);
xnor U1492 (N_1492,N_961,N_547);
or U1493 (N_1493,N_843,N_580);
nand U1494 (N_1494,N_922,N_695);
and U1495 (N_1495,N_605,N_868);
or U1496 (N_1496,N_620,N_549);
and U1497 (N_1497,N_996,N_648);
nand U1498 (N_1498,N_726,N_517);
or U1499 (N_1499,N_631,N_952);
nand U1500 (N_1500,N_1217,N_1440);
nor U1501 (N_1501,N_1020,N_1302);
xor U1502 (N_1502,N_1175,N_1163);
xor U1503 (N_1503,N_1180,N_1033);
and U1504 (N_1504,N_1077,N_1414);
nor U1505 (N_1505,N_1465,N_1203);
nand U1506 (N_1506,N_1073,N_1116);
nand U1507 (N_1507,N_1338,N_1395);
nor U1508 (N_1508,N_1131,N_1025);
nand U1509 (N_1509,N_1426,N_1165);
nand U1510 (N_1510,N_1321,N_1167);
or U1511 (N_1511,N_1053,N_1254);
and U1512 (N_1512,N_1011,N_1392);
nor U1513 (N_1513,N_1168,N_1119);
nand U1514 (N_1514,N_1322,N_1200);
or U1515 (N_1515,N_1120,N_1140);
and U1516 (N_1516,N_1156,N_1087);
nand U1517 (N_1517,N_1027,N_1271);
nor U1518 (N_1518,N_1155,N_1458);
and U1519 (N_1519,N_1037,N_1422);
nor U1520 (N_1520,N_1022,N_1247);
and U1521 (N_1521,N_1491,N_1361);
and U1522 (N_1522,N_1333,N_1295);
nor U1523 (N_1523,N_1215,N_1189);
and U1524 (N_1524,N_1026,N_1249);
or U1525 (N_1525,N_1086,N_1258);
nand U1526 (N_1526,N_1287,N_1107);
nor U1527 (N_1527,N_1494,N_1446);
or U1528 (N_1528,N_1473,N_1190);
nor U1529 (N_1529,N_1083,N_1010);
xor U1530 (N_1530,N_1496,N_1472);
and U1531 (N_1531,N_1490,N_1476);
and U1532 (N_1532,N_1199,N_1242);
nor U1533 (N_1533,N_1363,N_1207);
or U1534 (N_1534,N_1412,N_1463);
or U1535 (N_1535,N_1263,N_1124);
and U1536 (N_1536,N_1223,N_1157);
or U1537 (N_1537,N_1283,N_1404);
nor U1538 (N_1538,N_1499,N_1164);
or U1539 (N_1539,N_1014,N_1405);
and U1540 (N_1540,N_1208,N_1015);
nand U1541 (N_1541,N_1046,N_1234);
and U1542 (N_1542,N_1291,N_1311);
nor U1543 (N_1543,N_1399,N_1008);
or U1544 (N_1544,N_1276,N_1471);
nand U1545 (N_1545,N_1421,N_1103);
and U1546 (N_1546,N_1130,N_1147);
xor U1547 (N_1547,N_1460,N_1062);
nor U1548 (N_1548,N_1218,N_1349);
nand U1549 (N_1549,N_1019,N_1032);
and U1550 (N_1550,N_1100,N_1277);
or U1551 (N_1551,N_1372,N_1076);
and U1552 (N_1552,N_1005,N_1052);
nand U1553 (N_1553,N_1143,N_1396);
xor U1554 (N_1554,N_1160,N_1371);
and U1555 (N_1555,N_1012,N_1159);
nand U1556 (N_1556,N_1330,N_1222);
or U1557 (N_1557,N_1174,N_1357);
nor U1558 (N_1558,N_1031,N_1121);
or U1559 (N_1559,N_1055,N_1452);
nand U1560 (N_1560,N_1331,N_1497);
nor U1561 (N_1561,N_1065,N_1334);
nand U1562 (N_1562,N_1265,N_1098);
nor U1563 (N_1563,N_1398,N_1063);
and U1564 (N_1564,N_1042,N_1213);
nand U1565 (N_1565,N_1043,N_1454);
nor U1566 (N_1566,N_1212,N_1264);
nand U1567 (N_1567,N_1191,N_1113);
or U1568 (N_1568,N_1224,N_1352);
nor U1569 (N_1569,N_1112,N_1072);
or U1570 (N_1570,N_1133,N_1319);
or U1571 (N_1571,N_1182,N_1003);
nor U1572 (N_1572,N_1381,N_1050);
nand U1573 (N_1573,N_1006,N_1420);
xor U1574 (N_1574,N_1016,N_1141);
nand U1575 (N_1575,N_1267,N_1314);
nand U1576 (N_1576,N_1369,N_1275);
xor U1577 (N_1577,N_1281,N_1296);
or U1578 (N_1578,N_1248,N_1091);
nand U1579 (N_1579,N_1235,N_1310);
and U1580 (N_1580,N_1344,N_1188);
or U1581 (N_1581,N_1469,N_1244);
or U1582 (N_1582,N_1057,N_1260);
nor U1583 (N_1583,N_1435,N_1114);
and U1584 (N_1584,N_1362,N_1045);
nand U1585 (N_1585,N_1197,N_1401);
or U1586 (N_1586,N_1122,N_1376);
and U1587 (N_1587,N_1332,N_1000);
nor U1588 (N_1588,N_1092,N_1434);
or U1589 (N_1589,N_1255,N_1444);
or U1590 (N_1590,N_1206,N_1245);
xor U1591 (N_1591,N_1464,N_1241);
xnor U1592 (N_1592,N_1101,N_1411);
nand U1593 (N_1593,N_1198,N_1339);
nand U1594 (N_1594,N_1436,N_1298);
nand U1595 (N_1595,N_1451,N_1088);
and U1596 (N_1596,N_1109,N_1445);
xnor U1597 (N_1597,N_1069,N_1278);
nand U1598 (N_1598,N_1068,N_1232);
and U1599 (N_1599,N_1407,N_1138);
or U1600 (N_1600,N_1002,N_1024);
nor U1601 (N_1601,N_1326,N_1410);
nand U1602 (N_1602,N_1423,N_1177);
nor U1603 (N_1603,N_1450,N_1489);
or U1604 (N_1604,N_1449,N_1316);
nand U1605 (N_1605,N_1104,N_1237);
nand U1606 (N_1606,N_1300,N_1383);
nand U1607 (N_1607,N_1226,N_1134);
nand U1608 (N_1608,N_1253,N_1181);
nor U1609 (N_1609,N_1468,N_1129);
or U1610 (N_1610,N_1406,N_1259);
xnor U1611 (N_1611,N_1150,N_1048);
nand U1612 (N_1612,N_1211,N_1195);
nor U1613 (N_1613,N_1061,N_1257);
or U1614 (N_1614,N_1428,N_1419);
nor U1615 (N_1615,N_1183,N_1418);
and U1616 (N_1616,N_1059,N_1485);
nand U1617 (N_1617,N_1236,N_1082);
or U1618 (N_1618,N_1161,N_1273);
and U1619 (N_1619,N_1313,N_1417);
nand U1620 (N_1620,N_1151,N_1408);
nor U1621 (N_1621,N_1397,N_1096);
and U1622 (N_1622,N_1379,N_1293);
xor U1623 (N_1623,N_1488,N_1359);
xnor U1624 (N_1624,N_1290,N_1243);
nor U1625 (N_1625,N_1102,N_1060);
xor U1626 (N_1626,N_1084,N_1368);
nand U1627 (N_1627,N_1162,N_1013);
nor U1628 (N_1628,N_1185,N_1184);
nand U1629 (N_1629,N_1149,N_1474);
or U1630 (N_1630,N_1345,N_1085);
xor U1631 (N_1631,N_1374,N_1145);
or U1632 (N_1632,N_1400,N_1353);
nor U1633 (N_1633,N_1301,N_1481);
nor U1634 (N_1634,N_1461,N_1336);
nand U1635 (N_1635,N_1158,N_1169);
xor U1636 (N_1636,N_1038,N_1486);
or U1637 (N_1637,N_1036,N_1106);
and U1638 (N_1638,N_1456,N_1393);
nand U1639 (N_1639,N_1308,N_1462);
nand U1640 (N_1640,N_1210,N_1239);
nand U1641 (N_1641,N_1443,N_1288);
xor U1642 (N_1642,N_1035,N_1403);
xnor U1643 (N_1643,N_1146,N_1152);
or U1644 (N_1644,N_1266,N_1023);
or U1645 (N_1645,N_1386,N_1094);
or U1646 (N_1646,N_1268,N_1179);
and U1647 (N_1647,N_1216,N_1347);
or U1648 (N_1648,N_1039,N_1108);
or U1649 (N_1649,N_1303,N_1274);
nand U1650 (N_1650,N_1166,N_1367);
nor U1651 (N_1651,N_1132,N_1327);
nand U1652 (N_1652,N_1186,N_1390);
nor U1653 (N_1653,N_1312,N_1432);
xor U1654 (N_1654,N_1172,N_1009);
xor U1655 (N_1655,N_1286,N_1279);
and U1656 (N_1656,N_1227,N_1378);
and U1657 (N_1657,N_1343,N_1095);
and U1658 (N_1658,N_1079,N_1252);
or U1659 (N_1659,N_1358,N_1261);
nand U1660 (N_1660,N_1029,N_1136);
xnor U1661 (N_1661,N_1453,N_1430);
or U1662 (N_1662,N_1269,N_1317);
or U1663 (N_1663,N_1297,N_1416);
or U1664 (N_1664,N_1373,N_1034);
nor U1665 (N_1665,N_1004,N_1196);
and U1666 (N_1666,N_1388,N_1135);
nor U1667 (N_1667,N_1402,N_1256);
and U1668 (N_1668,N_1480,N_1346);
and U1669 (N_1669,N_1078,N_1441);
nand U1670 (N_1670,N_1364,N_1438);
nand U1671 (N_1671,N_1071,N_1429);
nor U1672 (N_1672,N_1054,N_1051);
nor U1673 (N_1673,N_1384,N_1220);
and U1674 (N_1674,N_1115,N_1251);
nand U1675 (N_1675,N_1306,N_1292);
or U1676 (N_1676,N_1228,N_1360);
and U1677 (N_1677,N_1457,N_1173);
or U1678 (N_1678,N_1382,N_1262);
nand U1679 (N_1679,N_1204,N_1477);
and U1680 (N_1680,N_1282,N_1437);
or U1681 (N_1681,N_1044,N_1470);
nand U1682 (N_1682,N_1294,N_1105);
and U1683 (N_1683,N_1448,N_1315);
or U1684 (N_1684,N_1233,N_1118);
or U1685 (N_1685,N_1018,N_1030);
nand U1686 (N_1686,N_1056,N_1483);
nor U1687 (N_1687,N_1366,N_1093);
and U1688 (N_1688,N_1495,N_1066);
nor U1689 (N_1689,N_1041,N_1067);
or U1690 (N_1690,N_1074,N_1272);
nand U1691 (N_1691,N_1123,N_1225);
or U1692 (N_1692,N_1205,N_1467);
nand U1693 (N_1693,N_1270,N_1375);
nor U1694 (N_1694,N_1370,N_1427);
or U1695 (N_1695,N_1304,N_1219);
nor U1696 (N_1696,N_1238,N_1425);
and U1697 (N_1697,N_1340,N_1089);
nor U1698 (N_1698,N_1459,N_1335);
nor U1699 (N_1699,N_1075,N_1309);
or U1700 (N_1700,N_1028,N_1176);
or U1701 (N_1701,N_1139,N_1221);
or U1702 (N_1702,N_1127,N_1229);
nand U1703 (N_1703,N_1111,N_1493);
nand U1704 (N_1704,N_1007,N_1466);
or U1705 (N_1705,N_1389,N_1377);
and U1706 (N_1706,N_1328,N_1170);
or U1707 (N_1707,N_1341,N_1154);
or U1708 (N_1708,N_1144,N_1246);
nand U1709 (N_1709,N_1231,N_1194);
nand U1710 (N_1710,N_1413,N_1058);
nand U1711 (N_1711,N_1081,N_1351);
nand U1712 (N_1712,N_1202,N_1350);
xnor U1713 (N_1713,N_1487,N_1455);
nor U1714 (N_1714,N_1307,N_1324);
or U1715 (N_1715,N_1492,N_1070);
nand U1716 (N_1716,N_1001,N_1090);
nand U1717 (N_1717,N_1355,N_1153);
nor U1718 (N_1718,N_1178,N_1475);
nand U1719 (N_1719,N_1171,N_1320);
nor U1720 (N_1720,N_1431,N_1117);
nor U1721 (N_1721,N_1299,N_1110);
nand U1722 (N_1722,N_1442,N_1017);
and U1723 (N_1723,N_1280,N_1285);
or U1724 (N_1724,N_1447,N_1337);
nor U1725 (N_1725,N_1250,N_1214);
nand U1726 (N_1726,N_1284,N_1064);
and U1727 (N_1727,N_1148,N_1365);
nand U1728 (N_1728,N_1380,N_1192);
nor U1729 (N_1729,N_1424,N_1479);
nand U1730 (N_1730,N_1049,N_1484);
xor U1731 (N_1731,N_1209,N_1498);
nor U1732 (N_1732,N_1342,N_1482);
nor U1733 (N_1733,N_1125,N_1394);
nand U1734 (N_1734,N_1128,N_1409);
nor U1735 (N_1735,N_1356,N_1305);
nand U1736 (N_1736,N_1325,N_1348);
or U1737 (N_1737,N_1040,N_1354);
nor U1738 (N_1738,N_1433,N_1099);
nor U1739 (N_1739,N_1240,N_1126);
and U1740 (N_1740,N_1329,N_1137);
or U1741 (N_1741,N_1097,N_1230);
nor U1742 (N_1742,N_1478,N_1323);
nand U1743 (N_1743,N_1187,N_1391);
or U1744 (N_1744,N_1193,N_1021);
and U1745 (N_1745,N_1387,N_1289);
nor U1746 (N_1746,N_1385,N_1415);
nand U1747 (N_1747,N_1318,N_1142);
nand U1748 (N_1748,N_1201,N_1439);
nor U1749 (N_1749,N_1080,N_1047);
and U1750 (N_1750,N_1259,N_1481);
or U1751 (N_1751,N_1393,N_1054);
and U1752 (N_1752,N_1457,N_1470);
nor U1753 (N_1753,N_1182,N_1474);
or U1754 (N_1754,N_1236,N_1146);
nor U1755 (N_1755,N_1276,N_1317);
nor U1756 (N_1756,N_1354,N_1177);
nor U1757 (N_1757,N_1118,N_1054);
or U1758 (N_1758,N_1279,N_1398);
nor U1759 (N_1759,N_1031,N_1187);
or U1760 (N_1760,N_1228,N_1402);
nor U1761 (N_1761,N_1254,N_1218);
nor U1762 (N_1762,N_1317,N_1421);
and U1763 (N_1763,N_1211,N_1076);
nor U1764 (N_1764,N_1282,N_1241);
and U1765 (N_1765,N_1081,N_1242);
xor U1766 (N_1766,N_1206,N_1469);
or U1767 (N_1767,N_1227,N_1246);
nand U1768 (N_1768,N_1215,N_1327);
or U1769 (N_1769,N_1361,N_1486);
nor U1770 (N_1770,N_1276,N_1483);
and U1771 (N_1771,N_1173,N_1463);
or U1772 (N_1772,N_1455,N_1258);
and U1773 (N_1773,N_1271,N_1205);
or U1774 (N_1774,N_1186,N_1041);
or U1775 (N_1775,N_1359,N_1445);
or U1776 (N_1776,N_1267,N_1202);
or U1777 (N_1777,N_1418,N_1375);
nor U1778 (N_1778,N_1485,N_1251);
and U1779 (N_1779,N_1466,N_1376);
and U1780 (N_1780,N_1188,N_1278);
nand U1781 (N_1781,N_1291,N_1023);
and U1782 (N_1782,N_1440,N_1398);
nor U1783 (N_1783,N_1424,N_1126);
and U1784 (N_1784,N_1385,N_1042);
or U1785 (N_1785,N_1064,N_1183);
nor U1786 (N_1786,N_1414,N_1158);
xor U1787 (N_1787,N_1458,N_1193);
or U1788 (N_1788,N_1422,N_1336);
and U1789 (N_1789,N_1217,N_1080);
and U1790 (N_1790,N_1364,N_1288);
or U1791 (N_1791,N_1003,N_1028);
nor U1792 (N_1792,N_1277,N_1147);
or U1793 (N_1793,N_1261,N_1414);
or U1794 (N_1794,N_1298,N_1475);
nand U1795 (N_1795,N_1041,N_1289);
or U1796 (N_1796,N_1163,N_1372);
and U1797 (N_1797,N_1234,N_1051);
or U1798 (N_1798,N_1423,N_1418);
and U1799 (N_1799,N_1286,N_1117);
nand U1800 (N_1800,N_1490,N_1023);
or U1801 (N_1801,N_1223,N_1280);
and U1802 (N_1802,N_1203,N_1158);
or U1803 (N_1803,N_1369,N_1250);
nor U1804 (N_1804,N_1464,N_1192);
nor U1805 (N_1805,N_1066,N_1362);
or U1806 (N_1806,N_1455,N_1215);
nor U1807 (N_1807,N_1475,N_1120);
xnor U1808 (N_1808,N_1018,N_1012);
xor U1809 (N_1809,N_1474,N_1063);
nor U1810 (N_1810,N_1293,N_1151);
or U1811 (N_1811,N_1375,N_1134);
or U1812 (N_1812,N_1226,N_1241);
nand U1813 (N_1813,N_1084,N_1066);
and U1814 (N_1814,N_1407,N_1154);
xor U1815 (N_1815,N_1479,N_1015);
nor U1816 (N_1816,N_1172,N_1349);
xor U1817 (N_1817,N_1419,N_1064);
nor U1818 (N_1818,N_1328,N_1337);
and U1819 (N_1819,N_1242,N_1339);
xor U1820 (N_1820,N_1160,N_1434);
or U1821 (N_1821,N_1471,N_1205);
nor U1822 (N_1822,N_1039,N_1319);
and U1823 (N_1823,N_1440,N_1396);
nor U1824 (N_1824,N_1195,N_1053);
and U1825 (N_1825,N_1441,N_1049);
nand U1826 (N_1826,N_1370,N_1094);
or U1827 (N_1827,N_1450,N_1188);
xor U1828 (N_1828,N_1117,N_1129);
nor U1829 (N_1829,N_1245,N_1080);
or U1830 (N_1830,N_1435,N_1248);
or U1831 (N_1831,N_1338,N_1239);
nor U1832 (N_1832,N_1149,N_1143);
nand U1833 (N_1833,N_1110,N_1470);
and U1834 (N_1834,N_1046,N_1433);
nand U1835 (N_1835,N_1248,N_1085);
and U1836 (N_1836,N_1068,N_1492);
xor U1837 (N_1837,N_1380,N_1462);
nand U1838 (N_1838,N_1013,N_1430);
and U1839 (N_1839,N_1423,N_1238);
or U1840 (N_1840,N_1216,N_1287);
and U1841 (N_1841,N_1085,N_1401);
nand U1842 (N_1842,N_1221,N_1202);
nand U1843 (N_1843,N_1396,N_1433);
and U1844 (N_1844,N_1174,N_1046);
nand U1845 (N_1845,N_1230,N_1495);
nand U1846 (N_1846,N_1454,N_1268);
xnor U1847 (N_1847,N_1401,N_1475);
and U1848 (N_1848,N_1259,N_1460);
xor U1849 (N_1849,N_1498,N_1451);
nand U1850 (N_1850,N_1079,N_1341);
nor U1851 (N_1851,N_1187,N_1318);
or U1852 (N_1852,N_1020,N_1080);
nand U1853 (N_1853,N_1079,N_1259);
nand U1854 (N_1854,N_1482,N_1380);
or U1855 (N_1855,N_1039,N_1443);
xnor U1856 (N_1856,N_1284,N_1147);
and U1857 (N_1857,N_1106,N_1245);
or U1858 (N_1858,N_1290,N_1088);
and U1859 (N_1859,N_1229,N_1488);
nand U1860 (N_1860,N_1427,N_1071);
nor U1861 (N_1861,N_1067,N_1383);
and U1862 (N_1862,N_1038,N_1477);
or U1863 (N_1863,N_1088,N_1432);
and U1864 (N_1864,N_1406,N_1301);
nor U1865 (N_1865,N_1495,N_1076);
nor U1866 (N_1866,N_1119,N_1152);
nor U1867 (N_1867,N_1478,N_1436);
xnor U1868 (N_1868,N_1386,N_1417);
nand U1869 (N_1869,N_1027,N_1181);
and U1870 (N_1870,N_1474,N_1315);
xnor U1871 (N_1871,N_1273,N_1460);
nor U1872 (N_1872,N_1427,N_1011);
nor U1873 (N_1873,N_1058,N_1087);
or U1874 (N_1874,N_1268,N_1465);
nand U1875 (N_1875,N_1285,N_1423);
or U1876 (N_1876,N_1107,N_1362);
or U1877 (N_1877,N_1283,N_1036);
xor U1878 (N_1878,N_1026,N_1180);
xnor U1879 (N_1879,N_1284,N_1316);
nand U1880 (N_1880,N_1274,N_1173);
nor U1881 (N_1881,N_1085,N_1145);
nand U1882 (N_1882,N_1307,N_1122);
nor U1883 (N_1883,N_1449,N_1247);
xor U1884 (N_1884,N_1138,N_1335);
nand U1885 (N_1885,N_1052,N_1369);
and U1886 (N_1886,N_1445,N_1443);
nand U1887 (N_1887,N_1432,N_1136);
or U1888 (N_1888,N_1467,N_1262);
nand U1889 (N_1889,N_1200,N_1009);
and U1890 (N_1890,N_1069,N_1048);
xor U1891 (N_1891,N_1386,N_1209);
nor U1892 (N_1892,N_1272,N_1284);
or U1893 (N_1893,N_1456,N_1090);
nand U1894 (N_1894,N_1136,N_1275);
nand U1895 (N_1895,N_1320,N_1279);
and U1896 (N_1896,N_1277,N_1023);
and U1897 (N_1897,N_1303,N_1014);
or U1898 (N_1898,N_1056,N_1445);
xnor U1899 (N_1899,N_1221,N_1416);
nor U1900 (N_1900,N_1155,N_1154);
or U1901 (N_1901,N_1481,N_1308);
nand U1902 (N_1902,N_1124,N_1285);
and U1903 (N_1903,N_1150,N_1487);
or U1904 (N_1904,N_1075,N_1206);
nand U1905 (N_1905,N_1354,N_1200);
and U1906 (N_1906,N_1282,N_1308);
and U1907 (N_1907,N_1250,N_1026);
xnor U1908 (N_1908,N_1174,N_1210);
nand U1909 (N_1909,N_1337,N_1028);
xor U1910 (N_1910,N_1057,N_1032);
or U1911 (N_1911,N_1210,N_1429);
nor U1912 (N_1912,N_1280,N_1439);
or U1913 (N_1913,N_1354,N_1459);
nand U1914 (N_1914,N_1485,N_1393);
nand U1915 (N_1915,N_1079,N_1354);
nor U1916 (N_1916,N_1098,N_1154);
nor U1917 (N_1917,N_1110,N_1369);
and U1918 (N_1918,N_1030,N_1447);
nand U1919 (N_1919,N_1380,N_1245);
xor U1920 (N_1920,N_1034,N_1139);
nor U1921 (N_1921,N_1400,N_1451);
nand U1922 (N_1922,N_1227,N_1239);
or U1923 (N_1923,N_1356,N_1498);
nand U1924 (N_1924,N_1253,N_1467);
nor U1925 (N_1925,N_1193,N_1361);
or U1926 (N_1926,N_1274,N_1266);
or U1927 (N_1927,N_1024,N_1307);
nor U1928 (N_1928,N_1315,N_1204);
and U1929 (N_1929,N_1462,N_1000);
nor U1930 (N_1930,N_1129,N_1021);
nand U1931 (N_1931,N_1100,N_1373);
and U1932 (N_1932,N_1287,N_1153);
xnor U1933 (N_1933,N_1372,N_1386);
nor U1934 (N_1934,N_1358,N_1276);
nand U1935 (N_1935,N_1068,N_1103);
or U1936 (N_1936,N_1110,N_1048);
and U1937 (N_1937,N_1125,N_1354);
nor U1938 (N_1938,N_1141,N_1477);
and U1939 (N_1939,N_1152,N_1479);
nor U1940 (N_1940,N_1189,N_1453);
or U1941 (N_1941,N_1357,N_1382);
and U1942 (N_1942,N_1444,N_1281);
nor U1943 (N_1943,N_1230,N_1019);
or U1944 (N_1944,N_1442,N_1481);
and U1945 (N_1945,N_1286,N_1150);
nand U1946 (N_1946,N_1349,N_1045);
xnor U1947 (N_1947,N_1388,N_1449);
nor U1948 (N_1948,N_1009,N_1004);
nor U1949 (N_1949,N_1490,N_1105);
nand U1950 (N_1950,N_1468,N_1481);
or U1951 (N_1951,N_1231,N_1214);
and U1952 (N_1952,N_1423,N_1291);
xnor U1953 (N_1953,N_1496,N_1125);
nor U1954 (N_1954,N_1459,N_1431);
and U1955 (N_1955,N_1145,N_1187);
or U1956 (N_1956,N_1495,N_1187);
nor U1957 (N_1957,N_1097,N_1471);
or U1958 (N_1958,N_1038,N_1376);
xor U1959 (N_1959,N_1247,N_1413);
and U1960 (N_1960,N_1105,N_1150);
and U1961 (N_1961,N_1408,N_1313);
nand U1962 (N_1962,N_1064,N_1156);
nor U1963 (N_1963,N_1439,N_1332);
or U1964 (N_1964,N_1391,N_1250);
or U1965 (N_1965,N_1158,N_1140);
nand U1966 (N_1966,N_1295,N_1451);
or U1967 (N_1967,N_1335,N_1472);
and U1968 (N_1968,N_1001,N_1357);
nor U1969 (N_1969,N_1428,N_1413);
nor U1970 (N_1970,N_1415,N_1280);
or U1971 (N_1971,N_1457,N_1040);
nor U1972 (N_1972,N_1400,N_1307);
or U1973 (N_1973,N_1297,N_1021);
nor U1974 (N_1974,N_1356,N_1446);
and U1975 (N_1975,N_1418,N_1205);
nor U1976 (N_1976,N_1092,N_1282);
nand U1977 (N_1977,N_1298,N_1163);
xnor U1978 (N_1978,N_1017,N_1206);
xnor U1979 (N_1979,N_1375,N_1490);
nor U1980 (N_1980,N_1006,N_1417);
and U1981 (N_1981,N_1190,N_1067);
nand U1982 (N_1982,N_1469,N_1376);
nor U1983 (N_1983,N_1038,N_1176);
nor U1984 (N_1984,N_1246,N_1081);
nand U1985 (N_1985,N_1298,N_1344);
nand U1986 (N_1986,N_1136,N_1238);
nand U1987 (N_1987,N_1336,N_1272);
nand U1988 (N_1988,N_1396,N_1176);
or U1989 (N_1989,N_1023,N_1401);
xor U1990 (N_1990,N_1156,N_1493);
nand U1991 (N_1991,N_1095,N_1127);
nor U1992 (N_1992,N_1122,N_1382);
or U1993 (N_1993,N_1078,N_1068);
nor U1994 (N_1994,N_1166,N_1296);
and U1995 (N_1995,N_1415,N_1074);
or U1996 (N_1996,N_1051,N_1451);
nor U1997 (N_1997,N_1475,N_1349);
nand U1998 (N_1998,N_1329,N_1464);
nand U1999 (N_1999,N_1243,N_1179);
and U2000 (N_2000,N_1829,N_1596);
and U2001 (N_2001,N_1666,N_1833);
xnor U2002 (N_2002,N_1562,N_1744);
xor U2003 (N_2003,N_1836,N_1823);
xor U2004 (N_2004,N_1582,N_1825);
and U2005 (N_2005,N_1884,N_1647);
nor U2006 (N_2006,N_1940,N_1640);
nand U2007 (N_2007,N_1765,N_1660);
nor U2008 (N_2008,N_1641,N_1990);
and U2009 (N_2009,N_1594,N_1506);
nor U2010 (N_2010,N_1948,N_1897);
or U2011 (N_2011,N_1993,N_1638);
and U2012 (N_2012,N_1642,N_1720);
nor U2013 (N_2013,N_1908,N_1900);
nor U2014 (N_2014,N_1922,N_1572);
nand U2015 (N_2015,N_1709,N_1956);
nor U2016 (N_2016,N_1882,N_1529);
xnor U2017 (N_2017,N_1970,N_1799);
and U2018 (N_2018,N_1834,N_1964);
nand U2019 (N_2019,N_1869,N_1512);
or U2020 (N_2020,N_1991,N_1602);
nand U2021 (N_2021,N_1946,N_1975);
nand U2022 (N_2022,N_1910,N_1706);
nand U2023 (N_2023,N_1729,N_1757);
or U2024 (N_2024,N_1894,N_1740);
nor U2025 (N_2025,N_1508,N_1541);
nand U2026 (N_2026,N_1779,N_1983);
nor U2027 (N_2027,N_1841,N_1864);
nor U2028 (N_2028,N_1742,N_1931);
nor U2029 (N_2029,N_1892,N_1756);
and U2030 (N_2030,N_1899,N_1616);
or U2031 (N_2031,N_1760,N_1817);
nand U2032 (N_2032,N_1697,N_1873);
xnor U2033 (N_2033,N_1805,N_1618);
nor U2034 (N_2034,N_1878,N_1976);
nand U2035 (N_2035,N_1928,N_1783);
nand U2036 (N_2036,N_1868,N_1840);
nor U2037 (N_2037,N_1958,N_1608);
or U2038 (N_2038,N_1780,N_1544);
nand U2039 (N_2039,N_1587,N_1674);
nor U2040 (N_2040,N_1906,N_1717);
and U2041 (N_2041,N_1947,N_1994);
or U2042 (N_2042,N_1627,N_1902);
nand U2043 (N_2043,N_1981,N_1909);
nor U2044 (N_2044,N_1664,N_1985);
nand U2045 (N_2045,N_1764,N_1672);
or U2046 (N_2046,N_1808,N_1730);
and U2047 (N_2047,N_1723,N_1896);
nand U2048 (N_2048,N_1622,N_1826);
and U2049 (N_2049,N_1696,N_1624);
xnor U2050 (N_2050,N_1832,N_1519);
or U2051 (N_2051,N_1962,N_1790);
and U2052 (N_2052,N_1597,N_1812);
and U2053 (N_2053,N_1574,N_1901);
xor U2054 (N_2054,N_1854,N_1858);
or U2055 (N_2055,N_1754,N_1793);
or U2056 (N_2056,N_1885,N_1677);
nor U2057 (N_2057,N_1626,N_1543);
or U2058 (N_2058,N_1557,N_1540);
and U2059 (N_2059,N_1671,N_1509);
and U2060 (N_2060,N_1684,N_1546);
nor U2061 (N_2061,N_1945,N_1815);
nand U2062 (N_2062,N_1609,N_1547);
nand U2063 (N_2063,N_1707,N_1781);
or U2064 (N_2064,N_1579,N_1814);
or U2065 (N_2065,N_1569,N_1934);
and U2066 (N_2066,N_1775,N_1704);
nor U2067 (N_2067,N_1789,N_1601);
or U2068 (N_2068,N_1804,N_1986);
or U2069 (N_2069,N_1728,N_1944);
and U2070 (N_2070,N_1849,N_1860);
or U2071 (N_2071,N_1938,N_1733);
nand U2072 (N_2072,N_1558,N_1842);
or U2073 (N_2073,N_1726,N_1731);
nand U2074 (N_2074,N_1987,N_1617);
nand U2075 (N_2075,N_1911,N_1598);
nand U2076 (N_2076,N_1939,N_1693);
nand U2077 (N_2077,N_1629,N_1984);
nor U2078 (N_2078,N_1969,N_1809);
nand U2079 (N_2079,N_1980,N_1850);
nand U2080 (N_2080,N_1563,N_1917);
xor U2081 (N_2081,N_1510,N_1505);
xnor U2082 (N_2082,N_1523,N_1504);
nor U2083 (N_2083,N_1904,N_1870);
or U2084 (N_2084,N_1941,N_1737);
nand U2085 (N_2085,N_1965,N_1988);
and U2086 (N_2086,N_1857,N_1797);
nand U2087 (N_2087,N_1611,N_1971);
xnor U2088 (N_2088,N_1914,N_1634);
or U2089 (N_2089,N_1875,N_1692);
or U2090 (N_2090,N_1531,N_1932);
or U2091 (N_2091,N_1796,N_1552);
or U2092 (N_2092,N_1585,N_1708);
or U2093 (N_2093,N_1998,N_1777);
or U2094 (N_2094,N_1863,N_1856);
xor U2095 (N_2095,N_1895,N_1646);
nor U2096 (N_2096,N_1798,N_1926);
xor U2097 (N_2097,N_1620,N_1800);
xnor U2098 (N_2098,N_1636,N_1650);
xor U2099 (N_2099,N_1891,N_1514);
nor U2100 (N_2100,N_1741,N_1542);
or U2101 (N_2101,N_1559,N_1745);
and U2102 (N_2102,N_1927,N_1912);
nand U2103 (N_2103,N_1584,N_1746);
and U2104 (N_2104,N_1581,N_1528);
nor U2105 (N_2105,N_1679,N_1643);
nor U2106 (N_2106,N_1853,N_1535);
and U2107 (N_2107,N_1923,N_1652);
and U2108 (N_2108,N_1950,N_1517);
nor U2109 (N_2109,N_1951,N_1577);
nor U2110 (N_2110,N_1952,N_1632);
xnor U2111 (N_2111,N_1607,N_1963);
xor U2112 (N_2112,N_1921,N_1802);
nand U2113 (N_2113,N_1848,N_1669);
or U2114 (N_2114,N_1750,N_1689);
xor U2115 (N_2115,N_1888,N_1773);
and U2116 (N_2116,N_1877,N_1612);
xor U2117 (N_2117,N_1893,N_1545);
or U2118 (N_2118,N_1661,N_1644);
and U2119 (N_2119,N_1819,N_1683);
and U2120 (N_2120,N_1957,N_1699);
and U2121 (N_2121,N_1516,N_1645);
or U2122 (N_2122,N_1924,N_1682);
nor U2123 (N_2123,N_1623,N_1613);
nor U2124 (N_2124,N_1806,N_1735);
and U2125 (N_2125,N_1759,N_1871);
xnor U2126 (N_2126,N_1816,N_1883);
nand U2127 (N_2127,N_1913,N_1656);
and U2128 (N_2128,N_1747,N_1734);
nand U2129 (N_2129,N_1570,N_1515);
xor U2130 (N_2130,N_1567,N_1818);
nor U2131 (N_2131,N_1979,N_1943);
nand U2132 (N_2132,N_1560,N_1678);
nand U2133 (N_2133,N_1905,N_1791);
or U2134 (N_2134,N_1530,N_1968);
xnor U2135 (N_2135,N_1992,N_1821);
and U2136 (N_2136,N_1625,N_1782);
nor U2137 (N_2137,N_1725,N_1880);
nand U2138 (N_2138,N_1847,N_1503);
nor U2139 (N_2139,N_1628,N_1722);
nor U2140 (N_2140,N_1554,N_1568);
or U2141 (N_2141,N_1500,N_1807);
and U2142 (N_2142,N_1685,N_1604);
or U2143 (N_2143,N_1691,N_1556);
and U2144 (N_2144,N_1845,N_1936);
or U2145 (N_2145,N_1942,N_1997);
or U2146 (N_2146,N_1758,N_1698);
nand U2147 (N_2147,N_1989,N_1837);
nor U2148 (N_2148,N_1710,N_1959);
or U2149 (N_2149,N_1724,N_1778);
or U2150 (N_2150,N_1824,N_1866);
or U2151 (N_2151,N_1960,N_1865);
and U2152 (N_2152,N_1953,N_1787);
nand U2153 (N_2153,N_1614,N_1839);
nor U2154 (N_2154,N_1580,N_1658);
nand U2155 (N_2155,N_1527,N_1651);
nor U2156 (N_2156,N_1772,N_1835);
nand U2157 (N_2157,N_1606,N_1846);
or U2158 (N_2158,N_1811,N_1955);
nor U2159 (N_2159,N_1702,N_1767);
nand U2160 (N_2160,N_1524,N_1705);
xnor U2161 (N_2161,N_1967,N_1714);
or U2162 (N_2162,N_1716,N_1501);
nand U2163 (N_2163,N_1550,N_1694);
and U2164 (N_2164,N_1820,N_1933);
nand U2165 (N_2165,N_1879,N_1571);
xnor U2166 (N_2166,N_1859,N_1553);
and U2167 (N_2167,N_1507,N_1827);
and U2168 (N_2168,N_1565,N_1768);
nor U2169 (N_2169,N_1522,N_1748);
nor U2170 (N_2170,N_1751,N_1794);
and U2171 (N_2171,N_1862,N_1536);
nand U2172 (N_2172,N_1639,N_1551);
nor U2173 (N_2173,N_1851,N_1762);
xor U2174 (N_2174,N_1534,N_1637);
xnor U2175 (N_2175,N_1513,N_1686);
nor U2176 (N_2176,N_1890,N_1649);
nand U2177 (N_2177,N_1761,N_1907);
nand U2178 (N_2178,N_1813,N_1786);
nand U2179 (N_2179,N_1918,N_1518);
and U2180 (N_2180,N_1681,N_1855);
xor U2181 (N_2181,N_1874,N_1738);
nand U2182 (N_2182,N_1715,N_1603);
nor U2183 (N_2183,N_1999,N_1774);
and U2184 (N_2184,N_1954,N_1776);
or U2185 (N_2185,N_1920,N_1511);
or U2186 (N_2186,N_1935,N_1831);
and U2187 (N_2187,N_1872,N_1752);
nand U2188 (N_2188,N_1695,N_1667);
or U2189 (N_2189,N_1668,N_1784);
nand U2190 (N_2190,N_1600,N_1919);
nor U2191 (N_2191,N_1732,N_1785);
and U2192 (N_2192,N_1711,N_1949);
and U2193 (N_2193,N_1770,N_1591);
nand U2194 (N_2194,N_1593,N_1803);
xor U2195 (N_2195,N_1903,N_1749);
nor U2196 (N_2196,N_1595,N_1727);
or U2197 (N_2197,N_1838,N_1532);
and U2198 (N_2198,N_1564,N_1755);
and U2199 (N_2199,N_1887,N_1599);
and U2200 (N_2200,N_1937,N_1712);
nand U2201 (N_2201,N_1589,N_1700);
and U2202 (N_2202,N_1788,N_1801);
and U2203 (N_2203,N_1713,N_1844);
nor U2204 (N_2204,N_1659,N_1619);
or U2205 (N_2205,N_1586,N_1578);
and U2206 (N_2206,N_1592,N_1654);
nor U2207 (N_2207,N_1548,N_1615);
nor U2208 (N_2208,N_1655,N_1526);
nand U2209 (N_2209,N_1867,N_1718);
nor U2210 (N_2210,N_1561,N_1843);
or U2211 (N_2211,N_1771,N_1690);
nor U2212 (N_2212,N_1573,N_1974);
or U2213 (N_2213,N_1670,N_1743);
and U2214 (N_2214,N_1898,N_1538);
nor U2215 (N_2215,N_1566,N_1889);
and U2216 (N_2216,N_1657,N_1810);
and U2217 (N_2217,N_1972,N_1703);
nand U2218 (N_2218,N_1995,N_1621);
or U2219 (N_2219,N_1576,N_1525);
or U2220 (N_2220,N_1916,N_1630);
or U2221 (N_2221,N_1753,N_1830);
nand U2222 (N_2222,N_1583,N_1588);
or U2223 (N_2223,N_1721,N_1828);
nand U2224 (N_2224,N_1886,N_1605);
nand U2225 (N_2225,N_1533,N_1687);
nor U2226 (N_2226,N_1739,N_1549);
and U2227 (N_2227,N_1653,N_1766);
xnor U2228 (N_2228,N_1881,N_1736);
and U2229 (N_2229,N_1610,N_1633);
or U2230 (N_2230,N_1680,N_1631);
and U2231 (N_2231,N_1795,N_1701);
nor U2232 (N_2232,N_1915,N_1978);
or U2233 (N_2233,N_1590,N_1861);
and U2234 (N_2234,N_1648,N_1676);
and U2235 (N_2235,N_1520,N_1663);
or U2236 (N_2236,N_1982,N_1635);
nor U2237 (N_2237,N_1977,N_1675);
and U2238 (N_2238,N_1688,N_1665);
and U2239 (N_2239,N_1769,N_1662);
and U2240 (N_2240,N_1719,N_1876);
nor U2241 (N_2241,N_1539,N_1502);
nand U2242 (N_2242,N_1961,N_1930);
xor U2243 (N_2243,N_1673,N_1925);
xnor U2244 (N_2244,N_1537,N_1852);
and U2245 (N_2245,N_1966,N_1521);
and U2246 (N_2246,N_1822,N_1973);
and U2247 (N_2247,N_1792,N_1575);
and U2248 (N_2248,N_1763,N_1929);
nor U2249 (N_2249,N_1555,N_1996);
nor U2250 (N_2250,N_1814,N_1596);
nor U2251 (N_2251,N_1922,N_1706);
nor U2252 (N_2252,N_1938,N_1508);
nand U2253 (N_2253,N_1852,N_1656);
or U2254 (N_2254,N_1925,N_1931);
nor U2255 (N_2255,N_1720,N_1546);
nand U2256 (N_2256,N_1919,N_1936);
nand U2257 (N_2257,N_1734,N_1918);
nand U2258 (N_2258,N_1961,N_1555);
or U2259 (N_2259,N_1722,N_1506);
and U2260 (N_2260,N_1769,N_1573);
nand U2261 (N_2261,N_1757,N_1709);
nor U2262 (N_2262,N_1569,N_1618);
and U2263 (N_2263,N_1873,N_1748);
and U2264 (N_2264,N_1653,N_1623);
nor U2265 (N_2265,N_1667,N_1528);
and U2266 (N_2266,N_1511,N_1998);
or U2267 (N_2267,N_1710,N_1820);
nor U2268 (N_2268,N_1500,N_1521);
nor U2269 (N_2269,N_1809,N_1976);
and U2270 (N_2270,N_1702,N_1891);
and U2271 (N_2271,N_1669,N_1699);
nor U2272 (N_2272,N_1603,N_1526);
nor U2273 (N_2273,N_1696,N_1980);
xor U2274 (N_2274,N_1724,N_1879);
nand U2275 (N_2275,N_1781,N_1599);
nand U2276 (N_2276,N_1698,N_1729);
nor U2277 (N_2277,N_1970,N_1813);
nor U2278 (N_2278,N_1814,N_1611);
and U2279 (N_2279,N_1751,N_1775);
nand U2280 (N_2280,N_1574,N_1866);
and U2281 (N_2281,N_1978,N_1590);
or U2282 (N_2282,N_1546,N_1545);
nor U2283 (N_2283,N_1820,N_1757);
nand U2284 (N_2284,N_1731,N_1572);
and U2285 (N_2285,N_1673,N_1969);
and U2286 (N_2286,N_1765,N_1931);
and U2287 (N_2287,N_1812,N_1750);
nor U2288 (N_2288,N_1997,N_1706);
or U2289 (N_2289,N_1617,N_1638);
xnor U2290 (N_2290,N_1892,N_1500);
nor U2291 (N_2291,N_1505,N_1642);
nor U2292 (N_2292,N_1517,N_1989);
and U2293 (N_2293,N_1522,N_1930);
nor U2294 (N_2294,N_1894,N_1931);
and U2295 (N_2295,N_1617,N_1785);
nor U2296 (N_2296,N_1869,N_1831);
and U2297 (N_2297,N_1871,N_1843);
or U2298 (N_2298,N_1561,N_1507);
nand U2299 (N_2299,N_1599,N_1646);
and U2300 (N_2300,N_1899,N_1686);
or U2301 (N_2301,N_1512,N_1604);
nor U2302 (N_2302,N_1726,N_1782);
nand U2303 (N_2303,N_1762,N_1819);
and U2304 (N_2304,N_1540,N_1751);
nand U2305 (N_2305,N_1731,N_1552);
nor U2306 (N_2306,N_1873,N_1761);
and U2307 (N_2307,N_1707,N_1853);
xor U2308 (N_2308,N_1816,N_1642);
nor U2309 (N_2309,N_1805,N_1848);
or U2310 (N_2310,N_1507,N_1514);
xor U2311 (N_2311,N_1817,N_1715);
nand U2312 (N_2312,N_1789,N_1524);
or U2313 (N_2313,N_1570,N_1500);
nor U2314 (N_2314,N_1945,N_1952);
nor U2315 (N_2315,N_1977,N_1810);
nand U2316 (N_2316,N_1835,N_1667);
nor U2317 (N_2317,N_1938,N_1966);
nand U2318 (N_2318,N_1974,N_1732);
nor U2319 (N_2319,N_1823,N_1522);
or U2320 (N_2320,N_1604,N_1646);
or U2321 (N_2321,N_1949,N_1502);
and U2322 (N_2322,N_1629,N_1658);
nor U2323 (N_2323,N_1882,N_1950);
nand U2324 (N_2324,N_1558,N_1543);
xnor U2325 (N_2325,N_1553,N_1872);
nand U2326 (N_2326,N_1666,N_1554);
and U2327 (N_2327,N_1732,N_1734);
nand U2328 (N_2328,N_1914,N_1980);
nand U2329 (N_2329,N_1665,N_1726);
and U2330 (N_2330,N_1801,N_1529);
and U2331 (N_2331,N_1592,N_1958);
nand U2332 (N_2332,N_1667,N_1715);
nor U2333 (N_2333,N_1609,N_1668);
nand U2334 (N_2334,N_1646,N_1719);
or U2335 (N_2335,N_1697,N_1628);
or U2336 (N_2336,N_1622,N_1694);
nor U2337 (N_2337,N_1593,N_1752);
nand U2338 (N_2338,N_1560,N_1704);
nor U2339 (N_2339,N_1885,N_1678);
or U2340 (N_2340,N_1723,N_1516);
and U2341 (N_2341,N_1961,N_1745);
or U2342 (N_2342,N_1629,N_1833);
nor U2343 (N_2343,N_1802,N_1507);
xor U2344 (N_2344,N_1854,N_1915);
nand U2345 (N_2345,N_1687,N_1573);
and U2346 (N_2346,N_1519,N_1721);
or U2347 (N_2347,N_1751,N_1606);
nand U2348 (N_2348,N_1624,N_1795);
and U2349 (N_2349,N_1503,N_1977);
nand U2350 (N_2350,N_1508,N_1630);
and U2351 (N_2351,N_1814,N_1790);
xnor U2352 (N_2352,N_1720,N_1559);
and U2353 (N_2353,N_1824,N_1950);
and U2354 (N_2354,N_1537,N_1824);
and U2355 (N_2355,N_1937,N_1955);
nand U2356 (N_2356,N_1744,N_1568);
nand U2357 (N_2357,N_1691,N_1689);
xnor U2358 (N_2358,N_1775,N_1544);
or U2359 (N_2359,N_1955,N_1787);
and U2360 (N_2360,N_1712,N_1709);
and U2361 (N_2361,N_1538,N_1683);
nor U2362 (N_2362,N_1616,N_1617);
or U2363 (N_2363,N_1929,N_1860);
nor U2364 (N_2364,N_1829,N_1719);
and U2365 (N_2365,N_1545,N_1897);
nor U2366 (N_2366,N_1997,N_1896);
nand U2367 (N_2367,N_1717,N_1582);
and U2368 (N_2368,N_1998,N_1722);
nor U2369 (N_2369,N_1682,N_1621);
nor U2370 (N_2370,N_1800,N_1731);
and U2371 (N_2371,N_1600,N_1817);
xor U2372 (N_2372,N_1784,N_1629);
or U2373 (N_2373,N_1838,N_1952);
and U2374 (N_2374,N_1779,N_1760);
and U2375 (N_2375,N_1661,N_1625);
and U2376 (N_2376,N_1900,N_1946);
nor U2377 (N_2377,N_1937,N_1779);
nand U2378 (N_2378,N_1606,N_1775);
or U2379 (N_2379,N_1667,N_1876);
nand U2380 (N_2380,N_1595,N_1643);
and U2381 (N_2381,N_1501,N_1641);
nand U2382 (N_2382,N_1851,N_1624);
and U2383 (N_2383,N_1969,N_1727);
and U2384 (N_2384,N_1937,N_1733);
nand U2385 (N_2385,N_1655,N_1848);
nor U2386 (N_2386,N_1915,N_1615);
and U2387 (N_2387,N_1972,N_1876);
or U2388 (N_2388,N_1526,N_1809);
and U2389 (N_2389,N_1643,N_1841);
and U2390 (N_2390,N_1524,N_1776);
nand U2391 (N_2391,N_1623,N_1673);
and U2392 (N_2392,N_1886,N_1851);
nor U2393 (N_2393,N_1993,N_1718);
or U2394 (N_2394,N_1529,N_1929);
and U2395 (N_2395,N_1807,N_1609);
nand U2396 (N_2396,N_1702,N_1751);
nor U2397 (N_2397,N_1514,N_1724);
nor U2398 (N_2398,N_1802,N_1816);
or U2399 (N_2399,N_1845,N_1573);
nor U2400 (N_2400,N_1625,N_1909);
or U2401 (N_2401,N_1806,N_1748);
nor U2402 (N_2402,N_1609,N_1525);
or U2403 (N_2403,N_1658,N_1901);
or U2404 (N_2404,N_1939,N_1502);
nor U2405 (N_2405,N_1905,N_1722);
xor U2406 (N_2406,N_1943,N_1989);
nor U2407 (N_2407,N_1598,N_1742);
or U2408 (N_2408,N_1507,N_1619);
nor U2409 (N_2409,N_1577,N_1591);
nand U2410 (N_2410,N_1892,N_1718);
or U2411 (N_2411,N_1545,N_1765);
nor U2412 (N_2412,N_1929,N_1764);
xnor U2413 (N_2413,N_1681,N_1913);
and U2414 (N_2414,N_1769,N_1648);
nand U2415 (N_2415,N_1851,N_1675);
nand U2416 (N_2416,N_1777,N_1918);
nand U2417 (N_2417,N_1602,N_1953);
or U2418 (N_2418,N_1708,N_1698);
or U2419 (N_2419,N_1982,N_1814);
or U2420 (N_2420,N_1651,N_1534);
nor U2421 (N_2421,N_1790,N_1789);
xor U2422 (N_2422,N_1534,N_1896);
and U2423 (N_2423,N_1790,N_1583);
nand U2424 (N_2424,N_1749,N_1517);
and U2425 (N_2425,N_1678,N_1559);
nor U2426 (N_2426,N_1871,N_1601);
xnor U2427 (N_2427,N_1902,N_1922);
or U2428 (N_2428,N_1657,N_1716);
nor U2429 (N_2429,N_1597,N_1827);
and U2430 (N_2430,N_1918,N_1861);
nor U2431 (N_2431,N_1762,N_1796);
xnor U2432 (N_2432,N_1646,N_1500);
and U2433 (N_2433,N_1535,N_1701);
and U2434 (N_2434,N_1554,N_1897);
nand U2435 (N_2435,N_1527,N_1972);
nor U2436 (N_2436,N_1966,N_1745);
nand U2437 (N_2437,N_1801,N_1815);
or U2438 (N_2438,N_1578,N_1871);
nand U2439 (N_2439,N_1880,N_1861);
nand U2440 (N_2440,N_1635,N_1727);
and U2441 (N_2441,N_1919,N_1942);
or U2442 (N_2442,N_1757,N_1677);
or U2443 (N_2443,N_1618,N_1736);
nor U2444 (N_2444,N_1640,N_1901);
nor U2445 (N_2445,N_1966,N_1875);
or U2446 (N_2446,N_1906,N_1949);
or U2447 (N_2447,N_1846,N_1881);
nor U2448 (N_2448,N_1541,N_1544);
nor U2449 (N_2449,N_1765,N_1879);
nor U2450 (N_2450,N_1834,N_1731);
and U2451 (N_2451,N_1644,N_1786);
nand U2452 (N_2452,N_1577,N_1760);
nor U2453 (N_2453,N_1544,N_1720);
nand U2454 (N_2454,N_1619,N_1740);
or U2455 (N_2455,N_1617,N_1714);
and U2456 (N_2456,N_1876,N_1766);
and U2457 (N_2457,N_1760,N_1571);
and U2458 (N_2458,N_1703,N_1773);
nor U2459 (N_2459,N_1677,N_1884);
nand U2460 (N_2460,N_1791,N_1659);
nand U2461 (N_2461,N_1780,N_1619);
nor U2462 (N_2462,N_1639,N_1661);
or U2463 (N_2463,N_1858,N_1880);
nand U2464 (N_2464,N_1633,N_1810);
or U2465 (N_2465,N_1903,N_1844);
nor U2466 (N_2466,N_1897,N_1784);
nor U2467 (N_2467,N_1863,N_1620);
nand U2468 (N_2468,N_1799,N_1737);
nand U2469 (N_2469,N_1873,N_1732);
or U2470 (N_2470,N_1628,N_1602);
and U2471 (N_2471,N_1548,N_1569);
xnor U2472 (N_2472,N_1772,N_1872);
nor U2473 (N_2473,N_1880,N_1970);
nor U2474 (N_2474,N_1584,N_1731);
xor U2475 (N_2475,N_1583,N_1843);
xor U2476 (N_2476,N_1710,N_1899);
or U2477 (N_2477,N_1980,N_1816);
or U2478 (N_2478,N_1630,N_1584);
nor U2479 (N_2479,N_1518,N_1982);
nand U2480 (N_2480,N_1882,N_1507);
and U2481 (N_2481,N_1870,N_1649);
or U2482 (N_2482,N_1960,N_1692);
and U2483 (N_2483,N_1826,N_1671);
nand U2484 (N_2484,N_1650,N_1857);
or U2485 (N_2485,N_1559,N_1761);
nor U2486 (N_2486,N_1976,N_1558);
xor U2487 (N_2487,N_1750,N_1540);
or U2488 (N_2488,N_1994,N_1760);
or U2489 (N_2489,N_1897,N_1743);
and U2490 (N_2490,N_1812,N_1884);
nand U2491 (N_2491,N_1745,N_1692);
and U2492 (N_2492,N_1511,N_1591);
nor U2493 (N_2493,N_1578,N_1570);
and U2494 (N_2494,N_1793,N_1909);
xor U2495 (N_2495,N_1603,N_1556);
nor U2496 (N_2496,N_1741,N_1921);
and U2497 (N_2497,N_1666,N_1573);
nand U2498 (N_2498,N_1758,N_1761);
xor U2499 (N_2499,N_1517,N_1604);
nor U2500 (N_2500,N_2365,N_2420);
and U2501 (N_2501,N_2096,N_2302);
or U2502 (N_2502,N_2104,N_2268);
or U2503 (N_2503,N_2241,N_2258);
nor U2504 (N_2504,N_2423,N_2329);
or U2505 (N_2505,N_2275,N_2361);
nand U2506 (N_2506,N_2196,N_2067);
or U2507 (N_2507,N_2491,N_2102);
and U2508 (N_2508,N_2356,N_2077);
or U2509 (N_2509,N_2229,N_2364);
and U2510 (N_2510,N_2457,N_2427);
xnor U2511 (N_2511,N_2011,N_2405);
nand U2512 (N_2512,N_2023,N_2123);
nor U2513 (N_2513,N_2492,N_2377);
nor U2514 (N_2514,N_2051,N_2373);
or U2515 (N_2515,N_2108,N_2174);
nand U2516 (N_2516,N_2433,N_2130);
or U2517 (N_2517,N_2325,N_2098);
nand U2518 (N_2518,N_2199,N_2015);
and U2519 (N_2519,N_2494,N_2343);
nor U2520 (N_2520,N_2039,N_2172);
and U2521 (N_2521,N_2291,N_2063);
and U2522 (N_2522,N_2212,N_2443);
nor U2523 (N_2523,N_2103,N_2141);
nand U2524 (N_2524,N_2266,N_2370);
and U2525 (N_2525,N_2121,N_2350);
nor U2526 (N_2526,N_2340,N_2382);
nor U2527 (N_2527,N_2150,N_2088);
nor U2528 (N_2528,N_2334,N_2101);
and U2529 (N_2529,N_2024,N_2442);
nand U2530 (N_2530,N_2120,N_2287);
and U2531 (N_2531,N_2472,N_2285);
nand U2532 (N_2532,N_2134,N_2019);
and U2533 (N_2533,N_2109,N_2110);
nand U2534 (N_2534,N_2487,N_2021);
nor U2535 (N_2535,N_2425,N_2380);
and U2536 (N_2536,N_2133,N_2489);
nor U2537 (N_2537,N_2301,N_2448);
and U2538 (N_2538,N_2034,N_2005);
and U2539 (N_2539,N_2112,N_2116);
or U2540 (N_2540,N_2157,N_2195);
nor U2541 (N_2541,N_2440,N_2453);
or U2542 (N_2542,N_2310,N_2092);
or U2543 (N_2543,N_2194,N_2056);
and U2544 (N_2544,N_2068,N_2048);
or U2545 (N_2545,N_2447,N_2483);
or U2546 (N_2546,N_2144,N_2324);
nand U2547 (N_2547,N_2086,N_2428);
nor U2548 (N_2548,N_2035,N_2115);
nand U2549 (N_2549,N_2210,N_2294);
and U2550 (N_2550,N_2486,N_2126);
nand U2551 (N_2551,N_2256,N_2010);
nor U2552 (N_2552,N_2259,N_2419);
nand U2553 (N_2553,N_2255,N_2192);
nand U2554 (N_2554,N_2100,N_2244);
or U2555 (N_2555,N_2330,N_2179);
nor U2556 (N_2556,N_2284,N_2355);
and U2557 (N_2557,N_2003,N_2017);
and U2558 (N_2558,N_2185,N_2461);
or U2559 (N_2559,N_2354,N_2416);
or U2560 (N_2560,N_2471,N_2452);
xor U2561 (N_2561,N_2415,N_2243);
nor U2562 (N_2562,N_2399,N_2065);
nand U2563 (N_2563,N_2135,N_2347);
nand U2564 (N_2564,N_2280,N_2279);
nand U2565 (N_2565,N_2468,N_2082);
nor U2566 (N_2566,N_2395,N_2213);
xor U2567 (N_2567,N_2114,N_2388);
and U2568 (N_2568,N_2436,N_2352);
nor U2569 (N_2569,N_2045,N_2408);
or U2570 (N_2570,N_2136,N_2218);
and U2571 (N_2571,N_2435,N_2239);
xnor U2572 (N_2572,N_2497,N_2252);
nand U2573 (N_2573,N_2418,N_2378);
nor U2574 (N_2574,N_2083,N_2317);
nand U2575 (N_2575,N_2495,N_2000);
or U2576 (N_2576,N_2277,N_2274);
xnor U2577 (N_2577,N_2152,N_2145);
and U2578 (N_2578,N_2223,N_2234);
and U2579 (N_2579,N_2177,N_2226);
and U2580 (N_2580,N_2331,N_2214);
nor U2581 (N_2581,N_2290,N_2394);
and U2582 (N_2582,N_2374,N_2156);
or U2583 (N_2583,N_2451,N_2446);
nor U2584 (N_2584,N_2375,N_2191);
or U2585 (N_2585,N_2411,N_2128);
or U2586 (N_2586,N_2161,N_2385);
nor U2587 (N_2587,N_2160,N_2458);
or U2588 (N_2588,N_2046,N_2188);
or U2589 (N_2589,N_2297,N_2455);
nor U2590 (N_2590,N_2078,N_2358);
nand U2591 (N_2591,N_2426,N_2403);
nor U2592 (N_2592,N_2469,N_2155);
or U2593 (N_2593,N_2311,N_2261);
nor U2594 (N_2594,N_2386,N_2032);
or U2595 (N_2595,N_2151,N_2404);
and U2596 (N_2596,N_2232,N_2193);
and U2597 (N_2597,N_2289,N_2307);
nand U2598 (N_2598,N_2147,N_2313);
and U2599 (N_2599,N_2478,N_2018);
or U2600 (N_2600,N_2037,N_2178);
or U2601 (N_2601,N_2075,N_2316);
nand U2602 (N_2602,N_2306,N_2070);
xnor U2603 (N_2603,N_2286,N_2066);
nor U2604 (N_2604,N_2189,N_2187);
and U2605 (N_2605,N_2421,N_2159);
xnor U2606 (N_2606,N_2139,N_2054);
nor U2607 (N_2607,N_2387,N_2476);
nand U2608 (N_2608,N_2233,N_2298);
nand U2609 (N_2609,N_2055,N_2413);
and U2610 (N_2610,N_2215,N_2182);
and U2611 (N_2611,N_2076,N_2367);
and U2612 (N_2612,N_2132,N_2398);
nor U2613 (N_2613,N_2273,N_2236);
nor U2614 (N_2614,N_2257,N_2203);
xor U2615 (N_2615,N_2376,N_2085);
or U2616 (N_2616,N_2009,N_2323);
and U2617 (N_2617,N_2235,N_2190);
nor U2618 (N_2618,N_2237,N_2389);
nand U2619 (N_2619,N_2475,N_2479);
or U2620 (N_2620,N_2049,N_2117);
nor U2621 (N_2621,N_2322,N_2062);
nor U2622 (N_2622,N_2119,N_2131);
or U2623 (N_2623,N_2296,N_2245);
nand U2624 (N_2624,N_2381,N_2064);
or U2625 (N_2625,N_2314,N_2168);
nand U2626 (N_2626,N_2366,N_2434);
xor U2627 (N_2627,N_2129,N_2344);
nand U2628 (N_2628,N_2022,N_2391);
nand U2629 (N_2629,N_2342,N_2118);
nor U2630 (N_2630,N_2407,N_2028);
and U2631 (N_2631,N_2014,N_2449);
or U2632 (N_2632,N_2300,N_2167);
or U2633 (N_2633,N_2205,N_2016);
nand U2634 (N_2634,N_2465,N_2484);
nand U2635 (N_2635,N_2463,N_2074);
nor U2636 (N_2636,N_2338,N_2047);
or U2637 (N_2637,N_2053,N_2059);
nor U2638 (N_2638,N_2216,N_2473);
and U2639 (N_2639,N_2246,N_2057);
nor U2640 (N_2640,N_2169,N_2201);
or U2641 (N_2641,N_2303,N_2309);
xnor U2642 (N_2642,N_2445,N_2397);
and U2643 (N_2643,N_2105,N_2211);
nor U2644 (N_2644,N_2345,N_2341);
and U2645 (N_2645,N_2271,N_2081);
xnor U2646 (N_2646,N_2142,N_2467);
nand U2647 (N_2647,N_2154,N_2173);
xor U2648 (N_2648,N_2013,N_2184);
nand U2649 (N_2649,N_2007,N_2304);
or U2650 (N_2650,N_2012,N_2071);
nand U2651 (N_2651,N_2320,N_2402);
and U2652 (N_2652,N_2200,N_2410);
and U2653 (N_2653,N_2165,N_2227);
nor U2654 (N_2654,N_2357,N_2025);
nor U2655 (N_2655,N_2464,N_2004);
and U2656 (N_2656,N_2401,N_2466);
nand U2657 (N_2657,N_2396,N_2459);
and U2658 (N_2658,N_2163,N_2470);
xnor U2659 (N_2659,N_2231,N_2153);
nor U2660 (N_2660,N_2496,N_2498);
or U2661 (N_2661,N_2400,N_2336);
nand U2662 (N_2662,N_2069,N_2371);
and U2663 (N_2663,N_2002,N_2346);
nor U2664 (N_2664,N_2499,N_2406);
and U2665 (N_2665,N_2043,N_2217);
nand U2666 (N_2666,N_2052,N_2033);
nand U2667 (N_2667,N_2293,N_2441);
nand U2668 (N_2668,N_2006,N_2369);
nor U2669 (N_2669,N_2444,N_2383);
nand U2670 (N_2670,N_2332,N_2209);
nand U2671 (N_2671,N_2084,N_2360);
and U2672 (N_2672,N_2044,N_2351);
or U2673 (N_2673,N_2230,N_2162);
nor U2674 (N_2674,N_2026,N_2372);
or U2675 (N_2675,N_2127,N_2422);
nor U2676 (N_2676,N_2138,N_2146);
or U2677 (N_2677,N_2242,N_2299);
nor U2678 (N_2678,N_2176,N_2094);
nand U2679 (N_2679,N_2030,N_2240);
and U2680 (N_2680,N_2321,N_2353);
and U2681 (N_2681,N_2267,N_2198);
nor U2682 (N_2682,N_2087,N_2140);
xnor U2683 (N_2683,N_2164,N_2327);
or U2684 (N_2684,N_2040,N_2143);
and U2685 (N_2685,N_2107,N_2253);
and U2686 (N_2686,N_2170,N_2008);
or U2687 (N_2687,N_2207,N_2238);
or U2688 (N_2688,N_2315,N_2482);
and U2689 (N_2689,N_2091,N_2456);
nand U2690 (N_2690,N_2001,N_2204);
nand U2691 (N_2691,N_2337,N_2073);
nand U2692 (N_2692,N_2412,N_2247);
nor U2693 (N_2693,N_2058,N_2020);
and U2694 (N_2694,N_2206,N_2312);
nor U2695 (N_2695,N_2137,N_2171);
or U2696 (N_2696,N_2430,N_2439);
nand U2697 (N_2697,N_2454,N_2248);
nor U2698 (N_2698,N_2339,N_2166);
xor U2699 (N_2699,N_2363,N_2197);
nor U2700 (N_2700,N_2254,N_2029);
or U2701 (N_2701,N_2265,N_2318);
and U2702 (N_2702,N_2249,N_2250);
nor U2703 (N_2703,N_2493,N_2432);
xor U2704 (N_2704,N_2060,N_2438);
nor U2705 (N_2705,N_2490,N_2379);
and U2706 (N_2706,N_2225,N_2281);
nand U2707 (N_2707,N_2149,N_2335);
or U2708 (N_2708,N_2090,N_2079);
nor U2709 (N_2709,N_2488,N_2175);
or U2710 (N_2710,N_2260,N_2462);
or U2711 (N_2711,N_2061,N_2148);
nand U2712 (N_2712,N_2208,N_2348);
or U2713 (N_2713,N_2481,N_2270);
and U2714 (N_2714,N_2278,N_2460);
or U2715 (N_2715,N_2362,N_2288);
or U2716 (N_2716,N_2437,N_2183);
xnor U2717 (N_2717,N_2295,N_2393);
nor U2718 (N_2718,N_2027,N_2263);
or U2719 (N_2719,N_2097,N_2042);
and U2720 (N_2720,N_2319,N_2269);
and U2721 (N_2721,N_2450,N_2264);
nand U2722 (N_2722,N_2262,N_2221);
or U2723 (N_2723,N_2480,N_2390);
nand U2724 (N_2724,N_2272,N_2429);
and U2725 (N_2725,N_2220,N_2036);
nand U2726 (N_2726,N_2222,N_2417);
nand U2727 (N_2727,N_2095,N_2219);
nand U2728 (N_2728,N_2158,N_2328);
xnor U2729 (N_2729,N_2122,N_2333);
or U2730 (N_2730,N_2186,N_2424);
and U2731 (N_2731,N_2093,N_2349);
nor U2732 (N_2732,N_2384,N_2368);
nand U2733 (N_2733,N_2124,N_2485);
nor U2734 (N_2734,N_2414,N_2113);
xnor U2735 (N_2735,N_2072,N_2359);
and U2736 (N_2736,N_2326,N_2292);
nand U2737 (N_2737,N_2089,N_2409);
nor U2738 (N_2738,N_2282,N_2038);
or U2739 (N_2739,N_2099,N_2392);
nor U2740 (N_2740,N_2031,N_2202);
nand U2741 (N_2741,N_2180,N_2181);
and U2742 (N_2742,N_2251,N_2080);
or U2743 (N_2743,N_2283,N_2474);
nor U2744 (N_2744,N_2228,N_2308);
nand U2745 (N_2745,N_2106,N_2041);
nor U2746 (N_2746,N_2111,N_2477);
nand U2747 (N_2747,N_2431,N_2224);
nor U2748 (N_2748,N_2305,N_2050);
or U2749 (N_2749,N_2125,N_2276);
nand U2750 (N_2750,N_2149,N_2120);
nor U2751 (N_2751,N_2300,N_2115);
and U2752 (N_2752,N_2481,N_2022);
and U2753 (N_2753,N_2178,N_2390);
nand U2754 (N_2754,N_2217,N_2316);
nor U2755 (N_2755,N_2297,N_2300);
nand U2756 (N_2756,N_2020,N_2189);
and U2757 (N_2757,N_2394,N_2475);
and U2758 (N_2758,N_2290,N_2372);
nand U2759 (N_2759,N_2337,N_2163);
nor U2760 (N_2760,N_2013,N_2200);
and U2761 (N_2761,N_2048,N_2351);
or U2762 (N_2762,N_2073,N_2260);
nand U2763 (N_2763,N_2368,N_2194);
or U2764 (N_2764,N_2372,N_2089);
or U2765 (N_2765,N_2044,N_2375);
nand U2766 (N_2766,N_2436,N_2103);
or U2767 (N_2767,N_2338,N_2042);
xor U2768 (N_2768,N_2361,N_2421);
nor U2769 (N_2769,N_2163,N_2336);
xnor U2770 (N_2770,N_2415,N_2124);
or U2771 (N_2771,N_2084,N_2337);
and U2772 (N_2772,N_2327,N_2295);
nor U2773 (N_2773,N_2045,N_2498);
or U2774 (N_2774,N_2406,N_2431);
and U2775 (N_2775,N_2373,N_2305);
nand U2776 (N_2776,N_2270,N_2053);
nor U2777 (N_2777,N_2012,N_2037);
or U2778 (N_2778,N_2309,N_2041);
xor U2779 (N_2779,N_2128,N_2198);
nor U2780 (N_2780,N_2235,N_2088);
and U2781 (N_2781,N_2008,N_2029);
nand U2782 (N_2782,N_2457,N_2438);
nor U2783 (N_2783,N_2361,N_2467);
nor U2784 (N_2784,N_2384,N_2445);
nand U2785 (N_2785,N_2248,N_2472);
and U2786 (N_2786,N_2390,N_2418);
nand U2787 (N_2787,N_2102,N_2397);
or U2788 (N_2788,N_2277,N_2026);
nor U2789 (N_2789,N_2163,N_2298);
and U2790 (N_2790,N_2120,N_2083);
and U2791 (N_2791,N_2314,N_2081);
or U2792 (N_2792,N_2370,N_2168);
nor U2793 (N_2793,N_2095,N_2266);
or U2794 (N_2794,N_2020,N_2386);
xnor U2795 (N_2795,N_2148,N_2081);
nand U2796 (N_2796,N_2329,N_2108);
nor U2797 (N_2797,N_2351,N_2132);
nand U2798 (N_2798,N_2167,N_2260);
or U2799 (N_2799,N_2074,N_2145);
nand U2800 (N_2800,N_2114,N_2415);
nor U2801 (N_2801,N_2468,N_2499);
or U2802 (N_2802,N_2451,N_2453);
nand U2803 (N_2803,N_2361,N_2338);
nand U2804 (N_2804,N_2007,N_2277);
nand U2805 (N_2805,N_2254,N_2047);
nand U2806 (N_2806,N_2155,N_2370);
and U2807 (N_2807,N_2236,N_2261);
and U2808 (N_2808,N_2027,N_2436);
or U2809 (N_2809,N_2198,N_2357);
nand U2810 (N_2810,N_2010,N_2052);
nand U2811 (N_2811,N_2478,N_2131);
or U2812 (N_2812,N_2433,N_2494);
or U2813 (N_2813,N_2482,N_2032);
or U2814 (N_2814,N_2141,N_2123);
nor U2815 (N_2815,N_2429,N_2028);
or U2816 (N_2816,N_2464,N_2007);
nor U2817 (N_2817,N_2327,N_2364);
and U2818 (N_2818,N_2008,N_2482);
nand U2819 (N_2819,N_2263,N_2433);
nand U2820 (N_2820,N_2182,N_2454);
or U2821 (N_2821,N_2430,N_2246);
nor U2822 (N_2822,N_2181,N_2259);
and U2823 (N_2823,N_2457,N_2166);
nand U2824 (N_2824,N_2082,N_2072);
nor U2825 (N_2825,N_2120,N_2254);
and U2826 (N_2826,N_2491,N_2431);
or U2827 (N_2827,N_2480,N_2448);
and U2828 (N_2828,N_2300,N_2311);
or U2829 (N_2829,N_2274,N_2327);
or U2830 (N_2830,N_2043,N_2279);
nor U2831 (N_2831,N_2337,N_2233);
or U2832 (N_2832,N_2461,N_2273);
and U2833 (N_2833,N_2172,N_2214);
nor U2834 (N_2834,N_2172,N_2007);
xor U2835 (N_2835,N_2067,N_2321);
xnor U2836 (N_2836,N_2224,N_2345);
or U2837 (N_2837,N_2383,N_2341);
and U2838 (N_2838,N_2249,N_2153);
xor U2839 (N_2839,N_2333,N_2383);
nor U2840 (N_2840,N_2135,N_2058);
or U2841 (N_2841,N_2180,N_2264);
nand U2842 (N_2842,N_2339,N_2075);
xor U2843 (N_2843,N_2198,N_2373);
nand U2844 (N_2844,N_2081,N_2201);
nand U2845 (N_2845,N_2004,N_2161);
and U2846 (N_2846,N_2368,N_2161);
xnor U2847 (N_2847,N_2390,N_2109);
and U2848 (N_2848,N_2062,N_2264);
nor U2849 (N_2849,N_2271,N_2197);
xnor U2850 (N_2850,N_2364,N_2132);
and U2851 (N_2851,N_2414,N_2489);
nand U2852 (N_2852,N_2089,N_2121);
nand U2853 (N_2853,N_2470,N_2465);
or U2854 (N_2854,N_2158,N_2007);
and U2855 (N_2855,N_2273,N_2339);
nor U2856 (N_2856,N_2320,N_2468);
nor U2857 (N_2857,N_2284,N_2127);
or U2858 (N_2858,N_2426,N_2066);
or U2859 (N_2859,N_2083,N_2101);
and U2860 (N_2860,N_2361,N_2292);
nand U2861 (N_2861,N_2213,N_2151);
nand U2862 (N_2862,N_2233,N_2469);
or U2863 (N_2863,N_2084,N_2247);
or U2864 (N_2864,N_2229,N_2016);
and U2865 (N_2865,N_2038,N_2377);
nand U2866 (N_2866,N_2446,N_2121);
nor U2867 (N_2867,N_2316,N_2266);
and U2868 (N_2868,N_2204,N_2498);
nor U2869 (N_2869,N_2102,N_2414);
and U2870 (N_2870,N_2100,N_2253);
and U2871 (N_2871,N_2090,N_2238);
nor U2872 (N_2872,N_2410,N_2485);
and U2873 (N_2873,N_2280,N_2383);
nor U2874 (N_2874,N_2228,N_2365);
and U2875 (N_2875,N_2197,N_2405);
and U2876 (N_2876,N_2087,N_2146);
xor U2877 (N_2877,N_2269,N_2122);
or U2878 (N_2878,N_2055,N_2329);
nor U2879 (N_2879,N_2176,N_2121);
or U2880 (N_2880,N_2303,N_2221);
and U2881 (N_2881,N_2156,N_2333);
and U2882 (N_2882,N_2106,N_2029);
and U2883 (N_2883,N_2120,N_2398);
or U2884 (N_2884,N_2110,N_2234);
nand U2885 (N_2885,N_2111,N_2473);
nor U2886 (N_2886,N_2387,N_2058);
or U2887 (N_2887,N_2495,N_2337);
or U2888 (N_2888,N_2179,N_2303);
xnor U2889 (N_2889,N_2277,N_2330);
and U2890 (N_2890,N_2353,N_2239);
and U2891 (N_2891,N_2249,N_2323);
nand U2892 (N_2892,N_2456,N_2244);
or U2893 (N_2893,N_2283,N_2333);
and U2894 (N_2894,N_2351,N_2075);
nor U2895 (N_2895,N_2427,N_2205);
and U2896 (N_2896,N_2425,N_2464);
or U2897 (N_2897,N_2133,N_2191);
and U2898 (N_2898,N_2090,N_2169);
nand U2899 (N_2899,N_2054,N_2040);
xor U2900 (N_2900,N_2292,N_2310);
nand U2901 (N_2901,N_2353,N_2147);
nand U2902 (N_2902,N_2471,N_2488);
nand U2903 (N_2903,N_2396,N_2493);
nor U2904 (N_2904,N_2212,N_2403);
nor U2905 (N_2905,N_2153,N_2460);
nor U2906 (N_2906,N_2117,N_2169);
or U2907 (N_2907,N_2350,N_2471);
nand U2908 (N_2908,N_2237,N_2098);
nor U2909 (N_2909,N_2307,N_2211);
or U2910 (N_2910,N_2130,N_2045);
and U2911 (N_2911,N_2358,N_2301);
xnor U2912 (N_2912,N_2098,N_2465);
nand U2913 (N_2913,N_2357,N_2499);
nor U2914 (N_2914,N_2067,N_2173);
and U2915 (N_2915,N_2240,N_2194);
or U2916 (N_2916,N_2008,N_2318);
xnor U2917 (N_2917,N_2335,N_2124);
nand U2918 (N_2918,N_2169,N_2373);
xnor U2919 (N_2919,N_2480,N_2309);
nand U2920 (N_2920,N_2241,N_2075);
nor U2921 (N_2921,N_2364,N_2120);
nor U2922 (N_2922,N_2499,N_2055);
xnor U2923 (N_2923,N_2188,N_2404);
and U2924 (N_2924,N_2064,N_2315);
xor U2925 (N_2925,N_2075,N_2301);
and U2926 (N_2926,N_2260,N_2134);
nor U2927 (N_2927,N_2097,N_2402);
xor U2928 (N_2928,N_2139,N_2074);
nand U2929 (N_2929,N_2128,N_2442);
nor U2930 (N_2930,N_2318,N_2386);
and U2931 (N_2931,N_2131,N_2073);
and U2932 (N_2932,N_2475,N_2355);
and U2933 (N_2933,N_2222,N_2325);
or U2934 (N_2934,N_2325,N_2188);
nor U2935 (N_2935,N_2393,N_2092);
nor U2936 (N_2936,N_2301,N_2068);
or U2937 (N_2937,N_2184,N_2179);
xnor U2938 (N_2938,N_2161,N_2163);
or U2939 (N_2939,N_2121,N_2322);
nor U2940 (N_2940,N_2399,N_2370);
nand U2941 (N_2941,N_2150,N_2058);
nand U2942 (N_2942,N_2428,N_2174);
or U2943 (N_2943,N_2062,N_2066);
or U2944 (N_2944,N_2259,N_2252);
and U2945 (N_2945,N_2259,N_2286);
nand U2946 (N_2946,N_2130,N_2310);
nand U2947 (N_2947,N_2215,N_2281);
xor U2948 (N_2948,N_2113,N_2402);
and U2949 (N_2949,N_2211,N_2230);
and U2950 (N_2950,N_2033,N_2190);
xnor U2951 (N_2951,N_2317,N_2393);
or U2952 (N_2952,N_2178,N_2320);
and U2953 (N_2953,N_2120,N_2404);
nor U2954 (N_2954,N_2065,N_2079);
nand U2955 (N_2955,N_2487,N_2485);
nand U2956 (N_2956,N_2185,N_2261);
nor U2957 (N_2957,N_2446,N_2461);
nor U2958 (N_2958,N_2334,N_2292);
nand U2959 (N_2959,N_2337,N_2405);
and U2960 (N_2960,N_2019,N_2182);
and U2961 (N_2961,N_2009,N_2180);
nor U2962 (N_2962,N_2050,N_2169);
nand U2963 (N_2963,N_2467,N_2117);
nor U2964 (N_2964,N_2051,N_2120);
and U2965 (N_2965,N_2082,N_2438);
and U2966 (N_2966,N_2313,N_2004);
and U2967 (N_2967,N_2253,N_2435);
nor U2968 (N_2968,N_2090,N_2324);
or U2969 (N_2969,N_2191,N_2152);
and U2970 (N_2970,N_2410,N_2486);
or U2971 (N_2971,N_2127,N_2286);
nand U2972 (N_2972,N_2107,N_2446);
nor U2973 (N_2973,N_2415,N_2284);
nand U2974 (N_2974,N_2251,N_2001);
nor U2975 (N_2975,N_2141,N_2007);
xnor U2976 (N_2976,N_2000,N_2281);
and U2977 (N_2977,N_2449,N_2119);
nand U2978 (N_2978,N_2304,N_2310);
nand U2979 (N_2979,N_2154,N_2155);
and U2980 (N_2980,N_2044,N_2397);
or U2981 (N_2981,N_2216,N_2187);
or U2982 (N_2982,N_2201,N_2437);
or U2983 (N_2983,N_2193,N_2077);
or U2984 (N_2984,N_2496,N_2254);
xor U2985 (N_2985,N_2387,N_2200);
or U2986 (N_2986,N_2345,N_2469);
or U2987 (N_2987,N_2207,N_2029);
or U2988 (N_2988,N_2370,N_2079);
nor U2989 (N_2989,N_2245,N_2495);
and U2990 (N_2990,N_2375,N_2198);
and U2991 (N_2991,N_2389,N_2087);
and U2992 (N_2992,N_2291,N_2342);
nor U2993 (N_2993,N_2048,N_2022);
nor U2994 (N_2994,N_2130,N_2182);
nand U2995 (N_2995,N_2280,N_2115);
or U2996 (N_2996,N_2479,N_2384);
xnor U2997 (N_2997,N_2407,N_2312);
xor U2998 (N_2998,N_2476,N_2027);
xor U2999 (N_2999,N_2334,N_2294);
or U3000 (N_3000,N_2862,N_2677);
nand U3001 (N_3001,N_2659,N_2924);
and U3002 (N_3002,N_2533,N_2841);
or U3003 (N_3003,N_2702,N_2519);
nand U3004 (N_3004,N_2856,N_2693);
nand U3005 (N_3005,N_2612,N_2925);
or U3006 (N_3006,N_2548,N_2880);
nor U3007 (N_3007,N_2776,N_2854);
nand U3008 (N_3008,N_2571,N_2797);
nor U3009 (N_3009,N_2564,N_2950);
nor U3010 (N_3010,N_2573,N_2584);
nor U3011 (N_3011,N_2994,N_2651);
and U3012 (N_3012,N_2608,N_2722);
or U3013 (N_3013,N_2923,N_2602);
nand U3014 (N_3014,N_2687,N_2648);
nand U3015 (N_3015,N_2511,N_2665);
and U3016 (N_3016,N_2973,N_2565);
and U3017 (N_3017,N_2739,N_2501);
nand U3018 (N_3018,N_2846,N_2765);
nand U3019 (N_3019,N_2538,N_2513);
and U3020 (N_3020,N_2509,N_2615);
or U3021 (N_3021,N_2874,N_2696);
nor U3022 (N_3022,N_2892,N_2670);
or U3023 (N_3023,N_2601,N_2760);
nor U3024 (N_3024,N_2627,N_2568);
and U3025 (N_3025,N_2577,N_2660);
xor U3026 (N_3026,N_2596,N_2764);
or U3027 (N_3027,N_2713,N_2691);
and U3028 (N_3028,N_2586,N_2837);
nor U3029 (N_3029,N_2530,N_2561);
nand U3030 (N_3030,N_2931,N_2575);
or U3031 (N_3031,N_2667,N_2685);
nor U3032 (N_3032,N_2801,N_2882);
or U3033 (N_3033,N_2743,N_2692);
and U3034 (N_3034,N_2542,N_2910);
or U3035 (N_3035,N_2682,N_2606);
nor U3036 (N_3036,N_2843,N_2671);
or U3037 (N_3037,N_2562,N_2644);
nor U3038 (N_3038,N_2832,N_2870);
and U3039 (N_3039,N_2942,N_2840);
nand U3040 (N_3040,N_2864,N_2547);
and U3041 (N_3041,N_2886,N_2588);
or U3042 (N_3042,N_2626,N_2933);
or U3043 (N_3043,N_2930,N_2728);
nand U3044 (N_3044,N_2723,N_2536);
and U3045 (N_3045,N_2850,N_2636);
or U3046 (N_3046,N_2907,N_2909);
nor U3047 (N_3047,N_2635,N_2617);
nor U3048 (N_3048,N_2629,N_2865);
nor U3049 (N_3049,N_2638,N_2855);
or U3050 (N_3050,N_2806,N_2947);
nand U3051 (N_3051,N_2952,N_2811);
nand U3052 (N_3052,N_2554,N_2639);
nand U3053 (N_3053,N_2594,N_2783);
and U3054 (N_3054,N_2553,N_2919);
and U3055 (N_3055,N_2642,N_2992);
or U3056 (N_3056,N_2695,N_2624);
and U3057 (N_3057,N_2675,N_2968);
nor U3058 (N_3058,N_2712,N_2830);
nand U3059 (N_3059,N_2911,N_2676);
and U3060 (N_3060,N_2936,N_2966);
xnor U3061 (N_3061,N_2767,N_2844);
or U3062 (N_3062,N_2944,N_2726);
nor U3063 (N_3063,N_2503,N_2578);
and U3064 (N_3064,N_2887,N_2831);
or U3065 (N_3065,N_2938,N_2515);
xnor U3066 (N_3066,N_2972,N_2535);
nor U3067 (N_3067,N_2522,N_2592);
nor U3068 (N_3068,N_2890,N_2585);
nor U3069 (N_3069,N_2860,N_2607);
or U3070 (N_3070,N_2512,N_2816);
xor U3071 (N_3071,N_2956,N_2786);
and U3072 (N_3072,N_2662,N_2859);
or U3073 (N_3073,N_2755,N_2842);
or U3074 (N_3074,N_2981,N_2746);
nor U3075 (N_3075,N_2745,N_2502);
or U3076 (N_3076,N_2807,N_2523);
nand U3077 (N_3077,N_2645,N_2725);
nor U3078 (N_3078,N_2967,N_2818);
nand U3079 (N_3079,N_2897,N_2759);
nor U3080 (N_3080,N_2766,N_2861);
and U3081 (N_3081,N_2836,N_2544);
or U3082 (N_3082,N_2657,N_2922);
nor U3083 (N_3083,N_2556,N_2681);
nor U3084 (N_3084,N_2731,N_2793);
and U3085 (N_3085,N_2876,N_2906);
nand U3086 (N_3086,N_2835,N_2918);
nand U3087 (N_3087,N_2893,N_2738);
xor U3088 (N_3088,N_2852,N_2970);
nor U3089 (N_3089,N_2805,N_2747);
xnor U3090 (N_3090,N_2965,N_2959);
nor U3091 (N_3091,N_2749,N_2913);
and U3092 (N_3092,N_2782,N_2754);
or U3093 (N_3093,N_2714,N_2845);
xor U3094 (N_3094,N_2704,N_2974);
nor U3095 (N_3095,N_2800,N_2684);
or U3096 (N_3096,N_2761,N_2748);
and U3097 (N_3097,N_2688,N_2888);
and U3098 (N_3098,N_2595,N_2998);
and U3099 (N_3099,N_2729,N_2809);
nor U3100 (N_3100,N_2543,N_2875);
nand U3101 (N_3101,N_2560,N_2650);
nand U3102 (N_3102,N_2799,N_2686);
and U3103 (N_3103,N_2590,N_2534);
nand U3104 (N_3104,N_2983,N_2914);
nor U3105 (N_3105,N_2709,N_2891);
and U3106 (N_3106,N_2796,N_2763);
nor U3107 (N_3107,N_2567,N_2661);
nor U3108 (N_3108,N_2904,N_2620);
nor U3109 (N_3109,N_2896,N_2504);
and U3110 (N_3110,N_2653,N_2654);
or U3111 (N_3111,N_2742,N_2507);
nor U3112 (N_3112,N_2508,N_2581);
xnor U3113 (N_3113,N_2991,N_2770);
xnor U3114 (N_3114,N_2785,N_2987);
xnor U3115 (N_3115,N_2795,N_2630);
nor U3116 (N_3116,N_2881,N_2540);
and U3117 (N_3117,N_2812,N_2658);
nand U3118 (N_3118,N_2762,N_2963);
nand U3119 (N_3119,N_2618,N_2736);
nand U3120 (N_3120,N_2622,N_2599);
nand U3121 (N_3121,N_2949,N_2741);
or U3122 (N_3122,N_2539,N_2699);
nor U3123 (N_3123,N_2955,N_2905);
nand U3124 (N_3124,N_2710,N_2999);
nor U3125 (N_3125,N_2640,N_2941);
nand U3126 (N_3126,N_2621,N_2825);
nand U3127 (N_3127,N_2819,N_2777);
nand U3128 (N_3128,N_2690,N_2719);
xor U3129 (N_3129,N_2802,N_2945);
or U3130 (N_3130,N_2853,N_2996);
xor U3131 (N_3131,N_2733,N_2813);
and U3132 (N_3132,N_2928,N_2737);
nand U3133 (N_3133,N_2788,N_2935);
and U3134 (N_3134,N_2866,N_2932);
xor U3135 (N_3135,N_2637,N_2781);
nor U3136 (N_3136,N_2868,N_2823);
xnor U3137 (N_3137,N_2758,N_2895);
or U3138 (N_3138,N_2940,N_2735);
and U3139 (N_3139,N_2500,N_2810);
nand U3140 (N_3140,N_2834,N_2851);
or U3141 (N_3141,N_2623,N_2871);
nand U3142 (N_3142,N_2744,N_2953);
nor U3143 (N_3143,N_2598,N_2948);
nand U3144 (N_3144,N_2525,N_2526);
or U3145 (N_3145,N_2903,N_2814);
nand U3146 (N_3146,N_2899,N_2926);
xor U3147 (N_3147,N_2984,N_2529);
and U3148 (N_3148,N_2555,N_2971);
xor U3149 (N_3149,N_2908,N_2934);
nand U3150 (N_3150,N_2943,N_2756);
and U3151 (N_3151,N_2647,N_2833);
and U3152 (N_3152,N_2773,N_2715);
and U3153 (N_3153,N_2669,N_2921);
and U3154 (N_3154,N_2927,N_2700);
or U3155 (N_3155,N_2790,N_2939);
nor U3156 (N_3156,N_2962,N_2779);
or U3157 (N_3157,N_2817,N_2957);
nand U3158 (N_3158,N_2873,N_2656);
or U3159 (N_3159,N_2663,N_2720);
or U3160 (N_3160,N_2976,N_2993);
or U3161 (N_3161,N_2558,N_2610);
or U3162 (N_3162,N_2701,N_2531);
or U3163 (N_3163,N_2877,N_2582);
nand U3164 (N_3164,N_2570,N_2532);
nor U3165 (N_3165,N_2827,N_2698);
or U3166 (N_3166,N_2668,N_2694);
nand U3167 (N_3167,N_2858,N_2917);
and U3168 (N_3168,N_2550,N_2774);
nand U3169 (N_3169,N_2697,N_2849);
and U3170 (N_3170,N_2863,N_2969);
nand U3171 (N_3171,N_2775,N_2505);
and U3172 (N_3172,N_2803,N_2997);
and U3173 (N_3173,N_2516,N_2520);
nor U3174 (N_3174,N_2619,N_2546);
and U3175 (N_3175,N_2826,N_2666);
nor U3176 (N_3176,N_2980,N_2557);
and U3177 (N_3177,N_2611,N_2528);
or U3178 (N_3178,N_2768,N_2683);
or U3179 (N_3179,N_2625,N_2900);
nand U3180 (N_3180,N_2808,N_2978);
nand U3181 (N_3181,N_2792,N_2829);
nor U3182 (N_3182,N_2679,N_2721);
or U3183 (N_3183,N_2705,N_2798);
nand U3184 (N_3184,N_2857,N_2847);
and U3185 (N_3185,N_2883,N_2632);
and U3186 (N_3186,N_2583,N_2951);
nand U3187 (N_3187,N_2521,N_2616);
xor U3188 (N_3188,N_2960,N_2757);
or U3189 (N_3189,N_2838,N_2605);
nand U3190 (N_3190,N_2631,N_2549);
nand U3191 (N_3191,N_2609,N_2824);
or U3192 (N_3192,N_2958,N_2664);
nand U3193 (N_3193,N_2655,N_2506);
nor U3194 (N_3194,N_2920,N_2989);
nand U3195 (N_3195,N_2672,N_2641);
and U3196 (N_3196,N_2514,N_2791);
and U3197 (N_3197,N_2678,N_2517);
and U3198 (N_3198,N_2649,N_2706);
xnor U3199 (N_3199,N_2794,N_2551);
and U3200 (N_3200,N_2784,N_2646);
nand U3201 (N_3201,N_2885,N_2977);
or U3202 (N_3202,N_2869,N_2717);
and U3203 (N_3203,N_2916,N_2878);
nor U3204 (N_3204,N_2559,N_2990);
xnor U3205 (N_3205,N_2674,N_2822);
nand U3206 (N_3206,N_2778,N_2894);
or U3207 (N_3207,N_2541,N_2789);
and U3208 (N_3208,N_2703,N_2982);
or U3209 (N_3209,N_2988,N_2740);
and U3210 (N_3210,N_2954,N_2937);
nand U3211 (N_3211,N_2634,N_2727);
or U3212 (N_3212,N_2566,N_2572);
nand U3213 (N_3213,N_2995,N_2839);
nand U3214 (N_3214,N_2527,N_2732);
xor U3215 (N_3215,N_2751,N_2884);
and U3216 (N_3216,N_2587,N_2753);
and U3217 (N_3217,N_2724,N_2769);
or U3218 (N_3218,N_2772,N_2591);
xor U3219 (N_3219,N_2603,N_2771);
nand U3220 (N_3220,N_2711,N_2633);
nand U3221 (N_3221,N_2689,N_2708);
and U3222 (N_3222,N_2867,N_2579);
and U3223 (N_3223,N_2750,N_2628);
nor U3224 (N_3224,N_2545,N_2821);
nand U3225 (N_3225,N_2912,N_2964);
nor U3226 (N_3226,N_2929,N_2879);
xnor U3227 (N_3227,N_2975,N_2597);
nor U3228 (N_3228,N_2820,N_2574);
nand U3229 (N_3229,N_2569,N_2510);
or U3230 (N_3230,N_2537,N_2518);
nor U3231 (N_3231,N_2716,N_2614);
xor U3232 (N_3232,N_2589,N_2828);
nor U3233 (N_3233,N_2848,N_2718);
nand U3234 (N_3234,N_2898,N_2986);
nor U3235 (N_3235,N_2804,N_2707);
nand U3236 (N_3236,N_2915,N_2889);
nand U3237 (N_3237,N_2580,N_2985);
xor U3238 (N_3238,N_2604,N_2652);
nor U3239 (N_3239,N_2872,N_2600);
and U3240 (N_3240,N_2552,N_2593);
nor U3241 (N_3241,N_2946,N_2780);
and U3242 (N_3242,N_2901,N_2730);
xor U3243 (N_3243,N_2613,N_2979);
nor U3244 (N_3244,N_2752,N_2524);
and U3245 (N_3245,N_2563,N_2680);
and U3246 (N_3246,N_2734,N_2643);
and U3247 (N_3247,N_2902,N_2961);
xor U3248 (N_3248,N_2673,N_2787);
nor U3249 (N_3249,N_2815,N_2576);
nor U3250 (N_3250,N_2525,N_2881);
nand U3251 (N_3251,N_2954,N_2570);
nor U3252 (N_3252,N_2844,N_2585);
xor U3253 (N_3253,N_2984,N_2999);
nor U3254 (N_3254,N_2977,N_2763);
or U3255 (N_3255,N_2795,N_2626);
and U3256 (N_3256,N_2737,N_2939);
and U3257 (N_3257,N_2909,N_2677);
or U3258 (N_3258,N_2582,N_2536);
xor U3259 (N_3259,N_2878,N_2950);
and U3260 (N_3260,N_2667,N_2966);
or U3261 (N_3261,N_2781,N_2922);
or U3262 (N_3262,N_2573,N_2750);
or U3263 (N_3263,N_2983,N_2676);
and U3264 (N_3264,N_2928,N_2741);
or U3265 (N_3265,N_2970,N_2550);
and U3266 (N_3266,N_2822,N_2996);
and U3267 (N_3267,N_2865,N_2930);
and U3268 (N_3268,N_2931,N_2935);
xnor U3269 (N_3269,N_2704,N_2637);
nand U3270 (N_3270,N_2684,N_2974);
nor U3271 (N_3271,N_2838,N_2677);
xnor U3272 (N_3272,N_2587,N_2575);
nand U3273 (N_3273,N_2875,N_2941);
nand U3274 (N_3274,N_2639,N_2573);
nand U3275 (N_3275,N_2890,N_2799);
nor U3276 (N_3276,N_2880,N_2766);
nor U3277 (N_3277,N_2891,N_2942);
nand U3278 (N_3278,N_2546,N_2584);
nor U3279 (N_3279,N_2948,N_2511);
nor U3280 (N_3280,N_2934,N_2619);
nor U3281 (N_3281,N_2883,N_2972);
nor U3282 (N_3282,N_2514,N_2869);
nand U3283 (N_3283,N_2701,N_2550);
nor U3284 (N_3284,N_2776,N_2527);
nand U3285 (N_3285,N_2786,N_2691);
or U3286 (N_3286,N_2970,N_2608);
nand U3287 (N_3287,N_2910,N_2630);
nor U3288 (N_3288,N_2906,N_2735);
or U3289 (N_3289,N_2778,N_2970);
or U3290 (N_3290,N_2960,N_2820);
nand U3291 (N_3291,N_2711,N_2527);
and U3292 (N_3292,N_2871,N_2653);
nor U3293 (N_3293,N_2515,N_2730);
xor U3294 (N_3294,N_2913,N_2501);
or U3295 (N_3295,N_2644,N_2859);
or U3296 (N_3296,N_2771,N_2649);
and U3297 (N_3297,N_2804,N_2715);
nand U3298 (N_3298,N_2939,N_2644);
nand U3299 (N_3299,N_2738,N_2949);
or U3300 (N_3300,N_2670,N_2791);
nand U3301 (N_3301,N_2656,N_2767);
and U3302 (N_3302,N_2836,N_2504);
or U3303 (N_3303,N_2523,N_2540);
and U3304 (N_3304,N_2506,N_2845);
and U3305 (N_3305,N_2698,N_2717);
xor U3306 (N_3306,N_2742,N_2957);
nand U3307 (N_3307,N_2925,N_2970);
xnor U3308 (N_3308,N_2648,N_2676);
nor U3309 (N_3309,N_2883,N_2818);
and U3310 (N_3310,N_2854,N_2725);
and U3311 (N_3311,N_2856,N_2612);
or U3312 (N_3312,N_2927,N_2666);
nand U3313 (N_3313,N_2950,N_2588);
or U3314 (N_3314,N_2510,N_2549);
xnor U3315 (N_3315,N_2707,N_2540);
nor U3316 (N_3316,N_2979,N_2761);
or U3317 (N_3317,N_2940,N_2726);
xnor U3318 (N_3318,N_2821,N_2595);
and U3319 (N_3319,N_2655,N_2788);
or U3320 (N_3320,N_2698,N_2570);
or U3321 (N_3321,N_2733,N_2633);
nor U3322 (N_3322,N_2936,N_2831);
and U3323 (N_3323,N_2725,N_2967);
or U3324 (N_3324,N_2606,N_2985);
nor U3325 (N_3325,N_2647,N_2913);
or U3326 (N_3326,N_2646,N_2724);
nor U3327 (N_3327,N_2840,N_2866);
nor U3328 (N_3328,N_2675,N_2503);
or U3329 (N_3329,N_2891,N_2889);
nor U3330 (N_3330,N_2971,N_2698);
or U3331 (N_3331,N_2925,N_2734);
nand U3332 (N_3332,N_2818,N_2657);
or U3333 (N_3333,N_2907,N_2544);
and U3334 (N_3334,N_2695,N_2974);
nand U3335 (N_3335,N_2772,N_2552);
nand U3336 (N_3336,N_2639,N_2581);
xor U3337 (N_3337,N_2734,N_2562);
nand U3338 (N_3338,N_2941,N_2868);
or U3339 (N_3339,N_2843,N_2995);
nor U3340 (N_3340,N_2506,N_2955);
nand U3341 (N_3341,N_2605,N_2929);
xor U3342 (N_3342,N_2908,N_2911);
nor U3343 (N_3343,N_2850,N_2776);
xnor U3344 (N_3344,N_2969,N_2701);
nor U3345 (N_3345,N_2978,N_2870);
nor U3346 (N_3346,N_2846,N_2633);
nor U3347 (N_3347,N_2512,N_2514);
nor U3348 (N_3348,N_2912,N_2997);
or U3349 (N_3349,N_2723,N_2566);
nor U3350 (N_3350,N_2673,N_2587);
or U3351 (N_3351,N_2857,N_2596);
nor U3352 (N_3352,N_2792,N_2586);
or U3353 (N_3353,N_2606,N_2622);
or U3354 (N_3354,N_2514,N_2873);
and U3355 (N_3355,N_2651,N_2794);
nor U3356 (N_3356,N_2655,N_2633);
nor U3357 (N_3357,N_2572,N_2756);
and U3358 (N_3358,N_2703,N_2644);
nor U3359 (N_3359,N_2949,N_2839);
nand U3360 (N_3360,N_2768,N_2934);
nor U3361 (N_3361,N_2671,N_2998);
nand U3362 (N_3362,N_2614,N_2889);
or U3363 (N_3363,N_2511,N_2795);
or U3364 (N_3364,N_2715,N_2614);
and U3365 (N_3365,N_2539,N_2811);
nand U3366 (N_3366,N_2508,N_2864);
nor U3367 (N_3367,N_2773,N_2824);
nor U3368 (N_3368,N_2543,N_2825);
nor U3369 (N_3369,N_2622,N_2618);
or U3370 (N_3370,N_2768,N_2962);
xor U3371 (N_3371,N_2501,N_2976);
or U3372 (N_3372,N_2533,N_2532);
and U3373 (N_3373,N_2844,N_2774);
or U3374 (N_3374,N_2659,N_2795);
and U3375 (N_3375,N_2723,N_2587);
nand U3376 (N_3376,N_2680,N_2708);
or U3377 (N_3377,N_2682,N_2723);
nor U3378 (N_3378,N_2856,N_2970);
or U3379 (N_3379,N_2745,N_2672);
nand U3380 (N_3380,N_2556,N_2761);
nor U3381 (N_3381,N_2966,N_2625);
or U3382 (N_3382,N_2761,N_2877);
and U3383 (N_3383,N_2692,N_2752);
and U3384 (N_3384,N_2971,N_2516);
nand U3385 (N_3385,N_2657,N_2659);
nand U3386 (N_3386,N_2989,N_2526);
nand U3387 (N_3387,N_2681,N_2823);
xnor U3388 (N_3388,N_2614,N_2750);
and U3389 (N_3389,N_2830,N_2656);
nand U3390 (N_3390,N_2801,N_2741);
xnor U3391 (N_3391,N_2814,N_2612);
and U3392 (N_3392,N_2785,N_2572);
or U3393 (N_3393,N_2783,N_2899);
nand U3394 (N_3394,N_2631,N_2899);
nand U3395 (N_3395,N_2809,N_2825);
nand U3396 (N_3396,N_2681,N_2734);
nand U3397 (N_3397,N_2620,N_2833);
or U3398 (N_3398,N_2508,N_2881);
and U3399 (N_3399,N_2596,N_2522);
or U3400 (N_3400,N_2568,N_2854);
nand U3401 (N_3401,N_2692,N_2939);
xnor U3402 (N_3402,N_2809,N_2877);
nor U3403 (N_3403,N_2616,N_2663);
nand U3404 (N_3404,N_2523,N_2890);
nand U3405 (N_3405,N_2877,N_2892);
or U3406 (N_3406,N_2961,N_2828);
or U3407 (N_3407,N_2846,N_2737);
nor U3408 (N_3408,N_2755,N_2663);
nor U3409 (N_3409,N_2898,N_2866);
and U3410 (N_3410,N_2519,N_2676);
and U3411 (N_3411,N_2628,N_2870);
nand U3412 (N_3412,N_2851,N_2813);
nor U3413 (N_3413,N_2938,N_2789);
nand U3414 (N_3414,N_2991,N_2735);
or U3415 (N_3415,N_2806,N_2780);
nand U3416 (N_3416,N_2653,N_2974);
or U3417 (N_3417,N_2782,N_2712);
nor U3418 (N_3418,N_2637,N_2712);
nor U3419 (N_3419,N_2588,N_2579);
and U3420 (N_3420,N_2877,N_2625);
nor U3421 (N_3421,N_2542,N_2673);
or U3422 (N_3422,N_2652,N_2849);
or U3423 (N_3423,N_2978,N_2952);
or U3424 (N_3424,N_2742,N_2823);
nor U3425 (N_3425,N_2886,N_2967);
or U3426 (N_3426,N_2632,N_2710);
nor U3427 (N_3427,N_2526,N_2630);
and U3428 (N_3428,N_2594,N_2725);
nor U3429 (N_3429,N_2689,N_2988);
or U3430 (N_3430,N_2806,N_2532);
or U3431 (N_3431,N_2536,N_2900);
and U3432 (N_3432,N_2795,N_2813);
and U3433 (N_3433,N_2636,N_2673);
nor U3434 (N_3434,N_2925,N_2514);
or U3435 (N_3435,N_2585,N_2704);
xnor U3436 (N_3436,N_2845,N_2716);
or U3437 (N_3437,N_2960,N_2604);
or U3438 (N_3438,N_2806,N_2738);
and U3439 (N_3439,N_2984,N_2693);
nor U3440 (N_3440,N_2880,N_2803);
and U3441 (N_3441,N_2717,N_2763);
or U3442 (N_3442,N_2751,N_2670);
or U3443 (N_3443,N_2860,N_2712);
or U3444 (N_3444,N_2580,N_2522);
nor U3445 (N_3445,N_2598,N_2936);
nor U3446 (N_3446,N_2862,N_2658);
and U3447 (N_3447,N_2661,N_2524);
and U3448 (N_3448,N_2601,N_2908);
or U3449 (N_3449,N_2988,N_2831);
xnor U3450 (N_3450,N_2767,N_2729);
and U3451 (N_3451,N_2640,N_2604);
nor U3452 (N_3452,N_2958,N_2858);
or U3453 (N_3453,N_2719,N_2796);
or U3454 (N_3454,N_2929,N_2762);
xor U3455 (N_3455,N_2639,N_2637);
or U3456 (N_3456,N_2579,N_2753);
nand U3457 (N_3457,N_2741,N_2909);
nand U3458 (N_3458,N_2719,N_2639);
or U3459 (N_3459,N_2547,N_2514);
nand U3460 (N_3460,N_2595,N_2721);
nand U3461 (N_3461,N_2725,N_2732);
or U3462 (N_3462,N_2866,N_2727);
or U3463 (N_3463,N_2977,N_2910);
nor U3464 (N_3464,N_2728,N_2505);
nor U3465 (N_3465,N_2906,N_2641);
nor U3466 (N_3466,N_2808,N_2633);
nand U3467 (N_3467,N_2982,N_2947);
and U3468 (N_3468,N_2554,N_2795);
xor U3469 (N_3469,N_2813,N_2846);
and U3470 (N_3470,N_2951,N_2697);
nor U3471 (N_3471,N_2558,N_2917);
or U3472 (N_3472,N_2546,N_2642);
nor U3473 (N_3473,N_2635,N_2859);
nand U3474 (N_3474,N_2730,N_2728);
and U3475 (N_3475,N_2828,N_2522);
nor U3476 (N_3476,N_2978,N_2986);
nor U3477 (N_3477,N_2647,N_2644);
and U3478 (N_3478,N_2608,N_2713);
and U3479 (N_3479,N_2697,N_2679);
or U3480 (N_3480,N_2727,N_2827);
nand U3481 (N_3481,N_2827,N_2749);
or U3482 (N_3482,N_2646,N_2721);
nor U3483 (N_3483,N_2885,N_2803);
or U3484 (N_3484,N_2995,N_2924);
and U3485 (N_3485,N_2889,N_2649);
or U3486 (N_3486,N_2535,N_2917);
or U3487 (N_3487,N_2601,N_2700);
and U3488 (N_3488,N_2807,N_2912);
nor U3489 (N_3489,N_2505,N_2508);
or U3490 (N_3490,N_2760,N_2553);
or U3491 (N_3491,N_2826,N_2847);
or U3492 (N_3492,N_2763,N_2975);
nor U3493 (N_3493,N_2857,N_2720);
nand U3494 (N_3494,N_2984,N_2857);
nor U3495 (N_3495,N_2785,N_2835);
or U3496 (N_3496,N_2868,N_2836);
nand U3497 (N_3497,N_2520,N_2670);
nand U3498 (N_3498,N_2924,N_2849);
nor U3499 (N_3499,N_2796,N_2809);
and U3500 (N_3500,N_3357,N_3093);
and U3501 (N_3501,N_3188,N_3365);
xnor U3502 (N_3502,N_3432,N_3355);
nor U3503 (N_3503,N_3098,N_3394);
and U3504 (N_3504,N_3439,N_3419);
nand U3505 (N_3505,N_3135,N_3158);
nor U3506 (N_3506,N_3195,N_3386);
or U3507 (N_3507,N_3463,N_3026);
xnor U3508 (N_3508,N_3452,N_3390);
or U3509 (N_3509,N_3495,N_3115);
and U3510 (N_3510,N_3297,N_3097);
or U3511 (N_3511,N_3054,N_3142);
and U3512 (N_3512,N_3404,N_3018);
and U3513 (N_3513,N_3215,N_3451);
nor U3514 (N_3514,N_3434,N_3028);
and U3515 (N_3515,N_3482,N_3176);
and U3516 (N_3516,N_3475,N_3414);
nand U3517 (N_3517,N_3042,N_3352);
nand U3518 (N_3518,N_3260,N_3116);
nand U3519 (N_3519,N_3445,N_3177);
nor U3520 (N_3520,N_3418,N_3429);
or U3521 (N_3521,N_3435,N_3038);
and U3522 (N_3522,N_3029,N_3347);
nor U3523 (N_3523,N_3460,N_3479);
and U3524 (N_3524,N_3001,N_3339);
or U3525 (N_3525,N_3413,N_3321);
and U3526 (N_3526,N_3275,N_3247);
and U3527 (N_3527,N_3335,N_3349);
and U3528 (N_3528,N_3372,N_3300);
or U3529 (N_3529,N_3229,N_3251);
nand U3530 (N_3530,N_3313,N_3428);
xnor U3531 (N_3531,N_3049,N_3249);
xor U3532 (N_3532,N_3104,N_3200);
nor U3533 (N_3533,N_3217,N_3287);
nand U3534 (N_3534,N_3170,N_3002);
and U3535 (N_3535,N_3148,N_3204);
nor U3536 (N_3536,N_3157,N_3112);
and U3537 (N_3537,N_3320,N_3137);
and U3538 (N_3538,N_3232,N_3131);
nor U3539 (N_3539,N_3324,N_3449);
xor U3540 (N_3540,N_3107,N_3015);
nor U3541 (N_3541,N_3318,N_3261);
nor U3542 (N_3542,N_3284,N_3470);
nand U3543 (N_3543,N_3253,N_3395);
nor U3544 (N_3544,N_3130,N_3020);
or U3545 (N_3545,N_3017,N_3491);
nand U3546 (N_3546,N_3367,N_3025);
nor U3547 (N_3547,N_3089,N_3455);
nor U3548 (N_3548,N_3466,N_3108);
and U3549 (N_3549,N_3279,N_3389);
and U3550 (N_3550,N_3123,N_3024);
nor U3551 (N_3551,N_3380,N_3457);
or U3552 (N_3552,N_3415,N_3443);
or U3553 (N_3553,N_3384,N_3333);
xnor U3554 (N_3554,N_3294,N_3139);
nand U3555 (N_3555,N_3114,N_3370);
nand U3556 (N_3556,N_3043,N_3173);
nand U3557 (N_3557,N_3012,N_3153);
or U3558 (N_3558,N_3231,N_3030);
xnor U3559 (N_3559,N_3224,N_3272);
or U3560 (N_3560,N_3239,N_3496);
nand U3561 (N_3561,N_3222,N_3174);
nand U3562 (N_3562,N_3143,N_3233);
or U3563 (N_3563,N_3181,N_3315);
or U3564 (N_3564,N_3314,N_3252);
xnor U3565 (N_3565,N_3085,N_3493);
and U3566 (N_3566,N_3250,N_3334);
or U3567 (N_3567,N_3296,N_3486);
or U3568 (N_3568,N_3122,N_3154);
or U3569 (N_3569,N_3442,N_3140);
nand U3570 (N_3570,N_3133,N_3169);
or U3571 (N_3571,N_3377,N_3151);
nand U3572 (N_3572,N_3437,N_3492);
xnor U3573 (N_3573,N_3156,N_3406);
nor U3574 (N_3574,N_3331,N_3218);
nand U3575 (N_3575,N_3034,N_3382);
nand U3576 (N_3576,N_3468,N_3109);
nand U3577 (N_3577,N_3110,N_3403);
xor U3578 (N_3578,N_3301,N_3149);
or U3579 (N_3579,N_3128,N_3059);
nand U3580 (N_3580,N_3362,N_3490);
nand U3581 (N_3581,N_3255,N_3117);
nand U3582 (N_3582,N_3219,N_3405);
or U3583 (N_3583,N_3411,N_3262);
nor U3584 (N_3584,N_3364,N_3424);
nor U3585 (N_3585,N_3193,N_3086);
nor U3586 (N_3586,N_3388,N_3202);
nor U3587 (N_3587,N_3146,N_3119);
or U3588 (N_3588,N_3423,N_3336);
nand U3589 (N_3589,N_3263,N_3161);
or U3590 (N_3590,N_3256,N_3243);
or U3591 (N_3591,N_3118,N_3011);
or U3592 (N_3592,N_3307,N_3329);
or U3593 (N_3593,N_3062,N_3044);
xor U3594 (N_3594,N_3317,N_3348);
and U3595 (N_3595,N_3425,N_3316);
nor U3596 (N_3596,N_3407,N_3494);
and U3597 (N_3597,N_3258,N_3196);
and U3598 (N_3598,N_3427,N_3354);
xor U3599 (N_3599,N_3292,N_3291);
and U3600 (N_3600,N_3088,N_3276);
or U3601 (N_3601,N_3068,N_3477);
nand U3602 (N_3602,N_3421,N_3409);
or U3603 (N_3603,N_3066,N_3402);
nand U3604 (N_3604,N_3003,N_3126);
nand U3605 (N_3605,N_3448,N_3120);
xnor U3606 (N_3606,N_3100,N_3350);
nor U3607 (N_3607,N_3216,N_3381);
or U3608 (N_3608,N_3270,N_3266);
nor U3609 (N_3609,N_3371,N_3323);
or U3610 (N_3610,N_3285,N_3374);
xor U3611 (N_3611,N_3376,N_3295);
nor U3612 (N_3612,N_3240,N_3487);
nor U3613 (N_3613,N_3473,N_3072);
and U3614 (N_3614,N_3484,N_3060);
xor U3615 (N_3615,N_3071,N_3091);
and U3616 (N_3616,N_3446,N_3178);
xor U3617 (N_3617,N_3076,N_3447);
and U3618 (N_3618,N_3326,N_3465);
nand U3619 (N_3619,N_3303,N_3440);
nand U3620 (N_3620,N_3081,N_3185);
or U3621 (N_3621,N_3078,N_3061);
nor U3622 (N_3622,N_3022,N_3172);
xnor U3623 (N_3623,N_3075,N_3064);
and U3624 (N_3624,N_3101,N_3194);
nand U3625 (N_3625,N_3192,N_3273);
nand U3626 (N_3626,N_3456,N_3467);
and U3627 (N_3627,N_3057,N_3006);
nor U3628 (N_3628,N_3052,N_3306);
and U3629 (N_3629,N_3016,N_3127);
nor U3630 (N_3630,N_3480,N_3410);
nor U3631 (N_3631,N_3027,N_3387);
nand U3632 (N_3632,N_3210,N_3308);
nor U3633 (N_3633,N_3264,N_3125);
nor U3634 (N_3634,N_3039,N_3454);
and U3635 (N_3635,N_3254,N_3037);
nand U3636 (N_3636,N_3469,N_3344);
and U3637 (N_3637,N_3293,N_3227);
nand U3638 (N_3638,N_3155,N_3385);
nand U3639 (N_3639,N_3168,N_3198);
nor U3640 (N_3640,N_3083,N_3069);
and U3641 (N_3641,N_3280,N_3408);
nand U3642 (N_3642,N_3444,N_3420);
nand U3643 (N_3643,N_3079,N_3373);
or U3644 (N_3644,N_3087,N_3189);
and U3645 (N_3645,N_3416,N_3211);
nor U3646 (N_3646,N_3214,N_3328);
xnor U3647 (N_3647,N_3004,N_3392);
and U3648 (N_3648,N_3165,N_3162);
and U3649 (N_3649,N_3286,N_3325);
and U3650 (N_3650,N_3090,N_3113);
and U3651 (N_3651,N_3186,N_3450);
and U3652 (N_3652,N_3383,N_3073);
and U3653 (N_3653,N_3332,N_3471);
nand U3654 (N_3654,N_3045,N_3041);
nor U3655 (N_3655,N_3008,N_3436);
or U3656 (N_3656,N_3077,N_3453);
or U3657 (N_3657,N_3281,N_3047);
nand U3658 (N_3658,N_3129,N_3274);
and U3659 (N_3659,N_3171,N_3074);
or U3660 (N_3660,N_3441,N_3191);
nand U3661 (N_3661,N_3267,N_3257);
and U3662 (N_3662,N_3055,N_3234);
nor U3663 (N_3663,N_3319,N_3141);
or U3664 (N_3664,N_3201,N_3488);
and U3665 (N_3665,N_3051,N_3094);
nor U3666 (N_3666,N_3132,N_3033);
nand U3667 (N_3667,N_3265,N_3311);
nand U3668 (N_3668,N_3180,N_3283);
nand U3669 (N_3669,N_3212,N_3304);
nor U3670 (N_3670,N_3175,N_3478);
nand U3671 (N_3671,N_3288,N_3431);
and U3672 (N_3672,N_3393,N_3082);
nor U3673 (N_3673,N_3351,N_3412);
and U3674 (N_3674,N_3322,N_3124);
nand U3675 (N_3675,N_3013,N_3343);
and U3676 (N_3676,N_3238,N_3379);
nand U3677 (N_3677,N_3035,N_3368);
nor U3678 (N_3678,N_3230,N_3268);
nand U3679 (N_3679,N_3197,N_3166);
nor U3680 (N_3680,N_3145,N_3401);
and U3681 (N_3681,N_3203,N_3040);
nand U3682 (N_3682,N_3228,N_3489);
nand U3683 (N_3683,N_3358,N_3167);
nand U3684 (N_3684,N_3430,N_3056);
or U3685 (N_3685,N_3023,N_3050);
nor U3686 (N_3686,N_3237,N_3341);
and U3687 (N_3687,N_3269,N_3209);
and U3688 (N_3688,N_3070,N_3103);
xnor U3689 (N_3689,N_3092,N_3063);
and U3690 (N_3690,N_3290,N_3363);
nor U3691 (N_3691,N_3474,N_3472);
or U3692 (N_3692,N_3244,N_3366);
and U3693 (N_3693,N_3058,N_3462);
or U3694 (N_3694,N_3134,N_3259);
nand U3695 (N_3695,N_3121,N_3369);
or U3696 (N_3696,N_3007,N_3356);
xor U3697 (N_3697,N_3036,N_3438);
and U3698 (N_3698,N_3391,N_3105);
nor U3699 (N_3699,N_3102,N_3236);
or U3700 (N_3700,N_3099,N_3220);
nand U3701 (N_3701,N_3426,N_3397);
nand U3702 (N_3702,N_3207,N_3282);
or U3703 (N_3703,N_3206,N_3241);
nor U3704 (N_3704,N_3422,N_3476);
nor U3705 (N_3705,N_3213,N_3159);
xor U3706 (N_3706,N_3400,N_3299);
nor U3707 (N_3707,N_3277,N_3248);
nor U3708 (N_3708,N_3021,N_3160);
and U3709 (N_3709,N_3226,N_3327);
nor U3710 (N_3710,N_3221,N_3375);
nor U3711 (N_3711,N_3096,N_3378);
nor U3712 (N_3712,N_3031,N_3340);
and U3713 (N_3713,N_3398,N_3278);
or U3714 (N_3714,N_3164,N_3190);
nor U3715 (N_3715,N_3150,N_3497);
xor U3716 (N_3716,N_3152,N_3289);
nor U3717 (N_3717,N_3302,N_3095);
and U3718 (N_3718,N_3242,N_3046);
and U3719 (N_3719,N_3399,N_3111);
or U3720 (N_3720,N_3338,N_3417);
nor U3721 (N_3721,N_3019,N_3499);
nor U3722 (N_3722,N_3183,N_3184);
nand U3723 (N_3723,N_3359,N_3048);
and U3724 (N_3724,N_3199,N_3084);
nand U3725 (N_3725,N_3483,N_3246);
nand U3726 (N_3726,N_3485,N_3305);
nand U3727 (N_3727,N_3342,N_3464);
nor U3728 (N_3728,N_3433,N_3346);
or U3729 (N_3729,N_3032,N_3065);
nand U3730 (N_3730,N_3179,N_3312);
nor U3731 (N_3731,N_3067,N_3461);
nand U3732 (N_3732,N_3235,N_3361);
nand U3733 (N_3733,N_3005,N_3053);
nand U3734 (N_3734,N_3225,N_3310);
xnor U3735 (N_3735,N_3010,N_3138);
or U3736 (N_3736,N_3208,N_3014);
or U3737 (N_3737,N_3337,N_3298);
xor U3738 (N_3738,N_3481,N_3271);
nand U3739 (N_3739,N_3223,N_3360);
and U3740 (N_3740,N_3136,N_3187);
nor U3741 (N_3741,N_3459,N_3498);
xnor U3742 (N_3742,N_3353,N_3144);
nor U3743 (N_3743,N_3163,N_3000);
nor U3744 (N_3744,N_3106,N_3458);
and U3745 (N_3745,N_3330,N_3147);
nor U3746 (N_3746,N_3205,N_3182);
xor U3747 (N_3747,N_3009,N_3080);
or U3748 (N_3748,N_3396,N_3245);
xnor U3749 (N_3749,N_3309,N_3345);
or U3750 (N_3750,N_3322,N_3052);
nor U3751 (N_3751,N_3199,N_3082);
nor U3752 (N_3752,N_3278,N_3010);
nor U3753 (N_3753,N_3173,N_3283);
and U3754 (N_3754,N_3070,N_3389);
or U3755 (N_3755,N_3104,N_3270);
or U3756 (N_3756,N_3280,N_3351);
or U3757 (N_3757,N_3130,N_3182);
xnor U3758 (N_3758,N_3267,N_3405);
xor U3759 (N_3759,N_3337,N_3275);
nand U3760 (N_3760,N_3129,N_3283);
or U3761 (N_3761,N_3481,N_3260);
or U3762 (N_3762,N_3435,N_3411);
xnor U3763 (N_3763,N_3281,N_3460);
xor U3764 (N_3764,N_3036,N_3424);
and U3765 (N_3765,N_3097,N_3298);
nand U3766 (N_3766,N_3008,N_3416);
nand U3767 (N_3767,N_3111,N_3274);
and U3768 (N_3768,N_3159,N_3380);
nand U3769 (N_3769,N_3191,N_3227);
nor U3770 (N_3770,N_3174,N_3173);
or U3771 (N_3771,N_3339,N_3103);
nand U3772 (N_3772,N_3435,N_3089);
and U3773 (N_3773,N_3223,N_3239);
and U3774 (N_3774,N_3259,N_3207);
or U3775 (N_3775,N_3214,N_3338);
nor U3776 (N_3776,N_3119,N_3092);
or U3777 (N_3777,N_3155,N_3486);
or U3778 (N_3778,N_3126,N_3085);
nand U3779 (N_3779,N_3328,N_3202);
xnor U3780 (N_3780,N_3224,N_3143);
nor U3781 (N_3781,N_3047,N_3362);
nand U3782 (N_3782,N_3092,N_3205);
nand U3783 (N_3783,N_3254,N_3487);
and U3784 (N_3784,N_3109,N_3324);
nor U3785 (N_3785,N_3018,N_3094);
and U3786 (N_3786,N_3204,N_3054);
and U3787 (N_3787,N_3118,N_3353);
and U3788 (N_3788,N_3136,N_3270);
or U3789 (N_3789,N_3281,N_3344);
nand U3790 (N_3790,N_3409,N_3230);
nor U3791 (N_3791,N_3051,N_3400);
nand U3792 (N_3792,N_3047,N_3382);
and U3793 (N_3793,N_3413,N_3470);
nor U3794 (N_3794,N_3340,N_3415);
or U3795 (N_3795,N_3082,N_3307);
nand U3796 (N_3796,N_3300,N_3275);
nand U3797 (N_3797,N_3165,N_3229);
or U3798 (N_3798,N_3280,N_3337);
xor U3799 (N_3799,N_3483,N_3067);
and U3800 (N_3800,N_3124,N_3381);
and U3801 (N_3801,N_3497,N_3459);
nand U3802 (N_3802,N_3186,N_3077);
nand U3803 (N_3803,N_3081,N_3427);
xnor U3804 (N_3804,N_3453,N_3266);
or U3805 (N_3805,N_3273,N_3255);
or U3806 (N_3806,N_3396,N_3358);
or U3807 (N_3807,N_3274,N_3280);
nand U3808 (N_3808,N_3330,N_3038);
nor U3809 (N_3809,N_3010,N_3448);
or U3810 (N_3810,N_3342,N_3281);
and U3811 (N_3811,N_3008,N_3074);
xor U3812 (N_3812,N_3040,N_3106);
nor U3813 (N_3813,N_3175,N_3473);
and U3814 (N_3814,N_3492,N_3082);
nor U3815 (N_3815,N_3473,N_3158);
nand U3816 (N_3816,N_3239,N_3128);
nand U3817 (N_3817,N_3007,N_3445);
and U3818 (N_3818,N_3122,N_3085);
nor U3819 (N_3819,N_3130,N_3164);
nor U3820 (N_3820,N_3187,N_3213);
or U3821 (N_3821,N_3398,N_3429);
and U3822 (N_3822,N_3443,N_3388);
or U3823 (N_3823,N_3281,N_3313);
nand U3824 (N_3824,N_3469,N_3296);
xnor U3825 (N_3825,N_3147,N_3313);
nand U3826 (N_3826,N_3327,N_3349);
nor U3827 (N_3827,N_3179,N_3246);
nand U3828 (N_3828,N_3420,N_3381);
nand U3829 (N_3829,N_3149,N_3459);
nor U3830 (N_3830,N_3489,N_3362);
nand U3831 (N_3831,N_3194,N_3221);
and U3832 (N_3832,N_3065,N_3320);
nand U3833 (N_3833,N_3427,N_3179);
and U3834 (N_3834,N_3291,N_3358);
nor U3835 (N_3835,N_3423,N_3256);
or U3836 (N_3836,N_3150,N_3151);
nor U3837 (N_3837,N_3029,N_3074);
nand U3838 (N_3838,N_3045,N_3313);
nand U3839 (N_3839,N_3312,N_3085);
and U3840 (N_3840,N_3296,N_3169);
nand U3841 (N_3841,N_3088,N_3092);
xnor U3842 (N_3842,N_3496,N_3065);
nor U3843 (N_3843,N_3420,N_3050);
nor U3844 (N_3844,N_3149,N_3498);
xnor U3845 (N_3845,N_3415,N_3143);
and U3846 (N_3846,N_3014,N_3197);
and U3847 (N_3847,N_3200,N_3092);
xor U3848 (N_3848,N_3329,N_3032);
xor U3849 (N_3849,N_3189,N_3242);
nand U3850 (N_3850,N_3351,N_3458);
nand U3851 (N_3851,N_3458,N_3028);
nand U3852 (N_3852,N_3177,N_3454);
nor U3853 (N_3853,N_3162,N_3343);
nor U3854 (N_3854,N_3263,N_3018);
nand U3855 (N_3855,N_3404,N_3379);
nor U3856 (N_3856,N_3453,N_3290);
nor U3857 (N_3857,N_3054,N_3216);
xnor U3858 (N_3858,N_3272,N_3412);
nor U3859 (N_3859,N_3078,N_3398);
nand U3860 (N_3860,N_3264,N_3163);
and U3861 (N_3861,N_3355,N_3435);
nor U3862 (N_3862,N_3346,N_3141);
nor U3863 (N_3863,N_3161,N_3102);
nor U3864 (N_3864,N_3001,N_3492);
nand U3865 (N_3865,N_3127,N_3373);
and U3866 (N_3866,N_3138,N_3088);
and U3867 (N_3867,N_3376,N_3458);
and U3868 (N_3868,N_3277,N_3193);
or U3869 (N_3869,N_3257,N_3215);
or U3870 (N_3870,N_3399,N_3032);
nand U3871 (N_3871,N_3449,N_3286);
or U3872 (N_3872,N_3309,N_3223);
nor U3873 (N_3873,N_3303,N_3159);
or U3874 (N_3874,N_3089,N_3108);
nand U3875 (N_3875,N_3262,N_3143);
or U3876 (N_3876,N_3357,N_3463);
nand U3877 (N_3877,N_3498,N_3132);
or U3878 (N_3878,N_3375,N_3257);
or U3879 (N_3879,N_3298,N_3340);
or U3880 (N_3880,N_3376,N_3274);
or U3881 (N_3881,N_3068,N_3425);
nor U3882 (N_3882,N_3155,N_3412);
nand U3883 (N_3883,N_3452,N_3028);
or U3884 (N_3884,N_3103,N_3473);
nand U3885 (N_3885,N_3008,N_3306);
nand U3886 (N_3886,N_3302,N_3127);
or U3887 (N_3887,N_3086,N_3450);
xor U3888 (N_3888,N_3181,N_3021);
and U3889 (N_3889,N_3464,N_3267);
nand U3890 (N_3890,N_3015,N_3175);
or U3891 (N_3891,N_3298,N_3243);
and U3892 (N_3892,N_3423,N_3322);
or U3893 (N_3893,N_3002,N_3443);
nor U3894 (N_3894,N_3079,N_3321);
and U3895 (N_3895,N_3062,N_3120);
or U3896 (N_3896,N_3259,N_3125);
or U3897 (N_3897,N_3376,N_3405);
or U3898 (N_3898,N_3235,N_3106);
or U3899 (N_3899,N_3293,N_3284);
nand U3900 (N_3900,N_3143,N_3384);
and U3901 (N_3901,N_3382,N_3399);
nand U3902 (N_3902,N_3113,N_3084);
or U3903 (N_3903,N_3093,N_3039);
nand U3904 (N_3904,N_3353,N_3469);
and U3905 (N_3905,N_3318,N_3449);
xor U3906 (N_3906,N_3401,N_3120);
nor U3907 (N_3907,N_3427,N_3038);
nor U3908 (N_3908,N_3393,N_3154);
or U3909 (N_3909,N_3276,N_3263);
and U3910 (N_3910,N_3376,N_3146);
nor U3911 (N_3911,N_3027,N_3032);
or U3912 (N_3912,N_3390,N_3309);
and U3913 (N_3913,N_3462,N_3454);
nor U3914 (N_3914,N_3271,N_3402);
nor U3915 (N_3915,N_3477,N_3272);
and U3916 (N_3916,N_3496,N_3010);
xnor U3917 (N_3917,N_3274,N_3237);
and U3918 (N_3918,N_3020,N_3184);
nand U3919 (N_3919,N_3417,N_3093);
nor U3920 (N_3920,N_3069,N_3342);
and U3921 (N_3921,N_3139,N_3032);
xnor U3922 (N_3922,N_3296,N_3265);
nor U3923 (N_3923,N_3386,N_3292);
and U3924 (N_3924,N_3277,N_3309);
and U3925 (N_3925,N_3271,N_3208);
or U3926 (N_3926,N_3180,N_3356);
or U3927 (N_3927,N_3244,N_3264);
or U3928 (N_3928,N_3418,N_3056);
xnor U3929 (N_3929,N_3494,N_3275);
or U3930 (N_3930,N_3352,N_3441);
nor U3931 (N_3931,N_3212,N_3150);
and U3932 (N_3932,N_3238,N_3442);
and U3933 (N_3933,N_3443,N_3157);
nand U3934 (N_3934,N_3481,N_3168);
xnor U3935 (N_3935,N_3311,N_3132);
and U3936 (N_3936,N_3331,N_3217);
or U3937 (N_3937,N_3253,N_3341);
or U3938 (N_3938,N_3195,N_3277);
or U3939 (N_3939,N_3157,N_3058);
or U3940 (N_3940,N_3484,N_3110);
nor U3941 (N_3941,N_3025,N_3037);
and U3942 (N_3942,N_3413,N_3468);
or U3943 (N_3943,N_3491,N_3442);
or U3944 (N_3944,N_3126,N_3333);
or U3945 (N_3945,N_3386,N_3345);
nand U3946 (N_3946,N_3461,N_3052);
and U3947 (N_3947,N_3052,N_3153);
or U3948 (N_3948,N_3129,N_3169);
nand U3949 (N_3949,N_3332,N_3171);
and U3950 (N_3950,N_3009,N_3325);
nand U3951 (N_3951,N_3033,N_3131);
nand U3952 (N_3952,N_3161,N_3492);
and U3953 (N_3953,N_3068,N_3423);
or U3954 (N_3954,N_3073,N_3044);
nor U3955 (N_3955,N_3092,N_3484);
nand U3956 (N_3956,N_3410,N_3319);
nor U3957 (N_3957,N_3262,N_3123);
or U3958 (N_3958,N_3370,N_3314);
and U3959 (N_3959,N_3485,N_3051);
nor U3960 (N_3960,N_3120,N_3033);
or U3961 (N_3961,N_3068,N_3064);
xnor U3962 (N_3962,N_3367,N_3088);
xnor U3963 (N_3963,N_3240,N_3063);
nand U3964 (N_3964,N_3312,N_3188);
xor U3965 (N_3965,N_3378,N_3119);
xnor U3966 (N_3966,N_3067,N_3264);
nand U3967 (N_3967,N_3272,N_3293);
nand U3968 (N_3968,N_3035,N_3026);
and U3969 (N_3969,N_3387,N_3344);
nor U3970 (N_3970,N_3196,N_3010);
and U3971 (N_3971,N_3045,N_3315);
and U3972 (N_3972,N_3122,N_3361);
nor U3973 (N_3973,N_3364,N_3174);
or U3974 (N_3974,N_3040,N_3190);
nand U3975 (N_3975,N_3457,N_3092);
xor U3976 (N_3976,N_3151,N_3370);
or U3977 (N_3977,N_3429,N_3361);
xnor U3978 (N_3978,N_3124,N_3299);
nand U3979 (N_3979,N_3244,N_3418);
or U3980 (N_3980,N_3141,N_3101);
and U3981 (N_3981,N_3264,N_3094);
or U3982 (N_3982,N_3497,N_3089);
and U3983 (N_3983,N_3284,N_3438);
nor U3984 (N_3984,N_3375,N_3154);
nor U3985 (N_3985,N_3109,N_3495);
or U3986 (N_3986,N_3142,N_3148);
nand U3987 (N_3987,N_3131,N_3453);
and U3988 (N_3988,N_3274,N_3489);
or U3989 (N_3989,N_3198,N_3381);
nand U3990 (N_3990,N_3460,N_3434);
nand U3991 (N_3991,N_3062,N_3458);
nor U3992 (N_3992,N_3378,N_3137);
nand U3993 (N_3993,N_3458,N_3461);
nor U3994 (N_3994,N_3345,N_3025);
or U3995 (N_3995,N_3389,N_3233);
or U3996 (N_3996,N_3111,N_3394);
nor U3997 (N_3997,N_3074,N_3196);
and U3998 (N_3998,N_3174,N_3335);
nand U3999 (N_3999,N_3232,N_3082);
and U4000 (N_4000,N_3523,N_3917);
and U4001 (N_4001,N_3576,N_3532);
and U4002 (N_4002,N_3707,N_3589);
and U4003 (N_4003,N_3887,N_3559);
nand U4004 (N_4004,N_3739,N_3876);
and U4005 (N_4005,N_3974,N_3776);
or U4006 (N_4006,N_3905,N_3964);
nand U4007 (N_4007,N_3697,N_3967);
nor U4008 (N_4008,N_3795,N_3823);
nand U4009 (N_4009,N_3954,N_3543);
and U4010 (N_4010,N_3839,N_3560);
or U4011 (N_4011,N_3835,N_3716);
nor U4012 (N_4012,N_3616,N_3551);
nand U4013 (N_4013,N_3761,N_3718);
or U4014 (N_4014,N_3965,N_3838);
nor U4015 (N_4015,N_3665,N_3524);
nand U4016 (N_4016,N_3908,N_3705);
and U4017 (N_4017,N_3787,N_3564);
or U4018 (N_4018,N_3521,N_3780);
nand U4019 (N_4019,N_3614,N_3683);
or U4020 (N_4020,N_3874,N_3599);
nand U4021 (N_4021,N_3734,N_3552);
and U4022 (N_4022,N_3775,N_3594);
nor U4023 (N_4023,N_3586,N_3726);
or U4024 (N_4024,N_3558,N_3990);
or U4025 (N_4025,N_3955,N_3582);
and U4026 (N_4026,N_3737,N_3746);
xor U4027 (N_4027,N_3538,N_3900);
and U4028 (N_4028,N_3617,N_3536);
nor U4029 (N_4029,N_3638,N_3960);
and U4030 (N_4030,N_3933,N_3983);
and U4031 (N_4031,N_3506,N_3592);
or U4032 (N_4032,N_3818,N_3744);
or U4033 (N_4033,N_3731,N_3914);
nor U4034 (N_4034,N_3676,N_3922);
and U4035 (N_4035,N_3939,N_3587);
nor U4036 (N_4036,N_3534,N_3685);
nand U4037 (N_4037,N_3843,N_3752);
xnor U4038 (N_4038,N_3958,N_3959);
xnor U4039 (N_4039,N_3608,N_3633);
nand U4040 (N_4040,N_3637,N_3711);
nor U4041 (N_4041,N_3831,N_3580);
nor U4042 (N_4042,N_3836,N_3710);
nand U4043 (N_4043,N_3845,N_3653);
or U4044 (N_4044,N_3590,N_3700);
xor U4045 (N_4045,N_3569,N_3813);
and U4046 (N_4046,N_3522,N_3973);
and U4047 (N_4047,N_3878,N_3913);
and U4048 (N_4048,N_3918,N_3751);
and U4049 (N_4049,N_3544,N_3798);
and U4050 (N_4050,N_3669,N_3858);
or U4051 (N_4051,N_3931,N_3722);
nor U4052 (N_4052,N_3791,N_3814);
or U4053 (N_4053,N_3745,N_3846);
or U4054 (N_4054,N_3689,N_3636);
and U4055 (N_4055,N_3598,N_3585);
nor U4056 (N_4056,N_3777,N_3565);
and U4057 (N_4057,N_3894,N_3794);
xnor U4058 (N_4058,N_3859,N_3597);
and U4059 (N_4059,N_3654,N_3850);
and U4060 (N_4060,N_3796,N_3934);
nor U4061 (N_4061,N_3873,N_3971);
nor U4062 (N_4062,N_3600,N_3588);
or U4063 (N_4063,N_3982,N_3574);
xnor U4064 (N_4064,N_3517,N_3822);
or U4065 (N_4065,N_3920,N_3889);
nand U4066 (N_4066,N_3748,N_3627);
or U4067 (N_4067,N_3531,N_3675);
nor U4068 (N_4068,N_3800,N_3852);
nand U4069 (N_4069,N_3735,N_3644);
and U4070 (N_4070,N_3789,N_3805);
or U4071 (N_4071,N_3528,N_3602);
or U4072 (N_4072,N_3634,N_3969);
or U4073 (N_4073,N_3884,N_3891);
nor U4074 (N_4074,N_3862,N_3540);
nor U4075 (N_4075,N_3757,N_3578);
nor U4076 (N_4076,N_3663,N_3773);
nor U4077 (N_4077,N_3994,N_3754);
or U4078 (N_4078,N_3662,N_3916);
and U4079 (N_4079,N_3961,N_3631);
nor U4080 (N_4080,N_3659,N_3952);
nand U4081 (N_4081,N_3962,N_3868);
nor U4082 (N_4082,N_3615,N_3504);
nand U4083 (N_4083,N_3713,N_3801);
xnor U4084 (N_4084,N_3628,N_3996);
nand U4085 (N_4085,N_3768,N_3643);
and U4086 (N_4086,N_3998,N_3925);
nand U4087 (N_4087,N_3696,N_3979);
nand U4088 (N_4088,N_3833,N_3886);
nor U4089 (N_4089,N_3949,N_3946);
xnor U4090 (N_4090,N_3826,N_3691);
nor U4091 (N_4091,N_3802,N_3968);
nand U4092 (N_4092,N_3724,N_3820);
and U4093 (N_4093,N_3537,N_3601);
or U4094 (N_4094,N_3812,N_3516);
nand U4095 (N_4095,N_3824,N_3661);
and U4096 (N_4096,N_3907,N_3561);
or U4097 (N_4097,N_3526,N_3834);
or U4098 (N_4098,N_3975,N_3674);
or U4099 (N_4099,N_3758,N_3603);
nor U4100 (N_4100,N_3658,N_3557);
nand U4101 (N_4101,N_3687,N_3869);
nor U4102 (N_4102,N_3810,N_3989);
nor U4103 (N_4103,N_3875,N_3942);
and U4104 (N_4104,N_3756,N_3732);
nor U4105 (N_4105,N_3511,N_3766);
and U4106 (N_4106,N_3575,N_3695);
and U4107 (N_4107,N_3699,N_3855);
nand U4108 (N_4108,N_3986,N_3945);
or U4109 (N_4109,N_3741,N_3844);
and U4110 (N_4110,N_3932,N_3510);
nor U4111 (N_4111,N_3577,N_3977);
or U4112 (N_4112,N_3803,N_3678);
and U4113 (N_4113,N_3503,N_3790);
xnor U4114 (N_4114,N_3611,N_3688);
nor U4115 (N_4115,N_3553,N_3623);
or U4116 (N_4116,N_3624,N_3879);
nand U4117 (N_4117,N_3743,N_3704);
and U4118 (N_4118,N_3893,N_3596);
and U4119 (N_4119,N_3515,N_3882);
nand U4120 (N_4120,N_3811,N_3672);
or U4121 (N_4121,N_3910,N_3657);
or U4122 (N_4122,N_3865,N_3840);
and U4123 (N_4123,N_3583,N_3618);
xor U4124 (N_4124,N_3930,N_3619);
nand U4125 (N_4125,N_3963,N_3926);
xnor U4126 (N_4126,N_3928,N_3815);
and U4127 (N_4127,N_3807,N_3613);
or U4128 (N_4128,N_3702,N_3727);
nand U4129 (N_4129,N_3548,N_3730);
or U4130 (N_4130,N_3866,N_3929);
and U4131 (N_4131,N_3682,N_3625);
nand U4132 (N_4132,N_3629,N_3648);
xor U4133 (N_4133,N_3539,N_3817);
nand U4134 (N_4134,N_3693,N_3857);
nor U4135 (N_4135,N_3966,N_3556);
and U4136 (N_4136,N_3924,N_3837);
and U4137 (N_4137,N_3830,N_3632);
or U4138 (N_4138,N_3686,N_3981);
or U4139 (N_4139,N_3976,N_3502);
nor U4140 (N_4140,N_3860,N_3991);
nand U4141 (N_4141,N_3750,N_3793);
nor U4142 (N_4142,N_3896,N_3867);
nor U4143 (N_4143,N_3806,N_3970);
nor U4144 (N_4144,N_3956,N_3980);
xor U4145 (N_4145,N_3808,N_3771);
nand U4146 (N_4146,N_3856,N_3892);
nor U4147 (N_4147,N_3546,N_3995);
nor U4148 (N_4148,N_3703,N_3880);
nor U4149 (N_4149,N_3783,N_3620);
nor U4150 (N_4150,N_3512,N_3717);
and U4151 (N_4151,N_3870,N_3904);
nor U4152 (N_4152,N_3725,N_3584);
nor U4153 (N_4153,N_3864,N_3909);
nand U4154 (N_4154,N_3753,N_3759);
nand U4155 (N_4155,N_3827,N_3919);
nor U4156 (N_4156,N_3505,N_3709);
nand U4157 (N_4157,N_3606,N_3667);
and U4158 (N_4158,N_3792,N_3719);
nor U4159 (N_4159,N_3819,N_3897);
nor U4160 (N_4160,N_3947,N_3572);
nand U4161 (N_4161,N_3728,N_3736);
and U4162 (N_4162,N_3677,N_3906);
nor U4163 (N_4163,N_3554,N_3591);
nand U4164 (N_4164,N_3579,N_3723);
xnor U4165 (N_4165,N_3530,N_3755);
xor U4166 (N_4166,N_3821,N_3849);
nor U4167 (N_4167,N_3635,N_3763);
or U4168 (N_4168,N_3993,N_3593);
nand U4169 (N_4169,N_3923,N_3733);
and U4170 (N_4170,N_3988,N_3936);
or U4171 (N_4171,N_3545,N_3640);
and U4172 (N_4172,N_3642,N_3652);
and U4173 (N_4173,N_3622,N_3927);
and U4174 (N_4174,N_3828,N_3851);
and U4175 (N_4175,N_3681,N_3568);
nor U4176 (N_4176,N_3694,N_3720);
nor U4177 (N_4177,N_3816,N_3533);
xor U4178 (N_4178,N_3872,N_3895);
and U4179 (N_4179,N_3951,N_3938);
nor U4180 (N_4180,N_3769,N_3649);
or U4181 (N_4181,N_3679,N_3604);
xnor U4182 (N_4182,N_3782,N_3680);
or U4183 (N_4183,N_3941,N_3525);
xor U4184 (N_4184,N_3809,N_3765);
nor U4185 (N_4185,N_3829,N_3890);
or U4186 (N_4186,N_3507,N_3549);
xnor U4187 (N_4187,N_3785,N_3854);
and U4188 (N_4188,N_3797,N_3784);
nor U4189 (N_4189,N_3671,N_3607);
and U4190 (N_4190,N_3563,N_3999);
or U4191 (N_4191,N_3901,N_3706);
and U4192 (N_4192,N_3562,N_3509);
nor U4193 (N_4193,N_3762,N_3985);
or U4194 (N_4194,N_3639,N_3921);
xor U4195 (N_4195,N_3647,N_3770);
nor U4196 (N_4196,N_3668,N_3935);
or U4197 (N_4197,N_3605,N_3595);
nor U4198 (N_4198,N_3774,N_3881);
nand U4199 (N_4199,N_3612,N_3641);
xor U4200 (N_4200,N_3764,N_3567);
nand U4201 (N_4201,N_3953,N_3804);
nor U4202 (N_4202,N_3684,N_3883);
or U4203 (N_4203,N_3863,N_3972);
nand U4204 (N_4204,N_3848,N_3767);
or U4205 (N_4205,N_3656,N_3626);
nor U4206 (N_4206,N_3853,N_3609);
nand U4207 (N_4207,N_3902,N_3573);
and U4208 (N_4208,N_3943,N_3708);
nand U4209 (N_4209,N_3721,N_3651);
and U4210 (N_4210,N_3948,N_3690);
nor U4211 (N_4211,N_3772,N_3666);
or U4212 (N_4212,N_3660,N_3714);
nand U4213 (N_4213,N_3729,N_3501);
nand U4214 (N_4214,N_3841,N_3978);
xor U4215 (N_4215,N_3911,N_3987);
nor U4216 (N_4216,N_3646,N_3547);
and U4217 (N_4217,N_3937,N_3738);
and U4218 (N_4218,N_3610,N_3747);
or U4219 (N_4219,N_3519,N_3566);
or U4220 (N_4220,N_3541,N_3555);
nor U4221 (N_4221,N_3899,N_3645);
and U4222 (N_4222,N_3779,N_3915);
xnor U4223 (N_4223,N_3514,N_3992);
nor U4224 (N_4224,N_3542,N_3997);
or U4225 (N_4225,N_3957,N_3701);
xnor U4226 (N_4226,N_3842,N_3571);
or U4227 (N_4227,N_3527,N_3799);
or U4228 (N_4228,N_3740,N_3749);
nor U4229 (N_4229,N_3535,N_3698);
and U4230 (N_4230,N_3786,N_3944);
nand U4231 (N_4231,N_3912,N_3781);
nand U4232 (N_4232,N_3898,N_3984);
or U4233 (N_4233,N_3861,N_3650);
and U4234 (N_4234,N_3570,N_3788);
nand U4235 (N_4235,N_3940,N_3655);
nor U4236 (N_4236,N_3621,N_3903);
nand U4237 (N_4237,N_3513,N_3885);
nand U4238 (N_4238,N_3550,N_3888);
and U4239 (N_4239,N_3670,N_3950);
nor U4240 (N_4240,N_3518,N_3520);
and U4241 (N_4241,N_3508,N_3847);
nor U4242 (N_4242,N_3630,N_3778);
nor U4243 (N_4243,N_3832,N_3712);
nor U4244 (N_4244,N_3529,N_3500);
xnor U4245 (N_4245,N_3664,N_3581);
nand U4246 (N_4246,N_3760,N_3673);
xor U4247 (N_4247,N_3825,N_3877);
nand U4248 (N_4248,N_3715,N_3692);
nor U4249 (N_4249,N_3742,N_3871);
nor U4250 (N_4250,N_3969,N_3636);
nor U4251 (N_4251,N_3785,N_3777);
or U4252 (N_4252,N_3959,N_3695);
or U4253 (N_4253,N_3568,N_3992);
or U4254 (N_4254,N_3579,N_3662);
nor U4255 (N_4255,N_3966,N_3540);
nor U4256 (N_4256,N_3548,N_3643);
nor U4257 (N_4257,N_3752,N_3552);
or U4258 (N_4258,N_3965,N_3945);
and U4259 (N_4259,N_3881,N_3648);
and U4260 (N_4260,N_3554,N_3983);
or U4261 (N_4261,N_3716,N_3679);
xnor U4262 (N_4262,N_3704,N_3979);
nor U4263 (N_4263,N_3861,N_3888);
nand U4264 (N_4264,N_3855,N_3796);
or U4265 (N_4265,N_3731,N_3843);
nand U4266 (N_4266,N_3851,N_3921);
nor U4267 (N_4267,N_3922,N_3900);
and U4268 (N_4268,N_3540,N_3946);
and U4269 (N_4269,N_3778,N_3539);
nor U4270 (N_4270,N_3951,N_3580);
nor U4271 (N_4271,N_3993,N_3575);
or U4272 (N_4272,N_3571,N_3604);
and U4273 (N_4273,N_3755,N_3750);
or U4274 (N_4274,N_3668,N_3932);
nand U4275 (N_4275,N_3827,N_3872);
nor U4276 (N_4276,N_3657,N_3676);
nand U4277 (N_4277,N_3959,N_3799);
nor U4278 (N_4278,N_3643,N_3611);
nor U4279 (N_4279,N_3999,N_3885);
and U4280 (N_4280,N_3529,N_3948);
or U4281 (N_4281,N_3602,N_3795);
and U4282 (N_4282,N_3898,N_3693);
nor U4283 (N_4283,N_3879,N_3759);
or U4284 (N_4284,N_3656,N_3641);
nand U4285 (N_4285,N_3688,N_3598);
nand U4286 (N_4286,N_3554,N_3612);
and U4287 (N_4287,N_3521,N_3949);
or U4288 (N_4288,N_3953,N_3918);
nor U4289 (N_4289,N_3720,N_3615);
and U4290 (N_4290,N_3757,N_3986);
and U4291 (N_4291,N_3580,N_3755);
and U4292 (N_4292,N_3648,N_3718);
nand U4293 (N_4293,N_3768,N_3937);
nor U4294 (N_4294,N_3987,N_3830);
nand U4295 (N_4295,N_3731,N_3933);
and U4296 (N_4296,N_3717,N_3964);
and U4297 (N_4297,N_3570,N_3851);
xor U4298 (N_4298,N_3852,N_3901);
or U4299 (N_4299,N_3852,N_3836);
and U4300 (N_4300,N_3799,N_3888);
or U4301 (N_4301,N_3618,N_3740);
nor U4302 (N_4302,N_3697,N_3966);
and U4303 (N_4303,N_3689,N_3668);
and U4304 (N_4304,N_3742,N_3886);
and U4305 (N_4305,N_3857,N_3735);
nor U4306 (N_4306,N_3613,N_3737);
nor U4307 (N_4307,N_3959,N_3522);
and U4308 (N_4308,N_3661,N_3569);
and U4309 (N_4309,N_3546,N_3775);
and U4310 (N_4310,N_3882,N_3708);
nor U4311 (N_4311,N_3798,N_3690);
nor U4312 (N_4312,N_3772,N_3544);
and U4313 (N_4313,N_3525,N_3968);
or U4314 (N_4314,N_3863,N_3965);
nand U4315 (N_4315,N_3607,N_3774);
nor U4316 (N_4316,N_3959,N_3705);
and U4317 (N_4317,N_3801,N_3718);
nand U4318 (N_4318,N_3638,N_3860);
nor U4319 (N_4319,N_3876,N_3708);
nand U4320 (N_4320,N_3598,N_3828);
and U4321 (N_4321,N_3726,N_3643);
nor U4322 (N_4322,N_3530,N_3811);
nand U4323 (N_4323,N_3674,N_3698);
xor U4324 (N_4324,N_3678,N_3744);
nor U4325 (N_4325,N_3732,N_3850);
and U4326 (N_4326,N_3975,N_3638);
nand U4327 (N_4327,N_3834,N_3704);
nand U4328 (N_4328,N_3838,N_3933);
or U4329 (N_4329,N_3685,N_3691);
xnor U4330 (N_4330,N_3524,N_3900);
nand U4331 (N_4331,N_3501,N_3540);
or U4332 (N_4332,N_3945,N_3645);
or U4333 (N_4333,N_3506,N_3903);
xor U4334 (N_4334,N_3821,N_3818);
and U4335 (N_4335,N_3599,N_3586);
or U4336 (N_4336,N_3632,N_3812);
and U4337 (N_4337,N_3654,N_3673);
or U4338 (N_4338,N_3673,N_3546);
nand U4339 (N_4339,N_3551,N_3783);
nor U4340 (N_4340,N_3548,N_3626);
and U4341 (N_4341,N_3941,N_3717);
or U4342 (N_4342,N_3512,N_3740);
nor U4343 (N_4343,N_3987,N_3557);
nor U4344 (N_4344,N_3872,N_3759);
or U4345 (N_4345,N_3896,N_3812);
or U4346 (N_4346,N_3529,N_3535);
nand U4347 (N_4347,N_3991,N_3649);
nor U4348 (N_4348,N_3728,N_3743);
or U4349 (N_4349,N_3603,N_3905);
nand U4350 (N_4350,N_3929,N_3731);
or U4351 (N_4351,N_3637,N_3994);
nand U4352 (N_4352,N_3600,N_3883);
and U4353 (N_4353,N_3794,N_3854);
and U4354 (N_4354,N_3793,N_3702);
xor U4355 (N_4355,N_3881,N_3853);
and U4356 (N_4356,N_3582,N_3846);
and U4357 (N_4357,N_3750,N_3587);
xor U4358 (N_4358,N_3888,N_3896);
nor U4359 (N_4359,N_3970,N_3856);
nor U4360 (N_4360,N_3847,N_3977);
and U4361 (N_4361,N_3724,N_3950);
nor U4362 (N_4362,N_3886,N_3508);
or U4363 (N_4363,N_3651,N_3756);
and U4364 (N_4364,N_3839,N_3640);
nand U4365 (N_4365,N_3508,N_3869);
and U4366 (N_4366,N_3854,N_3645);
or U4367 (N_4367,N_3826,N_3643);
or U4368 (N_4368,N_3958,N_3919);
or U4369 (N_4369,N_3687,N_3650);
nand U4370 (N_4370,N_3787,N_3900);
nor U4371 (N_4371,N_3806,N_3917);
and U4372 (N_4372,N_3748,N_3641);
nor U4373 (N_4373,N_3754,N_3979);
or U4374 (N_4374,N_3638,N_3672);
xnor U4375 (N_4375,N_3930,N_3631);
nand U4376 (N_4376,N_3562,N_3739);
and U4377 (N_4377,N_3753,N_3679);
or U4378 (N_4378,N_3818,N_3657);
nor U4379 (N_4379,N_3583,N_3606);
xnor U4380 (N_4380,N_3708,N_3538);
nand U4381 (N_4381,N_3519,N_3824);
nor U4382 (N_4382,N_3785,N_3807);
nand U4383 (N_4383,N_3954,N_3820);
and U4384 (N_4384,N_3544,N_3522);
or U4385 (N_4385,N_3852,N_3619);
and U4386 (N_4386,N_3694,N_3932);
or U4387 (N_4387,N_3532,N_3881);
or U4388 (N_4388,N_3555,N_3856);
nor U4389 (N_4389,N_3515,N_3742);
and U4390 (N_4390,N_3515,N_3627);
and U4391 (N_4391,N_3919,N_3807);
nor U4392 (N_4392,N_3732,N_3635);
and U4393 (N_4393,N_3807,N_3585);
nand U4394 (N_4394,N_3741,N_3637);
nand U4395 (N_4395,N_3614,N_3695);
nand U4396 (N_4396,N_3795,N_3569);
and U4397 (N_4397,N_3618,N_3615);
xnor U4398 (N_4398,N_3509,N_3791);
xnor U4399 (N_4399,N_3588,N_3960);
and U4400 (N_4400,N_3877,N_3523);
nor U4401 (N_4401,N_3817,N_3981);
and U4402 (N_4402,N_3528,N_3550);
or U4403 (N_4403,N_3730,N_3713);
or U4404 (N_4404,N_3711,N_3726);
nor U4405 (N_4405,N_3673,N_3553);
nor U4406 (N_4406,N_3931,N_3510);
or U4407 (N_4407,N_3881,N_3571);
or U4408 (N_4408,N_3777,N_3567);
nor U4409 (N_4409,N_3932,N_3509);
nand U4410 (N_4410,N_3584,N_3790);
nand U4411 (N_4411,N_3676,N_3517);
nand U4412 (N_4412,N_3958,N_3629);
xnor U4413 (N_4413,N_3653,N_3685);
nor U4414 (N_4414,N_3536,N_3576);
nand U4415 (N_4415,N_3636,N_3975);
nand U4416 (N_4416,N_3948,N_3507);
or U4417 (N_4417,N_3736,N_3887);
nand U4418 (N_4418,N_3901,N_3567);
nand U4419 (N_4419,N_3893,N_3781);
nand U4420 (N_4420,N_3734,N_3619);
and U4421 (N_4421,N_3625,N_3665);
nand U4422 (N_4422,N_3567,N_3737);
nor U4423 (N_4423,N_3671,N_3829);
nand U4424 (N_4424,N_3641,N_3996);
and U4425 (N_4425,N_3581,N_3891);
nand U4426 (N_4426,N_3792,N_3897);
nor U4427 (N_4427,N_3854,N_3707);
nand U4428 (N_4428,N_3577,N_3521);
or U4429 (N_4429,N_3620,N_3708);
and U4430 (N_4430,N_3653,N_3702);
and U4431 (N_4431,N_3641,N_3525);
nand U4432 (N_4432,N_3840,N_3883);
or U4433 (N_4433,N_3751,N_3547);
or U4434 (N_4434,N_3592,N_3843);
or U4435 (N_4435,N_3778,N_3785);
or U4436 (N_4436,N_3503,N_3637);
nand U4437 (N_4437,N_3763,N_3938);
nand U4438 (N_4438,N_3620,N_3841);
or U4439 (N_4439,N_3874,N_3861);
or U4440 (N_4440,N_3773,N_3754);
and U4441 (N_4441,N_3654,N_3610);
and U4442 (N_4442,N_3500,N_3986);
or U4443 (N_4443,N_3716,N_3525);
and U4444 (N_4444,N_3690,N_3894);
or U4445 (N_4445,N_3512,N_3627);
xor U4446 (N_4446,N_3896,N_3576);
nor U4447 (N_4447,N_3851,N_3947);
xnor U4448 (N_4448,N_3691,N_3618);
nor U4449 (N_4449,N_3806,N_3595);
and U4450 (N_4450,N_3791,N_3807);
nor U4451 (N_4451,N_3792,N_3501);
nand U4452 (N_4452,N_3677,N_3774);
nor U4453 (N_4453,N_3640,N_3993);
and U4454 (N_4454,N_3909,N_3876);
nand U4455 (N_4455,N_3737,N_3741);
nor U4456 (N_4456,N_3709,N_3950);
and U4457 (N_4457,N_3542,N_3659);
or U4458 (N_4458,N_3965,N_3510);
xnor U4459 (N_4459,N_3515,N_3790);
nand U4460 (N_4460,N_3969,N_3539);
and U4461 (N_4461,N_3972,N_3854);
nand U4462 (N_4462,N_3738,N_3584);
or U4463 (N_4463,N_3686,N_3533);
or U4464 (N_4464,N_3533,N_3952);
or U4465 (N_4465,N_3745,N_3588);
nor U4466 (N_4466,N_3590,N_3594);
or U4467 (N_4467,N_3825,N_3758);
or U4468 (N_4468,N_3703,N_3899);
nand U4469 (N_4469,N_3700,N_3833);
xor U4470 (N_4470,N_3858,N_3815);
nand U4471 (N_4471,N_3745,N_3999);
nand U4472 (N_4472,N_3631,N_3556);
or U4473 (N_4473,N_3826,N_3956);
or U4474 (N_4474,N_3813,N_3603);
or U4475 (N_4475,N_3627,N_3842);
or U4476 (N_4476,N_3645,N_3595);
nand U4477 (N_4477,N_3979,N_3640);
nand U4478 (N_4478,N_3817,N_3875);
xor U4479 (N_4479,N_3693,N_3629);
xor U4480 (N_4480,N_3780,N_3625);
or U4481 (N_4481,N_3563,N_3990);
or U4482 (N_4482,N_3598,N_3508);
nand U4483 (N_4483,N_3589,N_3879);
xnor U4484 (N_4484,N_3915,N_3586);
and U4485 (N_4485,N_3831,N_3853);
nand U4486 (N_4486,N_3501,N_3887);
xor U4487 (N_4487,N_3546,N_3958);
and U4488 (N_4488,N_3912,N_3780);
nor U4489 (N_4489,N_3728,N_3742);
nand U4490 (N_4490,N_3982,N_3821);
or U4491 (N_4491,N_3961,N_3920);
xor U4492 (N_4492,N_3998,N_3988);
and U4493 (N_4493,N_3857,N_3847);
nand U4494 (N_4494,N_3669,N_3572);
nor U4495 (N_4495,N_3769,N_3978);
and U4496 (N_4496,N_3689,N_3796);
nand U4497 (N_4497,N_3886,N_3831);
nand U4498 (N_4498,N_3507,N_3803);
or U4499 (N_4499,N_3742,N_3889);
nor U4500 (N_4500,N_4288,N_4037);
and U4501 (N_4501,N_4041,N_4058);
nor U4502 (N_4502,N_4307,N_4324);
and U4503 (N_4503,N_4151,N_4239);
nand U4504 (N_4504,N_4321,N_4488);
and U4505 (N_4505,N_4344,N_4070);
or U4506 (N_4506,N_4049,N_4407);
and U4507 (N_4507,N_4034,N_4461);
xnor U4508 (N_4508,N_4099,N_4458);
xnor U4509 (N_4509,N_4271,N_4095);
xnor U4510 (N_4510,N_4465,N_4101);
nor U4511 (N_4511,N_4399,N_4112);
nor U4512 (N_4512,N_4255,N_4451);
or U4513 (N_4513,N_4043,N_4483);
or U4514 (N_4514,N_4369,N_4357);
and U4515 (N_4515,N_4146,N_4349);
nor U4516 (N_4516,N_4150,N_4286);
nor U4517 (N_4517,N_4082,N_4012);
nand U4518 (N_4518,N_4092,N_4309);
nand U4519 (N_4519,N_4019,N_4044);
or U4520 (N_4520,N_4246,N_4148);
nor U4521 (N_4521,N_4475,N_4484);
nand U4522 (N_4522,N_4232,N_4218);
xor U4523 (N_4523,N_4200,N_4311);
nand U4524 (N_4524,N_4224,N_4259);
xnor U4525 (N_4525,N_4220,N_4040);
nor U4526 (N_4526,N_4030,N_4366);
nand U4527 (N_4527,N_4219,N_4069);
or U4528 (N_4528,N_4384,N_4116);
or U4529 (N_4529,N_4478,N_4157);
or U4530 (N_4530,N_4277,N_4121);
or U4531 (N_4531,N_4492,N_4308);
or U4532 (N_4532,N_4105,N_4430);
nand U4533 (N_4533,N_4310,N_4292);
or U4534 (N_4534,N_4236,N_4432);
and U4535 (N_4535,N_4173,N_4153);
nor U4536 (N_4536,N_4242,N_4108);
nor U4537 (N_4537,N_4325,N_4167);
xnor U4538 (N_4538,N_4390,N_4036);
and U4539 (N_4539,N_4193,N_4028);
xnor U4540 (N_4540,N_4360,N_4139);
and U4541 (N_4541,N_4001,N_4000);
and U4542 (N_4542,N_4210,N_4102);
or U4543 (N_4543,N_4206,N_4476);
or U4544 (N_4544,N_4493,N_4039);
and U4545 (N_4545,N_4053,N_4268);
xnor U4546 (N_4546,N_4184,N_4439);
and U4547 (N_4547,N_4107,N_4298);
xnor U4548 (N_4548,N_4133,N_4353);
nand U4549 (N_4549,N_4079,N_4134);
or U4550 (N_4550,N_4482,N_4051);
nor U4551 (N_4551,N_4245,N_4389);
nor U4552 (N_4552,N_4331,N_4033);
and U4553 (N_4553,N_4008,N_4428);
nand U4554 (N_4554,N_4472,N_4260);
and U4555 (N_4555,N_4191,N_4362);
and U4556 (N_4556,N_4229,N_4304);
or U4557 (N_4557,N_4328,N_4084);
nor U4558 (N_4558,N_4038,N_4382);
nor U4559 (N_4559,N_4186,N_4395);
nand U4560 (N_4560,N_4400,N_4122);
nor U4561 (N_4561,N_4050,N_4223);
nand U4562 (N_4562,N_4426,N_4266);
or U4563 (N_4563,N_4318,N_4067);
nand U4564 (N_4564,N_4119,N_4120);
or U4565 (N_4565,N_4446,N_4212);
nand U4566 (N_4566,N_4387,N_4348);
nand U4567 (N_4567,N_4383,N_4315);
xor U4568 (N_4568,N_4358,N_4449);
nor U4569 (N_4569,N_4241,N_4291);
and U4570 (N_4570,N_4083,N_4238);
nand U4571 (N_4571,N_4408,N_4335);
xnor U4572 (N_4572,N_4424,N_4284);
or U4573 (N_4573,N_4299,N_4368);
or U4574 (N_4574,N_4316,N_4339);
nand U4575 (N_4575,N_4152,N_4372);
and U4576 (N_4576,N_4171,N_4354);
xor U4577 (N_4577,N_4162,N_4042);
or U4578 (N_4578,N_4235,N_4179);
nand U4579 (N_4579,N_4345,N_4076);
xor U4580 (N_4580,N_4350,N_4135);
nor U4581 (N_4581,N_4330,N_4411);
xnor U4582 (N_4582,N_4234,N_4405);
nor U4583 (N_4583,N_4381,N_4275);
and U4584 (N_4584,N_4010,N_4340);
and U4585 (N_4585,N_4211,N_4161);
and U4586 (N_4586,N_4361,N_4197);
or U4587 (N_4587,N_4336,N_4087);
nor U4588 (N_4588,N_4429,N_4226);
nand U4589 (N_4589,N_4068,N_4002);
nor U4590 (N_4590,N_4454,N_4462);
nor U4591 (N_4591,N_4170,N_4305);
nand U4592 (N_4592,N_4293,N_4174);
xor U4593 (N_4593,N_4425,N_4443);
or U4594 (N_4594,N_4290,N_4440);
nor U4595 (N_4595,N_4427,N_4380);
nor U4596 (N_4596,N_4111,N_4205);
nand U4597 (N_4597,N_4251,N_4003);
or U4598 (N_4598,N_4208,N_4396);
and U4599 (N_4599,N_4355,N_4088);
nand U4600 (N_4600,N_4190,N_4160);
nand U4601 (N_4601,N_4257,N_4113);
and U4602 (N_4602,N_4185,N_4453);
or U4603 (N_4603,N_4320,N_4065);
nor U4604 (N_4604,N_4329,N_4237);
and U4605 (N_4605,N_4421,N_4231);
nor U4606 (N_4606,N_4202,N_4032);
or U4607 (N_4607,N_4109,N_4327);
and U4608 (N_4608,N_4142,N_4035);
and U4609 (N_4609,N_4163,N_4016);
or U4610 (N_4610,N_4064,N_4412);
nand U4611 (N_4611,N_4196,N_4464);
and U4612 (N_4612,N_4494,N_4386);
or U4613 (N_4613,N_4459,N_4341);
and U4614 (N_4614,N_4136,N_4233);
xnor U4615 (N_4615,N_4027,N_4436);
nor U4616 (N_4616,N_4061,N_4147);
and U4617 (N_4617,N_4378,N_4046);
nand U4618 (N_4618,N_4447,N_4129);
nand U4619 (N_4619,N_4303,N_4297);
nand U4620 (N_4620,N_4128,N_4183);
or U4621 (N_4621,N_4021,N_4401);
xnor U4622 (N_4622,N_4334,N_4302);
or U4623 (N_4623,N_4474,N_4256);
and U4624 (N_4624,N_4495,N_4086);
nor U4625 (N_4625,N_4269,N_4013);
and U4626 (N_4626,N_4370,N_4018);
or U4627 (N_4627,N_4228,N_4071);
and U4628 (N_4628,N_4056,N_4081);
nand U4629 (N_4629,N_4364,N_4254);
nand U4630 (N_4630,N_4244,N_4014);
and U4631 (N_4631,N_4463,N_4192);
and U4632 (N_4632,N_4419,N_4338);
and U4633 (N_4633,N_4486,N_4103);
and U4634 (N_4634,N_4417,N_4100);
and U4635 (N_4635,N_4031,N_4222);
nand U4636 (N_4636,N_4154,N_4204);
or U4637 (N_4637,N_4052,N_4029);
or U4638 (N_4638,N_4379,N_4442);
nor U4639 (N_4639,N_4434,N_4295);
or U4640 (N_4640,N_4047,N_4249);
nand U4641 (N_4641,N_4110,N_4282);
nand U4642 (N_4642,N_4470,N_4265);
nor U4643 (N_4643,N_4272,N_4248);
or U4644 (N_4644,N_4130,N_4481);
and U4645 (N_4645,N_4094,N_4393);
and U4646 (N_4646,N_4273,N_4227);
or U4647 (N_4647,N_4398,N_4015);
nor U4648 (N_4648,N_4422,N_4267);
nor U4649 (N_4649,N_4456,N_4199);
xnor U4650 (N_4650,N_4433,N_4416);
and U4651 (N_4651,N_4468,N_4312);
and U4652 (N_4652,N_4264,N_4352);
xnor U4653 (N_4653,N_4274,N_4326);
nor U4654 (N_4654,N_4406,N_4452);
or U4655 (N_4655,N_4073,N_4085);
xor U4656 (N_4656,N_4132,N_4356);
nor U4657 (N_4657,N_4300,N_4278);
xor U4658 (N_4658,N_4466,N_4156);
or U4659 (N_4659,N_4098,N_4004);
or U4660 (N_4660,N_4365,N_4024);
and U4661 (N_4661,N_4178,N_4490);
and U4662 (N_4662,N_4180,N_4479);
and U4663 (N_4663,N_4394,N_4498);
and U4664 (N_4664,N_4005,N_4009);
nand U4665 (N_4665,N_4346,N_4023);
or U4666 (N_4666,N_4025,N_4261);
or U4667 (N_4667,N_4491,N_4359);
nand U4668 (N_4668,N_4332,N_4322);
and U4669 (N_4669,N_4078,N_4062);
or U4670 (N_4670,N_4165,N_4169);
xor U4671 (N_4671,N_4319,N_4072);
nor U4672 (N_4672,N_4090,N_4438);
nand U4673 (N_4673,N_4203,N_4317);
nor U4674 (N_4674,N_4457,N_4323);
or U4675 (N_4675,N_4377,N_4477);
xnor U4676 (N_4676,N_4376,N_4054);
and U4677 (N_4677,N_4177,N_4418);
and U4678 (N_4678,N_4189,N_4011);
and U4679 (N_4679,N_4195,N_4176);
and U4680 (N_4680,N_4285,N_4181);
or U4681 (N_4681,N_4252,N_4287);
nand U4682 (N_4682,N_4258,N_4187);
nor U4683 (N_4683,N_4342,N_4240);
nand U4684 (N_4684,N_4333,N_4201);
and U4685 (N_4685,N_4216,N_4172);
nor U4686 (N_4686,N_4059,N_4091);
or U4687 (N_4687,N_4392,N_4351);
and U4688 (N_4688,N_4198,N_4409);
or U4689 (N_4689,N_4385,N_4283);
or U4690 (N_4690,N_4388,N_4155);
or U4691 (N_4691,N_4445,N_4455);
and U4692 (N_4692,N_4074,N_4022);
nand U4693 (N_4693,N_4168,N_4106);
or U4694 (N_4694,N_4281,N_4141);
and U4695 (N_4695,N_4347,N_4402);
xnor U4696 (N_4696,N_4117,N_4026);
nor U4697 (N_4697,N_4093,N_4230);
nand U4698 (N_4698,N_4209,N_4096);
nand U4699 (N_4699,N_4397,N_4471);
nand U4700 (N_4700,N_4118,N_4289);
nand U4701 (N_4701,N_4137,N_4247);
xnor U4702 (N_4702,N_4337,N_4045);
and U4703 (N_4703,N_4263,N_4207);
nand U4704 (N_4704,N_4140,N_4159);
and U4705 (N_4705,N_4164,N_4373);
nor U4706 (N_4706,N_4063,N_4127);
nand U4707 (N_4707,N_4055,N_4007);
nand U4708 (N_4708,N_4123,N_4262);
nor U4709 (N_4709,N_4080,N_4276);
nor U4710 (N_4710,N_4423,N_4473);
and U4711 (N_4711,N_4444,N_4485);
and U4712 (N_4712,N_4374,N_4448);
nor U4713 (N_4713,N_4048,N_4225);
nand U4714 (N_4714,N_4006,N_4060);
xnor U4715 (N_4715,N_4410,N_4391);
xor U4716 (N_4716,N_4250,N_4480);
or U4717 (N_4717,N_4075,N_4077);
or U4718 (N_4718,N_4363,N_4496);
nand U4719 (N_4719,N_4143,N_4188);
and U4720 (N_4720,N_4413,N_4057);
or U4721 (N_4721,N_4294,N_4343);
xnor U4722 (N_4722,N_4214,N_4144);
or U4723 (N_4723,N_4020,N_4124);
or U4724 (N_4724,N_4221,N_4497);
nor U4725 (N_4725,N_4460,N_4367);
xor U4726 (N_4726,N_4253,N_4499);
and U4727 (N_4727,N_4213,N_4182);
nand U4728 (N_4728,N_4467,N_4243);
and U4729 (N_4729,N_4487,N_4314);
nor U4730 (N_4730,N_4404,N_4469);
nor U4731 (N_4731,N_4066,N_4441);
nor U4732 (N_4732,N_4138,N_4437);
nand U4733 (N_4733,N_4158,N_4431);
or U4734 (N_4734,N_4420,N_4371);
nor U4735 (N_4735,N_4450,N_4217);
or U4736 (N_4736,N_4131,N_4313);
nor U4737 (N_4737,N_4114,N_4104);
or U4738 (N_4738,N_4125,N_4301);
and U4739 (N_4739,N_4270,N_4175);
nor U4740 (N_4740,N_4194,N_4215);
nand U4741 (N_4741,N_4489,N_4149);
nand U4742 (N_4742,N_4414,N_4306);
or U4743 (N_4743,N_4017,N_4435);
nor U4744 (N_4744,N_4145,N_4097);
or U4745 (N_4745,N_4115,N_4415);
nor U4746 (N_4746,N_4280,N_4403);
or U4747 (N_4747,N_4089,N_4375);
nor U4748 (N_4748,N_4166,N_4279);
nor U4749 (N_4749,N_4296,N_4126);
nor U4750 (N_4750,N_4001,N_4164);
xnor U4751 (N_4751,N_4377,N_4479);
or U4752 (N_4752,N_4460,N_4156);
or U4753 (N_4753,N_4444,N_4024);
nor U4754 (N_4754,N_4152,N_4112);
xor U4755 (N_4755,N_4155,N_4497);
nand U4756 (N_4756,N_4259,N_4169);
and U4757 (N_4757,N_4046,N_4147);
nand U4758 (N_4758,N_4332,N_4449);
nand U4759 (N_4759,N_4113,N_4058);
nand U4760 (N_4760,N_4471,N_4032);
or U4761 (N_4761,N_4429,N_4278);
nand U4762 (N_4762,N_4328,N_4038);
and U4763 (N_4763,N_4185,N_4372);
nor U4764 (N_4764,N_4188,N_4437);
nand U4765 (N_4765,N_4237,N_4228);
and U4766 (N_4766,N_4435,N_4271);
nor U4767 (N_4767,N_4182,N_4456);
xor U4768 (N_4768,N_4157,N_4136);
xnor U4769 (N_4769,N_4113,N_4466);
and U4770 (N_4770,N_4422,N_4226);
nand U4771 (N_4771,N_4348,N_4407);
nand U4772 (N_4772,N_4173,N_4296);
nand U4773 (N_4773,N_4381,N_4451);
or U4774 (N_4774,N_4010,N_4286);
xor U4775 (N_4775,N_4415,N_4105);
or U4776 (N_4776,N_4414,N_4208);
or U4777 (N_4777,N_4389,N_4469);
nor U4778 (N_4778,N_4092,N_4286);
nor U4779 (N_4779,N_4170,N_4440);
or U4780 (N_4780,N_4129,N_4491);
nand U4781 (N_4781,N_4448,N_4331);
or U4782 (N_4782,N_4314,N_4163);
nand U4783 (N_4783,N_4123,N_4120);
or U4784 (N_4784,N_4319,N_4099);
or U4785 (N_4785,N_4140,N_4414);
or U4786 (N_4786,N_4454,N_4203);
xor U4787 (N_4787,N_4063,N_4044);
nor U4788 (N_4788,N_4000,N_4194);
nor U4789 (N_4789,N_4358,N_4315);
xor U4790 (N_4790,N_4319,N_4287);
or U4791 (N_4791,N_4253,N_4195);
nand U4792 (N_4792,N_4300,N_4044);
nor U4793 (N_4793,N_4425,N_4315);
and U4794 (N_4794,N_4250,N_4131);
or U4795 (N_4795,N_4023,N_4265);
and U4796 (N_4796,N_4493,N_4158);
or U4797 (N_4797,N_4496,N_4488);
nor U4798 (N_4798,N_4092,N_4065);
and U4799 (N_4799,N_4237,N_4498);
or U4800 (N_4800,N_4124,N_4476);
nor U4801 (N_4801,N_4460,N_4167);
nor U4802 (N_4802,N_4131,N_4497);
nor U4803 (N_4803,N_4359,N_4394);
and U4804 (N_4804,N_4154,N_4304);
and U4805 (N_4805,N_4078,N_4463);
nor U4806 (N_4806,N_4403,N_4211);
and U4807 (N_4807,N_4196,N_4390);
and U4808 (N_4808,N_4002,N_4118);
nand U4809 (N_4809,N_4398,N_4349);
and U4810 (N_4810,N_4016,N_4153);
or U4811 (N_4811,N_4483,N_4190);
nor U4812 (N_4812,N_4454,N_4464);
nand U4813 (N_4813,N_4036,N_4000);
xor U4814 (N_4814,N_4043,N_4190);
and U4815 (N_4815,N_4391,N_4423);
nand U4816 (N_4816,N_4360,N_4459);
or U4817 (N_4817,N_4142,N_4456);
xnor U4818 (N_4818,N_4289,N_4263);
nand U4819 (N_4819,N_4054,N_4249);
nor U4820 (N_4820,N_4027,N_4169);
xnor U4821 (N_4821,N_4467,N_4297);
nand U4822 (N_4822,N_4183,N_4013);
nor U4823 (N_4823,N_4495,N_4144);
and U4824 (N_4824,N_4452,N_4475);
or U4825 (N_4825,N_4136,N_4016);
nand U4826 (N_4826,N_4291,N_4367);
or U4827 (N_4827,N_4432,N_4165);
nand U4828 (N_4828,N_4375,N_4285);
nor U4829 (N_4829,N_4184,N_4041);
nand U4830 (N_4830,N_4261,N_4140);
nor U4831 (N_4831,N_4136,N_4452);
or U4832 (N_4832,N_4020,N_4344);
nand U4833 (N_4833,N_4369,N_4180);
and U4834 (N_4834,N_4112,N_4244);
and U4835 (N_4835,N_4174,N_4314);
nand U4836 (N_4836,N_4364,N_4419);
xnor U4837 (N_4837,N_4124,N_4042);
nand U4838 (N_4838,N_4087,N_4228);
or U4839 (N_4839,N_4036,N_4025);
nor U4840 (N_4840,N_4081,N_4115);
xor U4841 (N_4841,N_4046,N_4161);
nor U4842 (N_4842,N_4259,N_4493);
nor U4843 (N_4843,N_4459,N_4488);
nor U4844 (N_4844,N_4307,N_4393);
xnor U4845 (N_4845,N_4273,N_4447);
nand U4846 (N_4846,N_4328,N_4217);
and U4847 (N_4847,N_4069,N_4272);
or U4848 (N_4848,N_4098,N_4426);
and U4849 (N_4849,N_4403,N_4357);
or U4850 (N_4850,N_4406,N_4432);
nor U4851 (N_4851,N_4429,N_4045);
nand U4852 (N_4852,N_4244,N_4392);
nor U4853 (N_4853,N_4396,N_4493);
xor U4854 (N_4854,N_4045,N_4499);
nor U4855 (N_4855,N_4070,N_4041);
nor U4856 (N_4856,N_4485,N_4351);
or U4857 (N_4857,N_4240,N_4092);
and U4858 (N_4858,N_4160,N_4115);
or U4859 (N_4859,N_4400,N_4111);
nand U4860 (N_4860,N_4276,N_4018);
nand U4861 (N_4861,N_4279,N_4028);
nand U4862 (N_4862,N_4346,N_4012);
or U4863 (N_4863,N_4090,N_4263);
or U4864 (N_4864,N_4205,N_4187);
nor U4865 (N_4865,N_4223,N_4251);
nor U4866 (N_4866,N_4199,N_4396);
nor U4867 (N_4867,N_4368,N_4013);
xnor U4868 (N_4868,N_4042,N_4402);
nand U4869 (N_4869,N_4378,N_4481);
nor U4870 (N_4870,N_4239,N_4245);
and U4871 (N_4871,N_4012,N_4370);
or U4872 (N_4872,N_4318,N_4469);
or U4873 (N_4873,N_4108,N_4448);
nor U4874 (N_4874,N_4080,N_4252);
and U4875 (N_4875,N_4229,N_4082);
nor U4876 (N_4876,N_4337,N_4173);
or U4877 (N_4877,N_4484,N_4276);
and U4878 (N_4878,N_4040,N_4278);
nor U4879 (N_4879,N_4021,N_4151);
xor U4880 (N_4880,N_4129,N_4157);
or U4881 (N_4881,N_4265,N_4045);
nand U4882 (N_4882,N_4170,N_4064);
nand U4883 (N_4883,N_4164,N_4044);
and U4884 (N_4884,N_4078,N_4343);
nor U4885 (N_4885,N_4487,N_4377);
nand U4886 (N_4886,N_4288,N_4266);
nor U4887 (N_4887,N_4494,N_4066);
or U4888 (N_4888,N_4362,N_4033);
nand U4889 (N_4889,N_4421,N_4483);
nand U4890 (N_4890,N_4253,N_4413);
xor U4891 (N_4891,N_4424,N_4342);
and U4892 (N_4892,N_4368,N_4057);
and U4893 (N_4893,N_4430,N_4153);
nor U4894 (N_4894,N_4052,N_4207);
nand U4895 (N_4895,N_4373,N_4386);
nand U4896 (N_4896,N_4303,N_4438);
or U4897 (N_4897,N_4297,N_4393);
or U4898 (N_4898,N_4209,N_4437);
xor U4899 (N_4899,N_4407,N_4271);
nor U4900 (N_4900,N_4174,N_4035);
or U4901 (N_4901,N_4476,N_4060);
xor U4902 (N_4902,N_4187,N_4058);
nand U4903 (N_4903,N_4363,N_4462);
or U4904 (N_4904,N_4375,N_4153);
nand U4905 (N_4905,N_4447,N_4019);
nor U4906 (N_4906,N_4169,N_4124);
and U4907 (N_4907,N_4003,N_4173);
xnor U4908 (N_4908,N_4352,N_4080);
xnor U4909 (N_4909,N_4102,N_4470);
nand U4910 (N_4910,N_4381,N_4312);
or U4911 (N_4911,N_4303,N_4344);
nand U4912 (N_4912,N_4374,N_4052);
or U4913 (N_4913,N_4092,N_4409);
nand U4914 (N_4914,N_4435,N_4413);
nand U4915 (N_4915,N_4307,N_4166);
nand U4916 (N_4916,N_4065,N_4442);
xnor U4917 (N_4917,N_4030,N_4272);
or U4918 (N_4918,N_4433,N_4033);
and U4919 (N_4919,N_4244,N_4166);
nor U4920 (N_4920,N_4328,N_4437);
nor U4921 (N_4921,N_4122,N_4071);
nand U4922 (N_4922,N_4317,N_4117);
or U4923 (N_4923,N_4368,N_4158);
or U4924 (N_4924,N_4263,N_4229);
or U4925 (N_4925,N_4052,N_4421);
and U4926 (N_4926,N_4238,N_4362);
nor U4927 (N_4927,N_4209,N_4491);
nand U4928 (N_4928,N_4399,N_4201);
nor U4929 (N_4929,N_4080,N_4363);
nor U4930 (N_4930,N_4364,N_4472);
and U4931 (N_4931,N_4400,N_4151);
and U4932 (N_4932,N_4326,N_4437);
or U4933 (N_4933,N_4361,N_4268);
nor U4934 (N_4934,N_4292,N_4278);
and U4935 (N_4935,N_4212,N_4341);
xnor U4936 (N_4936,N_4285,N_4113);
nor U4937 (N_4937,N_4114,N_4227);
xnor U4938 (N_4938,N_4237,N_4213);
or U4939 (N_4939,N_4032,N_4276);
or U4940 (N_4940,N_4326,N_4399);
nand U4941 (N_4941,N_4337,N_4225);
or U4942 (N_4942,N_4106,N_4493);
or U4943 (N_4943,N_4260,N_4003);
and U4944 (N_4944,N_4081,N_4387);
nand U4945 (N_4945,N_4165,N_4223);
nand U4946 (N_4946,N_4492,N_4108);
and U4947 (N_4947,N_4244,N_4431);
nand U4948 (N_4948,N_4414,N_4479);
and U4949 (N_4949,N_4277,N_4193);
nor U4950 (N_4950,N_4260,N_4435);
or U4951 (N_4951,N_4006,N_4352);
nor U4952 (N_4952,N_4182,N_4324);
xor U4953 (N_4953,N_4482,N_4411);
nand U4954 (N_4954,N_4067,N_4008);
xnor U4955 (N_4955,N_4352,N_4200);
or U4956 (N_4956,N_4127,N_4001);
and U4957 (N_4957,N_4332,N_4425);
xnor U4958 (N_4958,N_4286,N_4177);
nand U4959 (N_4959,N_4482,N_4436);
nand U4960 (N_4960,N_4461,N_4189);
nand U4961 (N_4961,N_4026,N_4194);
nand U4962 (N_4962,N_4303,N_4366);
nand U4963 (N_4963,N_4245,N_4388);
or U4964 (N_4964,N_4079,N_4262);
and U4965 (N_4965,N_4346,N_4303);
xnor U4966 (N_4966,N_4123,N_4035);
or U4967 (N_4967,N_4308,N_4064);
nor U4968 (N_4968,N_4026,N_4079);
or U4969 (N_4969,N_4236,N_4175);
nand U4970 (N_4970,N_4133,N_4080);
and U4971 (N_4971,N_4069,N_4200);
nor U4972 (N_4972,N_4242,N_4421);
nand U4973 (N_4973,N_4116,N_4329);
and U4974 (N_4974,N_4367,N_4349);
and U4975 (N_4975,N_4140,N_4195);
and U4976 (N_4976,N_4283,N_4414);
and U4977 (N_4977,N_4248,N_4456);
and U4978 (N_4978,N_4408,N_4216);
and U4979 (N_4979,N_4426,N_4143);
and U4980 (N_4980,N_4112,N_4088);
nor U4981 (N_4981,N_4017,N_4226);
or U4982 (N_4982,N_4361,N_4055);
nor U4983 (N_4983,N_4269,N_4063);
and U4984 (N_4984,N_4105,N_4405);
nand U4985 (N_4985,N_4154,N_4426);
and U4986 (N_4986,N_4183,N_4035);
nand U4987 (N_4987,N_4050,N_4359);
or U4988 (N_4988,N_4211,N_4456);
nand U4989 (N_4989,N_4464,N_4315);
nand U4990 (N_4990,N_4191,N_4478);
and U4991 (N_4991,N_4031,N_4399);
nand U4992 (N_4992,N_4360,N_4167);
and U4993 (N_4993,N_4425,N_4405);
nor U4994 (N_4994,N_4471,N_4475);
nand U4995 (N_4995,N_4427,N_4016);
nor U4996 (N_4996,N_4434,N_4082);
nand U4997 (N_4997,N_4000,N_4235);
nor U4998 (N_4998,N_4342,N_4218);
nor U4999 (N_4999,N_4254,N_4371);
xor U5000 (N_5000,N_4766,N_4572);
and U5001 (N_5001,N_4935,N_4652);
and U5002 (N_5002,N_4557,N_4970);
and U5003 (N_5003,N_4612,N_4747);
nor U5004 (N_5004,N_4639,N_4955);
nor U5005 (N_5005,N_4633,N_4725);
nand U5006 (N_5006,N_4928,N_4762);
or U5007 (N_5007,N_4655,N_4579);
nor U5008 (N_5008,N_4829,N_4558);
or U5009 (N_5009,N_4591,N_4830);
and U5010 (N_5010,N_4565,N_4711);
nor U5011 (N_5011,N_4776,N_4798);
or U5012 (N_5012,N_4919,N_4653);
xnor U5013 (N_5013,N_4743,N_4512);
nor U5014 (N_5014,N_4780,N_4944);
or U5015 (N_5015,N_4657,N_4936);
nand U5016 (N_5016,N_4744,N_4772);
or U5017 (N_5017,N_4905,N_4932);
or U5018 (N_5018,N_4745,N_4629);
or U5019 (N_5019,N_4883,N_4575);
nor U5020 (N_5020,N_4841,N_4686);
and U5021 (N_5021,N_4576,N_4690);
and U5022 (N_5022,N_4817,N_4615);
or U5023 (N_5023,N_4736,N_4902);
or U5024 (N_5024,N_4953,N_4869);
nand U5025 (N_5025,N_4625,N_4685);
and U5026 (N_5026,N_4804,N_4771);
or U5027 (N_5027,N_4834,N_4982);
nand U5028 (N_5028,N_4832,N_4887);
nand U5029 (N_5029,N_4989,N_4680);
and U5030 (N_5030,N_4994,N_4667);
and U5031 (N_5031,N_4514,N_4937);
nor U5032 (N_5032,N_4526,N_4527);
nand U5033 (N_5033,N_4952,N_4805);
and U5034 (N_5034,N_4785,N_4818);
or U5035 (N_5035,N_4654,N_4590);
or U5036 (N_5036,N_4899,N_4700);
nand U5037 (N_5037,N_4783,N_4607);
or U5038 (N_5038,N_4751,N_4746);
nor U5039 (N_5039,N_4675,N_4906);
or U5040 (N_5040,N_4934,N_4896);
nor U5041 (N_5041,N_4537,N_4687);
nor U5042 (N_5042,N_4695,N_4858);
and U5043 (N_5043,N_4597,N_4987);
nand U5044 (N_5044,N_4541,N_4813);
and U5045 (N_5045,N_4609,N_4912);
xnor U5046 (N_5046,N_4561,N_4578);
nand U5047 (N_5047,N_4918,N_4648);
or U5048 (N_5048,N_4574,N_4660);
nand U5049 (N_5049,N_4681,N_4656);
nor U5050 (N_5050,N_4956,N_4958);
xor U5051 (N_5051,N_4636,N_4594);
or U5052 (N_5052,N_4559,N_4645);
nor U5053 (N_5053,N_4671,N_4567);
or U5054 (N_5054,N_4616,N_4981);
or U5055 (N_5055,N_4506,N_4548);
nor U5056 (N_5056,N_4821,N_4861);
and U5057 (N_5057,N_4820,N_4778);
nand U5058 (N_5058,N_4809,N_4904);
nand U5059 (N_5059,N_4727,N_4707);
xor U5060 (N_5060,N_4968,N_4709);
nor U5061 (N_5061,N_4518,N_4717);
or U5062 (N_5062,N_4848,N_4699);
or U5063 (N_5063,N_4500,N_4913);
nor U5064 (N_5064,N_4917,N_4768);
nand U5065 (N_5065,N_4596,N_4697);
or U5066 (N_5066,N_4826,N_4640);
xor U5067 (N_5067,N_4856,N_4847);
and U5068 (N_5068,N_4642,N_4553);
nor U5069 (N_5069,N_4706,N_4903);
or U5070 (N_5070,N_4765,N_4679);
xor U5071 (N_5071,N_4692,N_4758);
and U5072 (N_5072,N_4501,N_4670);
or U5073 (N_5073,N_4814,N_4610);
and U5074 (N_5074,N_4613,N_4611);
nor U5075 (N_5075,N_4986,N_4603);
xnor U5076 (N_5076,N_4513,N_4757);
and U5077 (N_5077,N_4539,N_4517);
xor U5078 (N_5078,N_4938,N_4849);
nand U5079 (N_5079,N_4571,N_4885);
nor U5080 (N_5080,N_4593,N_4538);
and U5081 (N_5081,N_4983,N_4773);
or U5082 (N_5082,N_4601,N_4605);
nor U5083 (N_5083,N_4948,N_4698);
or U5084 (N_5084,N_4712,N_4844);
or U5085 (N_5085,N_4504,N_4967);
or U5086 (N_5086,N_4910,N_4569);
xnor U5087 (N_5087,N_4632,N_4560);
nor U5088 (N_5088,N_4728,N_4840);
xnor U5089 (N_5089,N_4855,N_4516);
and U5090 (N_5090,N_4879,N_4713);
nand U5091 (N_5091,N_4545,N_4749);
xor U5092 (N_5092,N_4801,N_4876);
xnor U5093 (N_5093,N_4731,N_4810);
or U5094 (N_5094,N_4886,N_4942);
xor U5095 (N_5095,N_4995,N_4877);
nor U5096 (N_5096,N_4833,N_4760);
nand U5097 (N_5097,N_4803,N_4750);
xor U5098 (N_5098,N_4650,N_4864);
xnor U5099 (N_5099,N_4975,N_4533);
or U5100 (N_5100,N_4872,N_4583);
and U5101 (N_5101,N_4852,N_4641);
nor U5102 (N_5102,N_4977,N_4889);
or U5103 (N_5103,N_4602,N_4900);
nor U5104 (N_5104,N_4867,N_4664);
nand U5105 (N_5105,N_4822,N_4988);
nand U5106 (N_5106,N_4523,N_4782);
nand U5107 (N_5107,N_4812,N_4756);
or U5108 (N_5108,N_4888,N_4684);
nand U5109 (N_5109,N_4550,N_4863);
nor U5110 (N_5110,N_4542,N_4505);
and U5111 (N_5111,N_4920,N_4960);
or U5112 (N_5112,N_4658,N_4819);
or U5113 (N_5113,N_4815,N_4828);
nand U5114 (N_5114,N_4528,N_4845);
or U5115 (N_5115,N_4666,N_4647);
and U5116 (N_5116,N_4683,N_4722);
xor U5117 (N_5117,N_4614,N_4908);
and U5118 (N_5118,N_4577,N_4769);
xor U5119 (N_5119,N_4965,N_4914);
and U5120 (N_5120,N_4898,N_4892);
or U5121 (N_5121,N_4691,N_4622);
xnor U5122 (N_5122,N_4868,N_4978);
nand U5123 (N_5123,N_4519,N_4677);
nand U5124 (N_5124,N_4825,N_4595);
or U5125 (N_5125,N_4882,N_4857);
and U5126 (N_5126,N_4945,N_4588);
or U5127 (N_5127,N_4922,N_4573);
nand U5128 (N_5128,N_4973,N_4663);
and U5129 (N_5129,N_4881,N_4676);
and U5130 (N_5130,N_4678,N_4570);
nor U5131 (N_5131,N_4532,N_4503);
nand U5132 (N_5132,N_4529,N_4703);
nor U5133 (N_5133,N_4754,N_4544);
nand U5134 (N_5134,N_4959,N_4586);
nand U5135 (N_5135,N_4950,N_4617);
nand U5136 (N_5136,N_4954,N_4907);
nand U5137 (N_5137,N_4726,N_4742);
and U5138 (N_5138,N_4897,N_4630);
xnor U5139 (N_5139,N_4556,N_4789);
and U5140 (N_5140,N_4669,N_4871);
xor U5141 (N_5141,N_4774,N_4974);
nand U5142 (N_5142,N_4748,N_4551);
nor U5143 (N_5143,N_4720,N_4962);
nor U5144 (N_5144,N_4716,N_4502);
or U5145 (N_5145,N_4816,N_4635);
nor U5146 (N_5146,N_4637,N_4659);
nor U5147 (N_5147,N_4719,N_4600);
nor U5148 (N_5148,N_4730,N_4587);
nand U5149 (N_5149,N_4668,N_4795);
nor U5150 (N_5150,N_4797,N_4939);
nand U5151 (N_5151,N_4672,N_4651);
nand U5152 (N_5152,N_4592,N_4930);
or U5153 (N_5153,N_4710,N_4835);
nand U5154 (N_5154,N_4643,N_4862);
or U5155 (N_5155,N_4916,N_4721);
xnor U5156 (N_5156,N_4991,N_4850);
nor U5157 (N_5157,N_4608,N_4555);
or U5158 (N_5158,N_4619,N_4638);
and U5159 (N_5159,N_4554,N_4624);
and U5160 (N_5160,N_4693,N_4997);
nor U5161 (N_5161,N_4839,N_4623);
xnor U5162 (N_5162,N_4599,N_4521);
or U5163 (N_5163,N_4915,N_4701);
xnor U5164 (N_5164,N_4562,N_4507);
xnor U5165 (N_5165,N_4784,N_4927);
nor U5166 (N_5166,N_4674,N_4740);
and U5167 (N_5167,N_4568,N_4984);
nor U5168 (N_5168,N_4999,N_4971);
and U5169 (N_5169,N_4598,N_4787);
nor U5170 (N_5170,N_4705,N_4843);
and U5171 (N_5171,N_4921,N_4866);
xnor U5172 (N_5172,N_4741,N_4729);
and U5173 (N_5173,N_4792,N_4794);
nand U5174 (N_5174,N_4520,N_4961);
and U5175 (N_5175,N_4715,N_4799);
and U5176 (N_5176,N_4564,N_4646);
nor U5177 (N_5177,N_4626,N_4972);
and U5178 (N_5178,N_4547,N_4884);
nand U5179 (N_5179,N_4708,N_4851);
nand U5180 (N_5180,N_4890,N_4793);
and U5181 (N_5181,N_4604,N_4770);
nand U5182 (N_5182,N_4786,N_4585);
xnor U5183 (N_5183,N_4764,N_4511);
and U5184 (N_5184,N_4893,N_4752);
nand U5185 (N_5185,N_4563,N_4673);
nor U5186 (N_5186,N_4933,N_4925);
nor U5187 (N_5187,N_4949,N_4581);
and U5188 (N_5188,N_4723,N_4846);
and U5189 (N_5189,N_4923,N_4824);
nand U5190 (N_5190,N_4837,N_4880);
nor U5191 (N_5191,N_4662,N_4929);
nand U5192 (N_5192,N_4531,N_4582);
nor U5193 (N_5193,N_4943,N_4689);
nor U5194 (N_5194,N_4940,N_4842);
nand U5195 (N_5195,N_4536,N_4901);
and U5196 (N_5196,N_4985,N_4524);
xnor U5197 (N_5197,N_4508,N_4775);
nand U5198 (N_5198,N_4509,N_4791);
or U5199 (N_5199,N_4644,N_4796);
nor U5200 (N_5200,N_4990,N_4628);
nor U5201 (N_5201,N_4800,N_4618);
or U5202 (N_5202,N_4827,N_4781);
or U5203 (N_5203,N_4755,N_4714);
xor U5204 (N_5204,N_4580,N_4566);
xor U5205 (N_5205,N_4926,N_4552);
nand U5206 (N_5206,N_4621,N_4732);
or U5207 (N_5207,N_4525,N_4702);
and U5208 (N_5208,N_4788,N_4976);
xor U5209 (N_5209,N_4546,N_4946);
nand U5210 (N_5210,N_4996,N_4853);
and U5211 (N_5211,N_4535,N_4530);
and U5212 (N_5212,N_4957,N_4924);
nor U5213 (N_5213,N_4584,N_4688);
nand U5214 (N_5214,N_4836,N_4767);
or U5215 (N_5215,N_4859,N_4704);
nor U5216 (N_5216,N_4870,N_4759);
nor U5217 (N_5217,N_4875,N_4891);
and U5218 (N_5218,N_4947,N_4779);
nand U5219 (N_5219,N_4665,N_4854);
and U5220 (N_5220,N_4761,N_4865);
and U5221 (N_5221,N_4941,N_4510);
and U5222 (N_5222,N_4694,N_4606);
and U5223 (N_5223,N_4777,N_4738);
nand U5224 (N_5224,N_4620,N_4969);
xnor U5225 (N_5225,N_4993,N_4807);
and U5226 (N_5226,N_4831,N_4737);
and U5227 (N_5227,N_4763,N_4631);
or U5228 (N_5228,N_4790,N_4682);
or U5229 (N_5229,N_4838,N_4909);
and U5230 (N_5230,N_4649,N_4534);
nand U5231 (N_5231,N_4963,N_4931);
xnor U5232 (N_5232,N_4724,N_4998);
xnor U5233 (N_5233,N_4894,N_4734);
or U5234 (N_5234,N_4980,N_4718);
xnor U5235 (N_5235,N_4873,N_4860);
nor U5236 (N_5236,N_4589,N_4992);
and U5237 (N_5237,N_4733,N_4823);
or U5238 (N_5238,N_4802,N_4540);
xor U5239 (N_5239,N_4549,N_4661);
or U5240 (N_5240,N_4739,N_4811);
nor U5241 (N_5241,N_4878,N_4634);
and U5242 (N_5242,N_4874,N_4808);
xor U5243 (N_5243,N_4522,N_4911);
nand U5244 (N_5244,N_4951,N_4966);
xnor U5245 (N_5245,N_4515,N_4964);
nor U5246 (N_5246,N_4806,N_4895);
or U5247 (N_5247,N_4543,N_4979);
and U5248 (N_5248,N_4696,N_4627);
nor U5249 (N_5249,N_4753,N_4735);
nand U5250 (N_5250,N_4593,N_4782);
nor U5251 (N_5251,N_4909,N_4910);
nand U5252 (N_5252,N_4892,N_4968);
or U5253 (N_5253,N_4523,N_4987);
nand U5254 (N_5254,N_4583,N_4639);
nor U5255 (N_5255,N_4503,N_4743);
and U5256 (N_5256,N_4749,N_4677);
nand U5257 (N_5257,N_4871,N_4997);
nand U5258 (N_5258,N_4936,N_4829);
and U5259 (N_5259,N_4591,N_4501);
xnor U5260 (N_5260,N_4528,N_4539);
nor U5261 (N_5261,N_4891,N_4874);
and U5262 (N_5262,N_4565,N_4640);
nand U5263 (N_5263,N_4586,N_4696);
nand U5264 (N_5264,N_4778,N_4508);
nand U5265 (N_5265,N_4526,N_4899);
xor U5266 (N_5266,N_4811,N_4807);
and U5267 (N_5267,N_4539,N_4889);
nor U5268 (N_5268,N_4733,N_4809);
xnor U5269 (N_5269,N_4607,N_4525);
and U5270 (N_5270,N_4596,N_4963);
and U5271 (N_5271,N_4672,N_4851);
or U5272 (N_5272,N_4528,N_4619);
nor U5273 (N_5273,N_4796,N_4961);
xnor U5274 (N_5274,N_4879,N_4684);
or U5275 (N_5275,N_4944,N_4795);
nor U5276 (N_5276,N_4616,N_4980);
or U5277 (N_5277,N_4987,N_4815);
nand U5278 (N_5278,N_4685,N_4689);
nor U5279 (N_5279,N_4647,N_4535);
and U5280 (N_5280,N_4925,N_4707);
and U5281 (N_5281,N_4607,N_4808);
or U5282 (N_5282,N_4621,N_4598);
nor U5283 (N_5283,N_4668,N_4694);
nor U5284 (N_5284,N_4652,N_4818);
or U5285 (N_5285,N_4633,N_4710);
nor U5286 (N_5286,N_4701,N_4644);
xnor U5287 (N_5287,N_4739,N_4954);
and U5288 (N_5288,N_4513,N_4916);
or U5289 (N_5289,N_4806,N_4740);
xnor U5290 (N_5290,N_4674,N_4963);
nand U5291 (N_5291,N_4937,N_4651);
or U5292 (N_5292,N_4759,N_4930);
or U5293 (N_5293,N_4570,N_4973);
and U5294 (N_5294,N_4645,N_4877);
xnor U5295 (N_5295,N_4989,N_4818);
and U5296 (N_5296,N_4657,N_4762);
nor U5297 (N_5297,N_4683,N_4758);
nand U5298 (N_5298,N_4603,N_4513);
and U5299 (N_5299,N_4877,N_4564);
nand U5300 (N_5300,N_4558,N_4676);
xor U5301 (N_5301,N_4776,N_4702);
and U5302 (N_5302,N_4581,N_4730);
or U5303 (N_5303,N_4717,N_4570);
and U5304 (N_5304,N_4670,N_4611);
or U5305 (N_5305,N_4994,N_4637);
or U5306 (N_5306,N_4893,N_4544);
xnor U5307 (N_5307,N_4622,N_4595);
xnor U5308 (N_5308,N_4551,N_4635);
nand U5309 (N_5309,N_4567,N_4556);
and U5310 (N_5310,N_4815,N_4565);
nor U5311 (N_5311,N_4537,N_4971);
and U5312 (N_5312,N_4901,N_4820);
or U5313 (N_5313,N_4689,N_4533);
xnor U5314 (N_5314,N_4528,N_4834);
and U5315 (N_5315,N_4849,N_4633);
and U5316 (N_5316,N_4924,N_4560);
nor U5317 (N_5317,N_4845,N_4573);
or U5318 (N_5318,N_4507,N_4914);
xor U5319 (N_5319,N_4700,N_4575);
nand U5320 (N_5320,N_4682,N_4816);
or U5321 (N_5321,N_4648,N_4718);
and U5322 (N_5322,N_4779,N_4653);
and U5323 (N_5323,N_4777,N_4901);
nor U5324 (N_5324,N_4554,N_4613);
or U5325 (N_5325,N_4978,N_4701);
nand U5326 (N_5326,N_4519,N_4567);
nand U5327 (N_5327,N_4668,N_4622);
or U5328 (N_5328,N_4930,N_4879);
nor U5329 (N_5329,N_4736,N_4840);
and U5330 (N_5330,N_4703,N_4714);
nand U5331 (N_5331,N_4739,N_4884);
or U5332 (N_5332,N_4847,N_4797);
nor U5333 (N_5333,N_4936,N_4695);
or U5334 (N_5334,N_4603,N_4653);
or U5335 (N_5335,N_4748,N_4893);
nand U5336 (N_5336,N_4515,N_4987);
or U5337 (N_5337,N_4768,N_4968);
or U5338 (N_5338,N_4844,N_4513);
nand U5339 (N_5339,N_4625,N_4719);
nor U5340 (N_5340,N_4666,N_4609);
or U5341 (N_5341,N_4637,N_4849);
nor U5342 (N_5342,N_4640,N_4981);
nand U5343 (N_5343,N_4840,N_4772);
nor U5344 (N_5344,N_4746,N_4995);
or U5345 (N_5345,N_4869,N_4819);
nor U5346 (N_5346,N_4652,N_4618);
or U5347 (N_5347,N_4828,N_4693);
or U5348 (N_5348,N_4615,N_4856);
nand U5349 (N_5349,N_4518,N_4953);
or U5350 (N_5350,N_4801,N_4971);
and U5351 (N_5351,N_4690,N_4830);
and U5352 (N_5352,N_4653,N_4983);
and U5353 (N_5353,N_4934,N_4715);
xor U5354 (N_5354,N_4770,N_4734);
or U5355 (N_5355,N_4565,N_4841);
nor U5356 (N_5356,N_4684,N_4520);
and U5357 (N_5357,N_4573,N_4512);
nor U5358 (N_5358,N_4875,N_4583);
nand U5359 (N_5359,N_4813,N_4696);
nand U5360 (N_5360,N_4664,N_4842);
and U5361 (N_5361,N_4855,N_4864);
and U5362 (N_5362,N_4639,N_4997);
nand U5363 (N_5363,N_4902,N_4615);
nand U5364 (N_5364,N_4820,N_4556);
xor U5365 (N_5365,N_4866,N_4753);
and U5366 (N_5366,N_4659,N_4519);
and U5367 (N_5367,N_4580,N_4850);
and U5368 (N_5368,N_4807,N_4567);
nand U5369 (N_5369,N_4506,N_4789);
xor U5370 (N_5370,N_4921,N_4857);
nor U5371 (N_5371,N_4556,N_4962);
and U5372 (N_5372,N_4529,N_4515);
or U5373 (N_5373,N_4632,N_4958);
or U5374 (N_5374,N_4726,N_4858);
nor U5375 (N_5375,N_4991,N_4934);
or U5376 (N_5376,N_4970,N_4652);
or U5377 (N_5377,N_4830,N_4666);
nand U5378 (N_5378,N_4601,N_4871);
nand U5379 (N_5379,N_4603,N_4990);
nand U5380 (N_5380,N_4619,N_4860);
and U5381 (N_5381,N_4611,N_4870);
or U5382 (N_5382,N_4778,N_4849);
or U5383 (N_5383,N_4820,N_4942);
nor U5384 (N_5384,N_4916,N_4564);
or U5385 (N_5385,N_4776,N_4860);
nand U5386 (N_5386,N_4743,N_4638);
nor U5387 (N_5387,N_4916,N_4667);
nor U5388 (N_5388,N_4655,N_4582);
xnor U5389 (N_5389,N_4962,N_4517);
or U5390 (N_5390,N_4610,N_4584);
xor U5391 (N_5391,N_4741,N_4912);
or U5392 (N_5392,N_4568,N_4658);
and U5393 (N_5393,N_4922,N_4997);
nand U5394 (N_5394,N_4927,N_4749);
and U5395 (N_5395,N_4855,N_4948);
xor U5396 (N_5396,N_4740,N_4541);
nor U5397 (N_5397,N_4551,N_4962);
or U5398 (N_5398,N_4980,N_4590);
xnor U5399 (N_5399,N_4724,N_4788);
and U5400 (N_5400,N_4600,N_4686);
xnor U5401 (N_5401,N_4654,N_4762);
or U5402 (N_5402,N_4981,N_4779);
xor U5403 (N_5403,N_4965,N_4926);
nor U5404 (N_5404,N_4831,N_4568);
nand U5405 (N_5405,N_4883,N_4634);
or U5406 (N_5406,N_4973,N_4729);
or U5407 (N_5407,N_4870,N_4764);
xor U5408 (N_5408,N_4883,N_4980);
nor U5409 (N_5409,N_4972,N_4577);
nor U5410 (N_5410,N_4643,N_4675);
nor U5411 (N_5411,N_4981,N_4534);
xor U5412 (N_5412,N_4742,N_4707);
xor U5413 (N_5413,N_4830,N_4713);
nand U5414 (N_5414,N_4779,N_4927);
nand U5415 (N_5415,N_4874,N_4909);
nand U5416 (N_5416,N_4936,N_4862);
nand U5417 (N_5417,N_4674,N_4985);
and U5418 (N_5418,N_4603,N_4567);
nor U5419 (N_5419,N_4784,N_4698);
nor U5420 (N_5420,N_4720,N_4635);
and U5421 (N_5421,N_4808,N_4989);
and U5422 (N_5422,N_4765,N_4683);
nor U5423 (N_5423,N_4618,N_4858);
and U5424 (N_5424,N_4582,N_4715);
nand U5425 (N_5425,N_4698,N_4543);
or U5426 (N_5426,N_4954,N_4827);
and U5427 (N_5427,N_4884,N_4809);
nor U5428 (N_5428,N_4650,N_4819);
nor U5429 (N_5429,N_4590,N_4714);
or U5430 (N_5430,N_4604,N_4527);
nand U5431 (N_5431,N_4790,N_4551);
and U5432 (N_5432,N_4705,N_4711);
nand U5433 (N_5433,N_4526,N_4540);
and U5434 (N_5434,N_4607,N_4549);
nand U5435 (N_5435,N_4541,N_4872);
or U5436 (N_5436,N_4956,N_4618);
or U5437 (N_5437,N_4508,N_4717);
nand U5438 (N_5438,N_4762,N_4642);
nand U5439 (N_5439,N_4731,N_4803);
nand U5440 (N_5440,N_4577,N_4619);
or U5441 (N_5441,N_4850,N_4751);
nand U5442 (N_5442,N_4728,N_4903);
and U5443 (N_5443,N_4921,N_4878);
nor U5444 (N_5444,N_4613,N_4822);
or U5445 (N_5445,N_4734,N_4601);
or U5446 (N_5446,N_4840,N_4739);
and U5447 (N_5447,N_4685,N_4991);
nand U5448 (N_5448,N_4974,N_4987);
nand U5449 (N_5449,N_4776,N_4775);
nand U5450 (N_5450,N_4823,N_4738);
or U5451 (N_5451,N_4666,N_4654);
nor U5452 (N_5452,N_4900,N_4501);
nand U5453 (N_5453,N_4831,N_4767);
nand U5454 (N_5454,N_4689,N_4963);
or U5455 (N_5455,N_4969,N_4629);
and U5456 (N_5456,N_4901,N_4583);
nor U5457 (N_5457,N_4989,N_4835);
nor U5458 (N_5458,N_4547,N_4678);
and U5459 (N_5459,N_4661,N_4670);
and U5460 (N_5460,N_4794,N_4542);
nand U5461 (N_5461,N_4689,N_4698);
nand U5462 (N_5462,N_4567,N_4622);
nor U5463 (N_5463,N_4889,N_4592);
nand U5464 (N_5464,N_4558,N_4574);
nand U5465 (N_5465,N_4867,N_4801);
nand U5466 (N_5466,N_4540,N_4881);
nor U5467 (N_5467,N_4713,N_4508);
nand U5468 (N_5468,N_4619,N_4586);
nand U5469 (N_5469,N_4857,N_4781);
or U5470 (N_5470,N_4694,N_4644);
or U5471 (N_5471,N_4831,N_4595);
or U5472 (N_5472,N_4550,N_4755);
xnor U5473 (N_5473,N_4871,N_4756);
nor U5474 (N_5474,N_4934,N_4664);
nand U5475 (N_5475,N_4584,N_4958);
nand U5476 (N_5476,N_4912,N_4535);
or U5477 (N_5477,N_4677,N_4652);
and U5478 (N_5478,N_4947,N_4848);
and U5479 (N_5479,N_4773,N_4987);
nor U5480 (N_5480,N_4912,N_4873);
and U5481 (N_5481,N_4845,N_4974);
or U5482 (N_5482,N_4881,N_4904);
nor U5483 (N_5483,N_4926,N_4858);
and U5484 (N_5484,N_4705,N_4601);
nand U5485 (N_5485,N_4584,N_4779);
and U5486 (N_5486,N_4892,N_4716);
nand U5487 (N_5487,N_4516,N_4989);
and U5488 (N_5488,N_4581,N_4866);
and U5489 (N_5489,N_4857,N_4975);
nor U5490 (N_5490,N_4923,N_4664);
nor U5491 (N_5491,N_4947,N_4633);
nor U5492 (N_5492,N_4655,N_4772);
nand U5493 (N_5493,N_4602,N_4649);
and U5494 (N_5494,N_4510,N_4979);
or U5495 (N_5495,N_4748,N_4953);
or U5496 (N_5496,N_4694,N_4690);
and U5497 (N_5497,N_4617,N_4827);
and U5498 (N_5498,N_4516,N_4543);
and U5499 (N_5499,N_4840,N_4680);
nor U5500 (N_5500,N_5448,N_5463);
xnor U5501 (N_5501,N_5038,N_5324);
and U5502 (N_5502,N_5300,N_5176);
or U5503 (N_5503,N_5061,N_5320);
or U5504 (N_5504,N_5455,N_5318);
nor U5505 (N_5505,N_5170,N_5007);
nand U5506 (N_5506,N_5309,N_5494);
xor U5507 (N_5507,N_5456,N_5270);
or U5508 (N_5508,N_5296,N_5069);
nor U5509 (N_5509,N_5364,N_5288);
nor U5510 (N_5510,N_5251,N_5020);
or U5511 (N_5511,N_5354,N_5247);
or U5512 (N_5512,N_5478,N_5352);
and U5513 (N_5513,N_5183,N_5186);
nand U5514 (N_5514,N_5053,N_5276);
or U5515 (N_5515,N_5245,N_5321);
nor U5516 (N_5516,N_5190,N_5400);
and U5517 (N_5517,N_5198,N_5060);
nand U5518 (N_5518,N_5173,N_5477);
and U5519 (N_5519,N_5389,N_5015);
or U5520 (N_5520,N_5114,N_5254);
nand U5521 (N_5521,N_5362,N_5342);
or U5522 (N_5522,N_5047,N_5048);
and U5523 (N_5523,N_5044,N_5171);
nor U5524 (N_5524,N_5002,N_5475);
and U5525 (N_5525,N_5192,N_5027);
or U5526 (N_5526,N_5262,N_5116);
nand U5527 (N_5527,N_5095,N_5444);
nor U5528 (N_5528,N_5272,N_5135);
and U5529 (N_5529,N_5366,N_5465);
or U5530 (N_5530,N_5297,N_5267);
or U5531 (N_5531,N_5392,N_5074);
nor U5532 (N_5532,N_5115,N_5089);
nor U5533 (N_5533,N_5483,N_5129);
nor U5534 (N_5534,N_5386,N_5435);
nand U5535 (N_5535,N_5265,N_5070);
nand U5536 (N_5536,N_5417,N_5088);
xnor U5537 (N_5537,N_5480,N_5368);
or U5538 (N_5538,N_5004,N_5216);
nor U5539 (N_5539,N_5429,N_5406);
and U5540 (N_5540,N_5237,N_5040);
nand U5541 (N_5541,N_5033,N_5025);
nand U5542 (N_5542,N_5204,N_5239);
xnor U5543 (N_5543,N_5246,N_5343);
nor U5544 (N_5544,N_5458,N_5075);
and U5545 (N_5545,N_5000,N_5420);
or U5546 (N_5546,N_5079,N_5283);
and U5547 (N_5547,N_5419,N_5144);
nand U5548 (N_5548,N_5096,N_5016);
nand U5549 (N_5549,N_5290,N_5100);
nor U5550 (N_5550,N_5168,N_5197);
xnor U5551 (N_5551,N_5145,N_5303);
or U5552 (N_5552,N_5488,N_5059);
nor U5553 (N_5553,N_5055,N_5453);
nor U5554 (N_5554,N_5311,N_5306);
and U5555 (N_5555,N_5019,N_5414);
and U5556 (N_5556,N_5383,N_5146);
nor U5557 (N_5557,N_5489,N_5426);
nor U5558 (N_5558,N_5193,N_5063);
nand U5559 (N_5559,N_5139,N_5295);
xnor U5560 (N_5560,N_5211,N_5011);
nor U5561 (N_5561,N_5117,N_5031);
nor U5562 (N_5562,N_5138,N_5166);
or U5563 (N_5563,N_5124,N_5225);
nor U5564 (N_5564,N_5172,N_5399);
and U5565 (N_5565,N_5314,N_5078);
and U5566 (N_5566,N_5361,N_5125);
and U5567 (N_5567,N_5334,N_5482);
or U5568 (N_5568,N_5330,N_5340);
or U5569 (N_5569,N_5006,N_5120);
xor U5570 (N_5570,N_5423,N_5136);
nand U5571 (N_5571,N_5119,N_5141);
or U5572 (N_5572,N_5372,N_5271);
or U5573 (N_5573,N_5083,N_5351);
or U5574 (N_5574,N_5091,N_5341);
nand U5575 (N_5575,N_5065,N_5133);
or U5576 (N_5576,N_5328,N_5499);
and U5577 (N_5577,N_5481,N_5244);
and U5578 (N_5578,N_5142,N_5355);
or U5579 (N_5579,N_5056,N_5263);
nand U5580 (N_5580,N_5408,N_5255);
nand U5581 (N_5581,N_5126,N_5495);
nand U5582 (N_5582,N_5252,N_5233);
xnor U5583 (N_5583,N_5285,N_5486);
and U5584 (N_5584,N_5442,N_5153);
or U5585 (N_5585,N_5161,N_5194);
or U5586 (N_5586,N_5106,N_5165);
and U5587 (N_5587,N_5101,N_5431);
nor U5588 (N_5588,N_5224,N_5325);
nor U5589 (N_5589,N_5424,N_5131);
nor U5590 (N_5590,N_5184,N_5035);
and U5591 (N_5591,N_5401,N_5085);
or U5592 (N_5592,N_5227,N_5159);
nor U5593 (N_5593,N_5461,N_5039);
or U5594 (N_5594,N_5185,N_5405);
and U5595 (N_5595,N_5460,N_5207);
or U5596 (N_5596,N_5337,N_5280);
and U5597 (N_5597,N_5284,N_5307);
nand U5598 (N_5598,N_5466,N_5279);
nor U5599 (N_5599,N_5215,N_5036);
nor U5600 (N_5600,N_5430,N_5416);
or U5601 (N_5601,N_5333,N_5257);
nand U5602 (N_5602,N_5396,N_5470);
or U5603 (N_5603,N_5043,N_5391);
and U5604 (N_5604,N_5313,N_5202);
nor U5605 (N_5605,N_5462,N_5370);
nor U5606 (N_5606,N_5118,N_5196);
and U5607 (N_5607,N_5380,N_5021);
nor U5608 (N_5608,N_5005,N_5397);
nand U5609 (N_5609,N_5322,N_5072);
nor U5610 (N_5610,N_5169,N_5450);
nand U5611 (N_5611,N_5437,N_5052);
and U5612 (N_5612,N_5022,N_5182);
nor U5613 (N_5613,N_5028,N_5206);
nand U5614 (N_5614,N_5199,N_5066);
and U5615 (N_5615,N_5108,N_5229);
and U5616 (N_5616,N_5317,N_5336);
nand U5617 (N_5617,N_5080,N_5107);
or U5618 (N_5618,N_5102,N_5130);
and U5619 (N_5619,N_5472,N_5098);
or U5620 (N_5620,N_5029,N_5228);
nor U5621 (N_5621,N_5382,N_5071);
and U5622 (N_5622,N_5238,N_5203);
nand U5623 (N_5623,N_5353,N_5447);
nand U5624 (N_5624,N_5127,N_5393);
or U5625 (N_5625,N_5212,N_5268);
nor U5626 (N_5626,N_5293,N_5433);
nor U5627 (N_5627,N_5479,N_5451);
nor U5628 (N_5628,N_5222,N_5162);
nor U5629 (N_5629,N_5104,N_5230);
nor U5630 (N_5630,N_5249,N_5058);
or U5631 (N_5631,N_5109,N_5167);
nor U5632 (N_5632,N_5454,N_5013);
nor U5633 (N_5633,N_5445,N_5250);
and U5634 (N_5634,N_5177,N_5086);
and U5635 (N_5635,N_5371,N_5221);
nor U5636 (N_5636,N_5347,N_5076);
and U5637 (N_5637,N_5260,N_5220);
and U5638 (N_5638,N_5217,N_5282);
nor U5639 (N_5639,N_5289,N_5189);
nand U5640 (N_5640,N_5443,N_5132);
nand U5641 (N_5641,N_5223,N_5385);
and U5642 (N_5642,N_5432,N_5157);
nor U5643 (N_5643,N_5274,N_5003);
nand U5644 (N_5644,N_5409,N_5344);
or U5645 (N_5645,N_5294,N_5110);
nand U5646 (N_5646,N_5026,N_5415);
nand U5647 (N_5647,N_5356,N_5374);
nand U5648 (N_5648,N_5112,N_5259);
nand U5649 (N_5649,N_5264,N_5087);
nand U5650 (N_5650,N_5329,N_5308);
xor U5651 (N_5651,N_5327,N_5493);
or U5652 (N_5652,N_5231,N_5441);
nand U5653 (N_5653,N_5160,N_5180);
xnor U5654 (N_5654,N_5137,N_5375);
xnor U5655 (N_5655,N_5150,N_5497);
and U5656 (N_5656,N_5474,N_5315);
and U5657 (N_5657,N_5310,N_5487);
and U5658 (N_5658,N_5277,N_5105);
and U5659 (N_5659,N_5484,N_5241);
xnor U5660 (N_5660,N_5292,N_5266);
or U5661 (N_5661,N_5248,N_5338);
nand U5662 (N_5662,N_5323,N_5094);
or U5663 (N_5663,N_5358,N_5111);
and U5664 (N_5664,N_5253,N_5034);
and U5665 (N_5665,N_5384,N_5331);
nand U5666 (N_5666,N_5084,N_5491);
nand U5667 (N_5667,N_5236,N_5049);
nand U5668 (N_5668,N_5210,N_5097);
nor U5669 (N_5669,N_5046,N_5149);
nor U5670 (N_5670,N_5410,N_5201);
nand U5671 (N_5671,N_5187,N_5093);
nand U5672 (N_5672,N_5226,N_5218);
and U5673 (N_5673,N_5395,N_5418);
and U5674 (N_5674,N_5068,N_5440);
nor U5675 (N_5675,N_5316,N_5359);
and U5676 (N_5676,N_5175,N_5350);
nor U5677 (N_5677,N_5164,N_5275);
or U5678 (N_5678,N_5348,N_5179);
and U5679 (N_5679,N_5024,N_5425);
and U5680 (N_5680,N_5054,N_5457);
or U5681 (N_5681,N_5261,N_5148);
or U5682 (N_5682,N_5009,N_5269);
nand U5683 (N_5683,N_5234,N_5335);
nand U5684 (N_5684,N_5134,N_5291);
or U5685 (N_5685,N_5001,N_5387);
xor U5686 (N_5686,N_5090,N_5143);
nor U5687 (N_5687,N_5398,N_5471);
xnor U5688 (N_5688,N_5032,N_5077);
nand U5689 (N_5689,N_5151,N_5379);
or U5690 (N_5690,N_5452,N_5195);
nor U5691 (N_5691,N_5449,N_5188);
xnor U5692 (N_5692,N_5412,N_5422);
nand U5693 (N_5693,N_5305,N_5394);
nor U5694 (N_5694,N_5273,N_5042);
and U5695 (N_5695,N_5388,N_5490);
and U5696 (N_5696,N_5156,N_5057);
xnor U5697 (N_5697,N_5099,N_5473);
nand U5698 (N_5698,N_5128,N_5081);
nand U5699 (N_5699,N_5492,N_5299);
or U5700 (N_5700,N_5339,N_5050);
nand U5701 (N_5701,N_5476,N_5073);
nand U5702 (N_5702,N_5018,N_5209);
or U5703 (N_5703,N_5155,N_5286);
nand U5704 (N_5704,N_5376,N_5434);
nand U5705 (N_5705,N_5496,N_5365);
nand U5706 (N_5706,N_5278,N_5312);
or U5707 (N_5707,N_5421,N_5367);
and U5708 (N_5708,N_5369,N_5381);
nor U5709 (N_5709,N_5152,N_5067);
nand U5710 (N_5710,N_5404,N_5163);
and U5711 (N_5711,N_5113,N_5302);
or U5712 (N_5712,N_5413,N_5468);
nor U5713 (N_5713,N_5174,N_5123);
and U5714 (N_5714,N_5037,N_5360);
and U5715 (N_5715,N_5030,N_5319);
or U5716 (N_5716,N_5023,N_5346);
or U5717 (N_5717,N_5498,N_5200);
nor U5718 (N_5718,N_5298,N_5178);
xor U5719 (N_5719,N_5158,N_5242);
nand U5720 (N_5720,N_5045,N_5438);
nor U5721 (N_5721,N_5140,N_5357);
xor U5722 (N_5722,N_5332,N_5439);
and U5723 (N_5723,N_5326,N_5082);
nor U5724 (N_5724,N_5301,N_5092);
xor U5725 (N_5725,N_5258,N_5436);
nor U5726 (N_5726,N_5411,N_5240);
nand U5727 (N_5727,N_5219,N_5402);
nand U5728 (N_5728,N_5017,N_5191);
nor U5729 (N_5729,N_5008,N_5014);
nor U5730 (N_5730,N_5345,N_5349);
and U5731 (N_5731,N_5363,N_5208);
and U5732 (N_5732,N_5062,N_5304);
nor U5733 (N_5733,N_5235,N_5010);
xnor U5734 (N_5734,N_5467,N_5154);
or U5735 (N_5735,N_5256,N_5121);
or U5736 (N_5736,N_5012,N_5213);
nand U5737 (N_5737,N_5378,N_5446);
and U5738 (N_5738,N_5403,N_5407);
xnor U5739 (N_5739,N_5051,N_5232);
and U5740 (N_5740,N_5373,N_5427);
nor U5741 (N_5741,N_5041,N_5485);
or U5742 (N_5742,N_5147,N_5464);
nor U5743 (N_5743,N_5428,N_5390);
or U5744 (N_5744,N_5214,N_5459);
xnor U5745 (N_5745,N_5103,N_5122);
nand U5746 (N_5746,N_5287,N_5064);
nor U5747 (N_5747,N_5243,N_5205);
nand U5748 (N_5748,N_5469,N_5181);
or U5749 (N_5749,N_5377,N_5281);
nor U5750 (N_5750,N_5353,N_5085);
nand U5751 (N_5751,N_5173,N_5022);
and U5752 (N_5752,N_5422,N_5345);
and U5753 (N_5753,N_5031,N_5228);
and U5754 (N_5754,N_5200,N_5092);
nand U5755 (N_5755,N_5285,N_5266);
nand U5756 (N_5756,N_5256,N_5310);
and U5757 (N_5757,N_5045,N_5067);
or U5758 (N_5758,N_5388,N_5298);
or U5759 (N_5759,N_5071,N_5249);
and U5760 (N_5760,N_5093,N_5151);
nand U5761 (N_5761,N_5370,N_5439);
and U5762 (N_5762,N_5406,N_5172);
nand U5763 (N_5763,N_5280,N_5209);
or U5764 (N_5764,N_5016,N_5141);
or U5765 (N_5765,N_5227,N_5420);
and U5766 (N_5766,N_5328,N_5068);
nand U5767 (N_5767,N_5157,N_5160);
or U5768 (N_5768,N_5447,N_5199);
and U5769 (N_5769,N_5439,N_5051);
and U5770 (N_5770,N_5072,N_5355);
nor U5771 (N_5771,N_5141,N_5098);
or U5772 (N_5772,N_5295,N_5470);
nor U5773 (N_5773,N_5103,N_5368);
or U5774 (N_5774,N_5183,N_5169);
and U5775 (N_5775,N_5418,N_5473);
or U5776 (N_5776,N_5260,N_5345);
nand U5777 (N_5777,N_5370,N_5332);
nand U5778 (N_5778,N_5167,N_5332);
nand U5779 (N_5779,N_5332,N_5266);
nand U5780 (N_5780,N_5385,N_5027);
or U5781 (N_5781,N_5201,N_5137);
or U5782 (N_5782,N_5424,N_5375);
or U5783 (N_5783,N_5439,N_5443);
nor U5784 (N_5784,N_5207,N_5165);
or U5785 (N_5785,N_5226,N_5266);
nor U5786 (N_5786,N_5114,N_5069);
and U5787 (N_5787,N_5152,N_5487);
nor U5788 (N_5788,N_5012,N_5074);
xor U5789 (N_5789,N_5228,N_5256);
or U5790 (N_5790,N_5120,N_5073);
nor U5791 (N_5791,N_5427,N_5171);
or U5792 (N_5792,N_5295,N_5385);
or U5793 (N_5793,N_5352,N_5012);
nor U5794 (N_5794,N_5135,N_5137);
xnor U5795 (N_5795,N_5395,N_5276);
or U5796 (N_5796,N_5198,N_5169);
nor U5797 (N_5797,N_5322,N_5079);
or U5798 (N_5798,N_5151,N_5136);
nand U5799 (N_5799,N_5387,N_5216);
and U5800 (N_5800,N_5043,N_5102);
nand U5801 (N_5801,N_5131,N_5353);
or U5802 (N_5802,N_5199,N_5420);
xnor U5803 (N_5803,N_5341,N_5447);
and U5804 (N_5804,N_5142,N_5475);
or U5805 (N_5805,N_5318,N_5280);
nand U5806 (N_5806,N_5008,N_5499);
or U5807 (N_5807,N_5354,N_5011);
and U5808 (N_5808,N_5149,N_5165);
or U5809 (N_5809,N_5272,N_5331);
or U5810 (N_5810,N_5365,N_5095);
nor U5811 (N_5811,N_5048,N_5144);
nor U5812 (N_5812,N_5472,N_5077);
nor U5813 (N_5813,N_5294,N_5087);
or U5814 (N_5814,N_5048,N_5430);
xor U5815 (N_5815,N_5489,N_5354);
nand U5816 (N_5816,N_5395,N_5080);
nor U5817 (N_5817,N_5492,N_5229);
and U5818 (N_5818,N_5312,N_5490);
or U5819 (N_5819,N_5334,N_5111);
or U5820 (N_5820,N_5275,N_5298);
nor U5821 (N_5821,N_5132,N_5467);
or U5822 (N_5822,N_5431,N_5475);
nor U5823 (N_5823,N_5396,N_5303);
nor U5824 (N_5824,N_5332,N_5102);
and U5825 (N_5825,N_5060,N_5413);
nand U5826 (N_5826,N_5214,N_5026);
and U5827 (N_5827,N_5456,N_5088);
or U5828 (N_5828,N_5308,N_5144);
nand U5829 (N_5829,N_5297,N_5018);
and U5830 (N_5830,N_5489,N_5056);
and U5831 (N_5831,N_5368,N_5437);
and U5832 (N_5832,N_5182,N_5117);
nor U5833 (N_5833,N_5487,N_5275);
nor U5834 (N_5834,N_5080,N_5339);
or U5835 (N_5835,N_5131,N_5493);
and U5836 (N_5836,N_5393,N_5282);
and U5837 (N_5837,N_5402,N_5359);
nor U5838 (N_5838,N_5044,N_5243);
xnor U5839 (N_5839,N_5427,N_5345);
nor U5840 (N_5840,N_5175,N_5006);
or U5841 (N_5841,N_5280,N_5374);
nor U5842 (N_5842,N_5047,N_5142);
nor U5843 (N_5843,N_5346,N_5413);
nor U5844 (N_5844,N_5459,N_5002);
or U5845 (N_5845,N_5146,N_5345);
nor U5846 (N_5846,N_5244,N_5396);
and U5847 (N_5847,N_5228,N_5199);
and U5848 (N_5848,N_5406,N_5482);
or U5849 (N_5849,N_5190,N_5268);
and U5850 (N_5850,N_5047,N_5333);
nor U5851 (N_5851,N_5029,N_5384);
nor U5852 (N_5852,N_5220,N_5018);
or U5853 (N_5853,N_5226,N_5235);
or U5854 (N_5854,N_5184,N_5174);
and U5855 (N_5855,N_5044,N_5232);
and U5856 (N_5856,N_5438,N_5352);
nand U5857 (N_5857,N_5246,N_5240);
and U5858 (N_5858,N_5469,N_5348);
xor U5859 (N_5859,N_5337,N_5201);
nand U5860 (N_5860,N_5292,N_5060);
or U5861 (N_5861,N_5158,N_5241);
nand U5862 (N_5862,N_5161,N_5312);
nor U5863 (N_5863,N_5054,N_5006);
and U5864 (N_5864,N_5141,N_5461);
nand U5865 (N_5865,N_5404,N_5100);
nand U5866 (N_5866,N_5065,N_5216);
nand U5867 (N_5867,N_5338,N_5344);
and U5868 (N_5868,N_5179,N_5345);
xnor U5869 (N_5869,N_5093,N_5178);
and U5870 (N_5870,N_5115,N_5120);
nand U5871 (N_5871,N_5152,N_5246);
nor U5872 (N_5872,N_5424,N_5177);
nor U5873 (N_5873,N_5100,N_5454);
xnor U5874 (N_5874,N_5490,N_5058);
or U5875 (N_5875,N_5043,N_5173);
nor U5876 (N_5876,N_5280,N_5126);
and U5877 (N_5877,N_5120,N_5386);
nor U5878 (N_5878,N_5101,N_5224);
nor U5879 (N_5879,N_5119,N_5224);
or U5880 (N_5880,N_5106,N_5029);
xnor U5881 (N_5881,N_5003,N_5497);
or U5882 (N_5882,N_5423,N_5148);
and U5883 (N_5883,N_5032,N_5295);
nor U5884 (N_5884,N_5036,N_5117);
nor U5885 (N_5885,N_5201,N_5068);
nand U5886 (N_5886,N_5248,N_5014);
xor U5887 (N_5887,N_5246,N_5045);
nor U5888 (N_5888,N_5010,N_5236);
nand U5889 (N_5889,N_5234,N_5339);
and U5890 (N_5890,N_5208,N_5480);
xnor U5891 (N_5891,N_5197,N_5433);
nor U5892 (N_5892,N_5014,N_5332);
and U5893 (N_5893,N_5426,N_5210);
xor U5894 (N_5894,N_5089,N_5054);
xnor U5895 (N_5895,N_5068,N_5248);
or U5896 (N_5896,N_5495,N_5163);
nor U5897 (N_5897,N_5189,N_5452);
xor U5898 (N_5898,N_5350,N_5332);
nand U5899 (N_5899,N_5078,N_5378);
or U5900 (N_5900,N_5211,N_5499);
nor U5901 (N_5901,N_5293,N_5312);
or U5902 (N_5902,N_5091,N_5110);
xor U5903 (N_5903,N_5412,N_5430);
or U5904 (N_5904,N_5348,N_5239);
xnor U5905 (N_5905,N_5443,N_5484);
nor U5906 (N_5906,N_5269,N_5282);
and U5907 (N_5907,N_5216,N_5163);
xnor U5908 (N_5908,N_5071,N_5173);
nor U5909 (N_5909,N_5270,N_5221);
nand U5910 (N_5910,N_5267,N_5049);
xnor U5911 (N_5911,N_5228,N_5364);
nand U5912 (N_5912,N_5112,N_5448);
and U5913 (N_5913,N_5275,N_5195);
and U5914 (N_5914,N_5394,N_5247);
nand U5915 (N_5915,N_5148,N_5167);
xor U5916 (N_5916,N_5400,N_5452);
nor U5917 (N_5917,N_5024,N_5384);
nand U5918 (N_5918,N_5321,N_5284);
xnor U5919 (N_5919,N_5229,N_5250);
nor U5920 (N_5920,N_5212,N_5129);
or U5921 (N_5921,N_5015,N_5456);
nor U5922 (N_5922,N_5378,N_5243);
nand U5923 (N_5923,N_5047,N_5096);
nand U5924 (N_5924,N_5345,N_5305);
and U5925 (N_5925,N_5241,N_5073);
or U5926 (N_5926,N_5397,N_5393);
and U5927 (N_5927,N_5368,N_5163);
xor U5928 (N_5928,N_5364,N_5430);
nor U5929 (N_5929,N_5155,N_5196);
or U5930 (N_5930,N_5493,N_5113);
nor U5931 (N_5931,N_5142,N_5240);
and U5932 (N_5932,N_5221,N_5087);
xor U5933 (N_5933,N_5093,N_5361);
or U5934 (N_5934,N_5110,N_5353);
nor U5935 (N_5935,N_5308,N_5250);
nand U5936 (N_5936,N_5063,N_5400);
and U5937 (N_5937,N_5107,N_5244);
xnor U5938 (N_5938,N_5328,N_5324);
or U5939 (N_5939,N_5147,N_5479);
or U5940 (N_5940,N_5196,N_5055);
and U5941 (N_5941,N_5259,N_5240);
nor U5942 (N_5942,N_5385,N_5374);
nor U5943 (N_5943,N_5301,N_5105);
and U5944 (N_5944,N_5109,N_5121);
nand U5945 (N_5945,N_5061,N_5180);
xnor U5946 (N_5946,N_5016,N_5211);
nand U5947 (N_5947,N_5271,N_5215);
nand U5948 (N_5948,N_5393,N_5143);
xnor U5949 (N_5949,N_5330,N_5338);
nor U5950 (N_5950,N_5078,N_5038);
nor U5951 (N_5951,N_5458,N_5154);
xnor U5952 (N_5952,N_5260,N_5495);
or U5953 (N_5953,N_5177,N_5117);
nand U5954 (N_5954,N_5371,N_5428);
or U5955 (N_5955,N_5495,N_5341);
nand U5956 (N_5956,N_5343,N_5384);
nor U5957 (N_5957,N_5003,N_5135);
nand U5958 (N_5958,N_5290,N_5488);
nand U5959 (N_5959,N_5186,N_5034);
xnor U5960 (N_5960,N_5043,N_5139);
and U5961 (N_5961,N_5240,N_5056);
nand U5962 (N_5962,N_5341,N_5160);
xor U5963 (N_5963,N_5326,N_5434);
and U5964 (N_5964,N_5417,N_5488);
xor U5965 (N_5965,N_5397,N_5097);
and U5966 (N_5966,N_5022,N_5330);
nor U5967 (N_5967,N_5174,N_5241);
nor U5968 (N_5968,N_5000,N_5036);
nand U5969 (N_5969,N_5251,N_5414);
nor U5970 (N_5970,N_5290,N_5058);
nand U5971 (N_5971,N_5033,N_5128);
nor U5972 (N_5972,N_5011,N_5432);
nor U5973 (N_5973,N_5006,N_5452);
and U5974 (N_5974,N_5165,N_5144);
or U5975 (N_5975,N_5188,N_5186);
or U5976 (N_5976,N_5302,N_5430);
or U5977 (N_5977,N_5005,N_5244);
or U5978 (N_5978,N_5005,N_5457);
or U5979 (N_5979,N_5324,N_5029);
or U5980 (N_5980,N_5180,N_5099);
and U5981 (N_5981,N_5348,N_5364);
or U5982 (N_5982,N_5355,N_5024);
nand U5983 (N_5983,N_5112,N_5078);
nand U5984 (N_5984,N_5272,N_5107);
xor U5985 (N_5985,N_5060,N_5031);
nand U5986 (N_5986,N_5047,N_5481);
xnor U5987 (N_5987,N_5463,N_5074);
nand U5988 (N_5988,N_5454,N_5432);
and U5989 (N_5989,N_5000,N_5018);
or U5990 (N_5990,N_5477,N_5108);
nand U5991 (N_5991,N_5269,N_5052);
and U5992 (N_5992,N_5183,N_5045);
nor U5993 (N_5993,N_5471,N_5079);
or U5994 (N_5994,N_5097,N_5136);
and U5995 (N_5995,N_5014,N_5406);
nand U5996 (N_5996,N_5115,N_5372);
and U5997 (N_5997,N_5414,N_5226);
nor U5998 (N_5998,N_5094,N_5058);
nor U5999 (N_5999,N_5294,N_5086);
nor U6000 (N_6000,N_5772,N_5580);
and U6001 (N_6001,N_5854,N_5989);
nor U6002 (N_6002,N_5906,N_5513);
nand U6003 (N_6003,N_5996,N_5931);
xnor U6004 (N_6004,N_5883,N_5961);
nand U6005 (N_6005,N_5503,N_5540);
and U6006 (N_6006,N_5602,N_5633);
and U6007 (N_6007,N_5599,N_5914);
or U6008 (N_6008,N_5848,N_5588);
nor U6009 (N_6009,N_5977,N_5617);
and U6010 (N_6010,N_5751,N_5620);
and U6011 (N_6011,N_5797,N_5900);
nand U6012 (N_6012,N_5539,N_5837);
and U6013 (N_6013,N_5892,N_5814);
and U6014 (N_6014,N_5622,N_5581);
nand U6015 (N_6015,N_5926,N_5861);
nand U6016 (N_6016,N_5946,N_5608);
and U6017 (N_6017,N_5598,N_5770);
nand U6018 (N_6018,N_5986,N_5919);
and U6019 (N_6019,N_5849,N_5653);
nor U6020 (N_6020,N_5865,N_5952);
or U6021 (N_6021,N_5727,N_5781);
xnor U6022 (N_6022,N_5839,N_5817);
and U6023 (N_6023,N_5857,N_5557);
or U6024 (N_6024,N_5582,N_5612);
nand U6025 (N_6025,N_5502,N_5877);
nand U6026 (N_6026,N_5956,N_5934);
nor U6027 (N_6027,N_5594,N_5871);
nand U6028 (N_6028,N_5940,N_5542);
nand U6029 (N_6029,N_5881,N_5525);
nor U6030 (N_6030,N_5569,N_5529);
nor U6031 (N_6031,N_5512,N_5759);
nand U6032 (N_6032,N_5745,N_5994);
or U6033 (N_6033,N_5568,N_5530);
nand U6034 (N_6034,N_5606,N_5693);
nor U6035 (N_6035,N_5974,N_5955);
nand U6036 (N_6036,N_5958,N_5951);
nand U6037 (N_6037,N_5761,N_5673);
nor U6038 (N_6038,N_5538,N_5532);
and U6039 (N_6039,N_5533,N_5687);
and U6040 (N_6040,N_5636,N_5647);
and U6041 (N_6041,N_5743,N_5853);
nor U6042 (N_6042,N_5784,N_5595);
nor U6043 (N_6043,N_5860,N_5935);
nor U6044 (N_6044,N_5765,N_5624);
and U6045 (N_6045,N_5713,N_5921);
nand U6046 (N_6046,N_5695,N_5771);
or U6047 (N_6047,N_5845,N_5941);
nor U6048 (N_6048,N_5630,N_5559);
and U6049 (N_6049,N_5916,N_5889);
nand U6050 (N_6050,N_5615,N_5783);
and U6051 (N_6051,N_5963,N_5516);
and U6052 (N_6052,N_5920,N_5721);
xnor U6053 (N_6053,N_5988,N_5555);
nor U6054 (N_6054,N_5894,N_5619);
or U6055 (N_6055,N_5739,N_5616);
nor U6056 (N_6056,N_5634,N_5810);
and U6057 (N_6057,N_5520,N_5524);
nor U6058 (N_6058,N_5717,N_5651);
and U6059 (N_6059,N_5950,N_5938);
or U6060 (N_6060,N_5790,N_5901);
or U6061 (N_6061,N_5782,N_5930);
xor U6062 (N_6062,N_5878,N_5862);
xor U6063 (N_6063,N_5815,N_5874);
or U6064 (N_6064,N_5800,N_5678);
nand U6065 (N_6065,N_5627,N_5789);
and U6066 (N_6066,N_5903,N_5980);
and U6067 (N_6067,N_5700,N_5546);
and U6068 (N_6068,N_5998,N_5644);
nand U6069 (N_6069,N_5689,N_5942);
or U6070 (N_6070,N_5613,N_5811);
nor U6071 (N_6071,N_5902,N_5666);
nand U6072 (N_6072,N_5749,N_5798);
nor U6073 (N_6073,N_5893,N_5600);
xor U6074 (N_6074,N_5614,N_5587);
and U6075 (N_6075,N_5913,N_5726);
nor U6076 (N_6076,N_5976,N_5688);
nand U6077 (N_6077,N_5631,N_5709);
and U6078 (N_6078,N_5589,N_5777);
nor U6079 (N_6079,N_5823,N_5659);
xor U6080 (N_6080,N_5758,N_5660);
xor U6081 (N_6081,N_5850,N_5668);
nand U6082 (N_6082,N_5718,N_5891);
or U6083 (N_6083,N_5866,N_5596);
nor U6084 (N_6084,N_5975,N_5623);
and U6085 (N_6085,N_5795,N_5820);
nor U6086 (N_6086,N_5957,N_5677);
or U6087 (N_6087,N_5869,N_5806);
nor U6088 (N_6088,N_5729,N_5775);
nor U6089 (N_6089,N_5640,N_5646);
nand U6090 (N_6090,N_5522,N_5933);
nand U6091 (N_6091,N_5698,N_5735);
xor U6092 (N_6092,N_5769,N_5887);
nor U6093 (N_6093,N_5551,N_5686);
xor U6094 (N_6094,N_5669,N_5740);
nor U6095 (N_6095,N_5899,N_5534);
xor U6096 (N_6096,N_5875,N_5995);
and U6097 (N_6097,N_5960,N_5697);
and U6098 (N_6098,N_5809,N_5791);
nand U6099 (N_6099,N_5564,N_5939);
nand U6100 (N_6100,N_5852,N_5964);
or U6101 (N_6101,N_5683,N_5936);
or U6102 (N_6102,N_5645,N_5872);
nor U6103 (N_6103,N_5999,N_5763);
or U6104 (N_6104,N_5937,N_5571);
or U6105 (N_6105,N_5734,N_5928);
or U6106 (N_6106,N_5954,N_5519);
nor U6107 (N_6107,N_5566,N_5609);
nand U6108 (N_6108,N_5641,N_5802);
or U6109 (N_6109,N_5774,N_5720);
or U6110 (N_6110,N_5707,N_5663);
nand U6111 (N_6111,N_5505,N_5573);
and U6112 (N_6112,N_5510,N_5703);
and U6113 (N_6113,N_5825,N_5738);
nor U6114 (N_6114,N_5842,N_5843);
xor U6115 (N_6115,N_5922,N_5731);
xor U6116 (N_6116,N_5808,N_5873);
nor U6117 (N_6117,N_5694,N_5927);
nor U6118 (N_6118,N_5674,N_5643);
and U6119 (N_6119,N_5741,N_5984);
or U6120 (N_6120,N_5511,N_5838);
and U6121 (N_6121,N_5544,N_5728);
nand U6122 (N_6122,N_5780,N_5671);
nor U6123 (N_6123,N_5699,N_5835);
nor U6124 (N_6124,N_5767,N_5805);
nand U6125 (N_6125,N_5621,N_5696);
nor U6126 (N_6126,N_5945,N_5563);
xor U6127 (N_6127,N_5679,N_5549);
and U6128 (N_6128,N_5685,N_5744);
or U6129 (N_6129,N_5545,N_5724);
nand U6130 (N_6130,N_5895,N_5792);
or U6131 (N_6131,N_5577,N_5670);
and U6132 (N_6132,N_5585,N_5796);
nand U6133 (N_6133,N_5509,N_5567);
nor U6134 (N_6134,N_5846,N_5658);
and U6135 (N_6135,N_5553,N_5905);
and U6136 (N_6136,N_5867,N_5526);
xor U6137 (N_6137,N_5704,N_5654);
xor U6138 (N_6138,N_5605,N_5982);
xnor U6139 (N_6139,N_5824,N_5822);
nand U6140 (N_6140,N_5932,N_5711);
nor U6141 (N_6141,N_5725,N_5924);
or U6142 (N_6142,N_5550,N_5672);
nand U6143 (N_6143,N_5650,N_5702);
nand U6144 (N_6144,N_5968,N_5884);
nand U6145 (N_6145,N_5722,N_5625);
nor U6146 (N_6146,N_5912,N_5818);
nor U6147 (N_6147,N_5821,N_5858);
and U6148 (N_6148,N_5909,N_5682);
nor U6149 (N_6149,N_5705,N_5570);
xor U6150 (N_6150,N_5528,N_5723);
or U6151 (N_6151,N_5742,N_5579);
and U6152 (N_6152,N_5890,N_5748);
nor U6153 (N_6153,N_5733,N_5779);
nand U6154 (N_6154,N_5736,N_5537);
nand U6155 (N_6155,N_5879,N_5925);
nor U6156 (N_6156,N_5870,N_5828);
and U6157 (N_6157,N_5863,N_5584);
xor U6158 (N_6158,N_5819,N_5959);
nor U6159 (N_6159,N_5886,N_5788);
and U6160 (N_6160,N_5506,N_5628);
xnor U6161 (N_6161,N_5990,N_5786);
or U6162 (N_6162,N_5969,N_5868);
nand U6163 (N_6163,N_5910,N_5943);
nor U6164 (N_6164,N_5991,N_5536);
nor U6165 (N_6165,N_5607,N_5755);
xnor U6166 (N_6166,N_5841,N_5799);
nand U6167 (N_6167,N_5592,N_5560);
xnor U6168 (N_6168,N_5514,N_5948);
or U6169 (N_6169,N_5970,N_5561);
nand U6170 (N_6170,N_5662,N_5649);
or U6171 (N_6171,N_5690,N_5701);
nor U6172 (N_6172,N_5665,N_5915);
and U6173 (N_6173,N_5541,N_5675);
or U6174 (N_6174,N_5543,N_5547);
and U6175 (N_6175,N_5527,N_5760);
and U6176 (N_6176,N_5898,N_5972);
nand U6177 (N_6177,N_5556,N_5642);
and U6178 (N_6178,N_5750,N_5766);
nor U6179 (N_6179,N_5629,N_5967);
or U6180 (N_6180,N_5656,N_5987);
nand U6181 (N_6181,N_5813,N_5856);
or U6182 (N_6182,N_5929,N_5876);
nand U6183 (N_6183,N_5586,N_5997);
nand U6184 (N_6184,N_5635,N_5712);
and U6185 (N_6185,N_5896,N_5501);
nand U6186 (N_6186,N_5716,N_5844);
and U6187 (N_6187,N_5680,N_5832);
nand U6188 (N_6188,N_5552,N_5554);
nand U6189 (N_6189,N_5667,N_5661);
or U6190 (N_6190,N_5637,N_5830);
nor U6191 (N_6191,N_5773,N_5639);
nor U6192 (N_6192,N_5985,N_5523);
or U6193 (N_6193,N_5993,N_5826);
nand U6194 (N_6194,N_5962,N_5710);
or U6195 (N_6195,N_5562,N_5953);
nor U6196 (N_6196,N_5804,N_5575);
nor U6197 (N_6197,N_5730,N_5973);
xor U6198 (N_6198,N_5840,N_5855);
or U6199 (N_6199,N_5882,N_5803);
nor U6200 (N_6200,N_5611,N_5508);
xnor U6201 (N_6201,N_5531,N_5746);
nand U6202 (N_6202,N_5632,N_5681);
nor U6203 (N_6203,N_5732,N_5518);
nor U6204 (N_6204,N_5708,N_5831);
and U6205 (N_6205,N_5923,N_5816);
and U6206 (N_6206,N_5715,N_5807);
and U6207 (N_6207,N_5747,N_5836);
and U6208 (N_6208,N_5603,N_5944);
and U6209 (N_6209,N_5983,N_5676);
nor U6210 (N_6210,N_5753,N_5572);
xnor U6211 (N_6211,N_5981,N_5979);
nor U6212 (N_6212,N_5500,N_5648);
xor U6213 (N_6213,N_5576,N_5578);
and U6214 (N_6214,N_5908,N_5827);
nor U6215 (N_6215,N_5719,N_5591);
or U6216 (N_6216,N_5911,N_5864);
nor U6217 (N_6217,N_5618,N_5558);
or U6218 (N_6218,N_5778,N_5978);
or U6219 (N_6219,N_5638,N_5655);
or U6220 (N_6220,N_5504,N_5664);
and U6221 (N_6221,N_5949,N_5657);
or U6222 (N_6222,N_5907,N_5992);
or U6223 (N_6223,N_5762,N_5764);
or U6224 (N_6224,N_5847,N_5583);
xor U6225 (N_6225,N_5601,N_5597);
and U6226 (N_6226,N_5917,N_5918);
and U6227 (N_6227,N_5851,N_5888);
nand U6228 (N_6228,N_5754,N_5829);
nor U6229 (N_6229,N_5785,N_5515);
and U6230 (N_6230,N_5684,N_5691);
nand U6231 (N_6231,N_5706,N_5971);
or U6232 (N_6232,N_5593,N_5517);
nor U6233 (N_6233,N_5507,N_5521);
nor U6234 (N_6234,N_5965,N_5610);
nor U6235 (N_6235,N_5626,N_5947);
or U6236 (N_6236,N_5833,N_5768);
and U6237 (N_6237,N_5757,N_5904);
and U6238 (N_6238,N_5590,N_5776);
nor U6239 (N_6239,N_5880,N_5859);
or U6240 (N_6240,N_5714,N_5794);
nor U6241 (N_6241,N_5692,N_5752);
nand U6242 (N_6242,N_5565,N_5793);
nor U6243 (N_6243,N_5812,N_5801);
or U6244 (N_6244,N_5897,N_5652);
nand U6245 (N_6245,N_5604,N_5737);
nand U6246 (N_6246,N_5548,N_5756);
nor U6247 (N_6247,N_5787,N_5574);
and U6248 (N_6248,N_5535,N_5834);
nand U6249 (N_6249,N_5885,N_5966);
nand U6250 (N_6250,N_5951,N_5914);
or U6251 (N_6251,N_5622,N_5769);
nand U6252 (N_6252,N_5995,N_5700);
or U6253 (N_6253,N_5779,N_5514);
and U6254 (N_6254,N_5891,N_5977);
or U6255 (N_6255,N_5521,N_5667);
nand U6256 (N_6256,N_5576,N_5597);
or U6257 (N_6257,N_5880,N_5820);
and U6258 (N_6258,N_5812,N_5649);
nand U6259 (N_6259,N_5880,N_5597);
or U6260 (N_6260,N_5547,N_5542);
and U6261 (N_6261,N_5977,N_5985);
or U6262 (N_6262,N_5866,N_5946);
nand U6263 (N_6263,N_5544,N_5858);
and U6264 (N_6264,N_5978,N_5644);
and U6265 (N_6265,N_5784,N_5893);
nor U6266 (N_6266,N_5871,N_5574);
xnor U6267 (N_6267,N_5849,N_5598);
and U6268 (N_6268,N_5747,N_5970);
nor U6269 (N_6269,N_5715,N_5939);
or U6270 (N_6270,N_5981,N_5651);
and U6271 (N_6271,N_5563,N_5836);
nor U6272 (N_6272,N_5880,N_5685);
nor U6273 (N_6273,N_5725,N_5876);
nand U6274 (N_6274,N_5504,N_5950);
and U6275 (N_6275,N_5571,N_5543);
xnor U6276 (N_6276,N_5938,N_5550);
nand U6277 (N_6277,N_5500,N_5707);
nand U6278 (N_6278,N_5901,N_5594);
xor U6279 (N_6279,N_5630,N_5821);
nor U6280 (N_6280,N_5547,N_5947);
nor U6281 (N_6281,N_5775,N_5861);
nor U6282 (N_6282,N_5597,N_5893);
or U6283 (N_6283,N_5620,N_5916);
nand U6284 (N_6284,N_5501,N_5864);
and U6285 (N_6285,N_5641,N_5979);
or U6286 (N_6286,N_5562,N_5533);
and U6287 (N_6287,N_5974,N_5640);
nor U6288 (N_6288,N_5824,N_5889);
and U6289 (N_6289,N_5842,N_5522);
xor U6290 (N_6290,N_5542,N_5784);
nor U6291 (N_6291,N_5652,N_5780);
nor U6292 (N_6292,N_5560,N_5936);
nor U6293 (N_6293,N_5870,N_5986);
or U6294 (N_6294,N_5569,N_5940);
or U6295 (N_6295,N_5763,N_5641);
xor U6296 (N_6296,N_5733,N_5546);
nand U6297 (N_6297,N_5777,N_5585);
xnor U6298 (N_6298,N_5856,N_5864);
or U6299 (N_6299,N_5819,N_5855);
xnor U6300 (N_6300,N_5566,N_5721);
nand U6301 (N_6301,N_5872,N_5987);
nand U6302 (N_6302,N_5595,N_5658);
or U6303 (N_6303,N_5564,N_5720);
nand U6304 (N_6304,N_5554,N_5522);
or U6305 (N_6305,N_5562,N_5932);
nand U6306 (N_6306,N_5866,N_5616);
xnor U6307 (N_6307,N_5871,N_5971);
or U6308 (N_6308,N_5739,N_5973);
and U6309 (N_6309,N_5659,N_5928);
or U6310 (N_6310,N_5654,N_5783);
nand U6311 (N_6311,N_5678,N_5953);
and U6312 (N_6312,N_5562,N_5882);
nand U6313 (N_6313,N_5913,N_5542);
xnor U6314 (N_6314,N_5529,N_5827);
and U6315 (N_6315,N_5924,N_5687);
nand U6316 (N_6316,N_5521,N_5931);
and U6317 (N_6317,N_5781,N_5671);
nand U6318 (N_6318,N_5503,N_5534);
and U6319 (N_6319,N_5707,N_5618);
nor U6320 (N_6320,N_5741,N_5927);
or U6321 (N_6321,N_5797,N_5612);
nor U6322 (N_6322,N_5639,N_5522);
and U6323 (N_6323,N_5506,N_5725);
xor U6324 (N_6324,N_5861,N_5520);
nor U6325 (N_6325,N_5984,N_5665);
and U6326 (N_6326,N_5764,N_5857);
nand U6327 (N_6327,N_5869,N_5873);
nor U6328 (N_6328,N_5654,N_5599);
nor U6329 (N_6329,N_5500,N_5636);
nor U6330 (N_6330,N_5951,N_5824);
nand U6331 (N_6331,N_5880,N_5637);
nor U6332 (N_6332,N_5568,N_5731);
nor U6333 (N_6333,N_5628,N_5816);
or U6334 (N_6334,N_5813,N_5917);
and U6335 (N_6335,N_5664,N_5944);
nor U6336 (N_6336,N_5543,N_5704);
or U6337 (N_6337,N_5897,N_5873);
and U6338 (N_6338,N_5815,N_5675);
nor U6339 (N_6339,N_5568,N_5768);
nor U6340 (N_6340,N_5886,N_5778);
nor U6341 (N_6341,N_5556,N_5656);
or U6342 (N_6342,N_5540,N_5772);
nand U6343 (N_6343,N_5885,N_5973);
and U6344 (N_6344,N_5690,N_5614);
or U6345 (N_6345,N_5702,N_5722);
nand U6346 (N_6346,N_5706,N_5961);
nor U6347 (N_6347,N_5975,N_5708);
nand U6348 (N_6348,N_5672,N_5660);
nor U6349 (N_6349,N_5984,N_5955);
nand U6350 (N_6350,N_5570,N_5763);
or U6351 (N_6351,N_5896,N_5512);
and U6352 (N_6352,N_5630,N_5617);
nand U6353 (N_6353,N_5959,N_5983);
nand U6354 (N_6354,N_5801,N_5625);
nand U6355 (N_6355,N_5960,N_5633);
and U6356 (N_6356,N_5718,N_5657);
or U6357 (N_6357,N_5890,N_5796);
and U6358 (N_6358,N_5880,N_5515);
nor U6359 (N_6359,N_5696,N_5587);
or U6360 (N_6360,N_5891,N_5558);
or U6361 (N_6361,N_5506,N_5919);
nand U6362 (N_6362,N_5695,N_5596);
and U6363 (N_6363,N_5747,N_5826);
or U6364 (N_6364,N_5511,N_5556);
nor U6365 (N_6365,N_5519,N_5993);
or U6366 (N_6366,N_5895,N_5546);
or U6367 (N_6367,N_5660,N_5503);
or U6368 (N_6368,N_5603,N_5662);
nor U6369 (N_6369,N_5628,N_5907);
nor U6370 (N_6370,N_5576,N_5807);
nor U6371 (N_6371,N_5698,N_5670);
and U6372 (N_6372,N_5593,N_5549);
nand U6373 (N_6373,N_5597,N_5897);
nand U6374 (N_6374,N_5804,N_5592);
nand U6375 (N_6375,N_5887,N_5943);
or U6376 (N_6376,N_5907,N_5751);
xnor U6377 (N_6377,N_5791,N_5789);
and U6378 (N_6378,N_5967,N_5692);
nor U6379 (N_6379,N_5741,N_5955);
xor U6380 (N_6380,N_5652,N_5606);
nor U6381 (N_6381,N_5867,N_5685);
nor U6382 (N_6382,N_5806,N_5560);
and U6383 (N_6383,N_5840,N_5680);
or U6384 (N_6384,N_5563,N_5630);
or U6385 (N_6385,N_5569,N_5677);
nor U6386 (N_6386,N_5647,N_5598);
nand U6387 (N_6387,N_5828,N_5846);
nor U6388 (N_6388,N_5614,N_5823);
or U6389 (N_6389,N_5533,N_5891);
xor U6390 (N_6390,N_5871,N_5845);
or U6391 (N_6391,N_5572,N_5935);
nor U6392 (N_6392,N_5803,N_5572);
or U6393 (N_6393,N_5518,N_5854);
nor U6394 (N_6394,N_5966,N_5710);
or U6395 (N_6395,N_5766,N_5538);
nand U6396 (N_6396,N_5605,N_5903);
nand U6397 (N_6397,N_5668,N_5561);
or U6398 (N_6398,N_5823,N_5999);
nand U6399 (N_6399,N_5877,N_5572);
or U6400 (N_6400,N_5876,N_5581);
and U6401 (N_6401,N_5848,N_5693);
nand U6402 (N_6402,N_5915,N_5773);
nand U6403 (N_6403,N_5520,N_5748);
nor U6404 (N_6404,N_5665,N_5789);
nand U6405 (N_6405,N_5859,N_5877);
or U6406 (N_6406,N_5754,N_5538);
or U6407 (N_6407,N_5611,N_5892);
nand U6408 (N_6408,N_5500,N_5689);
or U6409 (N_6409,N_5912,N_5693);
or U6410 (N_6410,N_5968,N_5876);
xnor U6411 (N_6411,N_5773,N_5583);
nand U6412 (N_6412,N_5861,N_5725);
nor U6413 (N_6413,N_5799,N_5862);
nor U6414 (N_6414,N_5892,N_5823);
nor U6415 (N_6415,N_5887,N_5930);
or U6416 (N_6416,N_5887,N_5610);
xnor U6417 (N_6417,N_5771,N_5587);
nand U6418 (N_6418,N_5974,N_5691);
nor U6419 (N_6419,N_5670,N_5751);
nor U6420 (N_6420,N_5890,N_5616);
xnor U6421 (N_6421,N_5534,N_5709);
and U6422 (N_6422,N_5639,N_5793);
or U6423 (N_6423,N_5518,N_5748);
or U6424 (N_6424,N_5725,N_5571);
and U6425 (N_6425,N_5841,N_5696);
nor U6426 (N_6426,N_5918,N_5629);
nor U6427 (N_6427,N_5877,N_5693);
or U6428 (N_6428,N_5816,N_5505);
nor U6429 (N_6429,N_5516,N_5642);
or U6430 (N_6430,N_5604,N_5525);
xor U6431 (N_6431,N_5560,N_5610);
nand U6432 (N_6432,N_5712,N_5581);
or U6433 (N_6433,N_5824,N_5767);
or U6434 (N_6434,N_5721,N_5523);
nand U6435 (N_6435,N_5873,N_5909);
or U6436 (N_6436,N_5980,N_5548);
and U6437 (N_6437,N_5528,N_5987);
nand U6438 (N_6438,N_5973,N_5718);
nor U6439 (N_6439,N_5905,N_5507);
nand U6440 (N_6440,N_5565,N_5625);
and U6441 (N_6441,N_5544,N_5932);
xor U6442 (N_6442,N_5827,N_5862);
nor U6443 (N_6443,N_5934,N_5836);
xnor U6444 (N_6444,N_5736,N_5982);
or U6445 (N_6445,N_5763,N_5503);
xnor U6446 (N_6446,N_5898,N_5600);
and U6447 (N_6447,N_5587,N_5812);
nand U6448 (N_6448,N_5537,N_5841);
and U6449 (N_6449,N_5755,N_5955);
nor U6450 (N_6450,N_5871,N_5839);
nor U6451 (N_6451,N_5557,N_5624);
and U6452 (N_6452,N_5723,N_5607);
xor U6453 (N_6453,N_5911,N_5700);
xnor U6454 (N_6454,N_5895,N_5552);
and U6455 (N_6455,N_5791,N_5749);
nand U6456 (N_6456,N_5596,N_5991);
nand U6457 (N_6457,N_5771,N_5667);
and U6458 (N_6458,N_5737,N_5610);
nor U6459 (N_6459,N_5572,N_5606);
or U6460 (N_6460,N_5617,N_5594);
nor U6461 (N_6461,N_5804,N_5935);
nand U6462 (N_6462,N_5772,N_5699);
or U6463 (N_6463,N_5879,N_5856);
or U6464 (N_6464,N_5770,N_5832);
or U6465 (N_6465,N_5786,N_5653);
and U6466 (N_6466,N_5986,N_5980);
nand U6467 (N_6467,N_5674,N_5585);
or U6468 (N_6468,N_5502,N_5884);
or U6469 (N_6469,N_5685,N_5911);
or U6470 (N_6470,N_5949,N_5708);
or U6471 (N_6471,N_5513,N_5902);
nor U6472 (N_6472,N_5523,N_5590);
nand U6473 (N_6473,N_5805,N_5753);
nor U6474 (N_6474,N_5530,N_5738);
and U6475 (N_6475,N_5562,N_5595);
and U6476 (N_6476,N_5719,N_5557);
nor U6477 (N_6477,N_5735,N_5998);
or U6478 (N_6478,N_5514,N_5855);
xnor U6479 (N_6479,N_5835,N_5671);
or U6480 (N_6480,N_5953,N_5965);
or U6481 (N_6481,N_5809,N_5794);
or U6482 (N_6482,N_5757,N_5888);
xnor U6483 (N_6483,N_5541,N_5633);
and U6484 (N_6484,N_5561,N_5873);
and U6485 (N_6485,N_5583,N_5951);
nor U6486 (N_6486,N_5883,N_5511);
nor U6487 (N_6487,N_5758,N_5568);
and U6488 (N_6488,N_5824,N_5780);
nor U6489 (N_6489,N_5908,N_5625);
nand U6490 (N_6490,N_5908,N_5881);
nor U6491 (N_6491,N_5901,N_5898);
xor U6492 (N_6492,N_5725,N_5807);
or U6493 (N_6493,N_5665,N_5631);
nor U6494 (N_6494,N_5989,N_5790);
nand U6495 (N_6495,N_5894,N_5553);
and U6496 (N_6496,N_5652,N_5514);
nand U6497 (N_6497,N_5788,N_5599);
nand U6498 (N_6498,N_5607,N_5916);
and U6499 (N_6499,N_5511,N_5793);
or U6500 (N_6500,N_6217,N_6020);
nand U6501 (N_6501,N_6259,N_6035);
xor U6502 (N_6502,N_6272,N_6188);
or U6503 (N_6503,N_6482,N_6422);
and U6504 (N_6504,N_6431,N_6483);
nor U6505 (N_6505,N_6164,N_6110);
xnor U6506 (N_6506,N_6372,N_6299);
xor U6507 (N_6507,N_6406,N_6173);
nand U6508 (N_6508,N_6413,N_6391);
nor U6509 (N_6509,N_6244,N_6425);
nand U6510 (N_6510,N_6092,N_6353);
or U6511 (N_6511,N_6449,N_6377);
nor U6512 (N_6512,N_6122,N_6388);
nor U6513 (N_6513,N_6415,N_6010);
nand U6514 (N_6514,N_6403,N_6338);
and U6515 (N_6515,N_6396,N_6261);
xnor U6516 (N_6516,N_6432,N_6202);
and U6517 (N_6517,N_6447,N_6079);
and U6518 (N_6518,N_6021,N_6038);
nand U6519 (N_6519,N_6424,N_6012);
or U6520 (N_6520,N_6118,N_6381);
nand U6521 (N_6521,N_6374,N_6446);
or U6522 (N_6522,N_6076,N_6210);
or U6523 (N_6523,N_6416,N_6102);
nor U6524 (N_6524,N_6354,N_6105);
or U6525 (N_6525,N_6114,N_6286);
and U6526 (N_6526,N_6480,N_6131);
and U6527 (N_6527,N_6022,N_6045);
or U6528 (N_6528,N_6086,N_6274);
and U6529 (N_6529,N_6130,N_6183);
xnor U6530 (N_6530,N_6078,N_6383);
nor U6531 (N_6531,N_6082,N_6247);
and U6532 (N_6532,N_6298,N_6084);
xor U6533 (N_6533,N_6484,N_6243);
nand U6534 (N_6534,N_6269,N_6225);
or U6535 (N_6535,N_6040,N_6313);
nor U6536 (N_6536,N_6072,N_6463);
nor U6537 (N_6537,N_6429,N_6124);
nor U6538 (N_6538,N_6363,N_6440);
nand U6539 (N_6539,N_6442,N_6062);
and U6540 (N_6540,N_6350,N_6435);
nor U6541 (N_6541,N_6113,N_6450);
nor U6542 (N_6542,N_6170,N_6264);
or U6543 (N_6543,N_6239,N_6467);
or U6544 (N_6544,N_6410,N_6158);
nor U6545 (N_6545,N_6250,N_6287);
nand U6546 (N_6546,N_6234,N_6224);
and U6547 (N_6547,N_6065,N_6461);
and U6548 (N_6548,N_6324,N_6481);
nand U6549 (N_6549,N_6074,N_6209);
and U6550 (N_6550,N_6211,N_6328);
nor U6551 (N_6551,N_6400,N_6077);
and U6552 (N_6552,N_6493,N_6491);
nand U6553 (N_6553,N_6140,N_6139);
nor U6554 (N_6554,N_6051,N_6266);
or U6555 (N_6555,N_6176,N_6218);
and U6556 (N_6556,N_6448,N_6094);
and U6557 (N_6557,N_6352,N_6312);
or U6558 (N_6558,N_6314,N_6276);
and U6559 (N_6559,N_6418,N_6223);
nand U6560 (N_6560,N_6064,N_6334);
or U6561 (N_6561,N_6121,N_6071);
nor U6562 (N_6562,N_6166,N_6154);
xnor U6563 (N_6563,N_6117,N_6115);
nand U6564 (N_6564,N_6497,N_6228);
and U6565 (N_6565,N_6364,N_6112);
nand U6566 (N_6566,N_6231,N_6143);
nand U6567 (N_6567,N_6123,N_6277);
and U6568 (N_6568,N_6411,N_6433);
or U6569 (N_6569,N_6219,N_6235);
nor U6570 (N_6570,N_6236,N_6392);
and U6571 (N_6571,N_6018,N_6355);
nand U6572 (N_6572,N_6394,N_6382);
nor U6573 (N_6573,N_6190,N_6376);
nor U6574 (N_6574,N_6428,N_6023);
nor U6575 (N_6575,N_6310,N_6362);
nor U6576 (N_6576,N_6007,N_6460);
and U6577 (N_6577,N_6050,N_6144);
nand U6578 (N_6578,N_6181,N_6241);
or U6579 (N_6579,N_6380,N_6260);
nand U6580 (N_6580,N_6329,N_6367);
and U6581 (N_6581,N_6061,N_6233);
and U6582 (N_6582,N_6060,N_6054);
nor U6583 (N_6583,N_6306,N_6301);
or U6584 (N_6584,N_6271,N_6280);
nand U6585 (N_6585,N_6366,N_6017);
nand U6586 (N_6586,N_6066,N_6304);
nand U6587 (N_6587,N_6308,N_6278);
or U6588 (N_6588,N_6436,N_6451);
or U6589 (N_6589,N_6297,N_6348);
or U6590 (N_6590,N_6152,N_6255);
or U6591 (N_6591,N_6098,N_6275);
nor U6592 (N_6592,N_6343,N_6133);
nor U6593 (N_6593,N_6437,N_6474);
or U6594 (N_6594,N_6052,N_6371);
xnor U6595 (N_6595,N_6330,N_6232);
xor U6596 (N_6596,N_6126,N_6254);
nor U6597 (N_6597,N_6387,N_6339);
and U6598 (N_6598,N_6138,N_6091);
nand U6599 (N_6599,N_6412,N_6470);
xnor U6600 (N_6600,N_6475,N_6195);
nand U6601 (N_6601,N_6466,N_6000);
xnor U6602 (N_6602,N_6373,N_6457);
xnor U6603 (N_6603,N_6057,N_6189);
or U6604 (N_6604,N_6002,N_6119);
or U6605 (N_6605,N_6495,N_6033);
or U6606 (N_6606,N_6423,N_6025);
nand U6607 (N_6607,N_6384,N_6081);
or U6608 (N_6608,N_6171,N_6162);
nand U6609 (N_6609,N_6014,N_6279);
or U6610 (N_6610,N_6351,N_6427);
and U6611 (N_6611,N_6494,N_6197);
or U6612 (N_6612,N_6193,N_6068);
nand U6613 (N_6613,N_6430,N_6016);
or U6614 (N_6614,N_6331,N_6032);
or U6615 (N_6615,N_6201,N_6159);
or U6616 (N_6616,N_6358,N_6095);
and U6617 (N_6617,N_6186,N_6284);
nand U6618 (N_6618,N_6004,N_6069);
or U6619 (N_6619,N_6393,N_6178);
and U6620 (N_6620,N_6125,N_6342);
nand U6621 (N_6621,N_6320,N_6359);
nand U6622 (N_6622,N_6325,N_6498);
xnor U6623 (N_6623,N_6456,N_6356);
nand U6624 (N_6624,N_6489,N_6281);
nand U6625 (N_6625,N_6473,N_6370);
nor U6626 (N_6626,N_6464,N_6408);
and U6627 (N_6627,N_6478,N_6097);
xor U6628 (N_6628,N_6345,N_6175);
xor U6629 (N_6629,N_6414,N_6289);
and U6630 (N_6630,N_6127,N_6208);
or U6631 (N_6631,N_6056,N_6246);
and U6632 (N_6632,N_6116,N_6379);
nor U6633 (N_6633,N_6398,N_6237);
and U6634 (N_6634,N_6177,N_6333);
nor U6635 (N_6635,N_6009,N_6222);
nor U6636 (N_6636,N_6147,N_6341);
and U6637 (N_6637,N_6439,N_6302);
xnor U6638 (N_6638,N_6469,N_6148);
xor U6639 (N_6639,N_6198,N_6088);
and U6640 (N_6640,N_6108,N_6137);
nand U6641 (N_6641,N_6245,N_6361);
xor U6642 (N_6642,N_6389,N_6141);
nand U6643 (N_6643,N_6047,N_6103);
nand U6644 (N_6644,N_6283,N_6323);
or U6645 (N_6645,N_6100,N_6317);
nand U6646 (N_6646,N_6340,N_6397);
or U6647 (N_6647,N_6149,N_6263);
and U6648 (N_6648,N_6434,N_6215);
and U6649 (N_6649,N_6042,N_6083);
and U6650 (N_6650,N_6150,N_6458);
nand U6651 (N_6651,N_6378,N_6167);
nand U6652 (N_6652,N_6292,N_6080);
nand U6653 (N_6653,N_6184,N_6368);
or U6654 (N_6654,N_6452,N_6180);
nand U6655 (N_6655,N_6347,N_6487);
and U6656 (N_6656,N_6142,N_6163);
nor U6657 (N_6657,N_6109,N_6043);
or U6658 (N_6658,N_6015,N_6029);
nand U6659 (N_6659,N_6207,N_6073);
nand U6660 (N_6660,N_6093,N_6156);
nor U6661 (N_6661,N_6268,N_6369);
and U6662 (N_6662,N_6337,N_6212);
xnor U6663 (N_6663,N_6036,N_6024);
and U6664 (N_6664,N_6265,N_6136);
and U6665 (N_6665,N_6305,N_6336);
nor U6666 (N_6666,N_6146,N_6034);
nor U6667 (N_6667,N_6300,N_6169);
nor U6668 (N_6668,N_6349,N_6303);
nand U6669 (N_6669,N_6058,N_6251);
and U6670 (N_6670,N_6226,N_6492);
and U6671 (N_6671,N_6438,N_6346);
or U6672 (N_6672,N_6485,N_6132);
nor U6673 (N_6673,N_6399,N_6238);
and U6674 (N_6674,N_6008,N_6168);
and U6675 (N_6675,N_6055,N_6059);
and U6676 (N_6676,N_6360,N_6153);
and U6677 (N_6677,N_6318,N_6011);
and U6678 (N_6678,N_6096,N_6089);
or U6679 (N_6679,N_6205,N_6214);
and U6680 (N_6680,N_6471,N_6293);
or U6681 (N_6681,N_6174,N_6309);
nor U6682 (N_6682,N_6315,N_6087);
xor U6683 (N_6683,N_6307,N_6120);
nor U6684 (N_6684,N_6101,N_6048);
and U6685 (N_6685,N_6477,N_6204);
or U6686 (N_6686,N_6462,N_6453);
nand U6687 (N_6687,N_6160,N_6402);
or U6688 (N_6688,N_6070,N_6295);
or U6689 (N_6689,N_6145,N_6322);
or U6690 (N_6690,N_6227,N_6443);
or U6691 (N_6691,N_6185,N_6157);
nand U6692 (N_6692,N_6257,N_6465);
and U6693 (N_6693,N_6417,N_6419);
nand U6694 (N_6694,N_6499,N_6134);
nor U6695 (N_6695,N_6490,N_6200);
and U6696 (N_6696,N_6006,N_6288);
and U6697 (N_6697,N_6407,N_6441);
and U6698 (N_6698,N_6192,N_6357);
or U6699 (N_6699,N_6179,N_6270);
and U6700 (N_6700,N_6316,N_6273);
or U6701 (N_6701,N_6488,N_6107);
and U6702 (N_6702,N_6030,N_6327);
nor U6703 (N_6703,N_6486,N_6199);
nor U6704 (N_6704,N_6063,N_6019);
nand U6705 (N_6705,N_6135,N_6344);
and U6706 (N_6706,N_6242,N_6472);
nor U6707 (N_6707,N_6335,N_6390);
nand U6708 (N_6708,N_6285,N_6294);
nor U6709 (N_6709,N_6258,N_6404);
nand U6710 (N_6710,N_6426,N_6172);
nor U6711 (N_6711,N_6240,N_6262);
or U6712 (N_6712,N_6326,N_6003);
or U6713 (N_6713,N_6290,N_6111);
nand U6714 (N_6714,N_6421,N_6476);
nand U6715 (N_6715,N_6128,N_6216);
nand U6716 (N_6716,N_6385,N_6206);
nor U6717 (N_6717,N_6187,N_6253);
and U6718 (N_6718,N_6191,N_6028);
and U6719 (N_6719,N_6319,N_6046);
nor U6720 (N_6720,N_6129,N_6049);
nor U6721 (N_6721,N_6455,N_6037);
and U6722 (N_6722,N_6106,N_6090);
nand U6723 (N_6723,N_6229,N_6445);
nor U6724 (N_6724,N_6282,N_6221);
xor U6725 (N_6725,N_6311,N_6454);
nor U6726 (N_6726,N_6296,N_6386);
nor U6727 (N_6727,N_6249,N_6248);
nor U6728 (N_6728,N_6099,N_6321);
or U6729 (N_6729,N_6496,N_6365);
or U6730 (N_6730,N_6067,N_6420);
or U6731 (N_6731,N_6165,N_6401);
and U6732 (N_6732,N_6027,N_6161);
or U6733 (N_6733,N_6468,N_6196);
nand U6734 (N_6734,N_6031,N_6044);
nor U6735 (N_6735,N_6220,N_6230);
nor U6736 (N_6736,N_6267,N_6291);
or U6737 (N_6737,N_6405,N_6005);
nand U6738 (N_6738,N_6479,N_6252);
or U6739 (N_6739,N_6459,N_6155);
nand U6740 (N_6740,N_6013,N_6001);
nor U6741 (N_6741,N_6409,N_6026);
or U6742 (N_6742,N_6053,N_6332);
nand U6743 (N_6743,N_6256,N_6203);
or U6744 (N_6744,N_6104,N_6085);
nand U6745 (N_6745,N_6444,N_6213);
and U6746 (N_6746,N_6182,N_6395);
xnor U6747 (N_6747,N_6041,N_6194);
or U6748 (N_6748,N_6375,N_6039);
and U6749 (N_6749,N_6075,N_6151);
and U6750 (N_6750,N_6062,N_6338);
nor U6751 (N_6751,N_6364,N_6033);
nor U6752 (N_6752,N_6133,N_6292);
nand U6753 (N_6753,N_6066,N_6001);
or U6754 (N_6754,N_6436,N_6479);
and U6755 (N_6755,N_6141,N_6227);
nor U6756 (N_6756,N_6038,N_6149);
and U6757 (N_6757,N_6371,N_6402);
nor U6758 (N_6758,N_6323,N_6060);
nand U6759 (N_6759,N_6275,N_6089);
and U6760 (N_6760,N_6338,N_6053);
or U6761 (N_6761,N_6387,N_6006);
nor U6762 (N_6762,N_6462,N_6449);
and U6763 (N_6763,N_6265,N_6231);
nand U6764 (N_6764,N_6013,N_6135);
and U6765 (N_6765,N_6142,N_6478);
xnor U6766 (N_6766,N_6492,N_6014);
or U6767 (N_6767,N_6269,N_6195);
nor U6768 (N_6768,N_6485,N_6431);
or U6769 (N_6769,N_6201,N_6409);
and U6770 (N_6770,N_6117,N_6457);
nand U6771 (N_6771,N_6337,N_6002);
nand U6772 (N_6772,N_6201,N_6324);
nor U6773 (N_6773,N_6139,N_6498);
or U6774 (N_6774,N_6197,N_6407);
nor U6775 (N_6775,N_6403,N_6478);
xor U6776 (N_6776,N_6155,N_6466);
xor U6777 (N_6777,N_6187,N_6026);
and U6778 (N_6778,N_6385,N_6373);
or U6779 (N_6779,N_6412,N_6213);
nor U6780 (N_6780,N_6437,N_6328);
xnor U6781 (N_6781,N_6080,N_6221);
or U6782 (N_6782,N_6190,N_6249);
nand U6783 (N_6783,N_6250,N_6054);
and U6784 (N_6784,N_6389,N_6250);
and U6785 (N_6785,N_6324,N_6448);
or U6786 (N_6786,N_6488,N_6239);
nor U6787 (N_6787,N_6154,N_6471);
xor U6788 (N_6788,N_6423,N_6463);
nand U6789 (N_6789,N_6192,N_6012);
and U6790 (N_6790,N_6467,N_6135);
or U6791 (N_6791,N_6350,N_6255);
nor U6792 (N_6792,N_6083,N_6499);
and U6793 (N_6793,N_6117,N_6009);
or U6794 (N_6794,N_6157,N_6394);
or U6795 (N_6795,N_6461,N_6087);
and U6796 (N_6796,N_6396,N_6163);
nor U6797 (N_6797,N_6269,N_6330);
nor U6798 (N_6798,N_6024,N_6234);
or U6799 (N_6799,N_6421,N_6001);
and U6800 (N_6800,N_6010,N_6495);
nand U6801 (N_6801,N_6137,N_6217);
and U6802 (N_6802,N_6468,N_6270);
and U6803 (N_6803,N_6039,N_6083);
and U6804 (N_6804,N_6028,N_6497);
nor U6805 (N_6805,N_6126,N_6217);
or U6806 (N_6806,N_6385,N_6150);
and U6807 (N_6807,N_6485,N_6418);
or U6808 (N_6808,N_6106,N_6334);
or U6809 (N_6809,N_6468,N_6155);
nand U6810 (N_6810,N_6495,N_6057);
nor U6811 (N_6811,N_6306,N_6273);
or U6812 (N_6812,N_6001,N_6400);
xnor U6813 (N_6813,N_6495,N_6364);
and U6814 (N_6814,N_6068,N_6462);
nor U6815 (N_6815,N_6442,N_6064);
and U6816 (N_6816,N_6201,N_6150);
and U6817 (N_6817,N_6469,N_6436);
nand U6818 (N_6818,N_6436,N_6466);
and U6819 (N_6819,N_6002,N_6136);
xor U6820 (N_6820,N_6227,N_6431);
or U6821 (N_6821,N_6273,N_6385);
nand U6822 (N_6822,N_6442,N_6134);
nor U6823 (N_6823,N_6302,N_6473);
or U6824 (N_6824,N_6485,N_6377);
or U6825 (N_6825,N_6294,N_6362);
nor U6826 (N_6826,N_6140,N_6268);
and U6827 (N_6827,N_6366,N_6466);
xor U6828 (N_6828,N_6094,N_6471);
or U6829 (N_6829,N_6402,N_6223);
or U6830 (N_6830,N_6432,N_6015);
nor U6831 (N_6831,N_6357,N_6277);
nand U6832 (N_6832,N_6400,N_6311);
nor U6833 (N_6833,N_6442,N_6391);
or U6834 (N_6834,N_6387,N_6074);
and U6835 (N_6835,N_6054,N_6271);
or U6836 (N_6836,N_6090,N_6423);
nor U6837 (N_6837,N_6308,N_6218);
nor U6838 (N_6838,N_6064,N_6481);
or U6839 (N_6839,N_6322,N_6470);
xor U6840 (N_6840,N_6100,N_6371);
nor U6841 (N_6841,N_6352,N_6331);
nor U6842 (N_6842,N_6097,N_6145);
or U6843 (N_6843,N_6286,N_6157);
xnor U6844 (N_6844,N_6495,N_6020);
nor U6845 (N_6845,N_6205,N_6051);
and U6846 (N_6846,N_6056,N_6480);
or U6847 (N_6847,N_6246,N_6174);
and U6848 (N_6848,N_6034,N_6229);
nand U6849 (N_6849,N_6192,N_6322);
nand U6850 (N_6850,N_6011,N_6251);
nand U6851 (N_6851,N_6149,N_6480);
or U6852 (N_6852,N_6197,N_6092);
xnor U6853 (N_6853,N_6089,N_6282);
and U6854 (N_6854,N_6135,N_6428);
or U6855 (N_6855,N_6233,N_6133);
nor U6856 (N_6856,N_6439,N_6480);
nor U6857 (N_6857,N_6029,N_6395);
or U6858 (N_6858,N_6048,N_6287);
nand U6859 (N_6859,N_6285,N_6127);
xor U6860 (N_6860,N_6297,N_6354);
nand U6861 (N_6861,N_6217,N_6105);
and U6862 (N_6862,N_6394,N_6226);
and U6863 (N_6863,N_6324,N_6147);
nor U6864 (N_6864,N_6150,N_6243);
xor U6865 (N_6865,N_6054,N_6203);
and U6866 (N_6866,N_6148,N_6326);
nor U6867 (N_6867,N_6030,N_6077);
and U6868 (N_6868,N_6238,N_6226);
or U6869 (N_6869,N_6160,N_6399);
and U6870 (N_6870,N_6193,N_6209);
nand U6871 (N_6871,N_6034,N_6301);
nand U6872 (N_6872,N_6082,N_6216);
nor U6873 (N_6873,N_6391,N_6323);
nor U6874 (N_6874,N_6222,N_6319);
or U6875 (N_6875,N_6074,N_6397);
or U6876 (N_6876,N_6057,N_6178);
or U6877 (N_6877,N_6450,N_6042);
nand U6878 (N_6878,N_6129,N_6295);
nand U6879 (N_6879,N_6057,N_6032);
and U6880 (N_6880,N_6080,N_6122);
xor U6881 (N_6881,N_6381,N_6457);
nand U6882 (N_6882,N_6094,N_6031);
or U6883 (N_6883,N_6432,N_6236);
xor U6884 (N_6884,N_6265,N_6120);
or U6885 (N_6885,N_6214,N_6282);
nor U6886 (N_6886,N_6448,N_6153);
and U6887 (N_6887,N_6240,N_6229);
nand U6888 (N_6888,N_6443,N_6146);
or U6889 (N_6889,N_6015,N_6128);
and U6890 (N_6890,N_6106,N_6354);
or U6891 (N_6891,N_6104,N_6092);
or U6892 (N_6892,N_6257,N_6003);
and U6893 (N_6893,N_6474,N_6473);
or U6894 (N_6894,N_6374,N_6279);
or U6895 (N_6895,N_6420,N_6186);
nand U6896 (N_6896,N_6247,N_6088);
or U6897 (N_6897,N_6448,N_6083);
or U6898 (N_6898,N_6215,N_6133);
and U6899 (N_6899,N_6006,N_6018);
nand U6900 (N_6900,N_6204,N_6150);
and U6901 (N_6901,N_6495,N_6084);
or U6902 (N_6902,N_6464,N_6014);
or U6903 (N_6903,N_6143,N_6433);
nand U6904 (N_6904,N_6247,N_6118);
nand U6905 (N_6905,N_6000,N_6345);
or U6906 (N_6906,N_6177,N_6323);
and U6907 (N_6907,N_6347,N_6479);
xnor U6908 (N_6908,N_6023,N_6124);
nand U6909 (N_6909,N_6303,N_6177);
nand U6910 (N_6910,N_6150,N_6089);
nor U6911 (N_6911,N_6071,N_6393);
or U6912 (N_6912,N_6281,N_6469);
nand U6913 (N_6913,N_6199,N_6416);
nand U6914 (N_6914,N_6229,N_6410);
nor U6915 (N_6915,N_6445,N_6432);
or U6916 (N_6916,N_6300,N_6097);
nor U6917 (N_6917,N_6091,N_6465);
or U6918 (N_6918,N_6390,N_6325);
or U6919 (N_6919,N_6159,N_6486);
nand U6920 (N_6920,N_6489,N_6103);
nand U6921 (N_6921,N_6335,N_6146);
or U6922 (N_6922,N_6090,N_6444);
nand U6923 (N_6923,N_6382,N_6332);
and U6924 (N_6924,N_6025,N_6320);
or U6925 (N_6925,N_6044,N_6410);
and U6926 (N_6926,N_6499,N_6166);
nor U6927 (N_6927,N_6487,N_6163);
and U6928 (N_6928,N_6383,N_6416);
and U6929 (N_6929,N_6474,N_6496);
and U6930 (N_6930,N_6392,N_6389);
nand U6931 (N_6931,N_6440,N_6184);
and U6932 (N_6932,N_6073,N_6155);
xor U6933 (N_6933,N_6123,N_6177);
or U6934 (N_6934,N_6307,N_6325);
or U6935 (N_6935,N_6436,N_6318);
or U6936 (N_6936,N_6051,N_6347);
or U6937 (N_6937,N_6240,N_6052);
nor U6938 (N_6938,N_6101,N_6192);
xor U6939 (N_6939,N_6355,N_6487);
and U6940 (N_6940,N_6399,N_6248);
or U6941 (N_6941,N_6474,N_6200);
and U6942 (N_6942,N_6299,N_6498);
nor U6943 (N_6943,N_6327,N_6421);
xnor U6944 (N_6944,N_6027,N_6249);
and U6945 (N_6945,N_6360,N_6095);
nor U6946 (N_6946,N_6025,N_6120);
xor U6947 (N_6947,N_6397,N_6411);
and U6948 (N_6948,N_6233,N_6466);
nand U6949 (N_6949,N_6410,N_6351);
xnor U6950 (N_6950,N_6320,N_6379);
or U6951 (N_6951,N_6081,N_6207);
or U6952 (N_6952,N_6187,N_6449);
xor U6953 (N_6953,N_6125,N_6371);
nor U6954 (N_6954,N_6403,N_6121);
nor U6955 (N_6955,N_6484,N_6458);
nand U6956 (N_6956,N_6002,N_6463);
and U6957 (N_6957,N_6032,N_6250);
and U6958 (N_6958,N_6033,N_6002);
or U6959 (N_6959,N_6183,N_6269);
or U6960 (N_6960,N_6330,N_6189);
nor U6961 (N_6961,N_6485,N_6235);
nor U6962 (N_6962,N_6149,N_6407);
nor U6963 (N_6963,N_6426,N_6019);
nor U6964 (N_6964,N_6046,N_6369);
nor U6965 (N_6965,N_6402,N_6220);
and U6966 (N_6966,N_6287,N_6210);
and U6967 (N_6967,N_6438,N_6358);
or U6968 (N_6968,N_6173,N_6256);
nor U6969 (N_6969,N_6267,N_6147);
or U6970 (N_6970,N_6282,N_6470);
nor U6971 (N_6971,N_6060,N_6243);
nor U6972 (N_6972,N_6337,N_6137);
nor U6973 (N_6973,N_6233,N_6326);
nand U6974 (N_6974,N_6226,N_6039);
or U6975 (N_6975,N_6361,N_6394);
or U6976 (N_6976,N_6491,N_6150);
nor U6977 (N_6977,N_6049,N_6241);
xnor U6978 (N_6978,N_6131,N_6390);
xnor U6979 (N_6979,N_6222,N_6288);
and U6980 (N_6980,N_6390,N_6098);
nor U6981 (N_6981,N_6218,N_6286);
and U6982 (N_6982,N_6293,N_6461);
xnor U6983 (N_6983,N_6295,N_6448);
or U6984 (N_6984,N_6444,N_6450);
nand U6985 (N_6985,N_6493,N_6059);
nand U6986 (N_6986,N_6003,N_6096);
and U6987 (N_6987,N_6137,N_6196);
and U6988 (N_6988,N_6184,N_6469);
and U6989 (N_6989,N_6347,N_6039);
nor U6990 (N_6990,N_6163,N_6223);
nand U6991 (N_6991,N_6059,N_6373);
nor U6992 (N_6992,N_6328,N_6038);
nor U6993 (N_6993,N_6304,N_6410);
or U6994 (N_6994,N_6412,N_6361);
nor U6995 (N_6995,N_6181,N_6014);
nand U6996 (N_6996,N_6411,N_6349);
nand U6997 (N_6997,N_6002,N_6281);
nor U6998 (N_6998,N_6232,N_6101);
nor U6999 (N_6999,N_6181,N_6311);
or U7000 (N_7000,N_6543,N_6970);
or U7001 (N_7001,N_6894,N_6679);
nand U7002 (N_7002,N_6812,N_6808);
or U7003 (N_7003,N_6503,N_6672);
or U7004 (N_7004,N_6795,N_6599);
or U7005 (N_7005,N_6993,N_6678);
nor U7006 (N_7006,N_6687,N_6942);
and U7007 (N_7007,N_6606,N_6588);
or U7008 (N_7008,N_6851,N_6916);
or U7009 (N_7009,N_6634,N_6883);
xnor U7010 (N_7010,N_6803,N_6936);
or U7011 (N_7011,N_6572,N_6875);
and U7012 (N_7012,N_6922,N_6522);
xor U7013 (N_7013,N_6733,N_6654);
nand U7014 (N_7014,N_6556,N_6537);
and U7015 (N_7015,N_6726,N_6782);
nand U7016 (N_7016,N_6590,N_6771);
nor U7017 (N_7017,N_6956,N_6737);
xor U7018 (N_7018,N_6793,N_6621);
or U7019 (N_7019,N_6960,N_6682);
nor U7020 (N_7020,N_6510,N_6871);
and U7021 (N_7021,N_6714,N_6767);
or U7022 (N_7022,N_6781,N_6809);
nand U7023 (N_7023,N_6536,N_6842);
nor U7024 (N_7024,N_6788,N_6866);
nand U7025 (N_7025,N_6535,N_6520);
nand U7026 (N_7026,N_6806,N_6921);
nor U7027 (N_7027,N_6651,N_6586);
or U7028 (N_7028,N_6691,N_6844);
nand U7029 (N_7029,N_6502,N_6841);
nor U7030 (N_7030,N_6903,N_6675);
nand U7031 (N_7031,N_6709,N_6593);
and U7032 (N_7032,N_6934,N_6619);
nor U7033 (N_7033,N_6995,N_6965);
or U7034 (N_7034,N_6648,N_6967);
nand U7035 (N_7035,N_6741,N_6707);
nor U7036 (N_7036,N_6983,N_6661);
nand U7037 (N_7037,N_6605,N_6591);
or U7038 (N_7038,N_6964,N_6656);
nor U7039 (N_7039,N_6930,N_6768);
nand U7040 (N_7040,N_6602,N_6973);
xnor U7041 (N_7041,N_6607,N_6669);
or U7042 (N_7042,N_6544,N_6953);
nand U7043 (N_7043,N_6533,N_6893);
and U7044 (N_7044,N_6990,N_6972);
nand U7045 (N_7045,N_6631,N_6689);
nand U7046 (N_7046,N_6924,N_6870);
nand U7047 (N_7047,N_6506,N_6914);
nand U7048 (N_7048,N_6928,N_6860);
or U7049 (N_7049,N_6596,N_6571);
nand U7050 (N_7050,N_6783,N_6530);
and U7051 (N_7051,N_6977,N_6697);
and U7052 (N_7052,N_6665,N_6872);
and U7053 (N_7053,N_6550,N_6854);
xor U7054 (N_7054,N_6861,N_6721);
nand U7055 (N_7055,N_6907,N_6579);
nor U7056 (N_7056,N_6974,N_6892);
and U7057 (N_7057,N_6904,N_6948);
xor U7058 (N_7058,N_6749,N_6676);
nand U7059 (N_7059,N_6670,N_6575);
nor U7060 (N_7060,N_6532,N_6864);
nor U7061 (N_7061,N_6702,N_6614);
xor U7062 (N_7062,N_6865,N_6869);
and U7063 (N_7063,N_6819,N_6755);
nor U7064 (N_7064,N_6762,N_6863);
nor U7065 (N_7065,N_6686,N_6896);
xor U7066 (N_7066,N_6719,N_6758);
nand U7067 (N_7067,N_6881,N_6730);
nor U7068 (N_7068,N_6852,N_6925);
or U7069 (N_7069,N_6816,N_6798);
xor U7070 (N_7070,N_6850,N_6565);
xor U7071 (N_7071,N_6640,N_6505);
or U7072 (N_7072,N_6722,N_6708);
xnor U7073 (N_7073,N_6978,N_6577);
and U7074 (N_7074,N_6745,N_6937);
nand U7075 (N_7075,N_6668,N_6932);
nor U7076 (N_7076,N_6703,N_6947);
and U7077 (N_7077,N_6815,N_6763);
and U7078 (N_7078,N_6878,N_6626);
and U7079 (N_7079,N_6601,N_6908);
nor U7080 (N_7080,N_6548,N_6569);
nand U7081 (N_7081,N_6962,N_6777);
or U7082 (N_7082,N_6552,N_6761);
xor U7083 (N_7083,N_6566,N_6994);
nor U7084 (N_7084,N_6635,N_6778);
nand U7085 (N_7085,N_6500,N_6929);
or U7086 (N_7086,N_6873,N_6666);
nand U7087 (N_7087,N_6935,N_6746);
nor U7088 (N_7088,N_6779,N_6647);
and U7089 (N_7089,N_6912,N_6775);
nand U7090 (N_7090,N_6582,N_6840);
and U7091 (N_7091,N_6531,N_6792);
nand U7092 (N_7092,N_6886,N_6825);
nand U7093 (N_7093,N_6658,N_6901);
nand U7094 (N_7094,N_6784,N_6772);
nand U7095 (N_7095,N_6827,N_6734);
and U7096 (N_7096,N_6988,N_6655);
nor U7097 (N_7097,N_6663,N_6646);
nand U7098 (N_7098,N_6701,N_6838);
and U7099 (N_7099,N_6835,N_6639);
and U7100 (N_7100,N_6546,N_6512);
nor U7101 (N_7101,N_6589,N_6727);
nand U7102 (N_7102,N_6905,N_6528);
nor U7103 (N_7103,N_6982,N_6927);
nand U7104 (N_7104,N_6828,N_6857);
or U7105 (N_7105,N_6629,N_6989);
nand U7106 (N_7106,N_6945,N_6644);
and U7107 (N_7107,N_6568,N_6876);
and U7108 (N_7108,N_6943,N_6969);
and U7109 (N_7109,N_6739,N_6829);
nand U7110 (N_7110,N_6616,N_6958);
and U7111 (N_7111,N_6917,N_6823);
nor U7112 (N_7112,N_6564,N_6902);
nand U7113 (N_7113,N_6756,N_6845);
and U7114 (N_7114,N_6799,N_6753);
and U7115 (N_7115,N_6509,N_6592);
xnor U7116 (N_7116,N_6743,N_6551);
nor U7117 (N_7117,N_6627,N_6547);
nor U7118 (N_7118,N_6711,N_6527);
nor U7119 (N_7119,N_6534,N_6765);
nand U7120 (N_7120,N_6740,N_6952);
xnor U7121 (N_7121,N_6773,N_6931);
nand U7122 (N_7122,N_6836,N_6649);
and U7123 (N_7123,N_6523,N_6736);
nand U7124 (N_7124,N_6889,N_6817);
or U7125 (N_7125,N_6738,N_6609);
or U7126 (N_7126,N_6963,N_6822);
nor U7127 (N_7127,N_6662,N_6692);
nand U7128 (N_7128,N_6538,N_6750);
nor U7129 (N_7129,N_6515,N_6660);
nor U7130 (N_7130,N_6624,N_6642);
or U7131 (N_7131,N_6517,N_6723);
or U7132 (N_7132,N_6884,N_6603);
xnor U7133 (N_7133,N_6833,N_6637);
nor U7134 (N_7134,N_6998,N_6744);
nor U7135 (N_7135,N_6712,N_6826);
nor U7136 (N_7136,N_6604,N_6976);
and U7137 (N_7137,N_6862,N_6559);
and U7138 (N_7138,N_6725,N_6879);
or U7139 (N_7139,N_6713,N_6975);
nor U7140 (N_7140,N_6834,N_6843);
nand U7141 (N_7141,N_6717,N_6754);
or U7142 (N_7142,N_6585,N_6807);
and U7143 (N_7143,N_6690,N_6511);
or U7144 (N_7144,N_6521,N_6940);
nor U7145 (N_7145,N_6683,N_6574);
xnor U7146 (N_7146,N_6821,N_6685);
nand U7147 (N_7147,N_6576,N_6797);
or U7148 (N_7148,N_6516,N_6769);
and U7149 (N_7149,N_6818,N_6805);
or U7150 (N_7150,N_6653,N_6785);
and U7151 (N_7151,N_6704,N_6831);
and U7152 (N_7152,N_6919,N_6580);
nor U7153 (N_7153,N_6659,N_6558);
or U7154 (N_7154,N_6729,N_6594);
or U7155 (N_7155,N_6877,N_6747);
and U7156 (N_7156,N_6830,N_6887);
nor U7157 (N_7157,N_6802,N_6780);
and U7158 (N_7158,N_6526,N_6652);
nand U7159 (N_7159,N_6909,N_6951);
or U7160 (N_7160,N_6911,N_6542);
or U7161 (N_7161,N_6600,N_6694);
or U7162 (N_7162,N_6824,N_6959);
nor U7163 (N_7163,N_6667,N_6553);
nor U7164 (N_7164,N_6837,N_6724);
nand U7165 (N_7165,N_6622,N_6849);
or U7166 (N_7166,N_6938,N_6997);
xor U7167 (N_7167,N_6561,N_6581);
and U7168 (N_7168,N_6570,N_6504);
nor U7169 (N_7169,N_6519,N_6996);
or U7170 (N_7170,N_6939,N_6557);
nand U7171 (N_7171,N_6874,N_6587);
and U7172 (N_7172,N_6562,N_6846);
nor U7173 (N_7173,N_6560,N_6966);
and U7174 (N_7174,N_6583,N_6541);
nand U7175 (N_7175,N_6955,N_6992);
and U7176 (N_7176,N_6987,N_6525);
or U7177 (N_7177,N_6698,N_6617);
or U7178 (N_7178,N_6981,N_6820);
nand U7179 (N_7179,N_6567,N_6787);
and U7180 (N_7180,N_6898,N_6748);
nor U7181 (N_7181,N_6984,N_6638);
nand U7182 (N_7182,N_6673,N_6518);
and U7183 (N_7183,N_6684,N_6979);
nor U7184 (N_7184,N_6832,N_6971);
nand U7185 (N_7185,N_6804,N_6732);
and U7186 (N_7186,N_6751,N_6980);
or U7187 (N_7187,N_6913,N_6545);
and U7188 (N_7188,N_6764,N_6664);
and U7189 (N_7189,N_6615,N_6858);
nand U7190 (N_7190,N_6643,N_6611);
or U7191 (N_7191,N_6760,N_6933);
nor U7192 (N_7192,N_6899,N_6618);
and U7193 (N_7193,N_6716,N_6796);
nor U7194 (N_7194,N_6941,N_6645);
xor U7195 (N_7195,N_6529,N_6801);
or U7196 (N_7196,N_6706,N_6735);
nand U7197 (N_7197,N_6794,N_6839);
xor U7198 (N_7198,N_6882,N_6688);
and U7199 (N_7199,N_6915,N_6718);
nand U7200 (N_7200,N_6859,N_6657);
nor U7201 (N_7201,N_6991,N_6891);
nand U7202 (N_7202,N_6856,N_6630);
nor U7203 (N_7203,N_6888,N_6610);
and U7204 (N_7204,N_6623,N_6693);
nand U7205 (N_7205,N_6598,N_6632);
nor U7206 (N_7206,N_6813,N_6855);
nand U7207 (N_7207,N_6923,N_6680);
nor U7208 (N_7208,N_6961,N_6949);
or U7209 (N_7209,N_6696,N_6946);
or U7210 (N_7210,N_6524,N_6906);
nand U7211 (N_7211,N_6514,N_6508);
nor U7212 (N_7212,N_6699,N_6513);
xor U7213 (N_7213,N_6578,N_6895);
or U7214 (N_7214,N_6728,N_6674);
or U7215 (N_7215,N_6926,N_6539);
nor U7216 (N_7216,N_6549,N_6985);
or U7217 (N_7217,N_6540,N_6900);
and U7218 (N_7218,N_6681,N_6742);
and U7219 (N_7219,N_6641,N_6847);
nand U7220 (N_7220,N_6563,N_6880);
nand U7221 (N_7221,N_6636,N_6810);
nand U7222 (N_7222,N_6613,N_6950);
nor U7223 (N_7223,N_6897,N_6731);
xnor U7224 (N_7224,N_6954,N_6885);
nand U7225 (N_7225,N_6650,N_6757);
nor U7226 (N_7226,N_6790,N_6944);
nand U7227 (N_7227,N_6770,N_6612);
nor U7228 (N_7228,N_6766,N_6752);
or U7229 (N_7229,N_6814,N_6867);
nand U7230 (N_7230,N_6811,N_6918);
nand U7231 (N_7231,N_6920,N_6628);
nand U7232 (N_7232,N_6791,N_6868);
nand U7233 (N_7233,N_6705,N_6595);
nand U7234 (N_7234,N_6625,N_6608);
nor U7235 (N_7235,N_6720,N_6620);
nor U7236 (N_7236,N_6848,N_6633);
nor U7237 (N_7237,N_6584,N_6986);
or U7238 (N_7238,N_6789,N_6910);
or U7239 (N_7239,N_6890,N_6700);
or U7240 (N_7240,N_6573,N_6774);
and U7241 (N_7241,N_6715,N_6507);
or U7242 (N_7242,N_6710,N_6776);
and U7243 (N_7243,N_6597,N_6999);
nor U7244 (N_7244,N_6786,N_6555);
and U7245 (N_7245,N_6501,N_6957);
xnor U7246 (N_7246,N_6695,N_6759);
nand U7247 (N_7247,N_6671,N_6853);
nor U7248 (N_7248,N_6554,N_6677);
or U7249 (N_7249,N_6800,N_6968);
nand U7250 (N_7250,N_6547,N_6773);
xor U7251 (N_7251,N_6578,N_6985);
nand U7252 (N_7252,N_6904,N_6637);
nor U7253 (N_7253,N_6545,N_6863);
nand U7254 (N_7254,N_6858,N_6620);
nand U7255 (N_7255,N_6572,N_6534);
xnor U7256 (N_7256,N_6818,N_6542);
nor U7257 (N_7257,N_6857,N_6666);
nor U7258 (N_7258,N_6817,N_6517);
nor U7259 (N_7259,N_6629,N_6650);
and U7260 (N_7260,N_6606,N_6762);
nor U7261 (N_7261,N_6841,N_6726);
or U7262 (N_7262,N_6804,N_6928);
or U7263 (N_7263,N_6967,N_6945);
and U7264 (N_7264,N_6838,N_6648);
or U7265 (N_7265,N_6976,N_6805);
nand U7266 (N_7266,N_6587,N_6707);
nor U7267 (N_7267,N_6631,N_6787);
or U7268 (N_7268,N_6529,N_6778);
and U7269 (N_7269,N_6841,N_6867);
nand U7270 (N_7270,N_6747,N_6613);
xor U7271 (N_7271,N_6716,N_6557);
or U7272 (N_7272,N_6896,N_6986);
xnor U7273 (N_7273,N_6733,N_6689);
nand U7274 (N_7274,N_6628,N_6805);
xnor U7275 (N_7275,N_6762,N_6902);
nor U7276 (N_7276,N_6616,N_6502);
or U7277 (N_7277,N_6842,N_6618);
or U7278 (N_7278,N_6533,N_6636);
and U7279 (N_7279,N_6980,N_6590);
nand U7280 (N_7280,N_6813,N_6959);
or U7281 (N_7281,N_6734,N_6748);
nor U7282 (N_7282,N_6897,N_6634);
or U7283 (N_7283,N_6746,N_6795);
nand U7284 (N_7284,N_6861,N_6972);
or U7285 (N_7285,N_6996,N_6691);
nor U7286 (N_7286,N_6697,N_6648);
xnor U7287 (N_7287,N_6687,N_6776);
xnor U7288 (N_7288,N_6603,N_6546);
and U7289 (N_7289,N_6996,N_6655);
nand U7290 (N_7290,N_6878,N_6744);
nor U7291 (N_7291,N_6604,N_6780);
or U7292 (N_7292,N_6509,N_6525);
or U7293 (N_7293,N_6715,N_6841);
nand U7294 (N_7294,N_6906,N_6875);
or U7295 (N_7295,N_6994,N_6914);
or U7296 (N_7296,N_6809,N_6585);
nor U7297 (N_7297,N_6634,N_6732);
xor U7298 (N_7298,N_6588,N_6769);
nor U7299 (N_7299,N_6977,N_6761);
or U7300 (N_7300,N_6580,N_6547);
and U7301 (N_7301,N_6845,N_6843);
nor U7302 (N_7302,N_6511,N_6555);
nand U7303 (N_7303,N_6875,N_6820);
nor U7304 (N_7304,N_6814,N_6935);
nor U7305 (N_7305,N_6992,N_6737);
or U7306 (N_7306,N_6761,N_6755);
xnor U7307 (N_7307,N_6523,N_6986);
and U7308 (N_7308,N_6783,N_6936);
and U7309 (N_7309,N_6979,N_6830);
or U7310 (N_7310,N_6550,N_6785);
and U7311 (N_7311,N_6599,N_6831);
and U7312 (N_7312,N_6821,N_6842);
nor U7313 (N_7313,N_6813,N_6752);
nand U7314 (N_7314,N_6936,N_6893);
nand U7315 (N_7315,N_6657,N_6662);
or U7316 (N_7316,N_6522,N_6840);
or U7317 (N_7317,N_6599,N_6976);
or U7318 (N_7318,N_6681,N_6602);
nor U7319 (N_7319,N_6957,N_6502);
nand U7320 (N_7320,N_6685,N_6558);
or U7321 (N_7321,N_6720,N_6671);
or U7322 (N_7322,N_6902,N_6655);
nand U7323 (N_7323,N_6946,N_6557);
nand U7324 (N_7324,N_6936,N_6876);
and U7325 (N_7325,N_6977,N_6511);
nand U7326 (N_7326,N_6507,N_6945);
and U7327 (N_7327,N_6634,N_6646);
xnor U7328 (N_7328,N_6624,N_6760);
nand U7329 (N_7329,N_6630,N_6978);
or U7330 (N_7330,N_6681,N_6651);
and U7331 (N_7331,N_6619,N_6682);
nand U7332 (N_7332,N_6635,N_6885);
nand U7333 (N_7333,N_6543,N_6836);
or U7334 (N_7334,N_6588,N_6823);
nand U7335 (N_7335,N_6562,N_6796);
or U7336 (N_7336,N_6521,N_6722);
nor U7337 (N_7337,N_6780,N_6858);
or U7338 (N_7338,N_6941,N_6636);
and U7339 (N_7339,N_6556,N_6885);
and U7340 (N_7340,N_6857,N_6871);
xor U7341 (N_7341,N_6903,N_6522);
and U7342 (N_7342,N_6698,N_6985);
or U7343 (N_7343,N_6881,N_6564);
nand U7344 (N_7344,N_6820,N_6644);
nand U7345 (N_7345,N_6824,N_6626);
or U7346 (N_7346,N_6872,N_6610);
and U7347 (N_7347,N_6530,N_6747);
nor U7348 (N_7348,N_6716,N_6993);
or U7349 (N_7349,N_6788,N_6510);
xor U7350 (N_7350,N_6916,N_6958);
nand U7351 (N_7351,N_6512,N_6632);
or U7352 (N_7352,N_6564,N_6593);
and U7353 (N_7353,N_6948,N_6520);
or U7354 (N_7354,N_6589,N_6652);
nand U7355 (N_7355,N_6872,N_6660);
nand U7356 (N_7356,N_6831,N_6508);
nand U7357 (N_7357,N_6640,N_6888);
and U7358 (N_7358,N_6540,N_6666);
or U7359 (N_7359,N_6665,N_6727);
nor U7360 (N_7360,N_6775,N_6946);
nand U7361 (N_7361,N_6911,N_6533);
and U7362 (N_7362,N_6668,N_6852);
nand U7363 (N_7363,N_6946,N_6992);
nand U7364 (N_7364,N_6572,N_6727);
nand U7365 (N_7365,N_6990,N_6843);
xor U7366 (N_7366,N_6731,N_6687);
and U7367 (N_7367,N_6520,N_6732);
nor U7368 (N_7368,N_6620,N_6599);
nand U7369 (N_7369,N_6669,N_6894);
and U7370 (N_7370,N_6634,N_6942);
or U7371 (N_7371,N_6737,N_6881);
nand U7372 (N_7372,N_6722,N_6852);
nor U7373 (N_7373,N_6974,N_6692);
or U7374 (N_7374,N_6851,N_6539);
and U7375 (N_7375,N_6836,N_6671);
and U7376 (N_7376,N_6736,N_6538);
xor U7377 (N_7377,N_6793,N_6780);
nor U7378 (N_7378,N_6961,N_6765);
nor U7379 (N_7379,N_6617,N_6515);
nand U7380 (N_7380,N_6527,N_6925);
nand U7381 (N_7381,N_6667,N_6803);
nor U7382 (N_7382,N_6961,N_6858);
nor U7383 (N_7383,N_6599,N_6933);
nor U7384 (N_7384,N_6866,N_6893);
and U7385 (N_7385,N_6867,N_6908);
nor U7386 (N_7386,N_6941,N_6715);
nand U7387 (N_7387,N_6632,N_6697);
and U7388 (N_7388,N_6857,N_6709);
nand U7389 (N_7389,N_6623,N_6742);
and U7390 (N_7390,N_6754,N_6804);
nand U7391 (N_7391,N_6828,N_6895);
and U7392 (N_7392,N_6541,N_6768);
nor U7393 (N_7393,N_6619,N_6907);
or U7394 (N_7394,N_6770,N_6703);
and U7395 (N_7395,N_6871,N_6773);
nand U7396 (N_7396,N_6997,N_6527);
and U7397 (N_7397,N_6733,N_6602);
or U7398 (N_7398,N_6500,N_6600);
nor U7399 (N_7399,N_6956,N_6554);
nand U7400 (N_7400,N_6988,N_6901);
nor U7401 (N_7401,N_6907,N_6530);
and U7402 (N_7402,N_6955,N_6530);
and U7403 (N_7403,N_6802,N_6898);
nor U7404 (N_7404,N_6743,N_6696);
or U7405 (N_7405,N_6961,N_6863);
and U7406 (N_7406,N_6779,N_6605);
nand U7407 (N_7407,N_6803,N_6961);
nand U7408 (N_7408,N_6776,N_6855);
or U7409 (N_7409,N_6591,N_6559);
nand U7410 (N_7410,N_6984,N_6507);
nand U7411 (N_7411,N_6720,N_6619);
nor U7412 (N_7412,N_6653,N_6974);
nor U7413 (N_7413,N_6589,N_6621);
or U7414 (N_7414,N_6573,N_6859);
xor U7415 (N_7415,N_6584,N_6533);
xnor U7416 (N_7416,N_6899,N_6729);
nor U7417 (N_7417,N_6907,N_6847);
nand U7418 (N_7418,N_6726,N_6504);
nor U7419 (N_7419,N_6710,N_6898);
and U7420 (N_7420,N_6765,N_6646);
and U7421 (N_7421,N_6721,N_6593);
nor U7422 (N_7422,N_6806,N_6526);
nand U7423 (N_7423,N_6752,N_6891);
nor U7424 (N_7424,N_6591,N_6943);
nand U7425 (N_7425,N_6838,N_6530);
or U7426 (N_7426,N_6789,N_6945);
nor U7427 (N_7427,N_6852,N_6819);
xnor U7428 (N_7428,N_6694,N_6701);
and U7429 (N_7429,N_6709,N_6605);
nand U7430 (N_7430,N_6689,N_6724);
or U7431 (N_7431,N_6598,N_6502);
or U7432 (N_7432,N_6585,N_6959);
and U7433 (N_7433,N_6759,N_6810);
nand U7434 (N_7434,N_6831,N_6699);
nand U7435 (N_7435,N_6976,N_6745);
nor U7436 (N_7436,N_6767,N_6761);
or U7437 (N_7437,N_6769,N_6800);
and U7438 (N_7438,N_6641,N_6958);
xnor U7439 (N_7439,N_6588,N_6672);
and U7440 (N_7440,N_6838,N_6600);
nand U7441 (N_7441,N_6700,N_6949);
nand U7442 (N_7442,N_6890,N_6819);
or U7443 (N_7443,N_6937,N_6829);
and U7444 (N_7444,N_6529,N_6817);
or U7445 (N_7445,N_6766,N_6825);
nor U7446 (N_7446,N_6809,N_6986);
and U7447 (N_7447,N_6622,N_6994);
nor U7448 (N_7448,N_6631,N_6742);
nand U7449 (N_7449,N_6845,N_6684);
or U7450 (N_7450,N_6791,N_6981);
or U7451 (N_7451,N_6800,N_6919);
nand U7452 (N_7452,N_6941,N_6717);
and U7453 (N_7453,N_6921,N_6784);
nor U7454 (N_7454,N_6720,N_6757);
and U7455 (N_7455,N_6667,N_6569);
nand U7456 (N_7456,N_6958,N_6865);
xor U7457 (N_7457,N_6547,N_6855);
nor U7458 (N_7458,N_6970,N_6881);
or U7459 (N_7459,N_6924,N_6842);
nor U7460 (N_7460,N_6856,N_6973);
and U7461 (N_7461,N_6706,N_6640);
xor U7462 (N_7462,N_6692,N_6869);
nor U7463 (N_7463,N_6531,N_6849);
or U7464 (N_7464,N_6992,N_6588);
and U7465 (N_7465,N_6885,N_6558);
nand U7466 (N_7466,N_6742,N_6969);
or U7467 (N_7467,N_6928,N_6775);
nor U7468 (N_7468,N_6625,N_6561);
nand U7469 (N_7469,N_6647,N_6864);
or U7470 (N_7470,N_6894,N_6671);
and U7471 (N_7471,N_6621,N_6961);
nand U7472 (N_7472,N_6954,N_6930);
nor U7473 (N_7473,N_6606,N_6671);
and U7474 (N_7474,N_6874,N_6827);
and U7475 (N_7475,N_6696,N_6613);
xnor U7476 (N_7476,N_6592,N_6573);
nor U7477 (N_7477,N_6931,N_6933);
nor U7478 (N_7478,N_6995,N_6830);
or U7479 (N_7479,N_6909,N_6509);
nor U7480 (N_7480,N_6844,N_6661);
nor U7481 (N_7481,N_6764,N_6981);
nor U7482 (N_7482,N_6767,N_6688);
nand U7483 (N_7483,N_6767,N_6683);
or U7484 (N_7484,N_6964,N_6704);
and U7485 (N_7485,N_6521,N_6639);
or U7486 (N_7486,N_6587,N_6558);
nand U7487 (N_7487,N_6920,N_6869);
and U7488 (N_7488,N_6845,N_6715);
nand U7489 (N_7489,N_6787,N_6940);
and U7490 (N_7490,N_6708,N_6866);
nand U7491 (N_7491,N_6510,N_6834);
and U7492 (N_7492,N_6694,N_6744);
and U7493 (N_7493,N_6594,N_6797);
nor U7494 (N_7494,N_6988,N_6587);
nor U7495 (N_7495,N_6576,N_6919);
nor U7496 (N_7496,N_6864,N_6856);
nand U7497 (N_7497,N_6764,N_6522);
and U7498 (N_7498,N_6507,N_6867);
or U7499 (N_7499,N_6524,N_6855);
and U7500 (N_7500,N_7005,N_7378);
nor U7501 (N_7501,N_7334,N_7263);
nand U7502 (N_7502,N_7440,N_7123);
xor U7503 (N_7503,N_7027,N_7267);
nand U7504 (N_7504,N_7314,N_7326);
nand U7505 (N_7505,N_7327,N_7274);
or U7506 (N_7506,N_7447,N_7370);
and U7507 (N_7507,N_7454,N_7246);
nor U7508 (N_7508,N_7418,N_7490);
and U7509 (N_7509,N_7339,N_7128);
nor U7510 (N_7510,N_7257,N_7036);
and U7511 (N_7511,N_7400,N_7238);
or U7512 (N_7512,N_7129,N_7282);
and U7513 (N_7513,N_7178,N_7059);
and U7514 (N_7514,N_7319,N_7459);
and U7515 (N_7515,N_7316,N_7394);
and U7516 (N_7516,N_7251,N_7083);
nor U7517 (N_7517,N_7439,N_7012);
nand U7518 (N_7518,N_7281,N_7458);
or U7519 (N_7519,N_7265,N_7283);
and U7520 (N_7520,N_7431,N_7289);
xor U7521 (N_7521,N_7402,N_7239);
and U7522 (N_7522,N_7428,N_7323);
xor U7523 (N_7523,N_7397,N_7057);
nand U7524 (N_7524,N_7338,N_7404);
xnor U7525 (N_7525,N_7030,N_7031);
or U7526 (N_7526,N_7214,N_7464);
or U7527 (N_7527,N_7469,N_7117);
nor U7528 (N_7528,N_7416,N_7291);
xnor U7529 (N_7529,N_7032,N_7318);
nand U7530 (N_7530,N_7375,N_7110);
and U7531 (N_7531,N_7357,N_7101);
or U7532 (N_7532,N_7009,N_7181);
and U7533 (N_7533,N_7371,N_7337);
and U7534 (N_7534,N_7149,N_7434);
or U7535 (N_7535,N_7138,N_7301);
nand U7536 (N_7536,N_7443,N_7218);
nor U7537 (N_7537,N_7259,N_7466);
nand U7538 (N_7538,N_7294,N_7461);
nor U7539 (N_7539,N_7079,N_7000);
nand U7540 (N_7540,N_7212,N_7328);
and U7541 (N_7541,N_7037,N_7125);
or U7542 (N_7542,N_7106,N_7237);
or U7543 (N_7543,N_7421,N_7054);
nand U7544 (N_7544,N_7011,N_7107);
or U7545 (N_7545,N_7056,N_7188);
nor U7546 (N_7546,N_7261,N_7279);
or U7547 (N_7547,N_7356,N_7325);
and U7548 (N_7548,N_7115,N_7450);
nor U7549 (N_7549,N_7286,N_7433);
nor U7550 (N_7550,N_7353,N_7432);
xor U7551 (N_7551,N_7304,N_7442);
nor U7552 (N_7552,N_7029,N_7383);
xnor U7553 (N_7553,N_7455,N_7494);
and U7554 (N_7554,N_7228,N_7199);
nor U7555 (N_7555,N_7063,N_7364);
nor U7556 (N_7556,N_7264,N_7345);
and U7557 (N_7557,N_7409,N_7350);
nor U7558 (N_7558,N_7476,N_7217);
nor U7559 (N_7559,N_7120,N_7290);
and U7560 (N_7560,N_7175,N_7422);
and U7561 (N_7561,N_7298,N_7122);
or U7562 (N_7562,N_7483,N_7213);
or U7563 (N_7563,N_7041,N_7025);
and U7564 (N_7564,N_7489,N_7379);
nor U7565 (N_7565,N_7189,N_7474);
xor U7566 (N_7566,N_7380,N_7077);
and U7567 (N_7567,N_7082,N_7358);
nor U7568 (N_7568,N_7448,N_7095);
and U7569 (N_7569,N_7068,N_7141);
xnor U7570 (N_7570,N_7241,N_7209);
nand U7571 (N_7571,N_7423,N_7044);
and U7572 (N_7572,N_7403,N_7463);
nand U7573 (N_7573,N_7162,N_7066);
nand U7574 (N_7574,N_7405,N_7254);
xnor U7575 (N_7575,N_7407,N_7196);
nand U7576 (N_7576,N_7295,N_7485);
nor U7577 (N_7577,N_7352,N_7412);
xor U7578 (N_7578,N_7411,N_7022);
and U7579 (N_7579,N_7406,N_7224);
nand U7580 (N_7580,N_7020,N_7441);
nand U7581 (N_7581,N_7361,N_7024);
nor U7582 (N_7582,N_7486,N_7023);
or U7583 (N_7583,N_7322,N_7135);
nand U7584 (N_7584,N_7437,N_7014);
nor U7585 (N_7585,N_7150,N_7146);
or U7586 (N_7586,N_7250,N_7275);
nand U7587 (N_7587,N_7293,N_7310);
or U7588 (N_7588,N_7258,N_7331);
nor U7589 (N_7589,N_7058,N_7108);
or U7590 (N_7590,N_7091,N_7478);
nand U7591 (N_7591,N_7090,N_7280);
nand U7592 (N_7592,N_7253,N_7396);
nand U7593 (N_7593,N_7419,N_7182);
xnor U7594 (N_7594,N_7157,N_7420);
xor U7595 (N_7595,N_7359,N_7131);
nor U7596 (N_7596,N_7010,N_7200);
nand U7597 (N_7597,N_7152,N_7417);
xor U7598 (N_7598,N_7481,N_7453);
nor U7599 (N_7599,N_7472,N_7477);
nor U7600 (N_7600,N_7343,N_7078);
nor U7601 (N_7601,N_7186,N_7013);
and U7602 (N_7602,N_7121,N_7114);
nand U7603 (N_7603,N_7424,N_7398);
xnor U7604 (N_7604,N_7360,N_7170);
and U7605 (N_7605,N_7071,N_7109);
nand U7606 (N_7606,N_7276,N_7161);
and U7607 (N_7607,N_7086,N_7296);
and U7608 (N_7608,N_7187,N_7127);
and U7609 (N_7609,N_7499,N_7329);
nor U7610 (N_7610,N_7244,N_7202);
and U7611 (N_7611,N_7446,N_7015);
nor U7612 (N_7612,N_7435,N_7302);
and U7613 (N_7613,N_7176,N_7102);
xor U7614 (N_7614,N_7093,N_7387);
nor U7615 (N_7615,N_7094,N_7355);
nor U7616 (N_7616,N_7073,N_7449);
nand U7617 (N_7617,N_7497,N_7206);
and U7618 (N_7618,N_7342,N_7307);
nand U7619 (N_7619,N_7415,N_7132);
nand U7620 (N_7620,N_7116,N_7171);
nor U7621 (N_7621,N_7236,N_7084);
nor U7622 (N_7622,N_7067,N_7235);
and U7623 (N_7623,N_7061,N_7179);
nor U7624 (N_7624,N_7330,N_7300);
nand U7625 (N_7625,N_7347,N_7484);
xnor U7626 (N_7626,N_7185,N_7016);
nor U7627 (N_7627,N_7229,N_7008);
or U7628 (N_7628,N_7388,N_7140);
and U7629 (N_7629,N_7098,N_7065);
and U7630 (N_7630,N_7156,N_7134);
or U7631 (N_7631,N_7018,N_7055);
and U7632 (N_7632,N_7382,N_7111);
xor U7633 (N_7633,N_7426,N_7096);
nand U7634 (N_7634,N_7362,N_7430);
xnor U7635 (N_7635,N_7221,N_7203);
or U7636 (N_7636,N_7321,N_7215);
and U7637 (N_7637,N_7045,N_7351);
nor U7638 (N_7638,N_7306,N_7308);
and U7639 (N_7639,N_7070,N_7451);
nand U7640 (N_7640,N_7220,N_7137);
or U7641 (N_7641,N_7226,N_7470);
or U7642 (N_7642,N_7180,N_7288);
xor U7643 (N_7643,N_7268,N_7104);
xor U7644 (N_7644,N_7482,N_7230);
and U7645 (N_7645,N_7376,N_7245);
nor U7646 (N_7646,N_7467,N_7475);
nor U7647 (N_7647,N_7354,N_7346);
or U7648 (N_7648,N_7194,N_7004);
nand U7649 (N_7649,N_7391,N_7126);
or U7650 (N_7650,N_7208,N_7193);
nand U7651 (N_7651,N_7373,N_7438);
nand U7652 (N_7652,N_7401,N_7197);
or U7653 (N_7653,N_7002,N_7313);
nor U7654 (N_7654,N_7173,N_7191);
or U7655 (N_7655,N_7192,N_7085);
and U7656 (N_7656,N_7174,N_7081);
or U7657 (N_7657,N_7427,N_7160);
nor U7658 (N_7658,N_7366,N_7492);
xnor U7659 (N_7659,N_7163,N_7344);
and U7660 (N_7660,N_7266,N_7075);
and U7661 (N_7661,N_7028,N_7017);
or U7662 (N_7662,N_7100,N_7271);
xor U7663 (N_7663,N_7048,N_7488);
nand U7664 (N_7664,N_7303,N_7205);
or U7665 (N_7665,N_7305,N_7053);
and U7666 (N_7666,N_7183,N_7069);
and U7667 (N_7667,N_7046,N_7113);
nor U7668 (N_7668,N_7247,N_7047);
or U7669 (N_7669,N_7335,N_7076);
or U7670 (N_7670,N_7363,N_7456);
and U7671 (N_7671,N_7277,N_7139);
nor U7672 (N_7672,N_7219,N_7386);
nor U7673 (N_7673,N_7487,N_7042);
xor U7674 (N_7674,N_7414,N_7292);
nor U7675 (N_7675,N_7341,N_7164);
and U7676 (N_7676,N_7260,N_7278);
xor U7677 (N_7677,N_7255,N_7201);
nand U7678 (N_7678,N_7393,N_7166);
nand U7679 (N_7679,N_7195,N_7413);
nand U7680 (N_7680,N_7001,N_7309);
xnor U7681 (N_7681,N_7033,N_7092);
and U7682 (N_7682,N_7311,N_7172);
nor U7683 (N_7683,N_7143,N_7367);
xor U7684 (N_7684,N_7495,N_7198);
and U7685 (N_7685,N_7231,N_7460);
nand U7686 (N_7686,N_7369,N_7007);
nand U7687 (N_7687,N_7471,N_7064);
and U7688 (N_7688,N_7384,N_7377);
or U7689 (N_7689,N_7177,N_7019);
or U7690 (N_7690,N_7315,N_7491);
or U7691 (N_7691,N_7052,N_7112);
nor U7692 (N_7692,N_7021,N_7269);
or U7693 (N_7693,N_7297,N_7272);
or U7694 (N_7694,N_7154,N_7252);
and U7695 (N_7695,N_7155,N_7262);
nor U7696 (N_7696,N_7299,N_7324);
nand U7697 (N_7697,N_7320,N_7038);
xor U7698 (N_7698,N_7240,N_7003);
nor U7699 (N_7699,N_7284,N_7043);
and U7700 (N_7700,N_7142,N_7144);
and U7701 (N_7701,N_7365,N_7368);
and U7702 (N_7702,N_7099,N_7234);
xnor U7703 (N_7703,N_7072,N_7227);
and U7704 (N_7704,N_7389,N_7381);
or U7705 (N_7705,N_7204,N_7216);
and U7706 (N_7706,N_7232,N_7317);
and U7707 (N_7707,N_7336,N_7452);
and U7708 (N_7708,N_7493,N_7089);
and U7709 (N_7709,N_7410,N_7408);
nand U7710 (N_7710,N_7087,N_7385);
or U7711 (N_7711,N_7153,N_7425);
and U7712 (N_7712,N_7399,N_7145);
and U7713 (N_7713,N_7158,N_7184);
or U7714 (N_7714,N_7374,N_7462);
or U7715 (N_7715,N_7136,N_7233);
and U7716 (N_7716,N_7287,N_7249);
and U7717 (N_7717,N_7256,N_7147);
or U7718 (N_7718,N_7050,N_7285);
xor U7719 (N_7719,N_7034,N_7468);
or U7720 (N_7720,N_7151,N_7480);
nand U7721 (N_7721,N_7390,N_7190);
xnor U7722 (N_7722,N_7496,N_7273);
nor U7723 (N_7723,N_7035,N_7457);
nand U7724 (N_7724,N_7105,N_7348);
nor U7725 (N_7725,N_7159,N_7340);
nand U7726 (N_7726,N_7133,N_7039);
nor U7727 (N_7727,N_7026,N_7207);
nand U7728 (N_7728,N_7080,N_7445);
and U7729 (N_7729,N_7210,N_7242);
nor U7730 (N_7730,N_7270,N_7062);
nor U7731 (N_7731,N_7223,N_7060);
nor U7732 (N_7732,N_7395,N_7006);
nand U7733 (N_7733,N_7498,N_7436);
xnor U7734 (N_7734,N_7312,N_7167);
or U7735 (N_7735,N_7074,N_7465);
or U7736 (N_7736,N_7222,N_7444);
nor U7737 (N_7737,N_7118,N_7168);
and U7738 (N_7738,N_7349,N_7088);
or U7739 (N_7739,N_7473,N_7165);
nor U7740 (N_7740,N_7333,N_7051);
nand U7741 (N_7741,N_7148,N_7211);
or U7742 (N_7742,N_7479,N_7103);
or U7743 (N_7743,N_7429,N_7097);
nand U7744 (N_7744,N_7119,N_7169);
or U7745 (N_7745,N_7225,N_7040);
and U7746 (N_7746,N_7332,N_7049);
nand U7747 (N_7747,N_7130,N_7248);
xor U7748 (N_7748,N_7124,N_7372);
nor U7749 (N_7749,N_7392,N_7243);
and U7750 (N_7750,N_7340,N_7234);
nor U7751 (N_7751,N_7357,N_7139);
and U7752 (N_7752,N_7082,N_7161);
or U7753 (N_7753,N_7039,N_7160);
nand U7754 (N_7754,N_7113,N_7097);
or U7755 (N_7755,N_7448,N_7318);
xnor U7756 (N_7756,N_7054,N_7330);
xnor U7757 (N_7757,N_7318,N_7043);
nor U7758 (N_7758,N_7455,N_7012);
and U7759 (N_7759,N_7080,N_7211);
nor U7760 (N_7760,N_7402,N_7249);
and U7761 (N_7761,N_7249,N_7345);
or U7762 (N_7762,N_7370,N_7143);
and U7763 (N_7763,N_7130,N_7166);
nand U7764 (N_7764,N_7064,N_7309);
nand U7765 (N_7765,N_7300,N_7265);
nand U7766 (N_7766,N_7054,N_7350);
nor U7767 (N_7767,N_7206,N_7075);
nand U7768 (N_7768,N_7330,N_7240);
xor U7769 (N_7769,N_7235,N_7378);
xor U7770 (N_7770,N_7032,N_7356);
xor U7771 (N_7771,N_7220,N_7234);
nand U7772 (N_7772,N_7083,N_7239);
and U7773 (N_7773,N_7063,N_7151);
nor U7774 (N_7774,N_7434,N_7312);
nand U7775 (N_7775,N_7028,N_7114);
xor U7776 (N_7776,N_7077,N_7260);
and U7777 (N_7777,N_7358,N_7205);
nor U7778 (N_7778,N_7360,N_7245);
and U7779 (N_7779,N_7164,N_7385);
and U7780 (N_7780,N_7435,N_7174);
nor U7781 (N_7781,N_7430,N_7304);
and U7782 (N_7782,N_7017,N_7176);
nand U7783 (N_7783,N_7062,N_7416);
or U7784 (N_7784,N_7066,N_7077);
or U7785 (N_7785,N_7200,N_7228);
and U7786 (N_7786,N_7147,N_7033);
and U7787 (N_7787,N_7070,N_7391);
nand U7788 (N_7788,N_7099,N_7457);
or U7789 (N_7789,N_7336,N_7046);
or U7790 (N_7790,N_7350,N_7213);
nor U7791 (N_7791,N_7379,N_7109);
and U7792 (N_7792,N_7424,N_7368);
or U7793 (N_7793,N_7296,N_7294);
and U7794 (N_7794,N_7298,N_7045);
and U7795 (N_7795,N_7077,N_7487);
nor U7796 (N_7796,N_7356,N_7018);
and U7797 (N_7797,N_7250,N_7267);
nand U7798 (N_7798,N_7399,N_7117);
nor U7799 (N_7799,N_7320,N_7401);
nor U7800 (N_7800,N_7077,N_7158);
and U7801 (N_7801,N_7440,N_7417);
nand U7802 (N_7802,N_7442,N_7242);
nand U7803 (N_7803,N_7372,N_7015);
nor U7804 (N_7804,N_7336,N_7059);
nand U7805 (N_7805,N_7376,N_7476);
nand U7806 (N_7806,N_7341,N_7137);
or U7807 (N_7807,N_7041,N_7145);
nor U7808 (N_7808,N_7071,N_7399);
and U7809 (N_7809,N_7331,N_7368);
nand U7810 (N_7810,N_7357,N_7298);
or U7811 (N_7811,N_7469,N_7137);
nor U7812 (N_7812,N_7227,N_7315);
or U7813 (N_7813,N_7477,N_7152);
and U7814 (N_7814,N_7426,N_7395);
and U7815 (N_7815,N_7429,N_7350);
and U7816 (N_7816,N_7392,N_7242);
xnor U7817 (N_7817,N_7083,N_7152);
nand U7818 (N_7818,N_7034,N_7241);
nor U7819 (N_7819,N_7037,N_7067);
or U7820 (N_7820,N_7113,N_7114);
and U7821 (N_7821,N_7184,N_7020);
or U7822 (N_7822,N_7016,N_7171);
nand U7823 (N_7823,N_7349,N_7065);
and U7824 (N_7824,N_7430,N_7480);
or U7825 (N_7825,N_7448,N_7119);
and U7826 (N_7826,N_7284,N_7352);
or U7827 (N_7827,N_7247,N_7111);
or U7828 (N_7828,N_7078,N_7218);
nor U7829 (N_7829,N_7277,N_7245);
and U7830 (N_7830,N_7042,N_7163);
or U7831 (N_7831,N_7476,N_7113);
or U7832 (N_7832,N_7269,N_7422);
nand U7833 (N_7833,N_7075,N_7295);
and U7834 (N_7834,N_7055,N_7155);
xor U7835 (N_7835,N_7247,N_7135);
nand U7836 (N_7836,N_7021,N_7429);
nor U7837 (N_7837,N_7392,N_7311);
or U7838 (N_7838,N_7450,N_7421);
nand U7839 (N_7839,N_7217,N_7287);
nand U7840 (N_7840,N_7363,N_7462);
and U7841 (N_7841,N_7012,N_7434);
xor U7842 (N_7842,N_7103,N_7421);
xnor U7843 (N_7843,N_7243,N_7206);
nand U7844 (N_7844,N_7428,N_7341);
nand U7845 (N_7845,N_7403,N_7113);
nand U7846 (N_7846,N_7445,N_7360);
and U7847 (N_7847,N_7355,N_7166);
and U7848 (N_7848,N_7194,N_7402);
nor U7849 (N_7849,N_7320,N_7452);
and U7850 (N_7850,N_7007,N_7197);
or U7851 (N_7851,N_7278,N_7327);
nand U7852 (N_7852,N_7366,N_7270);
nand U7853 (N_7853,N_7004,N_7369);
or U7854 (N_7854,N_7036,N_7123);
or U7855 (N_7855,N_7442,N_7308);
and U7856 (N_7856,N_7251,N_7091);
xnor U7857 (N_7857,N_7116,N_7414);
nor U7858 (N_7858,N_7239,N_7481);
or U7859 (N_7859,N_7198,N_7461);
and U7860 (N_7860,N_7362,N_7398);
or U7861 (N_7861,N_7088,N_7299);
and U7862 (N_7862,N_7288,N_7381);
nor U7863 (N_7863,N_7351,N_7369);
nand U7864 (N_7864,N_7268,N_7246);
nor U7865 (N_7865,N_7066,N_7160);
nor U7866 (N_7866,N_7250,N_7442);
nand U7867 (N_7867,N_7005,N_7061);
xnor U7868 (N_7868,N_7378,N_7116);
and U7869 (N_7869,N_7190,N_7202);
nor U7870 (N_7870,N_7360,N_7054);
nor U7871 (N_7871,N_7279,N_7175);
and U7872 (N_7872,N_7437,N_7387);
and U7873 (N_7873,N_7221,N_7361);
xor U7874 (N_7874,N_7379,N_7375);
nand U7875 (N_7875,N_7274,N_7326);
nand U7876 (N_7876,N_7336,N_7016);
or U7877 (N_7877,N_7299,N_7456);
xnor U7878 (N_7878,N_7167,N_7289);
nand U7879 (N_7879,N_7444,N_7056);
nor U7880 (N_7880,N_7270,N_7056);
and U7881 (N_7881,N_7233,N_7332);
nor U7882 (N_7882,N_7096,N_7383);
xnor U7883 (N_7883,N_7449,N_7385);
xnor U7884 (N_7884,N_7007,N_7059);
xnor U7885 (N_7885,N_7018,N_7362);
xnor U7886 (N_7886,N_7196,N_7319);
or U7887 (N_7887,N_7381,N_7028);
nor U7888 (N_7888,N_7335,N_7191);
and U7889 (N_7889,N_7209,N_7419);
nand U7890 (N_7890,N_7076,N_7389);
nand U7891 (N_7891,N_7342,N_7231);
and U7892 (N_7892,N_7377,N_7108);
nor U7893 (N_7893,N_7476,N_7150);
nand U7894 (N_7894,N_7275,N_7033);
and U7895 (N_7895,N_7202,N_7139);
and U7896 (N_7896,N_7214,N_7285);
or U7897 (N_7897,N_7052,N_7183);
or U7898 (N_7898,N_7055,N_7032);
nor U7899 (N_7899,N_7000,N_7017);
and U7900 (N_7900,N_7474,N_7454);
nand U7901 (N_7901,N_7171,N_7266);
and U7902 (N_7902,N_7486,N_7401);
or U7903 (N_7903,N_7413,N_7268);
nand U7904 (N_7904,N_7118,N_7194);
and U7905 (N_7905,N_7367,N_7224);
or U7906 (N_7906,N_7068,N_7375);
nor U7907 (N_7907,N_7110,N_7268);
nand U7908 (N_7908,N_7416,N_7016);
and U7909 (N_7909,N_7358,N_7135);
nor U7910 (N_7910,N_7381,N_7215);
nand U7911 (N_7911,N_7386,N_7230);
nand U7912 (N_7912,N_7229,N_7245);
nand U7913 (N_7913,N_7101,N_7088);
nand U7914 (N_7914,N_7416,N_7022);
nor U7915 (N_7915,N_7049,N_7111);
or U7916 (N_7916,N_7399,N_7321);
nand U7917 (N_7917,N_7438,N_7090);
or U7918 (N_7918,N_7288,N_7078);
and U7919 (N_7919,N_7353,N_7234);
and U7920 (N_7920,N_7069,N_7182);
and U7921 (N_7921,N_7301,N_7368);
or U7922 (N_7922,N_7451,N_7286);
nor U7923 (N_7923,N_7366,N_7398);
nor U7924 (N_7924,N_7426,N_7088);
nor U7925 (N_7925,N_7402,N_7216);
nor U7926 (N_7926,N_7408,N_7015);
nand U7927 (N_7927,N_7289,N_7488);
and U7928 (N_7928,N_7375,N_7131);
nand U7929 (N_7929,N_7215,N_7034);
or U7930 (N_7930,N_7213,N_7353);
or U7931 (N_7931,N_7425,N_7486);
and U7932 (N_7932,N_7147,N_7059);
xnor U7933 (N_7933,N_7490,N_7072);
xnor U7934 (N_7934,N_7169,N_7127);
nand U7935 (N_7935,N_7231,N_7309);
nand U7936 (N_7936,N_7353,N_7372);
nand U7937 (N_7937,N_7383,N_7180);
nand U7938 (N_7938,N_7051,N_7124);
xor U7939 (N_7939,N_7075,N_7463);
nand U7940 (N_7940,N_7047,N_7168);
nor U7941 (N_7941,N_7338,N_7263);
and U7942 (N_7942,N_7302,N_7498);
xnor U7943 (N_7943,N_7426,N_7230);
and U7944 (N_7944,N_7278,N_7368);
or U7945 (N_7945,N_7146,N_7017);
nor U7946 (N_7946,N_7090,N_7115);
nand U7947 (N_7947,N_7014,N_7448);
nor U7948 (N_7948,N_7446,N_7112);
or U7949 (N_7949,N_7448,N_7068);
or U7950 (N_7950,N_7323,N_7017);
and U7951 (N_7951,N_7089,N_7446);
nor U7952 (N_7952,N_7217,N_7051);
and U7953 (N_7953,N_7021,N_7451);
or U7954 (N_7954,N_7093,N_7459);
xnor U7955 (N_7955,N_7207,N_7022);
nor U7956 (N_7956,N_7409,N_7001);
or U7957 (N_7957,N_7354,N_7370);
and U7958 (N_7958,N_7418,N_7319);
nand U7959 (N_7959,N_7220,N_7412);
nand U7960 (N_7960,N_7164,N_7264);
and U7961 (N_7961,N_7390,N_7401);
and U7962 (N_7962,N_7343,N_7346);
and U7963 (N_7963,N_7077,N_7022);
nand U7964 (N_7964,N_7356,N_7024);
and U7965 (N_7965,N_7322,N_7393);
xnor U7966 (N_7966,N_7007,N_7101);
and U7967 (N_7967,N_7215,N_7382);
xor U7968 (N_7968,N_7313,N_7270);
nand U7969 (N_7969,N_7265,N_7062);
nor U7970 (N_7970,N_7275,N_7185);
nand U7971 (N_7971,N_7183,N_7272);
or U7972 (N_7972,N_7483,N_7105);
nor U7973 (N_7973,N_7118,N_7086);
nor U7974 (N_7974,N_7455,N_7438);
nand U7975 (N_7975,N_7043,N_7272);
nor U7976 (N_7976,N_7420,N_7489);
nand U7977 (N_7977,N_7322,N_7108);
or U7978 (N_7978,N_7185,N_7239);
xnor U7979 (N_7979,N_7377,N_7405);
nor U7980 (N_7980,N_7220,N_7289);
xnor U7981 (N_7981,N_7095,N_7071);
xnor U7982 (N_7982,N_7493,N_7227);
or U7983 (N_7983,N_7315,N_7355);
nand U7984 (N_7984,N_7363,N_7335);
nand U7985 (N_7985,N_7417,N_7188);
nand U7986 (N_7986,N_7478,N_7123);
nand U7987 (N_7987,N_7350,N_7236);
or U7988 (N_7988,N_7148,N_7230);
nor U7989 (N_7989,N_7077,N_7452);
nand U7990 (N_7990,N_7184,N_7013);
and U7991 (N_7991,N_7198,N_7320);
nand U7992 (N_7992,N_7395,N_7319);
nand U7993 (N_7993,N_7425,N_7220);
xor U7994 (N_7994,N_7098,N_7367);
and U7995 (N_7995,N_7213,N_7153);
nand U7996 (N_7996,N_7263,N_7326);
or U7997 (N_7997,N_7194,N_7352);
or U7998 (N_7998,N_7454,N_7069);
nand U7999 (N_7999,N_7121,N_7331);
and U8000 (N_8000,N_7711,N_7761);
or U8001 (N_8001,N_7743,N_7514);
nand U8002 (N_8002,N_7682,N_7715);
xor U8003 (N_8003,N_7591,N_7609);
nand U8004 (N_8004,N_7832,N_7595);
nor U8005 (N_8005,N_7838,N_7731);
and U8006 (N_8006,N_7974,N_7950);
xor U8007 (N_8007,N_7662,N_7678);
xnor U8008 (N_8008,N_7994,N_7569);
and U8009 (N_8009,N_7740,N_7987);
nor U8010 (N_8010,N_7957,N_7984);
and U8011 (N_8011,N_7566,N_7868);
nor U8012 (N_8012,N_7879,N_7791);
nor U8013 (N_8013,N_7976,N_7862);
nor U8014 (N_8014,N_7802,N_7511);
nand U8015 (N_8015,N_7540,N_7584);
and U8016 (N_8016,N_7773,N_7691);
nand U8017 (N_8017,N_7983,N_7606);
nor U8018 (N_8018,N_7846,N_7982);
nand U8019 (N_8019,N_7783,N_7860);
nor U8020 (N_8020,N_7754,N_7864);
and U8021 (N_8021,N_7794,N_7757);
nor U8022 (N_8022,N_7568,N_7737);
nand U8023 (N_8023,N_7718,N_7594);
or U8024 (N_8024,N_7938,N_7647);
nor U8025 (N_8025,N_7925,N_7643);
or U8026 (N_8026,N_7553,N_7671);
and U8027 (N_8027,N_7534,N_7932);
and U8028 (N_8028,N_7807,N_7755);
xor U8029 (N_8029,N_7923,N_7681);
and U8030 (N_8030,N_7687,N_7922);
or U8031 (N_8031,N_7583,N_7726);
xnor U8032 (N_8032,N_7676,N_7781);
or U8033 (N_8033,N_7702,N_7582);
nand U8034 (N_8034,N_7798,N_7750);
nand U8035 (N_8035,N_7572,N_7762);
nor U8036 (N_8036,N_7694,N_7552);
nand U8037 (N_8037,N_7690,N_7808);
and U8038 (N_8038,N_7632,N_7601);
or U8039 (N_8039,N_7823,N_7809);
or U8040 (N_8040,N_7847,N_7669);
nand U8041 (N_8041,N_7649,N_7544);
nand U8042 (N_8042,N_7622,N_7505);
nand U8043 (N_8043,N_7688,N_7863);
or U8044 (N_8044,N_7810,N_7557);
and U8045 (N_8045,N_7587,N_7875);
and U8046 (N_8046,N_7623,N_7975);
nand U8047 (N_8047,N_7893,N_7927);
nand U8048 (N_8048,N_7999,N_7765);
nor U8049 (N_8049,N_7789,N_7722);
or U8050 (N_8050,N_7924,N_7819);
xor U8051 (N_8051,N_7615,N_7656);
and U8052 (N_8052,N_7861,N_7996);
and U8053 (N_8053,N_7735,N_7536);
or U8054 (N_8054,N_7685,N_7747);
or U8055 (N_8055,N_7971,N_7532);
and U8056 (N_8056,N_7502,N_7659);
and U8057 (N_8057,N_7600,N_7736);
and U8058 (N_8058,N_7903,N_7709);
nor U8059 (N_8059,N_7954,N_7966);
nand U8060 (N_8060,N_7581,N_7633);
nor U8061 (N_8061,N_7817,N_7692);
or U8062 (N_8062,N_7792,N_7695);
and U8063 (N_8063,N_7889,N_7706);
nor U8064 (N_8064,N_7576,N_7666);
and U8065 (N_8065,N_7837,N_7995);
and U8066 (N_8066,N_7946,N_7831);
nor U8067 (N_8067,N_7992,N_7658);
nor U8068 (N_8068,N_7732,N_7652);
or U8069 (N_8069,N_7886,N_7697);
or U8070 (N_8070,N_7790,N_7844);
nor U8071 (N_8071,N_7801,N_7749);
nor U8072 (N_8072,N_7902,N_7962);
and U8073 (N_8073,N_7907,N_7657);
or U8074 (N_8074,N_7890,N_7836);
and U8075 (N_8075,N_7929,N_7805);
nand U8076 (N_8076,N_7812,N_7721);
nand U8077 (N_8077,N_7519,N_7895);
or U8078 (N_8078,N_7931,N_7788);
nor U8079 (N_8079,N_7611,N_7533);
nor U8080 (N_8080,N_7667,N_7851);
nor U8081 (N_8081,N_7934,N_7698);
and U8082 (N_8082,N_7745,N_7703);
nand U8083 (N_8083,N_7592,N_7752);
nor U8084 (N_8084,N_7855,N_7958);
nor U8085 (N_8085,N_7941,N_7727);
nor U8086 (N_8086,N_7642,N_7524);
nor U8087 (N_8087,N_7517,N_7835);
xor U8088 (N_8088,N_7869,N_7908);
nand U8089 (N_8089,N_7942,N_7588);
nor U8090 (N_8090,N_7503,N_7775);
or U8091 (N_8091,N_7604,N_7926);
xnor U8092 (N_8092,N_7822,N_7952);
xor U8093 (N_8093,N_7818,N_7738);
and U8094 (N_8094,N_7677,N_7548);
nand U8095 (N_8095,N_7693,N_7734);
nor U8096 (N_8096,N_7525,N_7526);
or U8097 (N_8097,N_7830,N_7547);
or U8098 (N_8098,N_7625,N_7521);
or U8099 (N_8099,N_7654,N_7631);
or U8100 (N_8100,N_7556,N_7977);
and U8101 (N_8101,N_7898,N_7870);
or U8102 (N_8102,N_7850,N_7651);
nand U8103 (N_8103,N_7779,N_7530);
xnor U8104 (N_8104,N_7575,N_7797);
nand U8105 (N_8105,N_7579,N_7515);
nor U8106 (N_8106,N_7916,N_7833);
nor U8107 (N_8107,N_7713,N_7683);
nand U8108 (N_8108,N_7930,N_7866);
nand U8109 (N_8109,N_7998,N_7626);
nor U8110 (N_8110,N_7959,N_7988);
and U8111 (N_8111,N_7763,N_7554);
nand U8112 (N_8112,N_7500,N_7627);
or U8113 (N_8113,N_7586,N_7674);
or U8114 (N_8114,N_7598,N_7529);
or U8115 (N_8115,N_7741,N_7558);
or U8116 (N_8116,N_7768,N_7904);
and U8117 (N_8117,N_7605,N_7778);
xnor U8118 (N_8118,N_7561,N_7949);
nand U8119 (N_8119,N_7624,N_7664);
and U8120 (N_8120,N_7522,N_7767);
xnor U8121 (N_8121,N_7739,N_7744);
xor U8122 (N_8122,N_7776,N_7764);
and U8123 (N_8123,N_7665,N_7986);
nand U8124 (N_8124,N_7585,N_7513);
or U8125 (N_8125,N_7634,N_7700);
or U8126 (N_8126,N_7896,N_7843);
nor U8127 (N_8127,N_7969,N_7888);
nand U8128 (N_8128,N_7759,N_7640);
nor U8129 (N_8129,N_7684,N_7840);
nand U8130 (N_8130,N_7965,N_7638);
nand U8131 (N_8131,N_7567,N_7865);
nand U8132 (N_8132,N_7804,N_7614);
xor U8133 (N_8133,N_7824,N_7539);
or U8134 (N_8134,N_7825,N_7639);
and U8135 (N_8135,N_7646,N_7520);
nor U8136 (N_8136,N_7915,N_7672);
xor U8137 (N_8137,N_7828,N_7508);
or U8138 (N_8138,N_7859,N_7748);
nor U8139 (N_8139,N_7590,N_7901);
nor U8140 (N_8140,N_7589,N_7644);
and U8141 (N_8141,N_7725,N_7538);
nand U8142 (N_8142,N_7786,N_7689);
nand U8143 (N_8143,N_7947,N_7680);
nand U8144 (N_8144,N_7973,N_7616);
nor U8145 (N_8145,N_7542,N_7723);
or U8146 (N_8146,N_7991,N_7774);
and U8147 (N_8147,N_7512,N_7653);
and U8148 (N_8148,N_7619,N_7968);
nor U8149 (N_8149,N_7636,N_7661);
nor U8150 (N_8150,N_7796,N_7724);
nand U8151 (N_8151,N_7820,N_7728);
and U8152 (N_8152,N_7849,N_7704);
and U8153 (N_8153,N_7880,N_7777);
and U8154 (N_8154,N_7878,N_7963);
nor U8155 (N_8155,N_7876,N_7937);
nand U8156 (N_8156,N_7979,N_7793);
or U8157 (N_8157,N_7760,N_7771);
nand U8158 (N_8158,N_7766,N_7673);
nor U8159 (N_8159,N_7772,N_7785);
or U8160 (N_8160,N_7603,N_7943);
nand U8161 (N_8161,N_7507,N_7972);
nor U8162 (N_8162,N_7892,N_7528);
or U8163 (N_8163,N_7596,N_7918);
nor U8164 (N_8164,N_7509,N_7978);
nand U8165 (N_8165,N_7546,N_7686);
and U8166 (N_8166,N_7821,N_7746);
xor U8167 (N_8167,N_7857,N_7910);
and U8168 (N_8168,N_7537,N_7990);
or U8169 (N_8169,N_7919,N_7853);
nand U8170 (N_8170,N_7602,N_7914);
and U8171 (N_8171,N_7571,N_7826);
nand U8172 (N_8172,N_7628,N_7608);
nor U8173 (N_8173,N_7897,N_7989);
xnor U8174 (N_8174,N_7578,N_7795);
nor U8175 (N_8175,N_7560,N_7610);
or U8176 (N_8176,N_7940,N_7559);
nor U8177 (N_8177,N_7629,N_7985);
or U8178 (N_8178,N_7708,N_7518);
and U8179 (N_8179,N_7716,N_7541);
nand U8180 (N_8180,N_7531,N_7617);
and U8181 (N_8181,N_7710,N_7580);
nand U8182 (N_8182,N_7881,N_7645);
nand U8183 (N_8183,N_7911,N_7980);
nand U8184 (N_8184,N_7648,N_7970);
nor U8185 (N_8185,N_7663,N_7501);
nand U8186 (N_8186,N_7555,N_7574);
and U8187 (N_8187,N_7597,N_7770);
nand U8188 (N_8188,N_7769,N_7900);
or U8189 (N_8189,N_7856,N_7806);
or U8190 (N_8190,N_7635,N_7696);
and U8191 (N_8191,N_7811,N_7917);
xnor U8192 (N_8192,N_7780,N_7621);
nand U8193 (N_8193,N_7936,N_7733);
xor U8194 (N_8194,N_7852,N_7799);
or U8195 (N_8195,N_7637,N_7841);
and U8196 (N_8196,N_7874,N_7871);
nor U8197 (N_8197,N_7858,N_7510);
and U8198 (N_8198,N_7742,N_7867);
xnor U8199 (N_8199,N_7803,N_7593);
xnor U8200 (N_8200,N_7877,N_7712);
or U8201 (N_8201,N_7670,N_7504);
and U8202 (N_8202,N_7707,N_7549);
nor U8203 (N_8203,N_7933,N_7730);
nand U8204 (N_8204,N_7939,N_7756);
nor U8205 (N_8205,N_7815,N_7787);
nand U8206 (N_8206,N_7945,N_7920);
and U8207 (N_8207,N_7891,N_7618);
nor U8208 (N_8208,N_7599,N_7527);
nor U8209 (N_8209,N_7535,N_7827);
nand U8210 (N_8210,N_7607,N_7997);
and U8211 (N_8211,N_7935,N_7854);
or U8212 (N_8212,N_7679,N_7570);
and U8213 (N_8213,N_7956,N_7506);
nor U8214 (N_8214,N_7758,N_7829);
nand U8215 (N_8215,N_7675,N_7620);
or U8216 (N_8216,N_7650,N_7848);
or U8217 (N_8217,N_7885,N_7953);
nand U8218 (N_8218,N_7955,N_7613);
and U8219 (N_8219,N_7928,N_7701);
or U8220 (N_8220,N_7612,N_7839);
and U8221 (N_8221,N_7550,N_7577);
xor U8222 (N_8222,N_7563,N_7719);
nand U8223 (N_8223,N_7814,N_7717);
nand U8224 (N_8224,N_7960,N_7699);
and U8225 (N_8225,N_7887,N_7714);
nand U8226 (N_8226,N_7884,N_7630);
or U8227 (N_8227,N_7545,N_7641);
nor U8228 (N_8228,N_7834,N_7912);
nor U8229 (N_8229,N_7816,N_7845);
xor U8230 (N_8230,N_7967,N_7981);
or U8231 (N_8231,N_7894,N_7562);
and U8232 (N_8232,N_7705,N_7899);
xor U8233 (N_8233,N_7913,N_7753);
nor U8234 (N_8234,N_7964,N_7784);
nand U8235 (N_8235,N_7944,N_7951);
nor U8236 (N_8236,N_7961,N_7872);
or U8237 (N_8237,N_7993,N_7782);
and U8238 (N_8238,N_7573,N_7660);
and U8239 (N_8239,N_7873,N_7564);
nor U8240 (N_8240,N_7883,N_7921);
nor U8241 (N_8241,N_7729,N_7906);
nand U8242 (N_8242,N_7813,N_7948);
nand U8243 (N_8243,N_7668,N_7523);
nor U8244 (N_8244,N_7543,N_7800);
and U8245 (N_8245,N_7655,N_7882);
nor U8246 (N_8246,N_7905,N_7842);
nand U8247 (N_8247,N_7720,N_7565);
nor U8248 (N_8248,N_7751,N_7909);
nand U8249 (N_8249,N_7551,N_7516);
nand U8250 (N_8250,N_7803,N_7670);
nor U8251 (N_8251,N_7593,N_7941);
and U8252 (N_8252,N_7519,N_7957);
and U8253 (N_8253,N_7554,N_7510);
nor U8254 (N_8254,N_7636,N_7939);
nor U8255 (N_8255,N_7732,N_7687);
or U8256 (N_8256,N_7591,N_7639);
or U8257 (N_8257,N_7887,N_7754);
nand U8258 (N_8258,N_7860,N_7949);
nor U8259 (N_8259,N_7854,N_7962);
and U8260 (N_8260,N_7513,N_7508);
and U8261 (N_8261,N_7615,N_7962);
nand U8262 (N_8262,N_7536,N_7910);
or U8263 (N_8263,N_7835,N_7857);
nand U8264 (N_8264,N_7513,N_7769);
and U8265 (N_8265,N_7920,N_7510);
or U8266 (N_8266,N_7586,N_7813);
or U8267 (N_8267,N_7769,N_7715);
and U8268 (N_8268,N_7803,N_7861);
nand U8269 (N_8269,N_7973,N_7599);
or U8270 (N_8270,N_7801,N_7728);
nand U8271 (N_8271,N_7985,N_7737);
xnor U8272 (N_8272,N_7740,N_7578);
or U8273 (N_8273,N_7728,N_7635);
nor U8274 (N_8274,N_7583,N_7571);
xor U8275 (N_8275,N_7905,N_7724);
nand U8276 (N_8276,N_7810,N_7759);
nand U8277 (N_8277,N_7809,N_7691);
nand U8278 (N_8278,N_7648,N_7642);
or U8279 (N_8279,N_7753,N_7580);
or U8280 (N_8280,N_7604,N_7987);
nand U8281 (N_8281,N_7566,N_7854);
or U8282 (N_8282,N_7545,N_7659);
or U8283 (N_8283,N_7979,N_7781);
xor U8284 (N_8284,N_7692,N_7915);
or U8285 (N_8285,N_7752,N_7870);
or U8286 (N_8286,N_7951,N_7594);
nor U8287 (N_8287,N_7781,N_7912);
xor U8288 (N_8288,N_7826,N_7672);
and U8289 (N_8289,N_7545,N_7899);
or U8290 (N_8290,N_7887,N_7581);
or U8291 (N_8291,N_7802,N_7527);
nand U8292 (N_8292,N_7782,N_7627);
xnor U8293 (N_8293,N_7953,N_7731);
nor U8294 (N_8294,N_7655,N_7633);
nand U8295 (N_8295,N_7506,N_7607);
nand U8296 (N_8296,N_7949,N_7848);
nand U8297 (N_8297,N_7787,N_7641);
xor U8298 (N_8298,N_7741,N_7735);
and U8299 (N_8299,N_7854,N_7781);
nand U8300 (N_8300,N_7804,N_7548);
nor U8301 (N_8301,N_7813,N_7872);
nor U8302 (N_8302,N_7961,N_7533);
xnor U8303 (N_8303,N_7664,N_7936);
nand U8304 (N_8304,N_7650,N_7503);
or U8305 (N_8305,N_7780,N_7861);
or U8306 (N_8306,N_7854,N_7702);
nand U8307 (N_8307,N_7917,N_7802);
nor U8308 (N_8308,N_7699,N_7917);
nand U8309 (N_8309,N_7620,N_7899);
and U8310 (N_8310,N_7607,N_7956);
and U8311 (N_8311,N_7873,N_7980);
or U8312 (N_8312,N_7676,N_7517);
nand U8313 (N_8313,N_7952,N_7934);
and U8314 (N_8314,N_7562,N_7623);
and U8315 (N_8315,N_7960,N_7834);
and U8316 (N_8316,N_7846,N_7761);
and U8317 (N_8317,N_7689,N_7970);
and U8318 (N_8318,N_7995,N_7663);
and U8319 (N_8319,N_7678,N_7878);
or U8320 (N_8320,N_7635,N_7833);
or U8321 (N_8321,N_7839,N_7714);
nand U8322 (N_8322,N_7612,N_7845);
nor U8323 (N_8323,N_7804,N_7878);
nand U8324 (N_8324,N_7650,N_7877);
nor U8325 (N_8325,N_7617,N_7835);
nand U8326 (N_8326,N_7854,N_7584);
or U8327 (N_8327,N_7853,N_7597);
nor U8328 (N_8328,N_7935,N_7619);
or U8329 (N_8329,N_7602,N_7777);
and U8330 (N_8330,N_7512,N_7994);
xor U8331 (N_8331,N_7851,N_7974);
or U8332 (N_8332,N_7586,N_7593);
and U8333 (N_8333,N_7739,N_7612);
xor U8334 (N_8334,N_7786,N_7764);
nor U8335 (N_8335,N_7970,N_7642);
xor U8336 (N_8336,N_7981,N_7866);
or U8337 (N_8337,N_7543,N_7905);
nand U8338 (N_8338,N_7529,N_7808);
and U8339 (N_8339,N_7540,N_7978);
nand U8340 (N_8340,N_7618,N_7978);
nor U8341 (N_8341,N_7671,N_7748);
xor U8342 (N_8342,N_7630,N_7617);
or U8343 (N_8343,N_7635,N_7982);
and U8344 (N_8344,N_7619,N_7910);
nor U8345 (N_8345,N_7554,N_7506);
and U8346 (N_8346,N_7511,N_7667);
xor U8347 (N_8347,N_7679,N_7810);
or U8348 (N_8348,N_7970,N_7936);
or U8349 (N_8349,N_7900,N_7782);
or U8350 (N_8350,N_7928,N_7865);
xor U8351 (N_8351,N_7969,N_7818);
nand U8352 (N_8352,N_7780,N_7670);
nand U8353 (N_8353,N_7711,N_7588);
and U8354 (N_8354,N_7741,N_7673);
nor U8355 (N_8355,N_7959,N_7586);
or U8356 (N_8356,N_7964,N_7562);
and U8357 (N_8357,N_7728,N_7563);
and U8358 (N_8358,N_7887,N_7935);
nor U8359 (N_8359,N_7947,N_7729);
and U8360 (N_8360,N_7591,N_7919);
nand U8361 (N_8361,N_7949,N_7618);
nor U8362 (N_8362,N_7902,N_7856);
or U8363 (N_8363,N_7595,N_7533);
nand U8364 (N_8364,N_7584,N_7642);
nor U8365 (N_8365,N_7607,N_7612);
nor U8366 (N_8366,N_7581,N_7669);
and U8367 (N_8367,N_7684,N_7614);
or U8368 (N_8368,N_7555,N_7527);
or U8369 (N_8369,N_7557,N_7993);
or U8370 (N_8370,N_7509,N_7608);
nor U8371 (N_8371,N_7749,N_7904);
xnor U8372 (N_8372,N_7744,N_7814);
and U8373 (N_8373,N_7576,N_7916);
or U8374 (N_8374,N_7757,N_7545);
nand U8375 (N_8375,N_7512,N_7584);
and U8376 (N_8376,N_7565,N_7673);
xnor U8377 (N_8377,N_7700,N_7596);
and U8378 (N_8378,N_7827,N_7737);
nor U8379 (N_8379,N_7713,N_7556);
xnor U8380 (N_8380,N_7554,N_7935);
and U8381 (N_8381,N_7856,N_7559);
xnor U8382 (N_8382,N_7536,N_7805);
nor U8383 (N_8383,N_7541,N_7927);
and U8384 (N_8384,N_7523,N_7990);
nor U8385 (N_8385,N_7717,N_7729);
and U8386 (N_8386,N_7787,N_7842);
and U8387 (N_8387,N_7699,N_7805);
and U8388 (N_8388,N_7571,N_7905);
nand U8389 (N_8389,N_7702,N_7548);
or U8390 (N_8390,N_7976,N_7602);
nor U8391 (N_8391,N_7958,N_7933);
nand U8392 (N_8392,N_7940,N_7520);
nand U8393 (N_8393,N_7928,N_7848);
or U8394 (N_8394,N_7894,N_7886);
nor U8395 (N_8395,N_7529,N_7743);
nor U8396 (N_8396,N_7957,N_7747);
and U8397 (N_8397,N_7846,N_7781);
and U8398 (N_8398,N_7624,N_7783);
xnor U8399 (N_8399,N_7503,N_7746);
or U8400 (N_8400,N_7836,N_7972);
or U8401 (N_8401,N_7526,N_7909);
and U8402 (N_8402,N_7821,N_7863);
or U8403 (N_8403,N_7508,N_7746);
and U8404 (N_8404,N_7885,N_7822);
or U8405 (N_8405,N_7506,N_7774);
nand U8406 (N_8406,N_7902,N_7724);
and U8407 (N_8407,N_7757,N_7822);
nand U8408 (N_8408,N_7933,N_7722);
or U8409 (N_8409,N_7763,N_7886);
or U8410 (N_8410,N_7956,N_7719);
and U8411 (N_8411,N_7515,N_7749);
or U8412 (N_8412,N_7583,N_7825);
or U8413 (N_8413,N_7571,N_7837);
nand U8414 (N_8414,N_7765,N_7749);
and U8415 (N_8415,N_7568,N_7791);
nand U8416 (N_8416,N_7542,N_7942);
nor U8417 (N_8417,N_7516,N_7958);
nand U8418 (N_8418,N_7589,N_7718);
or U8419 (N_8419,N_7828,N_7818);
nand U8420 (N_8420,N_7822,N_7967);
or U8421 (N_8421,N_7682,N_7991);
or U8422 (N_8422,N_7744,N_7573);
or U8423 (N_8423,N_7949,N_7682);
nor U8424 (N_8424,N_7726,N_7730);
nand U8425 (N_8425,N_7509,N_7982);
nand U8426 (N_8426,N_7600,N_7907);
and U8427 (N_8427,N_7889,N_7580);
xnor U8428 (N_8428,N_7872,N_7587);
or U8429 (N_8429,N_7826,N_7932);
and U8430 (N_8430,N_7627,N_7653);
nand U8431 (N_8431,N_7695,N_7754);
or U8432 (N_8432,N_7573,N_7803);
nor U8433 (N_8433,N_7780,N_7641);
xnor U8434 (N_8434,N_7733,N_7900);
or U8435 (N_8435,N_7921,N_7810);
nor U8436 (N_8436,N_7904,N_7795);
nor U8437 (N_8437,N_7793,N_7736);
nand U8438 (N_8438,N_7860,N_7673);
nor U8439 (N_8439,N_7830,N_7739);
nand U8440 (N_8440,N_7644,N_7941);
or U8441 (N_8441,N_7759,N_7886);
nand U8442 (N_8442,N_7884,N_7810);
or U8443 (N_8443,N_7931,N_7706);
nand U8444 (N_8444,N_7810,N_7693);
and U8445 (N_8445,N_7995,N_7644);
or U8446 (N_8446,N_7575,N_7727);
nor U8447 (N_8447,N_7655,N_7656);
nor U8448 (N_8448,N_7854,N_7643);
nor U8449 (N_8449,N_7755,N_7788);
or U8450 (N_8450,N_7654,N_7963);
nand U8451 (N_8451,N_7557,N_7712);
nor U8452 (N_8452,N_7879,N_7903);
or U8453 (N_8453,N_7610,N_7905);
nand U8454 (N_8454,N_7953,N_7807);
and U8455 (N_8455,N_7995,N_7714);
nor U8456 (N_8456,N_7784,N_7815);
or U8457 (N_8457,N_7888,N_7934);
nor U8458 (N_8458,N_7703,N_7667);
and U8459 (N_8459,N_7507,N_7649);
xor U8460 (N_8460,N_7697,N_7891);
or U8461 (N_8461,N_7947,N_7818);
nor U8462 (N_8462,N_7834,N_7518);
nor U8463 (N_8463,N_7558,N_7926);
and U8464 (N_8464,N_7723,N_7729);
nand U8465 (N_8465,N_7651,N_7607);
and U8466 (N_8466,N_7910,N_7715);
and U8467 (N_8467,N_7685,N_7593);
and U8468 (N_8468,N_7987,N_7675);
nand U8469 (N_8469,N_7915,N_7846);
nand U8470 (N_8470,N_7749,N_7576);
nand U8471 (N_8471,N_7740,N_7588);
nand U8472 (N_8472,N_7929,N_7831);
nand U8473 (N_8473,N_7988,N_7798);
nand U8474 (N_8474,N_7532,N_7745);
and U8475 (N_8475,N_7802,N_7754);
and U8476 (N_8476,N_7987,N_7788);
nand U8477 (N_8477,N_7568,N_7583);
nor U8478 (N_8478,N_7899,N_7579);
or U8479 (N_8479,N_7513,N_7889);
xor U8480 (N_8480,N_7906,N_7934);
nor U8481 (N_8481,N_7618,N_7530);
nor U8482 (N_8482,N_7707,N_7694);
or U8483 (N_8483,N_7789,N_7636);
and U8484 (N_8484,N_7975,N_7748);
and U8485 (N_8485,N_7831,N_7582);
and U8486 (N_8486,N_7834,N_7666);
nand U8487 (N_8487,N_7904,N_7632);
nor U8488 (N_8488,N_7708,N_7863);
or U8489 (N_8489,N_7922,N_7511);
nor U8490 (N_8490,N_7517,N_7807);
nor U8491 (N_8491,N_7574,N_7599);
or U8492 (N_8492,N_7589,N_7903);
xor U8493 (N_8493,N_7500,N_7676);
nand U8494 (N_8494,N_7642,N_7663);
nand U8495 (N_8495,N_7517,N_7743);
nand U8496 (N_8496,N_7710,N_7551);
nand U8497 (N_8497,N_7724,N_7897);
xor U8498 (N_8498,N_7967,N_7831);
xnor U8499 (N_8499,N_7849,N_7856);
and U8500 (N_8500,N_8293,N_8076);
nand U8501 (N_8501,N_8152,N_8222);
or U8502 (N_8502,N_8396,N_8304);
or U8503 (N_8503,N_8303,N_8103);
nand U8504 (N_8504,N_8278,N_8112);
or U8505 (N_8505,N_8419,N_8043);
nor U8506 (N_8506,N_8484,N_8317);
nand U8507 (N_8507,N_8178,N_8096);
xor U8508 (N_8508,N_8389,N_8149);
nand U8509 (N_8509,N_8124,N_8185);
or U8510 (N_8510,N_8032,N_8054);
nor U8511 (N_8511,N_8061,N_8221);
xor U8512 (N_8512,N_8497,N_8273);
nor U8513 (N_8513,N_8470,N_8340);
and U8514 (N_8514,N_8111,N_8362);
and U8515 (N_8515,N_8064,N_8405);
and U8516 (N_8516,N_8476,N_8066);
and U8517 (N_8517,N_8230,N_8176);
or U8518 (N_8518,N_8164,N_8198);
nand U8519 (N_8519,N_8018,N_8479);
and U8520 (N_8520,N_8426,N_8048);
nor U8521 (N_8521,N_8029,N_8408);
and U8522 (N_8522,N_8363,N_8355);
xor U8523 (N_8523,N_8006,N_8492);
nand U8524 (N_8524,N_8047,N_8243);
and U8525 (N_8525,N_8205,N_8137);
nor U8526 (N_8526,N_8282,N_8014);
or U8527 (N_8527,N_8429,N_8005);
and U8528 (N_8528,N_8296,N_8080);
or U8529 (N_8529,N_8219,N_8294);
nand U8530 (N_8530,N_8465,N_8057);
or U8531 (N_8531,N_8262,N_8068);
and U8532 (N_8532,N_8189,N_8079);
and U8533 (N_8533,N_8069,N_8349);
nand U8534 (N_8534,N_8095,N_8370);
and U8535 (N_8535,N_8000,N_8037);
or U8536 (N_8536,N_8352,N_8194);
or U8537 (N_8537,N_8255,N_8059);
and U8538 (N_8538,N_8093,N_8289);
and U8539 (N_8539,N_8428,N_8377);
and U8540 (N_8540,N_8175,N_8383);
nand U8541 (N_8541,N_8457,N_8224);
or U8542 (N_8542,N_8311,N_8186);
nand U8543 (N_8543,N_8280,N_8259);
or U8544 (N_8544,N_8239,N_8191);
nor U8545 (N_8545,N_8235,N_8078);
nor U8546 (N_8546,N_8237,N_8153);
and U8547 (N_8547,N_8168,N_8467);
and U8548 (N_8548,N_8385,N_8134);
nand U8549 (N_8549,N_8337,N_8441);
nand U8550 (N_8550,N_8107,N_8472);
nor U8551 (N_8551,N_8287,N_8358);
or U8552 (N_8552,N_8379,N_8253);
and U8553 (N_8553,N_8060,N_8240);
or U8554 (N_8554,N_8409,N_8143);
or U8555 (N_8555,N_8117,N_8157);
nor U8556 (N_8556,N_8391,N_8165);
and U8557 (N_8557,N_8114,N_8399);
and U8558 (N_8558,N_8147,N_8090);
or U8559 (N_8559,N_8241,N_8151);
nand U8560 (N_8560,N_8067,N_8110);
nor U8561 (N_8561,N_8142,N_8195);
and U8562 (N_8562,N_8085,N_8390);
nand U8563 (N_8563,N_8460,N_8245);
nor U8564 (N_8564,N_8403,N_8423);
nor U8565 (N_8565,N_8307,N_8169);
nor U8566 (N_8566,N_8021,N_8438);
nand U8567 (N_8567,N_8199,N_8430);
and U8568 (N_8568,N_8174,N_8321);
and U8569 (N_8569,N_8170,N_8433);
and U8570 (N_8570,N_8088,N_8368);
or U8571 (N_8571,N_8313,N_8468);
xnor U8572 (N_8572,N_8388,N_8410);
or U8573 (N_8573,N_8447,N_8402);
nor U8574 (N_8574,N_8083,N_8365);
xor U8575 (N_8575,N_8225,N_8133);
xnor U8576 (N_8576,N_8446,N_8361);
nor U8577 (N_8577,N_8486,N_8444);
nor U8578 (N_8578,N_8236,N_8373);
nand U8579 (N_8579,N_8381,N_8123);
and U8580 (N_8580,N_8306,N_8462);
nand U8581 (N_8581,N_8113,N_8172);
and U8582 (N_8582,N_8004,N_8188);
or U8583 (N_8583,N_8330,N_8250);
xor U8584 (N_8584,N_8351,N_8471);
nand U8585 (N_8585,N_8012,N_8279);
nor U8586 (N_8586,N_8331,N_8469);
or U8587 (N_8587,N_8380,N_8056);
or U8588 (N_8588,N_8285,N_8435);
and U8589 (N_8589,N_8334,N_8382);
nand U8590 (N_8590,N_8495,N_8466);
nor U8591 (N_8591,N_8427,N_8244);
xnor U8592 (N_8592,N_8291,N_8144);
nor U8593 (N_8593,N_8270,N_8415);
xor U8594 (N_8594,N_8378,N_8328);
or U8595 (N_8595,N_8455,N_8106);
nor U8596 (N_8596,N_8452,N_8081);
nand U8597 (N_8597,N_8101,N_8038);
or U8598 (N_8598,N_8338,N_8041);
and U8599 (N_8599,N_8102,N_8173);
or U8600 (N_8600,N_8261,N_8413);
nand U8601 (N_8601,N_8025,N_8442);
nand U8602 (N_8602,N_8275,N_8011);
and U8603 (N_8603,N_8281,N_8420);
and U8604 (N_8604,N_8267,N_8166);
and U8605 (N_8605,N_8336,N_8094);
or U8606 (N_8606,N_8477,N_8109);
nor U8607 (N_8607,N_8013,N_8118);
nand U8608 (N_8608,N_8202,N_8160);
xnor U8609 (N_8609,N_8007,N_8204);
nor U8610 (N_8610,N_8395,N_8009);
nor U8611 (N_8611,N_8269,N_8443);
and U8612 (N_8612,N_8499,N_8295);
and U8613 (N_8613,N_8210,N_8431);
and U8614 (N_8614,N_8422,N_8052);
and U8615 (N_8615,N_8372,N_8264);
or U8616 (N_8616,N_8159,N_8228);
and U8617 (N_8617,N_8329,N_8212);
and U8618 (N_8618,N_8461,N_8036);
nand U8619 (N_8619,N_8300,N_8196);
and U8620 (N_8620,N_8126,N_8322);
and U8621 (N_8621,N_8008,N_8148);
nand U8622 (N_8622,N_8028,N_8324);
and U8623 (N_8623,N_8364,N_8092);
and U8624 (N_8624,N_8254,N_8034);
nor U8625 (N_8625,N_8097,N_8211);
nand U8626 (N_8626,N_8203,N_8376);
nand U8627 (N_8627,N_8463,N_8432);
and U8628 (N_8628,N_8473,N_8354);
and U8629 (N_8629,N_8339,N_8020);
nand U8630 (N_8630,N_8348,N_8100);
xnor U8631 (N_8631,N_8122,N_8017);
nand U8632 (N_8632,N_8158,N_8125);
and U8633 (N_8633,N_8305,N_8485);
or U8634 (N_8634,N_8183,N_8258);
and U8635 (N_8635,N_8360,N_8404);
or U8636 (N_8636,N_8490,N_8286);
or U8637 (N_8637,N_8290,N_8045);
xor U8638 (N_8638,N_8049,N_8177);
or U8639 (N_8639,N_8180,N_8091);
nand U8640 (N_8640,N_8184,N_8042);
nand U8641 (N_8641,N_8016,N_8209);
nand U8642 (N_8642,N_8393,N_8356);
nand U8643 (N_8643,N_8163,N_8242);
xor U8644 (N_8644,N_8026,N_8121);
nor U8645 (N_8645,N_8299,N_8040);
nor U8646 (N_8646,N_8065,N_8496);
nor U8647 (N_8647,N_8150,N_8276);
and U8648 (N_8648,N_8182,N_8077);
or U8649 (N_8649,N_8246,N_8271);
nor U8650 (N_8650,N_8154,N_8437);
and U8651 (N_8651,N_8274,N_8206);
and U8652 (N_8652,N_8074,N_8448);
and U8653 (N_8653,N_8384,N_8314);
and U8654 (N_8654,N_8089,N_8283);
and U8655 (N_8655,N_8488,N_8058);
and U8656 (N_8656,N_8346,N_8141);
or U8657 (N_8657,N_8119,N_8084);
nor U8658 (N_8658,N_8247,N_8353);
nor U8659 (N_8659,N_8421,N_8003);
nand U8660 (N_8660,N_8087,N_8418);
xor U8661 (N_8661,N_8155,N_8335);
or U8662 (N_8662,N_8257,N_8193);
and U8663 (N_8663,N_8001,N_8318);
xor U8664 (N_8664,N_8098,N_8024);
or U8665 (N_8665,N_8398,N_8483);
or U8666 (N_8666,N_8310,N_8138);
and U8667 (N_8667,N_8319,N_8146);
and U8668 (N_8668,N_8343,N_8063);
or U8669 (N_8669,N_8071,N_8450);
nand U8670 (N_8670,N_8464,N_8302);
or U8671 (N_8671,N_8039,N_8207);
or U8672 (N_8672,N_8359,N_8449);
nor U8673 (N_8673,N_8400,N_8115);
nor U8674 (N_8674,N_8369,N_8053);
nor U8675 (N_8675,N_8232,N_8130);
nor U8676 (N_8676,N_8131,N_8375);
or U8677 (N_8677,N_8120,N_8190);
nand U8678 (N_8678,N_8451,N_8344);
and U8679 (N_8679,N_8082,N_8301);
and U8680 (N_8680,N_8325,N_8229);
or U8681 (N_8681,N_8482,N_8105);
and U8682 (N_8682,N_8387,N_8135);
nand U8683 (N_8683,N_8162,N_8347);
nand U8684 (N_8684,N_8374,N_8265);
or U8685 (N_8685,N_8213,N_8217);
nand U8686 (N_8686,N_8425,N_8424);
and U8687 (N_8687,N_8099,N_8249);
or U8688 (N_8688,N_8315,N_8233);
or U8689 (N_8689,N_8487,N_8139);
or U8690 (N_8690,N_8475,N_8341);
and U8691 (N_8691,N_8023,N_8434);
nand U8692 (N_8692,N_8035,N_8214);
xor U8693 (N_8693,N_8238,N_8268);
and U8694 (N_8694,N_8231,N_8104);
nand U8695 (N_8695,N_8031,N_8288);
xor U8696 (N_8696,N_8179,N_8223);
nor U8697 (N_8697,N_8456,N_8350);
nand U8698 (N_8698,N_8292,N_8248);
nor U8699 (N_8699,N_8326,N_8498);
or U8700 (N_8700,N_8072,N_8357);
xor U8701 (N_8701,N_8481,N_8411);
and U8702 (N_8702,N_8386,N_8308);
nor U8703 (N_8703,N_8327,N_8453);
nor U8704 (N_8704,N_8022,N_8073);
and U8705 (N_8705,N_8297,N_8284);
nand U8706 (N_8706,N_8167,N_8251);
and U8707 (N_8707,N_8171,N_8445);
nor U8708 (N_8708,N_8493,N_8200);
nand U8709 (N_8709,N_8256,N_8459);
xor U8710 (N_8710,N_8226,N_8366);
and U8711 (N_8711,N_8128,N_8489);
nand U8712 (N_8712,N_8116,N_8440);
and U8713 (N_8713,N_8046,N_8439);
nor U8714 (N_8714,N_8272,N_8062);
xor U8715 (N_8715,N_8458,N_8320);
or U8716 (N_8716,N_8263,N_8407);
nor U8717 (N_8717,N_8371,N_8136);
nor U8718 (N_8718,N_8491,N_8161);
nor U8719 (N_8719,N_8075,N_8234);
xnor U8720 (N_8720,N_8070,N_8201);
nand U8721 (N_8721,N_8323,N_8252);
and U8722 (N_8722,N_8216,N_8220);
nor U8723 (N_8723,N_8312,N_8394);
and U8724 (N_8724,N_8309,N_8227);
or U8725 (N_8725,N_8454,N_8277);
nor U8726 (N_8726,N_8132,N_8140);
or U8727 (N_8727,N_8345,N_8417);
nor U8728 (N_8728,N_8342,N_8044);
or U8729 (N_8729,N_8406,N_8108);
nand U8730 (N_8730,N_8367,N_8187);
or U8731 (N_8731,N_8478,N_8414);
nand U8732 (N_8732,N_8218,N_8192);
and U8733 (N_8733,N_8019,N_8416);
nor U8734 (N_8734,N_8412,N_8266);
nand U8735 (N_8735,N_8436,N_8260);
nor U8736 (N_8736,N_8332,N_8208);
or U8737 (N_8737,N_8145,N_8392);
nand U8738 (N_8738,N_8127,N_8002);
nand U8739 (N_8739,N_8401,N_8197);
xnor U8740 (N_8740,N_8298,N_8051);
nor U8741 (N_8741,N_8156,N_8215);
xor U8742 (N_8742,N_8316,N_8010);
xor U8743 (N_8743,N_8333,N_8474);
and U8744 (N_8744,N_8086,N_8055);
and U8745 (N_8745,N_8494,N_8397);
nand U8746 (N_8746,N_8015,N_8050);
nand U8747 (N_8747,N_8129,N_8033);
nand U8748 (N_8748,N_8030,N_8181);
nand U8749 (N_8749,N_8480,N_8027);
and U8750 (N_8750,N_8151,N_8158);
nor U8751 (N_8751,N_8145,N_8303);
nand U8752 (N_8752,N_8429,N_8281);
nand U8753 (N_8753,N_8472,N_8238);
and U8754 (N_8754,N_8260,N_8011);
and U8755 (N_8755,N_8142,N_8182);
nor U8756 (N_8756,N_8129,N_8496);
nand U8757 (N_8757,N_8473,N_8336);
and U8758 (N_8758,N_8342,N_8279);
xor U8759 (N_8759,N_8096,N_8242);
nand U8760 (N_8760,N_8366,N_8087);
and U8761 (N_8761,N_8460,N_8263);
nand U8762 (N_8762,N_8441,N_8404);
nor U8763 (N_8763,N_8257,N_8160);
and U8764 (N_8764,N_8157,N_8416);
nand U8765 (N_8765,N_8425,N_8247);
xnor U8766 (N_8766,N_8090,N_8284);
and U8767 (N_8767,N_8372,N_8390);
nand U8768 (N_8768,N_8236,N_8023);
and U8769 (N_8769,N_8191,N_8098);
or U8770 (N_8770,N_8240,N_8387);
xnor U8771 (N_8771,N_8462,N_8415);
or U8772 (N_8772,N_8100,N_8499);
nand U8773 (N_8773,N_8099,N_8167);
nor U8774 (N_8774,N_8385,N_8161);
xor U8775 (N_8775,N_8025,N_8012);
nand U8776 (N_8776,N_8151,N_8005);
nor U8777 (N_8777,N_8408,N_8201);
and U8778 (N_8778,N_8198,N_8314);
nor U8779 (N_8779,N_8011,N_8140);
or U8780 (N_8780,N_8122,N_8146);
or U8781 (N_8781,N_8129,N_8409);
nor U8782 (N_8782,N_8353,N_8212);
or U8783 (N_8783,N_8467,N_8085);
and U8784 (N_8784,N_8444,N_8282);
xnor U8785 (N_8785,N_8421,N_8029);
nor U8786 (N_8786,N_8044,N_8273);
or U8787 (N_8787,N_8135,N_8459);
nand U8788 (N_8788,N_8348,N_8036);
nand U8789 (N_8789,N_8347,N_8039);
nor U8790 (N_8790,N_8104,N_8082);
xor U8791 (N_8791,N_8223,N_8472);
and U8792 (N_8792,N_8027,N_8043);
or U8793 (N_8793,N_8008,N_8336);
or U8794 (N_8794,N_8199,N_8481);
nor U8795 (N_8795,N_8159,N_8498);
and U8796 (N_8796,N_8270,N_8321);
and U8797 (N_8797,N_8449,N_8430);
nor U8798 (N_8798,N_8295,N_8458);
nor U8799 (N_8799,N_8225,N_8430);
nand U8800 (N_8800,N_8394,N_8010);
or U8801 (N_8801,N_8065,N_8075);
or U8802 (N_8802,N_8069,N_8393);
or U8803 (N_8803,N_8475,N_8374);
nor U8804 (N_8804,N_8158,N_8156);
or U8805 (N_8805,N_8410,N_8362);
or U8806 (N_8806,N_8050,N_8217);
and U8807 (N_8807,N_8281,N_8191);
nand U8808 (N_8808,N_8456,N_8460);
nand U8809 (N_8809,N_8428,N_8086);
and U8810 (N_8810,N_8099,N_8215);
and U8811 (N_8811,N_8470,N_8003);
and U8812 (N_8812,N_8048,N_8327);
nor U8813 (N_8813,N_8025,N_8109);
nand U8814 (N_8814,N_8370,N_8170);
nand U8815 (N_8815,N_8261,N_8293);
nor U8816 (N_8816,N_8433,N_8230);
and U8817 (N_8817,N_8198,N_8256);
nand U8818 (N_8818,N_8149,N_8063);
nor U8819 (N_8819,N_8439,N_8137);
nand U8820 (N_8820,N_8115,N_8324);
or U8821 (N_8821,N_8450,N_8356);
nand U8822 (N_8822,N_8472,N_8194);
nor U8823 (N_8823,N_8373,N_8018);
and U8824 (N_8824,N_8138,N_8014);
nor U8825 (N_8825,N_8026,N_8384);
and U8826 (N_8826,N_8308,N_8423);
and U8827 (N_8827,N_8338,N_8049);
and U8828 (N_8828,N_8489,N_8211);
or U8829 (N_8829,N_8320,N_8180);
or U8830 (N_8830,N_8483,N_8186);
or U8831 (N_8831,N_8088,N_8266);
nand U8832 (N_8832,N_8309,N_8488);
nand U8833 (N_8833,N_8448,N_8395);
or U8834 (N_8834,N_8053,N_8486);
nand U8835 (N_8835,N_8162,N_8104);
xor U8836 (N_8836,N_8305,N_8329);
or U8837 (N_8837,N_8022,N_8015);
nor U8838 (N_8838,N_8368,N_8002);
and U8839 (N_8839,N_8106,N_8334);
or U8840 (N_8840,N_8269,N_8084);
nor U8841 (N_8841,N_8129,N_8096);
nand U8842 (N_8842,N_8018,N_8428);
nor U8843 (N_8843,N_8476,N_8266);
nand U8844 (N_8844,N_8383,N_8190);
or U8845 (N_8845,N_8235,N_8145);
and U8846 (N_8846,N_8290,N_8270);
nand U8847 (N_8847,N_8336,N_8449);
and U8848 (N_8848,N_8162,N_8051);
nand U8849 (N_8849,N_8246,N_8461);
xor U8850 (N_8850,N_8406,N_8286);
and U8851 (N_8851,N_8264,N_8137);
and U8852 (N_8852,N_8179,N_8366);
and U8853 (N_8853,N_8122,N_8220);
nand U8854 (N_8854,N_8098,N_8304);
and U8855 (N_8855,N_8157,N_8290);
and U8856 (N_8856,N_8153,N_8373);
and U8857 (N_8857,N_8185,N_8488);
nand U8858 (N_8858,N_8399,N_8313);
xnor U8859 (N_8859,N_8421,N_8488);
or U8860 (N_8860,N_8232,N_8135);
nor U8861 (N_8861,N_8444,N_8012);
or U8862 (N_8862,N_8177,N_8450);
nand U8863 (N_8863,N_8162,N_8389);
and U8864 (N_8864,N_8084,N_8490);
nor U8865 (N_8865,N_8230,N_8040);
xnor U8866 (N_8866,N_8184,N_8203);
and U8867 (N_8867,N_8437,N_8272);
xor U8868 (N_8868,N_8255,N_8063);
or U8869 (N_8869,N_8292,N_8489);
nor U8870 (N_8870,N_8189,N_8416);
xor U8871 (N_8871,N_8256,N_8328);
nand U8872 (N_8872,N_8089,N_8068);
nor U8873 (N_8873,N_8281,N_8023);
nand U8874 (N_8874,N_8147,N_8215);
nor U8875 (N_8875,N_8093,N_8087);
or U8876 (N_8876,N_8115,N_8474);
or U8877 (N_8877,N_8228,N_8348);
nor U8878 (N_8878,N_8072,N_8213);
or U8879 (N_8879,N_8309,N_8276);
or U8880 (N_8880,N_8117,N_8036);
and U8881 (N_8881,N_8204,N_8023);
nand U8882 (N_8882,N_8052,N_8236);
and U8883 (N_8883,N_8049,N_8427);
and U8884 (N_8884,N_8009,N_8129);
and U8885 (N_8885,N_8385,N_8314);
nor U8886 (N_8886,N_8198,N_8202);
xor U8887 (N_8887,N_8372,N_8001);
xnor U8888 (N_8888,N_8240,N_8298);
nand U8889 (N_8889,N_8229,N_8396);
nor U8890 (N_8890,N_8079,N_8495);
nand U8891 (N_8891,N_8414,N_8160);
or U8892 (N_8892,N_8427,N_8324);
nor U8893 (N_8893,N_8022,N_8492);
or U8894 (N_8894,N_8131,N_8064);
nand U8895 (N_8895,N_8047,N_8465);
nor U8896 (N_8896,N_8272,N_8289);
nor U8897 (N_8897,N_8351,N_8307);
nand U8898 (N_8898,N_8178,N_8029);
or U8899 (N_8899,N_8041,N_8389);
nand U8900 (N_8900,N_8181,N_8450);
nor U8901 (N_8901,N_8010,N_8173);
and U8902 (N_8902,N_8023,N_8253);
nand U8903 (N_8903,N_8044,N_8011);
nor U8904 (N_8904,N_8324,N_8316);
nor U8905 (N_8905,N_8487,N_8162);
nor U8906 (N_8906,N_8373,N_8184);
and U8907 (N_8907,N_8342,N_8104);
nand U8908 (N_8908,N_8373,N_8296);
xor U8909 (N_8909,N_8191,N_8393);
or U8910 (N_8910,N_8091,N_8241);
or U8911 (N_8911,N_8065,N_8379);
nand U8912 (N_8912,N_8270,N_8046);
nor U8913 (N_8913,N_8215,N_8072);
and U8914 (N_8914,N_8311,N_8211);
nor U8915 (N_8915,N_8186,N_8354);
and U8916 (N_8916,N_8360,N_8107);
nor U8917 (N_8917,N_8364,N_8022);
nor U8918 (N_8918,N_8336,N_8363);
nor U8919 (N_8919,N_8444,N_8322);
or U8920 (N_8920,N_8387,N_8163);
or U8921 (N_8921,N_8265,N_8102);
nor U8922 (N_8922,N_8347,N_8393);
nor U8923 (N_8923,N_8490,N_8381);
or U8924 (N_8924,N_8337,N_8035);
and U8925 (N_8925,N_8310,N_8315);
nand U8926 (N_8926,N_8309,N_8007);
nor U8927 (N_8927,N_8122,N_8223);
nand U8928 (N_8928,N_8013,N_8404);
nand U8929 (N_8929,N_8176,N_8378);
nor U8930 (N_8930,N_8434,N_8423);
or U8931 (N_8931,N_8377,N_8234);
and U8932 (N_8932,N_8168,N_8246);
and U8933 (N_8933,N_8074,N_8437);
nand U8934 (N_8934,N_8481,N_8499);
or U8935 (N_8935,N_8218,N_8157);
xnor U8936 (N_8936,N_8480,N_8398);
and U8937 (N_8937,N_8114,N_8398);
and U8938 (N_8938,N_8400,N_8352);
nor U8939 (N_8939,N_8137,N_8009);
nor U8940 (N_8940,N_8209,N_8495);
nor U8941 (N_8941,N_8082,N_8057);
nand U8942 (N_8942,N_8056,N_8462);
and U8943 (N_8943,N_8238,N_8098);
or U8944 (N_8944,N_8427,N_8475);
and U8945 (N_8945,N_8112,N_8163);
and U8946 (N_8946,N_8449,N_8478);
or U8947 (N_8947,N_8488,N_8293);
and U8948 (N_8948,N_8322,N_8375);
xor U8949 (N_8949,N_8465,N_8115);
nand U8950 (N_8950,N_8470,N_8084);
or U8951 (N_8951,N_8098,N_8104);
and U8952 (N_8952,N_8443,N_8130);
or U8953 (N_8953,N_8068,N_8416);
nor U8954 (N_8954,N_8434,N_8008);
or U8955 (N_8955,N_8146,N_8447);
xnor U8956 (N_8956,N_8043,N_8351);
xnor U8957 (N_8957,N_8317,N_8075);
nand U8958 (N_8958,N_8074,N_8418);
or U8959 (N_8959,N_8293,N_8379);
xor U8960 (N_8960,N_8267,N_8359);
and U8961 (N_8961,N_8066,N_8071);
and U8962 (N_8962,N_8349,N_8024);
or U8963 (N_8963,N_8040,N_8389);
or U8964 (N_8964,N_8264,N_8198);
nand U8965 (N_8965,N_8102,N_8350);
nand U8966 (N_8966,N_8391,N_8096);
and U8967 (N_8967,N_8190,N_8091);
nand U8968 (N_8968,N_8281,N_8198);
or U8969 (N_8969,N_8021,N_8292);
nand U8970 (N_8970,N_8195,N_8062);
nand U8971 (N_8971,N_8013,N_8040);
and U8972 (N_8972,N_8336,N_8494);
or U8973 (N_8973,N_8152,N_8251);
nor U8974 (N_8974,N_8017,N_8036);
or U8975 (N_8975,N_8257,N_8280);
nor U8976 (N_8976,N_8488,N_8296);
nor U8977 (N_8977,N_8239,N_8378);
nand U8978 (N_8978,N_8185,N_8447);
and U8979 (N_8979,N_8106,N_8028);
nand U8980 (N_8980,N_8079,N_8148);
nand U8981 (N_8981,N_8281,N_8373);
nand U8982 (N_8982,N_8374,N_8246);
nor U8983 (N_8983,N_8336,N_8322);
and U8984 (N_8984,N_8254,N_8320);
nand U8985 (N_8985,N_8035,N_8118);
nand U8986 (N_8986,N_8022,N_8303);
or U8987 (N_8987,N_8432,N_8300);
xor U8988 (N_8988,N_8252,N_8216);
nor U8989 (N_8989,N_8389,N_8278);
nand U8990 (N_8990,N_8021,N_8385);
nor U8991 (N_8991,N_8265,N_8259);
or U8992 (N_8992,N_8384,N_8188);
and U8993 (N_8993,N_8420,N_8345);
nand U8994 (N_8994,N_8344,N_8049);
and U8995 (N_8995,N_8461,N_8327);
nor U8996 (N_8996,N_8354,N_8067);
nor U8997 (N_8997,N_8495,N_8484);
xnor U8998 (N_8998,N_8047,N_8440);
nor U8999 (N_8999,N_8248,N_8314);
xnor U9000 (N_9000,N_8740,N_8503);
xnor U9001 (N_9001,N_8998,N_8607);
nor U9002 (N_9002,N_8839,N_8972);
and U9003 (N_9003,N_8721,N_8679);
or U9004 (N_9004,N_8953,N_8658);
or U9005 (N_9005,N_8927,N_8849);
nand U9006 (N_9006,N_8640,N_8549);
xnor U9007 (N_9007,N_8951,N_8556);
nor U9008 (N_9008,N_8564,N_8862);
nor U9009 (N_9009,N_8642,N_8838);
nor U9010 (N_9010,N_8584,N_8984);
or U9011 (N_9011,N_8594,N_8939);
or U9012 (N_9012,N_8614,N_8821);
or U9013 (N_9013,N_8676,N_8889);
or U9014 (N_9014,N_8778,N_8637);
nand U9015 (N_9015,N_8993,N_8990);
nor U9016 (N_9016,N_8651,N_8965);
nor U9017 (N_9017,N_8937,N_8566);
nand U9018 (N_9018,N_8709,N_8646);
nor U9019 (N_9019,N_8707,N_8923);
nor U9020 (N_9020,N_8970,N_8661);
nor U9021 (N_9021,N_8563,N_8559);
nand U9022 (N_9022,N_8659,N_8660);
nand U9023 (N_9023,N_8963,N_8724);
or U9024 (N_9024,N_8665,N_8797);
nand U9025 (N_9025,N_8766,N_8505);
or U9026 (N_9026,N_8866,N_8688);
or U9027 (N_9027,N_8896,N_8666);
nand U9028 (N_9028,N_8532,N_8996);
nor U9029 (N_9029,N_8576,N_8729);
or U9030 (N_9030,N_8882,N_8753);
or U9031 (N_9031,N_8975,N_8861);
xnor U9032 (N_9032,N_8734,N_8630);
nand U9033 (N_9033,N_8897,N_8940);
and U9034 (N_9034,N_8739,N_8760);
nor U9035 (N_9035,N_8905,N_8535);
nand U9036 (N_9036,N_8746,N_8978);
nand U9037 (N_9037,N_8690,N_8964);
xnor U9038 (N_9038,N_8588,N_8723);
nor U9039 (N_9039,N_8946,N_8592);
nor U9040 (N_9040,N_8852,N_8541);
or U9041 (N_9041,N_8769,N_8921);
nand U9042 (N_9042,N_8836,N_8545);
nand U9043 (N_9043,N_8810,N_8698);
nand U9044 (N_9044,N_8950,N_8622);
xor U9045 (N_9045,N_8969,N_8610);
or U9046 (N_9046,N_8612,N_8677);
or U9047 (N_9047,N_8888,N_8638);
nand U9048 (N_9048,N_8793,N_8593);
xnor U9049 (N_9049,N_8818,N_8992);
or U9050 (N_9050,N_8803,N_8597);
nor U9051 (N_9051,N_8682,N_8931);
and U9052 (N_9052,N_8641,N_8633);
or U9053 (N_9053,N_8546,N_8568);
xnor U9054 (N_9054,N_8554,N_8782);
nor U9055 (N_9055,N_8809,N_8713);
or U9056 (N_9056,N_8892,N_8987);
nor U9057 (N_9057,N_8741,N_8971);
nor U9058 (N_9058,N_8513,N_8579);
and U9059 (N_9059,N_8954,N_8664);
nor U9060 (N_9060,N_8786,N_8916);
nor U9061 (N_9061,N_8502,N_8945);
and U9062 (N_9062,N_8727,N_8865);
and U9063 (N_9063,N_8813,N_8697);
or U9064 (N_9064,N_8742,N_8781);
or U9065 (N_9065,N_8598,N_8764);
and U9066 (N_9066,N_8528,N_8999);
nand U9067 (N_9067,N_8645,N_8805);
nor U9068 (N_9068,N_8705,N_8562);
or U9069 (N_9069,N_8974,N_8920);
or U9070 (N_9070,N_8647,N_8935);
and U9071 (N_9071,N_8850,N_8828);
nand U9072 (N_9072,N_8518,N_8516);
or U9073 (N_9073,N_8620,N_8754);
and U9074 (N_9074,N_8982,N_8871);
nand U9075 (N_9075,N_8745,N_8900);
or U9076 (N_9076,N_8762,N_8807);
nand U9077 (N_9077,N_8913,N_8715);
nor U9078 (N_9078,N_8595,N_8833);
xnor U9079 (N_9079,N_8635,N_8625);
nand U9080 (N_9080,N_8878,N_8581);
nor U9081 (N_9081,N_8524,N_8843);
xnor U9082 (N_9082,N_8684,N_8577);
and U9083 (N_9083,N_8908,N_8624);
xor U9084 (N_9084,N_8874,N_8555);
xnor U9085 (N_9085,N_8605,N_8785);
or U9086 (N_9086,N_8795,N_8752);
and U9087 (N_9087,N_8673,N_8553);
nor U9088 (N_9088,N_8761,N_8501);
or U9089 (N_9089,N_8981,N_8934);
nand U9090 (N_9090,N_8617,N_8509);
nor U9091 (N_9091,N_8791,N_8800);
or U9092 (N_9092,N_8749,N_8979);
nor U9093 (N_9093,N_8648,N_8654);
nand U9094 (N_9094,N_8636,N_8956);
and U9095 (N_9095,N_8922,N_8985);
or U9096 (N_9096,N_8925,N_8575);
and U9097 (N_9097,N_8578,N_8519);
nand U9098 (N_9098,N_8768,N_8567);
and U9099 (N_9099,N_8829,N_8533);
or U9100 (N_9100,N_8655,N_8548);
nor U9101 (N_9101,N_8885,N_8538);
or U9102 (N_9102,N_8626,N_8986);
xnor U9103 (N_9103,N_8991,N_8907);
and U9104 (N_9104,N_8853,N_8710);
nor U9105 (N_9105,N_8904,N_8777);
xnor U9106 (N_9106,N_8687,N_8680);
or U9107 (N_9107,N_8542,N_8873);
nor U9108 (N_9108,N_8789,N_8557);
or U9109 (N_9109,N_8703,N_8717);
and U9110 (N_9110,N_8510,N_8919);
or U9111 (N_9111,N_8759,N_8726);
xor U9112 (N_9112,N_8751,N_8669);
xnor U9113 (N_9113,N_8776,N_8841);
and U9114 (N_9114,N_8737,N_8811);
nand U9115 (N_9115,N_8790,N_8947);
or U9116 (N_9116,N_8653,N_8787);
and U9117 (N_9117,N_8910,N_8846);
and U9118 (N_9118,N_8522,N_8860);
xor U9119 (N_9119,N_8718,N_8961);
or U9120 (N_9120,N_8894,N_8619);
and U9121 (N_9121,N_8539,N_8699);
nand U9122 (N_9122,N_8788,N_8608);
or U9123 (N_9123,N_8891,N_8962);
nor U9124 (N_9124,N_8870,N_8825);
xnor U9125 (N_9125,N_8890,N_8750);
nor U9126 (N_9126,N_8704,N_8570);
xnor U9127 (N_9127,N_8500,N_8526);
and U9128 (N_9128,N_8989,N_8623);
nor U9129 (N_9129,N_8767,N_8708);
nand U9130 (N_9130,N_8755,N_8571);
and U9131 (N_9131,N_8550,N_8822);
and U9132 (N_9132,N_8603,N_8942);
xor U9133 (N_9133,N_8508,N_8720);
nor U9134 (N_9134,N_8820,N_8823);
and U9135 (N_9135,N_8506,N_8618);
nor U9136 (N_9136,N_8774,N_8855);
and U9137 (N_9137,N_8859,N_8649);
nand U9138 (N_9138,N_8872,N_8763);
nor U9139 (N_9139,N_8929,N_8918);
nand U9140 (N_9140,N_8814,N_8558);
nand U9141 (N_9141,N_8585,N_8957);
nand U9142 (N_9142,N_8656,N_8731);
or U9143 (N_9143,N_8650,N_8663);
nor U9144 (N_9144,N_8604,N_8512);
xor U9145 (N_9145,N_8700,N_8844);
xnor U9146 (N_9146,N_8758,N_8840);
nor U9147 (N_9147,N_8531,N_8880);
and U9148 (N_9148,N_8504,N_8914);
and U9149 (N_9149,N_8932,N_8997);
xnor U9150 (N_9150,N_8976,N_8883);
xnor U9151 (N_9151,N_8574,N_8924);
nor U9152 (N_9152,N_8784,N_8815);
and U9153 (N_9153,N_8802,N_8692);
or U9154 (N_9154,N_8955,N_8770);
and U9155 (N_9155,N_8834,N_8599);
xnor U9156 (N_9156,N_8674,N_8507);
and U9157 (N_9157,N_8847,N_8543);
nand U9158 (N_9158,N_8590,N_8517);
xnor U9159 (N_9159,N_8689,N_8845);
or U9160 (N_9160,N_8672,N_8804);
and U9161 (N_9161,N_8792,N_8611);
nor U9162 (N_9162,N_8675,N_8826);
nand U9163 (N_9163,N_8779,N_8701);
xnor U9164 (N_9164,N_8959,N_8725);
or U9165 (N_9165,N_8601,N_8657);
and U9166 (N_9166,N_8893,N_8722);
or U9167 (N_9167,N_8854,N_8816);
xnor U9168 (N_9168,N_8948,N_8941);
nor U9169 (N_9169,N_8521,N_8652);
nor U9170 (N_9170,N_8714,N_8678);
or U9171 (N_9171,N_8552,N_8909);
nor U9172 (N_9172,N_8857,N_8903);
and U9173 (N_9173,N_8711,N_8627);
nand U9174 (N_9174,N_8602,N_8912);
nor U9175 (N_9175,N_8693,N_8628);
xor U9176 (N_9176,N_8799,N_8744);
and U9177 (N_9177,N_8899,N_8728);
nand U9178 (N_9178,N_8917,N_8561);
xnor U9179 (N_9179,N_8851,N_8671);
nand U9180 (N_9180,N_8606,N_8706);
and U9181 (N_9181,N_8743,N_8644);
xnor U9182 (N_9182,N_8968,N_8520);
nor U9183 (N_9183,N_8830,N_8773);
nand U9184 (N_9184,N_8685,N_8668);
xnor U9185 (N_9185,N_8933,N_8936);
nand U9186 (N_9186,N_8629,N_8943);
and U9187 (N_9187,N_8901,N_8949);
nand U9188 (N_9188,N_8796,N_8856);
and U9189 (N_9189,N_8757,N_8858);
and U9190 (N_9190,N_8587,N_8827);
nor U9191 (N_9191,N_8863,N_8591);
or U9192 (N_9192,N_8634,N_8616);
or U9193 (N_9193,N_8613,N_8869);
or U9194 (N_9194,N_8537,N_8832);
and U9195 (N_9195,N_8529,N_8527);
nand U9196 (N_9196,N_8780,N_8876);
or U9197 (N_9197,N_8867,N_8915);
nand U9198 (N_9198,N_8643,N_8632);
nor U9199 (N_9199,N_8596,N_8926);
nor U9200 (N_9200,N_8572,N_8686);
xnor U9201 (N_9201,N_8738,N_8569);
nand U9202 (N_9202,N_8756,N_8967);
nor U9203 (N_9203,N_8938,N_8514);
nand U9204 (N_9204,N_8842,N_8875);
nand U9205 (N_9205,N_8525,N_8702);
and U9206 (N_9206,N_8631,N_8583);
xnor U9207 (N_9207,N_8798,N_8733);
and U9208 (N_9208,N_8817,N_8819);
and U9209 (N_9209,N_8530,N_8952);
nor U9210 (N_9210,N_8973,N_8977);
or U9211 (N_9211,N_8848,N_8864);
xnor U9212 (N_9212,N_8783,N_8540);
nor U9213 (N_9213,N_8609,N_8515);
xor U9214 (N_9214,N_8944,N_8824);
nand U9215 (N_9215,N_8735,N_8831);
xor U9216 (N_9216,N_8868,N_8580);
nor U9217 (N_9217,N_8794,N_8716);
xnor U9218 (N_9218,N_8994,N_8732);
or U9219 (N_9219,N_8534,N_8886);
nor U9220 (N_9220,N_8995,N_8683);
or U9221 (N_9221,N_8730,N_8523);
and U9222 (N_9222,N_8691,N_8887);
and U9223 (N_9223,N_8547,N_8681);
nand U9224 (N_9224,N_8662,N_8667);
and U9225 (N_9225,N_8988,N_8615);
nand U9226 (N_9226,N_8895,N_8736);
or U9227 (N_9227,N_8670,N_8589);
nor U9228 (N_9228,N_8911,N_8775);
and U9229 (N_9229,N_8536,N_8806);
or U9230 (N_9230,N_8696,N_8712);
and U9231 (N_9231,N_8930,N_8808);
nand U9232 (N_9232,N_8582,N_8837);
and U9233 (N_9233,N_8565,N_8586);
nand U9234 (N_9234,N_8748,N_8928);
and U9235 (N_9235,N_8747,N_8771);
and U9236 (N_9236,N_8573,N_8639);
or U9237 (N_9237,N_8621,N_8906);
nand U9238 (N_9238,N_8801,N_8694);
or U9239 (N_9239,N_8879,N_8765);
nand U9240 (N_9240,N_8812,N_8877);
nand U9241 (N_9241,N_8560,N_8983);
or U9242 (N_9242,N_8980,N_8600);
and U9243 (N_9243,N_8898,N_8551);
nand U9244 (N_9244,N_8884,N_8835);
or U9245 (N_9245,N_8695,N_8511);
xnor U9246 (N_9246,N_8544,N_8772);
xnor U9247 (N_9247,N_8881,N_8902);
nand U9248 (N_9248,N_8719,N_8958);
nand U9249 (N_9249,N_8960,N_8966);
nor U9250 (N_9250,N_8842,N_8732);
and U9251 (N_9251,N_8507,N_8837);
or U9252 (N_9252,N_8937,N_8594);
nor U9253 (N_9253,N_8948,N_8737);
and U9254 (N_9254,N_8742,N_8565);
and U9255 (N_9255,N_8747,N_8731);
nor U9256 (N_9256,N_8860,N_8617);
or U9257 (N_9257,N_8955,N_8949);
and U9258 (N_9258,N_8836,N_8620);
and U9259 (N_9259,N_8755,N_8629);
xnor U9260 (N_9260,N_8626,N_8851);
nand U9261 (N_9261,N_8975,N_8686);
nand U9262 (N_9262,N_8903,N_8844);
and U9263 (N_9263,N_8893,N_8691);
or U9264 (N_9264,N_8606,N_8874);
nand U9265 (N_9265,N_8742,N_8779);
and U9266 (N_9266,N_8840,N_8886);
and U9267 (N_9267,N_8812,N_8876);
nand U9268 (N_9268,N_8858,N_8671);
nor U9269 (N_9269,N_8882,N_8746);
or U9270 (N_9270,N_8784,N_8801);
nand U9271 (N_9271,N_8884,N_8557);
and U9272 (N_9272,N_8641,N_8888);
and U9273 (N_9273,N_8602,N_8591);
or U9274 (N_9274,N_8805,N_8981);
nor U9275 (N_9275,N_8886,N_8891);
or U9276 (N_9276,N_8648,N_8795);
nor U9277 (N_9277,N_8951,N_8642);
nand U9278 (N_9278,N_8723,N_8599);
nand U9279 (N_9279,N_8952,N_8733);
nand U9280 (N_9280,N_8746,N_8998);
nor U9281 (N_9281,N_8534,N_8830);
nor U9282 (N_9282,N_8674,N_8776);
nor U9283 (N_9283,N_8965,N_8752);
or U9284 (N_9284,N_8549,N_8888);
xor U9285 (N_9285,N_8845,N_8932);
and U9286 (N_9286,N_8531,N_8615);
and U9287 (N_9287,N_8582,N_8661);
nor U9288 (N_9288,N_8551,N_8672);
or U9289 (N_9289,N_8697,N_8937);
and U9290 (N_9290,N_8545,N_8918);
nor U9291 (N_9291,N_8927,N_8842);
nand U9292 (N_9292,N_8866,N_8613);
nor U9293 (N_9293,N_8994,N_8926);
nand U9294 (N_9294,N_8819,N_8624);
and U9295 (N_9295,N_8786,N_8533);
or U9296 (N_9296,N_8507,N_8688);
nand U9297 (N_9297,N_8606,N_8679);
nor U9298 (N_9298,N_8619,N_8922);
nand U9299 (N_9299,N_8874,N_8931);
nor U9300 (N_9300,N_8936,N_8793);
nor U9301 (N_9301,N_8746,N_8597);
and U9302 (N_9302,N_8849,N_8827);
or U9303 (N_9303,N_8535,N_8794);
or U9304 (N_9304,N_8581,N_8570);
nor U9305 (N_9305,N_8854,N_8693);
nand U9306 (N_9306,N_8918,N_8590);
or U9307 (N_9307,N_8754,N_8846);
nand U9308 (N_9308,N_8598,N_8513);
nand U9309 (N_9309,N_8609,N_8831);
nor U9310 (N_9310,N_8739,N_8877);
nor U9311 (N_9311,N_8896,N_8857);
nand U9312 (N_9312,N_8741,N_8959);
or U9313 (N_9313,N_8577,N_8983);
nor U9314 (N_9314,N_8534,N_8740);
and U9315 (N_9315,N_8631,N_8990);
or U9316 (N_9316,N_8898,N_8613);
and U9317 (N_9317,N_8746,N_8646);
nand U9318 (N_9318,N_8626,N_8572);
or U9319 (N_9319,N_8970,N_8690);
and U9320 (N_9320,N_8667,N_8825);
nand U9321 (N_9321,N_8512,N_8992);
nor U9322 (N_9322,N_8872,N_8992);
and U9323 (N_9323,N_8906,N_8802);
nand U9324 (N_9324,N_8831,N_8771);
and U9325 (N_9325,N_8756,N_8597);
nand U9326 (N_9326,N_8527,N_8635);
nand U9327 (N_9327,N_8553,N_8612);
and U9328 (N_9328,N_8885,N_8616);
xnor U9329 (N_9329,N_8503,N_8516);
and U9330 (N_9330,N_8977,N_8644);
nor U9331 (N_9331,N_8954,N_8794);
and U9332 (N_9332,N_8723,N_8661);
and U9333 (N_9333,N_8897,N_8744);
nand U9334 (N_9334,N_8893,N_8555);
nand U9335 (N_9335,N_8976,N_8983);
nor U9336 (N_9336,N_8599,N_8606);
xor U9337 (N_9337,N_8729,N_8868);
nor U9338 (N_9338,N_8639,N_8716);
nand U9339 (N_9339,N_8823,N_8558);
nor U9340 (N_9340,N_8909,N_8704);
and U9341 (N_9341,N_8971,N_8963);
nor U9342 (N_9342,N_8803,N_8743);
nor U9343 (N_9343,N_8838,N_8853);
or U9344 (N_9344,N_8575,N_8886);
and U9345 (N_9345,N_8558,N_8726);
xor U9346 (N_9346,N_8526,N_8789);
xnor U9347 (N_9347,N_8616,N_8900);
or U9348 (N_9348,N_8943,N_8611);
nand U9349 (N_9349,N_8761,N_8895);
and U9350 (N_9350,N_8915,N_8823);
and U9351 (N_9351,N_8619,N_8757);
or U9352 (N_9352,N_8794,N_8667);
nor U9353 (N_9353,N_8527,N_8951);
and U9354 (N_9354,N_8949,N_8511);
and U9355 (N_9355,N_8831,N_8527);
nor U9356 (N_9356,N_8717,N_8788);
xnor U9357 (N_9357,N_8546,N_8903);
nand U9358 (N_9358,N_8895,N_8674);
nor U9359 (N_9359,N_8794,N_8647);
and U9360 (N_9360,N_8844,N_8662);
or U9361 (N_9361,N_8561,N_8802);
and U9362 (N_9362,N_8861,N_8823);
and U9363 (N_9363,N_8989,N_8944);
or U9364 (N_9364,N_8555,N_8985);
or U9365 (N_9365,N_8956,N_8992);
nand U9366 (N_9366,N_8831,N_8759);
or U9367 (N_9367,N_8765,N_8969);
nor U9368 (N_9368,N_8910,N_8916);
nand U9369 (N_9369,N_8548,N_8922);
nor U9370 (N_9370,N_8607,N_8966);
nor U9371 (N_9371,N_8527,N_8573);
nand U9372 (N_9372,N_8507,N_8697);
or U9373 (N_9373,N_8828,N_8536);
nor U9374 (N_9374,N_8562,N_8632);
or U9375 (N_9375,N_8606,N_8652);
nand U9376 (N_9376,N_8911,N_8598);
nand U9377 (N_9377,N_8654,N_8717);
nor U9378 (N_9378,N_8650,N_8578);
nand U9379 (N_9379,N_8944,N_8671);
or U9380 (N_9380,N_8891,N_8755);
and U9381 (N_9381,N_8937,N_8787);
nand U9382 (N_9382,N_8560,N_8716);
nor U9383 (N_9383,N_8769,N_8631);
or U9384 (N_9384,N_8703,N_8641);
nand U9385 (N_9385,N_8639,N_8735);
nor U9386 (N_9386,N_8952,N_8809);
xnor U9387 (N_9387,N_8950,N_8581);
and U9388 (N_9388,N_8559,N_8902);
nand U9389 (N_9389,N_8675,N_8711);
or U9390 (N_9390,N_8578,N_8927);
nor U9391 (N_9391,N_8765,N_8642);
and U9392 (N_9392,N_8590,N_8815);
nor U9393 (N_9393,N_8666,N_8606);
nor U9394 (N_9394,N_8966,N_8878);
nor U9395 (N_9395,N_8693,N_8702);
xnor U9396 (N_9396,N_8515,N_8767);
or U9397 (N_9397,N_8608,N_8536);
or U9398 (N_9398,N_8730,N_8991);
nor U9399 (N_9399,N_8898,N_8591);
or U9400 (N_9400,N_8874,N_8889);
xnor U9401 (N_9401,N_8533,N_8990);
nor U9402 (N_9402,N_8546,N_8827);
nor U9403 (N_9403,N_8620,N_8619);
and U9404 (N_9404,N_8612,N_8756);
and U9405 (N_9405,N_8616,N_8618);
nor U9406 (N_9406,N_8588,N_8782);
xor U9407 (N_9407,N_8926,N_8615);
or U9408 (N_9408,N_8813,N_8823);
nand U9409 (N_9409,N_8615,N_8661);
nor U9410 (N_9410,N_8720,N_8935);
or U9411 (N_9411,N_8532,N_8967);
nor U9412 (N_9412,N_8629,N_8614);
and U9413 (N_9413,N_8661,N_8558);
or U9414 (N_9414,N_8526,N_8835);
nand U9415 (N_9415,N_8939,N_8807);
or U9416 (N_9416,N_8917,N_8740);
nor U9417 (N_9417,N_8773,N_8608);
nand U9418 (N_9418,N_8657,N_8688);
nand U9419 (N_9419,N_8801,N_8860);
nand U9420 (N_9420,N_8675,N_8881);
and U9421 (N_9421,N_8734,N_8964);
xor U9422 (N_9422,N_8979,N_8730);
or U9423 (N_9423,N_8544,N_8626);
or U9424 (N_9424,N_8956,N_8961);
nor U9425 (N_9425,N_8680,N_8970);
nor U9426 (N_9426,N_8556,N_8612);
and U9427 (N_9427,N_8563,N_8679);
xor U9428 (N_9428,N_8994,N_8679);
nor U9429 (N_9429,N_8951,N_8884);
or U9430 (N_9430,N_8761,N_8606);
or U9431 (N_9431,N_8592,N_8502);
and U9432 (N_9432,N_8811,N_8578);
xor U9433 (N_9433,N_8951,N_8795);
or U9434 (N_9434,N_8898,N_8619);
nor U9435 (N_9435,N_8899,N_8695);
nor U9436 (N_9436,N_8902,N_8792);
nand U9437 (N_9437,N_8918,N_8573);
and U9438 (N_9438,N_8657,N_8932);
and U9439 (N_9439,N_8888,N_8518);
or U9440 (N_9440,N_8867,N_8573);
or U9441 (N_9441,N_8770,N_8557);
or U9442 (N_9442,N_8827,N_8635);
or U9443 (N_9443,N_8703,N_8547);
nor U9444 (N_9444,N_8577,N_8666);
and U9445 (N_9445,N_8643,N_8626);
nor U9446 (N_9446,N_8655,N_8502);
or U9447 (N_9447,N_8851,N_8739);
nor U9448 (N_9448,N_8928,N_8795);
nor U9449 (N_9449,N_8783,N_8786);
nand U9450 (N_9450,N_8643,N_8714);
xnor U9451 (N_9451,N_8930,N_8931);
and U9452 (N_9452,N_8717,N_8625);
and U9453 (N_9453,N_8743,N_8824);
and U9454 (N_9454,N_8990,N_8889);
nor U9455 (N_9455,N_8639,N_8919);
and U9456 (N_9456,N_8637,N_8639);
and U9457 (N_9457,N_8591,N_8834);
xor U9458 (N_9458,N_8905,N_8735);
or U9459 (N_9459,N_8501,N_8905);
and U9460 (N_9460,N_8958,N_8835);
and U9461 (N_9461,N_8533,N_8911);
nand U9462 (N_9462,N_8913,N_8881);
or U9463 (N_9463,N_8686,N_8960);
nand U9464 (N_9464,N_8622,N_8585);
nand U9465 (N_9465,N_8867,N_8923);
nor U9466 (N_9466,N_8955,N_8589);
nand U9467 (N_9467,N_8689,N_8573);
or U9468 (N_9468,N_8545,N_8783);
xnor U9469 (N_9469,N_8816,N_8698);
xnor U9470 (N_9470,N_8987,N_8983);
and U9471 (N_9471,N_8593,N_8803);
nand U9472 (N_9472,N_8932,N_8858);
nand U9473 (N_9473,N_8534,N_8604);
or U9474 (N_9474,N_8739,N_8530);
nor U9475 (N_9475,N_8564,N_8646);
nand U9476 (N_9476,N_8714,N_8969);
and U9477 (N_9477,N_8608,N_8741);
and U9478 (N_9478,N_8662,N_8780);
nand U9479 (N_9479,N_8560,N_8703);
or U9480 (N_9480,N_8636,N_8778);
and U9481 (N_9481,N_8923,N_8784);
and U9482 (N_9482,N_8620,N_8863);
nand U9483 (N_9483,N_8909,N_8526);
or U9484 (N_9484,N_8828,N_8862);
xor U9485 (N_9485,N_8630,N_8553);
nor U9486 (N_9486,N_8661,N_8561);
or U9487 (N_9487,N_8985,N_8906);
nand U9488 (N_9488,N_8847,N_8817);
and U9489 (N_9489,N_8544,N_8956);
nor U9490 (N_9490,N_8759,N_8974);
or U9491 (N_9491,N_8950,N_8550);
nor U9492 (N_9492,N_8838,N_8728);
and U9493 (N_9493,N_8940,N_8706);
and U9494 (N_9494,N_8665,N_8790);
nand U9495 (N_9495,N_8849,N_8505);
or U9496 (N_9496,N_8518,N_8893);
xor U9497 (N_9497,N_8854,N_8978);
nand U9498 (N_9498,N_8644,N_8564);
and U9499 (N_9499,N_8985,N_8731);
nor U9500 (N_9500,N_9080,N_9034);
or U9501 (N_9501,N_9443,N_9315);
nand U9502 (N_9502,N_9298,N_9299);
and U9503 (N_9503,N_9096,N_9106);
and U9504 (N_9504,N_9002,N_9097);
and U9505 (N_9505,N_9394,N_9091);
and U9506 (N_9506,N_9350,N_9090);
nor U9507 (N_9507,N_9488,N_9159);
and U9508 (N_9508,N_9463,N_9458);
nor U9509 (N_9509,N_9012,N_9473);
or U9510 (N_9510,N_9406,N_9476);
nor U9511 (N_9511,N_9059,N_9128);
nor U9512 (N_9512,N_9093,N_9172);
nor U9513 (N_9513,N_9494,N_9150);
and U9514 (N_9514,N_9317,N_9414);
and U9515 (N_9515,N_9353,N_9453);
or U9516 (N_9516,N_9135,N_9274);
or U9517 (N_9517,N_9191,N_9114);
and U9518 (N_9518,N_9492,N_9244);
xnor U9519 (N_9519,N_9115,N_9016);
nor U9520 (N_9520,N_9209,N_9204);
nand U9521 (N_9521,N_9491,N_9156);
or U9522 (N_9522,N_9457,N_9258);
nand U9523 (N_9523,N_9283,N_9264);
nand U9524 (N_9524,N_9027,N_9141);
or U9525 (N_9525,N_9247,N_9326);
or U9526 (N_9526,N_9266,N_9316);
nand U9527 (N_9527,N_9222,N_9278);
and U9528 (N_9528,N_9478,N_9388);
nor U9529 (N_9529,N_9177,N_9045);
nand U9530 (N_9530,N_9486,N_9065);
nand U9531 (N_9531,N_9270,N_9184);
nand U9532 (N_9532,N_9276,N_9286);
or U9533 (N_9533,N_9289,N_9238);
nand U9534 (N_9534,N_9195,N_9387);
nand U9535 (N_9535,N_9176,N_9143);
or U9536 (N_9536,N_9032,N_9261);
nor U9537 (N_9537,N_9461,N_9225);
and U9538 (N_9538,N_9066,N_9239);
and U9539 (N_9539,N_9446,N_9226);
or U9540 (N_9540,N_9487,N_9235);
or U9541 (N_9541,N_9181,N_9426);
nand U9542 (N_9542,N_9341,N_9448);
and U9543 (N_9543,N_9372,N_9237);
and U9544 (N_9544,N_9419,N_9173);
nand U9545 (N_9545,N_9241,N_9163);
nor U9546 (N_9546,N_9210,N_9355);
or U9547 (N_9547,N_9349,N_9004);
nand U9548 (N_9548,N_9440,N_9095);
nand U9549 (N_9549,N_9193,N_9409);
or U9550 (N_9550,N_9099,N_9134);
xnor U9551 (N_9551,N_9285,N_9309);
nand U9552 (N_9552,N_9380,N_9468);
nand U9553 (N_9553,N_9149,N_9370);
xor U9554 (N_9554,N_9190,N_9365);
xor U9555 (N_9555,N_9393,N_9399);
and U9556 (N_9556,N_9233,N_9232);
and U9557 (N_9557,N_9178,N_9101);
and U9558 (N_9558,N_9332,N_9021);
or U9559 (N_9559,N_9438,N_9146);
or U9560 (N_9560,N_9214,N_9078);
or U9561 (N_9561,N_9411,N_9329);
nand U9562 (N_9562,N_9382,N_9123);
and U9563 (N_9563,N_9073,N_9452);
nand U9564 (N_9564,N_9109,N_9416);
and U9565 (N_9565,N_9445,N_9312);
xor U9566 (N_9566,N_9250,N_9075);
nor U9567 (N_9567,N_9379,N_9265);
or U9568 (N_9568,N_9168,N_9052);
or U9569 (N_9569,N_9061,N_9144);
nor U9570 (N_9570,N_9484,N_9105);
nor U9571 (N_9571,N_9194,N_9389);
nand U9572 (N_9572,N_9104,N_9408);
nor U9573 (N_9573,N_9249,N_9088);
xor U9574 (N_9574,N_9174,N_9005);
or U9575 (N_9575,N_9364,N_9010);
or U9576 (N_9576,N_9152,N_9248);
and U9577 (N_9577,N_9122,N_9171);
nand U9578 (N_9578,N_9479,N_9040);
and U9579 (N_9579,N_9183,N_9424);
nand U9580 (N_9580,N_9398,N_9175);
nand U9581 (N_9581,N_9340,N_9337);
and U9582 (N_9582,N_9131,N_9142);
and U9583 (N_9583,N_9098,N_9369);
and U9584 (N_9584,N_9459,N_9023);
xnor U9585 (N_9585,N_9236,N_9068);
or U9586 (N_9586,N_9386,N_9475);
nand U9587 (N_9587,N_9102,N_9197);
or U9588 (N_9588,N_9138,N_9058);
and U9589 (N_9589,N_9344,N_9026);
and U9590 (N_9590,N_9334,N_9203);
nor U9591 (N_9591,N_9331,N_9162);
nor U9592 (N_9592,N_9219,N_9383);
or U9593 (N_9593,N_9018,N_9308);
or U9594 (N_9594,N_9303,N_9410);
or U9595 (N_9595,N_9067,N_9255);
and U9596 (N_9596,N_9240,N_9124);
nand U9597 (N_9597,N_9015,N_9116);
xor U9598 (N_9598,N_9467,N_9200);
and U9599 (N_9599,N_9215,N_9140);
or U9600 (N_9600,N_9043,N_9154);
or U9601 (N_9601,N_9199,N_9082);
and U9602 (N_9602,N_9218,N_9384);
or U9603 (N_9603,N_9480,N_9335);
nor U9604 (N_9604,N_9430,N_9437);
nand U9605 (N_9605,N_9413,N_9062);
and U9606 (N_9606,N_9420,N_9280);
xor U9607 (N_9607,N_9489,N_9187);
and U9608 (N_9608,N_9363,N_9381);
and U9609 (N_9609,N_9423,N_9305);
and U9610 (N_9610,N_9451,N_9050);
nor U9611 (N_9611,N_9338,N_9465);
nor U9612 (N_9612,N_9185,N_9092);
and U9613 (N_9613,N_9060,N_9361);
nand U9614 (N_9614,N_9390,N_9313);
and U9615 (N_9615,N_9330,N_9132);
nor U9616 (N_9616,N_9297,N_9160);
or U9617 (N_9617,N_9469,N_9396);
nand U9618 (N_9618,N_9000,N_9017);
xnor U9619 (N_9619,N_9495,N_9269);
nand U9620 (N_9620,N_9161,N_9454);
nand U9621 (N_9621,N_9311,N_9327);
and U9622 (N_9622,N_9301,N_9351);
nor U9623 (N_9623,N_9352,N_9014);
nand U9624 (N_9624,N_9107,N_9153);
nand U9625 (N_9625,N_9300,N_9339);
and U9626 (N_9626,N_9074,N_9253);
nand U9627 (N_9627,N_9063,N_9234);
nand U9628 (N_9628,N_9112,N_9378);
xnor U9629 (N_9629,N_9434,N_9356);
nand U9630 (N_9630,N_9007,N_9306);
nor U9631 (N_9631,N_9277,N_9125);
and U9632 (N_9632,N_9211,N_9366);
nor U9633 (N_9633,N_9466,N_9348);
nand U9634 (N_9634,N_9483,N_9165);
or U9635 (N_9635,N_9231,N_9385);
xor U9636 (N_9636,N_9296,N_9263);
and U9637 (N_9637,N_9456,N_9071);
xnor U9638 (N_9638,N_9011,N_9275);
or U9639 (N_9639,N_9288,N_9037);
or U9640 (N_9640,N_9496,N_9282);
or U9641 (N_9641,N_9243,N_9357);
or U9642 (N_9642,N_9431,N_9281);
and U9643 (N_9643,N_9039,N_9499);
nor U9644 (N_9644,N_9170,N_9217);
or U9645 (N_9645,N_9081,N_9262);
or U9646 (N_9646,N_9333,N_9103);
and U9647 (N_9647,N_9418,N_9498);
or U9648 (N_9648,N_9360,N_9442);
nor U9649 (N_9649,N_9208,N_9205);
or U9650 (N_9650,N_9460,N_9256);
or U9651 (N_9651,N_9164,N_9359);
nand U9652 (N_9652,N_9314,N_9148);
nand U9653 (N_9653,N_9345,N_9433);
nor U9654 (N_9654,N_9464,N_9375);
or U9655 (N_9655,N_9192,N_9323);
and U9656 (N_9656,N_9001,N_9425);
or U9657 (N_9657,N_9127,N_9358);
nor U9658 (N_9658,N_9048,N_9472);
and U9659 (N_9659,N_9242,N_9436);
nor U9660 (N_9660,N_9292,N_9428);
and U9661 (N_9661,N_9450,N_9415);
nand U9662 (N_9662,N_9343,N_9304);
or U9663 (N_9663,N_9158,N_9367);
nand U9664 (N_9664,N_9019,N_9259);
nand U9665 (N_9665,N_9049,N_9047);
or U9666 (N_9666,N_9167,N_9354);
nand U9667 (N_9667,N_9395,N_9076);
nor U9668 (N_9668,N_9252,N_9251);
or U9669 (N_9669,N_9377,N_9470);
or U9670 (N_9670,N_9402,N_9405);
and U9671 (N_9671,N_9121,N_9421);
nor U9672 (N_9672,N_9056,N_9441);
nand U9673 (N_9673,N_9042,N_9295);
nand U9674 (N_9674,N_9179,N_9051);
and U9675 (N_9675,N_9328,N_9145);
and U9676 (N_9676,N_9272,N_9287);
or U9677 (N_9677,N_9435,N_9432);
and U9678 (N_9678,N_9151,N_9257);
nor U9679 (N_9679,N_9346,N_9245);
or U9680 (N_9680,N_9033,N_9025);
nor U9681 (N_9681,N_9227,N_9212);
or U9682 (N_9682,N_9273,N_9485);
nor U9683 (N_9683,N_9284,N_9182);
nand U9684 (N_9684,N_9449,N_9024);
nand U9685 (N_9685,N_9188,N_9279);
xnor U9686 (N_9686,N_9412,N_9336);
nor U9687 (N_9687,N_9008,N_9035);
nand U9688 (N_9688,N_9302,N_9223);
and U9689 (N_9689,N_9447,N_9422);
nor U9690 (N_9690,N_9129,N_9044);
or U9691 (N_9691,N_9401,N_9130);
or U9692 (N_9692,N_9046,N_9079);
nand U9693 (N_9693,N_9224,N_9006);
nor U9694 (N_9694,N_9268,N_9342);
nand U9695 (N_9695,N_9147,N_9157);
nand U9696 (N_9696,N_9166,N_9371);
and U9697 (N_9697,N_9117,N_9089);
xor U9698 (N_9698,N_9009,N_9290);
or U9699 (N_9699,N_9403,N_9028);
xor U9700 (N_9700,N_9321,N_9490);
nand U9701 (N_9701,N_9029,N_9254);
nand U9702 (N_9702,N_9022,N_9201);
and U9703 (N_9703,N_9271,N_9221);
nor U9704 (N_9704,N_9110,N_9325);
nand U9705 (N_9705,N_9041,N_9155);
nor U9706 (N_9706,N_9213,N_9216);
nor U9707 (N_9707,N_9083,N_9020);
or U9708 (N_9708,N_9031,N_9444);
nor U9709 (N_9709,N_9230,N_9202);
and U9710 (N_9710,N_9113,N_9198);
or U9711 (N_9711,N_9220,N_9455);
nand U9712 (N_9712,N_9189,N_9482);
and U9713 (N_9713,N_9180,N_9206);
nor U9714 (N_9714,N_9094,N_9477);
nand U9715 (N_9715,N_9374,N_9310);
nand U9716 (N_9716,N_9347,N_9417);
nand U9717 (N_9717,N_9086,N_9186);
nor U9718 (N_9718,N_9319,N_9307);
xnor U9719 (N_9719,N_9376,N_9126);
nand U9720 (N_9720,N_9036,N_9397);
or U9721 (N_9721,N_9087,N_9139);
and U9722 (N_9722,N_9246,N_9493);
nand U9723 (N_9723,N_9072,N_9462);
or U9724 (N_9724,N_9324,N_9400);
or U9725 (N_9725,N_9038,N_9003);
nor U9726 (N_9726,N_9118,N_9057);
xnor U9727 (N_9727,N_9229,N_9069);
or U9728 (N_9728,N_9108,N_9260);
or U9729 (N_9729,N_9404,N_9196);
nor U9730 (N_9730,N_9119,N_9294);
nand U9731 (N_9731,N_9322,N_9362);
or U9732 (N_9732,N_9497,N_9320);
xor U9733 (N_9733,N_9427,N_9373);
nor U9734 (N_9734,N_9439,N_9391);
nand U9735 (N_9735,N_9407,N_9077);
or U9736 (N_9736,N_9137,N_9291);
nor U9737 (N_9737,N_9054,N_9120);
or U9738 (N_9738,N_9064,N_9053);
or U9739 (N_9739,N_9481,N_9429);
xor U9740 (N_9740,N_9169,N_9293);
and U9741 (N_9741,N_9013,N_9207);
nor U9742 (N_9742,N_9136,N_9070);
xor U9743 (N_9743,N_9133,N_9474);
and U9744 (N_9744,N_9392,N_9111);
and U9745 (N_9745,N_9318,N_9055);
nor U9746 (N_9746,N_9368,N_9100);
and U9747 (N_9747,N_9228,N_9085);
nor U9748 (N_9748,N_9471,N_9030);
and U9749 (N_9749,N_9084,N_9267);
nor U9750 (N_9750,N_9457,N_9084);
and U9751 (N_9751,N_9398,N_9079);
nand U9752 (N_9752,N_9197,N_9300);
nand U9753 (N_9753,N_9345,N_9091);
or U9754 (N_9754,N_9079,N_9380);
or U9755 (N_9755,N_9069,N_9467);
or U9756 (N_9756,N_9343,N_9066);
xor U9757 (N_9757,N_9072,N_9355);
nor U9758 (N_9758,N_9193,N_9157);
nand U9759 (N_9759,N_9457,N_9014);
or U9760 (N_9760,N_9197,N_9008);
nor U9761 (N_9761,N_9345,N_9148);
nand U9762 (N_9762,N_9026,N_9177);
or U9763 (N_9763,N_9387,N_9447);
and U9764 (N_9764,N_9460,N_9214);
and U9765 (N_9765,N_9382,N_9410);
nor U9766 (N_9766,N_9000,N_9087);
nor U9767 (N_9767,N_9123,N_9232);
nor U9768 (N_9768,N_9323,N_9325);
or U9769 (N_9769,N_9247,N_9105);
nand U9770 (N_9770,N_9052,N_9019);
or U9771 (N_9771,N_9278,N_9459);
nand U9772 (N_9772,N_9044,N_9452);
nand U9773 (N_9773,N_9024,N_9073);
nand U9774 (N_9774,N_9128,N_9184);
nand U9775 (N_9775,N_9081,N_9217);
nand U9776 (N_9776,N_9147,N_9181);
and U9777 (N_9777,N_9187,N_9362);
or U9778 (N_9778,N_9230,N_9098);
nand U9779 (N_9779,N_9047,N_9400);
nand U9780 (N_9780,N_9113,N_9451);
and U9781 (N_9781,N_9317,N_9270);
nand U9782 (N_9782,N_9370,N_9046);
nand U9783 (N_9783,N_9162,N_9493);
nand U9784 (N_9784,N_9278,N_9213);
and U9785 (N_9785,N_9074,N_9376);
nand U9786 (N_9786,N_9043,N_9267);
or U9787 (N_9787,N_9029,N_9117);
and U9788 (N_9788,N_9324,N_9362);
and U9789 (N_9789,N_9388,N_9375);
or U9790 (N_9790,N_9348,N_9305);
and U9791 (N_9791,N_9426,N_9063);
nor U9792 (N_9792,N_9446,N_9192);
nor U9793 (N_9793,N_9085,N_9324);
nand U9794 (N_9794,N_9291,N_9120);
or U9795 (N_9795,N_9182,N_9030);
or U9796 (N_9796,N_9214,N_9130);
xnor U9797 (N_9797,N_9158,N_9465);
nand U9798 (N_9798,N_9398,N_9168);
or U9799 (N_9799,N_9230,N_9350);
or U9800 (N_9800,N_9157,N_9284);
xnor U9801 (N_9801,N_9378,N_9380);
and U9802 (N_9802,N_9408,N_9420);
nor U9803 (N_9803,N_9063,N_9398);
or U9804 (N_9804,N_9040,N_9214);
and U9805 (N_9805,N_9496,N_9132);
nor U9806 (N_9806,N_9461,N_9189);
xnor U9807 (N_9807,N_9232,N_9412);
xor U9808 (N_9808,N_9226,N_9387);
nor U9809 (N_9809,N_9350,N_9015);
xnor U9810 (N_9810,N_9070,N_9155);
or U9811 (N_9811,N_9474,N_9174);
or U9812 (N_9812,N_9004,N_9443);
and U9813 (N_9813,N_9094,N_9435);
nor U9814 (N_9814,N_9132,N_9348);
or U9815 (N_9815,N_9144,N_9097);
nor U9816 (N_9816,N_9029,N_9132);
or U9817 (N_9817,N_9426,N_9403);
and U9818 (N_9818,N_9219,N_9334);
and U9819 (N_9819,N_9423,N_9394);
xnor U9820 (N_9820,N_9339,N_9399);
or U9821 (N_9821,N_9301,N_9417);
nand U9822 (N_9822,N_9231,N_9452);
or U9823 (N_9823,N_9057,N_9073);
and U9824 (N_9824,N_9132,N_9227);
or U9825 (N_9825,N_9081,N_9400);
or U9826 (N_9826,N_9037,N_9347);
xor U9827 (N_9827,N_9238,N_9096);
or U9828 (N_9828,N_9026,N_9044);
xor U9829 (N_9829,N_9020,N_9479);
nor U9830 (N_9830,N_9196,N_9472);
nor U9831 (N_9831,N_9453,N_9470);
nor U9832 (N_9832,N_9184,N_9214);
xnor U9833 (N_9833,N_9328,N_9114);
xor U9834 (N_9834,N_9260,N_9402);
and U9835 (N_9835,N_9359,N_9403);
or U9836 (N_9836,N_9200,N_9485);
xnor U9837 (N_9837,N_9474,N_9270);
nand U9838 (N_9838,N_9015,N_9025);
xor U9839 (N_9839,N_9420,N_9444);
nor U9840 (N_9840,N_9242,N_9284);
and U9841 (N_9841,N_9145,N_9394);
nand U9842 (N_9842,N_9361,N_9342);
nand U9843 (N_9843,N_9071,N_9337);
nand U9844 (N_9844,N_9065,N_9004);
or U9845 (N_9845,N_9455,N_9186);
xnor U9846 (N_9846,N_9133,N_9283);
nor U9847 (N_9847,N_9070,N_9260);
nor U9848 (N_9848,N_9155,N_9454);
nor U9849 (N_9849,N_9202,N_9357);
and U9850 (N_9850,N_9131,N_9323);
and U9851 (N_9851,N_9463,N_9384);
nor U9852 (N_9852,N_9075,N_9415);
nand U9853 (N_9853,N_9337,N_9195);
and U9854 (N_9854,N_9344,N_9179);
nand U9855 (N_9855,N_9263,N_9411);
or U9856 (N_9856,N_9261,N_9026);
nand U9857 (N_9857,N_9081,N_9351);
nor U9858 (N_9858,N_9027,N_9090);
or U9859 (N_9859,N_9162,N_9387);
or U9860 (N_9860,N_9214,N_9165);
nor U9861 (N_9861,N_9134,N_9121);
nor U9862 (N_9862,N_9146,N_9182);
or U9863 (N_9863,N_9450,N_9414);
and U9864 (N_9864,N_9142,N_9014);
xnor U9865 (N_9865,N_9366,N_9227);
and U9866 (N_9866,N_9238,N_9001);
nor U9867 (N_9867,N_9079,N_9059);
nand U9868 (N_9868,N_9331,N_9065);
nor U9869 (N_9869,N_9209,N_9075);
xnor U9870 (N_9870,N_9012,N_9059);
nand U9871 (N_9871,N_9317,N_9166);
nand U9872 (N_9872,N_9192,N_9251);
or U9873 (N_9873,N_9337,N_9051);
or U9874 (N_9874,N_9081,N_9301);
nand U9875 (N_9875,N_9496,N_9455);
and U9876 (N_9876,N_9374,N_9358);
nor U9877 (N_9877,N_9028,N_9120);
or U9878 (N_9878,N_9065,N_9097);
or U9879 (N_9879,N_9370,N_9029);
xor U9880 (N_9880,N_9442,N_9382);
xor U9881 (N_9881,N_9210,N_9181);
or U9882 (N_9882,N_9376,N_9402);
nor U9883 (N_9883,N_9040,N_9465);
nor U9884 (N_9884,N_9011,N_9151);
or U9885 (N_9885,N_9002,N_9272);
or U9886 (N_9886,N_9120,N_9448);
and U9887 (N_9887,N_9465,N_9028);
nand U9888 (N_9888,N_9020,N_9300);
nand U9889 (N_9889,N_9408,N_9404);
nand U9890 (N_9890,N_9406,N_9065);
or U9891 (N_9891,N_9279,N_9475);
or U9892 (N_9892,N_9309,N_9115);
nor U9893 (N_9893,N_9463,N_9074);
and U9894 (N_9894,N_9281,N_9499);
nand U9895 (N_9895,N_9009,N_9339);
nor U9896 (N_9896,N_9264,N_9066);
and U9897 (N_9897,N_9221,N_9396);
and U9898 (N_9898,N_9146,N_9030);
and U9899 (N_9899,N_9365,N_9200);
xor U9900 (N_9900,N_9289,N_9286);
or U9901 (N_9901,N_9070,N_9046);
and U9902 (N_9902,N_9175,N_9325);
or U9903 (N_9903,N_9390,N_9276);
and U9904 (N_9904,N_9366,N_9411);
and U9905 (N_9905,N_9103,N_9036);
or U9906 (N_9906,N_9447,N_9214);
nand U9907 (N_9907,N_9478,N_9355);
or U9908 (N_9908,N_9166,N_9411);
nand U9909 (N_9909,N_9165,N_9486);
xor U9910 (N_9910,N_9384,N_9246);
and U9911 (N_9911,N_9435,N_9074);
xor U9912 (N_9912,N_9191,N_9021);
nor U9913 (N_9913,N_9326,N_9419);
or U9914 (N_9914,N_9243,N_9419);
and U9915 (N_9915,N_9076,N_9048);
nand U9916 (N_9916,N_9334,N_9032);
and U9917 (N_9917,N_9147,N_9288);
or U9918 (N_9918,N_9336,N_9158);
nor U9919 (N_9919,N_9286,N_9166);
or U9920 (N_9920,N_9329,N_9284);
nand U9921 (N_9921,N_9251,N_9242);
xor U9922 (N_9922,N_9058,N_9325);
nand U9923 (N_9923,N_9119,N_9441);
nand U9924 (N_9924,N_9031,N_9317);
xor U9925 (N_9925,N_9056,N_9029);
nor U9926 (N_9926,N_9062,N_9423);
nor U9927 (N_9927,N_9378,N_9269);
nor U9928 (N_9928,N_9037,N_9085);
xnor U9929 (N_9929,N_9183,N_9244);
and U9930 (N_9930,N_9296,N_9185);
xnor U9931 (N_9931,N_9135,N_9319);
and U9932 (N_9932,N_9282,N_9263);
nand U9933 (N_9933,N_9071,N_9444);
and U9934 (N_9934,N_9354,N_9144);
and U9935 (N_9935,N_9067,N_9119);
nor U9936 (N_9936,N_9046,N_9450);
nand U9937 (N_9937,N_9477,N_9124);
nor U9938 (N_9938,N_9035,N_9235);
and U9939 (N_9939,N_9417,N_9010);
or U9940 (N_9940,N_9028,N_9100);
nor U9941 (N_9941,N_9017,N_9041);
nor U9942 (N_9942,N_9404,N_9183);
nand U9943 (N_9943,N_9303,N_9320);
nand U9944 (N_9944,N_9080,N_9173);
nor U9945 (N_9945,N_9088,N_9256);
and U9946 (N_9946,N_9064,N_9167);
nand U9947 (N_9947,N_9381,N_9479);
and U9948 (N_9948,N_9281,N_9326);
nor U9949 (N_9949,N_9082,N_9084);
nand U9950 (N_9950,N_9063,N_9307);
nor U9951 (N_9951,N_9091,N_9329);
or U9952 (N_9952,N_9381,N_9086);
or U9953 (N_9953,N_9443,N_9312);
or U9954 (N_9954,N_9450,N_9157);
xnor U9955 (N_9955,N_9205,N_9364);
and U9956 (N_9956,N_9258,N_9102);
nor U9957 (N_9957,N_9494,N_9154);
and U9958 (N_9958,N_9359,N_9236);
nand U9959 (N_9959,N_9392,N_9215);
nor U9960 (N_9960,N_9088,N_9494);
or U9961 (N_9961,N_9062,N_9163);
nand U9962 (N_9962,N_9203,N_9275);
nand U9963 (N_9963,N_9441,N_9448);
nand U9964 (N_9964,N_9350,N_9477);
and U9965 (N_9965,N_9278,N_9220);
and U9966 (N_9966,N_9369,N_9280);
or U9967 (N_9967,N_9274,N_9270);
xnor U9968 (N_9968,N_9263,N_9142);
nand U9969 (N_9969,N_9125,N_9416);
and U9970 (N_9970,N_9089,N_9379);
nand U9971 (N_9971,N_9052,N_9319);
nand U9972 (N_9972,N_9138,N_9048);
and U9973 (N_9973,N_9210,N_9241);
and U9974 (N_9974,N_9216,N_9415);
xor U9975 (N_9975,N_9054,N_9403);
or U9976 (N_9976,N_9253,N_9012);
nor U9977 (N_9977,N_9025,N_9303);
nand U9978 (N_9978,N_9024,N_9379);
nand U9979 (N_9979,N_9118,N_9360);
nor U9980 (N_9980,N_9013,N_9404);
or U9981 (N_9981,N_9285,N_9163);
and U9982 (N_9982,N_9323,N_9343);
or U9983 (N_9983,N_9002,N_9495);
nor U9984 (N_9984,N_9386,N_9389);
nor U9985 (N_9985,N_9014,N_9400);
or U9986 (N_9986,N_9354,N_9084);
and U9987 (N_9987,N_9390,N_9335);
or U9988 (N_9988,N_9383,N_9376);
nand U9989 (N_9989,N_9423,N_9437);
or U9990 (N_9990,N_9417,N_9261);
or U9991 (N_9991,N_9466,N_9270);
and U9992 (N_9992,N_9183,N_9285);
nor U9993 (N_9993,N_9109,N_9479);
nand U9994 (N_9994,N_9189,N_9260);
nor U9995 (N_9995,N_9290,N_9061);
or U9996 (N_9996,N_9045,N_9249);
nand U9997 (N_9997,N_9286,N_9059);
nand U9998 (N_9998,N_9300,N_9317);
nand U9999 (N_9999,N_9275,N_9290);
and U10000 (N_10000,N_9918,N_9945);
and U10001 (N_10001,N_9657,N_9916);
xor U10002 (N_10002,N_9723,N_9740);
and U10003 (N_10003,N_9807,N_9690);
and U10004 (N_10004,N_9583,N_9558);
or U10005 (N_10005,N_9813,N_9984);
nor U10006 (N_10006,N_9935,N_9570);
or U10007 (N_10007,N_9903,N_9981);
nand U10008 (N_10008,N_9697,N_9555);
and U10009 (N_10009,N_9760,N_9966);
xor U10010 (N_10010,N_9993,N_9861);
nand U10011 (N_10011,N_9609,N_9963);
and U10012 (N_10012,N_9602,N_9702);
or U10013 (N_10013,N_9736,N_9923);
and U10014 (N_10014,N_9961,N_9587);
or U10015 (N_10015,N_9634,N_9739);
nor U10016 (N_10016,N_9910,N_9548);
nor U10017 (N_10017,N_9643,N_9844);
and U10018 (N_10018,N_9667,N_9990);
xor U10019 (N_10019,N_9779,N_9573);
or U10020 (N_10020,N_9670,N_9591);
xor U10021 (N_10021,N_9825,N_9906);
nor U10022 (N_10022,N_9939,N_9654);
or U10023 (N_10023,N_9693,N_9630);
or U10024 (N_10024,N_9501,N_9970);
nand U10025 (N_10025,N_9783,N_9733);
nand U10026 (N_10026,N_9518,N_9873);
nand U10027 (N_10027,N_9732,N_9680);
and U10028 (N_10028,N_9784,N_9800);
and U10029 (N_10029,N_9526,N_9631);
or U10030 (N_10030,N_9824,N_9827);
and U10031 (N_10031,N_9930,N_9892);
nand U10032 (N_10032,N_9547,N_9545);
nand U10033 (N_10033,N_9994,N_9794);
nand U10034 (N_10034,N_9777,N_9705);
nand U10035 (N_10035,N_9729,N_9668);
and U10036 (N_10036,N_9589,N_9608);
and U10037 (N_10037,N_9864,N_9767);
nand U10038 (N_10038,N_9899,N_9720);
or U10039 (N_10039,N_9544,N_9940);
nand U10040 (N_10040,N_9571,N_9665);
and U10041 (N_10041,N_9623,N_9575);
nor U10042 (N_10042,N_9566,N_9572);
or U10043 (N_10043,N_9674,N_9941);
or U10044 (N_10044,N_9854,N_9673);
or U10045 (N_10045,N_9780,N_9655);
nand U10046 (N_10046,N_9817,N_9766);
nor U10047 (N_10047,N_9769,N_9770);
or U10048 (N_10048,N_9641,N_9848);
nand U10049 (N_10049,N_9815,N_9669);
nand U10050 (N_10050,N_9796,N_9836);
nor U10051 (N_10051,N_9682,N_9546);
nor U10052 (N_10052,N_9527,N_9746);
or U10053 (N_10053,N_9512,N_9859);
nor U10054 (N_10054,N_9958,N_9650);
or U10055 (N_10055,N_9709,N_9542);
or U10056 (N_10056,N_9600,N_9636);
or U10057 (N_10057,N_9831,N_9855);
and U10058 (N_10058,N_9754,N_9816);
nand U10059 (N_10059,N_9706,N_9964);
xnor U10060 (N_10060,N_9535,N_9627);
and U10061 (N_10061,N_9711,N_9744);
nor U10062 (N_10062,N_9637,N_9839);
nor U10063 (N_10063,N_9505,N_9778);
nand U10064 (N_10064,N_9771,N_9691);
xor U10065 (N_10065,N_9832,N_9624);
nand U10066 (N_10066,N_9629,N_9757);
or U10067 (N_10067,N_9722,N_9788);
nor U10068 (N_10068,N_9887,N_9793);
nand U10069 (N_10069,N_9974,N_9877);
xor U10070 (N_10070,N_9672,N_9536);
xor U10071 (N_10071,N_9897,N_9530);
nor U10072 (N_10072,N_9821,N_9504);
nand U10073 (N_10073,N_9797,N_9508);
and U10074 (N_10074,N_9590,N_9731);
and U10075 (N_10075,N_9931,N_9799);
or U10076 (N_10076,N_9612,N_9618);
nor U10077 (N_10077,N_9952,N_9648);
or U10078 (N_10078,N_9921,N_9912);
nor U10079 (N_10079,N_9528,N_9789);
or U10080 (N_10080,N_9932,N_9866);
nand U10081 (N_10081,N_9946,N_9606);
or U10082 (N_10082,N_9675,N_9726);
nand U10083 (N_10083,N_9653,N_9588);
nor U10084 (N_10084,N_9577,N_9886);
nand U10085 (N_10085,N_9878,N_9898);
and U10086 (N_10086,N_9805,N_9829);
and U10087 (N_10087,N_9947,N_9677);
or U10088 (N_10088,N_9696,N_9996);
nand U10089 (N_10089,N_9837,N_9911);
and U10090 (N_10090,N_9716,N_9664);
and U10091 (N_10091,N_9852,N_9721);
nor U10092 (N_10092,N_9534,N_9671);
or U10093 (N_10093,N_9632,N_9586);
nand U10094 (N_10094,N_9554,N_9728);
nor U10095 (N_10095,N_9895,N_9516);
or U10096 (N_10096,N_9986,N_9830);
nand U10097 (N_10097,N_9896,N_9810);
xnor U10098 (N_10098,N_9500,N_9870);
nor U10099 (N_10099,N_9568,N_9652);
nor U10100 (N_10100,N_9814,N_9510);
or U10101 (N_10101,N_9751,N_9642);
and U10102 (N_10102,N_9874,N_9734);
and U10103 (N_10103,N_9942,N_9742);
xor U10104 (N_10104,N_9978,N_9661);
xor U10105 (N_10105,N_9719,N_9663);
nand U10106 (N_10106,N_9714,N_9808);
nor U10107 (N_10107,N_9853,N_9578);
nor U10108 (N_10108,N_9552,N_9967);
or U10109 (N_10109,N_9871,N_9868);
xnor U10110 (N_10110,N_9698,N_9593);
nor U10111 (N_10111,N_9755,N_9803);
or U10112 (N_10112,N_9835,N_9781);
or U10113 (N_10113,N_9506,N_9743);
and U10114 (N_10114,N_9635,N_9948);
nand U10115 (N_10115,N_9867,N_9957);
xnor U10116 (N_10116,N_9764,N_9694);
nor U10117 (N_10117,N_9581,N_9953);
nand U10118 (N_10118,N_9900,N_9562);
nand U10119 (N_10119,N_9700,N_9532);
and U10120 (N_10120,N_9699,N_9934);
or U10121 (N_10121,N_9502,N_9750);
nor U10122 (N_10122,N_9782,N_9919);
and U10123 (N_10123,N_9620,N_9592);
nor U10124 (N_10124,N_9708,N_9598);
xor U10125 (N_10125,N_9791,N_9965);
nand U10126 (N_10126,N_9787,N_9882);
and U10127 (N_10127,N_9960,N_9718);
nand U10128 (N_10128,N_9869,N_9857);
nor U10129 (N_10129,N_9988,N_9768);
and U10130 (N_10130,N_9745,N_9975);
xor U10131 (N_10131,N_9991,N_9610);
nor U10132 (N_10132,N_9876,N_9804);
nand U10133 (N_10133,N_9891,N_9507);
nor U10134 (N_10134,N_9790,N_9724);
and U10135 (N_10135,N_9834,N_9759);
and U10136 (N_10136,N_9929,N_9601);
nand U10137 (N_10137,N_9617,N_9604);
nand U10138 (N_10138,N_9851,N_9905);
xor U10139 (N_10139,N_9968,N_9563);
and U10140 (N_10140,N_9543,N_9678);
nand U10141 (N_10141,N_9704,N_9713);
nor U10142 (N_10142,N_9893,N_9977);
or U10143 (N_10143,N_9614,N_9943);
nand U10144 (N_10144,N_9758,N_9594);
and U10145 (N_10145,N_9537,N_9540);
nand U10146 (N_10146,N_9687,N_9541);
nand U10147 (N_10147,N_9955,N_9599);
nor U10148 (N_10148,N_9828,N_9551);
or U10149 (N_10149,N_9569,N_9639);
nand U10150 (N_10150,N_9987,N_9515);
nand U10151 (N_10151,N_9725,N_9651);
and U10152 (N_10152,N_9607,N_9858);
xnor U10153 (N_10153,N_9884,N_9811);
or U10154 (N_10154,N_9904,N_9838);
and U10155 (N_10155,N_9511,N_9662);
or U10156 (N_10156,N_9514,N_9820);
or U10157 (N_10157,N_9951,N_9872);
nand U10158 (N_10158,N_9622,N_9956);
nand U10159 (N_10159,N_9765,N_9785);
or U10160 (N_10160,N_9559,N_9775);
xor U10161 (N_10161,N_9880,N_9936);
nor U10162 (N_10162,N_9525,N_9695);
nor U10163 (N_10163,N_9681,N_9860);
nand U10164 (N_10164,N_9626,N_9875);
nor U10165 (N_10165,N_9647,N_9688);
xor U10166 (N_10166,N_9567,N_9638);
nand U10167 (N_10167,N_9849,N_9944);
nand U10168 (N_10168,N_9727,N_9856);
and U10169 (N_10169,N_9850,N_9908);
nor U10170 (N_10170,N_9792,N_9761);
and U10171 (N_10171,N_9812,N_9596);
or U10172 (N_10172,N_9676,N_9863);
xor U10173 (N_10173,N_9881,N_9560);
nand U10174 (N_10174,N_9924,N_9841);
nor U10175 (N_10175,N_9922,N_9585);
nand U10176 (N_10176,N_9846,N_9616);
nand U10177 (N_10177,N_9801,N_9879);
nor U10178 (N_10178,N_9976,N_9749);
and U10179 (N_10179,N_9619,N_9818);
and U10180 (N_10180,N_9989,N_9628);
nor U10181 (N_10181,N_9692,N_9809);
nor U10182 (N_10182,N_9633,N_9640);
nand U10183 (N_10183,N_9972,N_9645);
or U10184 (N_10184,N_9579,N_9753);
or U10185 (N_10185,N_9533,N_9985);
nand U10186 (N_10186,N_9776,N_9995);
or U10187 (N_10187,N_9795,N_9524);
or U10188 (N_10188,N_9660,N_9938);
nor U10189 (N_10189,N_9703,N_9983);
and U10190 (N_10190,N_9920,N_9774);
and U10191 (N_10191,N_9520,N_9517);
xor U10192 (N_10192,N_9549,N_9747);
nor U10193 (N_10193,N_9576,N_9845);
nor U10194 (N_10194,N_9847,N_9580);
nor U10195 (N_10195,N_9683,N_9959);
or U10196 (N_10196,N_9752,N_9786);
and U10197 (N_10197,N_9584,N_9862);
or U10198 (N_10198,N_9658,N_9738);
nand U10199 (N_10199,N_9925,N_9605);
or U10200 (N_10200,N_9979,N_9603);
nand U10201 (N_10201,N_9865,N_9950);
or U10202 (N_10202,N_9522,N_9625);
and U10203 (N_10203,N_9842,N_9909);
nand U10204 (N_10204,N_9513,N_9521);
and U10205 (N_10205,N_9531,N_9762);
xnor U10206 (N_10206,N_9707,N_9756);
or U10207 (N_10207,N_9519,N_9806);
or U10208 (N_10208,N_9595,N_9644);
and U10209 (N_10209,N_9772,N_9763);
and U10210 (N_10210,N_9913,N_9689);
and U10211 (N_10211,N_9907,N_9937);
or U10212 (N_10212,N_9710,N_9915);
and U10213 (N_10213,N_9553,N_9890);
nor U10214 (N_10214,N_9659,N_9954);
nor U10215 (N_10215,N_9574,N_9894);
nor U10216 (N_10216,N_9730,N_9962);
and U10217 (N_10217,N_9914,N_9712);
nor U10218 (N_10218,N_9741,N_9529);
and U10219 (N_10219,N_9822,N_9523);
nand U10220 (N_10220,N_9798,N_9843);
or U10221 (N_10221,N_9611,N_9802);
nand U10222 (N_10222,N_9503,N_9889);
xnor U10223 (N_10223,N_9685,N_9597);
or U10224 (N_10224,N_9917,N_9735);
nor U10225 (N_10225,N_9715,N_9826);
and U10226 (N_10226,N_9883,N_9982);
or U10227 (N_10227,N_9717,N_9971);
xor U10228 (N_10228,N_9888,N_9748);
nand U10229 (N_10229,N_9998,N_9679);
and U10230 (N_10230,N_9550,N_9539);
and U10231 (N_10231,N_9901,N_9649);
and U10232 (N_10232,N_9928,N_9980);
xnor U10233 (N_10233,N_9933,N_9999);
or U10234 (N_10234,N_9561,N_9538);
xnor U10235 (N_10235,N_9926,N_9833);
or U10236 (N_10236,N_9737,N_9684);
and U10237 (N_10237,N_9666,N_9773);
and U10238 (N_10238,N_9509,N_9615);
nand U10239 (N_10239,N_9582,N_9701);
and U10240 (N_10240,N_9557,N_9564);
nand U10241 (N_10241,N_9949,N_9902);
and U10242 (N_10242,N_9840,N_9656);
nand U10243 (N_10243,N_9823,N_9621);
and U10244 (N_10244,N_9613,N_9973);
xor U10245 (N_10245,N_9969,N_9885);
nor U10246 (N_10246,N_9819,N_9992);
nor U10247 (N_10247,N_9927,N_9646);
nor U10248 (N_10248,N_9556,N_9565);
and U10249 (N_10249,N_9997,N_9686);
or U10250 (N_10250,N_9920,N_9679);
nand U10251 (N_10251,N_9921,N_9850);
and U10252 (N_10252,N_9570,N_9646);
or U10253 (N_10253,N_9725,N_9883);
nor U10254 (N_10254,N_9543,N_9520);
or U10255 (N_10255,N_9796,N_9955);
nor U10256 (N_10256,N_9860,N_9750);
nand U10257 (N_10257,N_9703,N_9643);
xnor U10258 (N_10258,N_9821,N_9718);
nor U10259 (N_10259,N_9794,N_9879);
and U10260 (N_10260,N_9744,N_9915);
or U10261 (N_10261,N_9797,N_9975);
or U10262 (N_10262,N_9642,N_9994);
nand U10263 (N_10263,N_9618,N_9923);
and U10264 (N_10264,N_9607,N_9975);
nand U10265 (N_10265,N_9576,N_9733);
xnor U10266 (N_10266,N_9610,N_9910);
or U10267 (N_10267,N_9988,N_9551);
xor U10268 (N_10268,N_9646,N_9580);
or U10269 (N_10269,N_9948,N_9648);
and U10270 (N_10270,N_9973,N_9854);
nand U10271 (N_10271,N_9950,N_9716);
nand U10272 (N_10272,N_9854,N_9738);
and U10273 (N_10273,N_9914,N_9689);
nand U10274 (N_10274,N_9689,N_9879);
nor U10275 (N_10275,N_9727,N_9901);
nor U10276 (N_10276,N_9972,N_9774);
nor U10277 (N_10277,N_9598,N_9595);
and U10278 (N_10278,N_9558,N_9544);
nand U10279 (N_10279,N_9543,N_9626);
nor U10280 (N_10280,N_9903,N_9769);
nor U10281 (N_10281,N_9508,N_9721);
or U10282 (N_10282,N_9551,N_9704);
nor U10283 (N_10283,N_9902,N_9955);
and U10284 (N_10284,N_9749,N_9600);
nand U10285 (N_10285,N_9750,N_9608);
nor U10286 (N_10286,N_9523,N_9851);
xnor U10287 (N_10287,N_9627,N_9613);
or U10288 (N_10288,N_9620,N_9697);
and U10289 (N_10289,N_9915,N_9595);
nor U10290 (N_10290,N_9587,N_9766);
nand U10291 (N_10291,N_9829,N_9669);
nand U10292 (N_10292,N_9504,N_9998);
and U10293 (N_10293,N_9842,N_9801);
nand U10294 (N_10294,N_9868,N_9879);
nor U10295 (N_10295,N_9570,N_9534);
nor U10296 (N_10296,N_9695,N_9866);
and U10297 (N_10297,N_9616,N_9566);
or U10298 (N_10298,N_9977,N_9531);
and U10299 (N_10299,N_9550,N_9701);
or U10300 (N_10300,N_9764,N_9700);
nor U10301 (N_10301,N_9985,N_9937);
or U10302 (N_10302,N_9841,N_9785);
and U10303 (N_10303,N_9513,N_9684);
nand U10304 (N_10304,N_9537,N_9604);
nand U10305 (N_10305,N_9834,N_9807);
nor U10306 (N_10306,N_9772,N_9744);
xnor U10307 (N_10307,N_9854,N_9835);
xnor U10308 (N_10308,N_9867,N_9736);
nand U10309 (N_10309,N_9656,N_9714);
or U10310 (N_10310,N_9995,N_9648);
or U10311 (N_10311,N_9503,N_9818);
or U10312 (N_10312,N_9556,N_9519);
xor U10313 (N_10313,N_9672,N_9656);
nor U10314 (N_10314,N_9647,N_9524);
or U10315 (N_10315,N_9542,N_9747);
nand U10316 (N_10316,N_9925,N_9931);
nor U10317 (N_10317,N_9897,N_9865);
nor U10318 (N_10318,N_9860,N_9654);
nor U10319 (N_10319,N_9863,N_9683);
or U10320 (N_10320,N_9561,N_9835);
or U10321 (N_10321,N_9726,N_9688);
nor U10322 (N_10322,N_9952,N_9625);
and U10323 (N_10323,N_9549,N_9721);
and U10324 (N_10324,N_9721,N_9735);
nand U10325 (N_10325,N_9910,N_9691);
nor U10326 (N_10326,N_9769,N_9711);
or U10327 (N_10327,N_9824,N_9688);
and U10328 (N_10328,N_9529,N_9900);
nor U10329 (N_10329,N_9906,N_9820);
and U10330 (N_10330,N_9973,N_9996);
and U10331 (N_10331,N_9586,N_9869);
nand U10332 (N_10332,N_9662,N_9895);
or U10333 (N_10333,N_9689,N_9886);
nor U10334 (N_10334,N_9553,N_9841);
nand U10335 (N_10335,N_9565,N_9983);
nand U10336 (N_10336,N_9526,N_9927);
xor U10337 (N_10337,N_9647,N_9678);
nor U10338 (N_10338,N_9647,N_9822);
xor U10339 (N_10339,N_9774,N_9891);
nand U10340 (N_10340,N_9917,N_9925);
nand U10341 (N_10341,N_9923,N_9528);
nand U10342 (N_10342,N_9816,N_9696);
or U10343 (N_10343,N_9832,N_9807);
or U10344 (N_10344,N_9547,N_9566);
or U10345 (N_10345,N_9548,N_9836);
nor U10346 (N_10346,N_9873,N_9596);
xor U10347 (N_10347,N_9578,N_9521);
nand U10348 (N_10348,N_9743,N_9769);
nor U10349 (N_10349,N_9917,N_9923);
xor U10350 (N_10350,N_9721,N_9594);
nand U10351 (N_10351,N_9584,N_9819);
nand U10352 (N_10352,N_9952,N_9510);
nand U10353 (N_10353,N_9833,N_9992);
nand U10354 (N_10354,N_9664,N_9835);
nand U10355 (N_10355,N_9804,N_9975);
or U10356 (N_10356,N_9524,N_9957);
xnor U10357 (N_10357,N_9789,N_9869);
xor U10358 (N_10358,N_9549,N_9613);
nor U10359 (N_10359,N_9984,N_9685);
nor U10360 (N_10360,N_9771,N_9974);
nor U10361 (N_10361,N_9704,N_9902);
nor U10362 (N_10362,N_9682,N_9605);
or U10363 (N_10363,N_9900,N_9584);
and U10364 (N_10364,N_9683,N_9914);
and U10365 (N_10365,N_9933,N_9603);
xnor U10366 (N_10366,N_9945,N_9968);
or U10367 (N_10367,N_9609,N_9520);
xnor U10368 (N_10368,N_9907,N_9680);
nor U10369 (N_10369,N_9837,N_9677);
or U10370 (N_10370,N_9657,N_9764);
or U10371 (N_10371,N_9841,N_9550);
nor U10372 (N_10372,N_9521,N_9635);
nor U10373 (N_10373,N_9860,N_9707);
nand U10374 (N_10374,N_9696,N_9920);
nor U10375 (N_10375,N_9994,N_9746);
or U10376 (N_10376,N_9787,N_9776);
and U10377 (N_10377,N_9783,N_9823);
nand U10378 (N_10378,N_9946,N_9625);
and U10379 (N_10379,N_9679,N_9724);
nor U10380 (N_10380,N_9577,N_9664);
or U10381 (N_10381,N_9926,N_9971);
and U10382 (N_10382,N_9624,N_9531);
nand U10383 (N_10383,N_9736,N_9927);
and U10384 (N_10384,N_9794,N_9587);
or U10385 (N_10385,N_9602,N_9869);
and U10386 (N_10386,N_9942,N_9615);
nand U10387 (N_10387,N_9698,N_9551);
xnor U10388 (N_10388,N_9772,N_9891);
and U10389 (N_10389,N_9543,N_9797);
nand U10390 (N_10390,N_9669,N_9645);
nand U10391 (N_10391,N_9569,N_9692);
or U10392 (N_10392,N_9793,N_9846);
nor U10393 (N_10393,N_9940,N_9949);
nor U10394 (N_10394,N_9782,N_9595);
xor U10395 (N_10395,N_9791,N_9713);
xnor U10396 (N_10396,N_9792,N_9508);
and U10397 (N_10397,N_9894,N_9996);
nand U10398 (N_10398,N_9539,N_9948);
nand U10399 (N_10399,N_9525,N_9670);
nand U10400 (N_10400,N_9684,N_9798);
nand U10401 (N_10401,N_9530,N_9584);
and U10402 (N_10402,N_9712,N_9913);
and U10403 (N_10403,N_9758,N_9861);
nand U10404 (N_10404,N_9763,N_9764);
or U10405 (N_10405,N_9744,N_9555);
nand U10406 (N_10406,N_9569,N_9537);
nor U10407 (N_10407,N_9889,N_9996);
nor U10408 (N_10408,N_9791,N_9658);
nand U10409 (N_10409,N_9564,N_9503);
nand U10410 (N_10410,N_9832,N_9540);
and U10411 (N_10411,N_9652,N_9799);
nor U10412 (N_10412,N_9511,N_9735);
and U10413 (N_10413,N_9919,N_9602);
nand U10414 (N_10414,N_9636,N_9536);
nor U10415 (N_10415,N_9561,N_9694);
and U10416 (N_10416,N_9587,N_9906);
xnor U10417 (N_10417,N_9835,N_9588);
and U10418 (N_10418,N_9720,N_9888);
and U10419 (N_10419,N_9844,N_9802);
nor U10420 (N_10420,N_9956,N_9826);
and U10421 (N_10421,N_9631,N_9977);
nor U10422 (N_10422,N_9715,N_9618);
nor U10423 (N_10423,N_9971,N_9930);
nor U10424 (N_10424,N_9859,N_9991);
and U10425 (N_10425,N_9880,N_9514);
nor U10426 (N_10426,N_9778,N_9579);
and U10427 (N_10427,N_9949,N_9628);
nand U10428 (N_10428,N_9846,N_9697);
nor U10429 (N_10429,N_9709,N_9783);
nand U10430 (N_10430,N_9789,N_9813);
nor U10431 (N_10431,N_9926,N_9894);
nand U10432 (N_10432,N_9945,N_9810);
and U10433 (N_10433,N_9944,N_9596);
nor U10434 (N_10434,N_9688,N_9861);
or U10435 (N_10435,N_9935,N_9727);
nor U10436 (N_10436,N_9884,N_9939);
xor U10437 (N_10437,N_9725,N_9955);
nor U10438 (N_10438,N_9515,N_9709);
nand U10439 (N_10439,N_9848,N_9637);
or U10440 (N_10440,N_9775,N_9562);
and U10441 (N_10441,N_9826,N_9936);
nor U10442 (N_10442,N_9892,N_9628);
xnor U10443 (N_10443,N_9521,N_9811);
or U10444 (N_10444,N_9903,N_9707);
xnor U10445 (N_10445,N_9906,N_9909);
and U10446 (N_10446,N_9950,N_9649);
or U10447 (N_10447,N_9610,N_9672);
and U10448 (N_10448,N_9717,N_9712);
and U10449 (N_10449,N_9818,N_9794);
xor U10450 (N_10450,N_9965,N_9691);
and U10451 (N_10451,N_9529,N_9867);
xnor U10452 (N_10452,N_9885,N_9703);
or U10453 (N_10453,N_9587,N_9702);
xnor U10454 (N_10454,N_9688,N_9505);
nor U10455 (N_10455,N_9629,N_9682);
nand U10456 (N_10456,N_9645,N_9828);
nor U10457 (N_10457,N_9668,N_9700);
and U10458 (N_10458,N_9880,N_9793);
or U10459 (N_10459,N_9561,N_9633);
nand U10460 (N_10460,N_9952,N_9902);
and U10461 (N_10461,N_9659,N_9583);
nor U10462 (N_10462,N_9904,N_9866);
and U10463 (N_10463,N_9761,N_9689);
nand U10464 (N_10464,N_9916,N_9767);
or U10465 (N_10465,N_9989,N_9619);
nand U10466 (N_10466,N_9565,N_9996);
nor U10467 (N_10467,N_9553,N_9659);
nand U10468 (N_10468,N_9966,N_9578);
nor U10469 (N_10469,N_9943,N_9894);
and U10470 (N_10470,N_9535,N_9981);
nor U10471 (N_10471,N_9929,N_9581);
nand U10472 (N_10472,N_9806,N_9750);
and U10473 (N_10473,N_9559,N_9788);
or U10474 (N_10474,N_9927,N_9596);
xor U10475 (N_10475,N_9634,N_9692);
nand U10476 (N_10476,N_9559,N_9700);
nand U10477 (N_10477,N_9750,N_9873);
xnor U10478 (N_10478,N_9984,N_9898);
or U10479 (N_10479,N_9984,N_9525);
and U10480 (N_10480,N_9712,N_9828);
xnor U10481 (N_10481,N_9556,N_9586);
or U10482 (N_10482,N_9747,N_9786);
or U10483 (N_10483,N_9926,N_9635);
nand U10484 (N_10484,N_9899,N_9618);
or U10485 (N_10485,N_9654,N_9914);
or U10486 (N_10486,N_9610,N_9740);
nor U10487 (N_10487,N_9874,N_9657);
xnor U10488 (N_10488,N_9586,N_9771);
nor U10489 (N_10489,N_9589,N_9970);
nand U10490 (N_10490,N_9671,N_9549);
xnor U10491 (N_10491,N_9943,N_9658);
and U10492 (N_10492,N_9661,N_9924);
nor U10493 (N_10493,N_9529,N_9892);
nand U10494 (N_10494,N_9826,N_9552);
nand U10495 (N_10495,N_9727,N_9697);
or U10496 (N_10496,N_9990,N_9645);
and U10497 (N_10497,N_9538,N_9548);
xor U10498 (N_10498,N_9865,N_9551);
and U10499 (N_10499,N_9838,N_9872);
nor U10500 (N_10500,N_10051,N_10371);
nor U10501 (N_10501,N_10482,N_10152);
or U10502 (N_10502,N_10093,N_10346);
or U10503 (N_10503,N_10187,N_10415);
nand U10504 (N_10504,N_10144,N_10169);
or U10505 (N_10505,N_10108,N_10357);
and U10506 (N_10506,N_10210,N_10280);
xor U10507 (N_10507,N_10476,N_10390);
nor U10508 (N_10508,N_10286,N_10030);
and U10509 (N_10509,N_10356,N_10201);
and U10510 (N_10510,N_10024,N_10004);
nand U10511 (N_10511,N_10066,N_10250);
or U10512 (N_10512,N_10011,N_10150);
nand U10513 (N_10513,N_10039,N_10479);
and U10514 (N_10514,N_10236,N_10249);
nand U10515 (N_10515,N_10370,N_10406);
or U10516 (N_10516,N_10361,N_10025);
or U10517 (N_10517,N_10149,N_10257);
nand U10518 (N_10518,N_10450,N_10486);
and U10519 (N_10519,N_10104,N_10261);
and U10520 (N_10520,N_10168,N_10422);
nand U10521 (N_10521,N_10136,N_10074);
nor U10522 (N_10522,N_10113,N_10192);
and U10523 (N_10523,N_10252,N_10374);
and U10524 (N_10524,N_10159,N_10239);
nand U10525 (N_10525,N_10404,N_10491);
nor U10526 (N_10526,N_10134,N_10148);
or U10527 (N_10527,N_10449,N_10340);
and U10528 (N_10528,N_10322,N_10133);
or U10529 (N_10529,N_10446,N_10130);
nand U10530 (N_10530,N_10316,N_10142);
or U10531 (N_10531,N_10348,N_10463);
nand U10532 (N_10532,N_10445,N_10345);
or U10533 (N_10533,N_10427,N_10253);
nor U10534 (N_10534,N_10031,N_10398);
or U10535 (N_10535,N_10315,N_10305);
xor U10536 (N_10536,N_10421,N_10010);
nand U10537 (N_10537,N_10197,N_10483);
or U10538 (N_10538,N_10419,N_10181);
or U10539 (N_10539,N_10417,N_10269);
nor U10540 (N_10540,N_10060,N_10441);
nor U10541 (N_10541,N_10347,N_10349);
and U10542 (N_10542,N_10260,N_10414);
xor U10543 (N_10543,N_10376,N_10462);
nor U10544 (N_10544,N_10412,N_10467);
nor U10545 (N_10545,N_10333,N_10175);
nor U10546 (N_10546,N_10151,N_10433);
nand U10547 (N_10547,N_10383,N_10284);
xnor U10548 (N_10548,N_10258,N_10331);
xnor U10549 (N_10549,N_10254,N_10232);
nand U10550 (N_10550,N_10263,N_10003);
nand U10551 (N_10551,N_10439,N_10082);
nand U10552 (N_10552,N_10460,N_10382);
xor U10553 (N_10553,N_10309,N_10073);
xnor U10554 (N_10554,N_10396,N_10381);
and U10555 (N_10555,N_10155,N_10310);
nor U10556 (N_10556,N_10424,N_10283);
or U10557 (N_10557,N_10163,N_10369);
nand U10558 (N_10558,N_10496,N_10266);
and U10559 (N_10559,N_10362,N_10043);
and U10560 (N_10560,N_10360,N_10437);
nor U10561 (N_10561,N_10470,N_10117);
nor U10562 (N_10562,N_10296,N_10202);
xor U10563 (N_10563,N_10455,N_10337);
nor U10564 (N_10564,N_10375,N_10311);
nor U10565 (N_10565,N_10457,N_10365);
or U10566 (N_10566,N_10265,N_10044);
nor U10567 (N_10567,N_10246,N_10292);
or U10568 (N_10568,N_10240,N_10288);
and U10569 (N_10569,N_10314,N_10334);
nor U10570 (N_10570,N_10139,N_10056);
or U10571 (N_10571,N_10154,N_10129);
nand U10572 (N_10572,N_10222,N_10173);
xor U10573 (N_10573,N_10198,N_10141);
and U10574 (N_10574,N_10488,N_10057);
or U10575 (N_10575,N_10413,N_10330);
and U10576 (N_10576,N_10058,N_10015);
and U10577 (N_10577,N_10268,N_10461);
and U10578 (N_10578,N_10220,N_10022);
nand U10579 (N_10579,N_10072,N_10095);
and U10580 (N_10580,N_10456,N_10402);
xnor U10581 (N_10581,N_10059,N_10238);
nand U10582 (N_10582,N_10270,N_10050);
xor U10583 (N_10583,N_10124,N_10205);
and U10584 (N_10584,N_10090,N_10185);
nor U10585 (N_10585,N_10013,N_10420);
or U10586 (N_10586,N_10126,N_10326);
nand U10587 (N_10587,N_10318,N_10490);
nand U10588 (N_10588,N_10400,N_10217);
or U10589 (N_10589,N_10418,N_10076);
nand U10590 (N_10590,N_10243,N_10285);
or U10591 (N_10591,N_10392,N_10435);
or U10592 (N_10592,N_10489,N_10196);
nand U10593 (N_10593,N_10171,N_10123);
nor U10594 (N_10594,N_10017,N_10294);
and U10595 (N_10595,N_10353,N_10247);
and U10596 (N_10596,N_10293,N_10453);
nand U10597 (N_10597,N_10048,N_10191);
nor U10598 (N_10598,N_10193,N_10298);
and U10599 (N_10599,N_10399,N_10194);
xnor U10600 (N_10600,N_10306,N_10475);
and U10601 (N_10601,N_10068,N_10052);
or U10602 (N_10602,N_10209,N_10484);
nand U10603 (N_10603,N_10276,N_10344);
and U10604 (N_10604,N_10228,N_10046);
nor U10605 (N_10605,N_10237,N_10227);
and U10606 (N_10606,N_10067,N_10105);
or U10607 (N_10607,N_10352,N_10018);
or U10608 (N_10608,N_10308,N_10324);
or U10609 (N_10609,N_10065,N_10119);
xor U10610 (N_10610,N_10416,N_10211);
or U10611 (N_10611,N_10341,N_10230);
or U10612 (N_10612,N_10471,N_10103);
nor U10613 (N_10613,N_10387,N_10055);
or U10614 (N_10614,N_10442,N_10088);
nand U10615 (N_10615,N_10397,N_10303);
nor U10616 (N_10616,N_10028,N_10170);
and U10617 (N_10617,N_10302,N_10367);
and U10618 (N_10618,N_10190,N_10118);
and U10619 (N_10619,N_10325,N_10338);
or U10620 (N_10620,N_10447,N_10388);
nor U10621 (N_10621,N_10213,N_10493);
xnor U10622 (N_10622,N_10177,N_10156);
or U10623 (N_10623,N_10206,N_10101);
xnor U10624 (N_10624,N_10212,N_10135);
nand U10625 (N_10625,N_10062,N_10287);
or U10626 (N_10626,N_10328,N_10221);
xnor U10627 (N_10627,N_10351,N_10497);
xnor U10628 (N_10628,N_10234,N_10033);
xor U10629 (N_10629,N_10029,N_10452);
nor U10630 (N_10630,N_10224,N_10146);
nand U10631 (N_10631,N_10120,N_10323);
and U10632 (N_10632,N_10219,N_10458);
and U10633 (N_10633,N_10373,N_10279);
nor U10634 (N_10634,N_10278,N_10026);
nor U10635 (N_10635,N_10480,N_10016);
or U10636 (N_10636,N_10186,N_10495);
and U10637 (N_10637,N_10248,N_10203);
nand U10638 (N_10638,N_10317,N_10273);
nor U10639 (N_10639,N_10385,N_10207);
and U10640 (N_10640,N_10157,N_10372);
and U10641 (N_10641,N_10121,N_10165);
nand U10642 (N_10642,N_10436,N_10199);
and U10643 (N_10643,N_10299,N_10454);
nor U10644 (N_10644,N_10083,N_10231);
nand U10645 (N_10645,N_10423,N_10487);
xnor U10646 (N_10646,N_10478,N_10368);
xnor U10647 (N_10647,N_10393,N_10377);
nor U10648 (N_10648,N_10301,N_10131);
xnor U10649 (N_10649,N_10354,N_10140);
nand U10650 (N_10650,N_10184,N_10320);
or U10651 (N_10651,N_10332,N_10096);
and U10652 (N_10652,N_10077,N_10465);
and U10653 (N_10653,N_10091,N_10327);
nor U10654 (N_10654,N_10178,N_10106);
or U10655 (N_10655,N_10242,N_10380);
xnor U10656 (N_10656,N_10366,N_10176);
nor U10657 (N_10657,N_10100,N_10473);
nor U10658 (N_10658,N_10281,N_10045);
or U10659 (N_10659,N_10038,N_10034);
nand U10660 (N_10660,N_10053,N_10443);
or U10661 (N_10661,N_10429,N_10023);
and U10662 (N_10662,N_10425,N_10407);
nor U10663 (N_10663,N_10438,N_10343);
nand U10664 (N_10664,N_10251,N_10160);
or U10665 (N_10665,N_10054,N_10000);
xnor U10666 (N_10666,N_10071,N_10291);
xnor U10667 (N_10667,N_10122,N_10092);
nand U10668 (N_10668,N_10075,N_10342);
xor U10669 (N_10669,N_10401,N_10114);
nor U10670 (N_10670,N_10289,N_10085);
nor U10671 (N_10671,N_10395,N_10432);
nand U10672 (N_10672,N_10115,N_10485);
and U10673 (N_10673,N_10218,N_10262);
nand U10674 (N_10674,N_10014,N_10183);
and U10675 (N_10675,N_10007,N_10020);
and U10676 (N_10676,N_10182,N_10472);
nor U10677 (N_10677,N_10125,N_10127);
or U10678 (N_10678,N_10403,N_10180);
nor U10679 (N_10679,N_10027,N_10440);
nor U10680 (N_10680,N_10070,N_10408);
nand U10681 (N_10681,N_10492,N_10110);
nand U10682 (N_10682,N_10195,N_10215);
and U10683 (N_10683,N_10112,N_10319);
or U10684 (N_10684,N_10132,N_10109);
or U10685 (N_10685,N_10275,N_10295);
nor U10686 (N_10686,N_10459,N_10267);
xor U10687 (N_10687,N_10047,N_10204);
and U10688 (N_10688,N_10097,N_10081);
nor U10689 (N_10689,N_10235,N_10179);
and U10690 (N_10690,N_10259,N_10255);
or U10691 (N_10691,N_10087,N_10256);
or U10692 (N_10692,N_10312,N_10145);
nor U10693 (N_10693,N_10498,N_10386);
or U10694 (N_10694,N_10188,N_10200);
nand U10695 (N_10695,N_10138,N_10005);
nand U10696 (N_10696,N_10158,N_10474);
nand U10697 (N_10697,N_10008,N_10431);
nor U10698 (N_10698,N_10464,N_10061);
xor U10699 (N_10699,N_10094,N_10389);
xnor U10700 (N_10700,N_10321,N_10174);
xnor U10701 (N_10701,N_10336,N_10107);
xor U10702 (N_10702,N_10297,N_10379);
and U10703 (N_10703,N_10147,N_10358);
nor U10704 (N_10704,N_10078,N_10378);
xnor U10705 (N_10705,N_10064,N_10102);
nand U10706 (N_10706,N_10272,N_10116);
and U10707 (N_10707,N_10189,N_10290);
xor U10708 (N_10708,N_10006,N_10428);
nand U10709 (N_10709,N_10477,N_10079);
and U10710 (N_10710,N_10244,N_10274);
nand U10711 (N_10711,N_10019,N_10271);
xnor U10712 (N_10712,N_10098,N_10335);
nand U10713 (N_10713,N_10499,N_10434);
or U10714 (N_10714,N_10063,N_10405);
or U10715 (N_10715,N_10128,N_10245);
nor U10716 (N_10716,N_10069,N_10037);
and U10717 (N_10717,N_10042,N_10430);
or U10718 (N_10718,N_10099,N_10161);
xnor U10719 (N_10719,N_10313,N_10214);
or U10720 (N_10720,N_10223,N_10277);
or U10721 (N_10721,N_10300,N_10359);
or U10722 (N_10722,N_10350,N_10084);
and U10723 (N_10723,N_10167,N_10329);
nor U10724 (N_10724,N_10229,N_10089);
xor U10725 (N_10725,N_10032,N_10282);
nor U10726 (N_10726,N_10384,N_10012);
nor U10727 (N_10727,N_10494,N_10241);
nand U10728 (N_10728,N_10021,N_10009);
nor U10729 (N_10729,N_10307,N_10172);
nand U10730 (N_10730,N_10137,N_10394);
and U10731 (N_10731,N_10035,N_10002);
and U10732 (N_10732,N_10216,N_10451);
nand U10733 (N_10733,N_10264,N_10041);
or U10734 (N_10734,N_10355,N_10409);
or U10735 (N_10735,N_10426,N_10049);
and U10736 (N_10736,N_10410,N_10226);
and U10737 (N_10737,N_10466,N_10469);
and U10738 (N_10738,N_10364,N_10040);
nand U10739 (N_10739,N_10086,N_10411);
and U10740 (N_10740,N_10225,N_10153);
or U10741 (N_10741,N_10111,N_10448);
nand U10742 (N_10742,N_10444,N_10304);
nand U10743 (N_10743,N_10391,N_10164);
nand U10744 (N_10744,N_10339,N_10001);
xor U10745 (N_10745,N_10481,N_10363);
nand U10746 (N_10746,N_10143,N_10036);
nor U10747 (N_10747,N_10166,N_10208);
and U10748 (N_10748,N_10468,N_10080);
nand U10749 (N_10749,N_10233,N_10162);
or U10750 (N_10750,N_10365,N_10148);
nor U10751 (N_10751,N_10116,N_10174);
and U10752 (N_10752,N_10317,N_10288);
nor U10753 (N_10753,N_10071,N_10454);
and U10754 (N_10754,N_10332,N_10302);
xnor U10755 (N_10755,N_10410,N_10030);
nand U10756 (N_10756,N_10496,N_10008);
or U10757 (N_10757,N_10198,N_10109);
nor U10758 (N_10758,N_10487,N_10183);
or U10759 (N_10759,N_10352,N_10138);
or U10760 (N_10760,N_10365,N_10175);
or U10761 (N_10761,N_10368,N_10342);
and U10762 (N_10762,N_10110,N_10207);
nor U10763 (N_10763,N_10113,N_10303);
nand U10764 (N_10764,N_10042,N_10088);
nand U10765 (N_10765,N_10324,N_10245);
and U10766 (N_10766,N_10343,N_10234);
and U10767 (N_10767,N_10455,N_10489);
nand U10768 (N_10768,N_10484,N_10267);
and U10769 (N_10769,N_10327,N_10226);
or U10770 (N_10770,N_10452,N_10431);
nor U10771 (N_10771,N_10019,N_10146);
or U10772 (N_10772,N_10049,N_10277);
and U10773 (N_10773,N_10188,N_10150);
or U10774 (N_10774,N_10196,N_10422);
or U10775 (N_10775,N_10270,N_10045);
and U10776 (N_10776,N_10033,N_10013);
nor U10777 (N_10777,N_10123,N_10055);
nor U10778 (N_10778,N_10471,N_10308);
or U10779 (N_10779,N_10155,N_10446);
xor U10780 (N_10780,N_10220,N_10272);
nor U10781 (N_10781,N_10000,N_10382);
nor U10782 (N_10782,N_10117,N_10346);
nor U10783 (N_10783,N_10214,N_10368);
or U10784 (N_10784,N_10238,N_10287);
and U10785 (N_10785,N_10002,N_10058);
or U10786 (N_10786,N_10006,N_10188);
xor U10787 (N_10787,N_10301,N_10360);
nor U10788 (N_10788,N_10273,N_10298);
and U10789 (N_10789,N_10214,N_10201);
or U10790 (N_10790,N_10401,N_10282);
nor U10791 (N_10791,N_10065,N_10150);
and U10792 (N_10792,N_10364,N_10457);
or U10793 (N_10793,N_10377,N_10171);
nor U10794 (N_10794,N_10405,N_10089);
and U10795 (N_10795,N_10053,N_10241);
or U10796 (N_10796,N_10257,N_10440);
nor U10797 (N_10797,N_10142,N_10061);
nand U10798 (N_10798,N_10485,N_10269);
and U10799 (N_10799,N_10332,N_10117);
nor U10800 (N_10800,N_10281,N_10416);
or U10801 (N_10801,N_10126,N_10318);
nand U10802 (N_10802,N_10482,N_10288);
xnor U10803 (N_10803,N_10040,N_10181);
xnor U10804 (N_10804,N_10205,N_10244);
nor U10805 (N_10805,N_10161,N_10122);
nor U10806 (N_10806,N_10195,N_10250);
nor U10807 (N_10807,N_10339,N_10085);
or U10808 (N_10808,N_10184,N_10014);
and U10809 (N_10809,N_10283,N_10041);
nor U10810 (N_10810,N_10205,N_10263);
or U10811 (N_10811,N_10247,N_10421);
or U10812 (N_10812,N_10469,N_10037);
nand U10813 (N_10813,N_10468,N_10405);
nand U10814 (N_10814,N_10137,N_10450);
and U10815 (N_10815,N_10242,N_10361);
nand U10816 (N_10816,N_10420,N_10254);
or U10817 (N_10817,N_10347,N_10490);
nor U10818 (N_10818,N_10192,N_10085);
nor U10819 (N_10819,N_10066,N_10409);
nand U10820 (N_10820,N_10108,N_10280);
and U10821 (N_10821,N_10452,N_10379);
nand U10822 (N_10822,N_10383,N_10135);
nand U10823 (N_10823,N_10024,N_10445);
or U10824 (N_10824,N_10125,N_10485);
nor U10825 (N_10825,N_10396,N_10171);
and U10826 (N_10826,N_10098,N_10185);
and U10827 (N_10827,N_10189,N_10171);
or U10828 (N_10828,N_10323,N_10006);
and U10829 (N_10829,N_10188,N_10398);
nor U10830 (N_10830,N_10397,N_10458);
nand U10831 (N_10831,N_10178,N_10410);
and U10832 (N_10832,N_10240,N_10060);
or U10833 (N_10833,N_10022,N_10166);
nor U10834 (N_10834,N_10197,N_10332);
nand U10835 (N_10835,N_10034,N_10493);
nand U10836 (N_10836,N_10117,N_10064);
nor U10837 (N_10837,N_10130,N_10023);
nor U10838 (N_10838,N_10367,N_10115);
nor U10839 (N_10839,N_10018,N_10157);
or U10840 (N_10840,N_10002,N_10425);
and U10841 (N_10841,N_10305,N_10279);
nand U10842 (N_10842,N_10439,N_10271);
xnor U10843 (N_10843,N_10349,N_10431);
nor U10844 (N_10844,N_10023,N_10140);
or U10845 (N_10845,N_10224,N_10360);
xor U10846 (N_10846,N_10472,N_10369);
and U10847 (N_10847,N_10349,N_10201);
nor U10848 (N_10848,N_10170,N_10275);
nand U10849 (N_10849,N_10086,N_10481);
nor U10850 (N_10850,N_10029,N_10359);
nor U10851 (N_10851,N_10029,N_10102);
xnor U10852 (N_10852,N_10375,N_10267);
or U10853 (N_10853,N_10412,N_10478);
or U10854 (N_10854,N_10182,N_10262);
nand U10855 (N_10855,N_10393,N_10275);
nand U10856 (N_10856,N_10276,N_10000);
nand U10857 (N_10857,N_10113,N_10204);
xnor U10858 (N_10858,N_10429,N_10019);
xnor U10859 (N_10859,N_10332,N_10023);
nand U10860 (N_10860,N_10437,N_10426);
or U10861 (N_10861,N_10017,N_10470);
nand U10862 (N_10862,N_10305,N_10120);
and U10863 (N_10863,N_10321,N_10176);
nor U10864 (N_10864,N_10360,N_10403);
nand U10865 (N_10865,N_10202,N_10323);
or U10866 (N_10866,N_10459,N_10056);
and U10867 (N_10867,N_10341,N_10050);
and U10868 (N_10868,N_10466,N_10477);
or U10869 (N_10869,N_10402,N_10261);
and U10870 (N_10870,N_10368,N_10422);
nor U10871 (N_10871,N_10264,N_10062);
nor U10872 (N_10872,N_10263,N_10009);
nor U10873 (N_10873,N_10274,N_10337);
or U10874 (N_10874,N_10065,N_10293);
nand U10875 (N_10875,N_10025,N_10026);
xnor U10876 (N_10876,N_10339,N_10254);
and U10877 (N_10877,N_10430,N_10358);
and U10878 (N_10878,N_10474,N_10257);
or U10879 (N_10879,N_10004,N_10256);
nand U10880 (N_10880,N_10169,N_10250);
nor U10881 (N_10881,N_10376,N_10394);
nor U10882 (N_10882,N_10180,N_10258);
or U10883 (N_10883,N_10463,N_10450);
nor U10884 (N_10884,N_10145,N_10442);
or U10885 (N_10885,N_10048,N_10420);
and U10886 (N_10886,N_10014,N_10457);
and U10887 (N_10887,N_10147,N_10229);
and U10888 (N_10888,N_10385,N_10029);
nand U10889 (N_10889,N_10235,N_10295);
or U10890 (N_10890,N_10104,N_10149);
or U10891 (N_10891,N_10301,N_10353);
nor U10892 (N_10892,N_10203,N_10000);
and U10893 (N_10893,N_10256,N_10394);
nand U10894 (N_10894,N_10357,N_10181);
nand U10895 (N_10895,N_10051,N_10003);
and U10896 (N_10896,N_10350,N_10115);
or U10897 (N_10897,N_10216,N_10302);
nor U10898 (N_10898,N_10329,N_10452);
and U10899 (N_10899,N_10179,N_10114);
nand U10900 (N_10900,N_10395,N_10365);
xor U10901 (N_10901,N_10223,N_10352);
nor U10902 (N_10902,N_10347,N_10043);
and U10903 (N_10903,N_10205,N_10272);
or U10904 (N_10904,N_10294,N_10422);
nand U10905 (N_10905,N_10416,N_10013);
nand U10906 (N_10906,N_10253,N_10274);
nand U10907 (N_10907,N_10333,N_10048);
nand U10908 (N_10908,N_10453,N_10071);
and U10909 (N_10909,N_10261,N_10111);
nand U10910 (N_10910,N_10348,N_10391);
nand U10911 (N_10911,N_10473,N_10340);
and U10912 (N_10912,N_10431,N_10412);
nand U10913 (N_10913,N_10054,N_10402);
nand U10914 (N_10914,N_10060,N_10348);
and U10915 (N_10915,N_10360,N_10479);
and U10916 (N_10916,N_10314,N_10184);
nor U10917 (N_10917,N_10098,N_10102);
and U10918 (N_10918,N_10377,N_10038);
or U10919 (N_10919,N_10451,N_10362);
xor U10920 (N_10920,N_10212,N_10053);
and U10921 (N_10921,N_10349,N_10351);
or U10922 (N_10922,N_10090,N_10370);
and U10923 (N_10923,N_10170,N_10119);
nor U10924 (N_10924,N_10348,N_10169);
and U10925 (N_10925,N_10457,N_10179);
nand U10926 (N_10926,N_10471,N_10174);
or U10927 (N_10927,N_10452,N_10050);
nand U10928 (N_10928,N_10254,N_10428);
nor U10929 (N_10929,N_10389,N_10464);
xor U10930 (N_10930,N_10297,N_10291);
and U10931 (N_10931,N_10329,N_10206);
and U10932 (N_10932,N_10233,N_10130);
nand U10933 (N_10933,N_10394,N_10293);
or U10934 (N_10934,N_10349,N_10094);
nor U10935 (N_10935,N_10131,N_10121);
nor U10936 (N_10936,N_10061,N_10492);
nand U10937 (N_10937,N_10073,N_10162);
nand U10938 (N_10938,N_10264,N_10147);
or U10939 (N_10939,N_10108,N_10492);
nor U10940 (N_10940,N_10277,N_10144);
nor U10941 (N_10941,N_10477,N_10339);
and U10942 (N_10942,N_10157,N_10418);
and U10943 (N_10943,N_10488,N_10216);
and U10944 (N_10944,N_10337,N_10298);
nor U10945 (N_10945,N_10299,N_10345);
and U10946 (N_10946,N_10120,N_10041);
nor U10947 (N_10947,N_10401,N_10336);
and U10948 (N_10948,N_10247,N_10280);
and U10949 (N_10949,N_10408,N_10046);
nand U10950 (N_10950,N_10414,N_10374);
nand U10951 (N_10951,N_10195,N_10387);
or U10952 (N_10952,N_10239,N_10294);
and U10953 (N_10953,N_10301,N_10148);
and U10954 (N_10954,N_10231,N_10008);
or U10955 (N_10955,N_10476,N_10012);
nand U10956 (N_10956,N_10403,N_10011);
nand U10957 (N_10957,N_10344,N_10498);
xor U10958 (N_10958,N_10069,N_10292);
and U10959 (N_10959,N_10190,N_10320);
nand U10960 (N_10960,N_10397,N_10437);
nand U10961 (N_10961,N_10022,N_10157);
nand U10962 (N_10962,N_10148,N_10443);
and U10963 (N_10963,N_10038,N_10232);
nor U10964 (N_10964,N_10442,N_10450);
nand U10965 (N_10965,N_10213,N_10365);
nor U10966 (N_10966,N_10045,N_10389);
nand U10967 (N_10967,N_10358,N_10155);
nor U10968 (N_10968,N_10373,N_10393);
and U10969 (N_10969,N_10433,N_10065);
and U10970 (N_10970,N_10252,N_10236);
and U10971 (N_10971,N_10477,N_10454);
nand U10972 (N_10972,N_10146,N_10318);
nor U10973 (N_10973,N_10206,N_10188);
or U10974 (N_10974,N_10357,N_10271);
or U10975 (N_10975,N_10051,N_10015);
nand U10976 (N_10976,N_10085,N_10127);
nand U10977 (N_10977,N_10457,N_10382);
nand U10978 (N_10978,N_10301,N_10129);
nor U10979 (N_10979,N_10389,N_10329);
nand U10980 (N_10980,N_10495,N_10491);
nand U10981 (N_10981,N_10255,N_10399);
nor U10982 (N_10982,N_10048,N_10334);
or U10983 (N_10983,N_10258,N_10398);
or U10984 (N_10984,N_10307,N_10116);
or U10985 (N_10985,N_10145,N_10389);
nor U10986 (N_10986,N_10352,N_10243);
nand U10987 (N_10987,N_10325,N_10198);
xor U10988 (N_10988,N_10253,N_10083);
nand U10989 (N_10989,N_10147,N_10173);
and U10990 (N_10990,N_10120,N_10409);
and U10991 (N_10991,N_10307,N_10194);
and U10992 (N_10992,N_10477,N_10102);
nand U10993 (N_10993,N_10450,N_10174);
nor U10994 (N_10994,N_10496,N_10020);
or U10995 (N_10995,N_10370,N_10403);
or U10996 (N_10996,N_10429,N_10295);
nand U10997 (N_10997,N_10143,N_10472);
nand U10998 (N_10998,N_10174,N_10148);
nor U10999 (N_10999,N_10105,N_10374);
and U11000 (N_11000,N_10950,N_10972);
or U11001 (N_11001,N_10593,N_10982);
nor U11002 (N_11002,N_10561,N_10869);
nand U11003 (N_11003,N_10526,N_10709);
nor U11004 (N_11004,N_10753,N_10796);
nand U11005 (N_11005,N_10559,N_10856);
nor U11006 (N_11006,N_10900,N_10532);
or U11007 (N_11007,N_10562,N_10914);
nor U11008 (N_11008,N_10953,N_10851);
and U11009 (N_11009,N_10588,N_10614);
and U11010 (N_11010,N_10591,N_10874);
nor U11011 (N_11011,N_10963,N_10902);
and U11012 (N_11012,N_10512,N_10955);
nand U11013 (N_11013,N_10524,N_10701);
nor U11014 (N_11014,N_10633,N_10766);
nor U11015 (N_11015,N_10711,N_10924);
nor U11016 (N_11016,N_10975,N_10678);
xor U11017 (N_11017,N_10626,N_10605);
xnor U11018 (N_11018,N_10739,N_10745);
nand U11019 (N_11019,N_10927,N_10871);
and U11020 (N_11020,N_10821,N_10572);
and U11021 (N_11021,N_10835,N_10989);
nor U11022 (N_11022,N_10746,N_10732);
or U11023 (N_11023,N_10798,N_10813);
nor U11024 (N_11024,N_10945,N_10685);
or U11025 (N_11025,N_10901,N_10954);
and U11026 (N_11026,N_10899,N_10819);
or U11027 (N_11027,N_10519,N_10878);
nand U11028 (N_11028,N_10543,N_10662);
nand U11029 (N_11029,N_10647,N_10848);
nand U11030 (N_11030,N_10707,N_10979);
and U11031 (N_11031,N_10797,N_10580);
and U11032 (N_11032,N_10781,N_10959);
and U11033 (N_11033,N_10875,N_10536);
and U11034 (N_11034,N_10936,N_10836);
or U11035 (N_11035,N_10585,N_10940);
nor U11036 (N_11036,N_10552,N_10834);
nand U11037 (N_11037,N_10948,N_10513);
and U11038 (N_11038,N_10557,N_10671);
xnor U11039 (N_11039,N_10812,N_10511);
or U11040 (N_11040,N_10713,N_10844);
and U11041 (N_11041,N_10853,N_10715);
nand U11042 (N_11042,N_10584,N_10547);
or U11043 (N_11043,N_10544,N_10699);
nand U11044 (N_11044,N_10700,N_10674);
or U11045 (N_11045,N_10981,N_10517);
nand U11046 (N_11046,N_10968,N_10632);
or U11047 (N_11047,N_10749,N_10799);
and U11048 (N_11048,N_10722,N_10931);
xor U11049 (N_11049,N_10881,N_10655);
and U11050 (N_11050,N_10560,N_10672);
and U11051 (N_11051,N_10744,N_10658);
nor U11052 (N_11052,N_10860,N_10758);
nor U11053 (N_11053,N_10503,N_10993);
and U11054 (N_11054,N_10515,N_10542);
nor U11055 (N_11055,N_10780,N_10965);
nand U11056 (N_11056,N_10582,N_10811);
or U11057 (N_11057,N_10830,N_10857);
or U11058 (N_11058,N_10618,N_10586);
nand U11059 (N_11059,N_10608,N_10828);
nor U11060 (N_11060,N_10894,N_10870);
nand U11061 (N_11061,N_10790,N_10666);
and U11062 (N_11062,N_10977,N_10535);
nor U11063 (N_11063,N_10641,N_10842);
and U11064 (N_11064,N_10893,N_10778);
nor U11065 (N_11065,N_10521,N_10695);
and U11066 (N_11066,N_10733,N_10533);
nor U11067 (N_11067,N_10809,N_10509);
and U11068 (N_11068,N_10537,N_10643);
and U11069 (N_11069,N_10941,N_10917);
nand U11070 (N_11070,N_10723,N_10958);
and U11071 (N_11071,N_10570,N_10861);
or U11072 (N_11072,N_10620,N_10508);
and U11073 (N_11073,N_10974,N_10743);
xnor U11074 (N_11074,N_10802,N_10872);
xnor U11075 (N_11075,N_10938,N_10852);
xnor U11076 (N_11076,N_10676,N_10581);
nand U11077 (N_11077,N_10688,N_10908);
and U11078 (N_11078,N_10510,N_10539);
xnor U11079 (N_11079,N_10976,N_10742);
and U11080 (N_11080,N_10642,N_10995);
xor U11081 (N_11081,N_10529,N_10998);
nor U11082 (N_11082,N_10978,N_10661);
nand U11083 (N_11083,N_10776,N_10578);
or U11084 (N_11084,N_10670,N_10720);
and U11085 (N_11085,N_10657,N_10841);
nand U11086 (N_11086,N_10712,N_10845);
nand U11087 (N_11087,N_10747,N_10736);
and U11088 (N_11088,N_10971,N_10592);
and U11089 (N_11089,N_10530,N_10942);
or U11090 (N_11090,N_10823,N_10805);
nor U11091 (N_11091,N_10926,N_10752);
nand U11092 (N_11092,N_10506,N_10595);
or U11093 (N_11093,N_10889,N_10849);
nand U11094 (N_11094,N_10859,N_10854);
nand U11095 (N_11095,N_10627,N_10654);
nor U11096 (N_11096,N_10935,N_10846);
or U11097 (N_11097,N_10531,N_10630);
or U11098 (N_11098,N_10667,N_10516);
or U11099 (N_11099,N_10691,N_10615);
nand U11100 (N_11100,N_10703,N_10887);
nor U11101 (N_11101,N_10782,N_10577);
nor U11102 (N_11102,N_10864,N_10690);
nor U11103 (N_11103,N_10774,N_10748);
xor U11104 (N_11104,N_10788,N_10787);
nor U11105 (N_11105,N_10610,N_10818);
and U11106 (N_11106,N_10937,N_10684);
or U11107 (N_11107,N_10612,N_10760);
nor U11108 (N_11108,N_10567,N_10505);
nor U11109 (N_11109,N_10741,N_10645);
and U11110 (N_11110,N_10772,N_10716);
and U11111 (N_11111,N_10984,N_10879);
and U11112 (N_11112,N_10946,N_10952);
and U11113 (N_11113,N_10623,N_10957);
or U11114 (N_11114,N_10783,N_10761);
nand U11115 (N_11115,N_10980,N_10934);
nand U11116 (N_11116,N_10682,N_10599);
and U11117 (N_11117,N_10904,N_10502);
and U11118 (N_11118,N_10563,N_10922);
xnor U11119 (N_11119,N_10644,N_10966);
nor U11120 (N_11120,N_10525,N_10576);
and U11121 (N_11121,N_10564,N_10669);
or U11122 (N_11122,N_10737,N_10652);
nand U11123 (N_11123,N_10762,N_10890);
nand U11124 (N_11124,N_10726,N_10597);
xnor U11125 (N_11125,N_10913,N_10873);
nor U11126 (N_11126,N_10755,N_10640);
nand U11127 (N_11127,N_10696,N_10888);
or U11128 (N_11128,N_10858,N_10613);
or U11129 (N_11129,N_10656,N_10628);
nor U11130 (N_11130,N_10638,N_10680);
and U11131 (N_11131,N_10912,N_10837);
nand U11132 (N_11132,N_10629,N_10565);
xnor U11133 (N_11133,N_10631,N_10994);
and U11134 (N_11134,N_10867,N_10863);
nor U11135 (N_11135,N_10768,N_10636);
and U11136 (N_11136,N_10775,N_10718);
or U11137 (N_11137,N_10735,N_10579);
or U11138 (N_11138,N_10897,N_10569);
or U11139 (N_11139,N_10639,N_10754);
nand U11140 (N_11140,N_10619,N_10725);
or U11141 (N_11141,N_10587,N_10604);
xor U11142 (N_11142,N_10548,N_10815);
and U11143 (N_11143,N_10816,N_10606);
and U11144 (N_11144,N_10550,N_10704);
and U11145 (N_11145,N_10730,N_10820);
or U11146 (N_11146,N_10877,N_10929);
and U11147 (N_11147,N_10764,N_10616);
or U11148 (N_11148,N_10770,N_10710);
or U11149 (N_11149,N_10892,N_10514);
nand U11150 (N_11150,N_10668,N_10895);
nor U11151 (N_11151,N_10589,N_10750);
and U11152 (N_11152,N_10686,N_10886);
nor U11153 (N_11153,N_10969,N_10600);
xnor U11154 (N_11154,N_10928,N_10689);
or U11155 (N_11155,N_10882,N_10765);
nand U11156 (N_11156,N_10907,N_10769);
nor U11157 (N_11157,N_10951,N_10826);
and U11158 (N_11158,N_10866,N_10829);
and U11159 (N_11159,N_10568,N_10649);
nor U11160 (N_11160,N_10991,N_10814);
nor U11161 (N_11161,N_10717,N_10808);
nand U11162 (N_11162,N_10804,N_10549);
nand U11163 (N_11163,N_10909,N_10973);
nand U11164 (N_11164,N_10862,N_10637);
nand U11165 (N_11165,N_10698,N_10683);
nor U11166 (N_11166,N_10687,N_10763);
and U11167 (N_11167,N_10624,N_10800);
or U11168 (N_11168,N_10944,N_10767);
nand U11169 (N_11169,N_10664,N_10898);
nor U11170 (N_11170,N_10729,N_10757);
or U11171 (N_11171,N_10617,N_10724);
nand U11172 (N_11172,N_10574,N_10556);
nor U11173 (N_11173,N_10540,N_10910);
xnor U11174 (N_11174,N_10596,N_10920);
and U11175 (N_11175,N_10635,N_10677);
nand U11176 (N_11176,N_10817,N_10827);
and U11177 (N_11177,N_10756,N_10500);
and U11178 (N_11178,N_10985,N_10602);
nor U11179 (N_11179,N_10838,N_10653);
or U11180 (N_11180,N_10997,N_10843);
nand U11181 (N_11181,N_10947,N_10706);
nor U11182 (N_11182,N_10786,N_10919);
and U11183 (N_11183,N_10806,N_10702);
nor U11184 (N_11184,N_10575,N_10967);
xnor U11185 (N_11185,N_10622,N_10918);
or U11186 (N_11186,N_10865,N_10807);
or U11187 (N_11187,N_10883,N_10905);
nand U11188 (N_11188,N_10956,N_10891);
nand U11189 (N_11189,N_10738,N_10970);
nor U11190 (N_11190,N_10553,N_10621);
xnor U11191 (N_11191,N_10607,N_10660);
nand U11192 (N_11192,N_10697,N_10847);
nand U11193 (N_11193,N_10566,N_10880);
xnor U11194 (N_11194,N_10708,N_10803);
nor U11195 (N_11195,N_10795,N_10609);
and U11196 (N_11196,N_10659,N_10527);
xnor U11197 (N_11197,N_10528,N_10694);
nand U11198 (N_11198,N_10840,N_10773);
and U11199 (N_11199,N_10793,N_10663);
nand U11200 (N_11200,N_10551,N_10523);
nor U11201 (N_11201,N_10885,N_10911);
nor U11202 (N_11202,N_10705,N_10986);
or U11203 (N_11203,N_10719,N_10558);
or U11204 (N_11204,N_10520,N_10990);
or U11205 (N_11205,N_10504,N_10992);
or U11206 (N_11206,N_10916,N_10932);
or U11207 (N_11207,N_10876,N_10679);
nor U11208 (N_11208,N_10681,N_10603);
or U11209 (N_11209,N_10714,N_10999);
nand U11210 (N_11210,N_10921,N_10583);
and U11211 (N_11211,N_10728,N_10810);
and U11212 (N_11212,N_10832,N_10923);
or U11213 (N_11213,N_10789,N_10779);
or U11214 (N_11214,N_10930,N_10996);
and U11215 (N_11215,N_10933,N_10731);
or U11216 (N_11216,N_10822,N_10545);
and U11217 (N_11217,N_10961,N_10801);
nor U11218 (N_11218,N_10665,N_10518);
nor U11219 (N_11219,N_10693,N_10824);
nand U11220 (N_11220,N_10850,N_10675);
nor U11221 (N_11221,N_10611,N_10939);
xnor U11222 (N_11222,N_10573,N_10884);
nor U11223 (N_11223,N_10625,N_10555);
or U11224 (N_11224,N_10501,N_10692);
or U11225 (N_11225,N_10791,N_10943);
or U11226 (N_11226,N_10833,N_10960);
or U11227 (N_11227,N_10925,N_10987);
nand U11228 (N_11228,N_10983,N_10590);
nor U11229 (N_11229,N_10546,N_10646);
nor U11230 (N_11230,N_10988,N_10777);
or U11231 (N_11231,N_10839,N_10541);
and U11232 (N_11232,N_10915,N_10785);
and U11233 (N_11233,N_10538,N_10962);
xnor U11234 (N_11234,N_10721,N_10794);
nor U11235 (N_11235,N_10825,N_10601);
nand U11236 (N_11236,N_10855,N_10634);
or U11237 (N_11237,N_10792,N_10784);
and U11238 (N_11238,N_10771,N_10594);
nand U11239 (N_11239,N_10734,N_10964);
and U11240 (N_11240,N_10727,N_10673);
and U11241 (N_11241,N_10648,N_10759);
or U11242 (N_11242,N_10896,N_10522);
or U11243 (N_11243,N_10554,N_10651);
or U11244 (N_11244,N_10903,N_10906);
or U11245 (N_11245,N_10740,N_10598);
or U11246 (N_11246,N_10751,N_10650);
nand U11247 (N_11247,N_10831,N_10507);
or U11248 (N_11248,N_10949,N_10534);
nand U11249 (N_11249,N_10868,N_10571);
xnor U11250 (N_11250,N_10806,N_10759);
nor U11251 (N_11251,N_10795,N_10622);
nor U11252 (N_11252,N_10991,N_10937);
nand U11253 (N_11253,N_10728,N_10848);
nand U11254 (N_11254,N_10502,N_10841);
or U11255 (N_11255,N_10501,N_10512);
nand U11256 (N_11256,N_10918,N_10536);
or U11257 (N_11257,N_10949,N_10624);
or U11258 (N_11258,N_10513,N_10927);
or U11259 (N_11259,N_10628,N_10997);
and U11260 (N_11260,N_10984,N_10644);
or U11261 (N_11261,N_10815,N_10789);
nor U11262 (N_11262,N_10939,N_10711);
and U11263 (N_11263,N_10513,N_10655);
and U11264 (N_11264,N_10542,N_10967);
and U11265 (N_11265,N_10682,N_10531);
nand U11266 (N_11266,N_10699,N_10729);
or U11267 (N_11267,N_10794,N_10559);
or U11268 (N_11268,N_10544,N_10681);
and U11269 (N_11269,N_10631,N_10903);
and U11270 (N_11270,N_10947,N_10677);
nand U11271 (N_11271,N_10881,N_10685);
or U11272 (N_11272,N_10867,N_10771);
nor U11273 (N_11273,N_10529,N_10741);
or U11274 (N_11274,N_10590,N_10948);
xor U11275 (N_11275,N_10531,N_10530);
and U11276 (N_11276,N_10747,N_10971);
or U11277 (N_11277,N_10555,N_10504);
and U11278 (N_11278,N_10550,N_10651);
nand U11279 (N_11279,N_10790,N_10649);
nand U11280 (N_11280,N_10564,N_10706);
xor U11281 (N_11281,N_10879,N_10999);
nor U11282 (N_11282,N_10622,N_10598);
and U11283 (N_11283,N_10652,N_10861);
nor U11284 (N_11284,N_10910,N_10770);
xor U11285 (N_11285,N_10816,N_10846);
and U11286 (N_11286,N_10684,N_10670);
nand U11287 (N_11287,N_10954,N_10872);
and U11288 (N_11288,N_10580,N_10628);
nor U11289 (N_11289,N_10636,N_10637);
or U11290 (N_11290,N_10674,N_10956);
and U11291 (N_11291,N_10919,N_10582);
nor U11292 (N_11292,N_10760,N_10721);
nor U11293 (N_11293,N_10605,N_10838);
xnor U11294 (N_11294,N_10630,N_10828);
or U11295 (N_11295,N_10925,N_10542);
and U11296 (N_11296,N_10988,N_10883);
nand U11297 (N_11297,N_10526,N_10848);
or U11298 (N_11298,N_10999,N_10997);
nand U11299 (N_11299,N_10913,N_10581);
nor U11300 (N_11300,N_10662,N_10778);
and U11301 (N_11301,N_10786,N_10662);
nand U11302 (N_11302,N_10814,N_10804);
and U11303 (N_11303,N_10700,N_10707);
xor U11304 (N_11304,N_10964,N_10733);
nand U11305 (N_11305,N_10910,N_10624);
xor U11306 (N_11306,N_10563,N_10890);
nor U11307 (N_11307,N_10609,N_10812);
or U11308 (N_11308,N_10843,N_10648);
or U11309 (N_11309,N_10697,N_10843);
and U11310 (N_11310,N_10974,N_10878);
and U11311 (N_11311,N_10786,N_10549);
or U11312 (N_11312,N_10900,N_10776);
and U11313 (N_11313,N_10781,N_10536);
and U11314 (N_11314,N_10991,N_10734);
or U11315 (N_11315,N_10904,N_10942);
nor U11316 (N_11316,N_10727,N_10584);
and U11317 (N_11317,N_10889,N_10970);
or U11318 (N_11318,N_10931,N_10832);
and U11319 (N_11319,N_10938,N_10755);
nand U11320 (N_11320,N_10604,N_10643);
nor U11321 (N_11321,N_10552,N_10713);
nor U11322 (N_11322,N_10626,N_10863);
xnor U11323 (N_11323,N_10755,N_10566);
xnor U11324 (N_11324,N_10841,N_10909);
nor U11325 (N_11325,N_10511,N_10538);
nor U11326 (N_11326,N_10925,N_10629);
nor U11327 (N_11327,N_10523,N_10739);
xor U11328 (N_11328,N_10526,N_10963);
or U11329 (N_11329,N_10948,N_10637);
or U11330 (N_11330,N_10907,N_10518);
and U11331 (N_11331,N_10517,N_10932);
xor U11332 (N_11332,N_10529,N_10607);
and U11333 (N_11333,N_10974,N_10531);
nor U11334 (N_11334,N_10869,N_10794);
and U11335 (N_11335,N_10608,N_10620);
or U11336 (N_11336,N_10876,N_10547);
nor U11337 (N_11337,N_10703,N_10508);
nor U11338 (N_11338,N_10986,N_10505);
xnor U11339 (N_11339,N_10770,N_10896);
nor U11340 (N_11340,N_10506,N_10639);
nand U11341 (N_11341,N_10582,N_10801);
xnor U11342 (N_11342,N_10561,N_10739);
or U11343 (N_11343,N_10862,N_10688);
or U11344 (N_11344,N_10942,N_10885);
or U11345 (N_11345,N_10720,N_10666);
xor U11346 (N_11346,N_10532,N_10903);
or U11347 (N_11347,N_10920,N_10842);
nand U11348 (N_11348,N_10835,N_10705);
nand U11349 (N_11349,N_10966,N_10876);
and U11350 (N_11350,N_10712,N_10571);
or U11351 (N_11351,N_10657,N_10994);
or U11352 (N_11352,N_10880,N_10523);
nand U11353 (N_11353,N_10725,N_10693);
nor U11354 (N_11354,N_10852,N_10893);
or U11355 (N_11355,N_10641,N_10862);
and U11356 (N_11356,N_10849,N_10614);
or U11357 (N_11357,N_10964,N_10823);
xor U11358 (N_11358,N_10617,N_10509);
nor U11359 (N_11359,N_10790,N_10785);
nor U11360 (N_11360,N_10994,N_10722);
and U11361 (N_11361,N_10731,N_10930);
nand U11362 (N_11362,N_10738,N_10836);
nor U11363 (N_11363,N_10811,N_10802);
nor U11364 (N_11364,N_10750,N_10933);
nand U11365 (N_11365,N_10850,N_10605);
nand U11366 (N_11366,N_10735,N_10723);
nand U11367 (N_11367,N_10978,N_10792);
xor U11368 (N_11368,N_10566,N_10959);
nor U11369 (N_11369,N_10650,N_10845);
nor U11370 (N_11370,N_10784,N_10913);
or U11371 (N_11371,N_10860,N_10703);
and U11372 (N_11372,N_10579,N_10554);
nor U11373 (N_11373,N_10623,N_10972);
nor U11374 (N_11374,N_10572,N_10568);
nand U11375 (N_11375,N_10820,N_10694);
nand U11376 (N_11376,N_10636,N_10891);
and U11377 (N_11377,N_10994,N_10781);
and U11378 (N_11378,N_10992,N_10526);
or U11379 (N_11379,N_10579,N_10654);
and U11380 (N_11380,N_10579,N_10817);
nand U11381 (N_11381,N_10760,N_10976);
and U11382 (N_11382,N_10814,N_10962);
nor U11383 (N_11383,N_10697,N_10753);
or U11384 (N_11384,N_10815,N_10668);
or U11385 (N_11385,N_10973,N_10866);
xnor U11386 (N_11386,N_10684,N_10866);
or U11387 (N_11387,N_10745,N_10656);
or U11388 (N_11388,N_10983,N_10595);
nor U11389 (N_11389,N_10591,N_10858);
nor U11390 (N_11390,N_10957,N_10516);
and U11391 (N_11391,N_10805,N_10899);
or U11392 (N_11392,N_10777,N_10604);
xor U11393 (N_11393,N_10601,N_10974);
xor U11394 (N_11394,N_10946,N_10903);
and U11395 (N_11395,N_10864,N_10823);
and U11396 (N_11396,N_10695,N_10926);
nand U11397 (N_11397,N_10658,N_10698);
or U11398 (N_11398,N_10651,N_10615);
nor U11399 (N_11399,N_10943,N_10676);
and U11400 (N_11400,N_10756,N_10682);
or U11401 (N_11401,N_10613,N_10890);
nor U11402 (N_11402,N_10628,N_10708);
or U11403 (N_11403,N_10682,N_10507);
or U11404 (N_11404,N_10841,N_10997);
or U11405 (N_11405,N_10713,N_10859);
nand U11406 (N_11406,N_10524,N_10909);
nor U11407 (N_11407,N_10667,N_10991);
nor U11408 (N_11408,N_10589,N_10761);
nor U11409 (N_11409,N_10608,N_10757);
nand U11410 (N_11410,N_10729,N_10581);
nand U11411 (N_11411,N_10794,N_10944);
or U11412 (N_11412,N_10706,N_10579);
nor U11413 (N_11413,N_10677,N_10911);
nand U11414 (N_11414,N_10699,N_10834);
nor U11415 (N_11415,N_10624,N_10762);
or U11416 (N_11416,N_10725,N_10984);
xnor U11417 (N_11417,N_10917,N_10599);
nor U11418 (N_11418,N_10795,N_10941);
and U11419 (N_11419,N_10951,N_10957);
and U11420 (N_11420,N_10709,N_10507);
nor U11421 (N_11421,N_10681,N_10726);
and U11422 (N_11422,N_10817,N_10764);
and U11423 (N_11423,N_10523,N_10895);
and U11424 (N_11424,N_10871,N_10921);
or U11425 (N_11425,N_10657,N_10870);
and U11426 (N_11426,N_10661,N_10733);
nand U11427 (N_11427,N_10964,N_10562);
and U11428 (N_11428,N_10991,N_10974);
nand U11429 (N_11429,N_10972,N_10930);
nand U11430 (N_11430,N_10748,N_10597);
xnor U11431 (N_11431,N_10735,N_10761);
nand U11432 (N_11432,N_10848,N_10512);
or U11433 (N_11433,N_10816,N_10624);
or U11434 (N_11434,N_10977,N_10897);
nor U11435 (N_11435,N_10875,N_10821);
and U11436 (N_11436,N_10945,N_10837);
nor U11437 (N_11437,N_10790,N_10920);
and U11438 (N_11438,N_10586,N_10516);
nor U11439 (N_11439,N_10574,N_10988);
xor U11440 (N_11440,N_10560,N_10860);
and U11441 (N_11441,N_10694,N_10991);
and U11442 (N_11442,N_10547,N_10822);
and U11443 (N_11443,N_10526,N_10521);
nor U11444 (N_11444,N_10849,N_10618);
nor U11445 (N_11445,N_10579,N_10886);
nand U11446 (N_11446,N_10993,N_10812);
nand U11447 (N_11447,N_10901,N_10541);
xor U11448 (N_11448,N_10871,N_10796);
nor U11449 (N_11449,N_10834,N_10858);
and U11450 (N_11450,N_10518,N_10790);
and U11451 (N_11451,N_10882,N_10860);
and U11452 (N_11452,N_10557,N_10904);
nand U11453 (N_11453,N_10696,N_10690);
nand U11454 (N_11454,N_10711,N_10540);
xor U11455 (N_11455,N_10721,N_10605);
nand U11456 (N_11456,N_10558,N_10737);
and U11457 (N_11457,N_10559,N_10524);
xnor U11458 (N_11458,N_10567,N_10609);
nor U11459 (N_11459,N_10549,N_10547);
nor U11460 (N_11460,N_10945,N_10511);
nand U11461 (N_11461,N_10923,N_10982);
nand U11462 (N_11462,N_10521,N_10954);
nor U11463 (N_11463,N_10993,N_10541);
or U11464 (N_11464,N_10942,N_10576);
and U11465 (N_11465,N_10982,N_10874);
nor U11466 (N_11466,N_10574,N_10892);
nand U11467 (N_11467,N_10732,N_10836);
or U11468 (N_11468,N_10660,N_10944);
and U11469 (N_11469,N_10690,N_10945);
or U11470 (N_11470,N_10704,N_10647);
or U11471 (N_11471,N_10592,N_10550);
nor U11472 (N_11472,N_10562,N_10810);
and U11473 (N_11473,N_10899,N_10562);
nand U11474 (N_11474,N_10800,N_10982);
or U11475 (N_11475,N_10993,N_10991);
nor U11476 (N_11476,N_10853,N_10511);
nor U11477 (N_11477,N_10714,N_10900);
or U11478 (N_11478,N_10896,N_10981);
nor U11479 (N_11479,N_10967,N_10643);
nor U11480 (N_11480,N_10643,N_10764);
nand U11481 (N_11481,N_10528,N_10705);
xor U11482 (N_11482,N_10966,N_10924);
or U11483 (N_11483,N_10963,N_10598);
or U11484 (N_11484,N_10610,N_10950);
or U11485 (N_11485,N_10841,N_10703);
or U11486 (N_11486,N_10809,N_10673);
or U11487 (N_11487,N_10810,N_10645);
and U11488 (N_11488,N_10666,N_10930);
nand U11489 (N_11489,N_10986,N_10920);
nor U11490 (N_11490,N_10810,N_10797);
or U11491 (N_11491,N_10897,N_10868);
and U11492 (N_11492,N_10553,N_10913);
xor U11493 (N_11493,N_10885,N_10838);
or U11494 (N_11494,N_10833,N_10818);
or U11495 (N_11495,N_10681,N_10662);
nor U11496 (N_11496,N_10850,N_10579);
or U11497 (N_11497,N_10699,N_10842);
nor U11498 (N_11498,N_10602,N_10930);
nor U11499 (N_11499,N_10519,N_10939);
and U11500 (N_11500,N_11073,N_11204);
or U11501 (N_11501,N_11130,N_11279);
nor U11502 (N_11502,N_11151,N_11415);
or U11503 (N_11503,N_11060,N_11387);
nor U11504 (N_11504,N_11406,N_11470);
and U11505 (N_11505,N_11260,N_11100);
nor U11506 (N_11506,N_11002,N_11286);
and U11507 (N_11507,N_11041,N_11444);
nand U11508 (N_11508,N_11135,N_11342);
and U11509 (N_11509,N_11178,N_11490);
nor U11510 (N_11510,N_11032,N_11142);
and U11511 (N_11511,N_11423,N_11085);
nand U11512 (N_11512,N_11416,N_11497);
nor U11513 (N_11513,N_11327,N_11217);
nor U11514 (N_11514,N_11303,N_11379);
or U11515 (N_11515,N_11484,N_11399);
and U11516 (N_11516,N_11143,N_11083);
or U11517 (N_11517,N_11499,N_11413);
nand U11518 (N_11518,N_11386,N_11312);
nor U11519 (N_11519,N_11113,N_11330);
or U11520 (N_11520,N_11350,N_11006);
and U11521 (N_11521,N_11426,N_11173);
nand U11522 (N_11522,N_11261,N_11369);
nand U11523 (N_11523,N_11468,N_11079);
nor U11524 (N_11524,N_11268,N_11007);
nor U11525 (N_11525,N_11114,N_11000);
nand U11526 (N_11526,N_11176,N_11337);
or U11527 (N_11527,N_11109,N_11466);
xor U11528 (N_11528,N_11152,N_11035);
nand U11529 (N_11529,N_11202,N_11192);
and U11530 (N_11530,N_11324,N_11424);
nand U11531 (N_11531,N_11485,N_11036);
nand U11532 (N_11532,N_11427,N_11056);
xnor U11533 (N_11533,N_11298,N_11281);
and U11534 (N_11534,N_11419,N_11317);
and U11535 (N_11535,N_11044,N_11263);
and U11536 (N_11536,N_11482,N_11012);
or U11537 (N_11537,N_11187,N_11095);
nor U11538 (N_11538,N_11272,N_11154);
and U11539 (N_11539,N_11471,N_11045);
or U11540 (N_11540,N_11163,N_11241);
or U11541 (N_11541,N_11216,N_11318);
nand U11542 (N_11542,N_11161,N_11137);
nand U11543 (N_11543,N_11206,N_11120);
and U11544 (N_11544,N_11400,N_11050);
and U11545 (N_11545,N_11365,N_11053);
or U11546 (N_11546,N_11134,N_11267);
nor U11547 (N_11547,N_11090,N_11183);
nand U11548 (N_11548,N_11244,N_11086);
nand U11549 (N_11549,N_11059,N_11066);
xor U11550 (N_11550,N_11165,N_11132);
or U11551 (N_11551,N_11401,N_11469);
nand U11552 (N_11552,N_11283,N_11333);
nand U11553 (N_11553,N_11474,N_11462);
nor U11554 (N_11554,N_11402,N_11326);
or U11555 (N_11555,N_11243,N_11184);
or U11556 (N_11556,N_11316,N_11384);
and U11557 (N_11557,N_11352,N_11069);
nor U11558 (N_11558,N_11033,N_11396);
and U11559 (N_11559,N_11203,N_11123);
or U11560 (N_11560,N_11037,N_11052);
and U11561 (N_11561,N_11221,N_11082);
or U11562 (N_11562,N_11408,N_11456);
or U11563 (N_11563,N_11453,N_11103);
or U11564 (N_11564,N_11201,N_11043);
or U11565 (N_11565,N_11273,N_11488);
nand U11566 (N_11566,N_11102,N_11025);
or U11567 (N_11567,N_11495,N_11382);
nor U11568 (N_11568,N_11160,N_11170);
xor U11569 (N_11569,N_11055,N_11277);
xnor U11570 (N_11570,N_11105,N_11167);
nor U11571 (N_11571,N_11451,N_11362);
nand U11572 (N_11572,N_11096,N_11332);
or U11573 (N_11573,N_11126,N_11275);
nand U11574 (N_11574,N_11015,N_11046);
and U11575 (N_11575,N_11486,N_11145);
nor U11576 (N_11576,N_11383,N_11129);
nand U11577 (N_11577,N_11254,N_11067);
nor U11578 (N_11578,N_11323,N_11226);
or U11579 (N_11579,N_11459,N_11230);
and U11580 (N_11580,N_11247,N_11348);
nor U11581 (N_11581,N_11224,N_11371);
or U11582 (N_11582,N_11321,N_11172);
or U11583 (N_11583,N_11262,N_11181);
and U11584 (N_11584,N_11021,N_11309);
or U11585 (N_11585,N_11122,N_11472);
nor U11586 (N_11586,N_11245,N_11403);
and U11587 (N_11587,N_11479,N_11271);
nor U11588 (N_11588,N_11011,N_11393);
or U11589 (N_11589,N_11162,N_11465);
or U11590 (N_11590,N_11363,N_11394);
xor U11591 (N_11591,N_11098,N_11099);
and U11592 (N_11592,N_11443,N_11106);
and U11593 (N_11593,N_11322,N_11213);
xor U11594 (N_11594,N_11346,N_11038);
or U11595 (N_11595,N_11421,N_11288);
nand U11596 (N_11596,N_11364,N_11158);
nor U11597 (N_11597,N_11237,N_11207);
or U11598 (N_11598,N_11040,N_11328);
nor U11599 (N_11599,N_11445,N_11392);
and U11600 (N_11600,N_11141,N_11039);
nand U11601 (N_11601,N_11084,N_11340);
or U11602 (N_11602,N_11496,N_11133);
nor U11603 (N_11603,N_11320,N_11344);
xnor U11604 (N_11604,N_11140,N_11013);
nor U11605 (N_11605,N_11477,N_11448);
nor U11606 (N_11606,N_11343,N_11212);
nor U11607 (N_11607,N_11433,N_11336);
nor U11608 (N_11608,N_11087,N_11194);
or U11609 (N_11609,N_11285,N_11068);
nand U11610 (N_11610,N_11308,N_11003);
or U11611 (N_11611,N_11205,N_11291);
or U11612 (N_11612,N_11048,N_11414);
nand U11613 (N_11613,N_11374,N_11397);
nand U11614 (N_11614,N_11420,N_11155);
nand U11615 (N_11615,N_11240,N_11351);
and U11616 (N_11616,N_11004,N_11492);
or U11617 (N_11617,N_11338,N_11347);
nand U11618 (N_11618,N_11229,N_11115);
or U11619 (N_11619,N_11460,N_11110);
or U11620 (N_11620,N_11009,N_11218);
nand U11621 (N_11621,N_11325,N_11047);
nor U11622 (N_11622,N_11255,N_11127);
nand U11623 (N_11623,N_11175,N_11425);
or U11624 (N_11624,N_11080,N_11353);
xnor U11625 (N_11625,N_11149,N_11131);
nor U11626 (N_11626,N_11051,N_11228);
or U11627 (N_11627,N_11071,N_11264);
and U11628 (N_11628,N_11016,N_11307);
xor U11629 (N_11629,N_11225,N_11014);
nand U11630 (N_11630,N_11375,N_11169);
nor U11631 (N_11631,N_11258,N_11447);
nor U11632 (N_11632,N_11431,N_11370);
nand U11633 (N_11633,N_11189,N_11372);
nor U11634 (N_11634,N_11180,N_11027);
xnor U11635 (N_11635,N_11250,N_11159);
nor U11636 (N_11636,N_11359,N_11199);
nand U11637 (N_11637,N_11315,N_11239);
nand U11638 (N_11638,N_11092,N_11491);
nand U11639 (N_11639,N_11434,N_11265);
and U11640 (N_11640,N_11390,N_11211);
and U11641 (N_11641,N_11437,N_11028);
or U11642 (N_11642,N_11058,N_11227);
nor U11643 (N_11643,N_11481,N_11295);
and U11644 (N_11644,N_11380,N_11215);
nor U11645 (N_11645,N_11449,N_11417);
and U11646 (N_11646,N_11138,N_11329);
nor U11647 (N_11647,N_11305,N_11168);
xor U11648 (N_11648,N_11024,N_11054);
nand U11649 (N_11649,N_11442,N_11026);
nor U11650 (N_11650,N_11253,N_11185);
nor U11651 (N_11651,N_11210,N_11008);
nand U11652 (N_11652,N_11197,N_11407);
and U11653 (N_11653,N_11269,N_11287);
xor U11654 (N_11654,N_11101,N_11065);
or U11655 (N_11655,N_11139,N_11428);
or U11656 (N_11656,N_11270,N_11182);
nand U11657 (N_11657,N_11422,N_11301);
nand U11658 (N_11658,N_11191,N_11061);
nand U11659 (N_11659,N_11251,N_11429);
nor U11660 (N_11660,N_11411,N_11404);
or U11661 (N_11661,N_11200,N_11467);
nand U11662 (N_11662,N_11432,N_11136);
nand U11663 (N_11663,N_11001,N_11223);
nor U11664 (N_11664,N_11311,N_11248);
or U11665 (N_11665,N_11121,N_11302);
and U11666 (N_11666,N_11062,N_11334);
nand U11667 (N_11667,N_11005,N_11112);
and U11668 (N_11668,N_11089,N_11299);
and U11669 (N_11669,N_11023,N_11331);
and U11670 (N_11670,N_11107,N_11118);
nand U11671 (N_11671,N_11124,N_11238);
nor U11672 (N_11672,N_11461,N_11487);
or U11673 (N_11673,N_11385,N_11042);
and U11674 (N_11674,N_11438,N_11310);
or U11675 (N_11675,N_11094,N_11018);
and U11676 (N_11676,N_11355,N_11398);
nand U11677 (N_11677,N_11171,N_11483);
and U11678 (N_11678,N_11235,N_11148);
nand U11679 (N_11679,N_11029,N_11358);
or U11680 (N_11680,N_11019,N_11360);
and U11681 (N_11681,N_11156,N_11439);
xnor U11682 (N_11682,N_11446,N_11441);
or U11683 (N_11683,N_11440,N_11246);
and U11684 (N_11684,N_11430,N_11473);
nor U11685 (N_11685,N_11147,N_11111);
or U11686 (N_11686,N_11164,N_11219);
nand U11687 (N_11687,N_11280,N_11234);
or U11688 (N_11688,N_11146,N_11208);
and U11689 (N_11689,N_11153,N_11074);
and U11690 (N_11690,N_11116,N_11341);
nor U11691 (N_11691,N_11489,N_11284);
nand U11692 (N_11692,N_11128,N_11242);
or U11693 (N_11693,N_11193,N_11405);
xor U11694 (N_11694,N_11150,N_11314);
and U11695 (N_11695,N_11233,N_11196);
nor U11696 (N_11696,N_11457,N_11498);
xnor U11697 (N_11697,N_11367,N_11020);
nor U11698 (N_11698,N_11373,N_11378);
and U11699 (N_11699,N_11034,N_11209);
or U11700 (N_11700,N_11377,N_11278);
xor U11701 (N_11701,N_11292,N_11010);
xnor U11702 (N_11702,N_11186,N_11361);
or U11703 (N_11703,N_11252,N_11409);
xnor U11704 (N_11704,N_11354,N_11188);
nor U11705 (N_11705,N_11368,N_11177);
nand U11706 (N_11706,N_11418,N_11088);
or U11707 (N_11707,N_11339,N_11174);
nand U11708 (N_11708,N_11195,N_11294);
and U11709 (N_11709,N_11455,N_11017);
nor U11710 (N_11710,N_11075,N_11293);
nand U11711 (N_11711,N_11464,N_11249);
nor U11712 (N_11712,N_11290,N_11117);
or U11713 (N_11713,N_11125,N_11266);
or U11714 (N_11714,N_11450,N_11144);
or U11715 (N_11715,N_11391,N_11157);
and U11716 (N_11716,N_11274,N_11436);
xnor U11717 (N_11717,N_11222,N_11214);
nand U11718 (N_11718,N_11296,N_11081);
xnor U11719 (N_11719,N_11077,N_11259);
nand U11720 (N_11720,N_11345,N_11412);
nand U11721 (N_11721,N_11349,N_11306);
nor U11722 (N_11722,N_11104,N_11097);
and U11723 (N_11723,N_11031,N_11166);
nand U11724 (N_11724,N_11480,N_11198);
nor U11725 (N_11725,N_11257,N_11313);
nor U11726 (N_11726,N_11022,N_11057);
nand U11727 (N_11727,N_11366,N_11476);
nand U11728 (N_11728,N_11282,N_11376);
nand U11729 (N_11729,N_11276,N_11458);
nor U11730 (N_11730,N_11049,N_11220);
and U11731 (N_11731,N_11395,N_11091);
or U11732 (N_11732,N_11389,N_11070);
or U11733 (N_11733,N_11356,N_11289);
xnor U11734 (N_11734,N_11319,N_11494);
or U11735 (N_11735,N_11236,N_11463);
and U11736 (N_11736,N_11179,N_11452);
nand U11737 (N_11737,N_11190,N_11357);
nor U11738 (N_11738,N_11381,N_11256);
nand U11739 (N_11739,N_11078,N_11435);
or U11740 (N_11740,N_11063,N_11232);
and U11741 (N_11741,N_11064,N_11072);
nand U11742 (N_11742,N_11493,N_11231);
nand U11743 (N_11743,N_11304,N_11300);
or U11744 (N_11744,N_11119,N_11410);
nor U11745 (N_11745,N_11454,N_11030);
nor U11746 (N_11746,N_11297,N_11388);
nor U11747 (N_11747,N_11475,N_11478);
or U11748 (N_11748,N_11335,N_11093);
nand U11749 (N_11749,N_11108,N_11076);
nor U11750 (N_11750,N_11012,N_11229);
and U11751 (N_11751,N_11420,N_11357);
nand U11752 (N_11752,N_11444,N_11141);
nand U11753 (N_11753,N_11084,N_11317);
or U11754 (N_11754,N_11321,N_11100);
nor U11755 (N_11755,N_11232,N_11122);
nand U11756 (N_11756,N_11340,N_11381);
nor U11757 (N_11757,N_11022,N_11365);
or U11758 (N_11758,N_11083,N_11467);
or U11759 (N_11759,N_11234,N_11200);
and U11760 (N_11760,N_11048,N_11049);
and U11761 (N_11761,N_11308,N_11257);
and U11762 (N_11762,N_11086,N_11386);
xor U11763 (N_11763,N_11487,N_11462);
nor U11764 (N_11764,N_11384,N_11268);
or U11765 (N_11765,N_11013,N_11162);
or U11766 (N_11766,N_11090,N_11225);
and U11767 (N_11767,N_11429,N_11214);
nor U11768 (N_11768,N_11378,N_11387);
xnor U11769 (N_11769,N_11174,N_11218);
nor U11770 (N_11770,N_11063,N_11130);
and U11771 (N_11771,N_11318,N_11392);
or U11772 (N_11772,N_11321,N_11496);
or U11773 (N_11773,N_11390,N_11256);
xnor U11774 (N_11774,N_11388,N_11213);
nand U11775 (N_11775,N_11412,N_11016);
nor U11776 (N_11776,N_11363,N_11029);
and U11777 (N_11777,N_11478,N_11101);
xnor U11778 (N_11778,N_11415,N_11135);
nand U11779 (N_11779,N_11151,N_11117);
or U11780 (N_11780,N_11109,N_11276);
nor U11781 (N_11781,N_11113,N_11031);
and U11782 (N_11782,N_11146,N_11021);
nand U11783 (N_11783,N_11299,N_11291);
or U11784 (N_11784,N_11099,N_11370);
nor U11785 (N_11785,N_11279,N_11241);
or U11786 (N_11786,N_11089,N_11163);
and U11787 (N_11787,N_11190,N_11235);
nor U11788 (N_11788,N_11168,N_11110);
xnor U11789 (N_11789,N_11449,N_11024);
or U11790 (N_11790,N_11199,N_11022);
and U11791 (N_11791,N_11389,N_11404);
nor U11792 (N_11792,N_11209,N_11286);
nand U11793 (N_11793,N_11066,N_11247);
or U11794 (N_11794,N_11002,N_11083);
or U11795 (N_11795,N_11031,N_11444);
nand U11796 (N_11796,N_11256,N_11025);
or U11797 (N_11797,N_11257,N_11051);
nor U11798 (N_11798,N_11236,N_11271);
nand U11799 (N_11799,N_11078,N_11141);
nand U11800 (N_11800,N_11459,N_11419);
or U11801 (N_11801,N_11139,N_11105);
nand U11802 (N_11802,N_11285,N_11209);
and U11803 (N_11803,N_11204,N_11047);
and U11804 (N_11804,N_11079,N_11338);
nor U11805 (N_11805,N_11326,N_11075);
and U11806 (N_11806,N_11187,N_11448);
or U11807 (N_11807,N_11032,N_11496);
nand U11808 (N_11808,N_11092,N_11240);
nor U11809 (N_11809,N_11347,N_11147);
nand U11810 (N_11810,N_11307,N_11481);
or U11811 (N_11811,N_11318,N_11466);
nand U11812 (N_11812,N_11227,N_11298);
xor U11813 (N_11813,N_11365,N_11203);
xnor U11814 (N_11814,N_11261,N_11196);
or U11815 (N_11815,N_11496,N_11341);
and U11816 (N_11816,N_11211,N_11253);
nand U11817 (N_11817,N_11311,N_11279);
nor U11818 (N_11818,N_11268,N_11350);
nor U11819 (N_11819,N_11081,N_11248);
nor U11820 (N_11820,N_11412,N_11262);
nor U11821 (N_11821,N_11087,N_11128);
or U11822 (N_11822,N_11089,N_11439);
or U11823 (N_11823,N_11464,N_11005);
and U11824 (N_11824,N_11154,N_11394);
and U11825 (N_11825,N_11066,N_11268);
xnor U11826 (N_11826,N_11426,N_11042);
nand U11827 (N_11827,N_11299,N_11158);
or U11828 (N_11828,N_11484,N_11134);
nor U11829 (N_11829,N_11358,N_11231);
nand U11830 (N_11830,N_11193,N_11093);
nor U11831 (N_11831,N_11109,N_11402);
or U11832 (N_11832,N_11482,N_11274);
and U11833 (N_11833,N_11481,N_11225);
xor U11834 (N_11834,N_11081,N_11164);
xnor U11835 (N_11835,N_11173,N_11227);
nand U11836 (N_11836,N_11097,N_11010);
or U11837 (N_11837,N_11128,N_11217);
nand U11838 (N_11838,N_11428,N_11393);
nor U11839 (N_11839,N_11491,N_11303);
or U11840 (N_11840,N_11119,N_11138);
or U11841 (N_11841,N_11422,N_11421);
xnor U11842 (N_11842,N_11180,N_11077);
nor U11843 (N_11843,N_11378,N_11161);
nand U11844 (N_11844,N_11376,N_11386);
and U11845 (N_11845,N_11334,N_11132);
or U11846 (N_11846,N_11162,N_11274);
and U11847 (N_11847,N_11175,N_11029);
nor U11848 (N_11848,N_11031,N_11185);
and U11849 (N_11849,N_11290,N_11429);
nand U11850 (N_11850,N_11298,N_11495);
and U11851 (N_11851,N_11319,N_11428);
and U11852 (N_11852,N_11091,N_11161);
or U11853 (N_11853,N_11314,N_11198);
nand U11854 (N_11854,N_11251,N_11415);
xnor U11855 (N_11855,N_11298,N_11190);
xnor U11856 (N_11856,N_11307,N_11154);
or U11857 (N_11857,N_11280,N_11476);
and U11858 (N_11858,N_11417,N_11116);
nand U11859 (N_11859,N_11366,N_11013);
or U11860 (N_11860,N_11347,N_11069);
nand U11861 (N_11861,N_11028,N_11449);
nor U11862 (N_11862,N_11192,N_11280);
xor U11863 (N_11863,N_11336,N_11219);
or U11864 (N_11864,N_11163,N_11284);
nor U11865 (N_11865,N_11475,N_11189);
nand U11866 (N_11866,N_11079,N_11137);
nand U11867 (N_11867,N_11093,N_11492);
nor U11868 (N_11868,N_11397,N_11408);
and U11869 (N_11869,N_11456,N_11315);
nor U11870 (N_11870,N_11328,N_11326);
xor U11871 (N_11871,N_11420,N_11116);
nand U11872 (N_11872,N_11476,N_11211);
nor U11873 (N_11873,N_11158,N_11350);
and U11874 (N_11874,N_11479,N_11135);
nand U11875 (N_11875,N_11417,N_11427);
nand U11876 (N_11876,N_11028,N_11308);
nand U11877 (N_11877,N_11117,N_11030);
or U11878 (N_11878,N_11143,N_11492);
nor U11879 (N_11879,N_11391,N_11308);
nand U11880 (N_11880,N_11165,N_11336);
or U11881 (N_11881,N_11014,N_11293);
nand U11882 (N_11882,N_11044,N_11046);
xnor U11883 (N_11883,N_11019,N_11300);
nand U11884 (N_11884,N_11223,N_11193);
or U11885 (N_11885,N_11437,N_11159);
nor U11886 (N_11886,N_11484,N_11111);
nor U11887 (N_11887,N_11461,N_11366);
nand U11888 (N_11888,N_11470,N_11365);
nor U11889 (N_11889,N_11477,N_11084);
nand U11890 (N_11890,N_11416,N_11187);
nor U11891 (N_11891,N_11057,N_11018);
xnor U11892 (N_11892,N_11438,N_11152);
and U11893 (N_11893,N_11369,N_11219);
xor U11894 (N_11894,N_11210,N_11411);
and U11895 (N_11895,N_11002,N_11415);
nor U11896 (N_11896,N_11012,N_11288);
nor U11897 (N_11897,N_11181,N_11075);
or U11898 (N_11898,N_11001,N_11351);
nand U11899 (N_11899,N_11040,N_11195);
nand U11900 (N_11900,N_11239,N_11025);
and U11901 (N_11901,N_11327,N_11079);
nor U11902 (N_11902,N_11338,N_11095);
or U11903 (N_11903,N_11457,N_11406);
nor U11904 (N_11904,N_11220,N_11018);
and U11905 (N_11905,N_11455,N_11442);
or U11906 (N_11906,N_11497,N_11428);
nand U11907 (N_11907,N_11422,N_11442);
nor U11908 (N_11908,N_11419,N_11068);
or U11909 (N_11909,N_11454,N_11291);
xnor U11910 (N_11910,N_11386,N_11036);
and U11911 (N_11911,N_11290,N_11326);
nor U11912 (N_11912,N_11159,N_11266);
nor U11913 (N_11913,N_11433,N_11021);
nand U11914 (N_11914,N_11365,N_11405);
or U11915 (N_11915,N_11336,N_11347);
nor U11916 (N_11916,N_11002,N_11025);
nor U11917 (N_11917,N_11258,N_11286);
and U11918 (N_11918,N_11000,N_11137);
and U11919 (N_11919,N_11037,N_11350);
and U11920 (N_11920,N_11233,N_11161);
nand U11921 (N_11921,N_11325,N_11153);
nand U11922 (N_11922,N_11411,N_11154);
or U11923 (N_11923,N_11399,N_11259);
nand U11924 (N_11924,N_11418,N_11360);
nand U11925 (N_11925,N_11042,N_11218);
and U11926 (N_11926,N_11125,N_11304);
and U11927 (N_11927,N_11422,N_11293);
nor U11928 (N_11928,N_11404,N_11336);
nand U11929 (N_11929,N_11096,N_11253);
nor U11930 (N_11930,N_11067,N_11133);
nor U11931 (N_11931,N_11142,N_11113);
nand U11932 (N_11932,N_11428,N_11338);
or U11933 (N_11933,N_11169,N_11105);
nor U11934 (N_11934,N_11132,N_11375);
nor U11935 (N_11935,N_11195,N_11496);
or U11936 (N_11936,N_11367,N_11223);
xor U11937 (N_11937,N_11498,N_11219);
nand U11938 (N_11938,N_11076,N_11443);
nor U11939 (N_11939,N_11290,N_11254);
nand U11940 (N_11940,N_11490,N_11276);
and U11941 (N_11941,N_11324,N_11216);
nand U11942 (N_11942,N_11273,N_11470);
xor U11943 (N_11943,N_11367,N_11229);
or U11944 (N_11944,N_11211,N_11258);
and U11945 (N_11945,N_11035,N_11301);
nor U11946 (N_11946,N_11440,N_11191);
nor U11947 (N_11947,N_11453,N_11266);
nor U11948 (N_11948,N_11493,N_11238);
nand U11949 (N_11949,N_11220,N_11217);
nand U11950 (N_11950,N_11233,N_11136);
and U11951 (N_11951,N_11382,N_11294);
nand U11952 (N_11952,N_11391,N_11183);
nor U11953 (N_11953,N_11348,N_11469);
nor U11954 (N_11954,N_11391,N_11218);
nor U11955 (N_11955,N_11010,N_11368);
xor U11956 (N_11956,N_11043,N_11417);
nand U11957 (N_11957,N_11196,N_11405);
or U11958 (N_11958,N_11072,N_11495);
or U11959 (N_11959,N_11178,N_11168);
and U11960 (N_11960,N_11457,N_11061);
and U11961 (N_11961,N_11320,N_11168);
nand U11962 (N_11962,N_11152,N_11477);
or U11963 (N_11963,N_11148,N_11122);
or U11964 (N_11964,N_11490,N_11488);
and U11965 (N_11965,N_11216,N_11238);
or U11966 (N_11966,N_11263,N_11053);
and U11967 (N_11967,N_11114,N_11165);
nand U11968 (N_11968,N_11356,N_11032);
nor U11969 (N_11969,N_11446,N_11193);
nor U11970 (N_11970,N_11479,N_11040);
nor U11971 (N_11971,N_11151,N_11045);
nand U11972 (N_11972,N_11052,N_11156);
nor U11973 (N_11973,N_11097,N_11195);
xnor U11974 (N_11974,N_11334,N_11201);
and U11975 (N_11975,N_11080,N_11190);
and U11976 (N_11976,N_11035,N_11025);
and U11977 (N_11977,N_11152,N_11380);
and U11978 (N_11978,N_11474,N_11189);
nand U11979 (N_11979,N_11363,N_11322);
or U11980 (N_11980,N_11271,N_11215);
nand U11981 (N_11981,N_11347,N_11480);
nor U11982 (N_11982,N_11159,N_11218);
nand U11983 (N_11983,N_11201,N_11270);
nand U11984 (N_11984,N_11331,N_11247);
and U11985 (N_11985,N_11463,N_11439);
or U11986 (N_11986,N_11499,N_11336);
nor U11987 (N_11987,N_11290,N_11460);
or U11988 (N_11988,N_11460,N_11198);
nor U11989 (N_11989,N_11288,N_11320);
nor U11990 (N_11990,N_11278,N_11279);
xor U11991 (N_11991,N_11493,N_11427);
nor U11992 (N_11992,N_11196,N_11171);
and U11993 (N_11993,N_11321,N_11133);
and U11994 (N_11994,N_11312,N_11127);
xor U11995 (N_11995,N_11016,N_11344);
and U11996 (N_11996,N_11080,N_11419);
and U11997 (N_11997,N_11063,N_11449);
or U11998 (N_11998,N_11374,N_11198);
or U11999 (N_11999,N_11286,N_11470);
or U12000 (N_12000,N_11935,N_11503);
nand U12001 (N_12001,N_11609,N_11994);
or U12002 (N_12002,N_11598,N_11651);
or U12003 (N_12003,N_11646,N_11642);
nand U12004 (N_12004,N_11560,N_11562);
nor U12005 (N_12005,N_11838,N_11600);
or U12006 (N_12006,N_11734,N_11908);
or U12007 (N_12007,N_11858,N_11707);
or U12008 (N_12008,N_11510,N_11763);
nor U12009 (N_12009,N_11686,N_11962);
nor U12010 (N_12010,N_11530,N_11957);
nand U12011 (N_12011,N_11783,N_11666);
xnor U12012 (N_12012,N_11737,N_11977);
nor U12013 (N_12013,N_11967,N_11717);
and U12014 (N_12014,N_11702,N_11703);
or U12015 (N_12015,N_11964,N_11552);
xor U12016 (N_12016,N_11509,N_11638);
nor U12017 (N_12017,N_11840,N_11541);
or U12018 (N_12018,N_11904,N_11695);
or U12019 (N_12019,N_11911,N_11831);
xnor U12020 (N_12020,N_11869,N_11889);
or U12021 (N_12021,N_11993,N_11513);
nand U12022 (N_12022,N_11821,N_11872);
nor U12023 (N_12023,N_11571,N_11898);
and U12024 (N_12024,N_11902,N_11755);
and U12025 (N_12025,N_11829,N_11584);
nor U12026 (N_12026,N_11713,N_11945);
or U12027 (N_12027,N_11801,N_11969);
or U12028 (N_12028,N_11820,N_11874);
nand U12029 (N_12029,N_11796,N_11777);
nor U12030 (N_12030,N_11819,N_11850);
and U12031 (N_12031,N_11657,N_11950);
xnor U12032 (N_12032,N_11611,N_11716);
xor U12033 (N_12033,N_11960,N_11572);
nand U12034 (N_12034,N_11832,N_11568);
nor U12035 (N_12035,N_11698,N_11573);
and U12036 (N_12036,N_11963,N_11797);
nor U12037 (N_12037,N_11735,N_11596);
and U12038 (N_12038,N_11738,N_11842);
xor U12039 (N_12039,N_11813,N_11655);
xnor U12040 (N_12040,N_11759,N_11949);
or U12041 (N_12041,N_11937,N_11885);
nand U12042 (N_12042,N_11604,N_11909);
nand U12043 (N_12043,N_11675,N_11507);
and U12044 (N_12044,N_11661,N_11711);
nor U12045 (N_12045,N_11585,N_11623);
nand U12046 (N_12046,N_11794,N_11606);
or U12047 (N_12047,N_11679,N_11762);
or U12048 (N_12048,N_11527,N_11750);
or U12049 (N_12049,N_11894,N_11860);
nor U12050 (N_12050,N_11896,N_11792);
and U12051 (N_12051,N_11757,N_11618);
and U12052 (N_12052,N_11617,N_11980);
or U12053 (N_12053,N_11859,N_11555);
or U12054 (N_12054,N_11929,N_11942);
nand U12055 (N_12055,N_11563,N_11628);
nand U12056 (N_12056,N_11536,N_11765);
nand U12057 (N_12057,N_11613,N_11981);
nor U12058 (N_12058,N_11932,N_11923);
nor U12059 (N_12059,N_11883,N_11636);
or U12060 (N_12060,N_11951,N_11982);
or U12061 (N_12061,N_11729,N_11799);
nand U12062 (N_12062,N_11812,N_11641);
and U12063 (N_12063,N_11927,N_11903);
and U12064 (N_12064,N_11660,N_11905);
or U12065 (N_12065,N_11870,N_11518);
nand U12066 (N_12066,N_11986,N_11540);
nor U12067 (N_12067,N_11658,N_11591);
and U12068 (N_12068,N_11997,N_11669);
nor U12069 (N_12069,N_11991,N_11543);
nor U12070 (N_12070,N_11815,N_11914);
or U12071 (N_12071,N_11793,N_11938);
or U12072 (N_12072,N_11549,N_11590);
nand U12073 (N_12073,N_11579,N_11728);
or U12074 (N_12074,N_11688,N_11545);
or U12075 (N_12075,N_11514,N_11682);
nand U12076 (N_12076,N_11913,N_11817);
nand U12077 (N_12077,N_11694,N_11972);
or U12078 (N_12078,N_11643,N_11798);
or U12079 (N_12079,N_11516,N_11745);
and U12080 (N_12080,N_11925,N_11630);
or U12081 (N_12081,N_11577,N_11683);
and U12082 (N_12082,N_11710,N_11715);
nor U12083 (N_12083,N_11625,N_11551);
nand U12084 (N_12084,N_11559,N_11578);
nand U12085 (N_12085,N_11833,N_11934);
and U12086 (N_12086,N_11827,N_11684);
nand U12087 (N_12087,N_11824,N_11924);
or U12088 (N_12088,N_11589,N_11721);
or U12089 (N_12089,N_11996,N_11887);
nand U12090 (N_12090,N_11848,N_11640);
and U12091 (N_12091,N_11802,N_11533);
or U12092 (N_12092,N_11546,N_11880);
nand U12093 (N_12093,N_11774,N_11693);
or U12094 (N_12094,N_11515,N_11569);
and U12095 (N_12095,N_11749,N_11839);
and U12096 (N_12096,N_11622,N_11878);
and U12097 (N_12097,N_11779,N_11770);
or U12098 (N_12098,N_11843,N_11955);
nand U12099 (N_12099,N_11989,N_11891);
or U12100 (N_12100,N_11588,N_11631);
xnor U12101 (N_12101,N_11998,N_11520);
or U12102 (N_12102,N_11856,N_11775);
nor U12103 (N_12103,N_11714,N_11603);
and U12104 (N_12104,N_11766,N_11768);
and U12105 (N_12105,N_11731,N_11940);
nor U12106 (N_12106,N_11992,N_11760);
xnor U12107 (N_12107,N_11849,N_11884);
nor U12108 (N_12108,N_11875,N_11825);
and U12109 (N_12109,N_11971,N_11550);
nand U12110 (N_12110,N_11814,N_11806);
nor U12111 (N_12111,N_11736,N_11795);
nor U12112 (N_12112,N_11685,N_11637);
or U12113 (N_12113,N_11649,N_11639);
and U12114 (N_12114,N_11751,N_11601);
and U12115 (N_12115,N_11882,N_11895);
nor U12116 (N_12116,N_11505,N_11519);
and U12117 (N_12117,N_11754,N_11784);
or U12118 (N_12118,N_11629,N_11855);
nor U12119 (N_12119,N_11633,N_11867);
or U12120 (N_12120,N_11916,N_11995);
or U12121 (N_12121,N_11746,N_11785);
nand U12122 (N_12122,N_11910,N_11594);
or U12123 (N_12123,N_11844,N_11761);
nor U12124 (N_12124,N_11906,N_11668);
nand U12125 (N_12125,N_11758,N_11567);
and U12126 (N_12126,N_11733,N_11958);
and U12127 (N_12127,N_11580,N_11803);
or U12128 (N_12128,N_11805,N_11724);
nor U12129 (N_12129,N_11608,N_11534);
nand U12130 (N_12130,N_11947,N_11930);
nor U12131 (N_12131,N_11922,N_11644);
and U12132 (N_12132,N_11808,N_11901);
nor U12133 (N_12133,N_11939,N_11502);
nand U12134 (N_12134,N_11593,N_11566);
xnor U12135 (N_12135,N_11772,N_11718);
or U12136 (N_12136,N_11501,N_11529);
and U12137 (N_12137,N_11897,N_11548);
xnor U12138 (N_12138,N_11809,N_11871);
nand U12139 (N_12139,N_11621,N_11586);
or U12140 (N_12140,N_11526,N_11570);
nand U12141 (N_12141,N_11893,N_11732);
and U12142 (N_12142,N_11965,N_11672);
and U12143 (N_12143,N_11861,N_11521);
and U12144 (N_12144,N_11730,N_11583);
and U12145 (N_12145,N_11961,N_11970);
and U12146 (N_12146,N_11575,N_11918);
and U12147 (N_12147,N_11953,N_11653);
or U12148 (N_12148,N_11946,N_11722);
or U12149 (N_12149,N_11767,N_11500);
nand U12150 (N_12150,N_11948,N_11807);
nand U12151 (N_12151,N_11787,N_11654);
or U12152 (N_12152,N_11615,N_11725);
nand U12153 (N_12153,N_11974,N_11727);
nand U12154 (N_12154,N_11769,N_11627);
nor U12155 (N_12155,N_11632,N_11720);
or U12156 (N_12156,N_11574,N_11565);
nand U12157 (N_12157,N_11976,N_11564);
or U12158 (N_12158,N_11508,N_11547);
or U12159 (N_12159,N_11665,N_11753);
nand U12160 (N_12160,N_11944,N_11741);
xnor U12161 (N_12161,N_11966,N_11719);
nand U12162 (N_12162,N_11558,N_11689);
and U12163 (N_12163,N_11742,N_11671);
and U12164 (N_12164,N_11764,N_11868);
and U12165 (N_12165,N_11811,N_11592);
xor U12166 (N_12166,N_11701,N_11708);
nand U12167 (N_12167,N_11670,N_11522);
or U12168 (N_12168,N_11862,N_11968);
nor U12169 (N_12169,N_11634,N_11973);
or U12170 (N_12170,N_11791,N_11771);
and U12171 (N_12171,N_11920,N_11692);
nor U12172 (N_12172,N_11851,N_11818);
nor U12173 (N_12173,N_11602,N_11709);
and U12174 (N_12174,N_11952,N_11978);
or U12175 (N_12175,N_11663,N_11773);
or U12176 (N_12176,N_11696,N_11557);
and U12177 (N_12177,N_11706,N_11863);
and U12178 (N_12178,N_11512,N_11919);
and U12179 (N_12179,N_11652,N_11677);
or U12180 (N_12180,N_11752,N_11866);
or U12181 (N_12181,N_11542,N_11595);
xnor U12182 (N_12182,N_11581,N_11699);
nor U12183 (N_12183,N_11726,N_11605);
or U12184 (N_12184,N_11888,N_11936);
nand U12185 (N_12185,N_11700,N_11554);
nand U12186 (N_12186,N_11876,N_11525);
nor U12187 (N_12187,N_11789,N_11678);
nor U12188 (N_12188,N_11739,N_11841);
or U12189 (N_12189,N_11528,N_11680);
or U12190 (N_12190,N_11857,N_11607);
xnor U12191 (N_12191,N_11975,N_11645);
nor U12192 (N_12192,N_11800,N_11659);
nand U12193 (N_12193,N_11690,N_11723);
nor U12194 (N_12194,N_11931,N_11847);
or U12195 (N_12195,N_11987,N_11597);
or U12196 (N_12196,N_11810,N_11790);
xor U12197 (N_12197,N_11999,N_11524);
and U12198 (N_12198,N_11933,N_11553);
xnor U12199 (N_12199,N_11781,N_11667);
nand U12200 (N_12200,N_11532,N_11582);
nand U12201 (N_12201,N_11619,N_11635);
nand U12202 (N_12202,N_11836,N_11676);
nand U12203 (N_12203,N_11740,N_11691);
or U12204 (N_12204,N_11743,N_11912);
xnor U12205 (N_12205,N_11504,N_11835);
xnor U12206 (N_12206,N_11531,N_11828);
or U12207 (N_12207,N_11873,N_11830);
or U12208 (N_12208,N_11926,N_11864);
nor U12209 (N_12209,N_11650,N_11826);
and U12210 (N_12210,N_11599,N_11776);
and U12211 (N_12211,N_11890,N_11614);
and U12212 (N_12212,N_11756,N_11845);
nor U12213 (N_12213,N_11941,N_11747);
nor U12214 (N_12214,N_11921,N_11886);
or U12215 (N_12215,N_11687,N_11899);
or U12216 (N_12216,N_11662,N_11979);
nor U12217 (N_12217,N_11780,N_11681);
or U12218 (N_12218,N_11956,N_11990);
and U12219 (N_12219,N_11523,N_11712);
and U12220 (N_12220,N_11544,N_11624);
nand U12221 (N_12221,N_11674,N_11816);
nor U12222 (N_12222,N_11647,N_11852);
nand U12223 (N_12223,N_11576,N_11984);
nand U12224 (N_12224,N_11561,N_11900);
or U12225 (N_12225,N_11928,N_11892);
nand U12226 (N_12226,N_11704,N_11881);
xor U12227 (N_12227,N_11673,N_11506);
and U12228 (N_12228,N_11988,N_11846);
and U12229 (N_12229,N_11744,N_11648);
and U12230 (N_12230,N_11822,N_11517);
nand U12231 (N_12231,N_11748,N_11853);
nor U12232 (N_12232,N_11786,N_11620);
and U12233 (N_12233,N_11778,N_11788);
nor U12234 (N_12234,N_11877,N_11656);
xnor U12235 (N_12235,N_11985,N_11834);
and U12236 (N_12236,N_11537,N_11612);
and U12237 (N_12237,N_11587,N_11879);
and U12238 (N_12238,N_11556,N_11610);
nand U12239 (N_12239,N_11616,N_11782);
nor U12240 (N_12240,N_11917,N_11664);
nor U12241 (N_12241,N_11865,N_11804);
nor U12242 (N_12242,N_11907,N_11697);
nand U12243 (N_12243,N_11959,N_11626);
xor U12244 (N_12244,N_11854,N_11954);
and U12245 (N_12245,N_11538,N_11837);
or U12246 (N_12246,N_11915,N_11705);
nand U12247 (N_12247,N_11823,N_11539);
nand U12248 (N_12248,N_11983,N_11943);
nand U12249 (N_12249,N_11535,N_11511);
nand U12250 (N_12250,N_11869,N_11870);
or U12251 (N_12251,N_11902,N_11761);
or U12252 (N_12252,N_11601,N_11637);
or U12253 (N_12253,N_11577,N_11603);
and U12254 (N_12254,N_11701,N_11666);
or U12255 (N_12255,N_11518,N_11603);
nor U12256 (N_12256,N_11930,N_11904);
or U12257 (N_12257,N_11905,N_11685);
and U12258 (N_12258,N_11702,N_11661);
nand U12259 (N_12259,N_11954,N_11728);
nand U12260 (N_12260,N_11912,N_11503);
and U12261 (N_12261,N_11517,N_11894);
or U12262 (N_12262,N_11923,N_11622);
or U12263 (N_12263,N_11753,N_11681);
or U12264 (N_12264,N_11888,N_11878);
nand U12265 (N_12265,N_11632,N_11940);
xnor U12266 (N_12266,N_11914,N_11837);
or U12267 (N_12267,N_11902,N_11920);
nand U12268 (N_12268,N_11946,N_11511);
nand U12269 (N_12269,N_11977,N_11619);
nand U12270 (N_12270,N_11855,N_11951);
and U12271 (N_12271,N_11875,N_11808);
nand U12272 (N_12272,N_11737,N_11573);
nor U12273 (N_12273,N_11900,N_11876);
xnor U12274 (N_12274,N_11822,N_11996);
nand U12275 (N_12275,N_11772,N_11773);
nand U12276 (N_12276,N_11975,N_11752);
or U12277 (N_12277,N_11917,N_11937);
or U12278 (N_12278,N_11977,N_11640);
nor U12279 (N_12279,N_11559,N_11739);
nor U12280 (N_12280,N_11996,N_11943);
nor U12281 (N_12281,N_11816,N_11889);
nor U12282 (N_12282,N_11532,N_11592);
and U12283 (N_12283,N_11561,N_11612);
nor U12284 (N_12284,N_11858,N_11945);
nor U12285 (N_12285,N_11831,N_11619);
xor U12286 (N_12286,N_11896,N_11870);
or U12287 (N_12287,N_11504,N_11967);
nand U12288 (N_12288,N_11513,N_11515);
or U12289 (N_12289,N_11941,N_11522);
xnor U12290 (N_12290,N_11773,N_11754);
nand U12291 (N_12291,N_11845,N_11744);
xor U12292 (N_12292,N_11644,N_11723);
nand U12293 (N_12293,N_11620,N_11979);
or U12294 (N_12294,N_11984,N_11968);
nand U12295 (N_12295,N_11979,N_11593);
and U12296 (N_12296,N_11549,N_11838);
or U12297 (N_12297,N_11656,N_11622);
or U12298 (N_12298,N_11979,N_11998);
nand U12299 (N_12299,N_11627,N_11625);
nor U12300 (N_12300,N_11657,N_11925);
nor U12301 (N_12301,N_11870,N_11838);
nor U12302 (N_12302,N_11747,N_11817);
nand U12303 (N_12303,N_11701,N_11573);
nand U12304 (N_12304,N_11719,N_11531);
or U12305 (N_12305,N_11593,N_11704);
xnor U12306 (N_12306,N_11741,N_11639);
nand U12307 (N_12307,N_11602,N_11901);
and U12308 (N_12308,N_11702,N_11534);
or U12309 (N_12309,N_11734,N_11711);
and U12310 (N_12310,N_11901,N_11943);
xnor U12311 (N_12311,N_11525,N_11642);
or U12312 (N_12312,N_11919,N_11830);
nand U12313 (N_12313,N_11993,N_11913);
and U12314 (N_12314,N_11903,N_11841);
nor U12315 (N_12315,N_11899,N_11523);
nand U12316 (N_12316,N_11873,N_11991);
nand U12317 (N_12317,N_11998,N_11820);
or U12318 (N_12318,N_11711,N_11653);
or U12319 (N_12319,N_11941,N_11754);
xor U12320 (N_12320,N_11868,N_11862);
nor U12321 (N_12321,N_11546,N_11622);
or U12322 (N_12322,N_11800,N_11585);
or U12323 (N_12323,N_11694,N_11669);
nand U12324 (N_12324,N_11926,N_11896);
xnor U12325 (N_12325,N_11961,N_11767);
nor U12326 (N_12326,N_11717,N_11667);
and U12327 (N_12327,N_11910,N_11690);
nor U12328 (N_12328,N_11625,N_11812);
nor U12329 (N_12329,N_11992,N_11546);
nand U12330 (N_12330,N_11717,N_11859);
nand U12331 (N_12331,N_11849,N_11513);
and U12332 (N_12332,N_11870,N_11946);
nand U12333 (N_12333,N_11924,N_11949);
or U12334 (N_12334,N_11628,N_11658);
nor U12335 (N_12335,N_11577,N_11608);
nand U12336 (N_12336,N_11925,N_11999);
xor U12337 (N_12337,N_11678,N_11994);
nand U12338 (N_12338,N_11959,N_11900);
nand U12339 (N_12339,N_11545,N_11597);
or U12340 (N_12340,N_11558,N_11751);
or U12341 (N_12341,N_11625,N_11953);
or U12342 (N_12342,N_11685,N_11831);
and U12343 (N_12343,N_11540,N_11830);
and U12344 (N_12344,N_11823,N_11550);
nand U12345 (N_12345,N_11571,N_11895);
and U12346 (N_12346,N_11803,N_11827);
or U12347 (N_12347,N_11668,N_11984);
and U12348 (N_12348,N_11685,N_11977);
or U12349 (N_12349,N_11923,N_11757);
nand U12350 (N_12350,N_11977,N_11551);
xor U12351 (N_12351,N_11937,N_11869);
nor U12352 (N_12352,N_11871,N_11843);
or U12353 (N_12353,N_11916,N_11893);
or U12354 (N_12354,N_11797,N_11545);
and U12355 (N_12355,N_11827,N_11722);
and U12356 (N_12356,N_11955,N_11725);
nor U12357 (N_12357,N_11611,N_11795);
or U12358 (N_12358,N_11624,N_11737);
xor U12359 (N_12359,N_11718,N_11764);
xor U12360 (N_12360,N_11621,N_11908);
nor U12361 (N_12361,N_11733,N_11810);
nor U12362 (N_12362,N_11771,N_11908);
or U12363 (N_12363,N_11627,N_11973);
and U12364 (N_12364,N_11971,N_11976);
and U12365 (N_12365,N_11785,N_11611);
nand U12366 (N_12366,N_11878,N_11528);
xor U12367 (N_12367,N_11982,N_11858);
and U12368 (N_12368,N_11836,N_11917);
nand U12369 (N_12369,N_11693,N_11761);
nor U12370 (N_12370,N_11922,N_11760);
or U12371 (N_12371,N_11839,N_11966);
nand U12372 (N_12372,N_11631,N_11805);
or U12373 (N_12373,N_11896,N_11819);
or U12374 (N_12374,N_11853,N_11795);
xor U12375 (N_12375,N_11774,N_11621);
nor U12376 (N_12376,N_11980,N_11807);
and U12377 (N_12377,N_11851,N_11618);
and U12378 (N_12378,N_11957,N_11694);
nor U12379 (N_12379,N_11807,N_11707);
nor U12380 (N_12380,N_11630,N_11623);
nand U12381 (N_12381,N_11754,N_11838);
xnor U12382 (N_12382,N_11631,N_11890);
nor U12383 (N_12383,N_11965,N_11585);
and U12384 (N_12384,N_11598,N_11700);
nand U12385 (N_12385,N_11654,N_11681);
and U12386 (N_12386,N_11998,N_11581);
and U12387 (N_12387,N_11695,N_11765);
nor U12388 (N_12388,N_11864,N_11705);
nor U12389 (N_12389,N_11509,N_11537);
and U12390 (N_12390,N_11502,N_11768);
and U12391 (N_12391,N_11643,N_11674);
nor U12392 (N_12392,N_11644,N_11961);
and U12393 (N_12393,N_11962,N_11848);
or U12394 (N_12394,N_11947,N_11730);
nand U12395 (N_12395,N_11978,N_11780);
nand U12396 (N_12396,N_11714,N_11777);
and U12397 (N_12397,N_11809,N_11665);
or U12398 (N_12398,N_11523,N_11843);
and U12399 (N_12399,N_11979,N_11715);
or U12400 (N_12400,N_11591,N_11759);
xnor U12401 (N_12401,N_11643,N_11637);
and U12402 (N_12402,N_11803,N_11541);
nand U12403 (N_12403,N_11843,N_11693);
and U12404 (N_12404,N_11500,N_11688);
and U12405 (N_12405,N_11656,N_11687);
nand U12406 (N_12406,N_11791,N_11680);
nor U12407 (N_12407,N_11772,N_11679);
xnor U12408 (N_12408,N_11762,N_11992);
nor U12409 (N_12409,N_11860,N_11795);
or U12410 (N_12410,N_11772,N_11560);
and U12411 (N_12411,N_11866,N_11572);
or U12412 (N_12412,N_11791,N_11635);
and U12413 (N_12413,N_11625,N_11570);
nor U12414 (N_12414,N_11788,N_11792);
or U12415 (N_12415,N_11749,N_11629);
or U12416 (N_12416,N_11572,N_11861);
xnor U12417 (N_12417,N_11769,N_11903);
nand U12418 (N_12418,N_11707,N_11849);
nor U12419 (N_12419,N_11672,N_11541);
nand U12420 (N_12420,N_11737,N_11633);
and U12421 (N_12421,N_11674,N_11583);
xor U12422 (N_12422,N_11905,N_11669);
nand U12423 (N_12423,N_11988,N_11640);
xnor U12424 (N_12424,N_11504,N_11848);
nand U12425 (N_12425,N_11678,N_11865);
nand U12426 (N_12426,N_11830,N_11702);
and U12427 (N_12427,N_11627,N_11743);
or U12428 (N_12428,N_11555,N_11763);
nor U12429 (N_12429,N_11840,N_11659);
nand U12430 (N_12430,N_11913,N_11517);
and U12431 (N_12431,N_11895,N_11551);
or U12432 (N_12432,N_11912,N_11575);
nor U12433 (N_12433,N_11745,N_11577);
nand U12434 (N_12434,N_11695,N_11945);
nand U12435 (N_12435,N_11825,N_11651);
and U12436 (N_12436,N_11740,N_11678);
and U12437 (N_12437,N_11949,N_11962);
nand U12438 (N_12438,N_11896,N_11803);
nor U12439 (N_12439,N_11949,N_11742);
nor U12440 (N_12440,N_11575,N_11654);
and U12441 (N_12441,N_11982,N_11545);
and U12442 (N_12442,N_11533,N_11810);
xnor U12443 (N_12443,N_11975,N_11689);
nor U12444 (N_12444,N_11804,N_11579);
nor U12445 (N_12445,N_11704,N_11656);
xnor U12446 (N_12446,N_11728,N_11572);
nand U12447 (N_12447,N_11691,N_11737);
nor U12448 (N_12448,N_11780,N_11660);
and U12449 (N_12449,N_11529,N_11765);
and U12450 (N_12450,N_11656,N_11757);
nor U12451 (N_12451,N_11884,N_11626);
nor U12452 (N_12452,N_11913,N_11785);
nor U12453 (N_12453,N_11792,N_11928);
or U12454 (N_12454,N_11898,N_11809);
or U12455 (N_12455,N_11733,N_11912);
nand U12456 (N_12456,N_11995,N_11920);
nand U12457 (N_12457,N_11837,N_11955);
and U12458 (N_12458,N_11802,N_11865);
xor U12459 (N_12459,N_11879,N_11847);
or U12460 (N_12460,N_11553,N_11673);
nor U12461 (N_12461,N_11993,N_11619);
or U12462 (N_12462,N_11960,N_11662);
xor U12463 (N_12463,N_11630,N_11851);
nor U12464 (N_12464,N_11685,N_11828);
and U12465 (N_12465,N_11735,N_11669);
nor U12466 (N_12466,N_11637,N_11850);
nand U12467 (N_12467,N_11880,N_11855);
nand U12468 (N_12468,N_11814,N_11815);
xor U12469 (N_12469,N_11918,N_11968);
or U12470 (N_12470,N_11543,N_11540);
nand U12471 (N_12471,N_11629,N_11951);
or U12472 (N_12472,N_11833,N_11700);
nor U12473 (N_12473,N_11951,N_11502);
nor U12474 (N_12474,N_11953,N_11623);
xor U12475 (N_12475,N_11660,N_11668);
xnor U12476 (N_12476,N_11778,N_11843);
nor U12477 (N_12477,N_11744,N_11665);
nor U12478 (N_12478,N_11933,N_11946);
xor U12479 (N_12479,N_11712,N_11945);
or U12480 (N_12480,N_11570,N_11721);
nor U12481 (N_12481,N_11786,N_11616);
and U12482 (N_12482,N_11589,N_11604);
nor U12483 (N_12483,N_11552,N_11818);
nor U12484 (N_12484,N_11875,N_11680);
or U12485 (N_12485,N_11910,N_11639);
nor U12486 (N_12486,N_11528,N_11844);
nor U12487 (N_12487,N_11678,N_11549);
and U12488 (N_12488,N_11683,N_11539);
and U12489 (N_12489,N_11698,N_11786);
nand U12490 (N_12490,N_11999,N_11858);
nand U12491 (N_12491,N_11904,N_11584);
nand U12492 (N_12492,N_11645,N_11765);
nand U12493 (N_12493,N_11781,N_11711);
or U12494 (N_12494,N_11986,N_11628);
or U12495 (N_12495,N_11760,N_11668);
nor U12496 (N_12496,N_11964,N_11533);
and U12497 (N_12497,N_11902,N_11659);
or U12498 (N_12498,N_11576,N_11579);
nand U12499 (N_12499,N_11741,N_11592);
xor U12500 (N_12500,N_12291,N_12382);
nor U12501 (N_12501,N_12015,N_12127);
nand U12502 (N_12502,N_12128,N_12087);
or U12503 (N_12503,N_12223,N_12268);
nand U12504 (N_12504,N_12316,N_12234);
nor U12505 (N_12505,N_12470,N_12424);
or U12506 (N_12506,N_12197,N_12454);
nand U12507 (N_12507,N_12373,N_12488);
or U12508 (N_12508,N_12134,N_12032);
nand U12509 (N_12509,N_12275,N_12473);
nand U12510 (N_12510,N_12031,N_12072);
xor U12511 (N_12511,N_12352,N_12126);
nand U12512 (N_12512,N_12188,N_12262);
xor U12513 (N_12513,N_12491,N_12025);
or U12514 (N_12514,N_12220,N_12034);
nor U12515 (N_12515,N_12091,N_12172);
or U12516 (N_12516,N_12350,N_12017);
or U12517 (N_12517,N_12214,N_12483);
nor U12518 (N_12518,N_12104,N_12313);
and U12519 (N_12519,N_12460,N_12187);
nor U12520 (N_12520,N_12252,N_12322);
nand U12521 (N_12521,N_12437,N_12293);
nor U12522 (N_12522,N_12137,N_12289);
and U12523 (N_12523,N_12173,N_12415);
nor U12524 (N_12524,N_12412,N_12113);
or U12525 (N_12525,N_12086,N_12056);
xnor U12526 (N_12526,N_12281,N_12122);
xor U12527 (N_12527,N_12013,N_12057);
or U12528 (N_12528,N_12431,N_12182);
xor U12529 (N_12529,N_12118,N_12273);
xnor U12530 (N_12530,N_12368,N_12452);
nor U12531 (N_12531,N_12230,N_12354);
xnor U12532 (N_12532,N_12084,N_12195);
or U12533 (N_12533,N_12233,N_12325);
or U12534 (N_12534,N_12458,N_12008);
and U12535 (N_12535,N_12436,N_12474);
nand U12536 (N_12536,N_12496,N_12097);
nor U12537 (N_12537,N_12406,N_12255);
nand U12538 (N_12538,N_12043,N_12472);
nand U12539 (N_12539,N_12090,N_12468);
xor U12540 (N_12540,N_12278,N_12124);
or U12541 (N_12541,N_12399,N_12475);
nor U12542 (N_12542,N_12400,N_12413);
and U12543 (N_12543,N_12235,N_12272);
nand U12544 (N_12544,N_12421,N_12184);
nor U12545 (N_12545,N_12001,N_12238);
nor U12546 (N_12546,N_12239,N_12283);
or U12547 (N_12547,N_12052,N_12408);
nand U12548 (N_12548,N_12388,N_12381);
and U12549 (N_12549,N_12221,N_12455);
nand U12550 (N_12550,N_12467,N_12242);
or U12551 (N_12551,N_12375,N_12355);
nand U12552 (N_12552,N_12147,N_12301);
nor U12553 (N_12553,N_12329,N_12027);
nor U12554 (N_12554,N_12318,N_12397);
nor U12555 (N_12555,N_12103,N_12170);
nor U12556 (N_12556,N_12411,N_12380);
xor U12557 (N_12557,N_12067,N_12246);
nand U12558 (N_12558,N_12088,N_12139);
or U12559 (N_12559,N_12304,N_12152);
nand U12560 (N_12560,N_12420,N_12277);
or U12561 (N_12561,N_12335,N_12331);
nor U12562 (N_12562,N_12306,N_12346);
nand U12563 (N_12563,N_12156,N_12100);
nand U12564 (N_12564,N_12218,N_12284);
nand U12565 (N_12565,N_12180,N_12059);
xnor U12566 (N_12566,N_12204,N_12224);
nor U12567 (N_12567,N_12058,N_12073);
xor U12568 (N_12568,N_12123,N_12146);
xnor U12569 (N_12569,N_12041,N_12256);
nand U12570 (N_12570,N_12495,N_12062);
xor U12571 (N_12571,N_12480,N_12226);
nand U12572 (N_12572,N_12111,N_12105);
nand U12573 (N_12573,N_12457,N_12066);
nand U12574 (N_12574,N_12063,N_12076);
xnor U12575 (N_12575,N_12045,N_12002);
or U12576 (N_12576,N_12075,N_12334);
xnor U12577 (N_12577,N_12494,N_12430);
nor U12578 (N_12578,N_12264,N_12393);
or U12579 (N_12579,N_12309,N_12130);
nand U12580 (N_12580,N_12083,N_12418);
xnor U12581 (N_12581,N_12014,N_12163);
or U12582 (N_12582,N_12094,N_12257);
or U12583 (N_12583,N_12006,N_12295);
and U12584 (N_12584,N_12328,N_12395);
or U12585 (N_12585,N_12243,N_12018);
nor U12586 (N_12586,N_12024,N_12080);
or U12587 (N_12587,N_12410,N_12282);
or U12588 (N_12588,N_12148,N_12074);
and U12589 (N_12589,N_12011,N_12225);
xnor U12590 (N_12590,N_12435,N_12198);
or U12591 (N_12591,N_12308,N_12070);
nand U12592 (N_12592,N_12336,N_12497);
and U12593 (N_12593,N_12287,N_12489);
and U12594 (N_12594,N_12106,N_12216);
nand U12595 (N_12595,N_12029,N_12060);
or U12596 (N_12596,N_12009,N_12093);
and U12597 (N_12597,N_12053,N_12349);
xnor U12598 (N_12598,N_12196,N_12324);
nor U12599 (N_12599,N_12244,N_12177);
nor U12600 (N_12600,N_12466,N_12033);
or U12601 (N_12601,N_12427,N_12389);
and U12602 (N_12602,N_12199,N_12071);
nand U12603 (N_12603,N_12299,N_12274);
nor U12604 (N_12604,N_12138,N_12432);
nor U12605 (N_12605,N_12000,N_12102);
nand U12606 (N_12606,N_12160,N_12020);
and U12607 (N_12607,N_12332,N_12116);
and U12608 (N_12608,N_12157,N_12377);
and U12609 (N_12609,N_12471,N_12323);
nor U12610 (N_12610,N_12085,N_12476);
nor U12611 (N_12611,N_12405,N_12099);
or U12612 (N_12612,N_12064,N_12108);
and U12613 (N_12613,N_12068,N_12231);
and U12614 (N_12614,N_12372,N_12341);
or U12615 (N_12615,N_12478,N_12181);
or U12616 (N_12616,N_12499,N_12171);
or U12617 (N_12617,N_12007,N_12167);
or U12618 (N_12618,N_12319,N_12327);
nand U12619 (N_12619,N_12178,N_12169);
and U12620 (N_12620,N_12036,N_12358);
or U12621 (N_12621,N_12485,N_12449);
and U12622 (N_12622,N_12433,N_12371);
nand U12623 (N_12623,N_12096,N_12054);
nor U12624 (N_12624,N_12311,N_12021);
or U12625 (N_12625,N_12426,N_12260);
or U12626 (N_12626,N_12151,N_12101);
nor U12627 (N_12627,N_12132,N_12343);
nand U12628 (N_12628,N_12205,N_12175);
nor U12629 (N_12629,N_12249,N_12383);
nor U12630 (N_12630,N_12445,N_12145);
and U12631 (N_12631,N_12237,N_12367);
and U12632 (N_12632,N_12398,N_12229);
and U12633 (N_12633,N_12303,N_12129);
nand U12634 (N_12634,N_12276,N_12114);
or U12635 (N_12635,N_12258,N_12360);
and U12636 (N_12636,N_12357,N_12493);
nor U12637 (N_12637,N_12125,N_12290);
nor U12638 (N_12638,N_12351,N_12241);
and U12639 (N_12639,N_12030,N_12259);
nand U12640 (N_12640,N_12403,N_12044);
nand U12641 (N_12641,N_12402,N_12285);
nor U12642 (N_12642,N_12210,N_12374);
xnor U12643 (N_12643,N_12247,N_12047);
xor U12644 (N_12644,N_12297,N_12463);
xnor U12645 (N_12645,N_12305,N_12442);
nor U12646 (N_12646,N_12370,N_12185);
or U12647 (N_12647,N_12330,N_12378);
nor U12648 (N_12648,N_12314,N_12340);
and U12649 (N_12649,N_12345,N_12046);
and U12650 (N_12650,N_12443,N_12095);
nand U12651 (N_12651,N_12166,N_12089);
and U12652 (N_12652,N_12191,N_12174);
or U12653 (N_12653,N_12004,N_12143);
nand U12654 (N_12654,N_12444,N_12190);
nor U12655 (N_12655,N_12207,N_12219);
nor U12656 (N_12656,N_12040,N_12019);
or U12657 (N_12657,N_12065,N_12133);
and U12658 (N_12658,N_12390,N_12016);
or U12659 (N_12659,N_12051,N_12194);
and U12660 (N_12660,N_12200,N_12456);
and U12661 (N_12661,N_12280,N_12356);
or U12662 (N_12662,N_12037,N_12212);
or U12663 (N_12663,N_12079,N_12055);
and U12664 (N_12664,N_12479,N_12213);
nand U12665 (N_12665,N_12447,N_12154);
or U12666 (N_12666,N_12337,N_12039);
nor U12667 (N_12667,N_12211,N_12179);
or U12668 (N_12668,N_12288,N_12161);
or U12669 (N_12669,N_12153,N_12344);
and U12670 (N_12670,N_12005,N_12441);
and U12671 (N_12671,N_12266,N_12158);
nor U12672 (N_12672,N_12168,N_12003);
and U12673 (N_12673,N_12369,N_12144);
or U12674 (N_12674,N_12365,N_12404);
and U12675 (N_12675,N_12164,N_12050);
and U12676 (N_12676,N_12379,N_12286);
nand U12677 (N_12677,N_12353,N_12092);
and U12678 (N_12678,N_12162,N_12081);
or U12679 (N_12679,N_12385,N_12119);
nor U12680 (N_12680,N_12135,N_12279);
and U12681 (N_12681,N_12326,N_12061);
or U12682 (N_12682,N_12296,N_12176);
xnor U12683 (N_12683,N_12098,N_12451);
nor U12684 (N_12684,N_12023,N_12010);
or U12685 (N_12685,N_12392,N_12348);
nor U12686 (N_12686,N_12434,N_12208);
and U12687 (N_12687,N_12416,N_12384);
nor U12688 (N_12688,N_12417,N_12267);
nor U12689 (N_12689,N_12333,N_12131);
or U12690 (N_12690,N_12265,N_12484);
and U12691 (N_12691,N_12469,N_12253);
and U12692 (N_12692,N_12407,N_12201);
and U12693 (N_12693,N_12109,N_12362);
and U12694 (N_12694,N_12142,N_12035);
nand U12695 (N_12695,N_12461,N_12248);
or U12696 (N_12696,N_12477,N_12387);
nand U12697 (N_12697,N_12361,N_12206);
or U12698 (N_12698,N_12183,N_12342);
nor U12699 (N_12699,N_12026,N_12302);
nor U12700 (N_12700,N_12165,N_12292);
nor U12701 (N_12701,N_12453,N_12481);
or U12702 (N_12702,N_12209,N_12077);
and U12703 (N_12703,N_12315,N_12121);
nand U12704 (N_12704,N_12347,N_12192);
nor U12705 (N_12705,N_12492,N_12446);
nand U12706 (N_12706,N_12320,N_12439);
or U12707 (N_12707,N_12391,N_12155);
nand U12708 (N_12708,N_12422,N_12269);
nor U12709 (N_12709,N_12498,N_12376);
or U12710 (N_12710,N_12112,N_12012);
or U12711 (N_12711,N_12310,N_12465);
or U12712 (N_12712,N_12240,N_12261);
nand U12713 (N_12713,N_12042,N_12366);
and U12714 (N_12714,N_12359,N_12082);
nor U12715 (N_12715,N_12312,N_12236);
or U12716 (N_12716,N_12186,N_12401);
nand U12717 (N_12717,N_12222,N_12217);
nor U12718 (N_12718,N_12450,N_12394);
or U12719 (N_12719,N_12189,N_12141);
or U12720 (N_12720,N_12423,N_12049);
or U12721 (N_12721,N_12202,N_12448);
xor U12722 (N_12722,N_12298,N_12364);
nand U12723 (N_12723,N_12300,N_12215);
nand U12724 (N_12724,N_12459,N_12232);
xnor U12725 (N_12725,N_12117,N_12120);
and U12726 (N_12726,N_12245,N_12321);
and U12727 (N_12727,N_12251,N_12363);
nor U12728 (N_12728,N_12294,N_12409);
or U12729 (N_12729,N_12428,N_12140);
nand U12730 (N_12730,N_12203,N_12317);
or U12731 (N_12731,N_12490,N_12107);
nor U12732 (N_12732,N_12038,N_12048);
and U12733 (N_12733,N_12078,N_12149);
nor U12734 (N_12734,N_12270,N_12115);
and U12735 (N_12735,N_12464,N_12396);
and U12736 (N_12736,N_12429,N_12271);
and U12737 (N_12737,N_12419,N_12386);
nand U12738 (N_12738,N_12028,N_12159);
xor U12739 (N_12739,N_12250,N_12414);
and U12740 (N_12740,N_12440,N_12022);
or U12741 (N_12741,N_12487,N_12069);
and U12742 (N_12742,N_12263,N_12339);
or U12743 (N_12743,N_12110,N_12254);
nor U12744 (N_12744,N_12462,N_12486);
nand U12745 (N_12745,N_12338,N_12227);
nor U12746 (N_12746,N_12482,N_12438);
nand U12747 (N_12747,N_12150,N_12136);
nor U12748 (N_12748,N_12193,N_12228);
nand U12749 (N_12749,N_12425,N_12307);
or U12750 (N_12750,N_12291,N_12180);
nand U12751 (N_12751,N_12173,N_12440);
and U12752 (N_12752,N_12211,N_12493);
and U12753 (N_12753,N_12022,N_12283);
or U12754 (N_12754,N_12255,N_12121);
nor U12755 (N_12755,N_12485,N_12230);
and U12756 (N_12756,N_12082,N_12261);
xor U12757 (N_12757,N_12293,N_12278);
xor U12758 (N_12758,N_12050,N_12173);
or U12759 (N_12759,N_12173,N_12353);
and U12760 (N_12760,N_12091,N_12394);
nand U12761 (N_12761,N_12431,N_12040);
nor U12762 (N_12762,N_12122,N_12340);
nor U12763 (N_12763,N_12297,N_12479);
or U12764 (N_12764,N_12039,N_12122);
nor U12765 (N_12765,N_12498,N_12063);
and U12766 (N_12766,N_12466,N_12250);
xnor U12767 (N_12767,N_12397,N_12488);
nor U12768 (N_12768,N_12256,N_12463);
xor U12769 (N_12769,N_12376,N_12134);
nand U12770 (N_12770,N_12179,N_12435);
nand U12771 (N_12771,N_12107,N_12489);
nand U12772 (N_12772,N_12169,N_12315);
nor U12773 (N_12773,N_12363,N_12324);
and U12774 (N_12774,N_12000,N_12377);
nor U12775 (N_12775,N_12470,N_12240);
nor U12776 (N_12776,N_12216,N_12041);
nor U12777 (N_12777,N_12173,N_12297);
nand U12778 (N_12778,N_12255,N_12134);
and U12779 (N_12779,N_12237,N_12100);
nor U12780 (N_12780,N_12380,N_12457);
and U12781 (N_12781,N_12475,N_12427);
nor U12782 (N_12782,N_12237,N_12378);
xor U12783 (N_12783,N_12082,N_12225);
or U12784 (N_12784,N_12444,N_12462);
or U12785 (N_12785,N_12453,N_12127);
and U12786 (N_12786,N_12287,N_12112);
nand U12787 (N_12787,N_12335,N_12383);
or U12788 (N_12788,N_12415,N_12477);
nor U12789 (N_12789,N_12148,N_12451);
nand U12790 (N_12790,N_12023,N_12025);
xnor U12791 (N_12791,N_12381,N_12182);
nand U12792 (N_12792,N_12348,N_12465);
and U12793 (N_12793,N_12229,N_12012);
nor U12794 (N_12794,N_12330,N_12404);
and U12795 (N_12795,N_12378,N_12259);
and U12796 (N_12796,N_12387,N_12175);
nand U12797 (N_12797,N_12327,N_12175);
and U12798 (N_12798,N_12334,N_12412);
or U12799 (N_12799,N_12417,N_12019);
nor U12800 (N_12800,N_12070,N_12203);
nand U12801 (N_12801,N_12304,N_12151);
nor U12802 (N_12802,N_12200,N_12448);
or U12803 (N_12803,N_12192,N_12070);
and U12804 (N_12804,N_12401,N_12333);
and U12805 (N_12805,N_12446,N_12193);
xor U12806 (N_12806,N_12143,N_12406);
and U12807 (N_12807,N_12349,N_12472);
and U12808 (N_12808,N_12089,N_12418);
nand U12809 (N_12809,N_12393,N_12280);
xor U12810 (N_12810,N_12186,N_12253);
nor U12811 (N_12811,N_12377,N_12022);
nand U12812 (N_12812,N_12365,N_12097);
nand U12813 (N_12813,N_12143,N_12050);
nor U12814 (N_12814,N_12218,N_12263);
nor U12815 (N_12815,N_12291,N_12024);
and U12816 (N_12816,N_12414,N_12416);
or U12817 (N_12817,N_12459,N_12127);
or U12818 (N_12818,N_12487,N_12169);
and U12819 (N_12819,N_12250,N_12074);
or U12820 (N_12820,N_12237,N_12356);
and U12821 (N_12821,N_12232,N_12356);
nand U12822 (N_12822,N_12460,N_12205);
or U12823 (N_12823,N_12343,N_12058);
nand U12824 (N_12824,N_12303,N_12072);
and U12825 (N_12825,N_12347,N_12047);
and U12826 (N_12826,N_12210,N_12234);
nor U12827 (N_12827,N_12296,N_12107);
or U12828 (N_12828,N_12101,N_12472);
or U12829 (N_12829,N_12240,N_12226);
or U12830 (N_12830,N_12185,N_12025);
xor U12831 (N_12831,N_12018,N_12483);
nor U12832 (N_12832,N_12423,N_12078);
and U12833 (N_12833,N_12096,N_12479);
xnor U12834 (N_12834,N_12146,N_12299);
nor U12835 (N_12835,N_12333,N_12397);
and U12836 (N_12836,N_12141,N_12407);
nand U12837 (N_12837,N_12288,N_12099);
or U12838 (N_12838,N_12281,N_12403);
or U12839 (N_12839,N_12257,N_12416);
or U12840 (N_12840,N_12492,N_12030);
or U12841 (N_12841,N_12464,N_12407);
or U12842 (N_12842,N_12375,N_12127);
and U12843 (N_12843,N_12161,N_12044);
nor U12844 (N_12844,N_12237,N_12073);
nor U12845 (N_12845,N_12026,N_12327);
xnor U12846 (N_12846,N_12086,N_12062);
or U12847 (N_12847,N_12059,N_12393);
or U12848 (N_12848,N_12268,N_12481);
nor U12849 (N_12849,N_12238,N_12206);
nor U12850 (N_12850,N_12294,N_12114);
nor U12851 (N_12851,N_12271,N_12315);
nor U12852 (N_12852,N_12367,N_12252);
and U12853 (N_12853,N_12330,N_12450);
nor U12854 (N_12854,N_12005,N_12473);
and U12855 (N_12855,N_12002,N_12300);
and U12856 (N_12856,N_12065,N_12119);
nand U12857 (N_12857,N_12109,N_12281);
nand U12858 (N_12858,N_12352,N_12083);
and U12859 (N_12859,N_12465,N_12356);
nor U12860 (N_12860,N_12051,N_12078);
nor U12861 (N_12861,N_12453,N_12244);
or U12862 (N_12862,N_12331,N_12145);
or U12863 (N_12863,N_12433,N_12044);
nor U12864 (N_12864,N_12378,N_12048);
nor U12865 (N_12865,N_12056,N_12006);
nand U12866 (N_12866,N_12239,N_12370);
nand U12867 (N_12867,N_12283,N_12137);
nand U12868 (N_12868,N_12241,N_12349);
or U12869 (N_12869,N_12237,N_12342);
nand U12870 (N_12870,N_12207,N_12087);
and U12871 (N_12871,N_12103,N_12067);
nand U12872 (N_12872,N_12446,N_12161);
and U12873 (N_12873,N_12497,N_12149);
and U12874 (N_12874,N_12370,N_12494);
or U12875 (N_12875,N_12063,N_12382);
or U12876 (N_12876,N_12458,N_12059);
and U12877 (N_12877,N_12105,N_12263);
nand U12878 (N_12878,N_12285,N_12253);
xnor U12879 (N_12879,N_12104,N_12358);
and U12880 (N_12880,N_12392,N_12432);
or U12881 (N_12881,N_12031,N_12009);
nor U12882 (N_12882,N_12181,N_12091);
and U12883 (N_12883,N_12361,N_12454);
nand U12884 (N_12884,N_12142,N_12294);
and U12885 (N_12885,N_12423,N_12454);
or U12886 (N_12886,N_12306,N_12029);
nor U12887 (N_12887,N_12182,N_12255);
and U12888 (N_12888,N_12073,N_12088);
nand U12889 (N_12889,N_12472,N_12272);
nor U12890 (N_12890,N_12418,N_12211);
or U12891 (N_12891,N_12315,N_12460);
nand U12892 (N_12892,N_12492,N_12088);
nand U12893 (N_12893,N_12069,N_12374);
xor U12894 (N_12894,N_12351,N_12325);
nor U12895 (N_12895,N_12218,N_12296);
and U12896 (N_12896,N_12177,N_12216);
xnor U12897 (N_12897,N_12150,N_12110);
and U12898 (N_12898,N_12008,N_12097);
nand U12899 (N_12899,N_12193,N_12217);
nand U12900 (N_12900,N_12164,N_12456);
or U12901 (N_12901,N_12296,N_12445);
nor U12902 (N_12902,N_12202,N_12001);
nor U12903 (N_12903,N_12207,N_12003);
xnor U12904 (N_12904,N_12154,N_12064);
nor U12905 (N_12905,N_12026,N_12439);
nor U12906 (N_12906,N_12012,N_12175);
and U12907 (N_12907,N_12099,N_12210);
nor U12908 (N_12908,N_12079,N_12307);
nor U12909 (N_12909,N_12386,N_12474);
xor U12910 (N_12910,N_12160,N_12059);
and U12911 (N_12911,N_12276,N_12083);
nand U12912 (N_12912,N_12113,N_12065);
xor U12913 (N_12913,N_12287,N_12142);
nor U12914 (N_12914,N_12406,N_12285);
xor U12915 (N_12915,N_12352,N_12096);
nor U12916 (N_12916,N_12060,N_12142);
and U12917 (N_12917,N_12422,N_12410);
nand U12918 (N_12918,N_12001,N_12227);
nor U12919 (N_12919,N_12432,N_12055);
and U12920 (N_12920,N_12419,N_12428);
and U12921 (N_12921,N_12397,N_12358);
or U12922 (N_12922,N_12305,N_12449);
and U12923 (N_12923,N_12364,N_12038);
or U12924 (N_12924,N_12145,N_12450);
or U12925 (N_12925,N_12338,N_12377);
xnor U12926 (N_12926,N_12248,N_12285);
nand U12927 (N_12927,N_12385,N_12213);
nor U12928 (N_12928,N_12184,N_12257);
nand U12929 (N_12929,N_12304,N_12173);
nor U12930 (N_12930,N_12197,N_12192);
nor U12931 (N_12931,N_12078,N_12337);
and U12932 (N_12932,N_12045,N_12346);
or U12933 (N_12933,N_12318,N_12235);
or U12934 (N_12934,N_12479,N_12469);
and U12935 (N_12935,N_12381,N_12236);
nor U12936 (N_12936,N_12355,N_12243);
nand U12937 (N_12937,N_12417,N_12116);
and U12938 (N_12938,N_12018,N_12375);
nand U12939 (N_12939,N_12263,N_12042);
and U12940 (N_12940,N_12394,N_12029);
or U12941 (N_12941,N_12131,N_12066);
nand U12942 (N_12942,N_12004,N_12476);
xor U12943 (N_12943,N_12328,N_12222);
xnor U12944 (N_12944,N_12378,N_12123);
or U12945 (N_12945,N_12075,N_12274);
xor U12946 (N_12946,N_12481,N_12260);
xnor U12947 (N_12947,N_12213,N_12054);
nor U12948 (N_12948,N_12241,N_12112);
nor U12949 (N_12949,N_12448,N_12113);
xnor U12950 (N_12950,N_12163,N_12355);
nand U12951 (N_12951,N_12202,N_12477);
nor U12952 (N_12952,N_12426,N_12133);
nor U12953 (N_12953,N_12429,N_12378);
nand U12954 (N_12954,N_12093,N_12259);
nor U12955 (N_12955,N_12242,N_12227);
or U12956 (N_12956,N_12485,N_12046);
nor U12957 (N_12957,N_12035,N_12247);
and U12958 (N_12958,N_12228,N_12090);
nand U12959 (N_12959,N_12389,N_12356);
and U12960 (N_12960,N_12210,N_12218);
xnor U12961 (N_12961,N_12144,N_12250);
nand U12962 (N_12962,N_12132,N_12056);
or U12963 (N_12963,N_12276,N_12375);
xor U12964 (N_12964,N_12053,N_12417);
or U12965 (N_12965,N_12492,N_12479);
or U12966 (N_12966,N_12192,N_12276);
nor U12967 (N_12967,N_12150,N_12225);
nand U12968 (N_12968,N_12192,N_12494);
xnor U12969 (N_12969,N_12003,N_12027);
xor U12970 (N_12970,N_12476,N_12293);
xnor U12971 (N_12971,N_12484,N_12094);
and U12972 (N_12972,N_12151,N_12234);
nor U12973 (N_12973,N_12109,N_12304);
nand U12974 (N_12974,N_12115,N_12386);
nand U12975 (N_12975,N_12092,N_12405);
xor U12976 (N_12976,N_12196,N_12494);
nor U12977 (N_12977,N_12256,N_12405);
nand U12978 (N_12978,N_12028,N_12318);
nand U12979 (N_12979,N_12349,N_12395);
nand U12980 (N_12980,N_12215,N_12434);
nand U12981 (N_12981,N_12419,N_12219);
nor U12982 (N_12982,N_12008,N_12306);
xor U12983 (N_12983,N_12177,N_12373);
nor U12984 (N_12984,N_12164,N_12189);
or U12985 (N_12985,N_12003,N_12101);
or U12986 (N_12986,N_12049,N_12088);
xor U12987 (N_12987,N_12251,N_12207);
and U12988 (N_12988,N_12471,N_12350);
nor U12989 (N_12989,N_12002,N_12284);
nand U12990 (N_12990,N_12421,N_12243);
nand U12991 (N_12991,N_12106,N_12448);
or U12992 (N_12992,N_12294,N_12006);
or U12993 (N_12993,N_12312,N_12233);
or U12994 (N_12994,N_12011,N_12449);
or U12995 (N_12995,N_12123,N_12352);
nand U12996 (N_12996,N_12061,N_12319);
nor U12997 (N_12997,N_12235,N_12244);
nand U12998 (N_12998,N_12095,N_12195);
nand U12999 (N_12999,N_12170,N_12025);
nand U13000 (N_13000,N_12758,N_12751);
or U13001 (N_13001,N_12975,N_12952);
nor U13002 (N_13002,N_12505,N_12523);
or U13003 (N_13003,N_12926,N_12675);
xor U13004 (N_13004,N_12599,N_12970);
nor U13005 (N_13005,N_12673,N_12663);
nor U13006 (N_13006,N_12982,N_12959);
or U13007 (N_13007,N_12942,N_12692);
nand U13008 (N_13008,N_12649,N_12911);
or U13009 (N_13009,N_12567,N_12923);
nand U13010 (N_13010,N_12813,N_12754);
nand U13011 (N_13011,N_12698,N_12576);
nand U13012 (N_13012,N_12527,N_12955);
nor U13013 (N_13013,N_12829,N_12973);
nor U13014 (N_13014,N_12849,N_12986);
nand U13015 (N_13015,N_12786,N_12680);
nor U13016 (N_13016,N_12723,N_12859);
nor U13017 (N_13017,N_12757,N_12634);
or U13018 (N_13018,N_12831,N_12655);
and U13019 (N_13019,N_12553,N_12857);
or U13020 (N_13020,N_12517,N_12594);
or U13021 (N_13021,N_12503,N_12795);
and U13022 (N_13022,N_12610,N_12854);
nand U13023 (N_13023,N_12941,N_12546);
or U13024 (N_13024,N_12860,N_12746);
and U13025 (N_13025,N_12668,N_12507);
nand U13026 (N_13026,N_12731,N_12619);
xnor U13027 (N_13027,N_12647,N_12685);
nor U13028 (N_13028,N_12824,N_12541);
nor U13029 (N_13029,N_12883,N_12889);
xnor U13030 (N_13030,N_12928,N_12865);
xor U13031 (N_13031,N_12686,N_12721);
and U13032 (N_13032,N_12535,N_12547);
and U13033 (N_13033,N_12598,N_12794);
and U13034 (N_13034,N_12738,N_12608);
or U13035 (N_13035,N_12729,N_12908);
xor U13036 (N_13036,N_12999,N_12814);
and U13037 (N_13037,N_12533,N_12819);
and U13038 (N_13038,N_12717,N_12585);
or U13039 (N_13039,N_12910,N_12569);
or U13040 (N_13040,N_12804,N_12590);
and U13041 (N_13041,N_12690,N_12994);
nor U13042 (N_13042,N_12519,N_12811);
nand U13043 (N_13043,N_12642,N_12932);
xor U13044 (N_13044,N_12631,N_12550);
nor U13045 (N_13045,N_12575,N_12909);
nor U13046 (N_13046,N_12633,N_12841);
nand U13047 (N_13047,N_12676,N_12895);
and U13048 (N_13048,N_12727,N_12753);
or U13049 (N_13049,N_12520,N_12666);
and U13050 (N_13050,N_12915,N_12810);
nand U13051 (N_13051,N_12630,N_12776);
and U13052 (N_13052,N_12705,N_12899);
or U13053 (N_13053,N_12874,N_12875);
nor U13054 (N_13054,N_12992,N_12635);
nand U13055 (N_13055,N_12760,N_12922);
and U13056 (N_13056,N_12584,N_12780);
and U13057 (N_13057,N_12512,N_12548);
nand U13058 (N_13058,N_12582,N_12769);
nor U13059 (N_13059,N_12848,N_12704);
xnor U13060 (N_13060,N_12531,N_12904);
nor U13061 (N_13061,N_12532,N_12715);
or U13062 (N_13062,N_12568,N_12924);
and U13063 (N_13063,N_12872,N_12658);
and U13064 (N_13064,N_12681,N_12591);
nand U13065 (N_13065,N_12534,N_12967);
or U13066 (N_13066,N_12894,N_12931);
nand U13067 (N_13067,N_12890,N_12913);
nor U13068 (N_13068,N_12595,N_12820);
nor U13069 (N_13069,N_12678,N_12544);
nor U13070 (N_13070,N_12998,N_12559);
or U13071 (N_13071,N_12993,N_12643);
nor U13072 (N_13072,N_12933,N_12538);
nand U13073 (N_13073,N_12748,N_12825);
or U13074 (N_13074,N_12656,N_12578);
and U13075 (N_13075,N_12732,N_12991);
and U13076 (N_13076,N_12510,N_12806);
nor U13077 (N_13077,N_12912,N_12718);
or U13078 (N_13078,N_12774,N_12525);
nand U13079 (N_13079,N_12834,N_12611);
and U13080 (N_13080,N_12867,N_12572);
or U13081 (N_13081,N_12793,N_12817);
nor U13082 (N_13082,N_12551,N_12801);
nand U13083 (N_13083,N_12522,N_12501);
nor U13084 (N_13084,N_12682,N_12963);
or U13085 (N_13085,N_12896,N_12845);
and U13086 (N_13086,N_12511,N_12798);
or U13087 (N_13087,N_12502,N_12981);
nor U13088 (N_13088,N_12773,N_12956);
nor U13089 (N_13089,N_12800,N_12891);
nand U13090 (N_13090,N_12778,N_12830);
nor U13091 (N_13091,N_12976,N_12962);
nor U13092 (N_13092,N_12871,N_12724);
and U13093 (N_13093,N_12927,N_12752);
nand U13094 (N_13094,N_12821,N_12742);
or U13095 (N_13095,N_12671,N_12636);
nor U13096 (N_13096,N_12638,N_12646);
or U13097 (N_13097,N_12518,N_12540);
nor U13098 (N_13098,N_12564,N_12737);
or U13099 (N_13099,N_12882,N_12526);
or U13100 (N_13100,N_12743,N_12697);
and U13101 (N_13101,N_12509,N_12648);
nand U13102 (N_13102,N_12897,N_12628);
or U13103 (N_13103,N_12949,N_12892);
xor U13104 (N_13104,N_12953,N_12900);
nand U13105 (N_13105,N_12528,N_12777);
nand U13106 (N_13106,N_12823,N_12818);
nor U13107 (N_13107,N_12625,N_12539);
nor U13108 (N_13108,N_12665,N_12609);
or U13109 (N_13109,N_12784,N_12852);
or U13110 (N_13110,N_12805,N_12688);
or U13111 (N_13111,N_12597,N_12974);
and U13112 (N_13112,N_12515,N_12878);
or U13113 (N_13113,N_12710,N_12736);
or U13114 (N_13114,N_12613,N_12921);
nand U13115 (N_13115,N_12652,N_12735);
and U13116 (N_13116,N_12935,N_12918);
nor U13117 (N_13117,N_12905,N_12902);
nor U13118 (N_13118,N_12529,N_12767);
or U13119 (N_13119,N_12542,N_12985);
nand U13120 (N_13120,N_12827,N_12653);
nor U13121 (N_13121,N_12556,N_12847);
nor U13122 (N_13122,N_12706,N_12851);
or U13123 (N_13123,N_12901,N_12920);
or U13124 (N_13124,N_12863,N_12898);
and U13125 (N_13125,N_12807,N_12712);
xnor U13126 (N_13126,N_12734,N_12775);
or U13127 (N_13127,N_12614,N_12988);
nand U13128 (N_13128,N_12659,N_12561);
nand U13129 (N_13129,N_12797,N_12691);
or U13130 (N_13130,N_12880,N_12888);
and U13131 (N_13131,N_12565,N_12850);
and U13132 (N_13132,N_12983,N_12979);
or U13133 (N_13133,N_12627,N_12978);
nand U13134 (N_13134,N_12654,N_12787);
nand U13135 (N_13135,N_12764,N_12870);
or U13136 (N_13136,N_12843,N_12966);
nor U13137 (N_13137,N_12560,N_12745);
nand U13138 (N_13138,N_12749,N_12917);
nand U13139 (N_13139,N_12700,N_12662);
or U13140 (N_13140,N_12733,N_12853);
xor U13141 (N_13141,N_12903,N_12968);
xnor U13142 (N_13142,N_12770,N_12683);
or U13143 (N_13143,N_12792,N_12596);
and U13144 (N_13144,N_12577,N_12660);
nand U13145 (N_13145,N_12809,N_12601);
and U13146 (N_13146,N_12637,N_12623);
or U13147 (N_13147,N_12783,N_12989);
nor U13148 (N_13148,N_12536,N_12803);
or U13149 (N_13149,N_12997,N_12722);
nor U13150 (N_13150,N_12677,N_12641);
nand U13151 (N_13151,N_12877,N_12944);
nand U13152 (N_13152,N_12580,N_12756);
nor U13153 (N_13153,N_12672,N_12971);
or U13154 (N_13154,N_12808,N_12586);
xnor U13155 (N_13155,N_12657,N_12771);
nor U13156 (N_13156,N_12930,N_12709);
nor U13157 (N_13157,N_12840,N_12925);
nor U13158 (N_13158,N_12980,N_12791);
nand U13159 (N_13159,N_12937,N_12951);
nand U13160 (N_13160,N_12763,N_12842);
nand U13161 (N_13161,N_12612,N_12708);
nand U13162 (N_13162,N_12916,N_12862);
or U13163 (N_13163,N_12947,N_12887);
nand U13164 (N_13164,N_12954,N_12615);
nand U13165 (N_13165,N_12632,N_12950);
or U13166 (N_13166,N_12602,N_12562);
and U13167 (N_13167,N_12624,N_12661);
or U13168 (N_13168,N_12939,N_12719);
or U13169 (N_13169,N_12566,N_12858);
nand U13170 (N_13170,N_12592,N_12765);
nand U13171 (N_13171,N_12855,N_12938);
and U13172 (N_13172,N_12788,N_12856);
or U13173 (N_13173,N_12747,N_12802);
nand U13174 (N_13174,N_12884,N_12674);
nand U13175 (N_13175,N_12626,N_12990);
nor U13176 (N_13176,N_12772,N_12521);
and U13177 (N_13177,N_12588,N_12816);
or U13178 (N_13178,N_12960,N_12669);
nor U13179 (N_13179,N_12885,N_12835);
and U13180 (N_13180,N_12741,N_12711);
nor U13181 (N_13181,N_12861,N_12508);
and U13182 (N_13182,N_12506,N_12603);
nand U13183 (N_13183,N_12755,N_12879);
and U13184 (N_13184,N_12964,N_12644);
nor U13185 (N_13185,N_12514,N_12573);
nand U13186 (N_13186,N_12936,N_12604);
nor U13187 (N_13187,N_12616,N_12593);
and U13188 (N_13188,N_12713,N_12779);
and U13189 (N_13189,N_12844,N_12869);
nand U13190 (N_13190,N_12969,N_12759);
nand U13191 (N_13191,N_12651,N_12881);
or U13192 (N_13192,N_12768,N_12945);
nand U13193 (N_13193,N_12622,N_12934);
or U13194 (N_13194,N_12876,N_12696);
and U13195 (N_13195,N_12730,N_12796);
or U13196 (N_13196,N_12687,N_12782);
nor U13197 (N_13197,N_12799,N_12504);
and U13198 (N_13198,N_12574,N_12650);
nor U13199 (N_13199,N_12762,N_12838);
xor U13200 (N_13200,N_12703,N_12725);
nor U13201 (N_13201,N_12785,N_12545);
and U13202 (N_13202,N_12699,N_12537);
nor U13203 (N_13203,N_12702,N_12866);
nand U13204 (N_13204,N_12739,N_12579);
nand U13205 (N_13205,N_12549,N_12948);
nand U13206 (N_13206,N_12664,N_12996);
nand U13207 (N_13207,N_12972,N_12554);
or U13208 (N_13208,N_12961,N_12789);
or U13209 (N_13209,N_12943,N_12836);
and U13210 (N_13210,N_12984,N_12886);
nor U13211 (N_13211,N_12832,N_12640);
nand U13212 (N_13212,N_12716,N_12684);
nand U13213 (N_13213,N_12621,N_12893);
nand U13214 (N_13214,N_12606,N_12645);
or U13215 (N_13215,N_12695,N_12907);
or U13216 (N_13216,N_12583,N_12873);
nor U13217 (N_13217,N_12761,N_12563);
nor U13218 (N_13218,N_12919,N_12965);
and U13219 (N_13219,N_12846,N_12558);
nand U13220 (N_13220,N_12605,N_12822);
nor U13221 (N_13221,N_12617,N_12868);
nand U13222 (N_13222,N_12500,N_12693);
nor U13223 (N_13223,N_12629,N_12958);
and U13224 (N_13224,N_12587,N_12766);
or U13225 (N_13225,N_12815,N_12543);
and U13226 (N_13226,N_12940,N_12839);
or U13227 (N_13227,N_12837,N_12714);
nor U13228 (N_13228,N_12750,N_12946);
and U13229 (N_13229,N_12977,N_12694);
or U13230 (N_13230,N_12607,N_12620);
nand U13231 (N_13231,N_12618,N_12740);
nor U13232 (N_13232,N_12728,N_12639);
nor U13233 (N_13233,N_12929,N_12812);
nand U13234 (N_13234,N_12600,N_12987);
nor U13235 (N_13235,N_12720,N_12689);
and U13236 (N_13236,N_12833,N_12530);
nor U13237 (N_13237,N_12581,N_12826);
nand U13238 (N_13238,N_12790,N_12957);
and U13239 (N_13239,N_12679,N_12707);
nor U13240 (N_13240,N_12914,N_12552);
nor U13241 (N_13241,N_12906,N_12557);
xnor U13242 (N_13242,N_12995,N_12513);
and U13243 (N_13243,N_12828,N_12524);
or U13244 (N_13244,N_12726,N_12670);
nor U13245 (N_13245,N_12555,N_12571);
or U13246 (N_13246,N_12744,N_12864);
or U13247 (N_13247,N_12781,N_12701);
nand U13248 (N_13248,N_12589,N_12516);
nor U13249 (N_13249,N_12570,N_12667);
and U13250 (N_13250,N_12622,N_12731);
nand U13251 (N_13251,N_12606,N_12726);
nand U13252 (N_13252,N_12505,N_12643);
or U13253 (N_13253,N_12547,N_12793);
or U13254 (N_13254,N_12761,N_12550);
and U13255 (N_13255,N_12928,N_12520);
or U13256 (N_13256,N_12685,N_12691);
nand U13257 (N_13257,N_12972,N_12601);
nor U13258 (N_13258,N_12865,N_12668);
nand U13259 (N_13259,N_12826,N_12515);
and U13260 (N_13260,N_12565,N_12684);
nand U13261 (N_13261,N_12955,N_12813);
nor U13262 (N_13262,N_12662,N_12874);
and U13263 (N_13263,N_12972,N_12889);
and U13264 (N_13264,N_12818,N_12751);
nor U13265 (N_13265,N_12889,N_12726);
nand U13266 (N_13266,N_12903,N_12687);
nor U13267 (N_13267,N_12886,N_12834);
nand U13268 (N_13268,N_12541,N_12718);
nor U13269 (N_13269,N_12733,N_12749);
or U13270 (N_13270,N_12868,N_12920);
nand U13271 (N_13271,N_12850,N_12563);
xor U13272 (N_13272,N_12779,N_12743);
nor U13273 (N_13273,N_12599,N_12873);
nor U13274 (N_13274,N_12793,N_12625);
nor U13275 (N_13275,N_12984,N_12934);
or U13276 (N_13276,N_12838,N_12667);
and U13277 (N_13277,N_12552,N_12638);
nand U13278 (N_13278,N_12979,N_12770);
or U13279 (N_13279,N_12730,N_12974);
nand U13280 (N_13280,N_12787,N_12834);
or U13281 (N_13281,N_12979,N_12594);
and U13282 (N_13282,N_12741,N_12583);
nor U13283 (N_13283,N_12961,N_12727);
nand U13284 (N_13284,N_12982,N_12963);
and U13285 (N_13285,N_12550,N_12725);
nand U13286 (N_13286,N_12827,N_12560);
xnor U13287 (N_13287,N_12914,N_12695);
and U13288 (N_13288,N_12918,N_12502);
or U13289 (N_13289,N_12663,N_12714);
and U13290 (N_13290,N_12811,N_12681);
nor U13291 (N_13291,N_12827,N_12789);
nor U13292 (N_13292,N_12720,N_12997);
nand U13293 (N_13293,N_12873,N_12689);
and U13294 (N_13294,N_12973,N_12512);
or U13295 (N_13295,N_12888,N_12948);
nor U13296 (N_13296,N_12540,N_12524);
and U13297 (N_13297,N_12507,N_12607);
nand U13298 (N_13298,N_12699,N_12760);
nand U13299 (N_13299,N_12537,N_12734);
nand U13300 (N_13300,N_12510,N_12759);
and U13301 (N_13301,N_12889,N_12542);
and U13302 (N_13302,N_12976,N_12779);
and U13303 (N_13303,N_12877,N_12922);
nand U13304 (N_13304,N_12814,N_12780);
or U13305 (N_13305,N_12751,N_12517);
nand U13306 (N_13306,N_12742,N_12939);
nor U13307 (N_13307,N_12672,N_12519);
or U13308 (N_13308,N_12940,N_12564);
nand U13309 (N_13309,N_12928,N_12596);
nand U13310 (N_13310,N_12630,N_12878);
or U13311 (N_13311,N_12693,N_12834);
and U13312 (N_13312,N_12694,N_12865);
nand U13313 (N_13313,N_12528,N_12783);
and U13314 (N_13314,N_12736,N_12576);
nand U13315 (N_13315,N_12579,N_12888);
nand U13316 (N_13316,N_12964,N_12782);
nand U13317 (N_13317,N_12862,N_12727);
nand U13318 (N_13318,N_12991,N_12833);
nor U13319 (N_13319,N_12799,N_12852);
nor U13320 (N_13320,N_12747,N_12594);
xor U13321 (N_13321,N_12711,N_12721);
or U13322 (N_13322,N_12971,N_12968);
or U13323 (N_13323,N_12655,N_12622);
or U13324 (N_13324,N_12923,N_12881);
xnor U13325 (N_13325,N_12845,N_12597);
xnor U13326 (N_13326,N_12782,N_12718);
xor U13327 (N_13327,N_12611,N_12833);
or U13328 (N_13328,N_12525,N_12770);
xor U13329 (N_13329,N_12574,N_12684);
nor U13330 (N_13330,N_12741,N_12954);
nand U13331 (N_13331,N_12820,N_12686);
nand U13332 (N_13332,N_12815,N_12572);
nor U13333 (N_13333,N_12892,N_12760);
nor U13334 (N_13334,N_12757,N_12648);
nand U13335 (N_13335,N_12551,N_12982);
or U13336 (N_13336,N_12579,N_12976);
nor U13337 (N_13337,N_12580,N_12895);
nor U13338 (N_13338,N_12609,N_12524);
nand U13339 (N_13339,N_12921,N_12682);
nand U13340 (N_13340,N_12532,N_12854);
nand U13341 (N_13341,N_12734,N_12749);
xor U13342 (N_13342,N_12643,N_12915);
nor U13343 (N_13343,N_12811,N_12542);
nor U13344 (N_13344,N_12811,N_12978);
and U13345 (N_13345,N_12908,N_12848);
nand U13346 (N_13346,N_12854,N_12642);
and U13347 (N_13347,N_12873,N_12526);
nor U13348 (N_13348,N_12710,N_12894);
nand U13349 (N_13349,N_12684,N_12699);
nand U13350 (N_13350,N_12835,N_12773);
nand U13351 (N_13351,N_12840,N_12856);
or U13352 (N_13352,N_12588,N_12607);
nor U13353 (N_13353,N_12877,N_12751);
or U13354 (N_13354,N_12811,N_12868);
nand U13355 (N_13355,N_12829,N_12955);
xnor U13356 (N_13356,N_12802,N_12798);
and U13357 (N_13357,N_12791,N_12671);
nor U13358 (N_13358,N_12829,N_12809);
and U13359 (N_13359,N_12544,N_12621);
or U13360 (N_13360,N_12538,N_12578);
nand U13361 (N_13361,N_12572,N_12915);
nor U13362 (N_13362,N_12796,N_12771);
and U13363 (N_13363,N_12748,N_12553);
or U13364 (N_13364,N_12614,N_12567);
and U13365 (N_13365,N_12842,N_12635);
xor U13366 (N_13366,N_12998,N_12865);
and U13367 (N_13367,N_12606,N_12671);
and U13368 (N_13368,N_12970,N_12692);
or U13369 (N_13369,N_12973,N_12912);
nor U13370 (N_13370,N_12827,N_12700);
and U13371 (N_13371,N_12832,N_12562);
xor U13372 (N_13372,N_12565,N_12552);
nand U13373 (N_13373,N_12979,N_12518);
and U13374 (N_13374,N_12635,N_12860);
or U13375 (N_13375,N_12721,N_12598);
or U13376 (N_13376,N_12631,N_12648);
nand U13377 (N_13377,N_12542,N_12732);
xnor U13378 (N_13378,N_12692,N_12567);
or U13379 (N_13379,N_12888,N_12692);
or U13380 (N_13380,N_12549,N_12557);
nor U13381 (N_13381,N_12537,N_12635);
nand U13382 (N_13382,N_12772,N_12659);
nor U13383 (N_13383,N_12539,N_12872);
nor U13384 (N_13384,N_12831,N_12778);
and U13385 (N_13385,N_12934,N_12911);
nand U13386 (N_13386,N_12519,N_12793);
and U13387 (N_13387,N_12979,N_12902);
nor U13388 (N_13388,N_12930,N_12999);
or U13389 (N_13389,N_12984,N_12503);
nand U13390 (N_13390,N_12513,N_12806);
or U13391 (N_13391,N_12659,N_12924);
nand U13392 (N_13392,N_12759,N_12546);
or U13393 (N_13393,N_12513,N_12575);
xnor U13394 (N_13394,N_12529,N_12922);
or U13395 (N_13395,N_12716,N_12558);
nand U13396 (N_13396,N_12535,N_12692);
or U13397 (N_13397,N_12875,N_12662);
or U13398 (N_13398,N_12998,N_12632);
nor U13399 (N_13399,N_12941,N_12776);
xnor U13400 (N_13400,N_12778,N_12966);
nor U13401 (N_13401,N_12919,N_12933);
and U13402 (N_13402,N_12538,N_12635);
nor U13403 (N_13403,N_12758,N_12686);
and U13404 (N_13404,N_12829,N_12543);
and U13405 (N_13405,N_12709,N_12741);
and U13406 (N_13406,N_12818,N_12758);
xnor U13407 (N_13407,N_12646,N_12793);
nand U13408 (N_13408,N_12690,N_12620);
nor U13409 (N_13409,N_12750,N_12660);
and U13410 (N_13410,N_12543,N_12621);
xor U13411 (N_13411,N_12886,N_12888);
nand U13412 (N_13412,N_12996,N_12849);
xor U13413 (N_13413,N_12615,N_12958);
and U13414 (N_13414,N_12503,N_12807);
and U13415 (N_13415,N_12763,N_12594);
nor U13416 (N_13416,N_12899,N_12546);
nand U13417 (N_13417,N_12605,N_12599);
nand U13418 (N_13418,N_12979,N_12774);
nand U13419 (N_13419,N_12623,N_12966);
nor U13420 (N_13420,N_12515,N_12959);
nor U13421 (N_13421,N_12769,N_12837);
nand U13422 (N_13422,N_12791,N_12632);
nand U13423 (N_13423,N_12809,N_12665);
nand U13424 (N_13424,N_12566,N_12740);
and U13425 (N_13425,N_12885,N_12587);
nand U13426 (N_13426,N_12545,N_12720);
and U13427 (N_13427,N_12769,N_12915);
and U13428 (N_13428,N_12574,N_12897);
xor U13429 (N_13429,N_12957,N_12958);
or U13430 (N_13430,N_12639,N_12750);
and U13431 (N_13431,N_12924,N_12682);
xnor U13432 (N_13432,N_12865,N_12959);
xnor U13433 (N_13433,N_12846,N_12512);
nand U13434 (N_13434,N_12525,N_12863);
nor U13435 (N_13435,N_12652,N_12602);
nor U13436 (N_13436,N_12606,N_12559);
xor U13437 (N_13437,N_12537,N_12886);
and U13438 (N_13438,N_12563,N_12862);
or U13439 (N_13439,N_12826,N_12967);
nand U13440 (N_13440,N_12946,N_12752);
and U13441 (N_13441,N_12717,N_12543);
and U13442 (N_13442,N_12757,N_12886);
or U13443 (N_13443,N_12624,N_12649);
or U13444 (N_13444,N_12703,N_12879);
xnor U13445 (N_13445,N_12619,N_12554);
and U13446 (N_13446,N_12560,N_12599);
or U13447 (N_13447,N_12849,N_12967);
nand U13448 (N_13448,N_12612,N_12714);
nand U13449 (N_13449,N_12949,N_12843);
nand U13450 (N_13450,N_12846,N_12676);
or U13451 (N_13451,N_12688,N_12785);
nor U13452 (N_13452,N_12906,N_12667);
xor U13453 (N_13453,N_12530,N_12759);
nand U13454 (N_13454,N_12635,N_12680);
nand U13455 (N_13455,N_12634,N_12629);
xnor U13456 (N_13456,N_12852,N_12828);
nor U13457 (N_13457,N_12847,N_12837);
nor U13458 (N_13458,N_12757,N_12735);
and U13459 (N_13459,N_12832,N_12946);
and U13460 (N_13460,N_12689,N_12622);
nand U13461 (N_13461,N_12828,N_12692);
nand U13462 (N_13462,N_12636,N_12500);
or U13463 (N_13463,N_12814,N_12861);
or U13464 (N_13464,N_12885,N_12807);
or U13465 (N_13465,N_12922,N_12740);
nand U13466 (N_13466,N_12654,N_12645);
and U13467 (N_13467,N_12510,N_12619);
nor U13468 (N_13468,N_12904,N_12853);
or U13469 (N_13469,N_12551,N_12744);
nand U13470 (N_13470,N_12542,N_12937);
nor U13471 (N_13471,N_12701,N_12727);
nor U13472 (N_13472,N_12659,N_12620);
nand U13473 (N_13473,N_12662,N_12944);
nand U13474 (N_13474,N_12980,N_12769);
nor U13475 (N_13475,N_12540,N_12514);
or U13476 (N_13476,N_12891,N_12889);
xnor U13477 (N_13477,N_12958,N_12655);
xor U13478 (N_13478,N_12890,N_12830);
or U13479 (N_13479,N_12594,N_12902);
or U13480 (N_13480,N_12530,N_12683);
nor U13481 (N_13481,N_12800,N_12522);
and U13482 (N_13482,N_12680,N_12699);
or U13483 (N_13483,N_12944,N_12633);
nand U13484 (N_13484,N_12953,N_12909);
or U13485 (N_13485,N_12625,N_12611);
and U13486 (N_13486,N_12655,N_12704);
nor U13487 (N_13487,N_12640,N_12813);
and U13488 (N_13488,N_12801,N_12700);
or U13489 (N_13489,N_12874,N_12635);
nand U13490 (N_13490,N_12792,N_12608);
or U13491 (N_13491,N_12968,N_12898);
nand U13492 (N_13492,N_12580,N_12635);
nand U13493 (N_13493,N_12649,N_12788);
nor U13494 (N_13494,N_12923,N_12988);
and U13495 (N_13495,N_12906,N_12785);
or U13496 (N_13496,N_12878,N_12969);
xnor U13497 (N_13497,N_12935,N_12826);
or U13498 (N_13498,N_12539,N_12891);
or U13499 (N_13499,N_12537,N_12696);
xor U13500 (N_13500,N_13243,N_13147);
and U13501 (N_13501,N_13401,N_13082);
xnor U13502 (N_13502,N_13431,N_13377);
and U13503 (N_13503,N_13167,N_13027);
nand U13504 (N_13504,N_13149,N_13326);
or U13505 (N_13505,N_13289,N_13451);
or U13506 (N_13506,N_13456,N_13179);
and U13507 (N_13507,N_13331,N_13443);
xnor U13508 (N_13508,N_13211,N_13154);
and U13509 (N_13509,N_13253,N_13303);
nand U13510 (N_13510,N_13004,N_13412);
and U13511 (N_13511,N_13187,N_13453);
xnor U13512 (N_13512,N_13051,N_13463);
and U13513 (N_13513,N_13310,N_13271);
and U13514 (N_13514,N_13348,N_13146);
and U13515 (N_13515,N_13089,N_13287);
or U13516 (N_13516,N_13069,N_13184);
nand U13517 (N_13517,N_13041,N_13044);
and U13518 (N_13518,N_13399,N_13371);
xor U13519 (N_13519,N_13432,N_13240);
or U13520 (N_13520,N_13319,N_13010);
or U13521 (N_13521,N_13021,N_13367);
nand U13522 (N_13522,N_13102,N_13402);
nand U13523 (N_13523,N_13378,N_13059);
nand U13524 (N_13524,N_13439,N_13291);
nor U13525 (N_13525,N_13449,N_13053);
nand U13526 (N_13526,N_13328,N_13267);
nor U13527 (N_13527,N_13118,N_13200);
nand U13528 (N_13528,N_13216,N_13174);
or U13529 (N_13529,N_13307,N_13337);
and U13530 (N_13530,N_13375,N_13352);
nand U13531 (N_13531,N_13300,N_13330);
nor U13532 (N_13532,N_13237,N_13086);
nor U13533 (N_13533,N_13441,N_13345);
nand U13534 (N_13534,N_13230,N_13272);
nand U13535 (N_13535,N_13383,N_13093);
xor U13536 (N_13536,N_13130,N_13101);
xnor U13537 (N_13537,N_13252,N_13424);
nor U13538 (N_13538,N_13366,N_13075);
or U13539 (N_13539,N_13478,N_13336);
nand U13540 (N_13540,N_13032,N_13056);
nand U13541 (N_13541,N_13162,N_13242);
and U13542 (N_13542,N_13031,N_13262);
and U13543 (N_13543,N_13062,N_13335);
xor U13544 (N_13544,N_13141,N_13065);
xor U13545 (N_13545,N_13195,N_13264);
nor U13546 (N_13546,N_13374,N_13046);
nor U13547 (N_13547,N_13293,N_13350);
xor U13548 (N_13548,N_13224,N_13384);
xnor U13549 (N_13549,N_13256,N_13040);
nor U13550 (N_13550,N_13329,N_13396);
xor U13551 (N_13551,N_13415,N_13100);
or U13552 (N_13552,N_13320,N_13098);
nor U13553 (N_13553,N_13039,N_13270);
nand U13554 (N_13554,N_13492,N_13340);
nor U13555 (N_13555,N_13493,N_13090);
nand U13556 (N_13556,N_13182,N_13382);
nand U13557 (N_13557,N_13254,N_13321);
and U13558 (N_13558,N_13160,N_13372);
or U13559 (N_13559,N_13338,N_13025);
and U13560 (N_13560,N_13007,N_13115);
nand U13561 (N_13561,N_13043,N_13426);
xor U13562 (N_13562,N_13128,N_13111);
nor U13563 (N_13563,N_13464,N_13088);
nor U13564 (N_13564,N_13324,N_13048);
or U13565 (N_13565,N_13356,N_13298);
and U13566 (N_13566,N_13061,N_13484);
nand U13567 (N_13567,N_13151,N_13116);
nor U13568 (N_13568,N_13099,N_13176);
or U13569 (N_13569,N_13064,N_13312);
and U13570 (N_13570,N_13076,N_13009);
nor U13571 (N_13571,N_13285,N_13346);
nand U13572 (N_13572,N_13411,N_13221);
nor U13573 (N_13573,N_13029,N_13016);
or U13574 (N_13574,N_13406,N_13097);
nand U13575 (N_13575,N_13306,N_13360);
nor U13576 (N_13576,N_13067,N_13436);
nand U13577 (N_13577,N_13333,N_13123);
or U13578 (N_13578,N_13214,N_13074);
or U13579 (N_13579,N_13060,N_13207);
or U13580 (N_13580,N_13481,N_13250);
xnor U13581 (N_13581,N_13072,N_13117);
nor U13582 (N_13582,N_13448,N_13175);
nor U13583 (N_13583,N_13398,N_13156);
or U13584 (N_13584,N_13132,N_13361);
xnor U13585 (N_13585,N_13071,N_13313);
nor U13586 (N_13586,N_13459,N_13477);
or U13587 (N_13587,N_13173,N_13433);
or U13588 (N_13588,N_13359,N_13213);
xnor U13589 (N_13589,N_13311,N_13024);
nand U13590 (N_13590,N_13479,N_13392);
nand U13591 (N_13591,N_13020,N_13472);
nor U13592 (N_13592,N_13419,N_13137);
and U13593 (N_13593,N_13486,N_13404);
and U13594 (N_13594,N_13084,N_13198);
nor U13595 (N_13595,N_13277,N_13414);
and U13596 (N_13596,N_13332,N_13466);
nand U13597 (N_13597,N_13379,N_13003);
and U13598 (N_13598,N_13259,N_13129);
and U13599 (N_13599,N_13019,N_13000);
nor U13600 (N_13600,N_13114,N_13322);
and U13601 (N_13601,N_13241,N_13085);
or U13602 (N_13602,N_13257,N_13255);
or U13603 (N_13603,N_13225,N_13140);
or U13604 (N_13604,N_13389,N_13273);
nor U13605 (N_13605,N_13236,N_13470);
or U13606 (N_13606,N_13410,N_13015);
and U13607 (N_13607,N_13217,N_13239);
nand U13608 (N_13608,N_13437,N_13425);
xor U13609 (N_13609,N_13229,N_13125);
or U13610 (N_13610,N_13301,N_13315);
nand U13611 (N_13611,N_13013,N_13138);
nor U13612 (N_13612,N_13033,N_13022);
nor U13613 (N_13613,N_13323,N_13394);
nand U13614 (N_13614,N_13421,N_13440);
and U13615 (N_13615,N_13457,N_13077);
xor U13616 (N_13616,N_13204,N_13142);
nand U13617 (N_13617,N_13327,N_13153);
xor U13618 (N_13618,N_13390,N_13483);
or U13619 (N_13619,N_13199,N_13473);
nor U13620 (N_13620,N_13028,N_13316);
nor U13621 (N_13621,N_13357,N_13244);
nor U13622 (N_13622,N_13317,N_13113);
xnor U13623 (N_13623,N_13011,N_13063);
xnor U13624 (N_13624,N_13249,N_13496);
xor U13625 (N_13625,N_13405,N_13026);
nor U13626 (N_13626,N_13388,N_13260);
or U13627 (N_13627,N_13054,N_13092);
nand U13628 (N_13628,N_13058,N_13023);
or U13629 (N_13629,N_13233,N_13124);
or U13630 (N_13630,N_13012,N_13280);
nand U13631 (N_13631,N_13017,N_13139);
or U13632 (N_13632,N_13127,N_13050);
and U13633 (N_13633,N_13418,N_13121);
xnor U13634 (N_13634,N_13276,N_13339);
nor U13635 (N_13635,N_13438,N_13001);
xor U13636 (N_13636,N_13362,N_13347);
nor U13637 (N_13637,N_13133,N_13381);
and U13638 (N_13638,N_13188,N_13261);
nand U13639 (N_13639,N_13209,N_13235);
nor U13640 (N_13640,N_13281,N_13365);
nand U13641 (N_13641,N_13251,N_13169);
or U13642 (N_13642,N_13126,N_13266);
or U13643 (N_13643,N_13091,N_13245);
or U13644 (N_13644,N_13037,N_13223);
or U13645 (N_13645,N_13487,N_13413);
nand U13646 (N_13646,N_13210,N_13228);
nor U13647 (N_13647,N_13192,N_13103);
nor U13648 (N_13648,N_13158,N_13447);
or U13649 (N_13649,N_13035,N_13191);
or U13650 (N_13650,N_13081,N_13181);
and U13651 (N_13651,N_13208,N_13434);
and U13652 (N_13652,N_13171,N_13430);
nand U13653 (N_13653,N_13417,N_13161);
and U13654 (N_13654,N_13386,N_13079);
or U13655 (N_13655,N_13480,N_13070);
nor U13656 (N_13656,N_13110,N_13247);
and U13657 (N_13657,N_13446,N_13458);
or U13658 (N_13658,N_13164,N_13109);
nor U13659 (N_13659,N_13096,N_13222);
or U13660 (N_13660,N_13364,N_13073);
and U13661 (N_13661,N_13269,N_13445);
nand U13662 (N_13662,N_13283,N_13219);
or U13663 (N_13663,N_13393,N_13442);
or U13664 (N_13664,N_13150,N_13258);
or U13665 (N_13665,N_13450,N_13148);
or U13666 (N_13666,N_13490,N_13353);
nor U13667 (N_13667,N_13295,N_13220);
and U13668 (N_13668,N_13452,N_13166);
nor U13669 (N_13669,N_13226,N_13408);
and U13670 (N_13670,N_13194,N_13052);
nor U13671 (N_13671,N_13363,N_13296);
or U13672 (N_13672,N_13047,N_13455);
xor U13673 (N_13673,N_13178,N_13429);
xor U13674 (N_13674,N_13427,N_13170);
nor U13675 (N_13675,N_13095,N_13469);
nor U13676 (N_13676,N_13334,N_13068);
and U13677 (N_13677,N_13038,N_13215);
and U13678 (N_13678,N_13314,N_13203);
or U13679 (N_13679,N_13395,N_13190);
or U13680 (N_13680,N_13005,N_13387);
nor U13681 (N_13681,N_13403,N_13197);
and U13682 (N_13682,N_13288,N_13152);
nand U13683 (N_13683,N_13369,N_13349);
nand U13684 (N_13684,N_13489,N_13342);
and U13685 (N_13685,N_13227,N_13177);
nand U13686 (N_13686,N_13196,N_13474);
and U13687 (N_13687,N_13159,N_13428);
and U13688 (N_13688,N_13143,N_13248);
nor U13689 (N_13689,N_13325,N_13358);
nor U13690 (N_13690,N_13423,N_13368);
or U13691 (N_13691,N_13465,N_13120);
or U13692 (N_13692,N_13488,N_13036);
or U13693 (N_13693,N_13119,N_13265);
nor U13694 (N_13694,N_13355,N_13193);
nor U13695 (N_13695,N_13416,N_13202);
nor U13696 (N_13696,N_13494,N_13461);
nor U13697 (N_13697,N_13263,N_13475);
and U13698 (N_13698,N_13292,N_13165);
xnor U13699 (N_13699,N_13183,N_13168);
nor U13700 (N_13700,N_13107,N_13305);
nor U13701 (N_13701,N_13163,N_13108);
and U13702 (N_13702,N_13180,N_13370);
nor U13703 (N_13703,N_13122,N_13485);
nor U13704 (N_13704,N_13131,N_13498);
or U13705 (N_13705,N_13476,N_13189);
and U13706 (N_13706,N_13422,N_13135);
or U13707 (N_13707,N_13309,N_13246);
nor U13708 (N_13708,N_13232,N_13391);
xor U13709 (N_13709,N_13268,N_13407);
or U13710 (N_13710,N_13157,N_13030);
xor U13711 (N_13711,N_13454,N_13284);
nor U13712 (N_13712,N_13397,N_13482);
nor U13713 (N_13713,N_13302,N_13499);
or U13714 (N_13714,N_13275,N_13144);
xnor U13715 (N_13715,N_13094,N_13106);
and U13716 (N_13716,N_13294,N_13400);
nand U13717 (N_13717,N_13008,N_13462);
and U13718 (N_13718,N_13468,N_13136);
and U13719 (N_13719,N_13460,N_13491);
or U13720 (N_13720,N_13155,N_13078);
or U13721 (N_13721,N_13341,N_13467);
xnor U13722 (N_13722,N_13083,N_13205);
nand U13723 (N_13723,N_13045,N_13497);
nor U13724 (N_13724,N_13105,N_13134);
and U13725 (N_13725,N_13238,N_13014);
nand U13726 (N_13726,N_13278,N_13234);
nor U13727 (N_13727,N_13380,N_13145);
xor U13728 (N_13728,N_13186,N_13104);
nand U13729 (N_13729,N_13354,N_13201);
xnor U13730 (N_13730,N_13351,N_13080);
or U13731 (N_13731,N_13049,N_13231);
and U13732 (N_13732,N_13297,N_13376);
nor U13733 (N_13733,N_13373,N_13282);
nor U13734 (N_13734,N_13344,N_13002);
or U13735 (N_13735,N_13304,N_13172);
nand U13736 (N_13736,N_13471,N_13343);
and U13737 (N_13737,N_13279,N_13435);
nor U13738 (N_13738,N_13055,N_13420);
nor U13739 (N_13739,N_13385,N_13006);
nand U13740 (N_13740,N_13066,N_13034);
or U13741 (N_13741,N_13112,N_13299);
nor U13742 (N_13742,N_13290,N_13212);
nor U13743 (N_13743,N_13409,N_13057);
nand U13744 (N_13744,N_13286,N_13308);
and U13745 (N_13745,N_13444,N_13185);
xor U13746 (N_13746,N_13087,N_13218);
nor U13747 (N_13747,N_13206,N_13042);
nor U13748 (N_13748,N_13274,N_13018);
nand U13749 (N_13749,N_13318,N_13495);
or U13750 (N_13750,N_13120,N_13109);
and U13751 (N_13751,N_13115,N_13014);
nor U13752 (N_13752,N_13049,N_13387);
or U13753 (N_13753,N_13077,N_13493);
nor U13754 (N_13754,N_13169,N_13351);
nand U13755 (N_13755,N_13337,N_13138);
or U13756 (N_13756,N_13339,N_13375);
nor U13757 (N_13757,N_13042,N_13208);
or U13758 (N_13758,N_13021,N_13009);
and U13759 (N_13759,N_13137,N_13341);
nand U13760 (N_13760,N_13040,N_13182);
and U13761 (N_13761,N_13486,N_13289);
xnor U13762 (N_13762,N_13101,N_13449);
and U13763 (N_13763,N_13226,N_13420);
nor U13764 (N_13764,N_13280,N_13410);
nand U13765 (N_13765,N_13175,N_13347);
xnor U13766 (N_13766,N_13299,N_13418);
and U13767 (N_13767,N_13266,N_13412);
xor U13768 (N_13768,N_13119,N_13294);
nor U13769 (N_13769,N_13457,N_13449);
xor U13770 (N_13770,N_13071,N_13400);
or U13771 (N_13771,N_13254,N_13304);
or U13772 (N_13772,N_13432,N_13487);
and U13773 (N_13773,N_13334,N_13295);
xnor U13774 (N_13774,N_13175,N_13084);
or U13775 (N_13775,N_13126,N_13140);
and U13776 (N_13776,N_13402,N_13086);
nor U13777 (N_13777,N_13487,N_13265);
and U13778 (N_13778,N_13208,N_13021);
nor U13779 (N_13779,N_13489,N_13208);
nand U13780 (N_13780,N_13170,N_13136);
and U13781 (N_13781,N_13448,N_13332);
nor U13782 (N_13782,N_13039,N_13129);
nand U13783 (N_13783,N_13057,N_13275);
nor U13784 (N_13784,N_13486,N_13244);
or U13785 (N_13785,N_13251,N_13176);
and U13786 (N_13786,N_13009,N_13084);
or U13787 (N_13787,N_13257,N_13177);
and U13788 (N_13788,N_13353,N_13473);
nand U13789 (N_13789,N_13311,N_13414);
nor U13790 (N_13790,N_13179,N_13205);
and U13791 (N_13791,N_13202,N_13291);
nand U13792 (N_13792,N_13474,N_13391);
nand U13793 (N_13793,N_13026,N_13114);
nand U13794 (N_13794,N_13153,N_13052);
and U13795 (N_13795,N_13128,N_13191);
nand U13796 (N_13796,N_13176,N_13470);
nand U13797 (N_13797,N_13056,N_13426);
nand U13798 (N_13798,N_13379,N_13214);
xor U13799 (N_13799,N_13025,N_13008);
nand U13800 (N_13800,N_13450,N_13429);
and U13801 (N_13801,N_13195,N_13424);
or U13802 (N_13802,N_13360,N_13185);
and U13803 (N_13803,N_13124,N_13296);
nand U13804 (N_13804,N_13120,N_13435);
nor U13805 (N_13805,N_13055,N_13052);
and U13806 (N_13806,N_13052,N_13117);
and U13807 (N_13807,N_13418,N_13069);
nand U13808 (N_13808,N_13366,N_13376);
nor U13809 (N_13809,N_13441,N_13073);
nor U13810 (N_13810,N_13080,N_13046);
nor U13811 (N_13811,N_13028,N_13285);
and U13812 (N_13812,N_13207,N_13498);
nand U13813 (N_13813,N_13422,N_13365);
or U13814 (N_13814,N_13228,N_13436);
nor U13815 (N_13815,N_13442,N_13250);
nor U13816 (N_13816,N_13003,N_13273);
or U13817 (N_13817,N_13459,N_13091);
and U13818 (N_13818,N_13412,N_13289);
nor U13819 (N_13819,N_13363,N_13148);
and U13820 (N_13820,N_13200,N_13059);
or U13821 (N_13821,N_13460,N_13439);
nor U13822 (N_13822,N_13310,N_13000);
nor U13823 (N_13823,N_13087,N_13399);
nor U13824 (N_13824,N_13312,N_13175);
and U13825 (N_13825,N_13441,N_13038);
nor U13826 (N_13826,N_13449,N_13470);
or U13827 (N_13827,N_13115,N_13123);
or U13828 (N_13828,N_13279,N_13413);
or U13829 (N_13829,N_13007,N_13017);
and U13830 (N_13830,N_13081,N_13366);
nand U13831 (N_13831,N_13248,N_13465);
nand U13832 (N_13832,N_13396,N_13458);
nor U13833 (N_13833,N_13418,N_13467);
xnor U13834 (N_13834,N_13159,N_13163);
or U13835 (N_13835,N_13146,N_13400);
and U13836 (N_13836,N_13457,N_13104);
nand U13837 (N_13837,N_13076,N_13284);
nand U13838 (N_13838,N_13462,N_13297);
and U13839 (N_13839,N_13119,N_13287);
and U13840 (N_13840,N_13214,N_13498);
and U13841 (N_13841,N_13473,N_13482);
and U13842 (N_13842,N_13348,N_13081);
or U13843 (N_13843,N_13012,N_13333);
nor U13844 (N_13844,N_13136,N_13270);
or U13845 (N_13845,N_13227,N_13241);
and U13846 (N_13846,N_13003,N_13123);
and U13847 (N_13847,N_13379,N_13498);
nand U13848 (N_13848,N_13257,N_13325);
nand U13849 (N_13849,N_13255,N_13196);
nand U13850 (N_13850,N_13096,N_13294);
and U13851 (N_13851,N_13391,N_13083);
xor U13852 (N_13852,N_13299,N_13402);
xor U13853 (N_13853,N_13065,N_13038);
nor U13854 (N_13854,N_13325,N_13287);
nor U13855 (N_13855,N_13200,N_13095);
nand U13856 (N_13856,N_13051,N_13176);
nand U13857 (N_13857,N_13089,N_13056);
xor U13858 (N_13858,N_13191,N_13357);
or U13859 (N_13859,N_13428,N_13493);
nand U13860 (N_13860,N_13012,N_13457);
nand U13861 (N_13861,N_13434,N_13023);
nor U13862 (N_13862,N_13088,N_13106);
nor U13863 (N_13863,N_13077,N_13193);
nand U13864 (N_13864,N_13078,N_13437);
or U13865 (N_13865,N_13168,N_13267);
xnor U13866 (N_13866,N_13484,N_13166);
xor U13867 (N_13867,N_13366,N_13440);
nor U13868 (N_13868,N_13098,N_13095);
and U13869 (N_13869,N_13402,N_13358);
nand U13870 (N_13870,N_13197,N_13360);
nand U13871 (N_13871,N_13036,N_13006);
nor U13872 (N_13872,N_13332,N_13286);
and U13873 (N_13873,N_13044,N_13095);
and U13874 (N_13874,N_13062,N_13224);
nor U13875 (N_13875,N_13015,N_13155);
nand U13876 (N_13876,N_13037,N_13457);
nor U13877 (N_13877,N_13450,N_13019);
nor U13878 (N_13878,N_13019,N_13358);
or U13879 (N_13879,N_13148,N_13219);
nor U13880 (N_13880,N_13119,N_13423);
nor U13881 (N_13881,N_13404,N_13348);
nand U13882 (N_13882,N_13124,N_13039);
or U13883 (N_13883,N_13078,N_13362);
nor U13884 (N_13884,N_13358,N_13063);
and U13885 (N_13885,N_13451,N_13380);
or U13886 (N_13886,N_13379,N_13189);
or U13887 (N_13887,N_13233,N_13200);
nor U13888 (N_13888,N_13490,N_13339);
or U13889 (N_13889,N_13136,N_13025);
nor U13890 (N_13890,N_13026,N_13101);
nor U13891 (N_13891,N_13489,N_13165);
and U13892 (N_13892,N_13126,N_13476);
or U13893 (N_13893,N_13228,N_13163);
and U13894 (N_13894,N_13385,N_13486);
or U13895 (N_13895,N_13122,N_13435);
or U13896 (N_13896,N_13260,N_13221);
nand U13897 (N_13897,N_13351,N_13310);
or U13898 (N_13898,N_13018,N_13233);
or U13899 (N_13899,N_13481,N_13030);
and U13900 (N_13900,N_13159,N_13323);
and U13901 (N_13901,N_13028,N_13360);
nor U13902 (N_13902,N_13062,N_13209);
nand U13903 (N_13903,N_13441,N_13018);
nand U13904 (N_13904,N_13073,N_13109);
nand U13905 (N_13905,N_13192,N_13410);
nor U13906 (N_13906,N_13481,N_13382);
or U13907 (N_13907,N_13288,N_13390);
and U13908 (N_13908,N_13135,N_13265);
xor U13909 (N_13909,N_13258,N_13187);
nand U13910 (N_13910,N_13184,N_13190);
nand U13911 (N_13911,N_13065,N_13210);
xnor U13912 (N_13912,N_13369,N_13352);
or U13913 (N_13913,N_13343,N_13357);
nand U13914 (N_13914,N_13478,N_13439);
or U13915 (N_13915,N_13242,N_13031);
xnor U13916 (N_13916,N_13202,N_13349);
and U13917 (N_13917,N_13100,N_13150);
nand U13918 (N_13918,N_13395,N_13067);
nand U13919 (N_13919,N_13255,N_13306);
and U13920 (N_13920,N_13332,N_13450);
and U13921 (N_13921,N_13219,N_13160);
nor U13922 (N_13922,N_13080,N_13476);
nand U13923 (N_13923,N_13331,N_13391);
and U13924 (N_13924,N_13103,N_13419);
nand U13925 (N_13925,N_13175,N_13418);
nand U13926 (N_13926,N_13131,N_13479);
and U13927 (N_13927,N_13462,N_13377);
and U13928 (N_13928,N_13206,N_13122);
and U13929 (N_13929,N_13027,N_13294);
xor U13930 (N_13930,N_13183,N_13164);
nand U13931 (N_13931,N_13007,N_13366);
nor U13932 (N_13932,N_13128,N_13120);
and U13933 (N_13933,N_13180,N_13214);
and U13934 (N_13934,N_13166,N_13340);
xnor U13935 (N_13935,N_13280,N_13321);
and U13936 (N_13936,N_13094,N_13174);
or U13937 (N_13937,N_13433,N_13189);
xor U13938 (N_13938,N_13332,N_13015);
nand U13939 (N_13939,N_13114,N_13131);
or U13940 (N_13940,N_13255,N_13241);
nand U13941 (N_13941,N_13431,N_13498);
nor U13942 (N_13942,N_13388,N_13496);
and U13943 (N_13943,N_13364,N_13077);
nand U13944 (N_13944,N_13494,N_13198);
and U13945 (N_13945,N_13223,N_13406);
and U13946 (N_13946,N_13290,N_13199);
nor U13947 (N_13947,N_13287,N_13037);
nor U13948 (N_13948,N_13063,N_13236);
or U13949 (N_13949,N_13487,N_13154);
or U13950 (N_13950,N_13190,N_13292);
and U13951 (N_13951,N_13454,N_13401);
nand U13952 (N_13952,N_13017,N_13072);
nand U13953 (N_13953,N_13351,N_13193);
and U13954 (N_13954,N_13040,N_13227);
and U13955 (N_13955,N_13144,N_13128);
nand U13956 (N_13956,N_13332,N_13049);
nand U13957 (N_13957,N_13303,N_13430);
or U13958 (N_13958,N_13288,N_13001);
xnor U13959 (N_13959,N_13039,N_13273);
nor U13960 (N_13960,N_13482,N_13475);
xnor U13961 (N_13961,N_13351,N_13235);
xnor U13962 (N_13962,N_13037,N_13060);
xor U13963 (N_13963,N_13034,N_13247);
or U13964 (N_13964,N_13248,N_13213);
xnor U13965 (N_13965,N_13095,N_13068);
and U13966 (N_13966,N_13350,N_13272);
nor U13967 (N_13967,N_13027,N_13233);
nor U13968 (N_13968,N_13318,N_13211);
and U13969 (N_13969,N_13304,N_13024);
or U13970 (N_13970,N_13311,N_13025);
and U13971 (N_13971,N_13459,N_13414);
or U13972 (N_13972,N_13013,N_13109);
nor U13973 (N_13973,N_13163,N_13304);
or U13974 (N_13974,N_13333,N_13232);
nor U13975 (N_13975,N_13149,N_13052);
nor U13976 (N_13976,N_13152,N_13131);
and U13977 (N_13977,N_13058,N_13243);
or U13978 (N_13978,N_13310,N_13293);
nand U13979 (N_13979,N_13295,N_13177);
nand U13980 (N_13980,N_13405,N_13477);
nand U13981 (N_13981,N_13406,N_13294);
nor U13982 (N_13982,N_13054,N_13490);
nand U13983 (N_13983,N_13145,N_13318);
and U13984 (N_13984,N_13341,N_13005);
and U13985 (N_13985,N_13354,N_13066);
nand U13986 (N_13986,N_13496,N_13192);
xor U13987 (N_13987,N_13000,N_13247);
nor U13988 (N_13988,N_13399,N_13077);
nor U13989 (N_13989,N_13461,N_13000);
nor U13990 (N_13990,N_13340,N_13434);
nand U13991 (N_13991,N_13133,N_13236);
nor U13992 (N_13992,N_13435,N_13495);
nor U13993 (N_13993,N_13383,N_13472);
nor U13994 (N_13994,N_13390,N_13322);
nor U13995 (N_13995,N_13035,N_13238);
nand U13996 (N_13996,N_13208,N_13499);
or U13997 (N_13997,N_13444,N_13450);
nor U13998 (N_13998,N_13389,N_13168);
or U13999 (N_13999,N_13398,N_13391);
or U14000 (N_14000,N_13745,N_13644);
nor U14001 (N_14001,N_13813,N_13865);
and U14002 (N_14002,N_13731,N_13962);
or U14003 (N_14003,N_13526,N_13572);
and U14004 (N_14004,N_13506,N_13741);
nand U14005 (N_14005,N_13970,N_13833);
nor U14006 (N_14006,N_13640,N_13571);
or U14007 (N_14007,N_13671,N_13637);
or U14008 (N_14008,N_13899,N_13854);
and U14009 (N_14009,N_13947,N_13593);
nand U14010 (N_14010,N_13752,N_13573);
and U14011 (N_14011,N_13558,N_13931);
or U14012 (N_14012,N_13955,N_13645);
and U14013 (N_14013,N_13673,N_13901);
nor U14014 (N_14014,N_13807,N_13896);
and U14015 (N_14015,N_13795,N_13714);
nand U14016 (N_14016,N_13706,N_13744);
and U14017 (N_14017,N_13621,N_13948);
and U14018 (N_14018,N_13918,N_13678);
xnor U14019 (N_14019,N_13654,N_13950);
or U14020 (N_14020,N_13909,N_13508);
or U14021 (N_14021,N_13863,N_13528);
nand U14022 (N_14022,N_13702,N_13521);
or U14023 (N_14023,N_13674,N_13589);
or U14024 (N_14024,N_13810,N_13597);
or U14025 (N_14025,N_13823,N_13728);
nor U14026 (N_14026,N_13834,N_13804);
nor U14027 (N_14027,N_13773,N_13539);
or U14028 (N_14028,N_13662,N_13746);
xnor U14029 (N_14029,N_13562,N_13542);
or U14030 (N_14030,N_13544,N_13545);
nor U14031 (N_14031,N_13825,N_13999);
or U14032 (N_14032,N_13519,N_13601);
nor U14033 (N_14033,N_13616,N_13697);
and U14034 (N_14034,N_13818,N_13740);
nand U14035 (N_14035,N_13657,N_13791);
or U14036 (N_14036,N_13839,N_13883);
or U14037 (N_14037,N_13996,N_13806);
and U14038 (N_14038,N_13965,N_13549);
and U14039 (N_14039,N_13705,N_13511);
and U14040 (N_14040,N_13869,N_13800);
nor U14041 (N_14041,N_13566,N_13775);
xor U14042 (N_14042,N_13503,N_13737);
nand U14043 (N_14043,N_13617,N_13720);
or U14044 (N_14044,N_13933,N_13792);
or U14045 (N_14045,N_13514,N_13591);
or U14046 (N_14046,N_13553,N_13525);
nand U14047 (N_14047,N_13864,N_13889);
or U14048 (N_14048,N_13577,N_13590);
and U14049 (N_14049,N_13935,N_13648);
nand U14050 (N_14050,N_13959,N_13556);
or U14051 (N_14051,N_13911,N_13672);
or U14052 (N_14052,N_13780,N_13788);
and U14053 (N_14053,N_13666,N_13533);
nor U14054 (N_14054,N_13599,N_13609);
nand U14055 (N_14055,N_13554,N_13582);
nor U14056 (N_14056,N_13504,N_13801);
or U14057 (N_14057,N_13820,N_13631);
nand U14058 (N_14058,N_13679,N_13595);
nand U14059 (N_14059,N_13915,N_13557);
xnor U14060 (N_14060,N_13634,N_13772);
or U14061 (N_14061,N_13707,N_13624);
and U14062 (N_14062,N_13829,N_13847);
or U14063 (N_14063,N_13567,N_13653);
and U14064 (N_14064,N_13994,N_13793);
nand U14065 (N_14065,N_13698,N_13765);
and U14066 (N_14066,N_13811,N_13874);
and U14067 (N_14067,N_13763,N_13650);
and U14068 (N_14068,N_13887,N_13622);
nand U14069 (N_14069,N_13749,N_13750);
nand U14070 (N_14070,N_13642,N_13560);
nor U14071 (N_14071,N_13734,N_13838);
nand U14072 (N_14072,N_13904,N_13636);
nor U14073 (N_14073,N_13578,N_13592);
and U14074 (N_14074,N_13665,N_13512);
nor U14075 (N_14075,N_13513,N_13778);
nand U14076 (N_14076,N_13532,N_13564);
nor U14077 (N_14077,N_13611,N_13912);
or U14078 (N_14078,N_13670,N_13689);
and U14079 (N_14079,N_13675,N_13574);
and U14080 (N_14080,N_13968,N_13951);
or U14081 (N_14081,N_13952,N_13808);
nor U14082 (N_14082,N_13894,N_13628);
and U14083 (N_14083,N_13934,N_13897);
nor U14084 (N_14084,N_13868,N_13692);
xnor U14085 (N_14085,N_13853,N_13727);
and U14086 (N_14086,N_13860,N_13957);
and U14087 (N_14087,N_13517,N_13880);
and U14088 (N_14088,N_13882,N_13659);
and U14089 (N_14089,N_13987,N_13747);
or U14090 (N_14090,N_13768,N_13633);
or U14091 (N_14091,N_13638,N_13523);
and U14092 (N_14092,N_13779,N_13843);
xor U14093 (N_14093,N_13585,N_13625);
nand U14094 (N_14094,N_13984,N_13607);
and U14095 (N_14095,N_13535,N_13836);
and U14096 (N_14096,N_13527,N_13992);
nor U14097 (N_14097,N_13682,N_13919);
and U14098 (N_14098,N_13726,N_13858);
nor U14099 (N_14099,N_13693,N_13849);
nand U14100 (N_14100,N_13939,N_13531);
nand U14101 (N_14101,N_13937,N_13852);
nand U14102 (N_14102,N_13717,N_13884);
or U14103 (N_14103,N_13976,N_13997);
nor U14104 (N_14104,N_13857,N_13776);
nand U14105 (N_14105,N_13835,N_13738);
nand U14106 (N_14106,N_13837,N_13991);
nor U14107 (N_14107,N_13651,N_13649);
xor U14108 (N_14108,N_13736,N_13784);
nor U14109 (N_14109,N_13958,N_13866);
or U14110 (N_14110,N_13753,N_13584);
nand U14111 (N_14111,N_13700,N_13719);
and U14112 (N_14112,N_13709,N_13695);
and U14113 (N_14113,N_13755,N_13522);
or U14114 (N_14114,N_13614,N_13930);
nand U14115 (N_14115,N_13711,N_13524);
nand U14116 (N_14116,N_13652,N_13623);
nand U14117 (N_14117,N_13660,N_13798);
nor U14118 (N_14118,N_13851,N_13774);
nor U14119 (N_14119,N_13600,N_13701);
and U14120 (N_14120,N_13536,N_13856);
nand U14121 (N_14121,N_13570,N_13579);
nor U14122 (N_14122,N_13677,N_13817);
nand U14123 (N_14123,N_13827,N_13938);
or U14124 (N_14124,N_13979,N_13981);
or U14125 (N_14125,N_13840,N_13803);
nand U14126 (N_14126,N_13832,N_13777);
nand U14127 (N_14127,N_13756,N_13664);
nand U14128 (N_14128,N_13949,N_13696);
nand U14129 (N_14129,N_13786,N_13893);
or U14130 (N_14130,N_13975,N_13739);
and U14131 (N_14131,N_13805,N_13748);
or U14132 (N_14132,N_13956,N_13646);
or U14133 (N_14133,N_13668,N_13501);
or U14134 (N_14134,N_13925,N_13555);
and U14135 (N_14135,N_13635,N_13867);
xnor U14136 (N_14136,N_13973,N_13723);
nor U14137 (N_14137,N_13615,N_13713);
nor U14138 (N_14138,N_13923,N_13961);
and U14139 (N_14139,N_13751,N_13708);
or U14140 (N_14140,N_13797,N_13985);
and U14141 (N_14141,N_13821,N_13977);
or U14142 (N_14142,N_13667,N_13690);
or U14143 (N_14143,N_13656,N_13940);
and U14144 (N_14144,N_13922,N_13790);
nand U14145 (N_14145,N_13841,N_13872);
or U14146 (N_14146,N_13781,N_13946);
or U14147 (N_14147,N_13538,N_13534);
nor U14148 (N_14148,N_13725,N_13855);
or U14149 (N_14149,N_13916,N_13641);
or U14150 (N_14150,N_13594,N_13581);
nor U14151 (N_14151,N_13760,N_13859);
nor U14152 (N_14152,N_13771,N_13966);
xnor U14153 (N_14153,N_13618,N_13926);
xnor U14154 (N_14154,N_13885,N_13878);
nor U14155 (N_14155,N_13518,N_13603);
nand U14156 (N_14156,N_13875,N_13782);
or U14157 (N_14157,N_13619,N_13809);
nor U14158 (N_14158,N_13565,N_13953);
and U14159 (N_14159,N_13643,N_13816);
and U14160 (N_14160,N_13908,N_13764);
nand U14161 (N_14161,N_13906,N_13972);
nand U14162 (N_14162,N_13815,N_13913);
and U14163 (N_14163,N_13569,N_13758);
or U14164 (N_14164,N_13543,N_13986);
nand U14165 (N_14165,N_13547,N_13932);
nor U14166 (N_14166,N_13612,N_13941);
nand U14167 (N_14167,N_13629,N_13954);
xor U14168 (N_14168,N_13561,N_13914);
xnor U14169 (N_14169,N_13710,N_13683);
or U14170 (N_14170,N_13620,N_13552);
nor U14171 (N_14171,N_13826,N_13982);
nor U14172 (N_14172,N_13530,N_13576);
or U14173 (N_14173,N_13694,N_13502);
nand U14174 (N_14174,N_13978,N_13548);
nand U14175 (N_14175,N_13681,N_13529);
nand U14176 (N_14176,N_13783,N_13845);
nor U14177 (N_14177,N_13550,N_13680);
xor U14178 (N_14178,N_13754,N_13730);
nand U14179 (N_14179,N_13828,N_13787);
nand U14180 (N_14180,N_13770,N_13830);
or U14181 (N_14181,N_13890,N_13691);
and U14182 (N_14182,N_13580,N_13732);
nor U14183 (N_14183,N_13546,N_13892);
and U14184 (N_14184,N_13895,N_13989);
nand U14185 (N_14185,N_13520,N_13924);
xor U14186 (N_14186,N_13743,N_13861);
nor U14187 (N_14187,N_13583,N_13742);
and U14188 (N_14188,N_13588,N_13718);
or U14189 (N_14189,N_13928,N_13990);
and U14190 (N_14190,N_13684,N_13850);
nor U14191 (N_14191,N_13888,N_13761);
nand U14192 (N_14192,N_13766,N_13862);
or U14193 (N_14193,N_13563,N_13735);
nand U14194 (N_14194,N_13812,N_13967);
or U14195 (N_14195,N_13964,N_13980);
or U14196 (N_14196,N_13669,N_13510);
or U14197 (N_14197,N_13983,N_13995);
nand U14198 (N_14198,N_13541,N_13802);
and U14199 (N_14199,N_13794,N_13630);
and U14200 (N_14200,N_13604,N_13627);
and U14201 (N_14201,N_13907,N_13685);
nor U14202 (N_14202,N_13876,N_13917);
xor U14203 (N_14203,N_13936,N_13814);
nand U14204 (N_14204,N_13505,N_13785);
nand U14205 (N_14205,N_13688,N_13699);
or U14206 (N_14206,N_13842,N_13613);
nor U14207 (N_14207,N_13799,N_13757);
nand U14208 (N_14208,N_13819,N_13846);
nand U14209 (N_14209,N_13626,N_13902);
and U14210 (N_14210,N_13960,N_13871);
nor U14211 (N_14211,N_13993,N_13929);
or U14212 (N_14212,N_13515,N_13759);
nand U14213 (N_14213,N_13715,N_13729);
nor U14214 (N_14214,N_13903,N_13598);
nand U14215 (N_14215,N_13639,N_13963);
xnor U14216 (N_14216,N_13831,N_13998);
xor U14217 (N_14217,N_13873,N_13703);
nor U14218 (N_14218,N_13724,N_13942);
nor U14219 (N_14219,N_13722,N_13551);
and U14220 (N_14220,N_13655,N_13769);
or U14221 (N_14221,N_13969,N_13898);
xor U14222 (N_14222,N_13661,N_13848);
or U14223 (N_14223,N_13721,N_13927);
or U14224 (N_14224,N_13762,N_13687);
nor U14225 (N_14225,N_13824,N_13988);
nand U14226 (N_14226,N_13537,N_13796);
nand U14227 (N_14227,N_13974,N_13879);
xnor U14228 (N_14228,N_13605,N_13704);
xnor U14229 (N_14229,N_13945,N_13910);
or U14230 (N_14230,N_13712,N_13608);
nand U14231 (N_14231,N_13575,N_13943);
nor U14232 (N_14232,N_13971,N_13658);
nand U14233 (N_14233,N_13559,N_13881);
nor U14234 (N_14234,N_13568,N_13606);
nor U14235 (N_14235,N_13586,N_13767);
nand U14236 (N_14236,N_13905,N_13540);
and U14237 (N_14237,N_13921,N_13647);
or U14238 (N_14238,N_13716,N_13877);
nor U14239 (N_14239,N_13944,N_13587);
and U14240 (N_14240,N_13596,N_13509);
and U14241 (N_14241,N_13610,N_13920);
or U14242 (N_14242,N_13891,N_13663);
or U14243 (N_14243,N_13676,N_13789);
and U14244 (N_14244,N_13870,N_13822);
nor U14245 (N_14245,N_13507,N_13844);
and U14246 (N_14246,N_13886,N_13900);
and U14247 (N_14247,N_13632,N_13686);
xnor U14248 (N_14248,N_13516,N_13733);
nand U14249 (N_14249,N_13500,N_13602);
nor U14250 (N_14250,N_13538,N_13610);
nor U14251 (N_14251,N_13771,N_13538);
and U14252 (N_14252,N_13518,N_13781);
and U14253 (N_14253,N_13559,N_13572);
nor U14254 (N_14254,N_13972,N_13707);
or U14255 (N_14255,N_13669,N_13880);
and U14256 (N_14256,N_13847,N_13560);
nor U14257 (N_14257,N_13807,N_13907);
or U14258 (N_14258,N_13722,N_13965);
nor U14259 (N_14259,N_13805,N_13865);
and U14260 (N_14260,N_13982,N_13568);
xnor U14261 (N_14261,N_13836,N_13800);
nor U14262 (N_14262,N_13750,N_13597);
nor U14263 (N_14263,N_13757,N_13952);
or U14264 (N_14264,N_13880,N_13514);
and U14265 (N_14265,N_13532,N_13573);
nand U14266 (N_14266,N_13715,N_13859);
and U14267 (N_14267,N_13759,N_13696);
and U14268 (N_14268,N_13982,N_13994);
xnor U14269 (N_14269,N_13798,N_13951);
or U14270 (N_14270,N_13782,N_13611);
or U14271 (N_14271,N_13747,N_13646);
nor U14272 (N_14272,N_13649,N_13993);
xnor U14273 (N_14273,N_13745,N_13501);
nor U14274 (N_14274,N_13854,N_13919);
nor U14275 (N_14275,N_13651,N_13901);
nand U14276 (N_14276,N_13732,N_13981);
and U14277 (N_14277,N_13696,N_13833);
nand U14278 (N_14278,N_13600,N_13995);
nor U14279 (N_14279,N_13989,N_13920);
or U14280 (N_14280,N_13620,N_13881);
or U14281 (N_14281,N_13972,N_13662);
nor U14282 (N_14282,N_13646,N_13784);
or U14283 (N_14283,N_13620,N_13611);
nand U14284 (N_14284,N_13865,N_13915);
xnor U14285 (N_14285,N_13607,N_13801);
or U14286 (N_14286,N_13884,N_13501);
xor U14287 (N_14287,N_13768,N_13790);
nand U14288 (N_14288,N_13862,N_13961);
nand U14289 (N_14289,N_13994,N_13915);
and U14290 (N_14290,N_13544,N_13823);
nand U14291 (N_14291,N_13712,N_13763);
and U14292 (N_14292,N_13811,N_13882);
and U14293 (N_14293,N_13629,N_13845);
or U14294 (N_14294,N_13685,N_13672);
nor U14295 (N_14295,N_13768,N_13678);
or U14296 (N_14296,N_13956,N_13836);
nand U14297 (N_14297,N_13546,N_13564);
and U14298 (N_14298,N_13582,N_13650);
nand U14299 (N_14299,N_13905,N_13710);
and U14300 (N_14300,N_13516,N_13935);
nor U14301 (N_14301,N_13840,N_13986);
nand U14302 (N_14302,N_13779,N_13607);
nand U14303 (N_14303,N_13902,N_13583);
and U14304 (N_14304,N_13598,N_13514);
nor U14305 (N_14305,N_13884,N_13571);
or U14306 (N_14306,N_13946,N_13822);
nor U14307 (N_14307,N_13541,N_13707);
or U14308 (N_14308,N_13613,N_13632);
and U14309 (N_14309,N_13609,N_13734);
xor U14310 (N_14310,N_13523,N_13503);
and U14311 (N_14311,N_13624,N_13574);
nor U14312 (N_14312,N_13524,N_13761);
nor U14313 (N_14313,N_13942,N_13997);
nand U14314 (N_14314,N_13511,N_13616);
or U14315 (N_14315,N_13881,N_13712);
nand U14316 (N_14316,N_13653,N_13972);
or U14317 (N_14317,N_13961,N_13632);
nor U14318 (N_14318,N_13782,N_13625);
xor U14319 (N_14319,N_13896,N_13918);
nor U14320 (N_14320,N_13570,N_13952);
nor U14321 (N_14321,N_13549,N_13695);
or U14322 (N_14322,N_13702,N_13580);
and U14323 (N_14323,N_13863,N_13501);
and U14324 (N_14324,N_13835,N_13806);
or U14325 (N_14325,N_13672,N_13924);
or U14326 (N_14326,N_13631,N_13835);
nand U14327 (N_14327,N_13508,N_13828);
nand U14328 (N_14328,N_13864,N_13866);
nor U14329 (N_14329,N_13613,N_13861);
and U14330 (N_14330,N_13826,N_13959);
nor U14331 (N_14331,N_13599,N_13955);
nand U14332 (N_14332,N_13883,N_13610);
xor U14333 (N_14333,N_13553,N_13829);
nand U14334 (N_14334,N_13679,N_13575);
nor U14335 (N_14335,N_13983,N_13904);
nand U14336 (N_14336,N_13899,N_13928);
and U14337 (N_14337,N_13554,N_13729);
or U14338 (N_14338,N_13570,N_13723);
nand U14339 (N_14339,N_13895,N_13574);
and U14340 (N_14340,N_13658,N_13788);
nor U14341 (N_14341,N_13950,N_13758);
nand U14342 (N_14342,N_13697,N_13726);
and U14343 (N_14343,N_13807,N_13581);
or U14344 (N_14344,N_13686,N_13918);
nor U14345 (N_14345,N_13909,N_13712);
nand U14346 (N_14346,N_13603,N_13851);
nor U14347 (N_14347,N_13618,N_13843);
nor U14348 (N_14348,N_13860,N_13909);
nand U14349 (N_14349,N_13790,N_13770);
or U14350 (N_14350,N_13696,N_13544);
nor U14351 (N_14351,N_13919,N_13933);
and U14352 (N_14352,N_13601,N_13683);
nor U14353 (N_14353,N_13565,N_13937);
nor U14354 (N_14354,N_13978,N_13794);
or U14355 (N_14355,N_13682,N_13718);
nand U14356 (N_14356,N_13956,N_13527);
and U14357 (N_14357,N_13708,N_13518);
or U14358 (N_14358,N_13527,N_13577);
nand U14359 (N_14359,N_13752,N_13674);
nand U14360 (N_14360,N_13882,N_13694);
or U14361 (N_14361,N_13973,N_13685);
and U14362 (N_14362,N_13801,N_13542);
nor U14363 (N_14363,N_13943,N_13786);
nor U14364 (N_14364,N_13977,N_13813);
nor U14365 (N_14365,N_13864,N_13930);
and U14366 (N_14366,N_13515,N_13969);
nand U14367 (N_14367,N_13616,N_13623);
nand U14368 (N_14368,N_13519,N_13889);
or U14369 (N_14369,N_13544,N_13748);
or U14370 (N_14370,N_13668,N_13714);
nor U14371 (N_14371,N_13923,N_13558);
and U14372 (N_14372,N_13567,N_13532);
xor U14373 (N_14373,N_13856,N_13773);
nor U14374 (N_14374,N_13832,N_13511);
or U14375 (N_14375,N_13592,N_13948);
nor U14376 (N_14376,N_13552,N_13884);
nor U14377 (N_14377,N_13846,N_13676);
or U14378 (N_14378,N_13708,N_13913);
nand U14379 (N_14379,N_13717,N_13743);
nand U14380 (N_14380,N_13948,N_13958);
xor U14381 (N_14381,N_13872,N_13689);
or U14382 (N_14382,N_13503,N_13992);
and U14383 (N_14383,N_13905,N_13774);
xnor U14384 (N_14384,N_13584,N_13655);
nand U14385 (N_14385,N_13736,N_13604);
and U14386 (N_14386,N_13924,N_13602);
nand U14387 (N_14387,N_13700,N_13622);
xnor U14388 (N_14388,N_13550,N_13507);
nand U14389 (N_14389,N_13591,N_13950);
nor U14390 (N_14390,N_13812,N_13832);
or U14391 (N_14391,N_13850,N_13954);
or U14392 (N_14392,N_13820,N_13535);
xnor U14393 (N_14393,N_13956,N_13686);
nor U14394 (N_14394,N_13592,N_13989);
and U14395 (N_14395,N_13554,N_13976);
or U14396 (N_14396,N_13797,N_13856);
nor U14397 (N_14397,N_13773,N_13723);
or U14398 (N_14398,N_13834,N_13632);
nand U14399 (N_14399,N_13733,N_13578);
and U14400 (N_14400,N_13784,N_13515);
nand U14401 (N_14401,N_13559,N_13719);
and U14402 (N_14402,N_13718,N_13698);
nand U14403 (N_14403,N_13873,N_13754);
and U14404 (N_14404,N_13945,N_13522);
or U14405 (N_14405,N_13748,N_13964);
or U14406 (N_14406,N_13901,N_13518);
nand U14407 (N_14407,N_13678,N_13722);
or U14408 (N_14408,N_13944,N_13887);
nand U14409 (N_14409,N_13851,N_13529);
nand U14410 (N_14410,N_13680,N_13585);
nand U14411 (N_14411,N_13661,N_13651);
nor U14412 (N_14412,N_13928,N_13749);
nor U14413 (N_14413,N_13568,N_13798);
and U14414 (N_14414,N_13625,N_13833);
nand U14415 (N_14415,N_13733,N_13555);
or U14416 (N_14416,N_13699,N_13966);
nor U14417 (N_14417,N_13796,N_13504);
and U14418 (N_14418,N_13667,N_13737);
and U14419 (N_14419,N_13904,N_13563);
and U14420 (N_14420,N_13854,N_13737);
nand U14421 (N_14421,N_13699,N_13956);
or U14422 (N_14422,N_13569,N_13521);
and U14423 (N_14423,N_13642,N_13677);
xor U14424 (N_14424,N_13680,N_13985);
and U14425 (N_14425,N_13865,N_13919);
and U14426 (N_14426,N_13744,N_13695);
nor U14427 (N_14427,N_13596,N_13579);
and U14428 (N_14428,N_13811,N_13914);
and U14429 (N_14429,N_13534,N_13710);
or U14430 (N_14430,N_13562,N_13540);
or U14431 (N_14431,N_13655,N_13856);
nor U14432 (N_14432,N_13849,N_13657);
or U14433 (N_14433,N_13860,N_13696);
or U14434 (N_14434,N_13928,N_13588);
nand U14435 (N_14435,N_13652,N_13602);
and U14436 (N_14436,N_13795,N_13617);
nand U14437 (N_14437,N_13608,N_13523);
nand U14438 (N_14438,N_13812,N_13639);
xor U14439 (N_14439,N_13910,N_13724);
or U14440 (N_14440,N_13841,N_13816);
nand U14441 (N_14441,N_13644,N_13621);
and U14442 (N_14442,N_13969,N_13743);
nor U14443 (N_14443,N_13778,N_13544);
xor U14444 (N_14444,N_13753,N_13931);
nand U14445 (N_14445,N_13675,N_13681);
or U14446 (N_14446,N_13856,N_13535);
and U14447 (N_14447,N_13758,N_13667);
nand U14448 (N_14448,N_13953,N_13922);
or U14449 (N_14449,N_13703,N_13893);
nor U14450 (N_14450,N_13829,N_13651);
nand U14451 (N_14451,N_13875,N_13665);
nand U14452 (N_14452,N_13675,N_13746);
nand U14453 (N_14453,N_13863,N_13986);
or U14454 (N_14454,N_13697,N_13557);
nor U14455 (N_14455,N_13690,N_13567);
or U14456 (N_14456,N_13634,N_13958);
nand U14457 (N_14457,N_13932,N_13769);
nor U14458 (N_14458,N_13574,N_13818);
or U14459 (N_14459,N_13849,N_13988);
or U14460 (N_14460,N_13581,N_13653);
and U14461 (N_14461,N_13730,N_13561);
nor U14462 (N_14462,N_13814,N_13899);
or U14463 (N_14463,N_13733,N_13539);
or U14464 (N_14464,N_13708,N_13567);
nand U14465 (N_14465,N_13874,N_13598);
or U14466 (N_14466,N_13592,N_13714);
and U14467 (N_14467,N_13688,N_13515);
and U14468 (N_14468,N_13518,N_13866);
xnor U14469 (N_14469,N_13839,N_13754);
or U14470 (N_14470,N_13865,N_13774);
and U14471 (N_14471,N_13533,N_13616);
nand U14472 (N_14472,N_13608,N_13620);
and U14473 (N_14473,N_13571,N_13992);
nand U14474 (N_14474,N_13902,N_13575);
xnor U14475 (N_14475,N_13757,N_13549);
nand U14476 (N_14476,N_13726,N_13791);
nand U14477 (N_14477,N_13923,N_13586);
or U14478 (N_14478,N_13671,N_13860);
nand U14479 (N_14479,N_13828,N_13666);
nor U14480 (N_14480,N_13902,N_13504);
nor U14481 (N_14481,N_13626,N_13650);
nand U14482 (N_14482,N_13640,N_13981);
or U14483 (N_14483,N_13993,N_13516);
nor U14484 (N_14484,N_13745,N_13952);
and U14485 (N_14485,N_13622,N_13854);
and U14486 (N_14486,N_13708,N_13996);
and U14487 (N_14487,N_13599,N_13967);
or U14488 (N_14488,N_13962,N_13733);
xnor U14489 (N_14489,N_13980,N_13821);
and U14490 (N_14490,N_13851,N_13911);
nor U14491 (N_14491,N_13898,N_13643);
nand U14492 (N_14492,N_13814,N_13798);
or U14493 (N_14493,N_13910,N_13927);
and U14494 (N_14494,N_13790,N_13731);
or U14495 (N_14495,N_13665,N_13913);
nor U14496 (N_14496,N_13711,N_13518);
nand U14497 (N_14497,N_13655,N_13568);
or U14498 (N_14498,N_13806,N_13978);
nor U14499 (N_14499,N_13953,N_13768);
nand U14500 (N_14500,N_14391,N_14239);
and U14501 (N_14501,N_14120,N_14401);
nand U14502 (N_14502,N_14040,N_14305);
and U14503 (N_14503,N_14408,N_14381);
nor U14504 (N_14504,N_14439,N_14331);
nand U14505 (N_14505,N_14290,N_14048);
xor U14506 (N_14506,N_14246,N_14483);
or U14507 (N_14507,N_14458,N_14077);
and U14508 (N_14508,N_14224,N_14463);
and U14509 (N_14509,N_14476,N_14413);
and U14510 (N_14510,N_14314,N_14378);
nand U14511 (N_14511,N_14111,N_14176);
or U14512 (N_14512,N_14299,N_14128);
and U14513 (N_14513,N_14345,N_14193);
xnor U14514 (N_14514,N_14219,N_14127);
nand U14515 (N_14515,N_14002,N_14234);
nor U14516 (N_14516,N_14230,N_14313);
and U14517 (N_14517,N_14223,N_14280);
nor U14518 (N_14518,N_14461,N_14045);
nand U14519 (N_14519,N_14088,N_14247);
or U14520 (N_14520,N_14312,N_14450);
and U14521 (N_14521,N_14183,N_14058);
or U14522 (N_14522,N_14472,N_14008);
or U14523 (N_14523,N_14116,N_14188);
or U14524 (N_14524,N_14470,N_14428);
nand U14525 (N_14525,N_14110,N_14392);
nand U14526 (N_14526,N_14468,N_14455);
nand U14527 (N_14527,N_14409,N_14168);
nand U14528 (N_14528,N_14155,N_14497);
nand U14529 (N_14529,N_14207,N_14028);
nor U14530 (N_14530,N_14306,N_14379);
nor U14531 (N_14531,N_14030,N_14484);
nor U14532 (N_14532,N_14109,N_14293);
nor U14533 (N_14533,N_14160,N_14426);
nor U14534 (N_14534,N_14274,N_14205);
and U14535 (N_14535,N_14380,N_14245);
and U14536 (N_14536,N_14418,N_14369);
nand U14537 (N_14537,N_14161,N_14236);
nor U14538 (N_14538,N_14137,N_14356);
or U14539 (N_14539,N_14022,N_14098);
or U14540 (N_14540,N_14441,N_14184);
or U14541 (N_14541,N_14003,N_14320);
and U14542 (N_14542,N_14318,N_14104);
xor U14543 (N_14543,N_14297,N_14327);
nor U14544 (N_14544,N_14208,N_14258);
or U14545 (N_14545,N_14482,N_14368);
nand U14546 (N_14546,N_14226,N_14210);
nand U14547 (N_14547,N_14475,N_14415);
or U14548 (N_14548,N_14198,N_14485);
xor U14549 (N_14549,N_14097,N_14201);
nor U14550 (N_14550,N_14112,N_14133);
nor U14551 (N_14551,N_14342,N_14481);
nand U14552 (N_14552,N_14304,N_14411);
nand U14553 (N_14553,N_14227,N_14140);
and U14554 (N_14554,N_14449,N_14324);
nand U14555 (N_14555,N_14195,N_14148);
and U14556 (N_14556,N_14326,N_14167);
nor U14557 (N_14557,N_14071,N_14412);
or U14558 (N_14558,N_14102,N_14059);
nor U14559 (N_14559,N_14351,N_14100);
nand U14560 (N_14560,N_14041,N_14020);
xnor U14561 (N_14561,N_14464,N_14374);
xor U14562 (N_14562,N_14339,N_14039);
nor U14563 (N_14563,N_14123,N_14420);
nand U14564 (N_14564,N_14103,N_14432);
nor U14565 (N_14565,N_14062,N_14444);
or U14566 (N_14566,N_14156,N_14284);
and U14567 (N_14567,N_14135,N_14422);
nor U14568 (N_14568,N_14129,N_14256);
nor U14569 (N_14569,N_14169,N_14005);
nor U14570 (N_14570,N_14163,N_14084);
xnor U14571 (N_14571,N_14240,N_14090);
or U14572 (N_14572,N_14174,N_14179);
and U14573 (N_14573,N_14189,N_14141);
and U14574 (N_14574,N_14122,N_14480);
nor U14575 (N_14575,N_14125,N_14091);
and U14576 (N_14576,N_14081,N_14465);
xor U14577 (N_14577,N_14253,N_14117);
xnor U14578 (N_14578,N_14213,N_14267);
nand U14579 (N_14579,N_14279,N_14488);
xor U14580 (N_14580,N_14332,N_14056);
nand U14581 (N_14581,N_14442,N_14093);
nor U14582 (N_14582,N_14429,N_14263);
nor U14583 (N_14583,N_14440,N_14399);
and U14584 (N_14584,N_14474,N_14437);
and U14585 (N_14585,N_14285,N_14158);
or U14586 (N_14586,N_14233,N_14114);
or U14587 (N_14587,N_14283,N_14347);
and U14588 (N_14588,N_14487,N_14036);
nand U14589 (N_14589,N_14004,N_14011);
or U14590 (N_14590,N_14144,N_14073);
or U14591 (N_14591,N_14268,N_14244);
and U14592 (N_14592,N_14473,N_14309);
nand U14593 (N_14593,N_14180,N_14322);
xor U14594 (N_14594,N_14007,N_14499);
nand U14595 (N_14595,N_14107,N_14453);
nand U14596 (N_14596,N_14275,N_14371);
or U14597 (N_14597,N_14452,N_14080);
and U14598 (N_14598,N_14178,N_14350);
or U14599 (N_14599,N_14038,N_14072);
xor U14600 (N_14600,N_14282,N_14251);
nor U14601 (N_14601,N_14043,N_14489);
nand U14602 (N_14602,N_14266,N_14433);
and U14603 (N_14603,N_14330,N_14291);
nor U14604 (N_14604,N_14096,N_14383);
or U14605 (N_14605,N_14301,N_14436);
or U14606 (N_14606,N_14199,N_14054);
or U14607 (N_14607,N_14134,N_14288);
and U14608 (N_14608,N_14185,N_14190);
nand U14609 (N_14609,N_14065,N_14343);
nand U14610 (N_14610,N_14145,N_14435);
nand U14611 (N_14611,N_14310,N_14490);
xor U14612 (N_14612,N_14311,N_14362);
or U14613 (N_14613,N_14298,N_14006);
nor U14614 (N_14614,N_14010,N_14231);
xor U14615 (N_14615,N_14060,N_14232);
and U14616 (N_14616,N_14064,N_14493);
and U14617 (N_14617,N_14260,N_14067);
or U14618 (N_14618,N_14300,N_14321);
and U14619 (N_14619,N_14106,N_14448);
nand U14620 (N_14620,N_14346,N_14074);
and U14621 (N_14621,N_14486,N_14353);
and U14622 (N_14622,N_14099,N_14361);
nor U14623 (N_14623,N_14445,N_14172);
nor U14624 (N_14624,N_14042,N_14241);
or U14625 (N_14625,N_14218,N_14024);
nand U14626 (N_14626,N_14365,N_14272);
or U14627 (N_14627,N_14295,N_14216);
and U14628 (N_14628,N_14287,N_14431);
nor U14629 (N_14629,N_14079,N_14358);
xor U14630 (N_14630,N_14469,N_14457);
nor U14631 (N_14631,N_14397,N_14419);
or U14632 (N_14632,N_14063,N_14276);
or U14633 (N_14633,N_14083,N_14215);
and U14634 (N_14634,N_14037,N_14078);
xnor U14635 (N_14635,N_14124,N_14398);
and U14636 (N_14636,N_14328,N_14498);
and U14637 (N_14637,N_14393,N_14211);
and U14638 (N_14638,N_14115,N_14026);
nand U14639 (N_14639,N_14402,N_14089);
xnor U14640 (N_14640,N_14095,N_14375);
and U14641 (N_14641,N_14136,N_14446);
nand U14642 (N_14642,N_14220,N_14286);
nand U14643 (N_14643,N_14403,N_14460);
and U14644 (N_14644,N_14235,N_14066);
and U14645 (N_14645,N_14221,N_14173);
xor U14646 (N_14646,N_14143,N_14162);
nor U14647 (N_14647,N_14495,N_14349);
or U14648 (N_14648,N_14018,N_14139);
and U14649 (N_14649,N_14447,N_14019);
and U14650 (N_14650,N_14000,N_14254);
nor U14651 (N_14651,N_14334,N_14242);
or U14652 (N_14652,N_14153,N_14278);
and U14653 (N_14653,N_14118,N_14259);
or U14654 (N_14654,N_14296,N_14146);
or U14655 (N_14655,N_14092,N_14108);
or U14656 (N_14656,N_14336,N_14410);
and U14657 (N_14657,N_14270,N_14434);
nand U14658 (N_14658,N_14255,N_14105);
nor U14659 (N_14659,N_14425,N_14191);
nor U14660 (N_14660,N_14491,N_14166);
or U14661 (N_14661,N_14204,N_14262);
nor U14662 (N_14662,N_14225,N_14170);
and U14663 (N_14663,N_14494,N_14055);
nor U14664 (N_14664,N_14335,N_14138);
xnor U14665 (N_14665,N_14212,N_14338);
xnor U14666 (N_14666,N_14049,N_14289);
and U14667 (N_14667,N_14407,N_14373);
or U14668 (N_14668,N_14243,N_14017);
and U14669 (N_14669,N_14113,N_14366);
and U14670 (N_14670,N_14033,N_14387);
nor U14671 (N_14671,N_14119,N_14222);
or U14672 (N_14672,N_14360,N_14386);
and U14673 (N_14673,N_14249,N_14023);
xnor U14674 (N_14674,N_14405,N_14325);
nand U14675 (N_14675,N_14237,N_14238);
xor U14676 (N_14676,N_14132,N_14376);
nor U14677 (N_14677,N_14151,N_14389);
nor U14678 (N_14678,N_14094,N_14196);
and U14679 (N_14679,N_14308,N_14150);
or U14680 (N_14680,N_14131,N_14404);
or U14681 (N_14681,N_14187,N_14016);
and U14682 (N_14682,N_14467,N_14029);
nor U14683 (N_14683,N_14307,N_14250);
or U14684 (N_14684,N_14027,N_14157);
or U14685 (N_14685,N_14229,N_14316);
nor U14686 (N_14686,N_14479,N_14101);
or U14687 (N_14687,N_14076,N_14477);
and U14688 (N_14688,N_14165,N_14388);
and U14689 (N_14689,N_14031,N_14082);
nor U14690 (N_14690,N_14175,N_14364);
and U14691 (N_14691,N_14044,N_14385);
xor U14692 (N_14692,N_14303,N_14206);
nor U14693 (N_14693,N_14032,N_14438);
and U14694 (N_14694,N_14035,N_14086);
or U14695 (N_14695,N_14394,N_14340);
and U14696 (N_14696,N_14069,N_14248);
or U14697 (N_14697,N_14430,N_14462);
nor U14698 (N_14698,N_14302,N_14152);
or U14699 (N_14699,N_14012,N_14214);
nor U14700 (N_14700,N_14478,N_14087);
nor U14701 (N_14701,N_14068,N_14363);
or U14702 (N_14702,N_14142,N_14203);
or U14703 (N_14703,N_14057,N_14015);
nand U14704 (N_14704,N_14421,N_14269);
and U14705 (N_14705,N_14281,N_14021);
xnor U14706 (N_14706,N_14417,N_14228);
nor U14707 (N_14707,N_14423,N_14454);
nand U14708 (N_14708,N_14341,N_14492);
nor U14709 (N_14709,N_14025,N_14271);
nand U14710 (N_14710,N_14277,N_14427);
xor U14711 (N_14711,N_14046,N_14384);
xnor U14712 (N_14712,N_14070,N_14451);
nand U14713 (N_14713,N_14406,N_14209);
nand U14714 (N_14714,N_14352,N_14182);
nand U14715 (N_14715,N_14085,N_14424);
or U14716 (N_14716,N_14466,N_14355);
nor U14717 (N_14717,N_14323,N_14001);
nor U14718 (N_14718,N_14329,N_14075);
or U14719 (N_14719,N_14443,N_14257);
nand U14720 (N_14720,N_14382,N_14186);
nand U14721 (N_14721,N_14292,N_14202);
xnor U14722 (N_14722,N_14192,N_14052);
xor U14723 (N_14723,N_14390,N_14459);
nand U14724 (N_14724,N_14456,N_14264);
and U14725 (N_14725,N_14265,N_14344);
xor U14726 (N_14726,N_14496,N_14273);
or U14727 (N_14727,N_14171,N_14014);
or U14728 (N_14728,N_14252,N_14181);
or U14729 (N_14729,N_14154,N_14333);
or U14730 (N_14730,N_14317,N_14471);
or U14731 (N_14731,N_14315,N_14400);
and U14732 (N_14732,N_14200,N_14414);
nand U14733 (N_14733,N_14009,N_14121);
or U14734 (N_14734,N_14034,N_14359);
nor U14735 (N_14735,N_14416,N_14367);
or U14736 (N_14736,N_14348,N_14377);
nand U14737 (N_14737,N_14194,N_14053);
nor U14738 (N_14738,N_14197,N_14051);
xor U14739 (N_14739,N_14149,N_14370);
nor U14740 (N_14740,N_14357,N_14013);
nor U14741 (N_14741,N_14372,N_14261);
or U14742 (N_14742,N_14294,N_14159);
and U14743 (N_14743,N_14217,N_14047);
and U14744 (N_14744,N_14130,N_14395);
xor U14745 (N_14745,N_14164,N_14319);
nand U14746 (N_14746,N_14050,N_14061);
nor U14747 (N_14747,N_14126,N_14354);
nor U14748 (N_14748,N_14147,N_14177);
or U14749 (N_14749,N_14337,N_14396);
nor U14750 (N_14750,N_14304,N_14286);
or U14751 (N_14751,N_14073,N_14238);
nand U14752 (N_14752,N_14069,N_14383);
nand U14753 (N_14753,N_14202,N_14273);
nor U14754 (N_14754,N_14200,N_14378);
xor U14755 (N_14755,N_14029,N_14419);
and U14756 (N_14756,N_14017,N_14437);
and U14757 (N_14757,N_14409,N_14359);
nand U14758 (N_14758,N_14338,N_14172);
nor U14759 (N_14759,N_14245,N_14198);
and U14760 (N_14760,N_14223,N_14405);
or U14761 (N_14761,N_14315,N_14077);
or U14762 (N_14762,N_14273,N_14149);
and U14763 (N_14763,N_14278,N_14266);
or U14764 (N_14764,N_14188,N_14458);
and U14765 (N_14765,N_14376,N_14488);
nand U14766 (N_14766,N_14308,N_14430);
nor U14767 (N_14767,N_14452,N_14084);
and U14768 (N_14768,N_14033,N_14167);
or U14769 (N_14769,N_14086,N_14410);
nand U14770 (N_14770,N_14217,N_14049);
xor U14771 (N_14771,N_14305,N_14379);
nor U14772 (N_14772,N_14350,N_14480);
nor U14773 (N_14773,N_14426,N_14163);
nor U14774 (N_14774,N_14259,N_14293);
and U14775 (N_14775,N_14370,N_14151);
nand U14776 (N_14776,N_14205,N_14254);
nor U14777 (N_14777,N_14187,N_14010);
nor U14778 (N_14778,N_14110,N_14348);
nor U14779 (N_14779,N_14020,N_14322);
nor U14780 (N_14780,N_14217,N_14207);
nand U14781 (N_14781,N_14087,N_14266);
or U14782 (N_14782,N_14177,N_14155);
or U14783 (N_14783,N_14245,N_14022);
nand U14784 (N_14784,N_14348,N_14075);
nand U14785 (N_14785,N_14423,N_14004);
and U14786 (N_14786,N_14196,N_14156);
and U14787 (N_14787,N_14483,N_14374);
and U14788 (N_14788,N_14273,N_14410);
or U14789 (N_14789,N_14405,N_14231);
xnor U14790 (N_14790,N_14475,N_14089);
nand U14791 (N_14791,N_14337,N_14107);
xor U14792 (N_14792,N_14183,N_14049);
or U14793 (N_14793,N_14060,N_14234);
or U14794 (N_14794,N_14491,N_14161);
nor U14795 (N_14795,N_14052,N_14039);
or U14796 (N_14796,N_14000,N_14444);
and U14797 (N_14797,N_14233,N_14343);
nand U14798 (N_14798,N_14215,N_14491);
or U14799 (N_14799,N_14333,N_14448);
nor U14800 (N_14800,N_14230,N_14226);
and U14801 (N_14801,N_14211,N_14295);
nor U14802 (N_14802,N_14163,N_14061);
or U14803 (N_14803,N_14133,N_14447);
nor U14804 (N_14804,N_14144,N_14054);
and U14805 (N_14805,N_14384,N_14168);
nand U14806 (N_14806,N_14003,N_14128);
nand U14807 (N_14807,N_14168,N_14333);
nor U14808 (N_14808,N_14257,N_14426);
or U14809 (N_14809,N_14337,N_14233);
nor U14810 (N_14810,N_14221,N_14128);
nand U14811 (N_14811,N_14144,N_14400);
nand U14812 (N_14812,N_14050,N_14432);
and U14813 (N_14813,N_14171,N_14380);
or U14814 (N_14814,N_14223,N_14007);
or U14815 (N_14815,N_14195,N_14398);
nor U14816 (N_14816,N_14215,N_14068);
nand U14817 (N_14817,N_14401,N_14057);
nand U14818 (N_14818,N_14458,N_14125);
and U14819 (N_14819,N_14344,N_14458);
or U14820 (N_14820,N_14347,N_14049);
xor U14821 (N_14821,N_14142,N_14129);
nor U14822 (N_14822,N_14466,N_14202);
or U14823 (N_14823,N_14348,N_14247);
nand U14824 (N_14824,N_14007,N_14466);
nor U14825 (N_14825,N_14012,N_14306);
xor U14826 (N_14826,N_14072,N_14182);
and U14827 (N_14827,N_14339,N_14207);
nor U14828 (N_14828,N_14428,N_14389);
nor U14829 (N_14829,N_14043,N_14033);
and U14830 (N_14830,N_14045,N_14218);
nand U14831 (N_14831,N_14321,N_14460);
nand U14832 (N_14832,N_14300,N_14367);
nand U14833 (N_14833,N_14038,N_14491);
or U14834 (N_14834,N_14112,N_14496);
nor U14835 (N_14835,N_14044,N_14414);
or U14836 (N_14836,N_14136,N_14351);
nand U14837 (N_14837,N_14230,N_14416);
or U14838 (N_14838,N_14466,N_14345);
nor U14839 (N_14839,N_14349,N_14426);
or U14840 (N_14840,N_14093,N_14284);
nand U14841 (N_14841,N_14418,N_14233);
or U14842 (N_14842,N_14156,N_14431);
and U14843 (N_14843,N_14140,N_14410);
and U14844 (N_14844,N_14489,N_14215);
nor U14845 (N_14845,N_14128,N_14372);
and U14846 (N_14846,N_14383,N_14399);
nor U14847 (N_14847,N_14290,N_14346);
and U14848 (N_14848,N_14304,N_14428);
or U14849 (N_14849,N_14409,N_14157);
and U14850 (N_14850,N_14169,N_14255);
and U14851 (N_14851,N_14360,N_14025);
nand U14852 (N_14852,N_14297,N_14171);
and U14853 (N_14853,N_14488,N_14023);
nor U14854 (N_14854,N_14168,N_14067);
xnor U14855 (N_14855,N_14209,N_14213);
nor U14856 (N_14856,N_14174,N_14131);
nor U14857 (N_14857,N_14109,N_14008);
and U14858 (N_14858,N_14095,N_14220);
xnor U14859 (N_14859,N_14433,N_14423);
xor U14860 (N_14860,N_14176,N_14197);
xor U14861 (N_14861,N_14499,N_14381);
or U14862 (N_14862,N_14402,N_14259);
nand U14863 (N_14863,N_14188,N_14387);
nand U14864 (N_14864,N_14260,N_14153);
or U14865 (N_14865,N_14177,N_14302);
and U14866 (N_14866,N_14157,N_14205);
nor U14867 (N_14867,N_14483,N_14429);
xnor U14868 (N_14868,N_14456,N_14094);
nor U14869 (N_14869,N_14436,N_14413);
nand U14870 (N_14870,N_14045,N_14400);
and U14871 (N_14871,N_14346,N_14296);
and U14872 (N_14872,N_14069,N_14391);
xnor U14873 (N_14873,N_14069,N_14200);
or U14874 (N_14874,N_14181,N_14353);
nand U14875 (N_14875,N_14170,N_14366);
nand U14876 (N_14876,N_14137,N_14348);
and U14877 (N_14877,N_14490,N_14471);
xnor U14878 (N_14878,N_14485,N_14036);
nand U14879 (N_14879,N_14208,N_14433);
or U14880 (N_14880,N_14003,N_14126);
nand U14881 (N_14881,N_14096,N_14346);
nand U14882 (N_14882,N_14071,N_14083);
or U14883 (N_14883,N_14027,N_14386);
or U14884 (N_14884,N_14432,N_14253);
or U14885 (N_14885,N_14202,N_14339);
nand U14886 (N_14886,N_14452,N_14473);
or U14887 (N_14887,N_14035,N_14346);
or U14888 (N_14888,N_14350,N_14392);
nor U14889 (N_14889,N_14089,N_14469);
and U14890 (N_14890,N_14425,N_14018);
nand U14891 (N_14891,N_14446,N_14418);
or U14892 (N_14892,N_14245,N_14033);
nand U14893 (N_14893,N_14084,N_14052);
or U14894 (N_14894,N_14122,N_14299);
or U14895 (N_14895,N_14148,N_14402);
xor U14896 (N_14896,N_14315,N_14117);
or U14897 (N_14897,N_14225,N_14485);
nor U14898 (N_14898,N_14057,N_14361);
nor U14899 (N_14899,N_14079,N_14386);
nor U14900 (N_14900,N_14184,N_14414);
and U14901 (N_14901,N_14474,N_14408);
nand U14902 (N_14902,N_14466,N_14330);
nor U14903 (N_14903,N_14240,N_14046);
nor U14904 (N_14904,N_14058,N_14251);
and U14905 (N_14905,N_14131,N_14082);
nor U14906 (N_14906,N_14153,N_14017);
and U14907 (N_14907,N_14324,N_14306);
and U14908 (N_14908,N_14430,N_14304);
nand U14909 (N_14909,N_14453,N_14393);
nor U14910 (N_14910,N_14295,N_14236);
nor U14911 (N_14911,N_14294,N_14306);
nor U14912 (N_14912,N_14091,N_14183);
and U14913 (N_14913,N_14408,N_14004);
or U14914 (N_14914,N_14298,N_14486);
or U14915 (N_14915,N_14182,N_14083);
nor U14916 (N_14916,N_14287,N_14457);
nand U14917 (N_14917,N_14082,N_14212);
or U14918 (N_14918,N_14127,N_14499);
or U14919 (N_14919,N_14347,N_14162);
nor U14920 (N_14920,N_14335,N_14444);
or U14921 (N_14921,N_14156,N_14430);
nand U14922 (N_14922,N_14138,N_14470);
nand U14923 (N_14923,N_14436,N_14254);
or U14924 (N_14924,N_14256,N_14213);
nand U14925 (N_14925,N_14074,N_14044);
and U14926 (N_14926,N_14390,N_14388);
nand U14927 (N_14927,N_14314,N_14057);
and U14928 (N_14928,N_14357,N_14019);
nor U14929 (N_14929,N_14474,N_14385);
or U14930 (N_14930,N_14238,N_14426);
or U14931 (N_14931,N_14217,N_14429);
and U14932 (N_14932,N_14163,N_14409);
nor U14933 (N_14933,N_14368,N_14158);
or U14934 (N_14934,N_14303,N_14148);
nor U14935 (N_14935,N_14438,N_14045);
and U14936 (N_14936,N_14053,N_14267);
nor U14937 (N_14937,N_14139,N_14176);
nand U14938 (N_14938,N_14058,N_14484);
and U14939 (N_14939,N_14459,N_14489);
nor U14940 (N_14940,N_14143,N_14059);
or U14941 (N_14941,N_14486,N_14267);
and U14942 (N_14942,N_14377,N_14457);
and U14943 (N_14943,N_14257,N_14246);
xor U14944 (N_14944,N_14034,N_14240);
nor U14945 (N_14945,N_14301,N_14420);
and U14946 (N_14946,N_14414,N_14001);
or U14947 (N_14947,N_14063,N_14136);
xnor U14948 (N_14948,N_14015,N_14082);
nand U14949 (N_14949,N_14003,N_14364);
nand U14950 (N_14950,N_14267,N_14436);
or U14951 (N_14951,N_14033,N_14140);
nand U14952 (N_14952,N_14188,N_14135);
nand U14953 (N_14953,N_14244,N_14090);
nand U14954 (N_14954,N_14179,N_14437);
and U14955 (N_14955,N_14299,N_14117);
and U14956 (N_14956,N_14166,N_14206);
nor U14957 (N_14957,N_14144,N_14200);
nand U14958 (N_14958,N_14450,N_14199);
and U14959 (N_14959,N_14128,N_14135);
nor U14960 (N_14960,N_14026,N_14405);
nor U14961 (N_14961,N_14431,N_14250);
and U14962 (N_14962,N_14014,N_14239);
or U14963 (N_14963,N_14102,N_14125);
or U14964 (N_14964,N_14219,N_14446);
xnor U14965 (N_14965,N_14317,N_14197);
xor U14966 (N_14966,N_14125,N_14425);
xor U14967 (N_14967,N_14297,N_14188);
or U14968 (N_14968,N_14437,N_14225);
nor U14969 (N_14969,N_14117,N_14166);
nand U14970 (N_14970,N_14325,N_14005);
or U14971 (N_14971,N_14409,N_14018);
or U14972 (N_14972,N_14221,N_14160);
nand U14973 (N_14973,N_14137,N_14493);
nand U14974 (N_14974,N_14092,N_14217);
nor U14975 (N_14975,N_14414,N_14284);
or U14976 (N_14976,N_14141,N_14304);
nand U14977 (N_14977,N_14053,N_14398);
and U14978 (N_14978,N_14378,N_14312);
nor U14979 (N_14979,N_14418,N_14237);
and U14980 (N_14980,N_14043,N_14130);
or U14981 (N_14981,N_14362,N_14473);
or U14982 (N_14982,N_14255,N_14259);
or U14983 (N_14983,N_14413,N_14475);
nor U14984 (N_14984,N_14199,N_14241);
nor U14985 (N_14985,N_14343,N_14017);
and U14986 (N_14986,N_14287,N_14011);
and U14987 (N_14987,N_14179,N_14473);
and U14988 (N_14988,N_14309,N_14146);
and U14989 (N_14989,N_14434,N_14478);
nand U14990 (N_14990,N_14488,N_14039);
nor U14991 (N_14991,N_14054,N_14384);
nand U14992 (N_14992,N_14170,N_14006);
nor U14993 (N_14993,N_14280,N_14493);
nand U14994 (N_14994,N_14095,N_14083);
nor U14995 (N_14995,N_14027,N_14175);
xor U14996 (N_14996,N_14221,N_14418);
nor U14997 (N_14997,N_14202,N_14423);
and U14998 (N_14998,N_14257,N_14249);
xnor U14999 (N_14999,N_14197,N_14386);
and UO_0 (O_0,N_14988,N_14576);
or UO_1 (O_1,N_14931,N_14985);
and UO_2 (O_2,N_14663,N_14643);
and UO_3 (O_3,N_14540,N_14513);
nor UO_4 (O_4,N_14873,N_14788);
xnor UO_5 (O_5,N_14564,N_14942);
nor UO_6 (O_6,N_14950,N_14972);
nor UO_7 (O_7,N_14568,N_14994);
or UO_8 (O_8,N_14516,N_14780);
xnor UO_9 (O_9,N_14782,N_14687);
nand UO_10 (O_10,N_14597,N_14562);
and UO_11 (O_11,N_14818,N_14758);
or UO_12 (O_12,N_14651,N_14908);
or UO_13 (O_13,N_14791,N_14830);
nand UO_14 (O_14,N_14677,N_14882);
nand UO_15 (O_15,N_14606,N_14550);
or UO_16 (O_16,N_14879,N_14593);
nand UO_17 (O_17,N_14583,N_14841);
or UO_18 (O_18,N_14948,N_14526);
nor UO_19 (O_19,N_14904,N_14610);
or UO_20 (O_20,N_14870,N_14525);
and UO_21 (O_21,N_14502,N_14536);
nor UO_22 (O_22,N_14871,N_14699);
or UO_23 (O_23,N_14921,N_14968);
nor UO_24 (O_24,N_14944,N_14505);
or UO_25 (O_25,N_14973,N_14746);
xor UO_26 (O_26,N_14855,N_14507);
nor UO_27 (O_27,N_14979,N_14567);
nand UO_28 (O_28,N_14509,N_14519);
and UO_29 (O_29,N_14869,N_14798);
and UO_30 (O_30,N_14611,N_14962);
nand UO_31 (O_31,N_14969,N_14572);
nor UO_32 (O_32,N_14660,N_14898);
or UO_33 (O_33,N_14963,N_14949);
nand UO_34 (O_34,N_14883,N_14637);
and UO_35 (O_35,N_14607,N_14551);
nor UO_36 (O_36,N_14807,N_14654);
or UO_37 (O_37,N_14534,N_14999);
and UO_38 (O_38,N_14947,N_14877);
nor UO_39 (O_39,N_14806,N_14813);
nor UO_40 (O_40,N_14679,N_14874);
nor UO_41 (O_41,N_14658,N_14613);
and UO_42 (O_42,N_14601,N_14899);
and UO_43 (O_43,N_14808,N_14965);
and UO_44 (O_44,N_14858,N_14638);
nor UO_45 (O_45,N_14903,N_14932);
nand UO_46 (O_46,N_14639,N_14835);
xnor UO_47 (O_47,N_14728,N_14723);
nand UO_48 (O_48,N_14569,N_14574);
nor UO_49 (O_49,N_14515,N_14853);
or UO_50 (O_50,N_14622,N_14795);
nand UO_51 (O_51,N_14749,N_14907);
or UO_52 (O_52,N_14784,N_14804);
nor UO_53 (O_53,N_14836,N_14681);
and UO_54 (O_54,N_14822,N_14900);
nor UO_55 (O_55,N_14765,N_14762);
and UO_56 (O_56,N_14840,N_14720);
nor UO_57 (O_57,N_14817,N_14916);
nor UO_58 (O_58,N_14744,N_14825);
xnor UO_59 (O_59,N_14716,N_14761);
nand UO_60 (O_60,N_14529,N_14794);
nand UO_61 (O_61,N_14545,N_14508);
and UO_62 (O_62,N_14919,N_14966);
nand UO_63 (O_63,N_14714,N_14546);
or UO_64 (O_64,N_14997,N_14700);
and UO_65 (O_65,N_14821,N_14575);
or UO_66 (O_66,N_14543,N_14960);
nand UO_67 (O_67,N_14920,N_14558);
or UO_68 (O_68,N_14838,N_14777);
nor UO_69 (O_69,N_14633,N_14629);
and UO_70 (O_70,N_14537,N_14987);
xor UO_71 (O_71,N_14748,N_14731);
nor UO_72 (O_72,N_14565,N_14696);
or UO_73 (O_73,N_14672,N_14937);
nand UO_74 (O_74,N_14646,N_14592);
xor UO_75 (O_75,N_14602,N_14938);
nor UO_76 (O_76,N_14880,N_14902);
or UO_77 (O_77,N_14834,N_14689);
or UO_78 (O_78,N_14781,N_14673);
or UO_79 (O_79,N_14630,N_14640);
or UO_80 (O_80,N_14741,N_14694);
xnor UO_81 (O_81,N_14952,N_14676);
xnor UO_82 (O_82,N_14770,N_14506);
nand UO_83 (O_83,N_14935,N_14512);
and UO_84 (O_84,N_14599,N_14998);
nor UO_85 (O_85,N_14905,N_14692);
xnor UO_86 (O_86,N_14789,N_14596);
and UO_87 (O_87,N_14589,N_14582);
nor UO_88 (O_88,N_14577,N_14895);
and UO_89 (O_89,N_14925,N_14605);
or UO_90 (O_90,N_14736,N_14740);
xor UO_91 (O_91,N_14738,N_14754);
nor UO_92 (O_92,N_14957,N_14984);
nand UO_93 (O_93,N_14786,N_14685);
or UO_94 (O_94,N_14612,N_14553);
nor UO_95 (O_95,N_14704,N_14678);
and UO_96 (O_96,N_14702,N_14655);
nand UO_97 (O_97,N_14839,N_14697);
or UO_98 (O_98,N_14636,N_14570);
or UO_99 (O_99,N_14632,N_14701);
or UO_100 (O_100,N_14620,N_14976);
or UO_101 (O_101,N_14983,N_14743);
and UO_102 (O_102,N_14800,N_14941);
xnor UO_103 (O_103,N_14946,N_14820);
xnor UO_104 (O_104,N_14524,N_14739);
xor UO_105 (O_105,N_14757,N_14707);
nor UO_106 (O_106,N_14766,N_14747);
nor UO_107 (O_107,N_14667,N_14772);
and UO_108 (O_108,N_14793,N_14527);
nand UO_109 (O_109,N_14811,N_14729);
nand UO_110 (O_110,N_14559,N_14971);
and UO_111 (O_111,N_14737,N_14730);
nor UO_112 (O_112,N_14974,N_14852);
or UO_113 (O_113,N_14913,N_14609);
xnor UO_114 (O_114,N_14859,N_14846);
nand UO_115 (O_115,N_14625,N_14719);
and UO_116 (O_116,N_14892,N_14764);
and UO_117 (O_117,N_14863,N_14554);
xnor UO_118 (O_118,N_14992,N_14563);
or UO_119 (O_119,N_14504,N_14889);
or UO_120 (O_120,N_14549,N_14671);
and UO_121 (O_121,N_14796,N_14929);
nand UO_122 (O_122,N_14649,N_14996);
and UO_123 (O_123,N_14684,N_14816);
nand UO_124 (O_124,N_14901,N_14652);
or UO_125 (O_125,N_14680,N_14928);
and UO_126 (O_126,N_14664,N_14893);
and UO_127 (O_127,N_14557,N_14862);
nand UO_128 (O_128,N_14724,N_14878);
and UO_129 (O_129,N_14691,N_14851);
and UO_130 (O_130,N_14734,N_14715);
and UO_131 (O_131,N_14939,N_14887);
xnor UO_132 (O_132,N_14587,N_14857);
and UO_133 (O_133,N_14964,N_14888);
nand UO_134 (O_134,N_14837,N_14531);
or UO_135 (O_135,N_14717,N_14805);
and UO_136 (O_136,N_14961,N_14849);
and UO_137 (O_137,N_14528,N_14521);
or UO_138 (O_138,N_14981,N_14539);
or UO_139 (O_139,N_14656,N_14756);
and UO_140 (O_140,N_14759,N_14867);
xnor UO_141 (O_141,N_14909,N_14922);
nor UO_142 (O_142,N_14769,N_14918);
or UO_143 (O_143,N_14912,N_14978);
nand UO_144 (O_144,N_14864,N_14634);
and UO_145 (O_145,N_14865,N_14991);
nand UO_146 (O_146,N_14631,N_14955);
nor UO_147 (O_147,N_14690,N_14647);
nand UO_148 (O_148,N_14683,N_14735);
nand UO_149 (O_149,N_14686,N_14866);
or UO_150 (O_150,N_14666,N_14624);
xnor UO_151 (O_151,N_14608,N_14911);
and UO_152 (O_152,N_14590,N_14580);
nor UO_153 (O_153,N_14617,N_14982);
nor UO_154 (O_154,N_14775,N_14668);
and UO_155 (O_155,N_14518,N_14776);
nand UO_156 (O_156,N_14532,N_14614);
or UO_157 (O_157,N_14819,N_14923);
xnor UO_158 (O_158,N_14986,N_14774);
or UO_159 (O_159,N_14659,N_14635);
or UO_160 (O_160,N_14522,N_14760);
and UO_161 (O_161,N_14560,N_14896);
or UO_162 (O_162,N_14779,N_14975);
and UO_163 (O_163,N_14915,N_14588);
and UO_164 (O_164,N_14885,N_14709);
nand UO_165 (O_165,N_14803,N_14586);
and UO_166 (O_166,N_14530,N_14773);
nor UO_167 (O_167,N_14872,N_14619);
and UO_168 (O_168,N_14967,N_14600);
nor UO_169 (O_169,N_14703,N_14827);
nand UO_170 (O_170,N_14875,N_14542);
and UO_171 (O_171,N_14732,N_14768);
nand UO_172 (O_172,N_14725,N_14641);
and UO_173 (O_173,N_14763,N_14675);
nand UO_174 (O_174,N_14812,N_14809);
nand UO_175 (O_175,N_14881,N_14850);
or UO_176 (O_176,N_14648,N_14712);
and UO_177 (O_177,N_14722,N_14706);
nor UO_178 (O_178,N_14644,N_14814);
nand UO_179 (O_179,N_14726,N_14848);
nand UO_180 (O_180,N_14603,N_14956);
nand UO_181 (O_181,N_14868,N_14933);
and UO_182 (O_182,N_14906,N_14626);
and UO_183 (O_183,N_14914,N_14894);
and UO_184 (O_184,N_14662,N_14801);
or UO_185 (O_185,N_14615,N_14934);
nand UO_186 (O_186,N_14833,N_14831);
or UO_187 (O_187,N_14510,N_14556);
xnor UO_188 (O_188,N_14594,N_14778);
or UO_189 (O_189,N_14854,N_14604);
nand UO_190 (O_190,N_14710,N_14823);
or UO_191 (O_191,N_14876,N_14653);
nor UO_192 (O_192,N_14520,N_14891);
or UO_193 (O_193,N_14733,N_14797);
nor UO_194 (O_194,N_14623,N_14936);
nor UO_195 (O_195,N_14787,N_14755);
nor UO_196 (O_196,N_14721,N_14753);
nor UO_197 (O_197,N_14541,N_14953);
nor UO_198 (O_198,N_14514,N_14977);
nand UO_199 (O_199,N_14552,N_14951);
or UO_200 (O_200,N_14943,N_14785);
or UO_201 (O_201,N_14897,N_14581);
xnor UO_202 (O_202,N_14860,N_14711);
nor UO_203 (O_203,N_14561,N_14555);
or UO_204 (O_204,N_14669,N_14566);
nand UO_205 (O_205,N_14705,N_14954);
and UO_206 (O_206,N_14799,N_14995);
nor UO_207 (O_207,N_14970,N_14815);
xnor UO_208 (O_208,N_14650,N_14958);
and UO_209 (O_209,N_14642,N_14548);
and UO_210 (O_210,N_14598,N_14616);
or UO_211 (O_211,N_14665,N_14628);
or UO_212 (O_212,N_14783,N_14674);
nand UO_213 (O_213,N_14727,N_14627);
nand UO_214 (O_214,N_14790,N_14945);
or UO_215 (O_215,N_14584,N_14591);
nand UO_216 (O_216,N_14752,N_14926);
or UO_217 (O_217,N_14856,N_14886);
nor UO_218 (O_218,N_14924,N_14890);
nand UO_219 (O_219,N_14573,N_14661);
or UO_220 (O_220,N_14501,N_14708);
nand UO_221 (O_221,N_14917,N_14861);
nor UO_222 (O_222,N_14989,N_14693);
and UO_223 (O_223,N_14578,N_14824);
or UO_224 (O_224,N_14845,N_14993);
nor UO_225 (O_225,N_14884,N_14792);
nor UO_226 (O_226,N_14802,N_14511);
nand UO_227 (O_227,N_14535,N_14980);
nand UO_228 (O_228,N_14523,N_14828);
or UO_229 (O_229,N_14930,N_14645);
or UO_230 (O_230,N_14595,N_14698);
nor UO_231 (O_231,N_14843,N_14910);
nand UO_232 (O_232,N_14751,N_14618);
or UO_233 (O_233,N_14829,N_14959);
and UO_234 (O_234,N_14621,N_14670);
and UO_235 (O_235,N_14844,N_14547);
or UO_236 (O_236,N_14927,N_14767);
and UO_237 (O_237,N_14533,N_14832);
nor UO_238 (O_238,N_14585,N_14745);
or UO_239 (O_239,N_14657,N_14750);
and UO_240 (O_240,N_14847,N_14538);
and UO_241 (O_241,N_14810,N_14771);
nand UO_242 (O_242,N_14990,N_14682);
or UO_243 (O_243,N_14579,N_14713);
nand UO_244 (O_244,N_14940,N_14718);
xnor UO_245 (O_245,N_14826,N_14503);
and UO_246 (O_246,N_14517,N_14571);
or UO_247 (O_247,N_14695,N_14544);
or UO_248 (O_248,N_14842,N_14688);
nor UO_249 (O_249,N_14742,N_14500);
and UO_250 (O_250,N_14594,N_14619);
or UO_251 (O_251,N_14634,N_14785);
or UO_252 (O_252,N_14818,N_14645);
and UO_253 (O_253,N_14887,N_14905);
xor UO_254 (O_254,N_14593,N_14575);
nand UO_255 (O_255,N_14971,N_14721);
xnor UO_256 (O_256,N_14782,N_14873);
and UO_257 (O_257,N_14646,N_14856);
nor UO_258 (O_258,N_14784,N_14717);
and UO_259 (O_259,N_14963,N_14883);
nand UO_260 (O_260,N_14738,N_14683);
and UO_261 (O_261,N_14502,N_14700);
nor UO_262 (O_262,N_14846,N_14540);
nand UO_263 (O_263,N_14897,N_14631);
and UO_264 (O_264,N_14824,N_14894);
and UO_265 (O_265,N_14652,N_14851);
nor UO_266 (O_266,N_14681,N_14995);
nor UO_267 (O_267,N_14833,N_14908);
nand UO_268 (O_268,N_14825,N_14616);
and UO_269 (O_269,N_14897,N_14602);
nand UO_270 (O_270,N_14844,N_14953);
nor UO_271 (O_271,N_14973,N_14767);
or UO_272 (O_272,N_14810,N_14980);
and UO_273 (O_273,N_14512,N_14823);
or UO_274 (O_274,N_14628,N_14967);
nor UO_275 (O_275,N_14888,N_14833);
or UO_276 (O_276,N_14778,N_14546);
or UO_277 (O_277,N_14863,N_14851);
nor UO_278 (O_278,N_14661,N_14987);
nor UO_279 (O_279,N_14927,N_14595);
or UO_280 (O_280,N_14578,N_14823);
nand UO_281 (O_281,N_14918,N_14573);
and UO_282 (O_282,N_14606,N_14514);
nor UO_283 (O_283,N_14638,N_14836);
and UO_284 (O_284,N_14830,N_14803);
nor UO_285 (O_285,N_14585,N_14896);
nor UO_286 (O_286,N_14671,N_14751);
nor UO_287 (O_287,N_14755,N_14779);
nand UO_288 (O_288,N_14998,N_14842);
nor UO_289 (O_289,N_14501,N_14709);
or UO_290 (O_290,N_14752,N_14537);
nand UO_291 (O_291,N_14501,N_14853);
nor UO_292 (O_292,N_14683,N_14889);
or UO_293 (O_293,N_14637,N_14504);
nor UO_294 (O_294,N_14639,N_14612);
nand UO_295 (O_295,N_14757,N_14977);
nand UO_296 (O_296,N_14792,N_14666);
nor UO_297 (O_297,N_14525,N_14877);
and UO_298 (O_298,N_14905,N_14854);
nand UO_299 (O_299,N_14913,N_14885);
nand UO_300 (O_300,N_14772,N_14991);
or UO_301 (O_301,N_14602,N_14949);
and UO_302 (O_302,N_14660,N_14694);
or UO_303 (O_303,N_14512,N_14965);
nand UO_304 (O_304,N_14766,N_14938);
and UO_305 (O_305,N_14681,N_14812);
xnor UO_306 (O_306,N_14742,N_14846);
nand UO_307 (O_307,N_14799,N_14820);
and UO_308 (O_308,N_14565,N_14647);
nand UO_309 (O_309,N_14631,N_14513);
or UO_310 (O_310,N_14987,N_14503);
or UO_311 (O_311,N_14752,N_14675);
xor UO_312 (O_312,N_14851,N_14778);
or UO_313 (O_313,N_14723,N_14856);
nand UO_314 (O_314,N_14847,N_14741);
and UO_315 (O_315,N_14616,N_14644);
nand UO_316 (O_316,N_14648,N_14541);
nand UO_317 (O_317,N_14601,N_14596);
nor UO_318 (O_318,N_14550,N_14788);
nor UO_319 (O_319,N_14572,N_14762);
and UO_320 (O_320,N_14648,N_14522);
nor UO_321 (O_321,N_14992,N_14952);
nand UO_322 (O_322,N_14692,N_14599);
nand UO_323 (O_323,N_14877,N_14919);
or UO_324 (O_324,N_14695,N_14805);
nand UO_325 (O_325,N_14673,N_14668);
nor UO_326 (O_326,N_14557,N_14506);
nor UO_327 (O_327,N_14735,N_14575);
nor UO_328 (O_328,N_14895,N_14996);
or UO_329 (O_329,N_14924,N_14636);
or UO_330 (O_330,N_14585,N_14867);
or UO_331 (O_331,N_14570,N_14565);
or UO_332 (O_332,N_14832,N_14994);
and UO_333 (O_333,N_14989,N_14960);
nand UO_334 (O_334,N_14650,N_14527);
or UO_335 (O_335,N_14590,N_14544);
and UO_336 (O_336,N_14905,N_14697);
or UO_337 (O_337,N_14502,N_14979);
and UO_338 (O_338,N_14806,N_14602);
or UO_339 (O_339,N_14730,N_14841);
nor UO_340 (O_340,N_14943,N_14632);
and UO_341 (O_341,N_14612,N_14660);
nor UO_342 (O_342,N_14771,N_14737);
and UO_343 (O_343,N_14509,N_14625);
and UO_344 (O_344,N_14914,N_14763);
or UO_345 (O_345,N_14523,N_14681);
xor UO_346 (O_346,N_14612,N_14780);
nand UO_347 (O_347,N_14600,N_14523);
nand UO_348 (O_348,N_14838,N_14671);
or UO_349 (O_349,N_14538,N_14955);
nor UO_350 (O_350,N_14911,N_14995);
nand UO_351 (O_351,N_14883,N_14729);
and UO_352 (O_352,N_14595,N_14659);
nor UO_353 (O_353,N_14940,N_14938);
nand UO_354 (O_354,N_14581,N_14990);
nor UO_355 (O_355,N_14839,N_14801);
xor UO_356 (O_356,N_14838,N_14831);
and UO_357 (O_357,N_14792,N_14510);
nor UO_358 (O_358,N_14699,N_14537);
or UO_359 (O_359,N_14834,N_14828);
and UO_360 (O_360,N_14546,N_14589);
and UO_361 (O_361,N_14957,N_14625);
or UO_362 (O_362,N_14981,N_14654);
or UO_363 (O_363,N_14548,N_14897);
nor UO_364 (O_364,N_14833,N_14756);
and UO_365 (O_365,N_14632,N_14797);
or UO_366 (O_366,N_14587,N_14698);
nand UO_367 (O_367,N_14820,N_14926);
or UO_368 (O_368,N_14985,N_14894);
or UO_369 (O_369,N_14888,N_14701);
nor UO_370 (O_370,N_14966,N_14720);
nor UO_371 (O_371,N_14853,N_14770);
or UO_372 (O_372,N_14641,N_14760);
or UO_373 (O_373,N_14939,N_14528);
xor UO_374 (O_374,N_14963,N_14782);
or UO_375 (O_375,N_14776,N_14802);
and UO_376 (O_376,N_14586,N_14509);
nand UO_377 (O_377,N_14854,N_14538);
and UO_378 (O_378,N_14948,N_14926);
nand UO_379 (O_379,N_14947,N_14687);
and UO_380 (O_380,N_14506,N_14838);
and UO_381 (O_381,N_14898,N_14640);
or UO_382 (O_382,N_14841,N_14722);
nor UO_383 (O_383,N_14575,N_14547);
or UO_384 (O_384,N_14892,N_14608);
and UO_385 (O_385,N_14779,N_14633);
nor UO_386 (O_386,N_14966,N_14527);
and UO_387 (O_387,N_14859,N_14860);
or UO_388 (O_388,N_14560,N_14593);
nand UO_389 (O_389,N_14656,N_14625);
nand UO_390 (O_390,N_14699,N_14875);
nand UO_391 (O_391,N_14651,N_14634);
or UO_392 (O_392,N_14565,N_14924);
or UO_393 (O_393,N_14974,N_14815);
and UO_394 (O_394,N_14775,N_14697);
xor UO_395 (O_395,N_14821,N_14736);
or UO_396 (O_396,N_14831,N_14657);
nor UO_397 (O_397,N_14641,N_14693);
and UO_398 (O_398,N_14960,N_14811);
nand UO_399 (O_399,N_14883,N_14573);
nor UO_400 (O_400,N_14650,N_14736);
nor UO_401 (O_401,N_14642,N_14992);
nand UO_402 (O_402,N_14824,N_14617);
nor UO_403 (O_403,N_14901,N_14729);
nand UO_404 (O_404,N_14854,N_14725);
nor UO_405 (O_405,N_14555,N_14771);
and UO_406 (O_406,N_14673,N_14701);
xnor UO_407 (O_407,N_14810,N_14672);
nand UO_408 (O_408,N_14941,N_14779);
or UO_409 (O_409,N_14842,N_14891);
or UO_410 (O_410,N_14883,N_14952);
nor UO_411 (O_411,N_14552,N_14542);
and UO_412 (O_412,N_14787,N_14797);
nor UO_413 (O_413,N_14951,N_14979);
nor UO_414 (O_414,N_14942,N_14789);
xnor UO_415 (O_415,N_14566,N_14698);
and UO_416 (O_416,N_14599,N_14676);
and UO_417 (O_417,N_14538,N_14992);
nand UO_418 (O_418,N_14811,N_14649);
nor UO_419 (O_419,N_14894,N_14683);
and UO_420 (O_420,N_14723,N_14702);
and UO_421 (O_421,N_14518,N_14719);
xnor UO_422 (O_422,N_14769,N_14979);
and UO_423 (O_423,N_14846,N_14988);
nand UO_424 (O_424,N_14854,N_14577);
nor UO_425 (O_425,N_14572,N_14993);
nor UO_426 (O_426,N_14597,N_14682);
nand UO_427 (O_427,N_14841,N_14859);
nand UO_428 (O_428,N_14924,N_14706);
and UO_429 (O_429,N_14563,N_14610);
nor UO_430 (O_430,N_14897,N_14573);
nand UO_431 (O_431,N_14869,N_14734);
or UO_432 (O_432,N_14501,N_14902);
or UO_433 (O_433,N_14515,N_14892);
and UO_434 (O_434,N_14554,N_14597);
nor UO_435 (O_435,N_14647,N_14674);
and UO_436 (O_436,N_14733,N_14681);
or UO_437 (O_437,N_14782,N_14991);
xnor UO_438 (O_438,N_14641,N_14898);
nand UO_439 (O_439,N_14525,N_14959);
or UO_440 (O_440,N_14756,N_14781);
xnor UO_441 (O_441,N_14828,N_14744);
nand UO_442 (O_442,N_14683,N_14993);
nor UO_443 (O_443,N_14944,N_14671);
nor UO_444 (O_444,N_14524,N_14741);
xnor UO_445 (O_445,N_14563,N_14815);
nand UO_446 (O_446,N_14968,N_14540);
xnor UO_447 (O_447,N_14917,N_14930);
and UO_448 (O_448,N_14570,N_14815);
xor UO_449 (O_449,N_14525,N_14884);
or UO_450 (O_450,N_14611,N_14982);
nor UO_451 (O_451,N_14806,N_14591);
and UO_452 (O_452,N_14555,N_14696);
or UO_453 (O_453,N_14577,N_14575);
and UO_454 (O_454,N_14804,N_14562);
and UO_455 (O_455,N_14591,N_14720);
or UO_456 (O_456,N_14560,N_14795);
and UO_457 (O_457,N_14998,N_14545);
nand UO_458 (O_458,N_14523,N_14532);
nor UO_459 (O_459,N_14778,N_14620);
nand UO_460 (O_460,N_14889,N_14939);
or UO_461 (O_461,N_14572,N_14904);
nor UO_462 (O_462,N_14547,N_14765);
and UO_463 (O_463,N_14511,N_14795);
and UO_464 (O_464,N_14909,N_14533);
nor UO_465 (O_465,N_14778,N_14808);
or UO_466 (O_466,N_14597,N_14852);
nand UO_467 (O_467,N_14575,N_14768);
xnor UO_468 (O_468,N_14812,N_14733);
or UO_469 (O_469,N_14701,N_14606);
or UO_470 (O_470,N_14891,N_14665);
or UO_471 (O_471,N_14754,N_14867);
or UO_472 (O_472,N_14621,N_14601);
nor UO_473 (O_473,N_14662,N_14512);
or UO_474 (O_474,N_14624,N_14662);
or UO_475 (O_475,N_14773,N_14923);
and UO_476 (O_476,N_14849,N_14809);
or UO_477 (O_477,N_14796,N_14819);
nor UO_478 (O_478,N_14740,N_14921);
or UO_479 (O_479,N_14845,N_14860);
nor UO_480 (O_480,N_14500,N_14992);
and UO_481 (O_481,N_14959,N_14989);
and UO_482 (O_482,N_14890,N_14793);
nand UO_483 (O_483,N_14604,N_14962);
or UO_484 (O_484,N_14945,N_14796);
and UO_485 (O_485,N_14979,N_14944);
and UO_486 (O_486,N_14588,N_14760);
or UO_487 (O_487,N_14916,N_14937);
or UO_488 (O_488,N_14902,N_14689);
xnor UO_489 (O_489,N_14746,N_14811);
nand UO_490 (O_490,N_14940,N_14951);
nor UO_491 (O_491,N_14843,N_14627);
nand UO_492 (O_492,N_14765,N_14744);
and UO_493 (O_493,N_14689,N_14722);
nor UO_494 (O_494,N_14752,N_14509);
nand UO_495 (O_495,N_14736,N_14993);
nand UO_496 (O_496,N_14581,N_14853);
or UO_497 (O_497,N_14605,N_14801);
nor UO_498 (O_498,N_14942,N_14534);
nor UO_499 (O_499,N_14700,N_14864);
or UO_500 (O_500,N_14971,N_14585);
nand UO_501 (O_501,N_14863,N_14998);
or UO_502 (O_502,N_14809,N_14576);
nand UO_503 (O_503,N_14520,N_14558);
nand UO_504 (O_504,N_14759,N_14623);
nor UO_505 (O_505,N_14690,N_14725);
xnor UO_506 (O_506,N_14706,N_14779);
nor UO_507 (O_507,N_14510,N_14973);
nor UO_508 (O_508,N_14941,N_14793);
or UO_509 (O_509,N_14927,N_14893);
nor UO_510 (O_510,N_14861,N_14940);
and UO_511 (O_511,N_14919,N_14907);
nor UO_512 (O_512,N_14676,N_14844);
nand UO_513 (O_513,N_14804,N_14723);
nor UO_514 (O_514,N_14853,N_14606);
or UO_515 (O_515,N_14639,N_14864);
nand UO_516 (O_516,N_14728,N_14506);
and UO_517 (O_517,N_14502,N_14908);
or UO_518 (O_518,N_14665,N_14858);
nand UO_519 (O_519,N_14692,N_14598);
and UO_520 (O_520,N_14794,N_14517);
nor UO_521 (O_521,N_14910,N_14821);
nor UO_522 (O_522,N_14779,N_14834);
and UO_523 (O_523,N_14984,N_14616);
nand UO_524 (O_524,N_14596,N_14900);
and UO_525 (O_525,N_14906,N_14736);
nor UO_526 (O_526,N_14618,N_14807);
nor UO_527 (O_527,N_14616,N_14848);
and UO_528 (O_528,N_14951,N_14528);
nor UO_529 (O_529,N_14554,N_14680);
or UO_530 (O_530,N_14889,N_14742);
nand UO_531 (O_531,N_14989,N_14791);
nand UO_532 (O_532,N_14538,N_14957);
and UO_533 (O_533,N_14746,N_14696);
nand UO_534 (O_534,N_14697,N_14853);
and UO_535 (O_535,N_14502,N_14781);
nand UO_536 (O_536,N_14702,N_14634);
nand UO_537 (O_537,N_14857,N_14721);
or UO_538 (O_538,N_14745,N_14993);
or UO_539 (O_539,N_14715,N_14852);
nor UO_540 (O_540,N_14827,N_14877);
nor UO_541 (O_541,N_14576,N_14734);
nand UO_542 (O_542,N_14908,N_14777);
or UO_543 (O_543,N_14763,N_14645);
nand UO_544 (O_544,N_14791,N_14803);
nor UO_545 (O_545,N_14514,N_14890);
nand UO_546 (O_546,N_14643,N_14512);
or UO_547 (O_547,N_14685,N_14963);
or UO_548 (O_548,N_14536,N_14952);
nand UO_549 (O_549,N_14511,N_14742);
or UO_550 (O_550,N_14804,N_14718);
nor UO_551 (O_551,N_14758,N_14734);
nand UO_552 (O_552,N_14888,N_14585);
and UO_553 (O_553,N_14821,N_14722);
and UO_554 (O_554,N_14537,N_14626);
nand UO_555 (O_555,N_14773,N_14593);
or UO_556 (O_556,N_14658,N_14522);
nand UO_557 (O_557,N_14699,N_14811);
nand UO_558 (O_558,N_14707,N_14722);
nor UO_559 (O_559,N_14675,N_14550);
or UO_560 (O_560,N_14738,N_14841);
and UO_561 (O_561,N_14865,N_14538);
nor UO_562 (O_562,N_14556,N_14525);
or UO_563 (O_563,N_14875,N_14649);
xor UO_564 (O_564,N_14781,N_14853);
nand UO_565 (O_565,N_14838,N_14686);
or UO_566 (O_566,N_14963,N_14505);
nand UO_567 (O_567,N_14980,N_14599);
or UO_568 (O_568,N_14894,N_14664);
nand UO_569 (O_569,N_14654,N_14751);
xnor UO_570 (O_570,N_14856,N_14882);
xnor UO_571 (O_571,N_14807,N_14949);
nand UO_572 (O_572,N_14580,N_14505);
nor UO_573 (O_573,N_14580,N_14991);
nand UO_574 (O_574,N_14500,N_14935);
and UO_575 (O_575,N_14720,N_14768);
or UO_576 (O_576,N_14644,N_14508);
nand UO_577 (O_577,N_14611,N_14899);
nor UO_578 (O_578,N_14623,N_14561);
and UO_579 (O_579,N_14545,N_14855);
xnor UO_580 (O_580,N_14757,N_14647);
nor UO_581 (O_581,N_14659,N_14975);
nor UO_582 (O_582,N_14708,N_14670);
or UO_583 (O_583,N_14961,N_14766);
nand UO_584 (O_584,N_14709,N_14631);
nand UO_585 (O_585,N_14502,N_14893);
and UO_586 (O_586,N_14624,N_14862);
and UO_587 (O_587,N_14694,N_14562);
or UO_588 (O_588,N_14921,N_14706);
and UO_589 (O_589,N_14655,N_14807);
xor UO_590 (O_590,N_14576,N_14631);
and UO_591 (O_591,N_14907,N_14779);
and UO_592 (O_592,N_14702,N_14986);
nor UO_593 (O_593,N_14778,N_14516);
and UO_594 (O_594,N_14997,N_14591);
nand UO_595 (O_595,N_14681,N_14626);
or UO_596 (O_596,N_14956,N_14835);
or UO_597 (O_597,N_14674,N_14628);
and UO_598 (O_598,N_14559,N_14573);
or UO_599 (O_599,N_14702,N_14925);
nor UO_600 (O_600,N_14839,N_14911);
and UO_601 (O_601,N_14909,N_14931);
or UO_602 (O_602,N_14749,N_14713);
or UO_603 (O_603,N_14834,N_14537);
or UO_604 (O_604,N_14581,N_14638);
or UO_605 (O_605,N_14633,N_14900);
xor UO_606 (O_606,N_14693,N_14982);
and UO_607 (O_607,N_14843,N_14538);
nand UO_608 (O_608,N_14828,N_14747);
nand UO_609 (O_609,N_14642,N_14750);
xnor UO_610 (O_610,N_14612,N_14609);
nand UO_611 (O_611,N_14735,N_14798);
nand UO_612 (O_612,N_14518,N_14997);
nor UO_613 (O_613,N_14889,N_14583);
nor UO_614 (O_614,N_14577,N_14524);
nor UO_615 (O_615,N_14785,N_14713);
nand UO_616 (O_616,N_14597,N_14774);
and UO_617 (O_617,N_14784,N_14569);
and UO_618 (O_618,N_14732,N_14849);
or UO_619 (O_619,N_14960,N_14687);
or UO_620 (O_620,N_14543,N_14823);
nor UO_621 (O_621,N_14882,N_14551);
or UO_622 (O_622,N_14532,N_14721);
and UO_623 (O_623,N_14744,N_14760);
nand UO_624 (O_624,N_14507,N_14865);
and UO_625 (O_625,N_14592,N_14625);
nor UO_626 (O_626,N_14766,N_14716);
nor UO_627 (O_627,N_14501,N_14825);
nand UO_628 (O_628,N_14712,N_14795);
and UO_629 (O_629,N_14780,N_14872);
or UO_630 (O_630,N_14902,N_14934);
xor UO_631 (O_631,N_14816,N_14789);
nand UO_632 (O_632,N_14825,N_14608);
and UO_633 (O_633,N_14958,N_14950);
and UO_634 (O_634,N_14537,N_14865);
or UO_635 (O_635,N_14869,N_14979);
and UO_636 (O_636,N_14783,N_14815);
or UO_637 (O_637,N_14884,N_14690);
nor UO_638 (O_638,N_14980,N_14883);
and UO_639 (O_639,N_14849,N_14785);
nor UO_640 (O_640,N_14508,N_14681);
nor UO_641 (O_641,N_14542,N_14672);
nand UO_642 (O_642,N_14939,N_14605);
nor UO_643 (O_643,N_14702,N_14913);
and UO_644 (O_644,N_14854,N_14829);
xor UO_645 (O_645,N_14596,N_14848);
xor UO_646 (O_646,N_14736,N_14863);
nor UO_647 (O_647,N_14713,N_14768);
xor UO_648 (O_648,N_14870,N_14533);
or UO_649 (O_649,N_14815,N_14674);
nand UO_650 (O_650,N_14722,N_14946);
nor UO_651 (O_651,N_14683,N_14939);
nand UO_652 (O_652,N_14611,N_14747);
nor UO_653 (O_653,N_14721,N_14544);
and UO_654 (O_654,N_14549,N_14756);
and UO_655 (O_655,N_14755,N_14567);
or UO_656 (O_656,N_14862,N_14782);
nand UO_657 (O_657,N_14553,N_14508);
nand UO_658 (O_658,N_14865,N_14994);
nand UO_659 (O_659,N_14640,N_14968);
and UO_660 (O_660,N_14507,N_14529);
and UO_661 (O_661,N_14593,N_14629);
or UO_662 (O_662,N_14700,N_14624);
or UO_663 (O_663,N_14579,N_14571);
nor UO_664 (O_664,N_14743,N_14573);
or UO_665 (O_665,N_14845,N_14713);
or UO_666 (O_666,N_14951,N_14821);
or UO_667 (O_667,N_14994,N_14757);
nand UO_668 (O_668,N_14706,N_14792);
and UO_669 (O_669,N_14569,N_14927);
nor UO_670 (O_670,N_14581,N_14718);
nor UO_671 (O_671,N_14610,N_14867);
and UO_672 (O_672,N_14779,N_14739);
and UO_673 (O_673,N_14695,N_14871);
nor UO_674 (O_674,N_14790,N_14604);
nand UO_675 (O_675,N_14533,N_14743);
nand UO_676 (O_676,N_14957,N_14767);
and UO_677 (O_677,N_14947,N_14869);
or UO_678 (O_678,N_14627,N_14964);
nor UO_679 (O_679,N_14604,N_14762);
nor UO_680 (O_680,N_14599,N_14743);
nor UO_681 (O_681,N_14550,N_14564);
or UO_682 (O_682,N_14596,N_14981);
or UO_683 (O_683,N_14876,N_14964);
or UO_684 (O_684,N_14502,N_14828);
and UO_685 (O_685,N_14977,N_14805);
nor UO_686 (O_686,N_14581,N_14547);
nand UO_687 (O_687,N_14581,N_14949);
or UO_688 (O_688,N_14586,N_14786);
nand UO_689 (O_689,N_14618,N_14597);
nand UO_690 (O_690,N_14818,N_14556);
nand UO_691 (O_691,N_14583,N_14671);
or UO_692 (O_692,N_14697,N_14759);
nor UO_693 (O_693,N_14865,N_14844);
nor UO_694 (O_694,N_14595,N_14712);
nor UO_695 (O_695,N_14614,N_14785);
and UO_696 (O_696,N_14981,N_14757);
xor UO_697 (O_697,N_14792,N_14650);
and UO_698 (O_698,N_14845,N_14706);
nor UO_699 (O_699,N_14846,N_14779);
and UO_700 (O_700,N_14993,N_14795);
nand UO_701 (O_701,N_14585,N_14690);
or UO_702 (O_702,N_14892,N_14546);
and UO_703 (O_703,N_14716,N_14506);
nor UO_704 (O_704,N_14803,N_14726);
nor UO_705 (O_705,N_14522,N_14921);
xnor UO_706 (O_706,N_14871,N_14955);
or UO_707 (O_707,N_14672,N_14613);
nor UO_708 (O_708,N_14953,N_14993);
nand UO_709 (O_709,N_14528,N_14918);
nand UO_710 (O_710,N_14634,N_14814);
nand UO_711 (O_711,N_14986,N_14625);
and UO_712 (O_712,N_14844,N_14905);
nor UO_713 (O_713,N_14651,N_14962);
and UO_714 (O_714,N_14509,N_14859);
and UO_715 (O_715,N_14755,N_14754);
or UO_716 (O_716,N_14868,N_14543);
nand UO_717 (O_717,N_14901,N_14968);
nand UO_718 (O_718,N_14925,N_14956);
nor UO_719 (O_719,N_14658,N_14906);
nand UO_720 (O_720,N_14615,N_14847);
nor UO_721 (O_721,N_14790,N_14640);
nand UO_722 (O_722,N_14961,N_14695);
nor UO_723 (O_723,N_14945,N_14562);
or UO_724 (O_724,N_14882,N_14736);
nand UO_725 (O_725,N_14512,N_14786);
nand UO_726 (O_726,N_14633,N_14989);
nor UO_727 (O_727,N_14571,N_14677);
or UO_728 (O_728,N_14550,N_14872);
nand UO_729 (O_729,N_14660,N_14680);
and UO_730 (O_730,N_14745,N_14519);
nand UO_731 (O_731,N_14727,N_14713);
and UO_732 (O_732,N_14568,N_14500);
nor UO_733 (O_733,N_14822,N_14800);
nand UO_734 (O_734,N_14860,N_14947);
or UO_735 (O_735,N_14562,N_14917);
or UO_736 (O_736,N_14925,N_14819);
nor UO_737 (O_737,N_14860,N_14513);
nor UO_738 (O_738,N_14850,N_14828);
nand UO_739 (O_739,N_14874,N_14899);
and UO_740 (O_740,N_14845,N_14905);
and UO_741 (O_741,N_14705,N_14870);
nand UO_742 (O_742,N_14581,N_14583);
nor UO_743 (O_743,N_14669,N_14858);
xor UO_744 (O_744,N_14654,N_14856);
xnor UO_745 (O_745,N_14942,N_14904);
or UO_746 (O_746,N_14766,N_14586);
nor UO_747 (O_747,N_14630,N_14516);
nand UO_748 (O_748,N_14550,N_14729);
or UO_749 (O_749,N_14620,N_14885);
nand UO_750 (O_750,N_14882,N_14946);
nand UO_751 (O_751,N_14531,N_14630);
nor UO_752 (O_752,N_14854,N_14793);
or UO_753 (O_753,N_14982,N_14767);
and UO_754 (O_754,N_14713,N_14669);
or UO_755 (O_755,N_14762,N_14711);
nor UO_756 (O_756,N_14509,N_14518);
nand UO_757 (O_757,N_14531,N_14667);
nand UO_758 (O_758,N_14792,N_14729);
or UO_759 (O_759,N_14654,N_14753);
or UO_760 (O_760,N_14955,N_14735);
and UO_761 (O_761,N_14997,N_14944);
or UO_762 (O_762,N_14782,N_14878);
and UO_763 (O_763,N_14957,N_14661);
xnor UO_764 (O_764,N_14705,N_14515);
nor UO_765 (O_765,N_14646,N_14819);
or UO_766 (O_766,N_14966,N_14993);
nor UO_767 (O_767,N_14503,N_14880);
nand UO_768 (O_768,N_14505,N_14885);
or UO_769 (O_769,N_14662,N_14866);
and UO_770 (O_770,N_14731,N_14840);
and UO_771 (O_771,N_14656,N_14770);
and UO_772 (O_772,N_14729,N_14659);
nor UO_773 (O_773,N_14706,N_14689);
nor UO_774 (O_774,N_14634,N_14868);
or UO_775 (O_775,N_14805,N_14978);
or UO_776 (O_776,N_14905,N_14583);
nor UO_777 (O_777,N_14712,N_14955);
or UO_778 (O_778,N_14889,N_14747);
nor UO_779 (O_779,N_14985,N_14594);
and UO_780 (O_780,N_14953,N_14871);
or UO_781 (O_781,N_14502,N_14820);
and UO_782 (O_782,N_14631,N_14579);
or UO_783 (O_783,N_14718,N_14522);
and UO_784 (O_784,N_14826,N_14924);
and UO_785 (O_785,N_14698,N_14721);
nor UO_786 (O_786,N_14668,N_14940);
and UO_787 (O_787,N_14773,N_14772);
xor UO_788 (O_788,N_14832,N_14806);
xnor UO_789 (O_789,N_14765,N_14649);
nand UO_790 (O_790,N_14645,N_14626);
nand UO_791 (O_791,N_14886,N_14887);
nor UO_792 (O_792,N_14709,N_14909);
xor UO_793 (O_793,N_14639,N_14804);
or UO_794 (O_794,N_14665,N_14678);
nor UO_795 (O_795,N_14800,N_14611);
and UO_796 (O_796,N_14929,N_14908);
nor UO_797 (O_797,N_14718,N_14704);
nand UO_798 (O_798,N_14628,N_14939);
nand UO_799 (O_799,N_14856,N_14556);
nand UO_800 (O_800,N_14519,N_14991);
nand UO_801 (O_801,N_14960,N_14958);
or UO_802 (O_802,N_14999,N_14817);
and UO_803 (O_803,N_14573,N_14742);
nand UO_804 (O_804,N_14737,N_14526);
or UO_805 (O_805,N_14558,N_14603);
or UO_806 (O_806,N_14940,N_14698);
and UO_807 (O_807,N_14637,N_14515);
nor UO_808 (O_808,N_14506,N_14614);
or UO_809 (O_809,N_14675,N_14898);
nand UO_810 (O_810,N_14573,N_14920);
nand UO_811 (O_811,N_14986,N_14739);
and UO_812 (O_812,N_14764,N_14885);
or UO_813 (O_813,N_14767,N_14748);
nor UO_814 (O_814,N_14731,N_14991);
nor UO_815 (O_815,N_14732,N_14682);
or UO_816 (O_816,N_14548,N_14604);
nor UO_817 (O_817,N_14560,N_14837);
or UO_818 (O_818,N_14811,N_14619);
and UO_819 (O_819,N_14999,N_14570);
or UO_820 (O_820,N_14860,N_14626);
nor UO_821 (O_821,N_14794,N_14583);
or UO_822 (O_822,N_14988,N_14749);
xor UO_823 (O_823,N_14963,N_14858);
nor UO_824 (O_824,N_14597,N_14879);
xnor UO_825 (O_825,N_14773,N_14679);
nor UO_826 (O_826,N_14656,N_14520);
nor UO_827 (O_827,N_14500,N_14991);
and UO_828 (O_828,N_14558,N_14687);
or UO_829 (O_829,N_14940,N_14706);
nor UO_830 (O_830,N_14967,N_14911);
nor UO_831 (O_831,N_14570,N_14743);
and UO_832 (O_832,N_14591,N_14908);
or UO_833 (O_833,N_14803,N_14903);
xnor UO_834 (O_834,N_14733,N_14575);
and UO_835 (O_835,N_14729,N_14705);
nor UO_836 (O_836,N_14641,N_14721);
nand UO_837 (O_837,N_14824,N_14637);
nand UO_838 (O_838,N_14928,N_14667);
xor UO_839 (O_839,N_14568,N_14875);
or UO_840 (O_840,N_14656,N_14569);
xnor UO_841 (O_841,N_14801,N_14508);
and UO_842 (O_842,N_14651,N_14501);
nand UO_843 (O_843,N_14702,N_14627);
or UO_844 (O_844,N_14500,N_14704);
nand UO_845 (O_845,N_14762,N_14958);
or UO_846 (O_846,N_14769,N_14906);
xnor UO_847 (O_847,N_14745,N_14513);
and UO_848 (O_848,N_14940,N_14887);
nor UO_849 (O_849,N_14943,N_14604);
or UO_850 (O_850,N_14970,N_14520);
or UO_851 (O_851,N_14834,N_14879);
or UO_852 (O_852,N_14932,N_14679);
nand UO_853 (O_853,N_14825,N_14588);
or UO_854 (O_854,N_14786,N_14632);
and UO_855 (O_855,N_14541,N_14590);
nand UO_856 (O_856,N_14643,N_14562);
nor UO_857 (O_857,N_14786,N_14894);
nor UO_858 (O_858,N_14522,N_14894);
nor UO_859 (O_859,N_14513,N_14934);
nor UO_860 (O_860,N_14852,N_14573);
and UO_861 (O_861,N_14926,N_14662);
and UO_862 (O_862,N_14897,N_14880);
and UO_863 (O_863,N_14578,N_14696);
and UO_864 (O_864,N_14614,N_14560);
xnor UO_865 (O_865,N_14935,N_14708);
xor UO_866 (O_866,N_14503,N_14878);
and UO_867 (O_867,N_14640,N_14508);
or UO_868 (O_868,N_14955,N_14976);
and UO_869 (O_869,N_14777,N_14743);
or UO_870 (O_870,N_14724,N_14654);
and UO_871 (O_871,N_14760,N_14770);
or UO_872 (O_872,N_14604,N_14858);
nand UO_873 (O_873,N_14594,N_14629);
or UO_874 (O_874,N_14989,N_14679);
nor UO_875 (O_875,N_14524,N_14880);
nor UO_876 (O_876,N_14729,N_14700);
nand UO_877 (O_877,N_14583,N_14691);
or UO_878 (O_878,N_14902,N_14929);
nand UO_879 (O_879,N_14775,N_14611);
and UO_880 (O_880,N_14642,N_14933);
and UO_881 (O_881,N_14737,N_14873);
and UO_882 (O_882,N_14504,N_14597);
and UO_883 (O_883,N_14861,N_14961);
and UO_884 (O_884,N_14899,N_14620);
and UO_885 (O_885,N_14960,N_14777);
and UO_886 (O_886,N_14847,N_14591);
nand UO_887 (O_887,N_14994,N_14720);
or UO_888 (O_888,N_14718,N_14606);
nor UO_889 (O_889,N_14925,N_14699);
nor UO_890 (O_890,N_14936,N_14901);
nor UO_891 (O_891,N_14508,N_14945);
or UO_892 (O_892,N_14654,N_14836);
nor UO_893 (O_893,N_14810,N_14905);
xor UO_894 (O_894,N_14789,N_14985);
nor UO_895 (O_895,N_14830,N_14826);
nor UO_896 (O_896,N_14871,N_14599);
and UO_897 (O_897,N_14982,N_14973);
nand UO_898 (O_898,N_14799,N_14769);
or UO_899 (O_899,N_14594,N_14615);
or UO_900 (O_900,N_14527,N_14693);
xnor UO_901 (O_901,N_14841,N_14520);
nor UO_902 (O_902,N_14814,N_14877);
xor UO_903 (O_903,N_14675,N_14531);
and UO_904 (O_904,N_14720,N_14767);
xor UO_905 (O_905,N_14783,N_14862);
nand UO_906 (O_906,N_14649,N_14778);
nor UO_907 (O_907,N_14631,N_14922);
nand UO_908 (O_908,N_14973,N_14552);
or UO_909 (O_909,N_14613,N_14994);
nor UO_910 (O_910,N_14762,N_14890);
nor UO_911 (O_911,N_14618,N_14988);
and UO_912 (O_912,N_14538,N_14904);
nor UO_913 (O_913,N_14925,N_14831);
or UO_914 (O_914,N_14783,N_14585);
nand UO_915 (O_915,N_14561,N_14742);
xnor UO_916 (O_916,N_14840,N_14733);
and UO_917 (O_917,N_14740,N_14747);
nand UO_918 (O_918,N_14663,N_14701);
and UO_919 (O_919,N_14589,N_14559);
nor UO_920 (O_920,N_14831,N_14658);
or UO_921 (O_921,N_14884,N_14769);
nor UO_922 (O_922,N_14620,N_14965);
nand UO_923 (O_923,N_14783,N_14800);
nor UO_924 (O_924,N_14850,N_14873);
nand UO_925 (O_925,N_14786,N_14950);
nor UO_926 (O_926,N_14988,N_14831);
and UO_927 (O_927,N_14807,N_14895);
and UO_928 (O_928,N_14682,N_14581);
and UO_929 (O_929,N_14733,N_14724);
nor UO_930 (O_930,N_14639,N_14847);
and UO_931 (O_931,N_14889,N_14946);
nor UO_932 (O_932,N_14820,N_14675);
or UO_933 (O_933,N_14887,N_14872);
xnor UO_934 (O_934,N_14860,N_14812);
and UO_935 (O_935,N_14575,N_14874);
nand UO_936 (O_936,N_14628,N_14905);
nor UO_937 (O_937,N_14546,N_14913);
nor UO_938 (O_938,N_14736,N_14572);
and UO_939 (O_939,N_14876,N_14959);
or UO_940 (O_940,N_14783,N_14829);
nor UO_941 (O_941,N_14658,N_14824);
and UO_942 (O_942,N_14582,N_14693);
and UO_943 (O_943,N_14722,N_14512);
nor UO_944 (O_944,N_14508,N_14630);
or UO_945 (O_945,N_14624,N_14884);
or UO_946 (O_946,N_14847,N_14976);
nor UO_947 (O_947,N_14974,N_14518);
xor UO_948 (O_948,N_14593,N_14927);
and UO_949 (O_949,N_14889,N_14709);
xnor UO_950 (O_950,N_14926,N_14866);
and UO_951 (O_951,N_14801,N_14726);
nand UO_952 (O_952,N_14781,N_14772);
and UO_953 (O_953,N_14725,N_14735);
xnor UO_954 (O_954,N_14629,N_14841);
or UO_955 (O_955,N_14536,N_14641);
nor UO_956 (O_956,N_14931,N_14531);
nor UO_957 (O_957,N_14859,N_14602);
and UO_958 (O_958,N_14505,N_14513);
nor UO_959 (O_959,N_14572,N_14590);
nand UO_960 (O_960,N_14819,N_14745);
or UO_961 (O_961,N_14964,N_14777);
and UO_962 (O_962,N_14549,N_14985);
xor UO_963 (O_963,N_14626,N_14648);
and UO_964 (O_964,N_14913,N_14631);
nand UO_965 (O_965,N_14553,N_14684);
nand UO_966 (O_966,N_14533,N_14898);
nand UO_967 (O_967,N_14814,N_14503);
nand UO_968 (O_968,N_14737,N_14606);
or UO_969 (O_969,N_14688,N_14542);
nand UO_970 (O_970,N_14659,N_14660);
or UO_971 (O_971,N_14582,N_14689);
and UO_972 (O_972,N_14646,N_14526);
nand UO_973 (O_973,N_14929,N_14717);
or UO_974 (O_974,N_14900,N_14871);
or UO_975 (O_975,N_14933,N_14671);
or UO_976 (O_976,N_14974,N_14674);
nand UO_977 (O_977,N_14607,N_14910);
and UO_978 (O_978,N_14730,N_14540);
nand UO_979 (O_979,N_14924,N_14524);
nor UO_980 (O_980,N_14556,N_14577);
nor UO_981 (O_981,N_14932,N_14738);
xor UO_982 (O_982,N_14540,N_14639);
nor UO_983 (O_983,N_14510,N_14743);
nand UO_984 (O_984,N_14647,N_14848);
nand UO_985 (O_985,N_14827,N_14529);
nand UO_986 (O_986,N_14763,N_14612);
nor UO_987 (O_987,N_14942,N_14877);
nor UO_988 (O_988,N_14995,N_14913);
or UO_989 (O_989,N_14789,N_14573);
and UO_990 (O_990,N_14990,N_14707);
xnor UO_991 (O_991,N_14790,N_14703);
nor UO_992 (O_992,N_14667,N_14584);
nor UO_993 (O_993,N_14692,N_14915);
or UO_994 (O_994,N_14971,N_14617);
nand UO_995 (O_995,N_14968,N_14910);
xnor UO_996 (O_996,N_14608,N_14613);
xor UO_997 (O_997,N_14695,N_14521);
nand UO_998 (O_998,N_14539,N_14715);
and UO_999 (O_999,N_14663,N_14906);
nor UO_1000 (O_1000,N_14516,N_14685);
nand UO_1001 (O_1001,N_14590,N_14962);
nor UO_1002 (O_1002,N_14729,N_14626);
and UO_1003 (O_1003,N_14963,N_14661);
xnor UO_1004 (O_1004,N_14743,N_14553);
nor UO_1005 (O_1005,N_14904,N_14836);
xor UO_1006 (O_1006,N_14988,N_14628);
nor UO_1007 (O_1007,N_14861,N_14923);
and UO_1008 (O_1008,N_14891,N_14732);
nor UO_1009 (O_1009,N_14978,N_14514);
xnor UO_1010 (O_1010,N_14523,N_14783);
or UO_1011 (O_1011,N_14528,N_14750);
xnor UO_1012 (O_1012,N_14658,N_14640);
or UO_1013 (O_1013,N_14504,N_14601);
nor UO_1014 (O_1014,N_14899,N_14733);
and UO_1015 (O_1015,N_14839,N_14546);
nor UO_1016 (O_1016,N_14882,N_14511);
nor UO_1017 (O_1017,N_14957,N_14798);
or UO_1018 (O_1018,N_14507,N_14546);
xor UO_1019 (O_1019,N_14552,N_14632);
and UO_1020 (O_1020,N_14512,N_14590);
or UO_1021 (O_1021,N_14617,N_14697);
nand UO_1022 (O_1022,N_14773,N_14967);
and UO_1023 (O_1023,N_14982,N_14838);
xnor UO_1024 (O_1024,N_14710,N_14852);
and UO_1025 (O_1025,N_14717,N_14831);
nand UO_1026 (O_1026,N_14821,N_14964);
nand UO_1027 (O_1027,N_14835,N_14529);
or UO_1028 (O_1028,N_14516,N_14613);
nand UO_1029 (O_1029,N_14579,N_14806);
nand UO_1030 (O_1030,N_14896,N_14898);
or UO_1031 (O_1031,N_14944,N_14824);
nand UO_1032 (O_1032,N_14824,N_14888);
nor UO_1033 (O_1033,N_14646,N_14975);
nor UO_1034 (O_1034,N_14701,N_14855);
nand UO_1035 (O_1035,N_14720,N_14946);
nor UO_1036 (O_1036,N_14934,N_14667);
or UO_1037 (O_1037,N_14578,N_14672);
nor UO_1038 (O_1038,N_14776,N_14562);
and UO_1039 (O_1039,N_14896,N_14970);
and UO_1040 (O_1040,N_14759,N_14799);
or UO_1041 (O_1041,N_14937,N_14902);
nor UO_1042 (O_1042,N_14671,N_14629);
or UO_1043 (O_1043,N_14672,N_14761);
and UO_1044 (O_1044,N_14737,N_14746);
or UO_1045 (O_1045,N_14504,N_14916);
nor UO_1046 (O_1046,N_14959,N_14925);
nand UO_1047 (O_1047,N_14679,N_14711);
or UO_1048 (O_1048,N_14613,N_14769);
nor UO_1049 (O_1049,N_14611,N_14765);
nand UO_1050 (O_1050,N_14613,N_14588);
or UO_1051 (O_1051,N_14788,N_14754);
nor UO_1052 (O_1052,N_14761,N_14889);
nand UO_1053 (O_1053,N_14689,N_14799);
and UO_1054 (O_1054,N_14866,N_14881);
nand UO_1055 (O_1055,N_14987,N_14554);
and UO_1056 (O_1056,N_14628,N_14775);
and UO_1057 (O_1057,N_14918,N_14585);
or UO_1058 (O_1058,N_14507,N_14750);
xnor UO_1059 (O_1059,N_14901,N_14569);
and UO_1060 (O_1060,N_14980,N_14802);
and UO_1061 (O_1061,N_14958,N_14857);
or UO_1062 (O_1062,N_14790,N_14874);
xnor UO_1063 (O_1063,N_14731,N_14628);
nor UO_1064 (O_1064,N_14573,N_14701);
and UO_1065 (O_1065,N_14718,N_14791);
and UO_1066 (O_1066,N_14906,N_14775);
nand UO_1067 (O_1067,N_14655,N_14833);
xnor UO_1068 (O_1068,N_14859,N_14818);
nor UO_1069 (O_1069,N_14646,N_14970);
xor UO_1070 (O_1070,N_14716,N_14697);
and UO_1071 (O_1071,N_14900,N_14775);
nand UO_1072 (O_1072,N_14737,N_14508);
or UO_1073 (O_1073,N_14715,N_14557);
nand UO_1074 (O_1074,N_14907,N_14810);
and UO_1075 (O_1075,N_14550,N_14503);
or UO_1076 (O_1076,N_14574,N_14739);
and UO_1077 (O_1077,N_14966,N_14758);
nand UO_1078 (O_1078,N_14543,N_14676);
or UO_1079 (O_1079,N_14510,N_14824);
and UO_1080 (O_1080,N_14964,N_14678);
nor UO_1081 (O_1081,N_14673,N_14796);
xnor UO_1082 (O_1082,N_14663,N_14870);
or UO_1083 (O_1083,N_14622,N_14778);
nand UO_1084 (O_1084,N_14987,N_14786);
nand UO_1085 (O_1085,N_14701,N_14605);
and UO_1086 (O_1086,N_14801,N_14678);
xor UO_1087 (O_1087,N_14991,N_14760);
nand UO_1088 (O_1088,N_14681,N_14787);
xor UO_1089 (O_1089,N_14931,N_14969);
and UO_1090 (O_1090,N_14547,N_14939);
nor UO_1091 (O_1091,N_14763,N_14704);
nand UO_1092 (O_1092,N_14598,N_14800);
nor UO_1093 (O_1093,N_14876,N_14801);
or UO_1094 (O_1094,N_14877,N_14903);
nor UO_1095 (O_1095,N_14716,N_14966);
xnor UO_1096 (O_1096,N_14980,N_14784);
or UO_1097 (O_1097,N_14553,N_14753);
nor UO_1098 (O_1098,N_14735,N_14967);
or UO_1099 (O_1099,N_14658,N_14759);
and UO_1100 (O_1100,N_14885,N_14859);
or UO_1101 (O_1101,N_14591,N_14653);
or UO_1102 (O_1102,N_14667,N_14856);
or UO_1103 (O_1103,N_14931,N_14634);
or UO_1104 (O_1104,N_14711,N_14678);
or UO_1105 (O_1105,N_14560,N_14836);
and UO_1106 (O_1106,N_14790,N_14670);
or UO_1107 (O_1107,N_14562,N_14752);
xor UO_1108 (O_1108,N_14894,N_14902);
xnor UO_1109 (O_1109,N_14707,N_14564);
nand UO_1110 (O_1110,N_14956,N_14562);
or UO_1111 (O_1111,N_14747,N_14703);
or UO_1112 (O_1112,N_14860,N_14761);
xnor UO_1113 (O_1113,N_14664,N_14572);
nor UO_1114 (O_1114,N_14867,N_14547);
nor UO_1115 (O_1115,N_14629,N_14728);
xnor UO_1116 (O_1116,N_14527,N_14613);
and UO_1117 (O_1117,N_14970,N_14895);
nor UO_1118 (O_1118,N_14946,N_14552);
or UO_1119 (O_1119,N_14707,N_14690);
nor UO_1120 (O_1120,N_14761,N_14713);
xnor UO_1121 (O_1121,N_14836,N_14890);
nor UO_1122 (O_1122,N_14567,N_14787);
nor UO_1123 (O_1123,N_14914,N_14907);
or UO_1124 (O_1124,N_14571,N_14520);
and UO_1125 (O_1125,N_14609,N_14703);
or UO_1126 (O_1126,N_14507,N_14861);
and UO_1127 (O_1127,N_14754,N_14542);
and UO_1128 (O_1128,N_14552,N_14660);
nor UO_1129 (O_1129,N_14526,N_14864);
and UO_1130 (O_1130,N_14802,N_14544);
and UO_1131 (O_1131,N_14924,N_14946);
nor UO_1132 (O_1132,N_14836,N_14983);
xnor UO_1133 (O_1133,N_14791,N_14682);
nor UO_1134 (O_1134,N_14697,N_14890);
or UO_1135 (O_1135,N_14765,N_14978);
nand UO_1136 (O_1136,N_14932,N_14594);
nor UO_1137 (O_1137,N_14927,N_14745);
xnor UO_1138 (O_1138,N_14503,N_14668);
nand UO_1139 (O_1139,N_14702,N_14930);
and UO_1140 (O_1140,N_14762,N_14788);
nor UO_1141 (O_1141,N_14944,N_14846);
nand UO_1142 (O_1142,N_14692,N_14863);
nand UO_1143 (O_1143,N_14547,N_14549);
nand UO_1144 (O_1144,N_14605,N_14702);
or UO_1145 (O_1145,N_14613,N_14637);
or UO_1146 (O_1146,N_14894,N_14912);
nand UO_1147 (O_1147,N_14853,N_14562);
nor UO_1148 (O_1148,N_14514,N_14982);
or UO_1149 (O_1149,N_14772,N_14883);
nand UO_1150 (O_1150,N_14624,N_14739);
xor UO_1151 (O_1151,N_14992,N_14662);
nand UO_1152 (O_1152,N_14667,N_14648);
nand UO_1153 (O_1153,N_14858,N_14629);
and UO_1154 (O_1154,N_14536,N_14587);
xor UO_1155 (O_1155,N_14786,N_14610);
nor UO_1156 (O_1156,N_14985,N_14739);
nand UO_1157 (O_1157,N_14746,N_14871);
or UO_1158 (O_1158,N_14697,N_14544);
or UO_1159 (O_1159,N_14712,N_14777);
or UO_1160 (O_1160,N_14726,N_14842);
and UO_1161 (O_1161,N_14885,N_14820);
and UO_1162 (O_1162,N_14535,N_14763);
nand UO_1163 (O_1163,N_14557,N_14695);
and UO_1164 (O_1164,N_14950,N_14994);
nor UO_1165 (O_1165,N_14655,N_14749);
nor UO_1166 (O_1166,N_14912,N_14733);
or UO_1167 (O_1167,N_14537,N_14978);
or UO_1168 (O_1168,N_14845,N_14510);
nand UO_1169 (O_1169,N_14748,N_14566);
and UO_1170 (O_1170,N_14633,N_14797);
nor UO_1171 (O_1171,N_14994,N_14546);
or UO_1172 (O_1172,N_14865,N_14799);
and UO_1173 (O_1173,N_14649,N_14648);
nor UO_1174 (O_1174,N_14678,N_14754);
or UO_1175 (O_1175,N_14685,N_14700);
xor UO_1176 (O_1176,N_14899,N_14635);
xnor UO_1177 (O_1177,N_14596,N_14859);
and UO_1178 (O_1178,N_14966,N_14784);
nand UO_1179 (O_1179,N_14554,N_14960);
and UO_1180 (O_1180,N_14760,N_14913);
nand UO_1181 (O_1181,N_14583,N_14760);
nand UO_1182 (O_1182,N_14690,N_14513);
xor UO_1183 (O_1183,N_14811,N_14934);
nor UO_1184 (O_1184,N_14844,N_14621);
or UO_1185 (O_1185,N_14686,N_14989);
nand UO_1186 (O_1186,N_14985,N_14625);
and UO_1187 (O_1187,N_14640,N_14964);
or UO_1188 (O_1188,N_14855,N_14900);
xor UO_1189 (O_1189,N_14770,N_14962);
or UO_1190 (O_1190,N_14781,N_14553);
nor UO_1191 (O_1191,N_14657,N_14820);
and UO_1192 (O_1192,N_14938,N_14671);
nand UO_1193 (O_1193,N_14597,N_14941);
nand UO_1194 (O_1194,N_14680,N_14563);
and UO_1195 (O_1195,N_14870,N_14602);
and UO_1196 (O_1196,N_14647,N_14569);
and UO_1197 (O_1197,N_14860,N_14710);
and UO_1198 (O_1198,N_14624,N_14973);
and UO_1199 (O_1199,N_14858,N_14803);
and UO_1200 (O_1200,N_14528,N_14636);
or UO_1201 (O_1201,N_14977,N_14774);
and UO_1202 (O_1202,N_14841,N_14857);
nor UO_1203 (O_1203,N_14891,N_14817);
and UO_1204 (O_1204,N_14827,N_14584);
nand UO_1205 (O_1205,N_14855,N_14772);
or UO_1206 (O_1206,N_14819,N_14668);
nand UO_1207 (O_1207,N_14970,N_14524);
nor UO_1208 (O_1208,N_14649,N_14976);
nand UO_1209 (O_1209,N_14627,N_14800);
nor UO_1210 (O_1210,N_14767,N_14785);
and UO_1211 (O_1211,N_14504,N_14996);
or UO_1212 (O_1212,N_14763,N_14863);
nor UO_1213 (O_1213,N_14981,N_14868);
nor UO_1214 (O_1214,N_14515,N_14944);
nand UO_1215 (O_1215,N_14766,N_14660);
nor UO_1216 (O_1216,N_14759,N_14890);
nor UO_1217 (O_1217,N_14849,N_14675);
xnor UO_1218 (O_1218,N_14941,N_14828);
or UO_1219 (O_1219,N_14621,N_14707);
xnor UO_1220 (O_1220,N_14523,N_14516);
or UO_1221 (O_1221,N_14567,N_14783);
nor UO_1222 (O_1222,N_14640,N_14780);
or UO_1223 (O_1223,N_14888,N_14948);
and UO_1224 (O_1224,N_14991,N_14567);
and UO_1225 (O_1225,N_14807,N_14566);
and UO_1226 (O_1226,N_14885,N_14627);
nor UO_1227 (O_1227,N_14532,N_14992);
nand UO_1228 (O_1228,N_14979,N_14683);
xnor UO_1229 (O_1229,N_14640,N_14715);
nor UO_1230 (O_1230,N_14825,N_14516);
nand UO_1231 (O_1231,N_14987,N_14760);
nand UO_1232 (O_1232,N_14638,N_14556);
xnor UO_1233 (O_1233,N_14984,N_14503);
nand UO_1234 (O_1234,N_14565,N_14956);
nor UO_1235 (O_1235,N_14546,N_14992);
nand UO_1236 (O_1236,N_14858,N_14608);
nor UO_1237 (O_1237,N_14952,N_14564);
nand UO_1238 (O_1238,N_14573,N_14783);
nand UO_1239 (O_1239,N_14854,N_14877);
and UO_1240 (O_1240,N_14563,N_14988);
and UO_1241 (O_1241,N_14766,N_14691);
nor UO_1242 (O_1242,N_14784,N_14525);
nor UO_1243 (O_1243,N_14823,N_14645);
xor UO_1244 (O_1244,N_14789,N_14943);
and UO_1245 (O_1245,N_14564,N_14570);
or UO_1246 (O_1246,N_14979,N_14689);
and UO_1247 (O_1247,N_14529,N_14658);
nor UO_1248 (O_1248,N_14902,N_14652);
and UO_1249 (O_1249,N_14737,N_14949);
and UO_1250 (O_1250,N_14732,N_14827);
or UO_1251 (O_1251,N_14838,N_14833);
or UO_1252 (O_1252,N_14544,N_14727);
and UO_1253 (O_1253,N_14781,N_14523);
or UO_1254 (O_1254,N_14770,N_14532);
nand UO_1255 (O_1255,N_14677,N_14990);
nor UO_1256 (O_1256,N_14615,N_14757);
nand UO_1257 (O_1257,N_14883,N_14984);
or UO_1258 (O_1258,N_14533,N_14777);
or UO_1259 (O_1259,N_14657,N_14760);
nor UO_1260 (O_1260,N_14930,N_14608);
and UO_1261 (O_1261,N_14702,N_14696);
and UO_1262 (O_1262,N_14559,N_14722);
or UO_1263 (O_1263,N_14950,N_14723);
nor UO_1264 (O_1264,N_14692,N_14727);
nor UO_1265 (O_1265,N_14643,N_14642);
nor UO_1266 (O_1266,N_14728,N_14582);
nand UO_1267 (O_1267,N_14644,N_14557);
nand UO_1268 (O_1268,N_14781,N_14876);
or UO_1269 (O_1269,N_14804,N_14563);
nor UO_1270 (O_1270,N_14724,N_14754);
nor UO_1271 (O_1271,N_14611,N_14695);
nand UO_1272 (O_1272,N_14581,N_14914);
nand UO_1273 (O_1273,N_14711,N_14836);
and UO_1274 (O_1274,N_14859,N_14918);
and UO_1275 (O_1275,N_14820,N_14615);
or UO_1276 (O_1276,N_14994,N_14812);
nand UO_1277 (O_1277,N_14865,N_14944);
or UO_1278 (O_1278,N_14952,N_14834);
and UO_1279 (O_1279,N_14552,N_14943);
nand UO_1280 (O_1280,N_14829,N_14579);
or UO_1281 (O_1281,N_14966,N_14765);
and UO_1282 (O_1282,N_14643,N_14606);
nand UO_1283 (O_1283,N_14991,N_14622);
nor UO_1284 (O_1284,N_14762,N_14575);
and UO_1285 (O_1285,N_14772,N_14666);
nor UO_1286 (O_1286,N_14535,N_14985);
nand UO_1287 (O_1287,N_14585,N_14654);
and UO_1288 (O_1288,N_14981,N_14966);
xor UO_1289 (O_1289,N_14946,N_14810);
xor UO_1290 (O_1290,N_14753,N_14762);
nor UO_1291 (O_1291,N_14800,N_14649);
xnor UO_1292 (O_1292,N_14871,N_14751);
xor UO_1293 (O_1293,N_14882,N_14827);
or UO_1294 (O_1294,N_14655,N_14999);
nor UO_1295 (O_1295,N_14917,N_14851);
nand UO_1296 (O_1296,N_14973,N_14579);
nand UO_1297 (O_1297,N_14687,N_14714);
xor UO_1298 (O_1298,N_14854,N_14875);
nand UO_1299 (O_1299,N_14775,N_14670);
nand UO_1300 (O_1300,N_14907,N_14507);
nor UO_1301 (O_1301,N_14694,N_14779);
or UO_1302 (O_1302,N_14609,N_14916);
or UO_1303 (O_1303,N_14675,N_14580);
nand UO_1304 (O_1304,N_14542,N_14867);
and UO_1305 (O_1305,N_14977,N_14794);
or UO_1306 (O_1306,N_14739,N_14725);
and UO_1307 (O_1307,N_14559,N_14583);
nand UO_1308 (O_1308,N_14877,N_14799);
and UO_1309 (O_1309,N_14673,N_14941);
nand UO_1310 (O_1310,N_14951,N_14628);
xor UO_1311 (O_1311,N_14656,N_14579);
and UO_1312 (O_1312,N_14546,N_14965);
nor UO_1313 (O_1313,N_14745,N_14952);
or UO_1314 (O_1314,N_14935,N_14644);
nor UO_1315 (O_1315,N_14973,N_14896);
and UO_1316 (O_1316,N_14624,N_14571);
xnor UO_1317 (O_1317,N_14540,N_14566);
or UO_1318 (O_1318,N_14824,N_14585);
and UO_1319 (O_1319,N_14501,N_14900);
nor UO_1320 (O_1320,N_14550,N_14598);
and UO_1321 (O_1321,N_14872,N_14906);
nor UO_1322 (O_1322,N_14619,N_14724);
nand UO_1323 (O_1323,N_14940,N_14834);
and UO_1324 (O_1324,N_14860,N_14543);
and UO_1325 (O_1325,N_14623,N_14766);
nand UO_1326 (O_1326,N_14693,N_14674);
and UO_1327 (O_1327,N_14648,N_14548);
nor UO_1328 (O_1328,N_14552,N_14905);
nor UO_1329 (O_1329,N_14850,N_14816);
nand UO_1330 (O_1330,N_14830,N_14808);
or UO_1331 (O_1331,N_14854,N_14988);
or UO_1332 (O_1332,N_14503,N_14829);
or UO_1333 (O_1333,N_14799,N_14530);
nand UO_1334 (O_1334,N_14500,N_14680);
nor UO_1335 (O_1335,N_14757,N_14747);
nand UO_1336 (O_1336,N_14825,N_14824);
or UO_1337 (O_1337,N_14643,N_14760);
nor UO_1338 (O_1338,N_14997,N_14515);
or UO_1339 (O_1339,N_14953,N_14639);
nand UO_1340 (O_1340,N_14583,N_14899);
nor UO_1341 (O_1341,N_14671,N_14678);
and UO_1342 (O_1342,N_14570,N_14588);
nor UO_1343 (O_1343,N_14524,N_14910);
or UO_1344 (O_1344,N_14697,N_14766);
nand UO_1345 (O_1345,N_14717,N_14915);
nand UO_1346 (O_1346,N_14836,N_14575);
or UO_1347 (O_1347,N_14836,N_14720);
nor UO_1348 (O_1348,N_14880,N_14952);
nand UO_1349 (O_1349,N_14766,N_14977);
nand UO_1350 (O_1350,N_14789,N_14649);
nor UO_1351 (O_1351,N_14849,N_14993);
and UO_1352 (O_1352,N_14617,N_14865);
and UO_1353 (O_1353,N_14821,N_14529);
and UO_1354 (O_1354,N_14759,N_14780);
xnor UO_1355 (O_1355,N_14645,N_14859);
and UO_1356 (O_1356,N_14941,N_14711);
nor UO_1357 (O_1357,N_14730,N_14630);
or UO_1358 (O_1358,N_14522,N_14853);
nand UO_1359 (O_1359,N_14870,N_14844);
nand UO_1360 (O_1360,N_14731,N_14970);
nor UO_1361 (O_1361,N_14687,N_14595);
and UO_1362 (O_1362,N_14816,N_14631);
and UO_1363 (O_1363,N_14780,N_14970);
or UO_1364 (O_1364,N_14865,N_14960);
or UO_1365 (O_1365,N_14594,N_14622);
xnor UO_1366 (O_1366,N_14944,N_14798);
nand UO_1367 (O_1367,N_14667,N_14860);
nor UO_1368 (O_1368,N_14521,N_14966);
nand UO_1369 (O_1369,N_14610,N_14990);
nor UO_1370 (O_1370,N_14728,N_14664);
or UO_1371 (O_1371,N_14593,N_14558);
and UO_1372 (O_1372,N_14562,N_14635);
nand UO_1373 (O_1373,N_14687,N_14735);
and UO_1374 (O_1374,N_14983,N_14608);
xor UO_1375 (O_1375,N_14858,N_14991);
and UO_1376 (O_1376,N_14549,N_14616);
nor UO_1377 (O_1377,N_14502,N_14562);
and UO_1378 (O_1378,N_14599,N_14981);
and UO_1379 (O_1379,N_14675,N_14806);
and UO_1380 (O_1380,N_14596,N_14716);
nand UO_1381 (O_1381,N_14880,N_14907);
and UO_1382 (O_1382,N_14611,N_14638);
xor UO_1383 (O_1383,N_14619,N_14925);
nand UO_1384 (O_1384,N_14829,N_14801);
and UO_1385 (O_1385,N_14844,N_14665);
or UO_1386 (O_1386,N_14939,N_14526);
nand UO_1387 (O_1387,N_14519,N_14562);
or UO_1388 (O_1388,N_14761,N_14671);
nand UO_1389 (O_1389,N_14556,N_14961);
or UO_1390 (O_1390,N_14679,N_14790);
or UO_1391 (O_1391,N_14868,N_14734);
nand UO_1392 (O_1392,N_14960,N_14647);
nor UO_1393 (O_1393,N_14563,N_14738);
nand UO_1394 (O_1394,N_14676,N_14879);
nand UO_1395 (O_1395,N_14777,N_14546);
and UO_1396 (O_1396,N_14924,N_14776);
xnor UO_1397 (O_1397,N_14541,N_14550);
or UO_1398 (O_1398,N_14906,N_14878);
and UO_1399 (O_1399,N_14661,N_14533);
and UO_1400 (O_1400,N_14685,N_14805);
or UO_1401 (O_1401,N_14783,N_14922);
nand UO_1402 (O_1402,N_14636,N_14848);
xor UO_1403 (O_1403,N_14862,N_14890);
and UO_1404 (O_1404,N_14712,N_14678);
nor UO_1405 (O_1405,N_14517,N_14934);
nor UO_1406 (O_1406,N_14698,N_14603);
nor UO_1407 (O_1407,N_14802,N_14907);
and UO_1408 (O_1408,N_14648,N_14859);
or UO_1409 (O_1409,N_14613,N_14643);
nor UO_1410 (O_1410,N_14984,N_14989);
nand UO_1411 (O_1411,N_14808,N_14903);
nand UO_1412 (O_1412,N_14776,N_14582);
nand UO_1413 (O_1413,N_14947,N_14835);
or UO_1414 (O_1414,N_14732,N_14877);
and UO_1415 (O_1415,N_14631,N_14704);
nor UO_1416 (O_1416,N_14750,N_14692);
nand UO_1417 (O_1417,N_14933,N_14507);
or UO_1418 (O_1418,N_14628,N_14906);
nor UO_1419 (O_1419,N_14701,N_14709);
nand UO_1420 (O_1420,N_14979,N_14801);
nand UO_1421 (O_1421,N_14797,N_14551);
nand UO_1422 (O_1422,N_14508,N_14981);
and UO_1423 (O_1423,N_14602,N_14562);
nand UO_1424 (O_1424,N_14569,N_14651);
nand UO_1425 (O_1425,N_14989,N_14619);
and UO_1426 (O_1426,N_14705,N_14767);
and UO_1427 (O_1427,N_14632,N_14735);
nand UO_1428 (O_1428,N_14995,N_14556);
nand UO_1429 (O_1429,N_14717,N_14976);
nor UO_1430 (O_1430,N_14785,N_14845);
or UO_1431 (O_1431,N_14788,N_14536);
or UO_1432 (O_1432,N_14660,N_14740);
and UO_1433 (O_1433,N_14520,N_14642);
nor UO_1434 (O_1434,N_14543,N_14570);
nand UO_1435 (O_1435,N_14794,N_14617);
nor UO_1436 (O_1436,N_14832,N_14522);
and UO_1437 (O_1437,N_14617,N_14661);
nand UO_1438 (O_1438,N_14638,N_14568);
or UO_1439 (O_1439,N_14711,N_14517);
nor UO_1440 (O_1440,N_14876,N_14586);
and UO_1441 (O_1441,N_14809,N_14780);
nor UO_1442 (O_1442,N_14666,N_14933);
or UO_1443 (O_1443,N_14827,N_14716);
nor UO_1444 (O_1444,N_14598,N_14886);
nor UO_1445 (O_1445,N_14663,N_14612);
nand UO_1446 (O_1446,N_14753,N_14678);
or UO_1447 (O_1447,N_14533,N_14760);
nand UO_1448 (O_1448,N_14553,N_14699);
and UO_1449 (O_1449,N_14670,N_14828);
nand UO_1450 (O_1450,N_14760,N_14558);
and UO_1451 (O_1451,N_14699,N_14572);
nor UO_1452 (O_1452,N_14805,N_14968);
nor UO_1453 (O_1453,N_14732,N_14615);
or UO_1454 (O_1454,N_14881,N_14526);
nand UO_1455 (O_1455,N_14741,N_14977);
nor UO_1456 (O_1456,N_14780,N_14581);
nand UO_1457 (O_1457,N_14692,N_14570);
or UO_1458 (O_1458,N_14846,N_14620);
nor UO_1459 (O_1459,N_14558,N_14720);
or UO_1460 (O_1460,N_14783,N_14513);
nor UO_1461 (O_1461,N_14607,N_14965);
nand UO_1462 (O_1462,N_14951,N_14878);
xnor UO_1463 (O_1463,N_14910,N_14610);
nand UO_1464 (O_1464,N_14564,N_14655);
xor UO_1465 (O_1465,N_14831,N_14991);
nand UO_1466 (O_1466,N_14780,N_14527);
and UO_1467 (O_1467,N_14852,N_14744);
or UO_1468 (O_1468,N_14561,N_14983);
and UO_1469 (O_1469,N_14792,N_14786);
or UO_1470 (O_1470,N_14914,N_14765);
xor UO_1471 (O_1471,N_14593,N_14884);
or UO_1472 (O_1472,N_14858,N_14567);
nand UO_1473 (O_1473,N_14729,N_14725);
xnor UO_1474 (O_1474,N_14646,N_14822);
nand UO_1475 (O_1475,N_14612,N_14857);
xnor UO_1476 (O_1476,N_14776,N_14645);
or UO_1477 (O_1477,N_14502,N_14911);
nor UO_1478 (O_1478,N_14711,N_14872);
nor UO_1479 (O_1479,N_14695,N_14759);
nor UO_1480 (O_1480,N_14704,N_14655);
or UO_1481 (O_1481,N_14665,N_14623);
nand UO_1482 (O_1482,N_14929,N_14856);
nor UO_1483 (O_1483,N_14536,N_14919);
nor UO_1484 (O_1484,N_14651,N_14946);
or UO_1485 (O_1485,N_14785,N_14999);
or UO_1486 (O_1486,N_14551,N_14625);
or UO_1487 (O_1487,N_14605,N_14612);
nand UO_1488 (O_1488,N_14662,N_14692);
and UO_1489 (O_1489,N_14528,N_14543);
and UO_1490 (O_1490,N_14509,N_14560);
nand UO_1491 (O_1491,N_14751,N_14634);
or UO_1492 (O_1492,N_14540,N_14581);
and UO_1493 (O_1493,N_14913,N_14696);
nor UO_1494 (O_1494,N_14677,N_14600);
or UO_1495 (O_1495,N_14874,N_14658);
nor UO_1496 (O_1496,N_14940,N_14762);
nor UO_1497 (O_1497,N_14973,N_14859);
xor UO_1498 (O_1498,N_14580,N_14579);
nor UO_1499 (O_1499,N_14988,N_14887);
or UO_1500 (O_1500,N_14873,N_14618);
nand UO_1501 (O_1501,N_14882,N_14760);
and UO_1502 (O_1502,N_14536,N_14713);
and UO_1503 (O_1503,N_14988,N_14839);
and UO_1504 (O_1504,N_14932,N_14564);
nand UO_1505 (O_1505,N_14518,N_14968);
or UO_1506 (O_1506,N_14820,N_14962);
nor UO_1507 (O_1507,N_14532,N_14783);
nor UO_1508 (O_1508,N_14961,N_14913);
xor UO_1509 (O_1509,N_14807,N_14553);
nand UO_1510 (O_1510,N_14581,N_14826);
nor UO_1511 (O_1511,N_14603,N_14681);
and UO_1512 (O_1512,N_14640,N_14582);
and UO_1513 (O_1513,N_14877,N_14800);
or UO_1514 (O_1514,N_14558,N_14643);
nand UO_1515 (O_1515,N_14589,N_14800);
or UO_1516 (O_1516,N_14822,N_14905);
nor UO_1517 (O_1517,N_14598,N_14887);
nor UO_1518 (O_1518,N_14817,N_14629);
nor UO_1519 (O_1519,N_14510,N_14517);
and UO_1520 (O_1520,N_14705,N_14710);
or UO_1521 (O_1521,N_14619,N_14904);
nor UO_1522 (O_1522,N_14894,N_14523);
or UO_1523 (O_1523,N_14917,N_14654);
nand UO_1524 (O_1524,N_14860,N_14765);
xor UO_1525 (O_1525,N_14706,N_14781);
nand UO_1526 (O_1526,N_14891,N_14552);
nor UO_1527 (O_1527,N_14959,N_14514);
or UO_1528 (O_1528,N_14929,N_14832);
and UO_1529 (O_1529,N_14813,N_14726);
nor UO_1530 (O_1530,N_14847,N_14988);
nor UO_1531 (O_1531,N_14524,N_14726);
and UO_1532 (O_1532,N_14946,N_14753);
nor UO_1533 (O_1533,N_14930,N_14886);
nand UO_1534 (O_1534,N_14521,N_14612);
or UO_1535 (O_1535,N_14835,N_14537);
nor UO_1536 (O_1536,N_14622,N_14792);
and UO_1537 (O_1537,N_14931,N_14968);
or UO_1538 (O_1538,N_14732,N_14708);
or UO_1539 (O_1539,N_14848,N_14731);
nor UO_1540 (O_1540,N_14660,N_14770);
or UO_1541 (O_1541,N_14677,N_14957);
and UO_1542 (O_1542,N_14634,N_14692);
nand UO_1543 (O_1543,N_14722,N_14784);
or UO_1544 (O_1544,N_14641,N_14596);
nand UO_1545 (O_1545,N_14562,N_14663);
xor UO_1546 (O_1546,N_14512,N_14644);
or UO_1547 (O_1547,N_14678,N_14662);
nand UO_1548 (O_1548,N_14790,N_14626);
nand UO_1549 (O_1549,N_14789,N_14761);
or UO_1550 (O_1550,N_14830,N_14960);
xor UO_1551 (O_1551,N_14919,N_14548);
and UO_1552 (O_1552,N_14841,N_14879);
and UO_1553 (O_1553,N_14976,N_14806);
xor UO_1554 (O_1554,N_14685,N_14938);
or UO_1555 (O_1555,N_14620,N_14556);
nor UO_1556 (O_1556,N_14559,N_14992);
nand UO_1557 (O_1557,N_14539,N_14927);
nand UO_1558 (O_1558,N_14973,N_14655);
xor UO_1559 (O_1559,N_14914,N_14972);
nor UO_1560 (O_1560,N_14753,N_14743);
or UO_1561 (O_1561,N_14965,N_14840);
xor UO_1562 (O_1562,N_14551,N_14834);
xnor UO_1563 (O_1563,N_14784,N_14537);
and UO_1564 (O_1564,N_14647,N_14699);
xor UO_1565 (O_1565,N_14860,N_14773);
or UO_1566 (O_1566,N_14597,N_14635);
xnor UO_1567 (O_1567,N_14683,N_14545);
and UO_1568 (O_1568,N_14688,N_14879);
nand UO_1569 (O_1569,N_14862,N_14597);
xnor UO_1570 (O_1570,N_14828,N_14879);
and UO_1571 (O_1571,N_14676,N_14862);
or UO_1572 (O_1572,N_14966,N_14933);
nor UO_1573 (O_1573,N_14588,N_14701);
and UO_1574 (O_1574,N_14857,N_14565);
nand UO_1575 (O_1575,N_14965,N_14756);
or UO_1576 (O_1576,N_14782,N_14724);
xor UO_1577 (O_1577,N_14649,N_14810);
nor UO_1578 (O_1578,N_14820,N_14902);
nor UO_1579 (O_1579,N_14771,N_14943);
nor UO_1580 (O_1580,N_14509,N_14517);
and UO_1581 (O_1581,N_14871,N_14633);
or UO_1582 (O_1582,N_14582,N_14611);
and UO_1583 (O_1583,N_14718,N_14539);
nor UO_1584 (O_1584,N_14559,N_14663);
and UO_1585 (O_1585,N_14730,N_14650);
and UO_1586 (O_1586,N_14624,N_14835);
and UO_1587 (O_1587,N_14835,N_14833);
nand UO_1588 (O_1588,N_14620,N_14661);
nor UO_1589 (O_1589,N_14647,N_14897);
nand UO_1590 (O_1590,N_14649,N_14632);
or UO_1591 (O_1591,N_14568,N_14856);
or UO_1592 (O_1592,N_14960,N_14931);
and UO_1593 (O_1593,N_14988,N_14905);
xor UO_1594 (O_1594,N_14910,N_14753);
xor UO_1595 (O_1595,N_14683,N_14927);
nor UO_1596 (O_1596,N_14851,N_14631);
and UO_1597 (O_1597,N_14828,N_14947);
nand UO_1598 (O_1598,N_14567,N_14711);
and UO_1599 (O_1599,N_14810,N_14706);
or UO_1600 (O_1600,N_14822,N_14870);
xnor UO_1601 (O_1601,N_14721,N_14944);
xnor UO_1602 (O_1602,N_14622,N_14591);
nor UO_1603 (O_1603,N_14825,N_14797);
xor UO_1604 (O_1604,N_14675,N_14742);
and UO_1605 (O_1605,N_14744,N_14989);
or UO_1606 (O_1606,N_14596,N_14992);
and UO_1607 (O_1607,N_14653,N_14836);
and UO_1608 (O_1608,N_14612,N_14826);
xor UO_1609 (O_1609,N_14941,N_14755);
nor UO_1610 (O_1610,N_14978,N_14812);
and UO_1611 (O_1611,N_14777,N_14972);
nor UO_1612 (O_1612,N_14835,N_14919);
and UO_1613 (O_1613,N_14904,N_14776);
and UO_1614 (O_1614,N_14954,N_14878);
and UO_1615 (O_1615,N_14945,N_14576);
and UO_1616 (O_1616,N_14953,N_14549);
and UO_1617 (O_1617,N_14867,N_14582);
nor UO_1618 (O_1618,N_14991,N_14535);
or UO_1619 (O_1619,N_14826,N_14869);
and UO_1620 (O_1620,N_14913,N_14861);
nand UO_1621 (O_1621,N_14578,N_14886);
or UO_1622 (O_1622,N_14904,N_14552);
or UO_1623 (O_1623,N_14588,N_14509);
and UO_1624 (O_1624,N_14845,N_14846);
nor UO_1625 (O_1625,N_14880,N_14776);
nor UO_1626 (O_1626,N_14664,N_14926);
nand UO_1627 (O_1627,N_14510,N_14603);
xnor UO_1628 (O_1628,N_14524,N_14733);
or UO_1629 (O_1629,N_14803,N_14747);
xnor UO_1630 (O_1630,N_14940,N_14850);
nor UO_1631 (O_1631,N_14683,N_14768);
nand UO_1632 (O_1632,N_14878,N_14739);
or UO_1633 (O_1633,N_14572,N_14959);
or UO_1634 (O_1634,N_14931,N_14957);
and UO_1635 (O_1635,N_14559,N_14928);
and UO_1636 (O_1636,N_14642,N_14509);
xor UO_1637 (O_1637,N_14965,N_14883);
or UO_1638 (O_1638,N_14666,N_14630);
or UO_1639 (O_1639,N_14527,N_14718);
nand UO_1640 (O_1640,N_14622,N_14869);
nor UO_1641 (O_1641,N_14618,N_14554);
nand UO_1642 (O_1642,N_14927,N_14699);
nand UO_1643 (O_1643,N_14773,N_14577);
nand UO_1644 (O_1644,N_14741,N_14873);
and UO_1645 (O_1645,N_14811,N_14878);
and UO_1646 (O_1646,N_14778,N_14536);
and UO_1647 (O_1647,N_14686,N_14824);
or UO_1648 (O_1648,N_14719,N_14553);
nand UO_1649 (O_1649,N_14536,N_14571);
and UO_1650 (O_1650,N_14720,N_14500);
or UO_1651 (O_1651,N_14733,N_14506);
nor UO_1652 (O_1652,N_14757,N_14644);
and UO_1653 (O_1653,N_14627,N_14876);
and UO_1654 (O_1654,N_14953,N_14976);
nand UO_1655 (O_1655,N_14733,N_14710);
nand UO_1656 (O_1656,N_14745,N_14791);
nand UO_1657 (O_1657,N_14917,N_14541);
nand UO_1658 (O_1658,N_14529,N_14512);
nand UO_1659 (O_1659,N_14762,N_14984);
xor UO_1660 (O_1660,N_14884,N_14630);
and UO_1661 (O_1661,N_14878,N_14546);
xnor UO_1662 (O_1662,N_14549,N_14518);
or UO_1663 (O_1663,N_14654,N_14599);
or UO_1664 (O_1664,N_14542,N_14643);
or UO_1665 (O_1665,N_14535,N_14608);
nor UO_1666 (O_1666,N_14820,N_14536);
xnor UO_1667 (O_1667,N_14865,N_14986);
nand UO_1668 (O_1668,N_14531,N_14865);
xnor UO_1669 (O_1669,N_14845,N_14683);
or UO_1670 (O_1670,N_14935,N_14941);
nor UO_1671 (O_1671,N_14816,N_14985);
xor UO_1672 (O_1672,N_14640,N_14689);
nand UO_1673 (O_1673,N_14766,N_14734);
and UO_1674 (O_1674,N_14950,N_14999);
nor UO_1675 (O_1675,N_14714,N_14775);
nor UO_1676 (O_1676,N_14678,N_14771);
nor UO_1677 (O_1677,N_14918,N_14959);
nand UO_1678 (O_1678,N_14848,N_14892);
or UO_1679 (O_1679,N_14946,N_14974);
nand UO_1680 (O_1680,N_14618,N_14544);
nor UO_1681 (O_1681,N_14537,N_14625);
and UO_1682 (O_1682,N_14562,N_14686);
nand UO_1683 (O_1683,N_14794,N_14848);
xor UO_1684 (O_1684,N_14587,N_14538);
and UO_1685 (O_1685,N_14877,N_14693);
nand UO_1686 (O_1686,N_14830,N_14620);
or UO_1687 (O_1687,N_14777,N_14842);
nor UO_1688 (O_1688,N_14527,N_14646);
or UO_1689 (O_1689,N_14535,N_14641);
nor UO_1690 (O_1690,N_14789,N_14978);
nand UO_1691 (O_1691,N_14515,N_14869);
or UO_1692 (O_1692,N_14948,N_14796);
and UO_1693 (O_1693,N_14997,N_14616);
nand UO_1694 (O_1694,N_14820,N_14817);
nand UO_1695 (O_1695,N_14892,N_14549);
or UO_1696 (O_1696,N_14993,N_14823);
and UO_1697 (O_1697,N_14885,N_14787);
and UO_1698 (O_1698,N_14677,N_14732);
nor UO_1699 (O_1699,N_14989,N_14979);
nor UO_1700 (O_1700,N_14661,N_14758);
nand UO_1701 (O_1701,N_14776,N_14611);
nor UO_1702 (O_1702,N_14876,N_14790);
nor UO_1703 (O_1703,N_14554,N_14753);
or UO_1704 (O_1704,N_14564,N_14567);
nand UO_1705 (O_1705,N_14917,N_14978);
or UO_1706 (O_1706,N_14878,N_14696);
and UO_1707 (O_1707,N_14969,N_14513);
xor UO_1708 (O_1708,N_14916,N_14747);
and UO_1709 (O_1709,N_14504,N_14737);
or UO_1710 (O_1710,N_14938,N_14862);
xnor UO_1711 (O_1711,N_14982,N_14828);
or UO_1712 (O_1712,N_14899,N_14643);
nand UO_1713 (O_1713,N_14943,N_14757);
xnor UO_1714 (O_1714,N_14603,N_14541);
and UO_1715 (O_1715,N_14732,N_14661);
or UO_1716 (O_1716,N_14749,N_14551);
nand UO_1717 (O_1717,N_14586,N_14746);
nand UO_1718 (O_1718,N_14929,N_14743);
nor UO_1719 (O_1719,N_14733,N_14721);
nor UO_1720 (O_1720,N_14622,N_14831);
xor UO_1721 (O_1721,N_14920,N_14955);
xor UO_1722 (O_1722,N_14614,N_14940);
or UO_1723 (O_1723,N_14642,N_14611);
nand UO_1724 (O_1724,N_14620,N_14672);
and UO_1725 (O_1725,N_14985,N_14764);
nor UO_1726 (O_1726,N_14934,N_14828);
or UO_1727 (O_1727,N_14612,N_14770);
nor UO_1728 (O_1728,N_14974,N_14630);
and UO_1729 (O_1729,N_14593,N_14682);
and UO_1730 (O_1730,N_14563,N_14573);
nor UO_1731 (O_1731,N_14558,N_14692);
and UO_1732 (O_1732,N_14636,N_14512);
or UO_1733 (O_1733,N_14915,N_14870);
nor UO_1734 (O_1734,N_14977,N_14853);
and UO_1735 (O_1735,N_14578,N_14708);
xnor UO_1736 (O_1736,N_14570,N_14537);
xor UO_1737 (O_1737,N_14786,N_14780);
nor UO_1738 (O_1738,N_14816,N_14663);
xnor UO_1739 (O_1739,N_14919,N_14960);
nand UO_1740 (O_1740,N_14793,N_14631);
xnor UO_1741 (O_1741,N_14519,N_14501);
nand UO_1742 (O_1742,N_14942,N_14774);
nand UO_1743 (O_1743,N_14884,N_14751);
nand UO_1744 (O_1744,N_14807,N_14932);
and UO_1745 (O_1745,N_14625,N_14972);
or UO_1746 (O_1746,N_14759,N_14855);
and UO_1747 (O_1747,N_14884,N_14709);
nand UO_1748 (O_1748,N_14596,N_14844);
xnor UO_1749 (O_1749,N_14675,N_14620);
xor UO_1750 (O_1750,N_14762,N_14713);
or UO_1751 (O_1751,N_14965,N_14967);
or UO_1752 (O_1752,N_14621,N_14632);
or UO_1753 (O_1753,N_14755,N_14582);
nand UO_1754 (O_1754,N_14956,N_14716);
and UO_1755 (O_1755,N_14845,N_14830);
and UO_1756 (O_1756,N_14980,N_14579);
and UO_1757 (O_1757,N_14750,N_14985);
and UO_1758 (O_1758,N_14695,N_14926);
or UO_1759 (O_1759,N_14907,N_14848);
xor UO_1760 (O_1760,N_14957,N_14649);
and UO_1761 (O_1761,N_14955,N_14725);
nor UO_1762 (O_1762,N_14769,N_14853);
nor UO_1763 (O_1763,N_14635,N_14528);
and UO_1764 (O_1764,N_14724,N_14583);
and UO_1765 (O_1765,N_14685,N_14584);
nor UO_1766 (O_1766,N_14553,N_14716);
and UO_1767 (O_1767,N_14723,N_14821);
nand UO_1768 (O_1768,N_14690,N_14658);
and UO_1769 (O_1769,N_14654,N_14738);
nor UO_1770 (O_1770,N_14846,N_14623);
and UO_1771 (O_1771,N_14849,N_14924);
or UO_1772 (O_1772,N_14583,N_14972);
or UO_1773 (O_1773,N_14532,N_14908);
nand UO_1774 (O_1774,N_14963,N_14864);
and UO_1775 (O_1775,N_14603,N_14506);
or UO_1776 (O_1776,N_14885,N_14608);
xnor UO_1777 (O_1777,N_14881,N_14733);
and UO_1778 (O_1778,N_14816,N_14625);
or UO_1779 (O_1779,N_14676,N_14748);
or UO_1780 (O_1780,N_14710,N_14737);
or UO_1781 (O_1781,N_14637,N_14755);
and UO_1782 (O_1782,N_14852,N_14836);
or UO_1783 (O_1783,N_14817,N_14827);
xor UO_1784 (O_1784,N_14969,N_14575);
nor UO_1785 (O_1785,N_14516,N_14660);
or UO_1786 (O_1786,N_14842,N_14568);
xnor UO_1787 (O_1787,N_14844,N_14939);
or UO_1788 (O_1788,N_14520,N_14971);
nor UO_1789 (O_1789,N_14546,N_14857);
xor UO_1790 (O_1790,N_14941,N_14862);
and UO_1791 (O_1791,N_14976,N_14658);
or UO_1792 (O_1792,N_14940,N_14934);
or UO_1793 (O_1793,N_14888,N_14643);
nor UO_1794 (O_1794,N_14668,N_14553);
and UO_1795 (O_1795,N_14682,N_14962);
nand UO_1796 (O_1796,N_14989,N_14757);
nor UO_1797 (O_1797,N_14956,N_14885);
nor UO_1798 (O_1798,N_14845,N_14527);
or UO_1799 (O_1799,N_14519,N_14721);
nand UO_1800 (O_1800,N_14779,N_14636);
or UO_1801 (O_1801,N_14768,N_14648);
or UO_1802 (O_1802,N_14776,N_14869);
nor UO_1803 (O_1803,N_14870,N_14832);
nand UO_1804 (O_1804,N_14715,N_14759);
nor UO_1805 (O_1805,N_14599,N_14620);
or UO_1806 (O_1806,N_14883,N_14719);
xnor UO_1807 (O_1807,N_14681,N_14871);
nor UO_1808 (O_1808,N_14872,N_14570);
or UO_1809 (O_1809,N_14575,N_14569);
or UO_1810 (O_1810,N_14920,N_14680);
or UO_1811 (O_1811,N_14551,N_14651);
nand UO_1812 (O_1812,N_14661,N_14723);
and UO_1813 (O_1813,N_14602,N_14972);
nor UO_1814 (O_1814,N_14725,N_14848);
nand UO_1815 (O_1815,N_14914,N_14705);
nand UO_1816 (O_1816,N_14952,N_14824);
nor UO_1817 (O_1817,N_14871,N_14616);
and UO_1818 (O_1818,N_14784,N_14879);
nand UO_1819 (O_1819,N_14964,N_14797);
nand UO_1820 (O_1820,N_14612,N_14522);
or UO_1821 (O_1821,N_14542,N_14815);
nor UO_1822 (O_1822,N_14623,N_14967);
or UO_1823 (O_1823,N_14835,N_14891);
or UO_1824 (O_1824,N_14885,N_14808);
nand UO_1825 (O_1825,N_14566,N_14915);
and UO_1826 (O_1826,N_14631,N_14743);
nand UO_1827 (O_1827,N_14632,N_14946);
and UO_1828 (O_1828,N_14584,N_14853);
nand UO_1829 (O_1829,N_14704,N_14748);
nor UO_1830 (O_1830,N_14541,N_14559);
or UO_1831 (O_1831,N_14599,N_14780);
nor UO_1832 (O_1832,N_14611,N_14998);
nand UO_1833 (O_1833,N_14633,N_14708);
nand UO_1834 (O_1834,N_14803,N_14945);
nor UO_1835 (O_1835,N_14692,N_14950);
and UO_1836 (O_1836,N_14722,N_14720);
nand UO_1837 (O_1837,N_14891,N_14948);
nand UO_1838 (O_1838,N_14838,N_14589);
nand UO_1839 (O_1839,N_14750,N_14670);
and UO_1840 (O_1840,N_14854,N_14711);
and UO_1841 (O_1841,N_14740,N_14635);
and UO_1842 (O_1842,N_14693,N_14842);
nand UO_1843 (O_1843,N_14519,N_14911);
xnor UO_1844 (O_1844,N_14653,N_14831);
nand UO_1845 (O_1845,N_14925,N_14818);
nor UO_1846 (O_1846,N_14612,N_14822);
or UO_1847 (O_1847,N_14758,N_14725);
nor UO_1848 (O_1848,N_14899,N_14713);
nor UO_1849 (O_1849,N_14854,N_14624);
or UO_1850 (O_1850,N_14772,N_14566);
nand UO_1851 (O_1851,N_14836,N_14874);
and UO_1852 (O_1852,N_14509,N_14606);
and UO_1853 (O_1853,N_14699,N_14756);
or UO_1854 (O_1854,N_14714,N_14682);
or UO_1855 (O_1855,N_14707,N_14822);
or UO_1856 (O_1856,N_14705,N_14978);
nor UO_1857 (O_1857,N_14869,N_14841);
nor UO_1858 (O_1858,N_14978,N_14794);
and UO_1859 (O_1859,N_14680,N_14795);
nand UO_1860 (O_1860,N_14520,N_14756);
or UO_1861 (O_1861,N_14754,N_14673);
xor UO_1862 (O_1862,N_14523,N_14953);
xor UO_1863 (O_1863,N_14518,N_14894);
and UO_1864 (O_1864,N_14746,N_14984);
and UO_1865 (O_1865,N_14611,N_14787);
nor UO_1866 (O_1866,N_14753,N_14783);
nor UO_1867 (O_1867,N_14598,N_14975);
nor UO_1868 (O_1868,N_14721,N_14633);
xor UO_1869 (O_1869,N_14501,N_14682);
nor UO_1870 (O_1870,N_14718,N_14576);
nor UO_1871 (O_1871,N_14756,N_14627);
and UO_1872 (O_1872,N_14699,N_14906);
nor UO_1873 (O_1873,N_14551,N_14916);
nand UO_1874 (O_1874,N_14671,N_14974);
or UO_1875 (O_1875,N_14777,N_14914);
nand UO_1876 (O_1876,N_14853,N_14726);
or UO_1877 (O_1877,N_14897,N_14688);
nand UO_1878 (O_1878,N_14566,N_14950);
and UO_1879 (O_1879,N_14524,N_14886);
nor UO_1880 (O_1880,N_14867,N_14779);
nand UO_1881 (O_1881,N_14883,N_14978);
and UO_1882 (O_1882,N_14971,N_14979);
and UO_1883 (O_1883,N_14998,N_14627);
and UO_1884 (O_1884,N_14994,N_14672);
nor UO_1885 (O_1885,N_14540,N_14577);
nand UO_1886 (O_1886,N_14817,N_14812);
and UO_1887 (O_1887,N_14822,N_14647);
xnor UO_1888 (O_1888,N_14543,N_14514);
nor UO_1889 (O_1889,N_14934,N_14725);
and UO_1890 (O_1890,N_14533,N_14706);
or UO_1891 (O_1891,N_14846,N_14750);
nor UO_1892 (O_1892,N_14823,N_14636);
nand UO_1893 (O_1893,N_14549,N_14848);
xnor UO_1894 (O_1894,N_14512,N_14562);
nand UO_1895 (O_1895,N_14867,N_14786);
or UO_1896 (O_1896,N_14538,N_14932);
and UO_1897 (O_1897,N_14763,N_14842);
and UO_1898 (O_1898,N_14577,N_14978);
or UO_1899 (O_1899,N_14802,N_14816);
and UO_1900 (O_1900,N_14791,N_14602);
nand UO_1901 (O_1901,N_14835,N_14736);
nor UO_1902 (O_1902,N_14886,N_14823);
nor UO_1903 (O_1903,N_14514,N_14702);
xnor UO_1904 (O_1904,N_14911,N_14735);
and UO_1905 (O_1905,N_14555,N_14958);
xor UO_1906 (O_1906,N_14720,N_14900);
or UO_1907 (O_1907,N_14730,N_14505);
nor UO_1908 (O_1908,N_14941,N_14917);
nor UO_1909 (O_1909,N_14855,N_14864);
nor UO_1910 (O_1910,N_14548,N_14670);
nand UO_1911 (O_1911,N_14867,N_14566);
nand UO_1912 (O_1912,N_14601,N_14760);
and UO_1913 (O_1913,N_14775,N_14938);
and UO_1914 (O_1914,N_14972,N_14680);
nand UO_1915 (O_1915,N_14639,N_14846);
nand UO_1916 (O_1916,N_14616,N_14780);
xor UO_1917 (O_1917,N_14530,N_14573);
nand UO_1918 (O_1918,N_14894,N_14515);
or UO_1919 (O_1919,N_14972,N_14813);
and UO_1920 (O_1920,N_14944,N_14892);
or UO_1921 (O_1921,N_14956,N_14561);
and UO_1922 (O_1922,N_14608,N_14889);
nor UO_1923 (O_1923,N_14871,N_14826);
and UO_1924 (O_1924,N_14857,N_14910);
and UO_1925 (O_1925,N_14967,N_14504);
and UO_1926 (O_1926,N_14619,N_14766);
and UO_1927 (O_1927,N_14933,N_14977);
nor UO_1928 (O_1928,N_14920,N_14515);
and UO_1929 (O_1929,N_14519,N_14531);
or UO_1930 (O_1930,N_14872,N_14689);
and UO_1931 (O_1931,N_14681,N_14952);
or UO_1932 (O_1932,N_14936,N_14738);
nor UO_1933 (O_1933,N_14641,N_14810);
or UO_1934 (O_1934,N_14703,N_14988);
and UO_1935 (O_1935,N_14861,N_14854);
nor UO_1936 (O_1936,N_14826,N_14751);
and UO_1937 (O_1937,N_14548,N_14502);
nor UO_1938 (O_1938,N_14891,N_14757);
nor UO_1939 (O_1939,N_14771,N_14762);
and UO_1940 (O_1940,N_14854,N_14516);
xor UO_1941 (O_1941,N_14912,N_14561);
nor UO_1942 (O_1942,N_14545,N_14530);
or UO_1943 (O_1943,N_14826,N_14746);
xnor UO_1944 (O_1944,N_14512,N_14714);
and UO_1945 (O_1945,N_14944,N_14927);
or UO_1946 (O_1946,N_14563,N_14718);
nor UO_1947 (O_1947,N_14935,N_14555);
or UO_1948 (O_1948,N_14898,N_14706);
or UO_1949 (O_1949,N_14815,N_14704);
or UO_1950 (O_1950,N_14909,N_14861);
nand UO_1951 (O_1951,N_14835,N_14817);
nor UO_1952 (O_1952,N_14910,N_14808);
nor UO_1953 (O_1953,N_14618,N_14883);
nor UO_1954 (O_1954,N_14564,N_14602);
nor UO_1955 (O_1955,N_14675,N_14572);
nand UO_1956 (O_1956,N_14852,N_14646);
nor UO_1957 (O_1957,N_14893,N_14597);
nor UO_1958 (O_1958,N_14894,N_14867);
nor UO_1959 (O_1959,N_14570,N_14534);
or UO_1960 (O_1960,N_14826,N_14965);
and UO_1961 (O_1961,N_14690,N_14886);
and UO_1962 (O_1962,N_14919,N_14611);
and UO_1963 (O_1963,N_14608,N_14521);
nor UO_1964 (O_1964,N_14776,N_14980);
nor UO_1965 (O_1965,N_14721,N_14634);
xor UO_1966 (O_1966,N_14652,N_14865);
and UO_1967 (O_1967,N_14600,N_14811);
nor UO_1968 (O_1968,N_14520,N_14562);
or UO_1969 (O_1969,N_14812,N_14871);
or UO_1970 (O_1970,N_14820,N_14760);
nand UO_1971 (O_1971,N_14830,N_14799);
xor UO_1972 (O_1972,N_14664,N_14887);
nand UO_1973 (O_1973,N_14945,N_14954);
xor UO_1974 (O_1974,N_14920,N_14977);
nand UO_1975 (O_1975,N_14773,N_14627);
xnor UO_1976 (O_1976,N_14914,N_14901);
nand UO_1977 (O_1977,N_14804,N_14703);
or UO_1978 (O_1978,N_14596,N_14602);
xor UO_1979 (O_1979,N_14740,N_14848);
or UO_1980 (O_1980,N_14602,N_14988);
nand UO_1981 (O_1981,N_14964,N_14682);
and UO_1982 (O_1982,N_14871,N_14969);
nand UO_1983 (O_1983,N_14921,N_14818);
nand UO_1984 (O_1984,N_14768,N_14987);
nand UO_1985 (O_1985,N_14920,N_14753);
nor UO_1986 (O_1986,N_14541,N_14853);
or UO_1987 (O_1987,N_14767,N_14630);
and UO_1988 (O_1988,N_14556,N_14673);
nand UO_1989 (O_1989,N_14609,N_14859);
nand UO_1990 (O_1990,N_14871,N_14939);
or UO_1991 (O_1991,N_14763,N_14985);
or UO_1992 (O_1992,N_14666,N_14890);
or UO_1993 (O_1993,N_14920,N_14732);
and UO_1994 (O_1994,N_14610,N_14700);
and UO_1995 (O_1995,N_14851,N_14810);
nor UO_1996 (O_1996,N_14917,N_14946);
or UO_1997 (O_1997,N_14773,N_14644);
nand UO_1998 (O_1998,N_14820,N_14909);
and UO_1999 (O_1999,N_14840,N_14847);
endmodule