module basic_500_3000_500_4_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_100,In_452);
and U1 (N_1,In_129,In_89);
nand U2 (N_2,In_324,In_363);
nor U3 (N_3,In_30,In_132);
and U4 (N_4,In_462,In_305);
nand U5 (N_5,In_329,In_242);
nand U6 (N_6,In_469,In_17);
nand U7 (N_7,In_133,In_116);
or U8 (N_8,In_451,In_63);
nand U9 (N_9,In_463,In_314);
nor U10 (N_10,In_176,In_230);
and U11 (N_11,In_7,In_39);
nand U12 (N_12,In_321,In_273);
xor U13 (N_13,In_361,In_486);
or U14 (N_14,In_69,In_115);
or U15 (N_15,In_343,In_299);
or U16 (N_16,In_415,In_281);
nor U17 (N_17,In_379,In_64);
or U18 (N_18,In_254,In_471);
and U19 (N_19,In_164,In_278);
and U20 (N_20,In_438,In_330);
or U21 (N_21,In_134,In_121);
and U22 (N_22,In_288,In_47);
and U23 (N_23,In_204,In_465);
nor U24 (N_24,In_177,In_218);
nor U25 (N_25,In_226,In_10);
nand U26 (N_26,In_456,In_90);
xor U27 (N_27,In_419,In_221);
or U28 (N_28,In_479,In_447);
nand U29 (N_29,In_280,In_464);
nand U30 (N_30,In_449,In_161);
nand U31 (N_31,In_398,In_61);
or U32 (N_32,In_215,In_388);
and U33 (N_33,In_406,In_458);
and U34 (N_34,In_453,In_411);
or U35 (N_35,In_24,In_78);
and U36 (N_36,In_207,In_118);
and U37 (N_37,In_228,In_189);
or U38 (N_38,In_171,In_274);
nand U39 (N_39,In_326,In_301);
or U40 (N_40,In_378,In_153);
nand U41 (N_41,In_184,In_444);
and U42 (N_42,In_422,In_131);
and U43 (N_43,In_202,In_498);
nor U44 (N_44,In_68,In_167);
nand U45 (N_45,In_428,In_491);
nand U46 (N_46,In_26,In_310);
nor U47 (N_47,In_147,In_474);
nand U48 (N_48,In_79,In_473);
nor U49 (N_49,In_200,In_284);
or U50 (N_50,In_99,In_331);
nand U51 (N_51,In_454,In_266);
and U52 (N_52,In_238,In_37);
or U53 (N_53,In_72,In_224);
nand U54 (N_54,In_32,In_103);
or U55 (N_55,In_159,In_29);
and U56 (N_56,In_381,In_31);
and U57 (N_57,In_359,In_225);
and U58 (N_58,In_76,In_125);
nand U59 (N_59,In_407,In_283);
nor U60 (N_60,In_23,In_259);
or U61 (N_61,In_57,In_107);
nor U62 (N_62,In_65,In_25);
or U63 (N_63,In_303,In_455);
nand U64 (N_64,In_442,In_44);
or U65 (N_65,In_272,In_145);
or U66 (N_66,In_353,In_162);
nor U67 (N_67,In_157,In_85);
or U68 (N_68,In_377,In_433);
and U69 (N_69,In_5,In_172);
and U70 (N_70,In_168,In_156);
or U71 (N_71,In_182,In_423);
nor U72 (N_72,In_470,In_128);
nand U73 (N_73,In_143,In_175);
or U74 (N_74,In_396,In_387);
nor U75 (N_75,In_246,In_41);
nor U76 (N_76,In_55,In_448);
nor U77 (N_77,In_234,In_389);
and U78 (N_78,In_190,In_249);
or U79 (N_79,In_136,In_276);
and U80 (N_80,In_193,In_466);
nor U81 (N_81,In_316,In_441);
and U82 (N_82,In_130,In_46);
or U83 (N_83,In_319,In_459);
nor U84 (N_84,In_122,In_142);
nand U85 (N_85,In_489,In_35);
or U86 (N_86,In_351,In_420);
nand U87 (N_87,In_210,In_251);
nor U88 (N_88,In_443,In_426);
nand U89 (N_89,In_374,In_252);
nand U90 (N_90,In_194,In_376);
or U91 (N_91,In_87,In_345);
nand U92 (N_92,In_302,In_139);
nand U93 (N_93,In_227,In_391);
nand U94 (N_94,In_430,In_279);
or U95 (N_95,In_82,In_109);
or U96 (N_96,In_220,In_113);
and U97 (N_97,In_102,In_320);
nor U98 (N_98,In_244,In_88);
nand U99 (N_99,In_337,In_309);
nand U100 (N_100,In_95,In_306);
nor U101 (N_101,In_27,In_154);
or U102 (N_102,In_327,In_21);
or U103 (N_103,In_360,In_339);
and U104 (N_104,In_372,In_492);
nand U105 (N_105,In_166,In_62);
nand U106 (N_106,In_20,In_98);
nand U107 (N_107,In_245,In_402);
or U108 (N_108,In_212,In_18);
or U109 (N_109,In_350,In_9);
nor U110 (N_110,In_185,In_105);
or U111 (N_111,In_148,In_385);
or U112 (N_112,In_120,In_290);
and U113 (N_113,In_83,In_257);
and U114 (N_114,In_400,In_155);
and U115 (N_115,In_181,In_293);
or U116 (N_116,In_275,In_137);
or U117 (N_117,In_219,In_412);
and U118 (N_118,In_261,In_174);
and U119 (N_119,In_267,In_341);
and U120 (N_120,In_141,In_483);
nor U121 (N_121,In_53,In_393);
nor U122 (N_122,In_28,In_467);
and U123 (N_123,In_253,In_362);
and U124 (N_124,In_386,In_186);
nor U125 (N_125,In_268,In_424);
and U126 (N_126,In_16,In_425);
nand U127 (N_127,In_344,In_373);
or U128 (N_128,In_66,In_262);
and U129 (N_129,In_269,In_36);
nand U130 (N_130,In_12,In_352);
nor U131 (N_131,In_265,In_52);
or U132 (N_132,In_3,In_50);
nor U133 (N_133,In_296,In_260);
or U134 (N_134,In_475,In_311);
and U135 (N_135,In_56,In_367);
nand U136 (N_136,In_356,In_255);
nor U137 (N_137,In_472,In_317);
nor U138 (N_138,In_71,In_188);
nor U139 (N_139,In_468,In_499);
nand U140 (N_140,In_355,In_446);
nor U141 (N_141,In_460,In_158);
nand U142 (N_142,In_110,In_308);
nor U143 (N_143,In_114,In_417);
nand U144 (N_144,In_410,In_497);
and U145 (N_145,In_409,In_282);
nor U146 (N_146,In_370,In_42);
and U147 (N_147,In_160,In_315);
nand U148 (N_148,In_432,In_233);
or U149 (N_149,In_271,In_96);
xor U150 (N_150,In_0,In_248);
and U151 (N_151,In_342,In_11);
and U152 (N_152,In_217,In_196);
nand U153 (N_153,In_146,In_322);
nor U154 (N_154,In_416,In_59);
and U155 (N_155,In_237,In_431);
or U156 (N_156,In_427,In_395);
nand U157 (N_157,In_332,In_49);
nor U158 (N_158,In_124,In_77);
nand U159 (N_159,In_384,In_394);
or U160 (N_160,In_476,In_364);
nand U161 (N_161,In_413,In_478);
and U162 (N_162,In_240,In_40);
and U163 (N_163,In_151,In_150);
nor U164 (N_164,In_22,In_323);
nor U165 (N_165,In_493,In_8);
nor U166 (N_166,In_169,In_232);
or U167 (N_167,In_33,In_418);
or U168 (N_168,In_357,In_199);
and U169 (N_169,In_91,In_73);
nor U170 (N_170,In_192,In_104);
nand U171 (N_171,In_484,In_354);
or U172 (N_172,In_457,In_440);
nand U173 (N_173,In_366,In_48);
and U174 (N_174,In_127,In_119);
and U175 (N_175,In_6,In_439);
or U176 (N_176,In_236,In_117);
nand U177 (N_177,In_365,In_383);
xor U178 (N_178,In_289,In_135);
and U179 (N_179,In_223,In_198);
and U180 (N_180,In_358,In_292);
and U181 (N_181,In_111,In_495);
nor U182 (N_182,In_318,In_216);
and U183 (N_183,In_173,In_206);
nand U184 (N_184,In_86,In_4);
or U185 (N_185,In_347,In_54);
and U186 (N_186,In_195,In_80);
and U187 (N_187,In_60,In_304);
nor U188 (N_188,In_399,In_93);
and U189 (N_189,In_461,In_371);
or U190 (N_190,In_15,In_229);
or U191 (N_191,In_434,In_138);
and U192 (N_192,In_34,In_397);
nor U193 (N_193,In_19,In_382);
nor U194 (N_194,In_403,In_336);
nor U195 (N_195,In_300,In_258);
nand U196 (N_196,In_298,In_297);
nor U197 (N_197,In_334,In_149);
nor U198 (N_198,In_70,In_94);
nor U199 (N_199,In_390,In_144);
and U200 (N_200,In_178,In_180);
xnor U201 (N_201,In_165,In_235);
or U202 (N_202,In_270,In_140);
nand U203 (N_203,In_101,In_286);
and U204 (N_204,In_287,In_201);
or U205 (N_205,In_163,In_312);
nor U206 (N_206,In_231,In_313);
nor U207 (N_207,In_263,In_74);
nand U208 (N_208,In_81,In_2);
and U209 (N_209,In_250,In_408);
nor U210 (N_210,In_214,In_106);
or U211 (N_211,In_436,In_429);
or U212 (N_212,In_295,In_277);
and U213 (N_213,In_437,In_191);
nor U214 (N_214,In_97,In_222);
or U215 (N_215,In_203,In_112);
or U216 (N_216,In_349,In_445);
nand U217 (N_217,In_209,In_392);
or U218 (N_218,In_338,In_494);
and U219 (N_219,In_123,In_92);
nand U220 (N_220,In_256,In_375);
and U221 (N_221,In_435,In_368);
or U222 (N_222,In_108,In_14);
nand U223 (N_223,In_51,In_208);
nand U224 (N_224,In_340,In_75);
and U225 (N_225,In_481,In_401);
or U226 (N_226,In_485,In_480);
nor U227 (N_227,In_307,In_179);
or U228 (N_228,In_414,In_405);
and U229 (N_229,In_264,In_325);
and U230 (N_230,In_496,In_213);
and U231 (N_231,In_43,In_241);
nor U232 (N_232,In_335,In_477);
or U233 (N_233,In_490,In_333);
or U234 (N_234,In_488,In_421);
and U235 (N_235,In_294,In_369);
nand U236 (N_236,In_243,In_346);
or U237 (N_237,In_348,In_247);
or U238 (N_238,In_450,In_45);
and U239 (N_239,In_380,In_84);
or U240 (N_240,In_328,In_211);
and U241 (N_241,In_58,In_205);
or U242 (N_242,In_197,In_170);
nand U243 (N_243,In_152,In_38);
nand U244 (N_244,In_13,In_404);
nor U245 (N_245,In_1,In_187);
xnor U246 (N_246,In_239,In_183);
nor U247 (N_247,In_487,In_285);
nor U248 (N_248,In_67,In_291);
nand U249 (N_249,In_126,In_482);
nand U250 (N_250,In_186,In_281);
or U251 (N_251,In_188,In_336);
nand U252 (N_252,In_231,In_192);
or U253 (N_253,In_146,In_127);
and U254 (N_254,In_171,In_345);
nor U255 (N_255,In_370,In_490);
or U256 (N_256,In_123,In_147);
nor U257 (N_257,In_484,In_141);
and U258 (N_258,In_233,In_478);
nand U259 (N_259,In_455,In_372);
nand U260 (N_260,In_477,In_471);
nand U261 (N_261,In_83,In_157);
and U262 (N_262,In_124,In_182);
nand U263 (N_263,In_479,In_344);
nand U264 (N_264,In_497,In_357);
or U265 (N_265,In_16,In_486);
or U266 (N_266,In_406,In_44);
nand U267 (N_267,In_10,In_219);
nor U268 (N_268,In_154,In_284);
and U269 (N_269,In_315,In_79);
or U270 (N_270,In_318,In_415);
nor U271 (N_271,In_114,In_380);
or U272 (N_272,In_456,In_112);
nor U273 (N_273,In_293,In_49);
nand U274 (N_274,In_362,In_10);
or U275 (N_275,In_69,In_94);
and U276 (N_276,In_367,In_163);
or U277 (N_277,In_40,In_295);
and U278 (N_278,In_393,In_117);
nor U279 (N_279,In_181,In_351);
nor U280 (N_280,In_48,In_451);
nand U281 (N_281,In_477,In_73);
nor U282 (N_282,In_376,In_451);
nor U283 (N_283,In_378,In_19);
or U284 (N_284,In_218,In_499);
nor U285 (N_285,In_335,In_15);
or U286 (N_286,In_364,In_401);
nor U287 (N_287,In_230,In_376);
and U288 (N_288,In_377,In_436);
or U289 (N_289,In_136,In_4);
nor U290 (N_290,In_486,In_207);
nor U291 (N_291,In_406,In_333);
nor U292 (N_292,In_48,In_262);
nor U293 (N_293,In_454,In_420);
and U294 (N_294,In_63,In_458);
nand U295 (N_295,In_258,In_498);
nor U296 (N_296,In_299,In_310);
nand U297 (N_297,In_461,In_472);
nand U298 (N_298,In_381,In_396);
or U299 (N_299,In_365,In_8);
or U300 (N_300,In_31,In_259);
nor U301 (N_301,In_225,In_416);
nor U302 (N_302,In_277,In_423);
and U303 (N_303,In_369,In_370);
nor U304 (N_304,In_169,In_343);
and U305 (N_305,In_202,In_100);
and U306 (N_306,In_309,In_168);
and U307 (N_307,In_246,In_118);
and U308 (N_308,In_470,In_455);
or U309 (N_309,In_285,In_266);
or U310 (N_310,In_254,In_176);
nor U311 (N_311,In_474,In_258);
nand U312 (N_312,In_114,In_284);
or U313 (N_313,In_126,In_200);
or U314 (N_314,In_238,In_303);
or U315 (N_315,In_462,In_148);
or U316 (N_316,In_312,In_33);
or U317 (N_317,In_367,In_386);
and U318 (N_318,In_311,In_1);
nor U319 (N_319,In_175,In_477);
or U320 (N_320,In_34,In_491);
nor U321 (N_321,In_348,In_400);
nor U322 (N_322,In_267,In_70);
nor U323 (N_323,In_202,In_382);
and U324 (N_324,In_257,In_446);
and U325 (N_325,In_434,In_61);
nand U326 (N_326,In_266,In_4);
or U327 (N_327,In_130,In_140);
and U328 (N_328,In_195,In_142);
nor U329 (N_329,In_487,In_433);
nand U330 (N_330,In_478,In_197);
nor U331 (N_331,In_343,In_304);
nand U332 (N_332,In_300,In_499);
or U333 (N_333,In_10,In_31);
nand U334 (N_334,In_426,In_499);
nor U335 (N_335,In_254,In_169);
nor U336 (N_336,In_102,In_418);
nand U337 (N_337,In_45,In_485);
nand U338 (N_338,In_143,In_298);
and U339 (N_339,In_428,In_365);
nor U340 (N_340,In_373,In_432);
nand U341 (N_341,In_9,In_455);
nor U342 (N_342,In_385,In_295);
nor U343 (N_343,In_435,In_125);
nand U344 (N_344,In_471,In_251);
and U345 (N_345,In_356,In_298);
nor U346 (N_346,In_356,In_374);
or U347 (N_347,In_292,In_413);
nor U348 (N_348,In_122,In_428);
or U349 (N_349,In_329,In_285);
and U350 (N_350,In_399,In_84);
or U351 (N_351,In_148,In_194);
or U352 (N_352,In_416,In_25);
nand U353 (N_353,In_71,In_334);
nor U354 (N_354,In_37,In_62);
or U355 (N_355,In_141,In_77);
or U356 (N_356,In_493,In_455);
or U357 (N_357,In_335,In_122);
or U358 (N_358,In_291,In_351);
and U359 (N_359,In_270,In_154);
or U360 (N_360,In_246,In_260);
nand U361 (N_361,In_407,In_311);
nand U362 (N_362,In_318,In_22);
nand U363 (N_363,In_402,In_270);
nand U364 (N_364,In_435,In_72);
nor U365 (N_365,In_369,In_394);
nand U366 (N_366,In_16,In_373);
nand U367 (N_367,In_330,In_10);
and U368 (N_368,In_233,In_188);
or U369 (N_369,In_484,In_311);
nor U370 (N_370,In_293,In_214);
nor U371 (N_371,In_235,In_334);
and U372 (N_372,In_230,In_216);
and U373 (N_373,In_168,In_391);
nor U374 (N_374,In_394,In_81);
nor U375 (N_375,In_332,In_300);
or U376 (N_376,In_167,In_490);
and U377 (N_377,In_495,In_240);
and U378 (N_378,In_387,In_82);
and U379 (N_379,In_439,In_64);
nor U380 (N_380,In_302,In_290);
nor U381 (N_381,In_108,In_270);
nor U382 (N_382,In_431,In_421);
nor U383 (N_383,In_221,In_449);
nor U384 (N_384,In_97,In_82);
or U385 (N_385,In_10,In_188);
nor U386 (N_386,In_128,In_10);
nor U387 (N_387,In_192,In_317);
and U388 (N_388,In_89,In_150);
nor U389 (N_389,In_239,In_163);
nor U390 (N_390,In_308,In_255);
or U391 (N_391,In_156,In_49);
nand U392 (N_392,In_60,In_45);
and U393 (N_393,In_127,In_205);
nand U394 (N_394,In_257,In_152);
xnor U395 (N_395,In_22,In_24);
and U396 (N_396,In_409,In_349);
and U397 (N_397,In_317,In_151);
or U398 (N_398,In_175,In_330);
nand U399 (N_399,In_405,In_322);
or U400 (N_400,In_359,In_294);
nand U401 (N_401,In_69,In_67);
or U402 (N_402,In_412,In_42);
nand U403 (N_403,In_200,In_79);
or U404 (N_404,In_414,In_425);
and U405 (N_405,In_244,In_207);
and U406 (N_406,In_18,In_162);
nor U407 (N_407,In_82,In_409);
nor U408 (N_408,In_450,In_247);
nand U409 (N_409,In_327,In_490);
and U410 (N_410,In_226,In_237);
or U411 (N_411,In_98,In_194);
or U412 (N_412,In_67,In_173);
nor U413 (N_413,In_423,In_198);
nor U414 (N_414,In_266,In_413);
and U415 (N_415,In_322,In_66);
and U416 (N_416,In_36,In_244);
nand U417 (N_417,In_479,In_37);
nor U418 (N_418,In_104,In_10);
nand U419 (N_419,In_95,In_178);
or U420 (N_420,In_226,In_14);
nand U421 (N_421,In_348,In_313);
and U422 (N_422,In_191,In_304);
nand U423 (N_423,In_86,In_323);
and U424 (N_424,In_191,In_261);
or U425 (N_425,In_497,In_235);
nand U426 (N_426,In_243,In_409);
nor U427 (N_427,In_240,In_338);
nand U428 (N_428,In_488,In_221);
nor U429 (N_429,In_93,In_365);
or U430 (N_430,In_228,In_107);
nor U431 (N_431,In_338,In_45);
or U432 (N_432,In_124,In_112);
or U433 (N_433,In_79,In_128);
nor U434 (N_434,In_371,In_221);
nor U435 (N_435,In_284,In_389);
or U436 (N_436,In_496,In_306);
nor U437 (N_437,In_52,In_451);
nand U438 (N_438,In_433,In_6);
and U439 (N_439,In_47,In_113);
nand U440 (N_440,In_0,In_446);
and U441 (N_441,In_225,In_181);
or U442 (N_442,In_165,In_51);
or U443 (N_443,In_264,In_497);
and U444 (N_444,In_65,In_410);
or U445 (N_445,In_256,In_181);
nor U446 (N_446,In_402,In_260);
nand U447 (N_447,In_220,In_331);
and U448 (N_448,In_185,In_66);
and U449 (N_449,In_74,In_401);
or U450 (N_450,In_246,In_3);
nand U451 (N_451,In_58,In_258);
or U452 (N_452,In_404,In_371);
or U453 (N_453,In_191,In_386);
or U454 (N_454,In_76,In_450);
and U455 (N_455,In_314,In_141);
or U456 (N_456,In_256,In_8);
and U457 (N_457,In_295,In_289);
or U458 (N_458,In_161,In_94);
nor U459 (N_459,In_245,In_181);
or U460 (N_460,In_11,In_166);
nand U461 (N_461,In_53,In_276);
nor U462 (N_462,In_81,In_64);
or U463 (N_463,In_476,In_75);
nand U464 (N_464,In_119,In_367);
nor U465 (N_465,In_445,In_173);
or U466 (N_466,In_442,In_49);
and U467 (N_467,In_300,In_484);
and U468 (N_468,In_350,In_80);
or U469 (N_469,In_441,In_44);
or U470 (N_470,In_201,In_445);
nand U471 (N_471,In_222,In_429);
and U472 (N_472,In_166,In_492);
nor U473 (N_473,In_86,In_247);
nor U474 (N_474,In_304,In_302);
and U475 (N_475,In_483,In_106);
nor U476 (N_476,In_248,In_314);
or U477 (N_477,In_410,In_265);
nor U478 (N_478,In_4,In_350);
nand U479 (N_479,In_174,In_393);
or U480 (N_480,In_396,In_408);
nand U481 (N_481,In_423,In_191);
nor U482 (N_482,In_169,In_462);
and U483 (N_483,In_280,In_144);
nand U484 (N_484,In_318,In_310);
nor U485 (N_485,In_391,In_431);
or U486 (N_486,In_26,In_363);
nor U487 (N_487,In_110,In_100);
nor U488 (N_488,In_366,In_470);
nor U489 (N_489,In_150,In_462);
or U490 (N_490,In_244,In_53);
nand U491 (N_491,In_419,In_164);
or U492 (N_492,In_96,In_213);
and U493 (N_493,In_16,In_161);
and U494 (N_494,In_183,In_191);
nand U495 (N_495,In_292,In_374);
or U496 (N_496,In_433,In_296);
or U497 (N_497,In_26,In_376);
or U498 (N_498,In_188,In_493);
and U499 (N_499,In_251,In_321);
nor U500 (N_500,In_343,In_422);
nor U501 (N_501,In_204,In_234);
or U502 (N_502,In_119,In_375);
nor U503 (N_503,In_438,In_470);
or U504 (N_504,In_167,In_437);
nor U505 (N_505,In_253,In_357);
nand U506 (N_506,In_270,In_131);
and U507 (N_507,In_240,In_268);
and U508 (N_508,In_299,In_322);
nor U509 (N_509,In_58,In_322);
nand U510 (N_510,In_426,In_332);
nor U511 (N_511,In_319,In_190);
nand U512 (N_512,In_345,In_354);
and U513 (N_513,In_135,In_376);
or U514 (N_514,In_172,In_472);
nand U515 (N_515,In_148,In_140);
or U516 (N_516,In_476,In_163);
or U517 (N_517,In_203,In_256);
and U518 (N_518,In_372,In_466);
nor U519 (N_519,In_406,In_323);
nand U520 (N_520,In_417,In_10);
or U521 (N_521,In_153,In_495);
or U522 (N_522,In_292,In_209);
nand U523 (N_523,In_373,In_358);
nor U524 (N_524,In_460,In_97);
nor U525 (N_525,In_160,In_134);
or U526 (N_526,In_265,In_187);
nor U527 (N_527,In_413,In_146);
and U528 (N_528,In_393,In_26);
and U529 (N_529,In_481,In_148);
nand U530 (N_530,In_80,In_136);
or U531 (N_531,In_408,In_374);
and U532 (N_532,In_418,In_450);
nor U533 (N_533,In_451,In_114);
and U534 (N_534,In_410,In_472);
nand U535 (N_535,In_436,In_138);
nor U536 (N_536,In_208,In_259);
or U537 (N_537,In_248,In_82);
or U538 (N_538,In_53,In_295);
nand U539 (N_539,In_424,In_409);
or U540 (N_540,In_389,In_203);
nor U541 (N_541,In_303,In_275);
nor U542 (N_542,In_387,In_298);
nor U543 (N_543,In_197,In_95);
xor U544 (N_544,In_263,In_393);
and U545 (N_545,In_8,In_436);
nor U546 (N_546,In_66,In_69);
or U547 (N_547,In_213,In_329);
nor U548 (N_548,In_102,In_95);
or U549 (N_549,In_443,In_113);
nand U550 (N_550,In_478,In_126);
or U551 (N_551,In_441,In_58);
or U552 (N_552,In_39,In_28);
nor U553 (N_553,In_121,In_199);
xnor U554 (N_554,In_451,In_463);
and U555 (N_555,In_100,In_448);
and U556 (N_556,In_395,In_114);
or U557 (N_557,In_197,In_115);
and U558 (N_558,In_451,In_87);
or U559 (N_559,In_134,In_461);
nand U560 (N_560,In_76,In_327);
and U561 (N_561,In_312,In_108);
and U562 (N_562,In_54,In_44);
nor U563 (N_563,In_466,In_70);
xor U564 (N_564,In_108,In_132);
nand U565 (N_565,In_224,In_380);
and U566 (N_566,In_163,In_337);
xor U567 (N_567,In_155,In_280);
nand U568 (N_568,In_77,In_277);
nor U569 (N_569,In_184,In_105);
and U570 (N_570,In_153,In_379);
and U571 (N_571,In_239,In_76);
nand U572 (N_572,In_94,In_449);
nor U573 (N_573,In_490,In_239);
and U574 (N_574,In_89,In_56);
and U575 (N_575,In_2,In_82);
and U576 (N_576,In_341,In_408);
and U577 (N_577,In_23,In_289);
nand U578 (N_578,In_317,In_343);
and U579 (N_579,In_431,In_196);
or U580 (N_580,In_56,In_223);
and U581 (N_581,In_499,In_357);
or U582 (N_582,In_375,In_125);
nand U583 (N_583,In_135,In_494);
or U584 (N_584,In_35,In_475);
and U585 (N_585,In_44,In_65);
or U586 (N_586,In_451,In_43);
and U587 (N_587,In_342,In_325);
nor U588 (N_588,In_112,In_153);
or U589 (N_589,In_25,In_63);
or U590 (N_590,In_190,In_420);
nand U591 (N_591,In_457,In_368);
nand U592 (N_592,In_459,In_108);
nand U593 (N_593,In_496,In_486);
nor U594 (N_594,In_236,In_14);
nand U595 (N_595,In_416,In_379);
nor U596 (N_596,In_282,In_330);
nor U597 (N_597,In_488,In_247);
and U598 (N_598,In_376,In_435);
nand U599 (N_599,In_364,In_420);
nor U600 (N_600,In_366,In_285);
and U601 (N_601,In_337,In_381);
nand U602 (N_602,In_339,In_148);
or U603 (N_603,In_29,In_464);
and U604 (N_604,In_375,In_195);
and U605 (N_605,In_48,In_480);
nor U606 (N_606,In_452,In_228);
and U607 (N_607,In_407,In_282);
nor U608 (N_608,In_83,In_287);
or U609 (N_609,In_254,In_348);
nor U610 (N_610,In_206,In_471);
and U611 (N_611,In_35,In_487);
or U612 (N_612,In_178,In_278);
and U613 (N_613,In_499,In_379);
or U614 (N_614,In_168,In_440);
and U615 (N_615,In_318,In_297);
nand U616 (N_616,In_289,In_435);
nor U617 (N_617,In_8,In_272);
or U618 (N_618,In_374,In_429);
or U619 (N_619,In_126,In_235);
nor U620 (N_620,In_307,In_457);
or U621 (N_621,In_254,In_47);
or U622 (N_622,In_485,In_184);
or U623 (N_623,In_211,In_418);
and U624 (N_624,In_149,In_18);
or U625 (N_625,In_469,In_165);
and U626 (N_626,In_239,In_103);
or U627 (N_627,In_202,In_131);
nor U628 (N_628,In_141,In_103);
and U629 (N_629,In_484,In_187);
or U630 (N_630,In_331,In_452);
nor U631 (N_631,In_104,In_146);
nor U632 (N_632,In_303,In_482);
or U633 (N_633,In_453,In_458);
or U634 (N_634,In_420,In_169);
and U635 (N_635,In_334,In_36);
nand U636 (N_636,In_346,In_427);
nor U637 (N_637,In_3,In_456);
and U638 (N_638,In_154,In_7);
nand U639 (N_639,In_418,In_213);
or U640 (N_640,In_442,In_68);
nor U641 (N_641,In_41,In_480);
nand U642 (N_642,In_478,In_194);
nand U643 (N_643,In_119,In_171);
nor U644 (N_644,In_176,In_420);
nand U645 (N_645,In_157,In_66);
nand U646 (N_646,In_165,In_111);
or U647 (N_647,In_442,In_39);
nand U648 (N_648,In_272,In_393);
or U649 (N_649,In_72,In_189);
and U650 (N_650,In_183,In_492);
or U651 (N_651,In_455,In_199);
or U652 (N_652,In_475,In_421);
and U653 (N_653,In_345,In_173);
nand U654 (N_654,In_9,In_11);
or U655 (N_655,In_476,In_9);
nor U656 (N_656,In_482,In_438);
and U657 (N_657,In_96,In_50);
nand U658 (N_658,In_390,In_6);
nor U659 (N_659,In_423,In_264);
nor U660 (N_660,In_497,In_494);
or U661 (N_661,In_163,In_387);
and U662 (N_662,In_417,In_90);
nand U663 (N_663,In_247,In_274);
nand U664 (N_664,In_359,In_80);
and U665 (N_665,In_268,In_339);
nand U666 (N_666,In_412,In_143);
nand U667 (N_667,In_306,In_463);
nand U668 (N_668,In_215,In_484);
or U669 (N_669,In_189,In_455);
or U670 (N_670,In_296,In_60);
and U671 (N_671,In_194,In_41);
nor U672 (N_672,In_453,In_119);
nand U673 (N_673,In_209,In_370);
nor U674 (N_674,In_144,In_89);
and U675 (N_675,In_120,In_43);
and U676 (N_676,In_337,In_348);
or U677 (N_677,In_69,In_407);
nand U678 (N_678,In_234,In_364);
nand U679 (N_679,In_467,In_119);
or U680 (N_680,In_448,In_390);
or U681 (N_681,In_72,In_141);
nand U682 (N_682,In_19,In_171);
nand U683 (N_683,In_288,In_313);
nor U684 (N_684,In_398,In_85);
nor U685 (N_685,In_195,In_117);
or U686 (N_686,In_29,In_222);
nand U687 (N_687,In_73,In_63);
nand U688 (N_688,In_60,In_8);
nor U689 (N_689,In_31,In_292);
or U690 (N_690,In_498,In_90);
nand U691 (N_691,In_432,In_55);
or U692 (N_692,In_52,In_341);
or U693 (N_693,In_430,In_149);
nand U694 (N_694,In_483,In_218);
or U695 (N_695,In_348,In_168);
nand U696 (N_696,In_301,In_478);
and U697 (N_697,In_116,In_154);
xor U698 (N_698,In_453,In_210);
and U699 (N_699,In_370,In_13);
and U700 (N_700,In_316,In_486);
nor U701 (N_701,In_304,In_467);
nand U702 (N_702,In_357,In_395);
xnor U703 (N_703,In_372,In_349);
nor U704 (N_704,In_338,In_76);
nand U705 (N_705,In_23,In_161);
or U706 (N_706,In_87,In_241);
and U707 (N_707,In_308,In_171);
nand U708 (N_708,In_435,In_106);
nand U709 (N_709,In_206,In_463);
or U710 (N_710,In_359,In_23);
nor U711 (N_711,In_245,In_68);
and U712 (N_712,In_491,In_464);
nand U713 (N_713,In_395,In_494);
and U714 (N_714,In_206,In_77);
nor U715 (N_715,In_153,In_241);
or U716 (N_716,In_332,In_473);
or U717 (N_717,In_24,In_237);
nand U718 (N_718,In_345,In_195);
nor U719 (N_719,In_142,In_242);
nor U720 (N_720,In_206,In_261);
nand U721 (N_721,In_54,In_498);
nand U722 (N_722,In_398,In_208);
or U723 (N_723,In_162,In_446);
or U724 (N_724,In_90,In_329);
nand U725 (N_725,In_309,In_98);
or U726 (N_726,In_248,In_385);
nand U727 (N_727,In_48,In_164);
nand U728 (N_728,In_215,In_312);
and U729 (N_729,In_486,In_68);
or U730 (N_730,In_280,In_96);
or U731 (N_731,In_53,In_401);
or U732 (N_732,In_480,In_67);
nand U733 (N_733,In_413,In_85);
nand U734 (N_734,In_356,In_175);
nor U735 (N_735,In_218,In_379);
or U736 (N_736,In_132,In_395);
and U737 (N_737,In_90,In_356);
nand U738 (N_738,In_267,In_50);
nand U739 (N_739,In_289,In_70);
nand U740 (N_740,In_282,In_492);
nand U741 (N_741,In_371,In_259);
nor U742 (N_742,In_301,In_151);
or U743 (N_743,In_433,In_417);
nor U744 (N_744,In_140,In_49);
nand U745 (N_745,In_21,In_31);
or U746 (N_746,In_213,In_272);
nand U747 (N_747,In_123,In_288);
nor U748 (N_748,In_209,In_123);
or U749 (N_749,In_174,In_314);
or U750 (N_750,N_195,N_681);
or U751 (N_751,N_539,N_502);
and U752 (N_752,N_395,N_376);
nand U753 (N_753,N_89,N_439);
nor U754 (N_754,N_206,N_216);
nand U755 (N_755,N_414,N_109);
and U756 (N_756,N_583,N_349);
nand U757 (N_757,N_279,N_440);
nor U758 (N_758,N_96,N_425);
and U759 (N_759,N_254,N_340);
nand U760 (N_760,N_586,N_198);
nand U761 (N_761,N_114,N_68);
nand U762 (N_762,N_541,N_239);
nand U763 (N_763,N_394,N_661);
nor U764 (N_764,N_515,N_323);
nand U765 (N_765,N_590,N_564);
and U766 (N_766,N_10,N_650);
nand U767 (N_767,N_692,N_468);
nor U768 (N_768,N_173,N_164);
xor U769 (N_769,N_458,N_303);
and U770 (N_770,N_192,N_626);
or U771 (N_771,N_603,N_683);
and U772 (N_772,N_120,N_483);
nand U773 (N_773,N_166,N_133);
nor U774 (N_774,N_506,N_627);
nor U775 (N_775,N_33,N_437);
or U776 (N_776,N_320,N_350);
nor U777 (N_777,N_451,N_208);
nor U778 (N_778,N_494,N_175);
and U779 (N_779,N_579,N_34);
and U780 (N_780,N_82,N_629);
and U781 (N_781,N_495,N_509);
and U782 (N_782,N_550,N_314);
nor U783 (N_783,N_296,N_40);
nand U784 (N_784,N_419,N_185);
nand U785 (N_785,N_0,N_156);
nand U786 (N_786,N_74,N_283);
nor U787 (N_787,N_469,N_3);
nor U788 (N_788,N_570,N_429);
and U789 (N_789,N_118,N_568);
or U790 (N_790,N_381,N_83);
or U791 (N_791,N_292,N_605);
nor U792 (N_792,N_746,N_310);
nor U793 (N_793,N_398,N_426);
and U794 (N_794,N_35,N_269);
or U795 (N_795,N_624,N_235);
or U796 (N_796,N_739,N_344);
and U797 (N_797,N_607,N_363);
and U798 (N_798,N_190,N_702);
nor U799 (N_799,N_546,N_687);
or U800 (N_800,N_551,N_115);
xor U801 (N_801,N_246,N_379);
nor U802 (N_802,N_393,N_97);
or U803 (N_803,N_717,N_105);
nand U804 (N_804,N_421,N_259);
or U805 (N_805,N_636,N_496);
nand U806 (N_806,N_667,N_284);
and U807 (N_807,N_703,N_336);
and U808 (N_808,N_13,N_189);
or U809 (N_809,N_405,N_364);
nand U810 (N_810,N_224,N_202);
nor U811 (N_811,N_174,N_578);
or U812 (N_812,N_697,N_662);
nand U813 (N_813,N_531,N_46);
nor U814 (N_814,N_428,N_203);
and U815 (N_815,N_80,N_598);
nand U816 (N_816,N_261,N_389);
nor U817 (N_817,N_54,N_481);
or U818 (N_818,N_176,N_6);
nor U819 (N_819,N_641,N_633);
or U820 (N_820,N_138,N_463);
and U821 (N_821,N_396,N_265);
and U822 (N_822,N_326,N_31);
nand U823 (N_823,N_334,N_286);
and U824 (N_824,N_62,N_26);
and U825 (N_825,N_49,N_562);
nor U826 (N_826,N_305,N_94);
or U827 (N_827,N_719,N_744);
nor U828 (N_828,N_15,N_709);
or U829 (N_829,N_613,N_300);
nor U830 (N_830,N_293,N_722);
or U831 (N_831,N_272,N_512);
or U832 (N_832,N_447,N_17);
nand U833 (N_833,N_228,N_153);
and U834 (N_834,N_162,N_242);
and U835 (N_835,N_136,N_124);
nor U836 (N_836,N_580,N_595);
nor U837 (N_837,N_637,N_172);
nand U838 (N_838,N_346,N_371);
nand U839 (N_839,N_47,N_77);
nor U840 (N_840,N_322,N_736);
nor U841 (N_841,N_701,N_545);
nand U842 (N_842,N_225,N_731);
nor U843 (N_843,N_184,N_591);
or U844 (N_844,N_245,N_402);
nand U845 (N_845,N_612,N_2);
and U846 (N_846,N_248,N_369);
nor U847 (N_847,N_362,N_378);
or U848 (N_848,N_342,N_125);
and U849 (N_849,N_585,N_178);
nand U850 (N_850,N_90,N_331);
nand U851 (N_851,N_524,N_312);
or U852 (N_852,N_392,N_680);
or U853 (N_853,N_298,N_465);
or U854 (N_854,N_304,N_20);
and U855 (N_855,N_623,N_199);
nand U856 (N_856,N_672,N_27);
and U857 (N_857,N_519,N_560);
nor U858 (N_858,N_219,N_724);
and U859 (N_859,N_694,N_457);
nand U860 (N_860,N_733,N_299);
or U861 (N_861,N_521,N_217);
nand U862 (N_862,N_60,N_107);
nor U863 (N_863,N_42,N_422);
and U864 (N_864,N_423,N_128);
nand U865 (N_865,N_664,N_500);
or U866 (N_866,N_88,N_123);
nor U867 (N_867,N_193,N_668);
or U868 (N_868,N_39,N_599);
nor U869 (N_869,N_18,N_448);
nor U870 (N_870,N_654,N_59);
nand U871 (N_871,N_729,N_537);
or U872 (N_872,N_146,N_732);
nor U873 (N_873,N_79,N_597);
nand U874 (N_874,N_655,N_726);
or U875 (N_875,N_533,N_45);
or U876 (N_876,N_142,N_517);
nor U877 (N_877,N_489,N_51);
nor U878 (N_878,N_14,N_163);
or U879 (N_879,N_148,N_470);
nand U880 (N_880,N_460,N_477);
or U881 (N_881,N_76,N_737);
and U882 (N_882,N_55,N_253);
nor U883 (N_883,N_713,N_182);
and U884 (N_884,N_520,N_526);
or U885 (N_885,N_659,N_93);
and U886 (N_886,N_708,N_514);
or U887 (N_887,N_532,N_368);
or U888 (N_888,N_547,N_252);
nand U889 (N_889,N_475,N_432);
or U890 (N_890,N_277,N_614);
and U891 (N_891,N_19,N_622);
nand U892 (N_892,N_61,N_157);
and U893 (N_893,N_171,N_601);
or U894 (N_894,N_611,N_615);
or U895 (N_895,N_691,N_635);
nor U896 (N_896,N_528,N_628);
or U897 (N_897,N_271,N_332);
nor U898 (N_898,N_390,N_718);
nand U899 (N_899,N_618,N_365);
or U900 (N_900,N_281,N_99);
and U901 (N_901,N_32,N_576);
or U902 (N_902,N_467,N_464);
and U903 (N_903,N_165,N_410);
or U904 (N_904,N_499,N_740);
nor U905 (N_905,N_418,N_745);
nand U906 (N_906,N_387,N_56);
or U907 (N_907,N_41,N_738);
nand U908 (N_908,N_316,N_669);
nor U909 (N_909,N_24,N_542);
nand U910 (N_910,N_501,N_101);
or U911 (N_911,N_705,N_335);
or U912 (N_912,N_431,N_442);
nand U913 (N_913,N_540,N_725);
or U914 (N_914,N_98,N_241);
nand U915 (N_915,N_536,N_313);
nand U916 (N_916,N_573,N_529);
xnor U917 (N_917,N_492,N_433);
or U918 (N_918,N_22,N_625);
nor U919 (N_919,N_119,N_516);
nor U920 (N_920,N_69,N_329);
and U921 (N_921,N_232,N_169);
nor U922 (N_922,N_478,N_511);
and U923 (N_923,N_205,N_436);
or U924 (N_924,N_518,N_572);
nor U925 (N_925,N_152,N_671);
nor U926 (N_926,N_473,N_482);
or U927 (N_927,N_236,N_554);
and U928 (N_928,N_243,N_676);
or U929 (N_929,N_237,N_324);
and U930 (N_930,N_452,N_63);
nor U931 (N_931,N_592,N_522);
and U932 (N_932,N_663,N_454);
and U933 (N_933,N_177,N_297);
or U934 (N_934,N_584,N_409);
nand U935 (N_935,N_723,N_294);
nor U936 (N_936,N_122,N_357);
or U937 (N_937,N_604,N_397);
or U938 (N_938,N_657,N_221);
and U939 (N_939,N_160,N_684);
nor U940 (N_940,N_290,N_534);
nor U941 (N_941,N_333,N_700);
nor U942 (N_942,N_58,N_704);
nor U943 (N_943,N_412,N_581);
or U944 (N_944,N_354,N_274);
or U945 (N_945,N_386,N_188);
and U946 (N_946,N_391,N_73);
or U947 (N_947,N_367,N_260);
and U948 (N_948,N_507,N_181);
nor U949 (N_949,N_92,N_81);
or U950 (N_950,N_459,N_404);
nand U951 (N_951,N_487,N_488);
nand U952 (N_952,N_491,N_508);
nand U953 (N_953,N_1,N_677);
nor U954 (N_954,N_558,N_65);
nand U955 (N_955,N_621,N_159);
or U956 (N_956,N_446,N_596);
nand U957 (N_957,N_696,N_154);
nor U958 (N_958,N_543,N_234);
nand U959 (N_959,N_38,N_427);
or U960 (N_960,N_229,N_309);
or U961 (N_961,N_710,N_295);
and U962 (N_962,N_466,N_352);
or U963 (N_963,N_43,N_72);
and U964 (N_964,N_291,N_504);
nand U965 (N_965,N_472,N_377);
nand U966 (N_966,N_630,N_653);
or U967 (N_967,N_689,N_44);
and U968 (N_968,N_556,N_453);
and U969 (N_969,N_327,N_498);
nor U970 (N_970,N_308,N_688);
or U971 (N_971,N_571,N_417);
or U972 (N_972,N_247,N_366);
nor U973 (N_973,N_187,N_110);
nand U974 (N_974,N_158,N_484);
or U975 (N_975,N_321,N_450);
or U976 (N_976,N_85,N_36);
nor U977 (N_977,N_267,N_220);
and U978 (N_978,N_651,N_319);
or U979 (N_979,N_682,N_330);
xor U980 (N_980,N_104,N_204);
and U981 (N_981,N_510,N_186);
nor U982 (N_982,N_563,N_339);
and U983 (N_983,N_608,N_686);
or U984 (N_984,N_212,N_144);
and U985 (N_985,N_530,N_582);
and U986 (N_986,N_587,N_191);
and U987 (N_987,N_372,N_456);
nand U988 (N_988,N_147,N_301);
and U989 (N_989,N_355,N_102);
nor U990 (N_990,N_513,N_384);
nand U991 (N_991,N_179,N_170);
nor U992 (N_992,N_400,N_679);
nand U993 (N_993,N_370,N_9);
nand U994 (N_994,N_643,N_721);
nand U995 (N_995,N_743,N_616);
nor U996 (N_996,N_449,N_287);
nand U997 (N_997,N_549,N_403);
and U998 (N_998,N_359,N_553);
or U999 (N_999,N_634,N_730);
or U1000 (N_1000,N_353,N_360);
nor U1001 (N_1001,N_268,N_233);
and U1002 (N_1002,N_649,N_538);
or U1003 (N_1003,N_276,N_289);
or U1004 (N_1004,N_645,N_222);
nor U1005 (N_1005,N_476,N_648);
nand U1006 (N_1006,N_64,N_411);
nand U1007 (N_1007,N_5,N_486);
nor U1008 (N_1008,N_445,N_196);
nand U1009 (N_1009,N_673,N_84);
or U1010 (N_1010,N_318,N_282);
or U1011 (N_1011,N_180,N_646);
nand U1012 (N_1012,N_345,N_201);
nand U1013 (N_1013,N_111,N_108);
nand U1014 (N_1014,N_712,N_210);
or U1015 (N_1015,N_632,N_430);
nor U1016 (N_1016,N_194,N_620);
nor U1017 (N_1017,N_127,N_639);
or U1018 (N_1018,N_161,N_238);
or U1019 (N_1019,N_307,N_749);
or U1020 (N_1020,N_78,N_71);
and U1021 (N_1021,N_341,N_249);
and U1022 (N_1022,N_589,N_407);
nand U1023 (N_1023,N_374,N_602);
and U1024 (N_1024,N_117,N_67);
or U1025 (N_1025,N_617,N_151);
nor U1026 (N_1026,N_474,N_631);
nor U1027 (N_1027,N_383,N_461);
and U1028 (N_1028,N_706,N_285);
and U1029 (N_1029,N_255,N_600);
nand U1030 (N_1030,N_656,N_347);
or U1031 (N_1031,N_112,N_28);
nor U1032 (N_1032,N_685,N_716);
xor U1033 (N_1033,N_555,N_131);
or U1034 (N_1034,N_741,N_441);
nand U1035 (N_1035,N_727,N_48);
and U1036 (N_1036,N_214,N_168);
nor U1037 (N_1037,N_462,N_12);
nand U1038 (N_1038,N_742,N_561);
nand U1039 (N_1039,N_720,N_140);
and U1040 (N_1040,N_302,N_134);
nor U1041 (N_1041,N_523,N_527);
nand U1042 (N_1042,N_103,N_575);
nand U1043 (N_1043,N_552,N_257);
nand U1044 (N_1044,N_317,N_135);
or U1045 (N_1045,N_438,N_86);
nor U1046 (N_1046,N_594,N_70);
nor U1047 (N_1047,N_215,N_747);
and U1048 (N_1048,N_29,N_4);
nor U1049 (N_1049,N_343,N_503);
nor U1050 (N_1050,N_150,N_565);
and U1051 (N_1051,N_275,N_569);
or U1052 (N_1052,N_351,N_338);
or U1053 (N_1053,N_497,N_493);
or U1054 (N_1054,N_273,N_66);
nand U1055 (N_1055,N_471,N_141);
nand U1056 (N_1056,N_695,N_52);
or U1057 (N_1057,N_106,N_8);
or U1058 (N_1058,N_660,N_735);
nand U1059 (N_1059,N_53,N_665);
nand U1060 (N_1060,N_256,N_479);
and U1061 (N_1061,N_525,N_444);
and U1062 (N_1062,N_57,N_640);
or U1063 (N_1063,N_356,N_385);
or U1064 (N_1064,N_588,N_139);
and U1065 (N_1065,N_574,N_609);
nor U1066 (N_1066,N_388,N_707);
or U1067 (N_1067,N_167,N_7);
nand U1068 (N_1068,N_644,N_358);
or U1069 (N_1069,N_490,N_424);
nand U1070 (N_1070,N_715,N_728);
nand U1071 (N_1071,N_666,N_251);
nand U1072 (N_1072,N_270,N_557);
or U1073 (N_1073,N_408,N_213);
and U1074 (N_1074,N_675,N_137);
nand U1075 (N_1075,N_223,N_100);
and U1076 (N_1076,N_258,N_209);
or U1077 (N_1077,N_348,N_250);
nor U1078 (N_1078,N_155,N_647);
nor U1079 (N_1079,N_325,N_435);
nor U1080 (N_1080,N_264,N_416);
nor U1081 (N_1081,N_306,N_113);
and U1082 (N_1082,N_714,N_658);
nand U1083 (N_1083,N_652,N_231);
nand U1084 (N_1084,N_21,N_226);
nor U1085 (N_1085,N_544,N_548);
or U1086 (N_1086,N_420,N_25);
nand U1087 (N_1087,N_382,N_693);
and U1088 (N_1088,N_37,N_129);
nand U1089 (N_1089,N_230,N_559);
nor U1090 (N_1090,N_262,N_748);
nor U1091 (N_1091,N_328,N_200);
nor U1092 (N_1092,N_183,N_218);
nand U1093 (N_1093,N_406,N_399);
or U1094 (N_1094,N_149,N_480);
nor U1095 (N_1095,N_670,N_211);
nor U1096 (N_1096,N_567,N_413);
and U1097 (N_1097,N_485,N_674);
or U1098 (N_1098,N_566,N_95);
nand U1099 (N_1099,N_50,N_337);
or U1100 (N_1100,N_455,N_280);
nand U1101 (N_1101,N_126,N_642);
and U1102 (N_1102,N_91,N_263);
or U1103 (N_1103,N_207,N_711);
xor U1104 (N_1104,N_30,N_401);
nor U1105 (N_1105,N_244,N_278);
nand U1106 (N_1106,N_227,N_678);
nor U1107 (N_1107,N_361,N_593);
and U1108 (N_1108,N_143,N_505);
or U1109 (N_1109,N_698,N_610);
and U1110 (N_1110,N_638,N_116);
nor U1111 (N_1111,N_577,N_266);
or U1112 (N_1112,N_443,N_87);
and U1113 (N_1113,N_699,N_121);
nand U1114 (N_1114,N_11,N_690);
or U1115 (N_1115,N_619,N_535);
nor U1116 (N_1116,N_315,N_240);
and U1117 (N_1117,N_197,N_311);
xor U1118 (N_1118,N_16,N_23);
and U1119 (N_1119,N_375,N_75);
or U1120 (N_1120,N_130,N_734);
nand U1121 (N_1121,N_380,N_606);
nand U1122 (N_1122,N_145,N_288);
nand U1123 (N_1123,N_434,N_415);
or U1124 (N_1124,N_373,N_132);
or U1125 (N_1125,N_229,N_521);
and U1126 (N_1126,N_738,N_553);
nand U1127 (N_1127,N_383,N_453);
nor U1128 (N_1128,N_695,N_612);
nand U1129 (N_1129,N_227,N_340);
or U1130 (N_1130,N_569,N_369);
nor U1131 (N_1131,N_119,N_126);
and U1132 (N_1132,N_394,N_68);
or U1133 (N_1133,N_272,N_494);
nand U1134 (N_1134,N_570,N_330);
nor U1135 (N_1135,N_43,N_693);
xnor U1136 (N_1136,N_236,N_267);
nor U1137 (N_1137,N_286,N_745);
and U1138 (N_1138,N_408,N_61);
or U1139 (N_1139,N_525,N_419);
or U1140 (N_1140,N_82,N_415);
or U1141 (N_1141,N_478,N_597);
nand U1142 (N_1142,N_431,N_234);
nand U1143 (N_1143,N_310,N_178);
and U1144 (N_1144,N_78,N_26);
nand U1145 (N_1145,N_591,N_658);
or U1146 (N_1146,N_230,N_678);
or U1147 (N_1147,N_665,N_263);
and U1148 (N_1148,N_24,N_83);
nand U1149 (N_1149,N_115,N_577);
or U1150 (N_1150,N_38,N_3);
xnor U1151 (N_1151,N_712,N_148);
nand U1152 (N_1152,N_383,N_380);
and U1153 (N_1153,N_602,N_377);
and U1154 (N_1154,N_206,N_370);
or U1155 (N_1155,N_706,N_497);
or U1156 (N_1156,N_670,N_483);
or U1157 (N_1157,N_641,N_364);
nor U1158 (N_1158,N_48,N_575);
nand U1159 (N_1159,N_665,N_621);
nand U1160 (N_1160,N_194,N_730);
nor U1161 (N_1161,N_304,N_342);
nor U1162 (N_1162,N_542,N_84);
nand U1163 (N_1163,N_340,N_674);
and U1164 (N_1164,N_191,N_684);
and U1165 (N_1165,N_559,N_735);
nor U1166 (N_1166,N_560,N_601);
nand U1167 (N_1167,N_670,N_413);
or U1168 (N_1168,N_432,N_159);
and U1169 (N_1169,N_184,N_255);
nor U1170 (N_1170,N_295,N_511);
or U1171 (N_1171,N_8,N_458);
and U1172 (N_1172,N_324,N_617);
nor U1173 (N_1173,N_461,N_610);
and U1174 (N_1174,N_88,N_670);
nor U1175 (N_1175,N_621,N_372);
and U1176 (N_1176,N_414,N_593);
and U1177 (N_1177,N_352,N_389);
or U1178 (N_1178,N_386,N_709);
nor U1179 (N_1179,N_697,N_226);
nor U1180 (N_1180,N_213,N_86);
and U1181 (N_1181,N_385,N_115);
nor U1182 (N_1182,N_453,N_384);
or U1183 (N_1183,N_677,N_593);
nor U1184 (N_1184,N_592,N_102);
and U1185 (N_1185,N_455,N_15);
nand U1186 (N_1186,N_67,N_334);
nor U1187 (N_1187,N_49,N_229);
and U1188 (N_1188,N_445,N_490);
nor U1189 (N_1189,N_93,N_205);
and U1190 (N_1190,N_404,N_320);
and U1191 (N_1191,N_15,N_718);
or U1192 (N_1192,N_82,N_8);
nor U1193 (N_1193,N_279,N_714);
or U1194 (N_1194,N_535,N_84);
nor U1195 (N_1195,N_503,N_342);
or U1196 (N_1196,N_735,N_318);
and U1197 (N_1197,N_667,N_449);
or U1198 (N_1198,N_37,N_141);
and U1199 (N_1199,N_331,N_613);
and U1200 (N_1200,N_737,N_375);
and U1201 (N_1201,N_612,N_644);
nor U1202 (N_1202,N_204,N_582);
or U1203 (N_1203,N_114,N_517);
and U1204 (N_1204,N_240,N_531);
nor U1205 (N_1205,N_285,N_715);
or U1206 (N_1206,N_385,N_73);
nand U1207 (N_1207,N_95,N_549);
nand U1208 (N_1208,N_296,N_594);
or U1209 (N_1209,N_26,N_400);
or U1210 (N_1210,N_244,N_368);
nand U1211 (N_1211,N_123,N_133);
or U1212 (N_1212,N_591,N_595);
nor U1213 (N_1213,N_443,N_129);
nor U1214 (N_1214,N_486,N_563);
or U1215 (N_1215,N_460,N_305);
nor U1216 (N_1216,N_471,N_655);
and U1217 (N_1217,N_80,N_283);
or U1218 (N_1218,N_321,N_339);
nor U1219 (N_1219,N_333,N_605);
nor U1220 (N_1220,N_114,N_593);
or U1221 (N_1221,N_704,N_631);
or U1222 (N_1222,N_735,N_474);
nor U1223 (N_1223,N_116,N_588);
and U1224 (N_1224,N_543,N_315);
nor U1225 (N_1225,N_39,N_30);
nor U1226 (N_1226,N_114,N_615);
nor U1227 (N_1227,N_267,N_271);
nand U1228 (N_1228,N_132,N_507);
and U1229 (N_1229,N_428,N_120);
or U1230 (N_1230,N_171,N_63);
nand U1231 (N_1231,N_95,N_669);
or U1232 (N_1232,N_376,N_734);
nor U1233 (N_1233,N_667,N_237);
or U1234 (N_1234,N_607,N_645);
or U1235 (N_1235,N_298,N_668);
nand U1236 (N_1236,N_671,N_147);
nand U1237 (N_1237,N_236,N_402);
or U1238 (N_1238,N_212,N_47);
nor U1239 (N_1239,N_404,N_660);
and U1240 (N_1240,N_631,N_540);
and U1241 (N_1241,N_164,N_194);
nor U1242 (N_1242,N_191,N_280);
or U1243 (N_1243,N_529,N_76);
nor U1244 (N_1244,N_581,N_730);
and U1245 (N_1245,N_307,N_396);
and U1246 (N_1246,N_719,N_271);
or U1247 (N_1247,N_564,N_118);
nand U1248 (N_1248,N_239,N_721);
or U1249 (N_1249,N_301,N_388);
nor U1250 (N_1250,N_224,N_446);
nand U1251 (N_1251,N_164,N_515);
nand U1252 (N_1252,N_540,N_649);
and U1253 (N_1253,N_425,N_175);
nor U1254 (N_1254,N_290,N_9);
nand U1255 (N_1255,N_617,N_140);
nand U1256 (N_1256,N_39,N_384);
nor U1257 (N_1257,N_651,N_10);
nor U1258 (N_1258,N_401,N_632);
and U1259 (N_1259,N_617,N_577);
xor U1260 (N_1260,N_428,N_204);
nand U1261 (N_1261,N_454,N_343);
and U1262 (N_1262,N_151,N_384);
nand U1263 (N_1263,N_434,N_679);
nand U1264 (N_1264,N_398,N_201);
nor U1265 (N_1265,N_196,N_740);
and U1266 (N_1266,N_190,N_684);
nand U1267 (N_1267,N_638,N_47);
nand U1268 (N_1268,N_569,N_225);
nor U1269 (N_1269,N_65,N_490);
or U1270 (N_1270,N_271,N_134);
nand U1271 (N_1271,N_467,N_400);
or U1272 (N_1272,N_13,N_691);
or U1273 (N_1273,N_567,N_602);
nor U1274 (N_1274,N_144,N_560);
nor U1275 (N_1275,N_646,N_52);
and U1276 (N_1276,N_694,N_241);
and U1277 (N_1277,N_566,N_86);
nand U1278 (N_1278,N_75,N_650);
nand U1279 (N_1279,N_583,N_535);
and U1280 (N_1280,N_489,N_537);
nor U1281 (N_1281,N_562,N_294);
or U1282 (N_1282,N_234,N_556);
nand U1283 (N_1283,N_361,N_246);
and U1284 (N_1284,N_315,N_433);
and U1285 (N_1285,N_254,N_111);
nor U1286 (N_1286,N_476,N_448);
or U1287 (N_1287,N_401,N_119);
nand U1288 (N_1288,N_288,N_436);
and U1289 (N_1289,N_252,N_478);
or U1290 (N_1290,N_41,N_25);
and U1291 (N_1291,N_31,N_318);
nand U1292 (N_1292,N_687,N_565);
nor U1293 (N_1293,N_281,N_569);
or U1294 (N_1294,N_294,N_713);
or U1295 (N_1295,N_45,N_582);
nor U1296 (N_1296,N_747,N_724);
and U1297 (N_1297,N_511,N_7);
and U1298 (N_1298,N_124,N_349);
nand U1299 (N_1299,N_446,N_263);
or U1300 (N_1300,N_75,N_670);
nor U1301 (N_1301,N_521,N_355);
or U1302 (N_1302,N_719,N_239);
nand U1303 (N_1303,N_146,N_235);
and U1304 (N_1304,N_59,N_408);
nand U1305 (N_1305,N_184,N_325);
nand U1306 (N_1306,N_633,N_196);
nor U1307 (N_1307,N_329,N_423);
nor U1308 (N_1308,N_719,N_364);
and U1309 (N_1309,N_170,N_333);
nor U1310 (N_1310,N_594,N_5);
nand U1311 (N_1311,N_68,N_400);
or U1312 (N_1312,N_121,N_462);
nor U1313 (N_1313,N_550,N_290);
and U1314 (N_1314,N_282,N_720);
nand U1315 (N_1315,N_106,N_57);
nand U1316 (N_1316,N_613,N_507);
nor U1317 (N_1317,N_654,N_292);
nor U1318 (N_1318,N_595,N_84);
nand U1319 (N_1319,N_299,N_612);
nand U1320 (N_1320,N_593,N_218);
or U1321 (N_1321,N_368,N_616);
and U1322 (N_1322,N_502,N_201);
nor U1323 (N_1323,N_538,N_316);
nand U1324 (N_1324,N_589,N_519);
and U1325 (N_1325,N_519,N_325);
nand U1326 (N_1326,N_602,N_226);
or U1327 (N_1327,N_718,N_339);
nand U1328 (N_1328,N_189,N_394);
and U1329 (N_1329,N_467,N_680);
nand U1330 (N_1330,N_409,N_442);
nand U1331 (N_1331,N_238,N_359);
nor U1332 (N_1332,N_370,N_660);
and U1333 (N_1333,N_477,N_192);
and U1334 (N_1334,N_322,N_275);
nor U1335 (N_1335,N_724,N_591);
nand U1336 (N_1336,N_713,N_628);
nand U1337 (N_1337,N_270,N_41);
nor U1338 (N_1338,N_727,N_694);
and U1339 (N_1339,N_650,N_720);
nand U1340 (N_1340,N_125,N_404);
and U1341 (N_1341,N_323,N_222);
or U1342 (N_1342,N_426,N_307);
or U1343 (N_1343,N_338,N_153);
nand U1344 (N_1344,N_88,N_561);
or U1345 (N_1345,N_35,N_28);
and U1346 (N_1346,N_539,N_421);
and U1347 (N_1347,N_407,N_335);
nand U1348 (N_1348,N_240,N_648);
nand U1349 (N_1349,N_349,N_448);
or U1350 (N_1350,N_428,N_610);
or U1351 (N_1351,N_631,N_570);
and U1352 (N_1352,N_349,N_321);
or U1353 (N_1353,N_367,N_681);
nor U1354 (N_1354,N_199,N_725);
or U1355 (N_1355,N_550,N_203);
nand U1356 (N_1356,N_126,N_103);
xnor U1357 (N_1357,N_346,N_132);
or U1358 (N_1358,N_79,N_645);
and U1359 (N_1359,N_261,N_625);
nor U1360 (N_1360,N_100,N_14);
nor U1361 (N_1361,N_404,N_46);
or U1362 (N_1362,N_574,N_637);
or U1363 (N_1363,N_494,N_74);
nor U1364 (N_1364,N_123,N_375);
nor U1365 (N_1365,N_167,N_572);
nor U1366 (N_1366,N_158,N_564);
nor U1367 (N_1367,N_720,N_318);
nand U1368 (N_1368,N_374,N_184);
and U1369 (N_1369,N_466,N_226);
and U1370 (N_1370,N_79,N_602);
and U1371 (N_1371,N_617,N_666);
or U1372 (N_1372,N_475,N_396);
and U1373 (N_1373,N_677,N_561);
and U1374 (N_1374,N_378,N_102);
or U1375 (N_1375,N_448,N_561);
or U1376 (N_1376,N_161,N_198);
and U1377 (N_1377,N_726,N_369);
nand U1378 (N_1378,N_254,N_58);
nor U1379 (N_1379,N_706,N_207);
or U1380 (N_1380,N_660,N_313);
and U1381 (N_1381,N_257,N_297);
and U1382 (N_1382,N_524,N_3);
and U1383 (N_1383,N_502,N_499);
nor U1384 (N_1384,N_183,N_458);
nor U1385 (N_1385,N_36,N_682);
or U1386 (N_1386,N_154,N_275);
and U1387 (N_1387,N_253,N_325);
and U1388 (N_1388,N_363,N_289);
and U1389 (N_1389,N_504,N_210);
nand U1390 (N_1390,N_520,N_731);
or U1391 (N_1391,N_289,N_455);
and U1392 (N_1392,N_655,N_636);
nor U1393 (N_1393,N_748,N_639);
nor U1394 (N_1394,N_702,N_633);
or U1395 (N_1395,N_362,N_22);
and U1396 (N_1396,N_629,N_651);
or U1397 (N_1397,N_228,N_460);
or U1398 (N_1398,N_6,N_461);
nor U1399 (N_1399,N_539,N_562);
nand U1400 (N_1400,N_418,N_728);
and U1401 (N_1401,N_149,N_444);
nand U1402 (N_1402,N_363,N_472);
and U1403 (N_1403,N_244,N_466);
nor U1404 (N_1404,N_401,N_15);
nand U1405 (N_1405,N_501,N_458);
or U1406 (N_1406,N_299,N_401);
and U1407 (N_1407,N_535,N_554);
nor U1408 (N_1408,N_86,N_26);
nor U1409 (N_1409,N_72,N_75);
nor U1410 (N_1410,N_128,N_275);
xnor U1411 (N_1411,N_181,N_443);
and U1412 (N_1412,N_0,N_91);
and U1413 (N_1413,N_63,N_465);
and U1414 (N_1414,N_427,N_10);
nand U1415 (N_1415,N_349,N_40);
nand U1416 (N_1416,N_456,N_327);
nand U1417 (N_1417,N_180,N_125);
nor U1418 (N_1418,N_280,N_586);
nor U1419 (N_1419,N_302,N_641);
and U1420 (N_1420,N_188,N_168);
nor U1421 (N_1421,N_568,N_495);
nand U1422 (N_1422,N_493,N_54);
nand U1423 (N_1423,N_377,N_274);
and U1424 (N_1424,N_647,N_459);
and U1425 (N_1425,N_645,N_509);
or U1426 (N_1426,N_655,N_36);
nor U1427 (N_1427,N_323,N_244);
or U1428 (N_1428,N_661,N_270);
or U1429 (N_1429,N_616,N_357);
and U1430 (N_1430,N_98,N_352);
or U1431 (N_1431,N_249,N_531);
nor U1432 (N_1432,N_95,N_266);
and U1433 (N_1433,N_25,N_370);
nor U1434 (N_1434,N_514,N_22);
nand U1435 (N_1435,N_572,N_247);
and U1436 (N_1436,N_206,N_196);
and U1437 (N_1437,N_189,N_629);
nand U1438 (N_1438,N_317,N_333);
or U1439 (N_1439,N_286,N_700);
nand U1440 (N_1440,N_201,N_596);
or U1441 (N_1441,N_421,N_160);
nor U1442 (N_1442,N_154,N_337);
and U1443 (N_1443,N_402,N_363);
and U1444 (N_1444,N_18,N_358);
nor U1445 (N_1445,N_488,N_122);
nor U1446 (N_1446,N_82,N_697);
and U1447 (N_1447,N_336,N_450);
or U1448 (N_1448,N_670,N_570);
nor U1449 (N_1449,N_243,N_177);
nor U1450 (N_1450,N_722,N_250);
nor U1451 (N_1451,N_41,N_356);
and U1452 (N_1452,N_141,N_255);
nor U1453 (N_1453,N_597,N_356);
and U1454 (N_1454,N_745,N_52);
nand U1455 (N_1455,N_25,N_463);
or U1456 (N_1456,N_689,N_741);
nand U1457 (N_1457,N_335,N_607);
or U1458 (N_1458,N_714,N_432);
or U1459 (N_1459,N_45,N_36);
and U1460 (N_1460,N_381,N_10);
nand U1461 (N_1461,N_101,N_91);
and U1462 (N_1462,N_150,N_302);
nor U1463 (N_1463,N_165,N_745);
and U1464 (N_1464,N_221,N_625);
nor U1465 (N_1465,N_42,N_204);
or U1466 (N_1466,N_718,N_651);
nor U1467 (N_1467,N_338,N_263);
and U1468 (N_1468,N_277,N_165);
or U1469 (N_1469,N_420,N_554);
and U1470 (N_1470,N_343,N_410);
nor U1471 (N_1471,N_339,N_144);
nor U1472 (N_1472,N_258,N_384);
nor U1473 (N_1473,N_521,N_642);
nor U1474 (N_1474,N_190,N_244);
nor U1475 (N_1475,N_644,N_479);
nor U1476 (N_1476,N_427,N_645);
or U1477 (N_1477,N_592,N_61);
or U1478 (N_1478,N_659,N_534);
and U1479 (N_1479,N_290,N_395);
and U1480 (N_1480,N_205,N_613);
and U1481 (N_1481,N_17,N_194);
nand U1482 (N_1482,N_278,N_15);
or U1483 (N_1483,N_114,N_497);
nand U1484 (N_1484,N_577,N_653);
or U1485 (N_1485,N_113,N_125);
nor U1486 (N_1486,N_232,N_18);
xnor U1487 (N_1487,N_224,N_409);
nand U1488 (N_1488,N_602,N_446);
or U1489 (N_1489,N_584,N_138);
nand U1490 (N_1490,N_171,N_310);
nor U1491 (N_1491,N_175,N_692);
and U1492 (N_1492,N_217,N_497);
nand U1493 (N_1493,N_358,N_281);
nor U1494 (N_1494,N_41,N_91);
and U1495 (N_1495,N_512,N_562);
and U1496 (N_1496,N_494,N_304);
and U1497 (N_1497,N_529,N_390);
and U1498 (N_1498,N_364,N_228);
nor U1499 (N_1499,N_660,N_161);
nand U1500 (N_1500,N_952,N_1331);
or U1501 (N_1501,N_1094,N_1200);
nand U1502 (N_1502,N_1190,N_1451);
or U1503 (N_1503,N_1147,N_984);
nand U1504 (N_1504,N_1436,N_1080);
nor U1505 (N_1505,N_802,N_1074);
nand U1506 (N_1506,N_983,N_1460);
nand U1507 (N_1507,N_1305,N_995);
or U1508 (N_1508,N_812,N_1426);
or U1509 (N_1509,N_845,N_1047);
nand U1510 (N_1510,N_835,N_969);
nor U1511 (N_1511,N_777,N_874);
nand U1512 (N_1512,N_1064,N_924);
nand U1513 (N_1513,N_1337,N_851);
nand U1514 (N_1514,N_914,N_1066);
or U1515 (N_1515,N_1497,N_904);
nand U1516 (N_1516,N_1093,N_973);
nand U1517 (N_1517,N_997,N_839);
and U1518 (N_1518,N_1007,N_1315);
or U1519 (N_1519,N_1281,N_1496);
or U1520 (N_1520,N_1117,N_1223);
xor U1521 (N_1521,N_1017,N_938);
nor U1522 (N_1522,N_1470,N_1052);
nor U1523 (N_1523,N_1078,N_1232);
and U1524 (N_1524,N_1151,N_1167);
nor U1525 (N_1525,N_963,N_1413);
and U1526 (N_1526,N_1224,N_1136);
and U1527 (N_1527,N_1448,N_1002);
and U1528 (N_1528,N_881,N_1242);
or U1529 (N_1529,N_1192,N_1063);
xor U1530 (N_1530,N_1272,N_1004);
nand U1531 (N_1531,N_987,N_1402);
or U1532 (N_1532,N_1444,N_836);
and U1533 (N_1533,N_822,N_1026);
and U1534 (N_1534,N_1209,N_1345);
nand U1535 (N_1535,N_1427,N_1018);
and U1536 (N_1536,N_915,N_1193);
nand U1537 (N_1537,N_813,N_1262);
and U1538 (N_1538,N_1457,N_1104);
and U1539 (N_1539,N_1067,N_853);
or U1540 (N_1540,N_1248,N_1332);
and U1541 (N_1541,N_1061,N_784);
nand U1542 (N_1542,N_1466,N_1022);
nor U1543 (N_1543,N_875,N_1241);
or U1544 (N_1544,N_787,N_1467);
or U1545 (N_1545,N_953,N_1035);
nor U1546 (N_1546,N_1418,N_1048);
and U1547 (N_1547,N_1082,N_872);
nand U1548 (N_1548,N_1255,N_1040);
nand U1549 (N_1549,N_1179,N_1428);
nor U1550 (N_1550,N_1180,N_1334);
nand U1551 (N_1551,N_1319,N_814);
or U1552 (N_1552,N_1073,N_1273);
nand U1553 (N_1553,N_794,N_1475);
and U1554 (N_1554,N_1172,N_1439);
or U1555 (N_1555,N_1422,N_1196);
nand U1556 (N_1556,N_1170,N_898);
and U1557 (N_1557,N_1020,N_1396);
nand U1558 (N_1558,N_951,N_1420);
nand U1559 (N_1559,N_950,N_1358);
or U1560 (N_1560,N_1181,N_1348);
nor U1561 (N_1561,N_1079,N_846);
xnor U1562 (N_1562,N_1154,N_764);
nand U1563 (N_1563,N_1363,N_935);
nor U1564 (N_1564,N_779,N_1355);
and U1565 (N_1565,N_1446,N_1398);
nor U1566 (N_1566,N_1060,N_1142);
and U1567 (N_1567,N_778,N_1031);
or U1568 (N_1568,N_797,N_1318);
nand U1569 (N_1569,N_1434,N_1486);
or U1570 (N_1570,N_1292,N_848);
nor U1571 (N_1571,N_1405,N_917);
nor U1572 (N_1572,N_1445,N_1127);
nand U1573 (N_1573,N_1086,N_838);
and U1574 (N_1574,N_1010,N_1473);
or U1575 (N_1575,N_801,N_913);
nand U1576 (N_1576,N_1263,N_966);
and U1577 (N_1577,N_1301,N_1347);
and U1578 (N_1578,N_830,N_1371);
and U1579 (N_1579,N_833,N_1099);
nor U1580 (N_1580,N_1354,N_1327);
or U1581 (N_1581,N_1085,N_768);
nand U1582 (N_1582,N_1478,N_1468);
nor U1583 (N_1583,N_970,N_1160);
and U1584 (N_1584,N_1210,N_923);
and U1585 (N_1585,N_781,N_971);
nor U1586 (N_1586,N_844,N_775);
and U1587 (N_1587,N_1175,N_1106);
or U1588 (N_1588,N_1032,N_1077);
nand U1589 (N_1589,N_1009,N_1463);
or U1590 (N_1590,N_1268,N_763);
xnor U1591 (N_1591,N_890,N_962);
nand U1592 (N_1592,N_1116,N_1430);
nand U1593 (N_1593,N_1366,N_885);
nand U1594 (N_1594,N_1459,N_1361);
and U1595 (N_1595,N_783,N_1295);
or U1596 (N_1596,N_1421,N_1050);
nand U1597 (N_1597,N_1286,N_1065);
nor U1598 (N_1598,N_829,N_1277);
nand U1599 (N_1599,N_903,N_1003);
or U1600 (N_1600,N_761,N_1051);
nor U1601 (N_1601,N_1177,N_807);
nand U1602 (N_1602,N_1499,N_1157);
and U1603 (N_1603,N_1492,N_1293);
nand U1604 (N_1604,N_1028,N_1222);
or U1605 (N_1605,N_918,N_873);
nor U1606 (N_1606,N_1495,N_1236);
xnor U1607 (N_1607,N_1344,N_1338);
nor U1608 (N_1608,N_799,N_926);
nand U1609 (N_1609,N_999,N_1280);
nand U1610 (N_1610,N_867,N_1137);
nor U1611 (N_1611,N_972,N_895);
nand U1612 (N_1612,N_1199,N_1424);
nand U1613 (N_1613,N_1414,N_1379);
and U1614 (N_1614,N_826,N_993);
nand U1615 (N_1615,N_1289,N_790);
xnor U1616 (N_1616,N_760,N_1226);
and U1617 (N_1617,N_896,N_1233);
nor U1618 (N_1618,N_905,N_868);
nor U1619 (N_1619,N_831,N_1215);
nor U1620 (N_1620,N_888,N_1055);
or U1621 (N_1621,N_916,N_1235);
or U1622 (N_1622,N_810,N_755);
nor U1623 (N_1623,N_1271,N_1118);
and U1624 (N_1624,N_1202,N_1034);
nor U1625 (N_1625,N_1423,N_1153);
and U1626 (N_1626,N_886,N_1163);
or U1627 (N_1627,N_1128,N_1364);
nand U1628 (N_1628,N_1217,N_1324);
or U1629 (N_1629,N_1244,N_1417);
nand U1630 (N_1630,N_908,N_1340);
or U1631 (N_1631,N_1493,N_823);
and U1632 (N_1632,N_1238,N_1432);
and U1633 (N_1633,N_1189,N_1112);
nor U1634 (N_1634,N_1419,N_765);
or U1635 (N_1635,N_1148,N_820);
nor U1636 (N_1636,N_1138,N_863);
and U1637 (N_1637,N_1351,N_1042);
nor U1638 (N_1638,N_1311,N_907);
xnor U1639 (N_1639,N_910,N_849);
nor U1640 (N_1640,N_850,N_1299);
or U1641 (N_1641,N_1382,N_1113);
nand U1642 (N_1642,N_1326,N_1015);
nor U1643 (N_1643,N_1485,N_1307);
nor U1644 (N_1644,N_1465,N_1229);
or U1645 (N_1645,N_782,N_1212);
nand U1646 (N_1646,N_988,N_1252);
nand U1647 (N_1647,N_1146,N_1266);
nor U1648 (N_1648,N_1440,N_1314);
and U1649 (N_1649,N_1494,N_1201);
nor U1650 (N_1650,N_1084,N_1464);
nand U1651 (N_1651,N_956,N_1247);
and U1652 (N_1652,N_865,N_791);
nor U1653 (N_1653,N_961,N_1365);
and U1654 (N_1654,N_759,N_939);
nand U1655 (N_1655,N_902,N_949);
nand U1656 (N_1656,N_1431,N_1208);
or U1657 (N_1657,N_841,N_1220);
or U1658 (N_1658,N_1110,N_1373);
nand U1659 (N_1659,N_1102,N_1105);
nand U1660 (N_1660,N_1474,N_1100);
nand U1661 (N_1661,N_1087,N_1412);
nand U1662 (N_1662,N_754,N_1168);
or U1663 (N_1663,N_1240,N_1409);
nand U1664 (N_1664,N_1033,N_1393);
nor U1665 (N_1665,N_780,N_818);
nand U1666 (N_1666,N_1498,N_751);
nand U1667 (N_1667,N_1343,N_1416);
or U1668 (N_1668,N_927,N_1243);
or U1669 (N_1669,N_1258,N_827);
nand U1670 (N_1670,N_1030,N_1141);
and U1671 (N_1671,N_1391,N_1390);
or U1672 (N_1672,N_1317,N_1225);
and U1673 (N_1673,N_1333,N_1049);
nand U1674 (N_1674,N_1452,N_1290);
or U1675 (N_1675,N_977,N_1041);
and U1676 (N_1676,N_756,N_870);
and U1677 (N_1677,N_1195,N_1429);
or U1678 (N_1678,N_1442,N_982);
and U1679 (N_1679,N_1198,N_842);
nand U1680 (N_1680,N_1069,N_1027);
nand U1681 (N_1681,N_941,N_933);
or U1682 (N_1682,N_1025,N_824);
and U1683 (N_1683,N_858,N_882);
or U1684 (N_1684,N_1265,N_1014);
and U1685 (N_1685,N_1090,N_1013);
or U1686 (N_1686,N_1375,N_1134);
and U1687 (N_1687,N_1058,N_1261);
nand U1688 (N_1688,N_1039,N_998);
nor U1689 (N_1689,N_1279,N_1339);
nor U1690 (N_1690,N_936,N_1166);
nand U1691 (N_1691,N_1288,N_1249);
or U1692 (N_1692,N_1120,N_1369);
nand U1693 (N_1693,N_1415,N_1231);
or U1694 (N_1694,N_1109,N_1384);
nand U1695 (N_1695,N_944,N_1346);
and U1696 (N_1696,N_1083,N_992);
or U1697 (N_1697,N_1159,N_1381);
and U1698 (N_1698,N_806,N_1152);
or U1699 (N_1699,N_1008,N_803);
and U1700 (N_1700,N_909,N_1021);
or U1701 (N_1701,N_1130,N_1045);
and U1702 (N_1702,N_1019,N_1400);
nand U1703 (N_1703,N_769,N_1095);
nor U1704 (N_1704,N_1135,N_1024);
nand U1705 (N_1705,N_832,N_1053);
nor U1706 (N_1706,N_1129,N_825);
nand U1707 (N_1707,N_1282,N_901);
and U1708 (N_1708,N_1389,N_837);
nor U1709 (N_1709,N_876,N_796);
or U1710 (N_1710,N_1378,N_789);
nor U1711 (N_1711,N_860,N_1367);
and U1712 (N_1712,N_1296,N_1435);
nand U1713 (N_1713,N_922,N_1246);
nand U1714 (N_1714,N_1205,N_854);
nor U1715 (N_1715,N_1313,N_1219);
and U1716 (N_1716,N_1174,N_800);
or U1717 (N_1717,N_792,N_1088);
and U1718 (N_1718,N_1036,N_1254);
nand U1719 (N_1719,N_1122,N_1075);
nor U1720 (N_1720,N_1211,N_1139);
and U1721 (N_1721,N_847,N_1357);
or U1722 (N_1722,N_1483,N_1479);
and U1723 (N_1723,N_1325,N_889);
or U1724 (N_1724,N_1089,N_991);
nand U1725 (N_1725,N_1191,N_1029);
or U1726 (N_1726,N_1230,N_967);
nor U1727 (N_1727,N_834,N_840);
or U1728 (N_1728,N_1490,N_1161);
nor U1729 (N_1729,N_1316,N_1341);
nand U1730 (N_1730,N_774,N_1356);
or U1731 (N_1731,N_980,N_883);
and U1732 (N_1732,N_857,N_866);
nor U1733 (N_1733,N_1385,N_1359);
or U1734 (N_1734,N_1336,N_968);
and U1735 (N_1735,N_1171,N_1342);
and U1736 (N_1736,N_1162,N_1216);
or U1737 (N_1737,N_762,N_862);
nand U1738 (N_1738,N_1491,N_1449);
nand U1739 (N_1739,N_1114,N_1126);
or U1740 (N_1740,N_1488,N_1387);
and U1741 (N_1741,N_1309,N_1443);
or U1742 (N_1742,N_1000,N_1329);
and U1743 (N_1743,N_1006,N_1441);
nor U1744 (N_1744,N_752,N_957);
and U1745 (N_1745,N_788,N_1267);
nor U1746 (N_1746,N_1044,N_1383);
nand U1747 (N_1747,N_819,N_1370);
nor U1748 (N_1748,N_1407,N_1098);
or U1749 (N_1749,N_1253,N_976);
nor U1750 (N_1750,N_1111,N_805);
nor U1751 (N_1751,N_809,N_1182);
nand U1752 (N_1752,N_1203,N_911);
nor U1753 (N_1753,N_1057,N_1304);
nor U1754 (N_1754,N_1092,N_1455);
nor U1755 (N_1755,N_1143,N_795);
nor U1756 (N_1756,N_981,N_1016);
or U1757 (N_1757,N_852,N_928);
or U1758 (N_1758,N_1257,N_1096);
and U1759 (N_1759,N_887,N_1227);
nor U1760 (N_1760,N_1321,N_900);
or U1761 (N_1761,N_856,N_1425);
nor U1762 (N_1762,N_1185,N_1251);
and U1763 (N_1763,N_942,N_815);
or U1764 (N_1764,N_1071,N_932);
nand U1765 (N_1765,N_1276,N_1308);
nand U1766 (N_1766,N_1300,N_793);
nor U1767 (N_1767,N_1294,N_1350);
and U1768 (N_1768,N_1453,N_1204);
nor U1769 (N_1769,N_871,N_1368);
or U1770 (N_1770,N_985,N_1264);
nor U1771 (N_1771,N_947,N_864);
nand U1772 (N_1772,N_1269,N_1081);
nor U1773 (N_1773,N_859,N_1132);
nor U1774 (N_1774,N_1218,N_943);
nand U1775 (N_1775,N_877,N_1176);
nand U1776 (N_1776,N_1103,N_897);
or U1777 (N_1777,N_1107,N_1458);
or U1778 (N_1778,N_808,N_974);
and U1779 (N_1779,N_894,N_1270);
and U1780 (N_1780,N_1234,N_1076);
and U1781 (N_1781,N_1477,N_878);
and U1782 (N_1782,N_1438,N_1484);
nand U1783 (N_1783,N_1140,N_828);
nand U1784 (N_1784,N_1186,N_1395);
nand U1785 (N_1785,N_1433,N_978);
nor U1786 (N_1786,N_1011,N_1149);
nor U1787 (N_1787,N_773,N_1437);
and U1788 (N_1788,N_1188,N_869);
or U1789 (N_1789,N_1194,N_785);
and U1790 (N_1790,N_816,N_945);
nand U1791 (N_1791,N_770,N_958);
and U1792 (N_1792,N_1133,N_861);
xor U1793 (N_1793,N_798,N_1068);
xnor U1794 (N_1794,N_1310,N_1376);
or U1795 (N_1795,N_929,N_1392);
nand U1796 (N_1796,N_879,N_1183);
nor U1797 (N_1797,N_1256,N_1169);
and U1798 (N_1798,N_1097,N_946);
and U1799 (N_1799,N_1353,N_1214);
or U1800 (N_1800,N_1377,N_1323);
nor U1801 (N_1801,N_1408,N_1245);
and U1802 (N_1802,N_1125,N_1487);
nand U1803 (N_1803,N_1173,N_906);
nand U1804 (N_1804,N_811,N_1285);
and U1805 (N_1805,N_1306,N_937);
and U1806 (N_1806,N_1360,N_1388);
or U1807 (N_1807,N_753,N_1207);
or U1808 (N_1808,N_1283,N_1164);
xnor U1809 (N_1809,N_1322,N_1394);
and U1810 (N_1810,N_1312,N_920);
nor U1811 (N_1811,N_1101,N_1119);
or U1812 (N_1812,N_1476,N_964);
xnor U1813 (N_1813,N_1228,N_1091);
or U1814 (N_1814,N_750,N_1397);
nor U1815 (N_1815,N_979,N_921);
and U1816 (N_1816,N_1237,N_1482);
and U1817 (N_1817,N_1178,N_1144);
and U1818 (N_1818,N_959,N_960);
xor U1819 (N_1819,N_1274,N_1275);
nor U1820 (N_1820,N_1362,N_994);
and U1821 (N_1821,N_934,N_1297);
and U1822 (N_1822,N_1335,N_975);
nor U1823 (N_1823,N_1206,N_1038);
nor U1824 (N_1824,N_1037,N_1291);
nand U1825 (N_1825,N_1352,N_1404);
or U1826 (N_1826,N_821,N_1070);
or U1827 (N_1827,N_1043,N_1150);
nor U1828 (N_1828,N_1123,N_1399);
and U1829 (N_1829,N_1456,N_1062);
or U1830 (N_1830,N_1259,N_843);
or U1831 (N_1831,N_1287,N_1046);
and U1832 (N_1832,N_1481,N_1410);
or U1833 (N_1833,N_1330,N_954);
nor U1834 (N_1834,N_766,N_1320);
and U1835 (N_1835,N_1374,N_1184);
nor U1836 (N_1836,N_1001,N_1213);
or U1837 (N_1837,N_948,N_1469);
nor U1838 (N_1838,N_1303,N_1328);
or U1839 (N_1839,N_1489,N_767);
and U1840 (N_1840,N_1450,N_1165);
and U1841 (N_1841,N_912,N_1386);
nand U1842 (N_1842,N_1298,N_1221);
and U1843 (N_1843,N_1005,N_1012);
or U1844 (N_1844,N_1124,N_1250);
or U1845 (N_1845,N_1349,N_1145);
xnor U1846 (N_1846,N_893,N_771);
nand U1847 (N_1847,N_1461,N_965);
and U1848 (N_1848,N_1372,N_1472);
nand U1849 (N_1849,N_919,N_989);
nor U1850 (N_1850,N_1197,N_1454);
nand U1851 (N_1851,N_891,N_817);
and U1852 (N_1852,N_1471,N_996);
or U1853 (N_1853,N_892,N_931);
nor U1854 (N_1854,N_1302,N_986);
nor U1855 (N_1855,N_1023,N_884);
nor U1856 (N_1856,N_776,N_758);
nor U1857 (N_1857,N_1187,N_1054);
or U1858 (N_1858,N_1406,N_1155);
nor U1859 (N_1859,N_804,N_786);
nor U1860 (N_1860,N_1278,N_1284);
nand U1861 (N_1861,N_1072,N_1480);
nand U1862 (N_1862,N_1059,N_1108);
nand U1863 (N_1863,N_955,N_990);
and U1864 (N_1864,N_1131,N_940);
and U1865 (N_1865,N_880,N_1156);
and U1866 (N_1866,N_1403,N_1239);
nand U1867 (N_1867,N_1447,N_1158);
xnor U1868 (N_1868,N_855,N_1115);
and U1869 (N_1869,N_772,N_1121);
nand U1870 (N_1870,N_1260,N_925);
nand U1871 (N_1871,N_899,N_1380);
or U1872 (N_1872,N_1411,N_1401);
nand U1873 (N_1873,N_1462,N_1056);
nand U1874 (N_1874,N_757,N_930);
nor U1875 (N_1875,N_767,N_802);
nor U1876 (N_1876,N_1183,N_797);
nor U1877 (N_1877,N_1356,N_917);
and U1878 (N_1878,N_1147,N_863);
or U1879 (N_1879,N_1394,N_900);
or U1880 (N_1880,N_1122,N_1024);
nand U1881 (N_1881,N_1245,N_940);
and U1882 (N_1882,N_1336,N_1184);
nor U1883 (N_1883,N_1216,N_992);
or U1884 (N_1884,N_1347,N_1217);
and U1885 (N_1885,N_1264,N_1254);
nand U1886 (N_1886,N_1469,N_1103);
nor U1887 (N_1887,N_1301,N_1208);
or U1888 (N_1888,N_772,N_1268);
and U1889 (N_1889,N_801,N_972);
nand U1890 (N_1890,N_1365,N_1089);
or U1891 (N_1891,N_1268,N_1476);
and U1892 (N_1892,N_1391,N_1148);
nor U1893 (N_1893,N_1145,N_1379);
or U1894 (N_1894,N_1019,N_950);
and U1895 (N_1895,N_1143,N_1315);
or U1896 (N_1896,N_891,N_755);
and U1897 (N_1897,N_1164,N_879);
or U1898 (N_1898,N_874,N_926);
and U1899 (N_1899,N_1298,N_1291);
nand U1900 (N_1900,N_1155,N_953);
nand U1901 (N_1901,N_1239,N_1117);
nor U1902 (N_1902,N_1320,N_1467);
or U1903 (N_1903,N_1144,N_1005);
nor U1904 (N_1904,N_986,N_1416);
or U1905 (N_1905,N_931,N_989);
or U1906 (N_1906,N_1187,N_1000);
nor U1907 (N_1907,N_1239,N_1031);
nand U1908 (N_1908,N_923,N_1297);
nor U1909 (N_1909,N_1498,N_905);
and U1910 (N_1910,N_1277,N_1133);
nor U1911 (N_1911,N_1308,N_1080);
nand U1912 (N_1912,N_928,N_890);
and U1913 (N_1913,N_952,N_949);
or U1914 (N_1914,N_784,N_1156);
and U1915 (N_1915,N_999,N_1045);
and U1916 (N_1916,N_1199,N_874);
nor U1917 (N_1917,N_1339,N_1475);
or U1918 (N_1918,N_1337,N_1307);
and U1919 (N_1919,N_804,N_913);
nor U1920 (N_1920,N_1044,N_1157);
nand U1921 (N_1921,N_1141,N_1043);
nor U1922 (N_1922,N_1450,N_1473);
nand U1923 (N_1923,N_867,N_1479);
nand U1924 (N_1924,N_920,N_876);
nor U1925 (N_1925,N_1420,N_997);
nor U1926 (N_1926,N_969,N_1319);
nor U1927 (N_1927,N_1303,N_1175);
or U1928 (N_1928,N_1000,N_1001);
nand U1929 (N_1929,N_1235,N_1132);
nand U1930 (N_1930,N_1464,N_1478);
and U1931 (N_1931,N_1482,N_1492);
or U1932 (N_1932,N_1339,N_1416);
nand U1933 (N_1933,N_928,N_1293);
nand U1934 (N_1934,N_1071,N_1145);
nand U1935 (N_1935,N_1014,N_1489);
and U1936 (N_1936,N_1214,N_1428);
or U1937 (N_1937,N_1382,N_758);
and U1938 (N_1938,N_1433,N_1093);
nand U1939 (N_1939,N_1323,N_1139);
or U1940 (N_1940,N_1113,N_1143);
or U1941 (N_1941,N_995,N_970);
or U1942 (N_1942,N_957,N_1020);
or U1943 (N_1943,N_810,N_1492);
or U1944 (N_1944,N_832,N_1257);
or U1945 (N_1945,N_751,N_1047);
or U1946 (N_1946,N_852,N_1017);
nor U1947 (N_1947,N_893,N_1232);
and U1948 (N_1948,N_1195,N_791);
nor U1949 (N_1949,N_1003,N_883);
nand U1950 (N_1950,N_1100,N_815);
nor U1951 (N_1951,N_761,N_1353);
nand U1952 (N_1952,N_1346,N_1292);
and U1953 (N_1953,N_1346,N_1477);
and U1954 (N_1954,N_1026,N_1350);
nand U1955 (N_1955,N_933,N_1114);
or U1956 (N_1956,N_1444,N_1174);
or U1957 (N_1957,N_1276,N_978);
or U1958 (N_1958,N_1218,N_820);
nor U1959 (N_1959,N_1491,N_1366);
nand U1960 (N_1960,N_1142,N_1027);
and U1961 (N_1961,N_938,N_1272);
and U1962 (N_1962,N_983,N_1050);
and U1963 (N_1963,N_1207,N_1006);
nor U1964 (N_1964,N_838,N_1335);
and U1965 (N_1965,N_804,N_880);
or U1966 (N_1966,N_1380,N_1193);
and U1967 (N_1967,N_1326,N_1443);
nor U1968 (N_1968,N_1225,N_1183);
nand U1969 (N_1969,N_1452,N_1408);
or U1970 (N_1970,N_1362,N_1121);
xnor U1971 (N_1971,N_1095,N_1168);
or U1972 (N_1972,N_937,N_1266);
nand U1973 (N_1973,N_1399,N_851);
or U1974 (N_1974,N_874,N_1128);
nor U1975 (N_1975,N_1005,N_808);
xnor U1976 (N_1976,N_1259,N_790);
or U1977 (N_1977,N_870,N_1147);
nor U1978 (N_1978,N_1118,N_815);
and U1979 (N_1979,N_1431,N_1403);
or U1980 (N_1980,N_1114,N_832);
nor U1981 (N_1981,N_991,N_809);
or U1982 (N_1982,N_966,N_1323);
nand U1983 (N_1983,N_1160,N_960);
nor U1984 (N_1984,N_1308,N_972);
xnor U1985 (N_1985,N_757,N_1399);
or U1986 (N_1986,N_1249,N_1323);
nand U1987 (N_1987,N_1133,N_1332);
nand U1988 (N_1988,N_780,N_1406);
and U1989 (N_1989,N_940,N_1160);
and U1990 (N_1990,N_1260,N_1398);
nor U1991 (N_1991,N_1487,N_922);
nand U1992 (N_1992,N_1138,N_1395);
nor U1993 (N_1993,N_971,N_1345);
nor U1994 (N_1994,N_1255,N_824);
nand U1995 (N_1995,N_958,N_1235);
nor U1996 (N_1996,N_819,N_1349);
and U1997 (N_1997,N_1096,N_1114);
or U1998 (N_1998,N_1140,N_963);
and U1999 (N_1999,N_930,N_1341);
or U2000 (N_2000,N_1081,N_1000);
nand U2001 (N_2001,N_756,N_866);
nor U2002 (N_2002,N_930,N_1195);
and U2003 (N_2003,N_1415,N_1401);
or U2004 (N_2004,N_1094,N_1191);
and U2005 (N_2005,N_1107,N_986);
and U2006 (N_2006,N_947,N_1433);
nor U2007 (N_2007,N_1156,N_1387);
or U2008 (N_2008,N_1118,N_1135);
nor U2009 (N_2009,N_1428,N_872);
and U2010 (N_2010,N_1281,N_942);
or U2011 (N_2011,N_924,N_1217);
nor U2012 (N_2012,N_1343,N_1475);
or U2013 (N_2013,N_996,N_915);
or U2014 (N_2014,N_910,N_1321);
nor U2015 (N_2015,N_1315,N_800);
nor U2016 (N_2016,N_1394,N_909);
or U2017 (N_2017,N_1459,N_1495);
or U2018 (N_2018,N_753,N_1355);
nor U2019 (N_2019,N_1020,N_912);
or U2020 (N_2020,N_1049,N_786);
or U2021 (N_2021,N_1220,N_834);
nand U2022 (N_2022,N_786,N_918);
or U2023 (N_2023,N_1343,N_967);
nor U2024 (N_2024,N_954,N_1401);
or U2025 (N_2025,N_845,N_967);
nor U2026 (N_2026,N_1076,N_1368);
or U2027 (N_2027,N_1360,N_1343);
and U2028 (N_2028,N_1462,N_1232);
and U2029 (N_2029,N_965,N_864);
or U2030 (N_2030,N_1248,N_855);
nor U2031 (N_2031,N_1383,N_826);
nand U2032 (N_2032,N_785,N_1131);
and U2033 (N_2033,N_1277,N_760);
nor U2034 (N_2034,N_760,N_1211);
and U2035 (N_2035,N_1348,N_975);
nor U2036 (N_2036,N_975,N_992);
or U2037 (N_2037,N_762,N_984);
and U2038 (N_2038,N_905,N_1451);
and U2039 (N_2039,N_993,N_1151);
nand U2040 (N_2040,N_753,N_837);
nand U2041 (N_2041,N_1401,N_843);
and U2042 (N_2042,N_1373,N_1017);
or U2043 (N_2043,N_1367,N_967);
nand U2044 (N_2044,N_1091,N_1423);
or U2045 (N_2045,N_1039,N_1012);
nor U2046 (N_2046,N_1231,N_1206);
nor U2047 (N_2047,N_985,N_1233);
nand U2048 (N_2048,N_1192,N_773);
or U2049 (N_2049,N_1335,N_1314);
nand U2050 (N_2050,N_1402,N_1469);
and U2051 (N_2051,N_1249,N_775);
nor U2052 (N_2052,N_1178,N_809);
or U2053 (N_2053,N_1492,N_1047);
or U2054 (N_2054,N_1348,N_1215);
nor U2055 (N_2055,N_1269,N_1354);
or U2056 (N_2056,N_1246,N_828);
nand U2057 (N_2057,N_994,N_757);
nor U2058 (N_2058,N_1175,N_1339);
nand U2059 (N_2059,N_1021,N_1438);
nor U2060 (N_2060,N_1286,N_1281);
and U2061 (N_2061,N_1094,N_1272);
and U2062 (N_2062,N_1026,N_826);
nor U2063 (N_2063,N_1052,N_1173);
and U2064 (N_2064,N_1398,N_1348);
and U2065 (N_2065,N_1054,N_1248);
nor U2066 (N_2066,N_1414,N_771);
and U2067 (N_2067,N_776,N_892);
and U2068 (N_2068,N_1169,N_1005);
and U2069 (N_2069,N_1172,N_804);
and U2070 (N_2070,N_773,N_994);
or U2071 (N_2071,N_1457,N_1077);
nor U2072 (N_2072,N_967,N_908);
or U2073 (N_2073,N_1245,N_1111);
or U2074 (N_2074,N_1434,N_1034);
or U2075 (N_2075,N_1361,N_789);
nand U2076 (N_2076,N_1086,N_1056);
or U2077 (N_2077,N_1240,N_920);
and U2078 (N_2078,N_1337,N_921);
nor U2079 (N_2079,N_1403,N_1059);
or U2080 (N_2080,N_879,N_1196);
and U2081 (N_2081,N_1493,N_1038);
nor U2082 (N_2082,N_1289,N_1255);
and U2083 (N_2083,N_898,N_1359);
and U2084 (N_2084,N_1451,N_1011);
or U2085 (N_2085,N_1162,N_1035);
nor U2086 (N_2086,N_1491,N_1271);
or U2087 (N_2087,N_1414,N_1152);
nor U2088 (N_2088,N_860,N_881);
or U2089 (N_2089,N_1009,N_1200);
or U2090 (N_2090,N_949,N_1257);
or U2091 (N_2091,N_790,N_1192);
and U2092 (N_2092,N_1383,N_1032);
nand U2093 (N_2093,N_1088,N_1367);
and U2094 (N_2094,N_1236,N_1375);
nand U2095 (N_2095,N_769,N_1207);
and U2096 (N_2096,N_1430,N_865);
nand U2097 (N_2097,N_1455,N_952);
and U2098 (N_2098,N_999,N_1418);
nor U2099 (N_2099,N_1457,N_1474);
nand U2100 (N_2100,N_755,N_859);
xnor U2101 (N_2101,N_794,N_994);
nand U2102 (N_2102,N_1398,N_1285);
and U2103 (N_2103,N_954,N_1412);
xnor U2104 (N_2104,N_1461,N_865);
nand U2105 (N_2105,N_882,N_972);
and U2106 (N_2106,N_1260,N_924);
and U2107 (N_2107,N_1315,N_1075);
and U2108 (N_2108,N_1430,N_973);
nor U2109 (N_2109,N_831,N_835);
nor U2110 (N_2110,N_1469,N_1446);
nor U2111 (N_2111,N_892,N_783);
nor U2112 (N_2112,N_1389,N_1274);
or U2113 (N_2113,N_1122,N_1399);
xor U2114 (N_2114,N_1254,N_1239);
nor U2115 (N_2115,N_1496,N_829);
and U2116 (N_2116,N_808,N_867);
or U2117 (N_2117,N_1454,N_858);
and U2118 (N_2118,N_1488,N_1070);
nor U2119 (N_2119,N_976,N_874);
or U2120 (N_2120,N_1194,N_936);
and U2121 (N_2121,N_1035,N_1145);
nor U2122 (N_2122,N_844,N_965);
and U2123 (N_2123,N_837,N_1361);
nor U2124 (N_2124,N_967,N_926);
nand U2125 (N_2125,N_882,N_1059);
nor U2126 (N_2126,N_1478,N_1004);
or U2127 (N_2127,N_860,N_1013);
or U2128 (N_2128,N_1218,N_970);
nand U2129 (N_2129,N_1327,N_1181);
nor U2130 (N_2130,N_1132,N_775);
and U2131 (N_2131,N_1291,N_1355);
nand U2132 (N_2132,N_770,N_1310);
or U2133 (N_2133,N_874,N_1460);
nand U2134 (N_2134,N_1443,N_1424);
or U2135 (N_2135,N_1320,N_1160);
or U2136 (N_2136,N_782,N_1155);
or U2137 (N_2137,N_1472,N_804);
nor U2138 (N_2138,N_1077,N_827);
or U2139 (N_2139,N_1069,N_1173);
or U2140 (N_2140,N_1194,N_1200);
nor U2141 (N_2141,N_1404,N_949);
and U2142 (N_2142,N_776,N_890);
nand U2143 (N_2143,N_1218,N_946);
nand U2144 (N_2144,N_926,N_1027);
nor U2145 (N_2145,N_929,N_806);
or U2146 (N_2146,N_1022,N_1155);
or U2147 (N_2147,N_1333,N_985);
or U2148 (N_2148,N_1152,N_1427);
or U2149 (N_2149,N_1377,N_755);
or U2150 (N_2150,N_904,N_909);
or U2151 (N_2151,N_1071,N_945);
and U2152 (N_2152,N_1280,N_1245);
nor U2153 (N_2153,N_1213,N_885);
or U2154 (N_2154,N_957,N_834);
nand U2155 (N_2155,N_1234,N_1059);
nor U2156 (N_2156,N_784,N_935);
and U2157 (N_2157,N_1329,N_1232);
nand U2158 (N_2158,N_860,N_1447);
nor U2159 (N_2159,N_1320,N_1255);
and U2160 (N_2160,N_966,N_847);
or U2161 (N_2161,N_788,N_822);
or U2162 (N_2162,N_1496,N_1298);
nand U2163 (N_2163,N_963,N_1131);
nand U2164 (N_2164,N_913,N_996);
nand U2165 (N_2165,N_1036,N_1284);
nand U2166 (N_2166,N_1065,N_760);
nand U2167 (N_2167,N_992,N_1101);
and U2168 (N_2168,N_1327,N_1217);
and U2169 (N_2169,N_1073,N_980);
xnor U2170 (N_2170,N_971,N_1367);
and U2171 (N_2171,N_1042,N_1345);
nand U2172 (N_2172,N_1174,N_973);
nand U2173 (N_2173,N_857,N_758);
nand U2174 (N_2174,N_1401,N_1467);
nand U2175 (N_2175,N_1266,N_1025);
nand U2176 (N_2176,N_1268,N_829);
and U2177 (N_2177,N_1326,N_1327);
nand U2178 (N_2178,N_852,N_1204);
nor U2179 (N_2179,N_1228,N_1380);
and U2180 (N_2180,N_1176,N_975);
nor U2181 (N_2181,N_1014,N_1417);
or U2182 (N_2182,N_1097,N_985);
or U2183 (N_2183,N_897,N_1312);
nor U2184 (N_2184,N_1260,N_1232);
and U2185 (N_2185,N_824,N_1179);
or U2186 (N_2186,N_830,N_858);
and U2187 (N_2187,N_1140,N_1351);
or U2188 (N_2188,N_1191,N_1260);
and U2189 (N_2189,N_1347,N_1174);
or U2190 (N_2190,N_1038,N_978);
and U2191 (N_2191,N_1420,N_1463);
and U2192 (N_2192,N_1044,N_1422);
and U2193 (N_2193,N_1395,N_1196);
nor U2194 (N_2194,N_916,N_1312);
nor U2195 (N_2195,N_1037,N_1446);
and U2196 (N_2196,N_1312,N_967);
or U2197 (N_2197,N_1191,N_881);
and U2198 (N_2198,N_1070,N_877);
nand U2199 (N_2199,N_1054,N_817);
or U2200 (N_2200,N_1113,N_855);
or U2201 (N_2201,N_1257,N_1240);
or U2202 (N_2202,N_1293,N_1299);
nand U2203 (N_2203,N_750,N_1315);
nor U2204 (N_2204,N_1013,N_832);
nand U2205 (N_2205,N_1467,N_1042);
nand U2206 (N_2206,N_1100,N_1296);
nor U2207 (N_2207,N_1225,N_1280);
nand U2208 (N_2208,N_982,N_1069);
nor U2209 (N_2209,N_1205,N_1435);
nand U2210 (N_2210,N_1428,N_833);
or U2211 (N_2211,N_911,N_1191);
or U2212 (N_2212,N_883,N_1196);
nor U2213 (N_2213,N_1021,N_816);
and U2214 (N_2214,N_1252,N_943);
or U2215 (N_2215,N_816,N_1002);
and U2216 (N_2216,N_1197,N_758);
and U2217 (N_2217,N_879,N_833);
and U2218 (N_2218,N_1169,N_1286);
and U2219 (N_2219,N_818,N_1379);
nand U2220 (N_2220,N_1180,N_865);
nand U2221 (N_2221,N_1417,N_1300);
and U2222 (N_2222,N_1428,N_1106);
nand U2223 (N_2223,N_935,N_1211);
nor U2224 (N_2224,N_825,N_1131);
nand U2225 (N_2225,N_1162,N_1384);
nand U2226 (N_2226,N_1347,N_883);
nand U2227 (N_2227,N_961,N_770);
nand U2228 (N_2228,N_935,N_1161);
nor U2229 (N_2229,N_798,N_1154);
nand U2230 (N_2230,N_811,N_1399);
or U2231 (N_2231,N_1050,N_893);
or U2232 (N_2232,N_1036,N_1056);
or U2233 (N_2233,N_1016,N_1329);
nand U2234 (N_2234,N_1279,N_768);
and U2235 (N_2235,N_830,N_841);
and U2236 (N_2236,N_1422,N_945);
nor U2237 (N_2237,N_1117,N_1236);
nor U2238 (N_2238,N_810,N_1199);
nand U2239 (N_2239,N_886,N_1438);
nand U2240 (N_2240,N_864,N_841);
nor U2241 (N_2241,N_1087,N_1304);
nand U2242 (N_2242,N_759,N_1282);
and U2243 (N_2243,N_808,N_1353);
nand U2244 (N_2244,N_990,N_1295);
or U2245 (N_2245,N_1118,N_1078);
nor U2246 (N_2246,N_1468,N_1284);
nor U2247 (N_2247,N_857,N_1343);
or U2248 (N_2248,N_1133,N_881);
or U2249 (N_2249,N_1460,N_852);
nor U2250 (N_2250,N_2048,N_1928);
nand U2251 (N_2251,N_2154,N_2167);
or U2252 (N_2252,N_1921,N_1787);
or U2253 (N_2253,N_1820,N_1797);
and U2254 (N_2254,N_1707,N_1557);
nor U2255 (N_2255,N_1728,N_2164);
or U2256 (N_2256,N_1576,N_2039);
nor U2257 (N_2257,N_2098,N_1609);
and U2258 (N_2258,N_1503,N_1941);
and U2259 (N_2259,N_2020,N_2058);
nand U2260 (N_2260,N_1993,N_1681);
nand U2261 (N_2261,N_1760,N_1960);
and U2262 (N_2262,N_1507,N_2231);
nand U2263 (N_2263,N_2147,N_1834);
nor U2264 (N_2264,N_2008,N_1781);
nor U2265 (N_2265,N_2171,N_1958);
nor U2266 (N_2266,N_2000,N_1725);
nor U2267 (N_2267,N_1513,N_1790);
and U2268 (N_2268,N_2223,N_1726);
and U2269 (N_2269,N_2091,N_1506);
nand U2270 (N_2270,N_1929,N_2036);
nand U2271 (N_2271,N_1897,N_2029);
nor U2272 (N_2272,N_1908,N_2001);
nor U2273 (N_2273,N_1989,N_2022);
nand U2274 (N_2274,N_1625,N_1717);
nor U2275 (N_2275,N_1919,N_2193);
nand U2276 (N_2276,N_1865,N_2227);
or U2277 (N_2277,N_1589,N_2212);
and U2278 (N_2278,N_2187,N_1679);
nand U2279 (N_2279,N_1899,N_1955);
nor U2280 (N_2280,N_1676,N_1549);
nand U2281 (N_2281,N_1501,N_1827);
nand U2282 (N_2282,N_1887,N_1907);
nor U2283 (N_2283,N_2120,N_1923);
or U2284 (N_2284,N_1977,N_1836);
and U2285 (N_2285,N_2135,N_2180);
nand U2286 (N_2286,N_1691,N_2224);
nor U2287 (N_2287,N_1646,N_1697);
or U2288 (N_2288,N_2159,N_1937);
nand U2289 (N_2289,N_2086,N_1532);
and U2290 (N_2290,N_1823,N_1537);
nor U2291 (N_2291,N_1565,N_1940);
or U2292 (N_2292,N_1570,N_1519);
nor U2293 (N_2293,N_2084,N_1642);
nor U2294 (N_2294,N_2109,N_1508);
or U2295 (N_2295,N_1879,N_1620);
and U2296 (N_2296,N_1866,N_1604);
or U2297 (N_2297,N_2133,N_1848);
and U2298 (N_2298,N_1802,N_1975);
or U2299 (N_2299,N_2131,N_1674);
or U2300 (N_2300,N_1767,N_2249);
nand U2301 (N_2301,N_1762,N_1988);
nand U2302 (N_2302,N_1952,N_2148);
or U2303 (N_2303,N_1886,N_1894);
and U2304 (N_2304,N_1706,N_1687);
nand U2305 (N_2305,N_1774,N_1518);
nor U2306 (N_2306,N_2194,N_1883);
nand U2307 (N_2307,N_1754,N_2181);
or U2308 (N_2308,N_2096,N_1548);
nand U2309 (N_2309,N_1577,N_1590);
nand U2310 (N_2310,N_1660,N_1587);
nor U2311 (N_2311,N_2178,N_1520);
nand U2312 (N_2312,N_1749,N_1634);
and U2313 (N_2313,N_1619,N_1505);
nor U2314 (N_2314,N_1873,N_1632);
and U2315 (N_2315,N_1949,N_1595);
nor U2316 (N_2316,N_1739,N_1543);
or U2317 (N_2317,N_1920,N_1771);
or U2318 (N_2318,N_1735,N_1740);
nand U2319 (N_2319,N_2248,N_1965);
nand U2320 (N_2320,N_2151,N_1708);
nand U2321 (N_2321,N_1715,N_1581);
or U2322 (N_2322,N_1611,N_1869);
nor U2323 (N_2323,N_2215,N_1963);
nor U2324 (N_2324,N_1783,N_1636);
or U2325 (N_2325,N_1773,N_1968);
and U2326 (N_2326,N_2114,N_1562);
nor U2327 (N_2327,N_1500,N_1881);
and U2328 (N_2328,N_1545,N_1554);
or U2329 (N_2329,N_1889,N_2002);
nand U2330 (N_2330,N_1525,N_1580);
nand U2331 (N_2331,N_1526,N_2014);
nand U2332 (N_2332,N_1705,N_1840);
xnor U2333 (N_2333,N_2204,N_2024);
or U2334 (N_2334,N_2129,N_1682);
nor U2335 (N_2335,N_1649,N_2240);
nand U2336 (N_2336,N_1806,N_2234);
and U2337 (N_2337,N_2182,N_2030);
nor U2338 (N_2338,N_2192,N_2044);
nand U2339 (N_2339,N_2062,N_2214);
or U2340 (N_2340,N_1668,N_1597);
and U2341 (N_2341,N_2064,N_1523);
and U2342 (N_2342,N_1855,N_1571);
and U2343 (N_2343,N_1807,N_1981);
or U2344 (N_2344,N_1901,N_1775);
and U2345 (N_2345,N_1838,N_1947);
and U2346 (N_2346,N_1568,N_1934);
or U2347 (N_2347,N_1831,N_1716);
nor U2348 (N_2348,N_2207,N_2203);
nor U2349 (N_2349,N_1942,N_1566);
nand U2350 (N_2350,N_2051,N_1796);
and U2351 (N_2351,N_1612,N_1556);
or U2352 (N_2352,N_2186,N_2222);
nor U2353 (N_2353,N_2169,N_2026);
or U2354 (N_2354,N_1585,N_1751);
and U2355 (N_2355,N_1527,N_1885);
and U2356 (N_2356,N_1995,N_1644);
and U2357 (N_2357,N_1758,N_2218);
nor U2358 (N_2358,N_1786,N_1986);
nor U2359 (N_2359,N_1969,N_1628);
nor U2360 (N_2360,N_2225,N_1766);
nand U2361 (N_2361,N_2093,N_1584);
and U2362 (N_2362,N_1791,N_1623);
xor U2363 (N_2363,N_1524,N_1509);
nand U2364 (N_2364,N_1748,N_1677);
and U2365 (N_2365,N_1666,N_1852);
and U2366 (N_2366,N_2208,N_2177);
or U2367 (N_2367,N_1910,N_2073);
nor U2368 (N_2368,N_1756,N_2195);
xnor U2369 (N_2369,N_1645,N_1872);
nor U2370 (N_2370,N_1830,N_2099);
or U2371 (N_2371,N_1882,N_2111);
and U2372 (N_2372,N_1712,N_1971);
nor U2373 (N_2373,N_2165,N_2142);
nand U2374 (N_2374,N_2055,N_1829);
or U2375 (N_2375,N_1851,N_1978);
nor U2376 (N_2376,N_2170,N_2127);
and U2377 (N_2377,N_1946,N_1976);
and U2378 (N_2378,N_2088,N_1832);
or U2379 (N_2379,N_1994,N_2102);
nor U2380 (N_2380,N_1985,N_1983);
nor U2381 (N_2381,N_1877,N_1616);
nand U2382 (N_2382,N_1938,N_1864);
nand U2383 (N_2383,N_1945,N_1534);
and U2384 (N_2384,N_2143,N_1962);
nor U2385 (N_2385,N_1615,N_2191);
and U2386 (N_2386,N_1780,N_2247);
nand U2387 (N_2387,N_1973,N_1546);
and U2388 (N_2388,N_1922,N_1633);
nand U2389 (N_2389,N_1927,N_1710);
nor U2390 (N_2390,N_2105,N_2035);
nand U2391 (N_2391,N_1690,N_2027);
nor U2392 (N_2392,N_1732,N_1722);
nor U2393 (N_2393,N_2232,N_1853);
and U2394 (N_2394,N_1950,N_1809);
and U2395 (N_2395,N_1930,N_1640);
nor U2396 (N_2396,N_1770,N_1800);
nor U2397 (N_2397,N_2090,N_1782);
nand U2398 (N_2398,N_1730,N_1918);
nand U2399 (N_2399,N_2157,N_2217);
or U2400 (N_2400,N_2092,N_1573);
nand U2401 (N_2401,N_1794,N_1559);
nor U2402 (N_2402,N_1586,N_1972);
or U2403 (N_2403,N_1892,N_2172);
or U2404 (N_2404,N_1598,N_2005);
nand U2405 (N_2405,N_2118,N_2107);
and U2406 (N_2406,N_1997,N_1673);
nor U2407 (N_2407,N_1667,N_1542);
nor U2408 (N_2408,N_2040,N_1936);
and U2409 (N_2409,N_1992,N_1884);
nand U2410 (N_2410,N_1821,N_1639);
or U2411 (N_2411,N_1713,N_2059);
nand U2412 (N_2412,N_1828,N_1747);
nand U2413 (N_2413,N_1727,N_2095);
nor U2414 (N_2414,N_1544,N_1504);
and U2415 (N_2415,N_1530,N_1635);
nand U2416 (N_2416,N_2082,N_1689);
nand U2417 (N_2417,N_1629,N_2141);
nand U2418 (N_2418,N_1657,N_2072);
and U2419 (N_2419,N_1594,N_1755);
nor U2420 (N_2420,N_1601,N_2197);
nor U2421 (N_2421,N_2125,N_1763);
nand U2422 (N_2422,N_2126,N_1711);
and U2423 (N_2423,N_2243,N_1718);
or U2424 (N_2424,N_2079,N_1627);
or U2425 (N_2425,N_2056,N_1618);
nor U2426 (N_2426,N_2113,N_1729);
or U2427 (N_2427,N_2206,N_1630);
and U2428 (N_2428,N_1719,N_1822);
and U2429 (N_2429,N_2017,N_2015);
or U2430 (N_2430,N_2063,N_1964);
nor U2431 (N_2431,N_1582,N_1931);
nor U2432 (N_2432,N_2032,N_1656);
nand U2433 (N_2433,N_1647,N_2210);
nor U2434 (N_2434,N_2221,N_2067);
and U2435 (N_2435,N_2166,N_1599);
nand U2436 (N_2436,N_2046,N_1954);
nand U2437 (N_2437,N_1538,N_1777);
nor U2438 (N_2438,N_2031,N_2047);
nor U2439 (N_2439,N_1811,N_2028);
and U2440 (N_2440,N_1761,N_2117);
and U2441 (N_2441,N_1804,N_1675);
nand U2442 (N_2442,N_1815,N_1558);
nand U2443 (N_2443,N_2061,N_1704);
nor U2444 (N_2444,N_1979,N_1607);
nor U2445 (N_2445,N_2219,N_1696);
nor U2446 (N_2446,N_1933,N_1650);
and U2447 (N_2447,N_1734,N_2188);
and U2448 (N_2448,N_2034,N_2101);
or U2449 (N_2449,N_1810,N_1529);
nand U2450 (N_2450,N_2244,N_2176);
xor U2451 (N_2451,N_2119,N_1841);
or U2452 (N_2452,N_1970,N_1913);
or U2453 (N_2453,N_1880,N_1917);
and U2454 (N_2454,N_1798,N_1753);
or U2455 (N_2455,N_2163,N_2065);
nor U2456 (N_2456,N_1843,N_2081);
or U2457 (N_2457,N_2042,N_1561);
or U2458 (N_2458,N_2155,N_1890);
nor U2459 (N_2459,N_2077,N_2239);
or U2460 (N_2460,N_2033,N_2189);
xor U2461 (N_2461,N_2211,N_1914);
and U2462 (N_2462,N_1915,N_1870);
and U2463 (N_2463,N_1961,N_2076);
and U2464 (N_2464,N_2116,N_1847);
nor U2465 (N_2465,N_1515,N_2140);
and U2466 (N_2466,N_2123,N_2175);
and U2467 (N_2467,N_1539,N_1661);
or U2468 (N_2468,N_1805,N_1895);
or U2469 (N_2469,N_1891,N_1731);
nor U2470 (N_2470,N_2242,N_1874);
and U2471 (N_2471,N_1816,N_1860);
nor U2472 (N_2472,N_1700,N_1813);
nor U2473 (N_2473,N_1693,N_1614);
and U2474 (N_2474,N_1555,N_1833);
nor U2475 (N_2475,N_1665,N_1808);
and U2476 (N_2476,N_1757,N_2122);
nor U2477 (N_2477,N_1839,N_1511);
and U2478 (N_2478,N_2112,N_1745);
and U2479 (N_2479,N_1984,N_1621);
or U2480 (N_2480,N_1662,N_2237);
or U2481 (N_2481,N_1871,N_1846);
or U2482 (N_2482,N_1522,N_1898);
or U2483 (N_2483,N_2074,N_1521);
or U2484 (N_2484,N_1854,N_2241);
and U2485 (N_2485,N_1737,N_1622);
and U2486 (N_2486,N_1709,N_1610);
nor U2487 (N_2487,N_1684,N_2202);
nor U2488 (N_2488,N_1998,N_2132);
or U2489 (N_2489,N_2115,N_2054);
nand U2490 (N_2490,N_1654,N_2134);
nor U2491 (N_2491,N_2085,N_1641);
or U2492 (N_2492,N_2018,N_1624);
or U2493 (N_2493,N_2007,N_1959);
nand U2494 (N_2494,N_1743,N_1765);
nor U2495 (N_2495,N_2233,N_2216);
or U2496 (N_2496,N_1999,N_1778);
and U2497 (N_2497,N_1552,N_1912);
and U2498 (N_2498,N_1670,N_1550);
or U2499 (N_2499,N_2230,N_1678);
or U2500 (N_2500,N_1746,N_2213);
nor U2501 (N_2501,N_2236,N_2045);
and U2502 (N_2502,N_1502,N_1699);
and U2503 (N_2503,N_1904,N_2128);
and U2504 (N_2504,N_2144,N_1987);
or U2505 (N_2505,N_2190,N_1799);
or U2506 (N_2506,N_2075,N_1768);
or U2507 (N_2507,N_1916,N_2153);
and U2508 (N_2508,N_1835,N_1772);
nor U2509 (N_2509,N_1593,N_2013);
or U2510 (N_2510,N_1900,N_1888);
nand U2511 (N_2511,N_1720,N_1547);
nand U2512 (N_2512,N_1738,N_2130);
and U2513 (N_2513,N_2246,N_2106);
nand U2514 (N_2514,N_2220,N_2226);
nor U2515 (N_2515,N_1643,N_2010);
nand U2516 (N_2516,N_1535,N_1626);
nor U2517 (N_2517,N_1857,N_1974);
nor U2518 (N_2518,N_2168,N_1574);
nand U2519 (N_2519,N_1849,N_2071);
or U2520 (N_2520,N_1578,N_1868);
and U2521 (N_2521,N_1683,N_2185);
nand U2522 (N_2522,N_2078,N_1944);
nand U2523 (N_2523,N_1801,N_1563);
nand U2524 (N_2524,N_1569,N_1685);
or U2525 (N_2525,N_1596,N_2137);
or U2526 (N_2526,N_1564,N_1605);
or U2527 (N_2527,N_2228,N_2083);
nand U2528 (N_2528,N_1567,N_2161);
or U2529 (N_2529,N_1867,N_1652);
nand U2530 (N_2530,N_2198,N_1789);
or U2531 (N_2531,N_1896,N_1856);
or U2532 (N_2532,N_1911,N_1858);
nor U2533 (N_2533,N_1935,N_1638);
or U2534 (N_2534,N_1909,N_1551);
and U2535 (N_2535,N_2160,N_1669);
and U2536 (N_2536,N_2209,N_1842);
nand U2537 (N_2537,N_2053,N_2136);
nor U2538 (N_2538,N_1991,N_2066);
or U2539 (N_2539,N_2012,N_1990);
and U2540 (N_2540,N_1608,N_2184);
nor U2541 (N_2541,N_1876,N_2179);
xnor U2542 (N_2542,N_2050,N_1517);
and U2543 (N_2543,N_1659,N_1818);
nand U2544 (N_2544,N_2060,N_1824);
nor U2545 (N_2545,N_2205,N_1583);
nand U2546 (N_2546,N_2023,N_1592);
nor U2547 (N_2547,N_1982,N_1812);
and U2548 (N_2548,N_2174,N_1540);
nor U2549 (N_2549,N_1863,N_1902);
nand U2550 (N_2550,N_1966,N_2139);
or U2551 (N_2551,N_1943,N_2037);
or U2552 (N_2552,N_1663,N_1814);
or U2553 (N_2553,N_1631,N_2100);
nor U2554 (N_2554,N_2110,N_1906);
nand U2555 (N_2555,N_2173,N_1953);
nand U2556 (N_2556,N_1541,N_2156);
nor U2557 (N_2557,N_1686,N_1837);
nor U2558 (N_2558,N_2162,N_1721);
nor U2559 (N_2559,N_1702,N_1996);
nor U2560 (N_2560,N_1512,N_2043);
nand U2561 (N_2561,N_1878,N_1939);
nand U2562 (N_2562,N_1613,N_1957);
or U2563 (N_2563,N_2103,N_1588);
nor U2564 (N_2564,N_1764,N_1826);
or U2565 (N_2565,N_2229,N_2158);
nand U2566 (N_2566,N_1924,N_2138);
or U2567 (N_2567,N_1528,N_1967);
or U2568 (N_2568,N_1701,N_1723);
and U2569 (N_2569,N_1560,N_1579);
or U2570 (N_2570,N_2003,N_1862);
nor U2571 (N_2571,N_2094,N_1658);
nor U2572 (N_2572,N_1637,N_1844);
or U2573 (N_2573,N_2183,N_1572);
nand U2574 (N_2574,N_2070,N_2087);
nand U2575 (N_2575,N_1536,N_1672);
nand U2576 (N_2576,N_1776,N_1703);
and U2577 (N_2577,N_1792,N_2069);
nand U2578 (N_2578,N_1850,N_2041);
nand U2579 (N_2579,N_1750,N_2121);
and U2580 (N_2580,N_1692,N_2057);
and U2581 (N_2581,N_1698,N_1516);
or U2582 (N_2582,N_1510,N_1903);
nand U2583 (N_2583,N_1779,N_2104);
and U2584 (N_2584,N_1733,N_2049);
nor U2585 (N_2585,N_1553,N_1741);
and U2586 (N_2586,N_1664,N_2150);
nand U2587 (N_2587,N_1514,N_1714);
or U2588 (N_2588,N_1736,N_1531);
or U2589 (N_2589,N_1926,N_2006);
nor U2590 (N_2590,N_1742,N_2235);
or U2591 (N_2591,N_2152,N_1533);
nand U2592 (N_2592,N_1680,N_2238);
nor U2593 (N_2593,N_1602,N_1825);
and U2594 (N_2594,N_1784,N_2145);
and U2595 (N_2595,N_1648,N_1951);
nand U2596 (N_2596,N_1617,N_1893);
nor U2597 (N_2597,N_1655,N_2089);
nor U2598 (N_2598,N_2016,N_1695);
nand U2599 (N_2599,N_1752,N_2021);
and U2600 (N_2600,N_1875,N_2196);
or U2601 (N_2601,N_2019,N_1769);
or U2602 (N_2602,N_1980,N_2108);
nand U2603 (N_2603,N_1575,N_1785);
and U2604 (N_2604,N_2149,N_1653);
nor U2605 (N_2605,N_1948,N_2068);
or U2606 (N_2606,N_1671,N_1788);
nor U2607 (N_2607,N_1651,N_1759);
nand U2608 (N_2608,N_1793,N_2200);
nor U2609 (N_2609,N_1591,N_1694);
or U2610 (N_2610,N_1861,N_2201);
and U2611 (N_2611,N_1817,N_1803);
or U2612 (N_2612,N_2124,N_2009);
and U2613 (N_2613,N_2245,N_1744);
or U2614 (N_2614,N_1600,N_1905);
and U2615 (N_2615,N_2080,N_1956);
nand U2616 (N_2616,N_1925,N_2004);
and U2617 (N_2617,N_1688,N_2011);
or U2618 (N_2618,N_2025,N_1845);
or U2619 (N_2619,N_2146,N_1606);
or U2620 (N_2620,N_1819,N_1795);
nor U2621 (N_2621,N_2199,N_2052);
nor U2622 (N_2622,N_1932,N_1603);
nand U2623 (N_2623,N_2038,N_1724);
or U2624 (N_2624,N_1859,N_2097);
and U2625 (N_2625,N_1629,N_1870);
and U2626 (N_2626,N_2165,N_1842);
and U2627 (N_2627,N_2111,N_1676);
and U2628 (N_2628,N_1643,N_2158);
or U2629 (N_2629,N_1554,N_1991);
nand U2630 (N_2630,N_1707,N_2076);
nand U2631 (N_2631,N_1778,N_2005);
or U2632 (N_2632,N_2180,N_1591);
nor U2633 (N_2633,N_2121,N_1729);
and U2634 (N_2634,N_2124,N_1902);
and U2635 (N_2635,N_1965,N_1623);
or U2636 (N_2636,N_1580,N_1906);
or U2637 (N_2637,N_1615,N_1509);
and U2638 (N_2638,N_2178,N_1979);
or U2639 (N_2639,N_1721,N_1843);
or U2640 (N_2640,N_1993,N_2140);
and U2641 (N_2641,N_2005,N_1615);
and U2642 (N_2642,N_2069,N_1749);
nand U2643 (N_2643,N_1612,N_1871);
and U2644 (N_2644,N_1896,N_2020);
or U2645 (N_2645,N_2052,N_1554);
or U2646 (N_2646,N_1886,N_1953);
and U2647 (N_2647,N_2033,N_1753);
nor U2648 (N_2648,N_2142,N_1659);
nor U2649 (N_2649,N_1747,N_1995);
nor U2650 (N_2650,N_1691,N_1617);
nor U2651 (N_2651,N_1830,N_1659);
or U2652 (N_2652,N_1712,N_1503);
or U2653 (N_2653,N_2026,N_1571);
nor U2654 (N_2654,N_1530,N_1972);
and U2655 (N_2655,N_1709,N_1547);
or U2656 (N_2656,N_2128,N_1629);
and U2657 (N_2657,N_1764,N_1920);
or U2658 (N_2658,N_2133,N_2052);
and U2659 (N_2659,N_1531,N_1801);
or U2660 (N_2660,N_1845,N_1945);
nor U2661 (N_2661,N_1789,N_1768);
or U2662 (N_2662,N_1579,N_2041);
nor U2663 (N_2663,N_2013,N_2182);
or U2664 (N_2664,N_1724,N_1763);
or U2665 (N_2665,N_1704,N_1626);
nand U2666 (N_2666,N_1523,N_2038);
nor U2667 (N_2667,N_2218,N_2065);
nand U2668 (N_2668,N_1923,N_1893);
or U2669 (N_2669,N_1989,N_1927);
nor U2670 (N_2670,N_1562,N_1881);
and U2671 (N_2671,N_2173,N_1551);
or U2672 (N_2672,N_1730,N_1932);
or U2673 (N_2673,N_1939,N_1738);
and U2674 (N_2674,N_1504,N_1721);
nor U2675 (N_2675,N_2139,N_1616);
or U2676 (N_2676,N_1985,N_2018);
or U2677 (N_2677,N_1616,N_1684);
or U2678 (N_2678,N_1682,N_1673);
or U2679 (N_2679,N_1658,N_1615);
nor U2680 (N_2680,N_2210,N_2047);
or U2681 (N_2681,N_1508,N_1557);
or U2682 (N_2682,N_2098,N_1939);
and U2683 (N_2683,N_2117,N_1686);
nor U2684 (N_2684,N_1690,N_2047);
or U2685 (N_2685,N_2090,N_1867);
xor U2686 (N_2686,N_2194,N_1833);
or U2687 (N_2687,N_2031,N_1780);
or U2688 (N_2688,N_2212,N_2080);
and U2689 (N_2689,N_1751,N_1560);
nand U2690 (N_2690,N_1821,N_1543);
nand U2691 (N_2691,N_1905,N_1640);
or U2692 (N_2692,N_1807,N_2077);
and U2693 (N_2693,N_2018,N_1948);
nor U2694 (N_2694,N_2192,N_2111);
nand U2695 (N_2695,N_1801,N_1521);
nand U2696 (N_2696,N_1785,N_1768);
or U2697 (N_2697,N_2007,N_2116);
nor U2698 (N_2698,N_2130,N_2010);
nand U2699 (N_2699,N_1525,N_1545);
xnor U2700 (N_2700,N_2019,N_1845);
nor U2701 (N_2701,N_1549,N_1633);
nor U2702 (N_2702,N_1818,N_1762);
nand U2703 (N_2703,N_2228,N_1757);
xor U2704 (N_2704,N_2123,N_1942);
nand U2705 (N_2705,N_2241,N_2010);
or U2706 (N_2706,N_2233,N_2058);
nand U2707 (N_2707,N_1521,N_2240);
nor U2708 (N_2708,N_2073,N_2128);
and U2709 (N_2709,N_2139,N_2020);
nor U2710 (N_2710,N_1693,N_1889);
or U2711 (N_2711,N_2133,N_2163);
nor U2712 (N_2712,N_2121,N_1760);
nor U2713 (N_2713,N_1580,N_1829);
nor U2714 (N_2714,N_1543,N_1503);
nand U2715 (N_2715,N_1699,N_1592);
and U2716 (N_2716,N_2203,N_2160);
or U2717 (N_2717,N_1978,N_1942);
nor U2718 (N_2718,N_1832,N_2173);
or U2719 (N_2719,N_1780,N_1712);
and U2720 (N_2720,N_2076,N_1625);
nor U2721 (N_2721,N_2072,N_1812);
nor U2722 (N_2722,N_1865,N_2231);
and U2723 (N_2723,N_1794,N_1514);
nand U2724 (N_2724,N_1817,N_2173);
nand U2725 (N_2725,N_2154,N_1767);
nand U2726 (N_2726,N_1613,N_1652);
nand U2727 (N_2727,N_2177,N_2209);
nor U2728 (N_2728,N_1687,N_1840);
nor U2729 (N_2729,N_1979,N_2171);
nand U2730 (N_2730,N_2235,N_2024);
or U2731 (N_2731,N_1804,N_1566);
nor U2732 (N_2732,N_1681,N_2129);
and U2733 (N_2733,N_1652,N_2032);
and U2734 (N_2734,N_1736,N_1761);
nand U2735 (N_2735,N_1576,N_1896);
and U2736 (N_2736,N_1564,N_2163);
nand U2737 (N_2737,N_1793,N_1777);
and U2738 (N_2738,N_2011,N_1713);
or U2739 (N_2739,N_1908,N_1626);
and U2740 (N_2740,N_2105,N_1529);
nor U2741 (N_2741,N_1971,N_2033);
xor U2742 (N_2742,N_2201,N_2207);
and U2743 (N_2743,N_1660,N_2191);
or U2744 (N_2744,N_1551,N_1650);
nand U2745 (N_2745,N_1746,N_2013);
nor U2746 (N_2746,N_1828,N_2221);
nor U2747 (N_2747,N_1971,N_2157);
or U2748 (N_2748,N_2021,N_1694);
nor U2749 (N_2749,N_2088,N_2209);
and U2750 (N_2750,N_1778,N_1741);
nand U2751 (N_2751,N_1624,N_1894);
nor U2752 (N_2752,N_1699,N_2083);
and U2753 (N_2753,N_1836,N_1938);
nor U2754 (N_2754,N_1576,N_1531);
and U2755 (N_2755,N_2172,N_1577);
and U2756 (N_2756,N_2040,N_1998);
nand U2757 (N_2757,N_2235,N_1762);
and U2758 (N_2758,N_1689,N_1601);
nor U2759 (N_2759,N_2088,N_2138);
and U2760 (N_2760,N_1922,N_1848);
or U2761 (N_2761,N_2036,N_2221);
nand U2762 (N_2762,N_1860,N_1554);
nor U2763 (N_2763,N_1579,N_1837);
nor U2764 (N_2764,N_2050,N_2014);
and U2765 (N_2765,N_1532,N_2094);
nor U2766 (N_2766,N_2162,N_1528);
and U2767 (N_2767,N_1628,N_2059);
or U2768 (N_2768,N_1856,N_1701);
nor U2769 (N_2769,N_1622,N_2112);
or U2770 (N_2770,N_2019,N_1594);
nand U2771 (N_2771,N_1843,N_2020);
nor U2772 (N_2772,N_2180,N_2150);
nor U2773 (N_2773,N_1597,N_1658);
and U2774 (N_2774,N_1585,N_2229);
or U2775 (N_2775,N_1602,N_2120);
or U2776 (N_2776,N_2132,N_1897);
nor U2777 (N_2777,N_1632,N_2217);
and U2778 (N_2778,N_2185,N_1895);
nor U2779 (N_2779,N_2127,N_1999);
nand U2780 (N_2780,N_1833,N_1565);
and U2781 (N_2781,N_2012,N_2189);
or U2782 (N_2782,N_1693,N_1647);
nand U2783 (N_2783,N_1995,N_1841);
or U2784 (N_2784,N_1718,N_1812);
and U2785 (N_2785,N_1801,N_1667);
and U2786 (N_2786,N_1907,N_1711);
nand U2787 (N_2787,N_1702,N_2092);
nand U2788 (N_2788,N_2183,N_1586);
nand U2789 (N_2789,N_1779,N_1961);
nand U2790 (N_2790,N_1547,N_2138);
and U2791 (N_2791,N_1572,N_2086);
or U2792 (N_2792,N_2245,N_1506);
or U2793 (N_2793,N_1911,N_1984);
or U2794 (N_2794,N_2167,N_2170);
nand U2795 (N_2795,N_1682,N_2086);
or U2796 (N_2796,N_1643,N_1706);
nor U2797 (N_2797,N_1557,N_1761);
nand U2798 (N_2798,N_2216,N_1957);
nor U2799 (N_2799,N_1834,N_1614);
and U2800 (N_2800,N_2152,N_1768);
and U2801 (N_2801,N_2167,N_2161);
nor U2802 (N_2802,N_1970,N_1753);
or U2803 (N_2803,N_1609,N_1621);
nor U2804 (N_2804,N_1543,N_1957);
nor U2805 (N_2805,N_2053,N_1831);
nand U2806 (N_2806,N_1960,N_1851);
nor U2807 (N_2807,N_1763,N_1912);
or U2808 (N_2808,N_1977,N_2122);
nand U2809 (N_2809,N_1589,N_1967);
nand U2810 (N_2810,N_2041,N_2209);
and U2811 (N_2811,N_2142,N_1707);
nor U2812 (N_2812,N_1663,N_2187);
or U2813 (N_2813,N_1684,N_1958);
and U2814 (N_2814,N_1839,N_1665);
or U2815 (N_2815,N_1647,N_2074);
nand U2816 (N_2816,N_2147,N_1536);
and U2817 (N_2817,N_2188,N_1535);
nor U2818 (N_2818,N_1907,N_1928);
or U2819 (N_2819,N_2063,N_1853);
nand U2820 (N_2820,N_2130,N_1640);
nor U2821 (N_2821,N_1732,N_1761);
or U2822 (N_2822,N_2209,N_1669);
nor U2823 (N_2823,N_1889,N_1697);
nand U2824 (N_2824,N_2009,N_1532);
nand U2825 (N_2825,N_1995,N_1792);
and U2826 (N_2826,N_1894,N_1749);
and U2827 (N_2827,N_1686,N_2235);
nor U2828 (N_2828,N_1748,N_1973);
and U2829 (N_2829,N_1559,N_1567);
and U2830 (N_2830,N_1576,N_1524);
nor U2831 (N_2831,N_1991,N_1644);
nand U2832 (N_2832,N_1999,N_1532);
nor U2833 (N_2833,N_2103,N_2207);
nand U2834 (N_2834,N_1736,N_1694);
and U2835 (N_2835,N_1597,N_1840);
nand U2836 (N_2836,N_2053,N_2245);
and U2837 (N_2837,N_2043,N_2185);
and U2838 (N_2838,N_2213,N_2080);
or U2839 (N_2839,N_1808,N_1857);
nor U2840 (N_2840,N_1957,N_1905);
nor U2841 (N_2841,N_1919,N_1680);
nand U2842 (N_2842,N_2057,N_2152);
nor U2843 (N_2843,N_1945,N_1915);
or U2844 (N_2844,N_1760,N_1755);
or U2845 (N_2845,N_1595,N_2210);
nand U2846 (N_2846,N_1962,N_2006);
xnor U2847 (N_2847,N_2131,N_2245);
nor U2848 (N_2848,N_1806,N_1587);
or U2849 (N_2849,N_1736,N_2176);
nand U2850 (N_2850,N_1830,N_1946);
and U2851 (N_2851,N_2032,N_1594);
or U2852 (N_2852,N_1792,N_1895);
or U2853 (N_2853,N_1886,N_1866);
or U2854 (N_2854,N_1765,N_2141);
nor U2855 (N_2855,N_1841,N_1989);
nor U2856 (N_2856,N_2154,N_1531);
nand U2857 (N_2857,N_2091,N_1880);
nor U2858 (N_2858,N_1845,N_1625);
and U2859 (N_2859,N_1552,N_1999);
nor U2860 (N_2860,N_2097,N_2169);
and U2861 (N_2861,N_1928,N_1697);
nor U2862 (N_2862,N_2170,N_1587);
and U2863 (N_2863,N_1596,N_1992);
and U2864 (N_2864,N_1910,N_2121);
nor U2865 (N_2865,N_1536,N_1862);
and U2866 (N_2866,N_1704,N_2036);
or U2867 (N_2867,N_2248,N_2189);
nor U2868 (N_2868,N_2108,N_1958);
nand U2869 (N_2869,N_2159,N_1647);
nor U2870 (N_2870,N_2059,N_2094);
nor U2871 (N_2871,N_2199,N_1539);
or U2872 (N_2872,N_1905,N_1507);
nor U2873 (N_2873,N_1863,N_2126);
nand U2874 (N_2874,N_1829,N_1947);
and U2875 (N_2875,N_1529,N_1738);
nor U2876 (N_2876,N_1536,N_1979);
or U2877 (N_2877,N_2243,N_2088);
nor U2878 (N_2878,N_1511,N_2002);
and U2879 (N_2879,N_2115,N_2107);
and U2880 (N_2880,N_1616,N_2045);
or U2881 (N_2881,N_1633,N_1797);
or U2882 (N_2882,N_1699,N_1973);
and U2883 (N_2883,N_1771,N_2231);
and U2884 (N_2884,N_1859,N_2231);
and U2885 (N_2885,N_1970,N_1982);
or U2886 (N_2886,N_2206,N_1760);
nand U2887 (N_2887,N_1803,N_1539);
nand U2888 (N_2888,N_1839,N_1588);
and U2889 (N_2889,N_1884,N_1598);
and U2890 (N_2890,N_1775,N_2006);
or U2891 (N_2891,N_1706,N_2247);
and U2892 (N_2892,N_2142,N_1784);
nand U2893 (N_2893,N_2037,N_1870);
nand U2894 (N_2894,N_1988,N_1829);
xor U2895 (N_2895,N_1940,N_1758);
or U2896 (N_2896,N_1816,N_2099);
nor U2897 (N_2897,N_1885,N_1747);
and U2898 (N_2898,N_1670,N_1950);
nor U2899 (N_2899,N_2040,N_1823);
and U2900 (N_2900,N_2232,N_1525);
and U2901 (N_2901,N_1971,N_1715);
nand U2902 (N_2902,N_2130,N_1773);
nor U2903 (N_2903,N_1894,N_1632);
xnor U2904 (N_2904,N_2202,N_1796);
nor U2905 (N_2905,N_1541,N_2005);
nand U2906 (N_2906,N_2052,N_2248);
or U2907 (N_2907,N_1540,N_1649);
and U2908 (N_2908,N_1672,N_1847);
nand U2909 (N_2909,N_1591,N_1660);
nand U2910 (N_2910,N_2218,N_2034);
and U2911 (N_2911,N_2069,N_2174);
and U2912 (N_2912,N_1927,N_1544);
nor U2913 (N_2913,N_2018,N_1958);
or U2914 (N_2914,N_2206,N_1593);
nor U2915 (N_2915,N_1890,N_1501);
or U2916 (N_2916,N_1807,N_1513);
or U2917 (N_2917,N_2025,N_1866);
nand U2918 (N_2918,N_2053,N_2174);
and U2919 (N_2919,N_1605,N_1604);
nand U2920 (N_2920,N_1918,N_2122);
nand U2921 (N_2921,N_1983,N_1745);
nor U2922 (N_2922,N_1930,N_1959);
or U2923 (N_2923,N_1689,N_2036);
xnor U2924 (N_2924,N_1929,N_2225);
and U2925 (N_2925,N_1975,N_1810);
nand U2926 (N_2926,N_2039,N_2070);
or U2927 (N_2927,N_1889,N_1909);
nand U2928 (N_2928,N_2019,N_1740);
or U2929 (N_2929,N_2140,N_2198);
nand U2930 (N_2930,N_2179,N_1542);
and U2931 (N_2931,N_1831,N_2176);
nor U2932 (N_2932,N_1984,N_1922);
nor U2933 (N_2933,N_1987,N_1620);
nand U2934 (N_2934,N_2238,N_1876);
nor U2935 (N_2935,N_1887,N_1872);
nand U2936 (N_2936,N_2019,N_1833);
nor U2937 (N_2937,N_1842,N_1680);
or U2938 (N_2938,N_1695,N_1638);
nor U2939 (N_2939,N_1975,N_1788);
nand U2940 (N_2940,N_1593,N_1543);
and U2941 (N_2941,N_2181,N_1504);
nand U2942 (N_2942,N_2064,N_1983);
or U2943 (N_2943,N_1951,N_2017);
nor U2944 (N_2944,N_1992,N_1974);
nand U2945 (N_2945,N_2119,N_2240);
or U2946 (N_2946,N_1969,N_2216);
nor U2947 (N_2947,N_2144,N_1513);
nor U2948 (N_2948,N_2041,N_2110);
nor U2949 (N_2949,N_2091,N_1760);
or U2950 (N_2950,N_1646,N_1545);
or U2951 (N_2951,N_1750,N_1754);
or U2952 (N_2952,N_2172,N_1697);
and U2953 (N_2953,N_2018,N_1810);
or U2954 (N_2954,N_2033,N_1647);
and U2955 (N_2955,N_1563,N_1781);
or U2956 (N_2956,N_1930,N_2147);
or U2957 (N_2957,N_1615,N_2041);
nor U2958 (N_2958,N_2190,N_1762);
nor U2959 (N_2959,N_1784,N_1798);
nor U2960 (N_2960,N_1845,N_2047);
or U2961 (N_2961,N_2175,N_2075);
nand U2962 (N_2962,N_2138,N_2064);
and U2963 (N_2963,N_2046,N_1950);
and U2964 (N_2964,N_1832,N_1584);
and U2965 (N_2965,N_1870,N_1582);
nor U2966 (N_2966,N_1676,N_2198);
nand U2967 (N_2967,N_1891,N_1958);
nand U2968 (N_2968,N_1970,N_1911);
and U2969 (N_2969,N_1849,N_1966);
and U2970 (N_2970,N_1928,N_2202);
nor U2971 (N_2971,N_2192,N_2166);
or U2972 (N_2972,N_1864,N_1561);
and U2973 (N_2973,N_1959,N_2186);
and U2974 (N_2974,N_1527,N_1586);
and U2975 (N_2975,N_1846,N_1522);
or U2976 (N_2976,N_1609,N_1983);
and U2977 (N_2977,N_1871,N_1827);
or U2978 (N_2978,N_1691,N_2130);
and U2979 (N_2979,N_1627,N_2147);
nand U2980 (N_2980,N_1510,N_1809);
nand U2981 (N_2981,N_1560,N_1964);
and U2982 (N_2982,N_1552,N_1691);
or U2983 (N_2983,N_1968,N_1950);
and U2984 (N_2984,N_1874,N_2228);
nand U2985 (N_2985,N_1907,N_1849);
nand U2986 (N_2986,N_2132,N_1857);
nand U2987 (N_2987,N_1978,N_1887);
or U2988 (N_2988,N_1595,N_2162);
nand U2989 (N_2989,N_1948,N_1734);
or U2990 (N_2990,N_1518,N_1660);
nand U2991 (N_2991,N_1625,N_2014);
nor U2992 (N_2992,N_2149,N_1777);
or U2993 (N_2993,N_1670,N_1633);
nor U2994 (N_2994,N_1947,N_2056);
nor U2995 (N_2995,N_1773,N_2055);
and U2996 (N_2996,N_2001,N_2208);
or U2997 (N_2997,N_1748,N_1521);
nor U2998 (N_2998,N_2046,N_1674);
and U2999 (N_2999,N_2063,N_1785);
nand UO_0 (O_0,N_2346,N_2799);
nor UO_1 (O_1,N_2617,N_2338);
nor UO_2 (O_2,N_2357,N_2405);
nor UO_3 (O_3,N_2531,N_2560);
nand UO_4 (O_4,N_2948,N_2507);
and UO_5 (O_5,N_2317,N_2668);
nor UO_6 (O_6,N_2651,N_2425);
xor UO_7 (O_7,N_2774,N_2902);
or UO_8 (O_8,N_2616,N_2546);
nor UO_9 (O_9,N_2390,N_2622);
or UO_10 (O_10,N_2536,N_2772);
and UO_11 (O_11,N_2904,N_2387);
or UO_12 (O_12,N_2587,N_2377);
nor UO_13 (O_13,N_2938,N_2918);
nand UO_14 (O_14,N_2978,N_2694);
or UO_15 (O_15,N_2707,N_2399);
or UO_16 (O_16,N_2781,N_2964);
nand UO_17 (O_17,N_2987,N_2514);
nor UO_18 (O_18,N_2613,N_2788);
nor UO_19 (O_19,N_2813,N_2720);
and UO_20 (O_20,N_2309,N_2701);
or UO_21 (O_21,N_2812,N_2595);
nand UO_22 (O_22,N_2322,N_2517);
nand UO_23 (O_23,N_2401,N_2796);
and UO_24 (O_24,N_2581,N_2940);
or UO_25 (O_25,N_2681,N_2873);
nand UO_26 (O_26,N_2300,N_2751);
nand UO_27 (O_27,N_2963,N_2807);
xnor UO_28 (O_28,N_2974,N_2254);
or UO_29 (O_29,N_2883,N_2474);
or UO_30 (O_30,N_2965,N_2336);
or UO_31 (O_31,N_2422,N_2716);
and UO_32 (O_32,N_2747,N_2782);
and UO_33 (O_33,N_2342,N_2618);
nor UO_34 (O_34,N_2693,N_2915);
nand UO_35 (O_35,N_2828,N_2705);
and UO_36 (O_36,N_2732,N_2424);
nand UO_37 (O_37,N_2733,N_2495);
nor UO_38 (O_38,N_2354,N_2385);
and UO_39 (O_39,N_2262,N_2848);
nand UO_40 (O_40,N_2988,N_2870);
nor UO_41 (O_41,N_2440,N_2593);
and UO_42 (O_42,N_2416,N_2480);
and UO_43 (O_43,N_2676,N_2910);
nor UO_44 (O_44,N_2833,N_2543);
nor UO_45 (O_45,N_2599,N_2626);
and UO_46 (O_46,N_2684,N_2430);
nand UO_47 (O_47,N_2816,N_2648);
nand UO_48 (O_48,N_2961,N_2370);
nor UO_49 (O_49,N_2559,N_2468);
and UO_50 (O_50,N_2927,N_2291);
nor UO_51 (O_51,N_2650,N_2327);
and UO_52 (O_52,N_2276,N_2880);
nor UO_53 (O_53,N_2275,N_2995);
nand UO_54 (O_54,N_2689,N_2408);
nor UO_55 (O_55,N_2836,N_2766);
or UO_56 (O_56,N_2257,N_2742);
and UO_57 (O_57,N_2889,N_2516);
nor UO_58 (O_58,N_2971,N_2597);
or UO_59 (O_59,N_2420,N_2548);
nor UO_60 (O_60,N_2897,N_2578);
nor UO_61 (O_61,N_2312,N_2955);
nand UO_62 (O_62,N_2643,N_2875);
nor UO_63 (O_63,N_2361,N_2515);
and UO_64 (O_64,N_2922,N_2809);
nand UO_65 (O_65,N_2538,N_2951);
and UO_66 (O_66,N_2724,N_2776);
nand UO_67 (O_67,N_2339,N_2662);
or UO_68 (O_68,N_2803,N_2784);
nor UO_69 (O_69,N_2590,N_2690);
or UO_70 (O_70,N_2646,N_2448);
or UO_71 (O_71,N_2944,N_2350);
or UO_72 (O_72,N_2632,N_2274);
nor UO_73 (O_73,N_2804,N_2786);
and UO_74 (O_74,N_2400,N_2564);
and UO_75 (O_75,N_2638,N_2523);
and UO_76 (O_76,N_2872,N_2509);
nor UO_77 (O_77,N_2310,N_2612);
and UO_78 (O_78,N_2982,N_2697);
nand UO_79 (O_79,N_2834,N_2759);
nor UO_80 (O_80,N_2882,N_2688);
and UO_81 (O_81,N_2271,N_2823);
or UO_82 (O_82,N_2905,N_2476);
or UO_83 (O_83,N_2925,N_2885);
or UO_84 (O_84,N_2343,N_2952);
nand UO_85 (O_85,N_2455,N_2976);
nor UO_86 (O_86,N_2734,N_2421);
and UO_87 (O_87,N_2829,N_2996);
or UO_88 (O_88,N_2403,N_2798);
nand UO_89 (O_89,N_2534,N_2535);
and UO_90 (O_90,N_2969,N_2550);
or UO_91 (O_91,N_2447,N_2749);
or UO_92 (O_92,N_2364,N_2903);
and UO_93 (O_93,N_2777,N_2606);
nor UO_94 (O_94,N_2737,N_2344);
nor UO_95 (O_95,N_2436,N_2609);
nor UO_96 (O_96,N_2859,N_2417);
nand UO_97 (O_97,N_2864,N_2544);
or UO_98 (O_98,N_2847,N_2877);
nand UO_99 (O_99,N_2814,N_2503);
nand UO_100 (O_100,N_2946,N_2849);
and UO_101 (O_101,N_2950,N_2696);
nand UO_102 (O_102,N_2414,N_2497);
nand UO_103 (O_103,N_2710,N_2579);
or UO_104 (O_104,N_2673,N_2529);
and UO_105 (O_105,N_2522,N_2375);
nand UO_106 (O_106,N_2450,N_2429);
or UO_107 (O_107,N_2585,N_2819);
and UO_108 (O_108,N_2933,N_2661);
or UO_109 (O_109,N_2332,N_2261);
nor UO_110 (O_110,N_2469,N_2947);
and UO_111 (O_111,N_2610,N_2325);
nand UO_112 (O_112,N_2319,N_2934);
and UO_113 (O_113,N_2901,N_2504);
or UO_114 (O_114,N_2380,N_2820);
nand UO_115 (O_115,N_2753,N_2482);
nor UO_116 (O_116,N_2827,N_2392);
nand UO_117 (O_117,N_2574,N_2633);
and UO_118 (O_118,N_2491,N_2333);
or UO_119 (O_119,N_2962,N_2444);
and UO_120 (O_120,N_2348,N_2349);
nor UO_121 (O_121,N_2323,N_2306);
nor UO_122 (O_122,N_2499,N_2711);
nor UO_123 (O_123,N_2506,N_2647);
nor UO_124 (O_124,N_2808,N_2556);
nand UO_125 (O_125,N_2605,N_2252);
and UO_126 (O_126,N_2384,N_2973);
or UO_127 (O_127,N_2869,N_2473);
nand UO_128 (O_128,N_2727,N_2362);
or UO_129 (O_129,N_2841,N_2663);
and UO_130 (O_130,N_2551,N_2467);
nand UO_131 (O_131,N_2260,N_2966);
or UO_132 (O_132,N_2360,N_2998);
nor UO_133 (O_133,N_2908,N_2914);
and UO_134 (O_134,N_2815,N_2671);
nor UO_135 (O_135,N_2975,N_2328);
nand UO_136 (O_136,N_2537,N_2715);
nor UO_137 (O_137,N_2459,N_2582);
and UO_138 (O_138,N_2958,N_2856);
or UO_139 (O_139,N_2764,N_2866);
and UO_140 (O_140,N_2717,N_2899);
nand UO_141 (O_141,N_2657,N_2780);
nor UO_142 (O_142,N_2685,N_2383);
and UO_143 (O_143,N_2294,N_2972);
and UO_144 (O_144,N_2528,N_2394);
nand UO_145 (O_145,N_2907,N_2505);
xnor UO_146 (O_146,N_2852,N_2817);
or UO_147 (O_147,N_2960,N_2708);
nor UO_148 (O_148,N_2992,N_2270);
nand UO_149 (O_149,N_2356,N_2431);
and UO_150 (O_150,N_2921,N_2519);
nand UO_151 (O_151,N_2674,N_2494);
nand UO_152 (O_152,N_2340,N_2412);
nor UO_153 (O_153,N_2686,N_2532);
and UO_154 (O_154,N_2396,N_2754);
nand UO_155 (O_155,N_2454,N_2884);
and UO_156 (O_156,N_2266,N_2586);
or UO_157 (O_157,N_2267,N_2959);
nand UO_158 (O_158,N_2572,N_2418);
nand UO_159 (O_159,N_2939,N_2824);
or UO_160 (O_160,N_2743,N_2863);
nor UO_161 (O_161,N_2488,N_2943);
and UO_162 (O_162,N_2700,N_2839);
nor UO_163 (O_163,N_2890,N_2789);
and UO_164 (O_164,N_2862,N_2576);
xor UO_165 (O_165,N_2453,N_2462);
or UO_166 (O_166,N_2712,N_2288);
and UO_167 (O_167,N_2264,N_2457);
or UO_168 (O_168,N_2845,N_2787);
and UO_169 (O_169,N_2888,N_2744);
and UO_170 (O_170,N_2296,N_2466);
or UO_171 (O_171,N_2680,N_2692);
nor UO_172 (O_172,N_2793,N_2860);
or UO_173 (O_173,N_2896,N_2575);
nor UO_174 (O_174,N_2320,N_2871);
nand UO_175 (O_175,N_2278,N_2561);
nand UO_176 (O_176,N_2463,N_2533);
nand UO_177 (O_177,N_2985,N_2893);
nor UO_178 (O_178,N_2381,N_2659);
nor UO_179 (O_179,N_2917,N_2378);
and UO_180 (O_180,N_2486,N_2409);
and UO_181 (O_181,N_2299,N_2580);
or UO_182 (O_182,N_2750,N_2555);
nand UO_183 (O_183,N_2351,N_2855);
and UO_184 (O_184,N_2930,N_2801);
and UO_185 (O_185,N_2876,N_2878);
and UO_186 (O_186,N_2990,N_2567);
xor UO_187 (O_187,N_2513,N_2314);
nor UO_188 (O_188,N_2916,N_2675);
nand UO_189 (O_189,N_2695,N_2725);
nand UO_190 (O_190,N_2308,N_2968);
nor UO_191 (O_191,N_2746,N_2602);
or UO_192 (O_192,N_2691,N_2280);
or UO_193 (O_193,N_2376,N_2379);
or UO_194 (O_194,N_2667,N_2924);
or UO_195 (O_195,N_2830,N_2584);
nand UO_196 (O_196,N_2837,N_2923);
nor UO_197 (O_197,N_2778,N_2398);
nor UO_198 (O_198,N_2557,N_2986);
or UO_199 (O_199,N_2524,N_2954);
and UO_200 (O_200,N_2769,N_2989);
or UO_201 (O_201,N_2500,N_2838);
and UO_202 (O_202,N_2891,N_2620);
and UO_203 (O_203,N_2723,N_2573);
nand UO_204 (O_204,N_2371,N_2931);
nand UO_205 (O_205,N_2832,N_2779);
nor UO_206 (O_206,N_2419,N_2461);
and UO_207 (O_207,N_2645,N_2679);
nand UO_208 (O_208,N_2324,N_2406);
nor UO_209 (O_209,N_2337,N_2740);
nor UO_210 (O_210,N_2552,N_2826);
nand UO_211 (O_211,N_2365,N_2977);
xor UO_212 (O_212,N_2775,N_2570);
nor UO_213 (O_213,N_2683,N_2490);
nor UO_214 (O_214,N_2911,N_2670);
or UO_215 (O_215,N_2635,N_2352);
nand UO_216 (O_216,N_2472,N_2452);
and UO_217 (O_217,N_2372,N_2304);
and UO_218 (O_218,N_2331,N_2456);
nor UO_219 (O_219,N_2255,N_2843);
nor UO_220 (O_220,N_2525,N_2434);
nor UO_221 (O_221,N_2539,N_2442);
nand UO_222 (O_222,N_2677,N_2449);
and UO_223 (O_223,N_2251,N_2664);
or UO_224 (O_224,N_2660,N_2687);
nand UO_225 (O_225,N_2854,N_2588);
nor UO_226 (O_226,N_2404,N_2485);
or UO_227 (O_227,N_2993,N_2920);
nor UO_228 (O_228,N_2757,N_2991);
nand UO_229 (O_229,N_2393,N_2512);
or UO_230 (O_230,N_2805,N_2566);
or UO_231 (O_231,N_2530,N_2835);
nor UO_232 (O_232,N_2526,N_2496);
or UO_233 (O_233,N_2821,N_2407);
nand UO_234 (O_234,N_2840,N_2790);
nand UO_235 (O_235,N_2831,N_2460);
nand UO_236 (O_236,N_2865,N_2928);
nor UO_237 (O_237,N_2281,N_2699);
or UO_238 (O_238,N_2297,N_2912);
and UO_239 (O_239,N_2983,N_2762);
nor UO_240 (O_240,N_2756,N_2967);
and UO_241 (O_241,N_2373,N_2748);
or UO_242 (O_242,N_2458,N_2721);
nor UO_243 (O_243,N_2432,N_2761);
nor UO_244 (O_244,N_2621,N_2795);
nand UO_245 (O_245,N_2604,N_2636);
nor UO_246 (O_246,N_2624,N_2886);
nor UO_247 (O_247,N_2678,N_2438);
and UO_248 (O_248,N_2942,N_2366);
or UO_249 (O_249,N_2510,N_2501);
or UO_250 (O_250,N_2284,N_2825);
and UO_251 (O_251,N_2311,N_2481);
and UO_252 (O_252,N_2984,N_2415);
or UO_253 (O_253,N_2895,N_2722);
or UO_254 (O_254,N_2511,N_2554);
nor UO_255 (O_255,N_2439,N_2359);
and UO_256 (O_256,N_2818,N_2521);
or UO_257 (O_257,N_2731,N_2303);
nand UO_258 (O_258,N_2881,N_2253);
or UO_259 (O_259,N_2850,N_2773);
nor UO_260 (O_260,N_2611,N_2286);
and UO_261 (O_261,N_2771,N_2316);
nand UO_262 (O_262,N_2464,N_2487);
nor UO_263 (O_263,N_2791,N_2806);
nand UO_264 (O_264,N_2713,N_2427);
or UO_265 (O_265,N_2479,N_2601);
nor UO_266 (O_266,N_2335,N_2637);
and UO_267 (O_267,N_2298,N_2752);
nand UO_268 (O_268,N_2250,N_2282);
nor UO_269 (O_269,N_2493,N_2368);
nor UO_270 (O_270,N_2642,N_2802);
or UO_271 (O_271,N_2549,N_2568);
or UO_272 (O_272,N_2811,N_2330);
and UO_273 (O_273,N_2656,N_2935);
nand UO_274 (O_274,N_2545,N_2639);
nand UO_275 (O_275,N_2341,N_2956);
nor UO_276 (O_276,N_2857,N_2861);
nand UO_277 (O_277,N_2402,N_2269);
nand UO_278 (O_278,N_2290,N_2594);
and UO_279 (O_279,N_2589,N_2413);
nand UO_280 (O_280,N_2329,N_2600);
nand UO_281 (O_281,N_2313,N_2718);
nor UO_282 (O_282,N_2738,N_2706);
and UO_283 (O_283,N_2489,N_2936);
and UO_284 (O_284,N_2614,N_2669);
nor UO_285 (O_285,N_2492,N_2653);
or UO_286 (O_286,N_2665,N_2388);
nor UO_287 (O_287,N_2446,N_2293);
or UO_288 (O_288,N_2334,N_2318);
nor UO_289 (O_289,N_2547,N_2358);
and UO_290 (O_290,N_2906,N_2728);
and UO_291 (O_291,N_2726,N_2760);
nand UO_292 (O_292,N_2471,N_2979);
and UO_293 (O_293,N_2397,N_2592);
or UO_294 (O_294,N_2265,N_2997);
or UO_295 (O_295,N_2879,N_2435);
and UO_296 (O_296,N_2672,N_2714);
nor UO_297 (O_297,N_2465,N_2623);
or UO_298 (O_298,N_2758,N_2355);
or UO_299 (O_299,N_2596,N_2391);
nand UO_300 (O_300,N_2794,N_2563);
nand UO_301 (O_301,N_2478,N_2287);
or UO_302 (O_302,N_2520,N_2553);
or UO_303 (O_303,N_2631,N_2347);
or UO_304 (O_304,N_2851,N_2326);
nor UO_305 (O_305,N_2792,N_2315);
nand UO_306 (O_306,N_2562,N_2268);
nand UO_307 (O_307,N_2702,N_2698);
nand UO_308 (O_308,N_2628,N_2745);
nor UO_309 (O_309,N_2445,N_2625);
nand UO_310 (O_310,N_2981,N_2258);
nand UO_311 (O_311,N_2542,N_2949);
or UO_312 (O_312,N_2797,N_2929);
or UO_313 (O_313,N_2867,N_2844);
and UO_314 (O_314,N_2598,N_2709);
nand UO_315 (O_315,N_2898,N_2703);
or UO_316 (O_316,N_2367,N_2767);
nand UO_317 (O_317,N_2498,N_2874);
and UO_318 (O_318,N_2649,N_2259);
nor UO_319 (O_319,N_2437,N_2846);
and UO_320 (O_320,N_2634,N_2704);
nand UO_321 (O_321,N_2518,N_2423);
or UO_322 (O_322,N_2540,N_2272);
nor UO_323 (O_323,N_2443,N_2256);
or UO_324 (O_324,N_2302,N_2652);
or UO_325 (O_325,N_2741,N_2800);
or UO_326 (O_326,N_2654,N_2369);
or UO_327 (O_327,N_2426,N_2382);
nor UO_328 (O_328,N_2591,N_2629);
and UO_329 (O_329,N_2627,N_2603);
nor UO_330 (O_330,N_2953,N_2353);
or UO_331 (O_331,N_2433,N_2345);
nor UO_332 (O_332,N_2301,N_2941);
or UO_333 (O_333,N_2842,N_2451);
nand UO_334 (O_334,N_2900,N_2735);
nand UO_335 (O_335,N_2729,N_2441);
and UO_336 (O_336,N_2909,N_2508);
nand UO_337 (O_337,N_2785,N_2892);
nor UO_338 (O_338,N_2428,N_2926);
nor UO_339 (O_339,N_2768,N_2571);
nand UO_340 (O_340,N_2307,N_2755);
and UO_341 (O_341,N_2957,N_2763);
or UO_342 (O_342,N_2887,N_2527);
nand UO_343 (O_343,N_2395,N_2810);
nor UO_344 (O_344,N_2363,N_2736);
or UO_345 (O_345,N_2640,N_2644);
and UO_346 (O_346,N_2283,N_2894);
and UO_347 (O_347,N_2630,N_2483);
and UO_348 (O_348,N_2484,N_2583);
or UO_349 (O_349,N_2608,N_2932);
nand UO_350 (O_350,N_2658,N_2666);
nand UO_351 (O_351,N_2765,N_2945);
and UO_352 (O_352,N_2937,N_2739);
nor UO_353 (O_353,N_2619,N_2277);
nand UO_354 (O_354,N_2292,N_2682);
or UO_355 (O_355,N_2999,N_2411);
and UO_356 (O_356,N_2565,N_2321);
and UO_357 (O_357,N_2783,N_2477);
nand UO_358 (O_358,N_2305,N_2719);
and UO_359 (O_359,N_2822,N_2263);
and UO_360 (O_360,N_2386,N_2913);
nor UO_361 (O_361,N_2569,N_2374);
nor UO_362 (O_362,N_2858,N_2994);
nor UO_363 (O_363,N_2853,N_2615);
nor UO_364 (O_364,N_2502,N_2980);
or UO_365 (O_365,N_2577,N_2770);
nor UO_366 (O_366,N_2475,N_2289);
nor UO_367 (O_367,N_2607,N_2970);
or UO_368 (O_368,N_2279,N_2541);
or UO_369 (O_369,N_2919,N_2641);
or UO_370 (O_370,N_2730,N_2410);
and UO_371 (O_371,N_2273,N_2389);
and UO_372 (O_372,N_2655,N_2295);
nand UO_373 (O_373,N_2868,N_2558);
nor UO_374 (O_374,N_2470,N_2285);
nor UO_375 (O_375,N_2810,N_2818);
nor UO_376 (O_376,N_2662,N_2530);
and UO_377 (O_377,N_2538,N_2624);
nand UO_378 (O_378,N_2924,N_2901);
nor UO_379 (O_379,N_2712,N_2811);
nor UO_380 (O_380,N_2658,N_2582);
nand UO_381 (O_381,N_2523,N_2819);
nor UO_382 (O_382,N_2437,N_2418);
and UO_383 (O_383,N_2329,N_2523);
nand UO_384 (O_384,N_2612,N_2916);
and UO_385 (O_385,N_2986,N_2787);
and UO_386 (O_386,N_2888,N_2515);
or UO_387 (O_387,N_2997,N_2922);
nor UO_388 (O_388,N_2869,N_2484);
nand UO_389 (O_389,N_2497,N_2280);
nor UO_390 (O_390,N_2631,N_2653);
and UO_391 (O_391,N_2905,N_2856);
or UO_392 (O_392,N_2652,N_2583);
and UO_393 (O_393,N_2331,N_2390);
nor UO_394 (O_394,N_2989,N_2679);
nor UO_395 (O_395,N_2963,N_2965);
or UO_396 (O_396,N_2654,N_2674);
nor UO_397 (O_397,N_2946,N_2255);
and UO_398 (O_398,N_2971,N_2487);
nor UO_399 (O_399,N_2674,N_2263);
or UO_400 (O_400,N_2500,N_2495);
nand UO_401 (O_401,N_2771,N_2708);
and UO_402 (O_402,N_2788,N_2989);
nor UO_403 (O_403,N_2925,N_2549);
or UO_404 (O_404,N_2825,N_2321);
nor UO_405 (O_405,N_2358,N_2418);
nor UO_406 (O_406,N_2493,N_2264);
nor UO_407 (O_407,N_2748,N_2943);
or UO_408 (O_408,N_2803,N_2276);
nand UO_409 (O_409,N_2552,N_2671);
nand UO_410 (O_410,N_2456,N_2387);
or UO_411 (O_411,N_2388,N_2692);
and UO_412 (O_412,N_2392,N_2779);
nor UO_413 (O_413,N_2589,N_2786);
or UO_414 (O_414,N_2797,N_2681);
nor UO_415 (O_415,N_2416,N_2719);
and UO_416 (O_416,N_2826,N_2577);
or UO_417 (O_417,N_2565,N_2474);
nor UO_418 (O_418,N_2404,N_2601);
and UO_419 (O_419,N_2316,N_2556);
nand UO_420 (O_420,N_2336,N_2691);
and UO_421 (O_421,N_2373,N_2825);
nand UO_422 (O_422,N_2918,N_2255);
and UO_423 (O_423,N_2867,N_2550);
nand UO_424 (O_424,N_2853,N_2465);
and UO_425 (O_425,N_2441,N_2623);
nor UO_426 (O_426,N_2377,N_2290);
nand UO_427 (O_427,N_2808,N_2291);
nand UO_428 (O_428,N_2437,N_2736);
and UO_429 (O_429,N_2401,N_2886);
or UO_430 (O_430,N_2718,N_2891);
xnor UO_431 (O_431,N_2789,N_2363);
nor UO_432 (O_432,N_2444,N_2317);
nand UO_433 (O_433,N_2732,N_2688);
nand UO_434 (O_434,N_2913,N_2308);
nand UO_435 (O_435,N_2524,N_2904);
and UO_436 (O_436,N_2734,N_2896);
and UO_437 (O_437,N_2885,N_2321);
nand UO_438 (O_438,N_2884,N_2807);
or UO_439 (O_439,N_2754,N_2486);
nand UO_440 (O_440,N_2754,N_2953);
nand UO_441 (O_441,N_2446,N_2969);
nand UO_442 (O_442,N_2624,N_2777);
and UO_443 (O_443,N_2720,N_2736);
xor UO_444 (O_444,N_2658,N_2575);
nor UO_445 (O_445,N_2477,N_2732);
or UO_446 (O_446,N_2905,N_2533);
nand UO_447 (O_447,N_2523,N_2805);
or UO_448 (O_448,N_2286,N_2743);
or UO_449 (O_449,N_2543,N_2946);
and UO_450 (O_450,N_2695,N_2318);
nor UO_451 (O_451,N_2796,N_2690);
nor UO_452 (O_452,N_2657,N_2319);
nor UO_453 (O_453,N_2680,N_2402);
or UO_454 (O_454,N_2420,N_2320);
and UO_455 (O_455,N_2605,N_2775);
and UO_456 (O_456,N_2685,N_2719);
and UO_457 (O_457,N_2527,N_2808);
or UO_458 (O_458,N_2856,N_2252);
and UO_459 (O_459,N_2396,N_2599);
nor UO_460 (O_460,N_2268,N_2889);
nand UO_461 (O_461,N_2951,N_2370);
nor UO_462 (O_462,N_2369,N_2533);
nor UO_463 (O_463,N_2454,N_2979);
and UO_464 (O_464,N_2440,N_2811);
nor UO_465 (O_465,N_2912,N_2496);
nor UO_466 (O_466,N_2735,N_2683);
or UO_467 (O_467,N_2804,N_2988);
or UO_468 (O_468,N_2339,N_2880);
nand UO_469 (O_469,N_2432,N_2806);
nor UO_470 (O_470,N_2700,N_2954);
and UO_471 (O_471,N_2796,N_2337);
nand UO_472 (O_472,N_2356,N_2770);
or UO_473 (O_473,N_2508,N_2590);
and UO_474 (O_474,N_2309,N_2938);
nor UO_475 (O_475,N_2689,N_2648);
or UO_476 (O_476,N_2853,N_2920);
or UO_477 (O_477,N_2886,N_2989);
nor UO_478 (O_478,N_2655,N_2632);
nor UO_479 (O_479,N_2415,N_2812);
or UO_480 (O_480,N_2712,N_2467);
nand UO_481 (O_481,N_2340,N_2719);
nand UO_482 (O_482,N_2899,N_2954);
or UO_483 (O_483,N_2509,N_2857);
or UO_484 (O_484,N_2276,N_2424);
and UO_485 (O_485,N_2361,N_2770);
nor UO_486 (O_486,N_2849,N_2784);
and UO_487 (O_487,N_2593,N_2823);
nor UO_488 (O_488,N_2730,N_2482);
and UO_489 (O_489,N_2921,N_2397);
or UO_490 (O_490,N_2406,N_2947);
nor UO_491 (O_491,N_2492,N_2957);
nand UO_492 (O_492,N_2653,N_2337);
nand UO_493 (O_493,N_2737,N_2802);
or UO_494 (O_494,N_2781,N_2258);
nand UO_495 (O_495,N_2387,N_2480);
nor UO_496 (O_496,N_2455,N_2881);
and UO_497 (O_497,N_2908,N_2633);
or UO_498 (O_498,N_2992,N_2708);
nand UO_499 (O_499,N_2566,N_2663);
endmodule