module basic_500_3000_500_5_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_251,In_378);
nand U1 (N_1,In_107,In_229);
or U2 (N_2,In_11,In_418);
and U3 (N_3,In_397,In_256);
nand U4 (N_4,In_128,In_263);
or U5 (N_5,In_3,In_350);
nand U6 (N_6,In_476,In_247);
and U7 (N_7,In_351,In_66);
nor U8 (N_8,In_360,In_477);
nor U9 (N_9,In_322,In_432);
nor U10 (N_10,In_490,In_284);
nor U11 (N_11,In_405,In_177);
or U12 (N_12,In_118,In_352);
or U13 (N_13,In_52,In_441);
nand U14 (N_14,In_224,In_345);
or U15 (N_15,In_292,In_121);
xor U16 (N_16,In_148,In_278);
nor U17 (N_17,In_357,In_421);
nor U18 (N_18,In_87,In_40);
nor U19 (N_19,In_23,In_41);
nand U20 (N_20,In_364,In_387);
nor U21 (N_21,In_400,In_275);
nor U22 (N_22,In_457,In_332);
and U23 (N_23,In_102,In_307);
nor U24 (N_24,In_17,In_4);
and U25 (N_25,In_283,In_460);
nand U26 (N_26,In_308,In_205);
nor U27 (N_27,In_424,In_346);
nand U28 (N_28,In_185,In_150);
or U29 (N_29,In_51,In_15);
and U30 (N_30,In_483,In_172);
and U31 (N_31,In_295,In_59);
or U32 (N_32,In_272,In_134);
and U33 (N_33,In_184,In_138);
or U34 (N_34,In_39,In_237);
nor U35 (N_35,In_293,In_402);
or U36 (N_36,In_214,In_57);
and U37 (N_37,In_408,In_60);
nand U38 (N_38,In_277,In_190);
nor U39 (N_39,In_16,In_238);
nand U40 (N_40,In_88,In_252);
or U41 (N_41,In_474,In_62);
nor U42 (N_42,In_69,In_494);
and U43 (N_43,In_200,In_149);
nor U44 (N_44,In_393,In_93);
nand U45 (N_45,In_168,In_466);
nor U46 (N_46,In_188,In_489);
and U47 (N_47,In_246,In_426);
nand U48 (N_48,In_410,In_367);
nand U49 (N_49,In_442,In_161);
nor U50 (N_50,In_5,In_314);
nor U51 (N_51,In_199,In_461);
nor U52 (N_52,In_266,In_279);
nand U53 (N_53,In_301,In_430);
or U54 (N_54,In_320,In_427);
nand U55 (N_55,In_328,In_486);
nor U56 (N_56,In_89,In_13);
and U57 (N_57,In_385,In_217);
or U58 (N_58,In_10,In_201);
or U59 (N_59,In_376,In_108);
and U60 (N_60,In_287,In_395);
nor U61 (N_61,In_222,In_250);
nor U62 (N_62,In_499,In_319);
xor U63 (N_63,In_428,In_475);
nor U64 (N_64,In_331,In_115);
xor U65 (N_65,In_32,In_303);
or U66 (N_66,In_391,In_80);
nor U67 (N_67,In_288,In_249);
and U68 (N_68,In_462,In_392);
nor U69 (N_69,In_174,In_416);
nor U70 (N_70,In_338,In_68);
and U71 (N_71,In_167,In_198);
and U72 (N_72,In_409,In_9);
and U73 (N_73,In_194,In_444);
or U74 (N_74,In_152,In_182);
and U75 (N_75,In_139,In_132);
nand U76 (N_76,In_339,In_459);
and U77 (N_77,In_223,In_101);
xor U78 (N_78,In_452,In_248);
or U79 (N_79,In_226,In_349);
or U80 (N_80,In_12,In_394);
and U81 (N_81,In_470,In_389);
nor U82 (N_82,In_267,In_404);
and U83 (N_83,In_358,In_29);
and U84 (N_84,In_333,In_24);
or U85 (N_85,In_334,In_342);
nand U86 (N_86,In_35,In_463);
nor U87 (N_87,In_82,In_399);
nor U88 (N_88,In_264,In_329);
or U89 (N_89,In_173,In_56);
nor U90 (N_90,In_326,In_330);
or U91 (N_91,In_47,In_240);
and U92 (N_92,In_99,In_305);
or U93 (N_93,In_407,In_160);
nand U94 (N_94,In_197,In_91);
nor U95 (N_95,In_135,In_164);
and U96 (N_96,In_276,In_242);
and U97 (N_97,In_447,In_294);
or U98 (N_98,In_218,In_163);
and U99 (N_99,In_96,In_372);
xor U100 (N_100,In_370,In_144);
and U101 (N_101,In_95,In_113);
and U102 (N_102,In_245,In_335);
or U103 (N_103,In_493,In_44);
and U104 (N_104,In_210,In_344);
or U105 (N_105,In_446,In_384);
and U106 (N_106,In_481,In_46);
nor U107 (N_107,In_285,In_336);
or U108 (N_108,In_316,In_231);
and U109 (N_109,In_390,In_317);
nor U110 (N_110,In_123,In_219);
and U111 (N_111,In_371,In_431);
nor U112 (N_112,In_73,In_383);
nor U113 (N_113,In_196,In_497);
or U114 (N_114,In_20,In_171);
nor U115 (N_115,In_122,In_456);
nand U116 (N_116,In_398,In_154);
nand U117 (N_117,In_420,In_380);
nand U118 (N_118,In_175,In_147);
or U119 (N_119,In_119,In_103);
nand U120 (N_120,In_162,In_45);
or U121 (N_121,In_449,In_443);
and U122 (N_122,In_232,In_465);
or U123 (N_123,In_487,In_221);
nor U124 (N_124,In_381,In_236);
and U125 (N_125,In_243,In_469);
nand U126 (N_126,In_419,In_77);
or U127 (N_127,In_100,In_327);
nand U128 (N_128,In_433,In_270);
or U129 (N_129,In_348,In_434);
nand U130 (N_130,In_300,In_120);
nor U131 (N_131,In_206,In_58);
nand U132 (N_132,In_435,In_453);
nand U133 (N_133,In_53,In_268);
nand U134 (N_134,In_362,In_423);
nor U135 (N_135,In_299,In_67);
or U136 (N_136,In_480,In_176);
or U137 (N_137,In_124,In_425);
or U138 (N_138,In_208,In_366);
and U139 (N_139,In_417,In_415);
and U140 (N_140,In_166,In_216);
or U141 (N_141,In_396,In_375);
or U142 (N_142,In_125,In_233);
or U143 (N_143,In_359,In_63);
nand U144 (N_144,In_261,In_323);
nand U145 (N_145,In_356,In_92);
nor U146 (N_146,In_178,In_450);
nor U147 (N_147,In_141,In_215);
nor U148 (N_148,In_186,In_413);
and U149 (N_149,In_290,In_157);
nand U150 (N_150,In_255,In_187);
nor U151 (N_151,In_72,In_145);
nor U152 (N_152,In_355,In_43);
and U153 (N_153,In_491,In_2);
nand U154 (N_154,In_155,In_311);
and U155 (N_155,In_281,In_22);
and U156 (N_156,In_259,In_455);
nor U157 (N_157,In_153,In_468);
or U158 (N_158,In_126,In_291);
nand U159 (N_159,In_209,In_191);
nor U160 (N_160,In_297,In_71);
and U161 (N_161,In_225,In_78);
nand U162 (N_162,In_28,In_373);
and U163 (N_163,In_386,In_492);
nor U164 (N_164,In_239,In_65);
or U165 (N_165,In_411,In_273);
or U166 (N_166,In_143,In_298);
and U167 (N_167,In_388,In_340);
nor U168 (N_168,In_106,In_439);
nand U169 (N_169,In_429,In_484);
nand U170 (N_170,In_265,In_36);
and U171 (N_171,In_79,In_488);
nor U172 (N_172,In_158,In_70);
or U173 (N_173,In_37,In_136);
nor U174 (N_174,In_485,In_84);
xnor U175 (N_175,In_230,In_165);
and U176 (N_176,In_254,In_74);
nor U177 (N_177,In_412,In_61);
nand U178 (N_178,In_271,In_347);
or U179 (N_179,In_104,In_33);
or U180 (N_180,In_114,In_309);
nand U181 (N_181,In_129,In_90);
nand U182 (N_182,In_94,In_26);
nor U183 (N_183,In_133,In_195);
nand U184 (N_184,In_156,In_354);
and U185 (N_185,In_289,In_280);
nand U186 (N_186,In_109,In_207);
or U187 (N_187,In_105,In_81);
or U188 (N_188,In_25,In_262);
nand U189 (N_189,In_151,In_437);
or U190 (N_190,In_498,In_181);
nand U191 (N_191,In_286,In_377);
or U192 (N_192,In_7,In_18);
nor U193 (N_193,In_495,In_50);
nand U194 (N_194,In_142,In_253);
and U195 (N_195,In_54,In_315);
or U196 (N_196,In_260,In_192);
nand U197 (N_197,In_472,In_48);
and U198 (N_198,In_83,In_235);
nand U199 (N_199,In_274,In_14);
xor U200 (N_200,In_30,In_422);
nand U201 (N_201,In_296,In_170);
nand U202 (N_202,In_0,In_21);
nor U203 (N_203,In_130,In_341);
nor U204 (N_204,In_304,In_111);
or U205 (N_205,In_34,In_169);
nand U206 (N_206,In_479,In_343);
and U207 (N_207,In_31,In_179);
nor U208 (N_208,In_76,In_228);
nor U209 (N_209,In_193,In_86);
and U210 (N_210,In_27,In_353);
xor U211 (N_211,In_8,In_258);
nand U212 (N_212,In_306,In_471);
or U213 (N_213,In_365,In_302);
and U214 (N_214,In_213,In_55);
and U215 (N_215,In_440,In_42);
or U216 (N_216,In_401,In_451);
or U217 (N_217,In_203,In_478);
and U218 (N_218,In_212,In_445);
and U219 (N_219,In_382,In_241);
or U220 (N_220,In_180,In_98);
or U221 (N_221,In_202,In_482);
or U222 (N_222,In_436,In_448);
nand U223 (N_223,In_137,In_473);
nand U224 (N_224,In_146,In_75);
and U225 (N_225,In_467,In_313);
or U226 (N_226,In_183,In_282);
nand U227 (N_227,In_97,In_379);
nor U228 (N_228,In_110,In_64);
or U229 (N_229,In_227,In_189);
nand U230 (N_230,In_116,In_318);
nand U231 (N_231,In_244,In_127);
and U232 (N_232,In_406,In_324);
or U233 (N_233,In_369,In_112);
nand U234 (N_234,In_454,In_374);
or U235 (N_235,In_85,In_458);
or U236 (N_236,In_325,In_310);
nand U237 (N_237,In_269,In_312);
nor U238 (N_238,In_361,In_414);
nand U239 (N_239,In_403,In_131);
and U240 (N_240,In_117,In_321);
nor U241 (N_241,In_140,In_257);
or U242 (N_242,In_220,In_368);
or U243 (N_243,In_38,In_19);
xor U244 (N_244,In_496,In_337);
nand U245 (N_245,In_438,In_49);
nand U246 (N_246,In_204,In_6);
or U247 (N_247,In_363,In_159);
nand U248 (N_248,In_464,In_234);
nand U249 (N_249,In_211,In_1);
or U250 (N_250,In_318,In_73);
and U251 (N_251,In_371,In_93);
nor U252 (N_252,In_129,In_52);
or U253 (N_253,In_208,In_239);
and U254 (N_254,In_422,In_37);
nor U255 (N_255,In_7,In_194);
nor U256 (N_256,In_133,In_364);
nor U257 (N_257,In_479,In_496);
xnor U258 (N_258,In_140,In_162);
nand U259 (N_259,In_214,In_292);
and U260 (N_260,In_183,In_200);
nand U261 (N_261,In_253,In_312);
nor U262 (N_262,In_81,In_253);
and U263 (N_263,In_16,In_44);
nand U264 (N_264,In_186,In_406);
or U265 (N_265,In_473,In_255);
nand U266 (N_266,In_349,In_163);
nand U267 (N_267,In_456,In_236);
or U268 (N_268,In_328,In_109);
or U269 (N_269,In_274,In_438);
nor U270 (N_270,In_90,In_491);
nand U271 (N_271,In_192,In_443);
and U272 (N_272,In_127,In_380);
nor U273 (N_273,In_189,In_1);
and U274 (N_274,In_134,In_353);
xnor U275 (N_275,In_42,In_217);
and U276 (N_276,In_79,In_152);
nor U277 (N_277,In_147,In_49);
or U278 (N_278,In_301,In_426);
or U279 (N_279,In_143,In_0);
or U280 (N_280,In_130,In_277);
xnor U281 (N_281,In_107,In_454);
and U282 (N_282,In_235,In_103);
or U283 (N_283,In_145,In_418);
or U284 (N_284,In_411,In_496);
and U285 (N_285,In_39,In_313);
or U286 (N_286,In_240,In_94);
nor U287 (N_287,In_294,In_412);
nor U288 (N_288,In_12,In_152);
xnor U289 (N_289,In_300,In_349);
nand U290 (N_290,In_478,In_417);
or U291 (N_291,In_46,In_8);
nor U292 (N_292,In_153,In_172);
and U293 (N_293,In_103,In_475);
nor U294 (N_294,In_296,In_19);
nor U295 (N_295,In_40,In_280);
and U296 (N_296,In_307,In_35);
nor U297 (N_297,In_143,In_413);
and U298 (N_298,In_198,In_218);
and U299 (N_299,In_314,In_298);
nor U300 (N_300,In_381,In_231);
and U301 (N_301,In_281,In_33);
nor U302 (N_302,In_126,In_231);
or U303 (N_303,In_358,In_457);
or U304 (N_304,In_344,In_209);
nor U305 (N_305,In_19,In_336);
and U306 (N_306,In_17,In_469);
or U307 (N_307,In_199,In_11);
and U308 (N_308,In_332,In_459);
nand U309 (N_309,In_272,In_103);
and U310 (N_310,In_117,In_191);
nor U311 (N_311,In_344,In_449);
and U312 (N_312,In_260,In_14);
nor U313 (N_313,In_376,In_296);
or U314 (N_314,In_75,In_399);
nand U315 (N_315,In_391,In_425);
nand U316 (N_316,In_320,In_117);
or U317 (N_317,In_370,In_372);
or U318 (N_318,In_388,In_45);
or U319 (N_319,In_177,In_174);
nor U320 (N_320,In_329,In_199);
or U321 (N_321,In_322,In_95);
nand U322 (N_322,In_116,In_86);
nand U323 (N_323,In_411,In_192);
xor U324 (N_324,In_209,In_400);
xnor U325 (N_325,In_270,In_386);
nand U326 (N_326,In_291,In_258);
and U327 (N_327,In_49,In_315);
or U328 (N_328,In_347,In_189);
nand U329 (N_329,In_196,In_296);
and U330 (N_330,In_407,In_350);
or U331 (N_331,In_436,In_119);
and U332 (N_332,In_453,In_66);
and U333 (N_333,In_173,In_161);
nand U334 (N_334,In_172,In_202);
nand U335 (N_335,In_442,In_137);
nor U336 (N_336,In_135,In_277);
nor U337 (N_337,In_56,In_441);
nor U338 (N_338,In_188,In_224);
and U339 (N_339,In_436,In_427);
or U340 (N_340,In_395,In_469);
or U341 (N_341,In_334,In_228);
and U342 (N_342,In_439,In_39);
nor U343 (N_343,In_20,In_396);
or U344 (N_344,In_57,In_420);
or U345 (N_345,In_173,In_445);
nor U346 (N_346,In_118,In_408);
or U347 (N_347,In_249,In_475);
and U348 (N_348,In_32,In_294);
and U349 (N_349,In_361,In_47);
and U350 (N_350,In_195,In_31);
nand U351 (N_351,In_434,In_65);
and U352 (N_352,In_125,In_246);
nor U353 (N_353,In_389,In_327);
nand U354 (N_354,In_139,In_419);
or U355 (N_355,In_240,In_423);
and U356 (N_356,In_305,In_345);
nand U357 (N_357,In_327,In_123);
and U358 (N_358,In_488,In_441);
nand U359 (N_359,In_373,In_147);
nor U360 (N_360,In_272,In_87);
nor U361 (N_361,In_40,In_302);
nor U362 (N_362,In_438,In_286);
and U363 (N_363,In_318,In_276);
nand U364 (N_364,In_438,In_417);
nor U365 (N_365,In_395,In_397);
and U366 (N_366,In_300,In_159);
nor U367 (N_367,In_70,In_409);
and U368 (N_368,In_71,In_27);
or U369 (N_369,In_199,In_398);
or U370 (N_370,In_367,In_493);
nor U371 (N_371,In_484,In_411);
or U372 (N_372,In_480,In_260);
nor U373 (N_373,In_412,In_290);
nand U374 (N_374,In_134,In_347);
and U375 (N_375,In_139,In_83);
or U376 (N_376,In_52,In_475);
xor U377 (N_377,In_401,In_109);
and U378 (N_378,In_458,In_81);
or U379 (N_379,In_444,In_8);
or U380 (N_380,In_99,In_285);
xnor U381 (N_381,In_475,In_3);
or U382 (N_382,In_18,In_44);
and U383 (N_383,In_201,In_448);
or U384 (N_384,In_7,In_27);
or U385 (N_385,In_307,In_161);
or U386 (N_386,In_140,In_342);
and U387 (N_387,In_34,In_174);
or U388 (N_388,In_492,In_62);
nor U389 (N_389,In_180,In_335);
or U390 (N_390,In_248,In_179);
nand U391 (N_391,In_407,In_5);
nor U392 (N_392,In_76,In_11);
and U393 (N_393,In_331,In_186);
nand U394 (N_394,In_28,In_288);
and U395 (N_395,In_393,In_203);
and U396 (N_396,In_400,In_337);
and U397 (N_397,In_207,In_5);
nand U398 (N_398,In_346,In_402);
nor U399 (N_399,In_456,In_140);
or U400 (N_400,In_38,In_145);
nand U401 (N_401,In_403,In_41);
and U402 (N_402,In_139,In_71);
or U403 (N_403,In_135,In_202);
and U404 (N_404,In_278,In_420);
or U405 (N_405,In_482,In_258);
or U406 (N_406,In_153,In_250);
and U407 (N_407,In_330,In_449);
xor U408 (N_408,In_298,In_206);
nor U409 (N_409,In_28,In_384);
or U410 (N_410,In_0,In_342);
and U411 (N_411,In_453,In_275);
nor U412 (N_412,In_236,In_329);
nor U413 (N_413,In_211,In_112);
and U414 (N_414,In_468,In_471);
or U415 (N_415,In_385,In_136);
or U416 (N_416,In_275,In_346);
and U417 (N_417,In_184,In_372);
and U418 (N_418,In_269,In_384);
and U419 (N_419,In_278,In_79);
and U420 (N_420,In_349,In_467);
and U421 (N_421,In_4,In_97);
nor U422 (N_422,In_444,In_259);
and U423 (N_423,In_90,In_292);
nand U424 (N_424,In_256,In_80);
and U425 (N_425,In_498,In_169);
and U426 (N_426,In_262,In_1);
nor U427 (N_427,In_429,In_131);
or U428 (N_428,In_489,In_339);
or U429 (N_429,In_298,In_441);
nand U430 (N_430,In_326,In_262);
and U431 (N_431,In_275,In_485);
nand U432 (N_432,In_359,In_38);
nor U433 (N_433,In_336,In_361);
or U434 (N_434,In_266,In_285);
nand U435 (N_435,In_266,In_16);
and U436 (N_436,In_412,In_21);
or U437 (N_437,In_236,In_96);
and U438 (N_438,In_454,In_234);
nor U439 (N_439,In_97,In_80);
nand U440 (N_440,In_318,In_489);
or U441 (N_441,In_212,In_317);
and U442 (N_442,In_278,In_117);
nor U443 (N_443,In_277,In_343);
nand U444 (N_444,In_136,In_333);
nand U445 (N_445,In_348,In_185);
and U446 (N_446,In_427,In_343);
or U447 (N_447,In_170,In_371);
or U448 (N_448,In_225,In_89);
or U449 (N_449,In_482,In_252);
and U450 (N_450,In_25,In_38);
nor U451 (N_451,In_30,In_200);
xnor U452 (N_452,In_420,In_106);
nor U453 (N_453,In_126,In_257);
nor U454 (N_454,In_81,In_484);
nor U455 (N_455,In_286,In_456);
nor U456 (N_456,In_266,In_496);
nand U457 (N_457,In_100,In_392);
and U458 (N_458,In_478,In_492);
and U459 (N_459,In_391,In_153);
or U460 (N_460,In_186,In_404);
and U461 (N_461,In_306,In_181);
and U462 (N_462,In_2,In_238);
nor U463 (N_463,In_69,In_352);
or U464 (N_464,In_456,In_295);
nor U465 (N_465,In_151,In_334);
nor U466 (N_466,In_206,In_485);
nor U467 (N_467,In_125,In_17);
and U468 (N_468,In_258,In_480);
and U469 (N_469,In_345,In_275);
or U470 (N_470,In_331,In_432);
xnor U471 (N_471,In_277,In_317);
or U472 (N_472,In_282,In_338);
and U473 (N_473,In_164,In_281);
and U474 (N_474,In_95,In_231);
nand U475 (N_475,In_24,In_295);
or U476 (N_476,In_464,In_303);
nand U477 (N_477,In_230,In_272);
nor U478 (N_478,In_343,In_383);
nor U479 (N_479,In_95,In_423);
nor U480 (N_480,In_222,In_13);
nor U481 (N_481,In_311,In_152);
and U482 (N_482,In_58,In_251);
and U483 (N_483,In_14,In_336);
and U484 (N_484,In_463,In_76);
and U485 (N_485,In_450,In_482);
nor U486 (N_486,In_77,In_53);
and U487 (N_487,In_206,In_204);
nor U488 (N_488,In_362,In_492);
or U489 (N_489,In_370,In_129);
nor U490 (N_490,In_193,In_90);
nand U491 (N_491,In_212,In_408);
nand U492 (N_492,In_412,In_321);
nor U493 (N_493,In_377,In_498);
and U494 (N_494,In_366,In_342);
or U495 (N_495,In_461,In_459);
xnor U496 (N_496,In_90,In_314);
or U497 (N_497,In_113,In_370);
xnor U498 (N_498,In_23,In_117);
nand U499 (N_499,In_406,In_164);
and U500 (N_500,In_465,In_270);
nor U501 (N_501,In_331,In_48);
or U502 (N_502,In_75,In_32);
nor U503 (N_503,In_469,In_374);
nand U504 (N_504,In_357,In_374);
and U505 (N_505,In_358,In_368);
xnor U506 (N_506,In_141,In_487);
nor U507 (N_507,In_477,In_251);
nor U508 (N_508,In_147,In_95);
and U509 (N_509,In_366,In_439);
and U510 (N_510,In_453,In_303);
nand U511 (N_511,In_183,In_201);
nor U512 (N_512,In_317,In_188);
nor U513 (N_513,In_369,In_378);
nand U514 (N_514,In_463,In_247);
nor U515 (N_515,In_445,In_164);
and U516 (N_516,In_198,In_247);
nor U517 (N_517,In_65,In_363);
nor U518 (N_518,In_484,In_48);
or U519 (N_519,In_396,In_298);
and U520 (N_520,In_235,In_461);
or U521 (N_521,In_139,In_180);
nor U522 (N_522,In_306,In_162);
and U523 (N_523,In_301,In_40);
and U524 (N_524,In_64,In_242);
and U525 (N_525,In_420,In_240);
nor U526 (N_526,In_94,In_33);
and U527 (N_527,In_336,In_104);
nand U528 (N_528,In_130,In_362);
nor U529 (N_529,In_371,In_174);
nand U530 (N_530,In_498,In_175);
or U531 (N_531,In_416,In_444);
or U532 (N_532,In_8,In_396);
nand U533 (N_533,In_18,In_255);
or U534 (N_534,In_457,In_272);
nor U535 (N_535,In_109,In_173);
and U536 (N_536,In_32,In_438);
or U537 (N_537,In_15,In_131);
or U538 (N_538,In_389,In_118);
nor U539 (N_539,In_285,In_294);
and U540 (N_540,In_92,In_135);
nand U541 (N_541,In_230,In_10);
and U542 (N_542,In_376,In_464);
or U543 (N_543,In_458,In_347);
and U544 (N_544,In_430,In_21);
nand U545 (N_545,In_109,In_331);
nor U546 (N_546,In_305,In_314);
nor U547 (N_547,In_300,In_117);
nor U548 (N_548,In_188,In_391);
nand U549 (N_549,In_300,In_447);
or U550 (N_550,In_461,In_251);
or U551 (N_551,In_496,In_302);
nor U552 (N_552,In_193,In_337);
or U553 (N_553,In_206,In_116);
nand U554 (N_554,In_274,In_80);
and U555 (N_555,In_42,In_446);
and U556 (N_556,In_91,In_152);
and U557 (N_557,In_372,In_71);
nand U558 (N_558,In_438,In_268);
nor U559 (N_559,In_140,In_330);
nor U560 (N_560,In_155,In_106);
nand U561 (N_561,In_130,In_385);
nor U562 (N_562,In_131,In_238);
and U563 (N_563,In_87,In_318);
nand U564 (N_564,In_35,In_168);
or U565 (N_565,In_65,In_133);
nand U566 (N_566,In_277,In_390);
and U567 (N_567,In_125,In_137);
or U568 (N_568,In_42,In_165);
nand U569 (N_569,In_487,In_173);
or U570 (N_570,In_134,In_178);
and U571 (N_571,In_407,In_368);
nor U572 (N_572,In_320,In_468);
nor U573 (N_573,In_273,In_9);
xor U574 (N_574,In_382,In_343);
nand U575 (N_575,In_69,In_98);
nor U576 (N_576,In_357,In_265);
nand U577 (N_577,In_73,In_199);
or U578 (N_578,In_392,In_195);
nor U579 (N_579,In_381,In_9);
nor U580 (N_580,In_44,In_405);
or U581 (N_581,In_127,In_248);
and U582 (N_582,In_226,In_409);
nor U583 (N_583,In_458,In_357);
xnor U584 (N_584,In_371,In_280);
and U585 (N_585,In_27,In_43);
and U586 (N_586,In_403,In_304);
nor U587 (N_587,In_301,In_382);
nor U588 (N_588,In_283,In_87);
nor U589 (N_589,In_493,In_116);
nand U590 (N_590,In_337,In_121);
and U591 (N_591,In_97,In_361);
nand U592 (N_592,In_238,In_319);
and U593 (N_593,In_427,In_440);
xnor U594 (N_594,In_40,In_365);
nand U595 (N_595,In_425,In_24);
and U596 (N_596,In_69,In_167);
and U597 (N_597,In_97,In_367);
and U598 (N_598,In_494,In_246);
nor U599 (N_599,In_140,In_322);
and U600 (N_600,N_540,N_228);
or U601 (N_601,N_437,N_492);
nor U602 (N_602,N_290,N_533);
or U603 (N_603,N_346,N_377);
and U604 (N_604,N_269,N_335);
nand U605 (N_605,N_587,N_68);
or U606 (N_606,N_327,N_454);
or U607 (N_607,N_300,N_432);
nor U608 (N_608,N_347,N_312);
nor U609 (N_609,N_419,N_283);
xor U610 (N_610,N_317,N_134);
nand U611 (N_611,N_567,N_241);
or U612 (N_612,N_385,N_339);
nor U613 (N_613,N_400,N_93);
nand U614 (N_614,N_445,N_135);
xnor U615 (N_615,N_167,N_13);
or U616 (N_616,N_5,N_364);
or U617 (N_617,N_548,N_491);
and U618 (N_618,N_514,N_158);
nor U619 (N_619,N_395,N_331);
nor U620 (N_620,N_41,N_599);
or U621 (N_621,N_554,N_442);
and U622 (N_622,N_176,N_74);
nor U623 (N_623,N_150,N_114);
nor U624 (N_624,N_305,N_531);
nand U625 (N_625,N_577,N_596);
nand U626 (N_626,N_45,N_69);
nor U627 (N_627,N_108,N_537);
or U628 (N_628,N_368,N_384);
nor U629 (N_629,N_91,N_512);
and U630 (N_630,N_387,N_80);
or U631 (N_631,N_482,N_382);
and U632 (N_632,N_216,N_354);
or U633 (N_633,N_280,N_133);
nand U634 (N_634,N_575,N_55);
or U635 (N_635,N_120,N_325);
nand U636 (N_636,N_594,N_304);
nand U637 (N_637,N_337,N_15);
and U638 (N_638,N_408,N_62);
or U639 (N_639,N_536,N_566);
nand U640 (N_640,N_348,N_527);
nand U641 (N_641,N_119,N_397);
and U642 (N_642,N_451,N_379);
nand U643 (N_643,N_414,N_8);
and U644 (N_644,N_574,N_593);
and U645 (N_645,N_205,N_388);
and U646 (N_646,N_38,N_417);
or U647 (N_647,N_281,N_488);
and U648 (N_648,N_207,N_340);
and U649 (N_649,N_350,N_195);
nand U650 (N_650,N_155,N_362);
and U651 (N_651,N_56,N_129);
and U652 (N_652,N_591,N_507);
or U653 (N_653,N_77,N_39);
nor U654 (N_654,N_374,N_505);
or U655 (N_655,N_578,N_213);
nor U656 (N_656,N_440,N_433);
nor U657 (N_657,N_307,N_265);
and U658 (N_658,N_394,N_84);
or U659 (N_659,N_495,N_321);
and U660 (N_660,N_296,N_209);
and U661 (N_661,N_423,N_163);
nand U662 (N_662,N_494,N_65);
nand U663 (N_663,N_552,N_588);
nor U664 (N_664,N_34,N_324);
nand U665 (N_665,N_226,N_7);
or U666 (N_666,N_219,N_571);
and U667 (N_667,N_192,N_510);
or U668 (N_668,N_376,N_351);
or U669 (N_669,N_366,N_358);
nor U670 (N_670,N_30,N_378);
and U671 (N_671,N_391,N_272);
nand U672 (N_672,N_220,N_54);
nand U673 (N_673,N_130,N_137);
and U674 (N_674,N_489,N_421);
xnor U675 (N_675,N_48,N_76);
and U676 (N_676,N_590,N_123);
or U677 (N_677,N_284,N_581);
nand U678 (N_678,N_103,N_586);
or U679 (N_679,N_106,N_457);
or U680 (N_680,N_169,N_122);
and U681 (N_681,N_263,N_172);
or U682 (N_682,N_323,N_89);
or U683 (N_683,N_401,N_22);
nor U684 (N_684,N_233,N_341);
nand U685 (N_685,N_439,N_496);
nand U686 (N_686,N_471,N_246);
and U687 (N_687,N_199,N_411);
nor U688 (N_688,N_383,N_334);
or U689 (N_689,N_273,N_203);
nor U690 (N_690,N_434,N_493);
nand U691 (N_691,N_144,N_124);
or U692 (N_692,N_259,N_468);
nor U693 (N_693,N_565,N_483);
nand U694 (N_694,N_201,N_486);
nor U695 (N_695,N_168,N_298);
nor U696 (N_696,N_239,N_550);
nand U697 (N_697,N_63,N_118);
nand U698 (N_698,N_478,N_104);
or U699 (N_699,N_452,N_18);
nand U700 (N_700,N_35,N_345);
and U701 (N_701,N_184,N_116);
nand U702 (N_702,N_36,N_474);
xnor U703 (N_703,N_243,N_287);
or U704 (N_704,N_245,N_174);
nand U705 (N_705,N_85,N_266);
nand U706 (N_706,N_412,N_198);
nor U707 (N_707,N_541,N_240);
or U708 (N_708,N_82,N_186);
and U709 (N_709,N_557,N_589);
or U710 (N_710,N_465,N_110);
or U711 (N_711,N_210,N_534);
nand U712 (N_712,N_399,N_185);
or U713 (N_713,N_293,N_470);
or U714 (N_714,N_420,N_154);
nor U715 (N_715,N_299,N_227);
or U716 (N_716,N_455,N_173);
xnor U717 (N_717,N_458,N_326);
nor U718 (N_718,N_515,N_329);
nand U719 (N_719,N_128,N_285);
nor U720 (N_720,N_232,N_592);
or U721 (N_721,N_583,N_2);
and U722 (N_722,N_328,N_171);
or U723 (N_723,N_286,N_214);
and U724 (N_724,N_490,N_431);
and U725 (N_725,N_224,N_70);
or U726 (N_726,N_279,N_102);
nor U727 (N_727,N_136,N_509);
nor U728 (N_728,N_121,N_462);
and U729 (N_729,N_142,N_559);
nand U730 (N_730,N_161,N_314);
or U731 (N_731,N_436,N_398);
or U732 (N_732,N_464,N_26);
and U733 (N_733,N_407,N_59);
and U734 (N_734,N_258,N_107);
nor U735 (N_735,N_125,N_278);
nand U736 (N_736,N_0,N_276);
nor U737 (N_737,N_580,N_369);
and U738 (N_738,N_200,N_543);
nor U739 (N_739,N_160,N_37);
and U740 (N_740,N_242,N_572);
xor U741 (N_741,N_4,N_211);
nor U742 (N_742,N_373,N_126);
or U743 (N_743,N_149,N_547);
nand U744 (N_744,N_99,N_585);
nand U745 (N_745,N_367,N_532);
nor U746 (N_746,N_513,N_381);
or U747 (N_747,N_526,N_560);
or U748 (N_748,N_179,N_556);
nor U749 (N_749,N_467,N_579);
or U750 (N_750,N_310,N_569);
nor U751 (N_751,N_426,N_257);
nand U752 (N_752,N_389,N_318);
and U753 (N_753,N_487,N_271);
and U754 (N_754,N_197,N_429);
nor U755 (N_755,N_44,N_562);
xnor U756 (N_756,N_180,N_223);
nand U757 (N_757,N_217,N_584);
nand U758 (N_758,N_274,N_191);
nor U759 (N_759,N_222,N_415);
nor U760 (N_760,N_444,N_520);
xnor U761 (N_761,N_294,N_42);
and U762 (N_762,N_375,N_143);
nand U763 (N_763,N_58,N_189);
nand U764 (N_764,N_29,N_190);
nand U765 (N_765,N_88,N_275);
and U766 (N_766,N_525,N_81);
and U767 (N_767,N_320,N_11);
nand U768 (N_768,N_109,N_98);
and U769 (N_769,N_270,N_450);
and U770 (N_770,N_162,N_582);
or U771 (N_771,N_316,N_221);
nand U772 (N_772,N_477,N_338);
and U773 (N_773,N_466,N_313);
or U774 (N_774,N_459,N_508);
or U775 (N_775,N_268,N_16);
or U776 (N_776,N_9,N_255);
nand U777 (N_777,N_32,N_469);
or U778 (N_778,N_256,N_563);
and U779 (N_779,N_315,N_24);
and U780 (N_780,N_46,N_502);
xor U781 (N_781,N_595,N_261);
nor U782 (N_782,N_330,N_542);
or U783 (N_783,N_21,N_31);
nor U784 (N_784,N_441,N_598);
or U785 (N_785,N_430,N_500);
or U786 (N_786,N_164,N_178);
and U787 (N_787,N_343,N_40);
or U788 (N_788,N_427,N_518);
nand U789 (N_789,N_237,N_402);
or U790 (N_790,N_472,N_75);
and U791 (N_791,N_396,N_19);
nand U792 (N_792,N_524,N_139);
or U793 (N_793,N_530,N_175);
nor U794 (N_794,N_64,N_66);
and U795 (N_795,N_561,N_1);
nor U796 (N_796,N_208,N_410);
and U797 (N_797,N_342,N_292);
nand U798 (N_798,N_576,N_244);
nand U799 (N_799,N_3,N_463);
or U800 (N_800,N_511,N_28);
xnor U801 (N_801,N_253,N_181);
or U802 (N_802,N_60,N_86);
nor U803 (N_803,N_87,N_115);
nor U804 (N_804,N_83,N_359);
nor U805 (N_805,N_202,N_460);
nor U806 (N_806,N_188,N_504);
and U807 (N_807,N_117,N_165);
nand U808 (N_808,N_564,N_10);
or U809 (N_809,N_302,N_476);
or U810 (N_810,N_418,N_61);
nand U811 (N_811,N_353,N_573);
or U812 (N_812,N_33,N_52);
nor U813 (N_813,N_291,N_438);
or U814 (N_814,N_344,N_473);
and U815 (N_815,N_73,N_308);
nand U816 (N_816,N_355,N_236);
nor U817 (N_817,N_204,N_425);
and U818 (N_818,N_146,N_311);
and U819 (N_819,N_235,N_523);
and U820 (N_820,N_132,N_360);
and U821 (N_821,N_424,N_53);
nand U822 (N_822,N_157,N_538);
nand U823 (N_823,N_372,N_371);
or U824 (N_824,N_282,N_306);
or U825 (N_825,N_141,N_262);
xor U826 (N_826,N_447,N_72);
or U827 (N_827,N_558,N_250);
nand U828 (N_828,N_303,N_295);
and U829 (N_829,N_156,N_551);
nor U830 (N_830,N_416,N_481);
nand U831 (N_831,N_361,N_101);
or U832 (N_832,N_230,N_79);
and U833 (N_833,N_322,N_349);
and U834 (N_834,N_229,N_506);
or U835 (N_835,N_529,N_297);
and U836 (N_836,N_96,N_249);
and U837 (N_837,N_71,N_446);
nor U838 (N_838,N_461,N_553);
and U839 (N_839,N_597,N_555);
nand U840 (N_840,N_428,N_333);
and U841 (N_841,N_409,N_545);
or U842 (N_842,N_570,N_549);
xor U843 (N_843,N_159,N_215);
nor U844 (N_844,N_365,N_100);
nand U845 (N_845,N_544,N_568);
nor U846 (N_846,N_138,N_153);
nor U847 (N_847,N_51,N_519);
nor U848 (N_848,N_539,N_497);
or U849 (N_849,N_480,N_131);
nor U850 (N_850,N_499,N_252);
nand U851 (N_851,N_498,N_196);
nor U852 (N_852,N_289,N_112);
or U853 (N_853,N_43,N_264);
nor U854 (N_854,N_435,N_521);
nor U855 (N_855,N_503,N_363);
and U856 (N_856,N_288,N_95);
nor U857 (N_857,N_248,N_78);
and U858 (N_858,N_166,N_92);
nand U859 (N_859,N_17,N_522);
and U860 (N_860,N_145,N_127);
nor U861 (N_861,N_111,N_475);
nor U862 (N_862,N_251,N_50);
and U863 (N_863,N_443,N_27);
or U864 (N_864,N_247,N_456);
and U865 (N_865,N_6,N_151);
nor U866 (N_866,N_218,N_309);
nand U867 (N_867,N_140,N_113);
nor U868 (N_868,N_393,N_182);
and U869 (N_869,N_234,N_301);
and U870 (N_870,N_23,N_206);
nand U871 (N_871,N_267,N_453);
nor U872 (N_872,N_336,N_332);
nand U873 (N_873,N_194,N_485);
or U874 (N_874,N_528,N_516);
or U875 (N_875,N_413,N_277);
xnor U876 (N_876,N_14,N_448);
or U877 (N_877,N_170,N_422);
or U878 (N_878,N_193,N_57);
nand U879 (N_879,N_254,N_148);
nor U880 (N_880,N_183,N_20);
nand U881 (N_881,N_535,N_386);
nor U882 (N_882,N_94,N_212);
nor U883 (N_883,N_405,N_90);
or U884 (N_884,N_152,N_231);
nand U885 (N_885,N_238,N_25);
nand U886 (N_886,N_352,N_356);
nor U887 (N_887,N_380,N_187);
nor U888 (N_888,N_319,N_392);
or U889 (N_889,N_546,N_357);
nand U890 (N_890,N_177,N_225);
nor U891 (N_891,N_449,N_260);
and U892 (N_892,N_404,N_67);
or U893 (N_893,N_484,N_406);
and U894 (N_894,N_49,N_517);
nand U895 (N_895,N_105,N_403);
nand U896 (N_896,N_147,N_12);
nand U897 (N_897,N_47,N_370);
nand U898 (N_898,N_501,N_390);
nand U899 (N_899,N_479,N_97);
nor U900 (N_900,N_118,N_529);
or U901 (N_901,N_142,N_539);
and U902 (N_902,N_221,N_244);
nand U903 (N_903,N_574,N_415);
nor U904 (N_904,N_545,N_439);
nand U905 (N_905,N_35,N_481);
or U906 (N_906,N_521,N_427);
nor U907 (N_907,N_412,N_258);
or U908 (N_908,N_496,N_561);
nor U909 (N_909,N_406,N_384);
and U910 (N_910,N_471,N_210);
nor U911 (N_911,N_542,N_32);
or U912 (N_912,N_158,N_87);
nand U913 (N_913,N_506,N_457);
nor U914 (N_914,N_33,N_371);
or U915 (N_915,N_73,N_582);
or U916 (N_916,N_542,N_497);
nor U917 (N_917,N_365,N_226);
nand U918 (N_918,N_122,N_250);
and U919 (N_919,N_283,N_395);
and U920 (N_920,N_438,N_186);
or U921 (N_921,N_432,N_83);
or U922 (N_922,N_456,N_212);
and U923 (N_923,N_87,N_381);
nand U924 (N_924,N_532,N_403);
or U925 (N_925,N_256,N_73);
or U926 (N_926,N_329,N_501);
or U927 (N_927,N_382,N_312);
nand U928 (N_928,N_20,N_338);
or U929 (N_929,N_414,N_530);
and U930 (N_930,N_424,N_123);
or U931 (N_931,N_355,N_7);
and U932 (N_932,N_484,N_459);
or U933 (N_933,N_596,N_187);
and U934 (N_934,N_248,N_221);
and U935 (N_935,N_103,N_294);
nand U936 (N_936,N_204,N_360);
or U937 (N_937,N_325,N_433);
or U938 (N_938,N_302,N_154);
nor U939 (N_939,N_491,N_110);
or U940 (N_940,N_91,N_495);
and U941 (N_941,N_483,N_365);
and U942 (N_942,N_405,N_574);
and U943 (N_943,N_387,N_544);
nand U944 (N_944,N_468,N_383);
nand U945 (N_945,N_267,N_237);
nor U946 (N_946,N_141,N_466);
nor U947 (N_947,N_492,N_498);
and U948 (N_948,N_431,N_415);
xnor U949 (N_949,N_438,N_564);
nor U950 (N_950,N_491,N_298);
and U951 (N_951,N_404,N_265);
nor U952 (N_952,N_160,N_175);
nor U953 (N_953,N_66,N_559);
and U954 (N_954,N_443,N_157);
and U955 (N_955,N_126,N_24);
nand U956 (N_956,N_200,N_9);
nor U957 (N_957,N_296,N_481);
nand U958 (N_958,N_181,N_185);
nor U959 (N_959,N_507,N_392);
and U960 (N_960,N_435,N_334);
or U961 (N_961,N_494,N_260);
nand U962 (N_962,N_361,N_153);
nand U963 (N_963,N_81,N_530);
or U964 (N_964,N_573,N_455);
or U965 (N_965,N_170,N_73);
or U966 (N_966,N_521,N_148);
nor U967 (N_967,N_216,N_187);
nor U968 (N_968,N_90,N_42);
nor U969 (N_969,N_191,N_159);
nand U970 (N_970,N_209,N_122);
and U971 (N_971,N_172,N_189);
nor U972 (N_972,N_566,N_479);
or U973 (N_973,N_291,N_517);
nor U974 (N_974,N_232,N_478);
or U975 (N_975,N_392,N_321);
and U976 (N_976,N_500,N_363);
nor U977 (N_977,N_41,N_391);
nand U978 (N_978,N_309,N_114);
nand U979 (N_979,N_544,N_554);
or U980 (N_980,N_398,N_337);
nand U981 (N_981,N_532,N_366);
nand U982 (N_982,N_473,N_242);
nand U983 (N_983,N_15,N_420);
or U984 (N_984,N_519,N_402);
nor U985 (N_985,N_121,N_301);
or U986 (N_986,N_401,N_314);
or U987 (N_987,N_522,N_457);
nor U988 (N_988,N_180,N_326);
and U989 (N_989,N_190,N_561);
and U990 (N_990,N_148,N_474);
or U991 (N_991,N_491,N_279);
and U992 (N_992,N_105,N_554);
nand U993 (N_993,N_42,N_108);
and U994 (N_994,N_36,N_388);
or U995 (N_995,N_345,N_259);
nor U996 (N_996,N_265,N_592);
nand U997 (N_997,N_27,N_382);
nor U998 (N_998,N_221,N_412);
or U999 (N_999,N_139,N_514);
or U1000 (N_1000,N_42,N_258);
and U1001 (N_1001,N_387,N_468);
nor U1002 (N_1002,N_254,N_2);
or U1003 (N_1003,N_248,N_232);
nand U1004 (N_1004,N_599,N_443);
nor U1005 (N_1005,N_224,N_132);
nor U1006 (N_1006,N_334,N_329);
or U1007 (N_1007,N_25,N_390);
and U1008 (N_1008,N_494,N_513);
and U1009 (N_1009,N_46,N_491);
nor U1010 (N_1010,N_533,N_489);
nand U1011 (N_1011,N_435,N_346);
nor U1012 (N_1012,N_126,N_315);
nand U1013 (N_1013,N_340,N_310);
and U1014 (N_1014,N_65,N_193);
and U1015 (N_1015,N_213,N_394);
and U1016 (N_1016,N_447,N_131);
nor U1017 (N_1017,N_370,N_123);
nor U1018 (N_1018,N_496,N_417);
or U1019 (N_1019,N_200,N_248);
nor U1020 (N_1020,N_540,N_560);
and U1021 (N_1021,N_144,N_469);
nor U1022 (N_1022,N_347,N_588);
and U1023 (N_1023,N_129,N_132);
nand U1024 (N_1024,N_47,N_199);
and U1025 (N_1025,N_211,N_404);
and U1026 (N_1026,N_186,N_309);
nand U1027 (N_1027,N_219,N_420);
or U1028 (N_1028,N_507,N_201);
nand U1029 (N_1029,N_213,N_81);
or U1030 (N_1030,N_263,N_233);
and U1031 (N_1031,N_242,N_25);
or U1032 (N_1032,N_203,N_165);
nor U1033 (N_1033,N_101,N_493);
and U1034 (N_1034,N_102,N_162);
nand U1035 (N_1035,N_593,N_211);
xor U1036 (N_1036,N_227,N_52);
nor U1037 (N_1037,N_123,N_322);
or U1038 (N_1038,N_418,N_273);
or U1039 (N_1039,N_99,N_4);
xor U1040 (N_1040,N_149,N_151);
nor U1041 (N_1041,N_230,N_191);
and U1042 (N_1042,N_18,N_69);
nor U1043 (N_1043,N_423,N_300);
nand U1044 (N_1044,N_503,N_444);
and U1045 (N_1045,N_554,N_86);
and U1046 (N_1046,N_261,N_112);
nor U1047 (N_1047,N_122,N_573);
and U1048 (N_1048,N_229,N_199);
and U1049 (N_1049,N_291,N_34);
and U1050 (N_1050,N_135,N_149);
or U1051 (N_1051,N_1,N_416);
nor U1052 (N_1052,N_419,N_280);
or U1053 (N_1053,N_217,N_216);
or U1054 (N_1054,N_318,N_376);
nor U1055 (N_1055,N_126,N_502);
or U1056 (N_1056,N_53,N_301);
or U1057 (N_1057,N_215,N_264);
nor U1058 (N_1058,N_201,N_589);
and U1059 (N_1059,N_87,N_478);
nand U1060 (N_1060,N_570,N_494);
or U1061 (N_1061,N_187,N_548);
or U1062 (N_1062,N_479,N_180);
nand U1063 (N_1063,N_295,N_482);
or U1064 (N_1064,N_9,N_467);
or U1065 (N_1065,N_392,N_493);
and U1066 (N_1066,N_510,N_28);
or U1067 (N_1067,N_220,N_223);
and U1068 (N_1068,N_434,N_566);
or U1069 (N_1069,N_51,N_419);
nor U1070 (N_1070,N_518,N_585);
nand U1071 (N_1071,N_178,N_435);
nor U1072 (N_1072,N_154,N_555);
nand U1073 (N_1073,N_268,N_385);
nand U1074 (N_1074,N_106,N_400);
nor U1075 (N_1075,N_129,N_382);
or U1076 (N_1076,N_66,N_442);
or U1077 (N_1077,N_452,N_17);
nor U1078 (N_1078,N_437,N_466);
nor U1079 (N_1079,N_472,N_499);
nand U1080 (N_1080,N_499,N_357);
nor U1081 (N_1081,N_210,N_19);
nand U1082 (N_1082,N_94,N_469);
nand U1083 (N_1083,N_23,N_147);
or U1084 (N_1084,N_230,N_364);
nand U1085 (N_1085,N_380,N_431);
nor U1086 (N_1086,N_546,N_396);
nand U1087 (N_1087,N_200,N_484);
nand U1088 (N_1088,N_192,N_485);
nor U1089 (N_1089,N_78,N_237);
and U1090 (N_1090,N_19,N_261);
or U1091 (N_1091,N_109,N_586);
nand U1092 (N_1092,N_493,N_494);
nor U1093 (N_1093,N_134,N_178);
or U1094 (N_1094,N_355,N_163);
nor U1095 (N_1095,N_386,N_523);
or U1096 (N_1096,N_492,N_321);
xnor U1097 (N_1097,N_451,N_244);
and U1098 (N_1098,N_135,N_494);
and U1099 (N_1099,N_29,N_158);
nand U1100 (N_1100,N_478,N_246);
nor U1101 (N_1101,N_33,N_554);
xnor U1102 (N_1102,N_573,N_271);
nand U1103 (N_1103,N_64,N_240);
and U1104 (N_1104,N_230,N_103);
and U1105 (N_1105,N_584,N_236);
nand U1106 (N_1106,N_517,N_563);
or U1107 (N_1107,N_324,N_250);
or U1108 (N_1108,N_488,N_35);
nor U1109 (N_1109,N_320,N_337);
nand U1110 (N_1110,N_435,N_516);
nand U1111 (N_1111,N_549,N_99);
and U1112 (N_1112,N_249,N_234);
nand U1113 (N_1113,N_40,N_306);
and U1114 (N_1114,N_535,N_192);
nor U1115 (N_1115,N_191,N_107);
nand U1116 (N_1116,N_519,N_510);
or U1117 (N_1117,N_505,N_530);
nor U1118 (N_1118,N_452,N_319);
nor U1119 (N_1119,N_357,N_587);
nand U1120 (N_1120,N_518,N_281);
nor U1121 (N_1121,N_11,N_215);
nor U1122 (N_1122,N_244,N_322);
and U1123 (N_1123,N_171,N_513);
nor U1124 (N_1124,N_214,N_147);
and U1125 (N_1125,N_386,N_261);
and U1126 (N_1126,N_341,N_197);
nand U1127 (N_1127,N_385,N_222);
and U1128 (N_1128,N_469,N_584);
xor U1129 (N_1129,N_330,N_221);
and U1130 (N_1130,N_74,N_245);
or U1131 (N_1131,N_321,N_541);
or U1132 (N_1132,N_422,N_348);
nor U1133 (N_1133,N_507,N_253);
and U1134 (N_1134,N_3,N_84);
nor U1135 (N_1135,N_327,N_236);
nand U1136 (N_1136,N_516,N_496);
nand U1137 (N_1137,N_298,N_413);
xor U1138 (N_1138,N_32,N_412);
nor U1139 (N_1139,N_178,N_49);
nor U1140 (N_1140,N_31,N_431);
xor U1141 (N_1141,N_472,N_29);
or U1142 (N_1142,N_550,N_86);
nand U1143 (N_1143,N_188,N_241);
or U1144 (N_1144,N_76,N_174);
nor U1145 (N_1145,N_341,N_559);
or U1146 (N_1146,N_346,N_439);
nand U1147 (N_1147,N_53,N_468);
nand U1148 (N_1148,N_585,N_566);
nand U1149 (N_1149,N_5,N_509);
and U1150 (N_1150,N_377,N_282);
nand U1151 (N_1151,N_118,N_171);
nand U1152 (N_1152,N_358,N_579);
nor U1153 (N_1153,N_59,N_360);
or U1154 (N_1154,N_393,N_305);
or U1155 (N_1155,N_83,N_264);
nor U1156 (N_1156,N_137,N_285);
and U1157 (N_1157,N_548,N_560);
or U1158 (N_1158,N_108,N_300);
nor U1159 (N_1159,N_396,N_572);
nor U1160 (N_1160,N_429,N_333);
nor U1161 (N_1161,N_43,N_122);
nor U1162 (N_1162,N_553,N_485);
and U1163 (N_1163,N_232,N_178);
or U1164 (N_1164,N_282,N_270);
nand U1165 (N_1165,N_510,N_220);
nand U1166 (N_1166,N_591,N_45);
and U1167 (N_1167,N_64,N_587);
nor U1168 (N_1168,N_521,N_86);
nand U1169 (N_1169,N_131,N_461);
nor U1170 (N_1170,N_403,N_411);
and U1171 (N_1171,N_420,N_87);
nand U1172 (N_1172,N_84,N_90);
nand U1173 (N_1173,N_407,N_343);
and U1174 (N_1174,N_6,N_62);
and U1175 (N_1175,N_36,N_66);
nor U1176 (N_1176,N_276,N_77);
nor U1177 (N_1177,N_35,N_36);
nand U1178 (N_1178,N_435,N_245);
and U1179 (N_1179,N_409,N_450);
nand U1180 (N_1180,N_298,N_302);
xor U1181 (N_1181,N_357,N_194);
or U1182 (N_1182,N_288,N_133);
nand U1183 (N_1183,N_572,N_116);
nor U1184 (N_1184,N_289,N_554);
nor U1185 (N_1185,N_102,N_107);
and U1186 (N_1186,N_494,N_546);
nand U1187 (N_1187,N_466,N_294);
nand U1188 (N_1188,N_242,N_355);
and U1189 (N_1189,N_4,N_74);
nand U1190 (N_1190,N_353,N_79);
nor U1191 (N_1191,N_352,N_300);
or U1192 (N_1192,N_114,N_375);
nand U1193 (N_1193,N_427,N_223);
nand U1194 (N_1194,N_279,N_333);
and U1195 (N_1195,N_302,N_141);
nor U1196 (N_1196,N_412,N_577);
nand U1197 (N_1197,N_488,N_257);
and U1198 (N_1198,N_370,N_186);
and U1199 (N_1199,N_7,N_239);
nor U1200 (N_1200,N_978,N_840);
and U1201 (N_1201,N_1099,N_1163);
and U1202 (N_1202,N_1123,N_1168);
or U1203 (N_1203,N_875,N_1166);
nor U1204 (N_1204,N_638,N_873);
nor U1205 (N_1205,N_929,N_830);
or U1206 (N_1206,N_699,N_755);
nor U1207 (N_1207,N_1136,N_603);
nor U1208 (N_1208,N_611,N_807);
or U1209 (N_1209,N_885,N_957);
nor U1210 (N_1210,N_734,N_744);
nor U1211 (N_1211,N_672,N_738);
or U1212 (N_1212,N_1010,N_720);
nand U1213 (N_1213,N_976,N_851);
nor U1214 (N_1214,N_891,N_1079);
nor U1215 (N_1215,N_844,N_1024);
nand U1216 (N_1216,N_617,N_691);
nor U1217 (N_1217,N_739,N_650);
xor U1218 (N_1218,N_1185,N_618);
nand U1219 (N_1219,N_605,N_654);
and U1220 (N_1220,N_1021,N_751);
nor U1221 (N_1221,N_1009,N_764);
nor U1222 (N_1222,N_943,N_1091);
nand U1223 (N_1223,N_810,N_1051);
nor U1224 (N_1224,N_722,N_705);
or U1225 (N_1225,N_661,N_860);
nand U1226 (N_1226,N_833,N_653);
and U1227 (N_1227,N_643,N_1146);
nand U1228 (N_1228,N_856,N_754);
nor U1229 (N_1229,N_781,N_817);
or U1230 (N_1230,N_906,N_1018);
nor U1231 (N_1231,N_736,N_786);
nor U1232 (N_1232,N_1191,N_1101);
and U1233 (N_1233,N_850,N_1031);
or U1234 (N_1234,N_766,N_780);
and U1235 (N_1235,N_793,N_1043);
or U1236 (N_1236,N_721,N_763);
nand U1237 (N_1237,N_1150,N_1134);
nor U1238 (N_1238,N_948,N_1077);
nor U1239 (N_1239,N_623,N_1037);
nand U1240 (N_1240,N_905,N_1030);
xor U1241 (N_1241,N_852,N_1190);
nand U1242 (N_1242,N_797,N_1180);
nor U1243 (N_1243,N_953,N_1175);
nand U1244 (N_1244,N_629,N_1182);
xnor U1245 (N_1245,N_637,N_1165);
nand U1246 (N_1246,N_1068,N_1036);
and U1247 (N_1247,N_811,N_973);
or U1248 (N_1248,N_995,N_1071);
or U1249 (N_1249,N_765,N_1120);
and U1250 (N_1250,N_1129,N_1049);
nand U1251 (N_1251,N_1118,N_994);
and U1252 (N_1252,N_771,N_774);
or U1253 (N_1253,N_698,N_874);
or U1254 (N_1254,N_701,N_677);
or U1255 (N_1255,N_1003,N_937);
nand U1256 (N_1256,N_748,N_879);
nand U1257 (N_1257,N_612,N_1194);
or U1258 (N_1258,N_839,N_1046);
or U1259 (N_1259,N_675,N_1032);
nor U1260 (N_1260,N_846,N_990);
and U1261 (N_1261,N_1193,N_1139);
or U1262 (N_1262,N_951,N_1104);
nor U1263 (N_1263,N_1112,N_1029);
and U1264 (N_1264,N_824,N_1074);
and U1265 (N_1265,N_655,N_950);
or U1266 (N_1266,N_858,N_750);
xnor U1267 (N_1267,N_892,N_903);
and U1268 (N_1268,N_1196,N_967);
or U1269 (N_1269,N_652,N_855);
nor U1270 (N_1270,N_831,N_1064);
nor U1271 (N_1271,N_782,N_986);
and U1272 (N_1272,N_659,N_845);
nor U1273 (N_1273,N_923,N_998);
nand U1274 (N_1274,N_620,N_883);
or U1275 (N_1275,N_1177,N_902);
nor U1276 (N_1276,N_1159,N_932);
or U1277 (N_1277,N_886,N_788);
or U1278 (N_1278,N_895,N_709);
and U1279 (N_1279,N_982,N_684);
or U1280 (N_1280,N_685,N_727);
nor U1281 (N_1281,N_640,N_801);
and U1282 (N_1282,N_627,N_1167);
and U1283 (N_1283,N_1137,N_1189);
or U1284 (N_1284,N_938,N_884);
or U1285 (N_1285,N_799,N_970);
nand U1286 (N_1286,N_899,N_1173);
nor U1287 (N_1287,N_634,N_1063);
nor U1288 (N_1288,N_835,N_1174);
and U1289 (N_1289,N_1170,N_616);
nor U1290 (N_1290,N_1039,N_822);
or U1291 (N_1291,N_1153,N_619);
nand U1292 (N_1292,N_991,N_1069);
or U1293 (N_1293,N_1103,N_604);
nand U1294 (N_1294,N_707,N_1157);
and U1295 (N_1295,N_926,N_912);
nor U1296 (N_1296,N_1087,N_1106);
nor U1297 (N_1297,N_869,N_749);
nand U1298 (N_1298,N_924,N_778);
nor U1299 (N_1299,N_1090,N_731);
nand U1300 (N_1300,N_742,N_1001);
nand U1301 (N_1301,N_683,N_815);
or U1302 (N_1302,N_714,N_1131);
or U1303 (N_1303,N_897,N_882);
or U1304 (N_1304,N_857,N_954);
or U1305 (N_1305,N_1109,N_608);
nor U1306 (N_1306,N_662,N_633);
nor U1307 (N_1307,N_706,N_665);
nor U1308 (N_1308,N_1124,N_800);
nand U1309 (N_1309,N_768,N_942);
nor U1310 (N_1310,N_1078,N_1122);
and U1311 (N_1311,N_1085,N_696);
or U1312 (N_1312,N_1130,N_1006);
and U1313 (N_1313,N_651,N_798);
and U1314 (N_1314,N_915,N_1033);
or U1315 (N_1315,N_1015,N_1056);
nor U1316 (N_1316,N_896,N_1184);
and U1317 (N_1317,N_1028,N_779);
and U1318 (N_1318,N_642,N_743);
nor U1319 (N_1319,N_796,N_1050);
nand U1320 (N_1320,N_802,N_862);
nor U1321 (N_1321,N_1192,N_1080);
nor U1322 (N_1322,N_894,N_645);
xor U1323 (N_1323,N_787,N_890);
nand U1324 (N_1324,N_1045,N_966);
and U1325 (N_1325,N_854,N_1012);
or U1326 (N_1326,N_631,N_1070);
or U1327 (N_1327,N_1156,N_1114);
nand U1328 (N_1328,N_747,N_911);
nor U1329 (N_1329,N_1172,N_909);
and U1330 (N_1330,N_772,N_1000);
or U1331 (N_1331,N_717,N_1005);
and U1332 (N_1332,N_803,N_1048);
or U1333 (N_1333,N_1143,N_745);
and U1334 (N_1334,N_1075,N_834);
or U1335 (N_1335,N_690,N_925);
xor U1336 (N_1336,N_988,N_1017);
or U1337 (N_1337,N_1144,N_961);
and U1338 (N_1338,N_726,N_1089);
and U1339 (N_1339,N_814,N_907);
or U1340 (N_1340,N_1055,N_1007);
nor U1341 (N_1341,N_992,N_1195);
nand U1342 (N_1342,N_939,N_700);
or U1343 (N_1343,N_1096,N_901);
nand U1344 (N_1344,N_1082,N_945);
nand U1345 (N_1345,N_692,N_838);
nor U1346 (N_1346,N_1086,N_681);
and U1347 (N_1347,N_1110,N_1047);
nand U1348 (N_1348,N_1038,N_1142);
and U1349 (N_1349,N_861,N_917);
or U1350 (N_1350,N_1187,N_671);
and U1351 (N_1351,N_732,N_622);
or U1352 (N_1352,N_859,N_723);
nand U1353 (N_1353,N_1040,N_872);
nand U1354 (N_1354,N_713,N_777);
and U1355 (N_1355,N_1161,N_687);
or U1356 (N_1356,N_1095,N_997);
or U1357 (N_1357,N_794,N_636);
and U1358 (N_1358,N_607,N_1088);
nor U1359 (N_1359,N_1147,N_600);
or U1360 (N_1360,N_962,N_809);
or U1361 (N_1361,N_1171,N_1119);
nand U1362 (N_1362,N_843,N_919);
nand U1363 (N_1363,N_656,N_975);
and U1364 (N_1364,N_1140,N_989);
or U1365 (N_1365,N_1061,N_1162);
nor U1366 (N_1366,N_1011,N_1081);
nand U1367 (N_1367,N_759,N_648);
or U1368 (N_1368,N_718,N_985);
xnor U1369 (N_1369,N_613,N_737);
or U1370 (N_1370,N_770,N_870);
xnor U1371 (N_1371,N_1155,N_1111);
nand U1372 (N_1372,N_783,N_876);
nand U1373 (N_1373,N_1164,N_712);
and U1374 (N_1374,N_639,N_647);
or U1375 (N_1375,N_660,N_670);
and U1376 (N_1376,N_791,N_1102);
and U1377 (N_1377,N_848,N_746);
nand U1378 (N_1378,N_711,N_646);
and U1379 (N_1379,N_947,N_868);
nand U1380 (N_1380,N_1145,N_898);
nand U1381 (N_1381,N_628,N_1135);
nand U1382 (N_1382,N_1023,N_694);
nor U1383 (N_1383,N_716,N_1148);
nor U1384 (N_1384,N_1098,N_624);
and U1385 (N_1385,N_1019,N_740);
or U1386 (N_1386,N_1188,N_1020);
and U1387 (N_1387,N_1067,N_1062);
and U1388 (N_1388,N_724,N_601);
and U1389 (N_1389,N_626,N_974);
nor U1390 (N_1390,N_849,N_941);
nand U1391 (N_1391,N_669,N_1132);
and U1392 (N_1392,N_674,N_865);
nand U1393 (N_1393,N_728,N_1169);
or U1394 (N_1394,N_1093,N_993);
or U1395 (N_1395,N_880,N_1092);
nand U1396 (N_1396,N_1141,N_940);
nor U1397 (N_1397,N_676,N_959);
nand U1398 (N_1398,N_668,N_914);
nand U1399 (N_1399,N_863,N_649);
nand U1400 (N_1400,N_877,N_969);
or U1401 (N_1401,N_821,N_635);
or U1402 (N_1402,N_1022,N_708);
and U1403 (N_1403,N_826,N_952);
and U1404 (N_1404,N_792,N_980);
and U1405 (N_1405,N_1044,N_1154);
nor U1406 (N_1406,N_1034,N_933);
nor U1407 (N_1407,N_864,N_679);
nand U1408 (N_1408,N_680,N_789);
and U1409 (N_1409,N_808,N_686);
or U1410 (N_1410,N_730,N_1083);
or U1411 (N_1411,N_1027,N_602);
and U1412 (N_1412,N_666,N_725);
nor U1413 (N_1413,N_1008,N_735);
nor U1414 (N_1414,N_644,N_1054);
nor U1415 (N_1415,N_867,N_741);
and U1416 (N_1416,N_832,N_908);
and U1417 (N_1417,N_828,N_1002);
and U1418 (N_1418,N_987,N_1108);
or U1419 (N_1419,N_812,N_968);
nand U1420 (N_1420,N_813,N_641);
nand U1421 (N_1421,N_931,N_818);
or U1422 (N_1422,N_913,N_1149);
nand U1423 (N_1423,N_1042,N_936);
nand U1424 (N_1424,N_1053,N_1097);
or U1425 (N_1425,N_804,N_965);
nand U1426 (N_1426,N_625,N_888);
nand U1427 (N_1427,N_922,N_1057);
or U1428 (N_1428,N_775,N_1183);
and U1429 (N_1429,N_693,N_1115);
and U1430 (N_1430,N_983,N_1107);
or U1431 (N_1431,N_958,N_1127);
or U1432 (N_1432,N_893,N_729);
nand U1433 (N_1433,N_984,N_1041);
nand U1434 (N_1434,N_1116,N_773);
or U1435 (N_1435,N_1158,N_752);
nor U1436 (N_1436,N_1016,N_853);
nor U1437 (N_1437,N_767,N_1004);
or U1438 (N_1438,N_1125,N_1138);
nor U1439 (N_1439,N_964,N_1121);
and U1440 (N_1440,N_769,N_1052);
and U1441 (N_1441,N_1179,N_881);
or U1442 (N_1442,N_632,N_795);
and U1443 (N_1443,N_667,N_1065);
or U1444 (N_1444,N_910,N_847);
and U1445 (N_1445,N_614,N_1105);
nor U1446 (N_1446,N_1128,N_918);
or U1447 (N_1447,N_1199,N_825);
nand U1448 (N_1448,N_928,N_920);
nand U1449 (N_1449,N_695,N_1025);
and U1450 (N_1450,N_1198,N_827);
and U1451 (N_1451,N_921,N_610);
nor U1452 (N_1452,N_971,N_760);
nand U1453 (N_1453,N_842,N_819);
nand U1454 (N_1454,N_806,N_823);
and U1455 (N_1455,N_889,N_955);
or U1456 (N_1456,N_678,N_621);
nand U1457 (N_1457,N_900,N_1084);
and U1458 (N_1458,N_606,N_790);
and U1459 (N_1459,N_972,N_1073);
or U1460 (N_1460,N_934,N_871);
or U1461 (N_1461,N_977,N_981);
nor U1462 (N_1462,N_1035,N_1066);
and U1463 (N_1463,N_837,N_663);
xor U1464 (N_1464,N_784,N_887);
and U1465 (N_1465,N_1151,N_1117);
xor U1466 (N_1466,N_1059,N_689);
or U1467 (N_1467,N_776,N_702);
nor U1468 (N_1468,N_960,N_1026);
and U1469 (N_1469,N_904,N_1072);
or U1470 (N_1470,N_1100,N_682);
nand U1471 (N_1471,N_704,N_1176);
and U1472 (N_1472,N_697,N_805);
nor U1473 (N_1473,N_673,N_820);
nand U1474 (N_1474,N_935,N_1060);
nand U1475 (N_1475,N_949,N_1186);
nand U1476 (N_1476,N_757,N_829);
or U1477 (N_1477,N_761,N_996);
and U1478 (N_1478,N_719,N_1058);
nor U1479 (N_1479,N_878,N_1181);
and U1480 (N_1480,N_979,N_836);
nand U1481 (N_1481,N_1094,N_866);
and U1482 (N_1482,N_944,N_756);
and U1483 (N_1483,N_946,N_733);
nor U1484 (N_1484,N_710,N_1014);
and U1485 (N_1485,N_1197,N_963);
and U1486 (N_1486,N_1076,N_916);
nor U1487 (N_1487,N_930,N_715);
nand U1488 (N_1488,N_1160,N_816);
or U1489 (N_1489,N_630,N_762);
nor U1490 (N_1490,N_657,N_1013);
nor U1491 (N_1491,N_664,N_999);
nand U1492 (N_1492,N_688,N_1113);
or U1493 (N_1493,N_956,N_615);
or U1494 (N_1494,N_1178,N_609);
nand U1495 (N_1495,N_753,N_927);
nor U1496 (N_1496,N_1152,N_1126);
nand U1497 (N_1497,N_658,N_841);
and U1498 (N_1498,N_785,N_703);
nor U1499 (N_1499,N_1133,N_758);
nor U1500 (N_1500,N_853,N_900);
nand U1501 (N_1501,N_648,N_841);
and U1502 (N_1502,N_940,N_1187);
xnor U1503 (N_1503,N_781,N_887);
nand U1504 (N_1504,N_974,N_929);
nand U1505 (N_1505,N_1178,N_631);
or U1506 (N_1506,N_1005,N_736);
or U1507 (N_1507,N_1187,N_809);
nor U1508 (N_1508,N_1073,N_805);
nor U1509 (N_1509,N_814,N_857);
or U1510 (N_1510,N_985,N_1137);
and U1511 (N_1511,N_1064,N_690);
and U1512 (N_1512,N_967,N_803);
nand U1513 (N_1513,N_1160,N_899);
nor U1514 (N_1514,N_1009,N_655);
or U1515 (N_1515,N_1038,N_857);
xor U1516 (N_1516,N_732,N_759);
nand U1517 (N_1517,N_720,N_1100);
nand U1518 (N_1518,N_866,N_997);
nand U1519 (N_1519,N_1112,N_1179);
and U1520 (N_1520,N_781,N_665);
or U1521 (N_1521,N_695,N_893);
or U1522 (N_1522,N_618,N_919);
nor U1523 (N_1523,N_704,N_1179);
nand U1524 (N_1524,N_1099,N_853);
or U1525 (N_1525,N_1155,N_1182);
nand U1526 (N_1526,N_763,N_649);
nor U1527 (N_1527,N_1033,N_661);
or U1528 (N_1528,N_696,N_1101);
nor U1529 (N_1529,N_742,N_641);
xor U1530 (N_1530,N_896,N_1050);
nand U1531 (N_1531,N_982,N_948);
and U1532 (N_1532,N_671,N_662);
and U1533 (N_1533,N_684,N_769);
and U1534 (N_1534,N_647,N_665);
nor U1535 (N_1535,N_684,N_778);
and U1536 (N_1536,N_964,N_617);
nand U1537 (N_1537,N_1027,N_869);
or U1538 (N_1538,N_1135,N_853);
nor U1539 (N_1539,N_925,N_622);
nand U1540 (N_1540,N_773,N_908);
nand U1541 (N_1541,N_941,N_763);
nand U1542 (N_1542,N_639,N_1019);
nand U1543 (N_1543,N_1199,N_897);
nand U1544 (N_1544,N_626,N_1004);
nand U1545 (N_1545,N_1053,N_870);
nand U1546 (N_1546,N_806,N_680);
nand U1547 (N_1547,N_1076,N_884);
nand U1548 (N_1548,N_690,N_767);
nand U1549 (N_1549,N_1122,N_830);
or U1550 (N_1550,N_657,N_1050);
and U1551 (N_1551,N_1151,N_817);
or U1552 (N_1552,N_810,N_737);
nor U1553 (N_1553,N_665,N_605);
and U1554 (N_1554,N_885,N_1165);
nor U1555 (N_1555,N_727,N_983);
nand U1556 (N_1556,N_740,N_953);
nor U1557 (N_1557,N_1004,N_685);
or U1558 (N_1558,N_977,N_620);
nor U1559 (N_1559,N_737,N_720);
and U1560 (N_1560,N_689,N_821);
nand U1561 (N_1561,N_807,N_961);
nor U1562 (N_1562,N_1102,N_1123);
or U1563 (N_1563,N_785,N_684);
or U1564 (N_1564,N_654,N_1105);
nor U1565 (N_1565,N_1199,N_1008);
or U1566 (N_1566,N_707,N_1043);
nor U1567 (N_1567,N_1102,N_755);
nand U1568 (N_1568,N_955,N_865);
nand U1569 (N_1569,N_901,N_681);
or U1570 (N_1570,N_910,N_684);
or U1571 (N_1571,N_1131,N_1180);
and U1572 (N_1572,N_1114,N_848);
and U1573 (N_1573,N_1122,N_937);
or U1574 (N_1574,N_661,N_734);
or U1575 (N_1575,N_663,N_1166);
nor U1576 (N_1576,N_970,N_699);
nor U1577 (N_1577,N_1103,N_1157);
or U1578 (N_1578,N_870,N_886);
and U1579 (N_1579,N_1101,N_863);
or U1580 (N_1580,N_615,N_1155);
nand U1581 (N_1581,N_848,N_606);
and U1582 (N_1582,N_895,N_1023);
nor U1583 (N_1583,N_652,N_1187);
or U1584 (N_1584,N_616,N_622);
nor U1585 (N_1585,N_739,N_790);
and U1586 (N_1586,N_972,N_880);
or U1587 (N_1587,N_627,N_767);
nand U1588 (N_1588,N_646,N_877);
or U1589 (N_1589,N_876,N_1078);
nand U1590 (N_1590,N_603,N_798);
nor U1591 (N_1591,N_1027,N_1126);
nor U1592 (N_1592,N_1169,N_1033);
or U1593 (N_1593,N_781,N_1049);
nand U1594 (N_1594,N_890,N_1070);
and U1595 (N_1595,N_816,N_640);
or U1596 (N_1596,N_835,N_840);
and U1597 (N_1597,N_853,N_1164);
and U1598 (N_1598,N_720,N_653);
and U1599 (N_1599,N_1081,N_650);
nand U1600 (N_1600,N_917,N_850);
and U1601 (N_1601,N_728,N_838);
nand U1602 (N_1602,N_1081,N_607);
and U1603 (N_1603,N_1164,N_1011);
and U1604 (N_1604,N_808,N_946);
nor U1605 (N_1605,N_1112,N_813);
or U1606 (N_1606,N_1167,N_635);
nand U1607 (N_1607,N_1025,N_834);
xnor U1608 (N_1608,N_934,N_692);
and U1609 (N_1609,N_1038,N_1195);
nand U1610 (N_1610,N_853,N_1123);
nor U1611 (N_1611,N_1124,N_1136);
nor U1612 (N_1612,N_941,N_613);
nand U1613 (N_1613,N_912,N_947);
or U1614 (N_1614,N_701,N_670);
or U1615 (N_1615,N_1067,N_1116);
nand U1616 (N_1616,N_1144,N_1160);
nor U1617 (N_1617,N_907,N_726);
nand U1618 (N_1618,N_1198,N_916);
nand U1619 (N_1619,N_673,N_1106);
nor U1620 (N_1620,N_862,N_666);
nor U1621 (N_1621,N_1004,N_633);
or U1622 (N_1622,N_1075,N_1115);
or U1623 (N_1623,N_822,N_1186);
and U1624 (N_1624,N_1120,N_1037);
or U1625 (N_1625,N_800,N_821);
nand U1626 (N_1626,N_920,N_619);
nand U1627 (N_1627,N_861,N_703);
nand U1628 (N_1628,N_821,N_666);
nand U1629 (N_1629,N_1145,N_924);
and U1630 (N_1630,N_945,N_1167);
nor U1631 (N_1631,N_752,N_921);
xor U1632 (N_1632,N_929,N_1111);
nand U1633 (N_1633,N_735,N_1066);
nand U1634 (N_1634,N_778,N_1169);
nor U1635 (N_1635,N_702,N_762);
nand U1636 (N_1636,N_639,N_625);
or U1637 (N_1637,N_729,N_971);
or U1638 (N_1638,N_1093,N_1005);
or U1639 (N_1639,N_839,N_955);
and U1640 (N_1640,N_758,N_1019);
or U1641 (N_1641,N_1161,N_1123);
nand U1642 (N_1642,N_666,N_962);
nor U1643 (N_1643,N_918,N_1064);
nand U1644 (N_1644,N_660,N_1039);
nand U1645 (N_1645,N_624,N_1043);
nand U1646 (N_1646,N_748,N_1084);
and U1647 (N_1647,N_648,N_1172);
nor U1648 (N_1648,N_842,N_809);
or U1649 (N_1649,N_1095,N_993);
or U1650 (N_1650,N_780,N_671);
nor U1651 (N_1651,N_803,N_808);
and U1652 (N_1652,N_1167,N_1033);
and U1653 (N_1653,N_794,N_960);
or U1654 (N_1654,N_643,N_1064);
nand U1655 (N_1655,N_651,N_1067);
nand U1656 (N_1656,N_1087,N_1136);
and U1657 (N_1657,N_894,N_839);
and U1658 (N_1658,N_737,N_601);
or U1659 (N_1659,N_868,N_760);
nand U1660 (N_1660,N_892,N_829);
nor U1661 (N_1661,N_1163,N_613);
nand U1662 (N_1662,N_809,N_648);
and U1663 (N_1663,N_882,N_866);
and U1664 (N_1664,N_1024,N_899);
nor U1665 (N_1665,N_966,N_836);
and U1666 (N_1666,N_634,N_859);
and U1667 (N_1667,N_947,N_1029);
and U1668 (N_1668,N_999,N_1092);
nand U1669 (N_1669,N_685,N_839);
nor U1670 (N_1670,N_919,N_684);
nor U1671 (N_1671,N_915,N_685);
or U1672 (N_1672,N_994,N_1012);
or U1673 (N_1673,N_1138,N_1096);
nor U1674 (N_1674,N_672,N_1128);
and U1675 (N_1675,N_870,N_1015);
and U1676 (N_1676,N_1028,N_644);
and U1677 (N_1677,N_896,N_640);
or U1678 (N_1678,N_1007,N_613);
nand U1679 (N_1679,N_869,N_1198);
and U1680 (N_1680,N_1017,N_921);
or U1681 (N_1681,N_786,N_768);
nor U1682 (N_1682,N_600,N_753);
or U1683 (N_1683,N_842,N_869);
nor U1684 (N_1684,N_636,N_773);
xnor U1685 (N_1685,N_1027,N_913);
xor U1686 (N_1686,N_959,N_1150);
or U1687 (N_1687,N_766,N_672);
nor U1688 (N_1688,N_626,N_1016);
nand U1689 (N_1689,N_901,N_649);
or U1690 (N_1690,N_933,N_675);
nor U1691 (N_1691,N_943,N_1058);
nor U1692 (N_1692,N_928,N_656);
nand U1693 (N_1693,N_1199,N_991);
and U1694 (N_1694,N_641,N_983);
nand U1695 (N_1695,N_748,N_856);
nor U1696 (N_1696,N_1082,N_1018);
xnor U1697 (N_1697,N_1038,N_687);
or U1698 (N_1698,N_837,N_995);
or U1699 (N_1699,N_1144,N_912);
or U1700 (N_1700,N_758,N_1149);
nand U1701 (N_1701,N_1061,N_1169);
or U1702 (N_1702,N_674,N_1178);
nor U1703 (N_1703,N_726,N_1160);
and U1704 (N_1704,N_838,N_1075);
or U1705 (N_1705,N_954,N_1041);
or U1706 (N_1706,N_1120,N_646);
and U1707 (N_1707,N_865,N_1063);
and U1708 (N_1708,N_1081,N_772);
nand U1709 (N_1709,N_819,N_1121);
and U1710 (N_1710,N_952,N_872);
or U1711 (N_1711,N_1140,N_624);
and U1712 (N_1712,N_815,N_973);
or U1713 (N_1713,N_765,N_808);
or U1714 (N_1714,N_618,N_1165);
or U1715 (N_1715,N_705,N_1004);
and U1716 (N_1716,N_952,N_791);
or U1717 (N_1717,N_729,N_1181);
nor U1718 (N_1718,N_880,N_1042);
or U1719 (N_1719,N_1148,N_1101);
or U1720 (N_1720,N_693,N_909);
or U1721 (N_1721,N_1115,N_644);
nor U1722 (N_1722,N_1156,N_950);
or U1723 (N_1723,N_815,N_1022);
and U1724 (N_1724,N_738,N_602);
xnor U1725 (N_1725,N_863,N_693);
or U1726 (N_1726,N_1090,N_1035);
and U1727 (N_1727,N_1002,N_1127);
nand U1728 (N_1728,N_743,N_1188);
nand U1729 (N_1729,N_814,N_675);
nor U1730 (N_1730,N_671,N_921);
xor U1731 (N_1731,N_1186,N_768);
nand U1732 (N_1732,N_686,N_847);
or U1733 (N_1733,N_896,N_619);
nor U1734 (N_1734,N_937,N_1080);
or U1735 (N_1735,N_780,N_687);
and U1736 (N_1736,N_782,N_605);
nand U1737 (N_1737,N_816,N_1187);
or U1738 (N_1738,N_1148,N_880);
nor U1739 (N_1739,N_908,N_729);
and U1740 (N_1740,N_709,N_638);
nand U1741 (N_1741,N_891,N_675);
nand U1742 (N_1742,N_1198,N_645);
nand U1743 (N_1743,N_740,N_1198);
nand U1744 (N_1744,N_699,N_1175);
xor U1745 (N_1745,N_1152,N_686);
xor U1746 (N_1746,N_964,N_781);
nand U1747 (N_1747,N_763,N_1152);
or U1748 (N_1748,N_792,N_1043);
and U1749 (N_1749,N_922,N_1180);
nor U1750 (N_1750,N_613,N_772);
nand U1751 (N_1751,N_923,N_684);
nand U1752 (N_1752,N_909,N_783);
or U1753 (N_1753,N_607,N_674);
nor U1754 (N_1754,N_851,N_810);
or U1755 (N_1755,N_1159,N_946);
and U1756 (N_1756,N_682,N_713);
nand U1757 (N_1757,N_1150,N_972);
or U1758 (N_1758,N_645,N_774);
nor U1759 (N_1759,N_694,N_1109);
nor U1760 (N_1760,N_853,N_759);
and U1761 (N_1761,N_830,N_978);
and U1762 (N_1762,N_1070,N_1087);
and U1763 (N_1763,N_1072,N_625);
nor U1764 (N_1764,N_848,N_709);
nand U1765 (N_1765,N_1074,N_931);
or U1766 (N_1766,N_1150,N_617);
nor U1767 (N_1767,N_1183,N_1021);
and U1768 (N_1768,N_686,N_886);
or U1769 (N_1769,N_986,N_1195);
nand U1770 (N_1770,N_801,N_858);
or U1771 (N_1771,N_727,N_1082);
and U1772 (N_1772,N_758,N_1060);
and U1773 (N_1773,N_1174,N_1045);
nand U1774 (N_1774,N_638,N_734);
or U1775 (N_1775,N_1084,N_731);
nand U1776 (N_1776,N_665,N_989);
nand U1777 (N_1777,N_1003,N_726);
or U1778 (N_1778,N_891,N_1138);
or U1779 (N_1779,N_1027,N_1022);
nand U1780 (N_1780,N_800,N_927);
or U1781 (N_1781,N_983,N_1098);
nor U1782 (N_1782,N_773,N_771);
nor U1783 (N_1783,N_659,N_677);
nor U1784 (N_1784,N_752,N_814);
or U1785 (N_1785,N_1076,N_769);
and U1786 (N_1786,N_612,N_691);
or U1787 (N_1787,N_771,N_1140);
nor U1788 (N_1788,N_819,N_690);
and U1789 (N_1789,N_1147,N_720);
or U1790 (N_1790,N_1197,N_1082);
or U1791 (N_1791,N_1136,N_884);
nor U1792 (N_1792,N_958,N_832);
nand U1793 (N_1793,N_1162,N_991);
or U1794 (N_1794,N_651,N_864);
nand U1795 (N_1795,N_893,N_1065);
nand U1796 (N_1796,N_979,N_864);
or U1797 (N_1797,N_1119,N_676);
and U1798 (N_1798,N_950,N_1008);
nand U1799 (N_1799,N_1129,N_926);
nand U1800 (N_1800,N_1579,N_1642);
nor U1801 (N_1801,N_1666,N_1210);
nand U1802 (N_1802,N_1396,N_1526);
or U1803 (N_1803,N_1541,N_1301);
nand U1804 (N_1804,N_1467,N_1319);
nor U1805 (N_1805,N_1281,N_1653);
nor U1806 (N_1806,N_1392,N_1787);
nand U1807 (N_1807,N_1625,N_1223);
and U1808 (N_1808,N_1659,N_1326);
and U1809 (N_1809,N_1631,N_1593);
or U1810 (N_1810,N_1643,N_1456);
nand U1811 (N_1811,N_1548,N_1349);
nor U1812 (N_1812,N_1338,N_1604);
nand U1813 (N_1813,N_1283,N_1294);
nand U1814 (N_1814,N_1328,N_1245);
nor U1815 (N_1815,N_1644,N_1201);
nand U1816 (N_1816,N_1617,N_1655);
nand U1817 (N_1817,N_1410,N_1718);
nor U1818 (N_1818,N_1404,N_1499);
and U1819 (N_1819,N_1699,N_1424);
or U1820 (N_1820,N_1475,N_1364);
nand U1821 (N_1821,N_1569,N_1209);
or U1822 (N_1822,N_1566,N_1514);
or U1823 (N_1823,N_1639,N_1448);
and U1824 (N_1824,N_1553,N_1204);
or U1825 (N_1825,N_1583,N_1276);
and U1826 (N_1826,N_1490,N_1397);
and U1827 (N_1827,N_1473,N_1563);
nand U1828 (N_1828,N_1369,N_1314);
nor U1829 (N_1829,N_1251,N_1411);
nor U1830 (N_1830,N_1446,N_1612);
and U1831 (N_1831,N_1280,N_1670);
or U1832 (N_1832,N_1698,N_1632);
nand U1833 (N_1833,N_1669,N_1752);
nand U1834 (N_1834,N_1431,N_1322);
nor U1835 (N_1835,N_1623,N_1320);
nand U1836 (N_1836,N_1444,N_1596);
nand U1837 (N_1837,N_1324,N_1292);
nand U1838 (N_1838,N_1504,N_1359);
nand U1839 (N_1839,N_1736,N_1496);
or U1840 (N_1840,N_1620,N_1224);
and U1841 (N_1841,N_1724,N_1225);
nor U1842 (N_1842,N_1489,N_1272);
nand U1843 (N_1843,N_1524,N_1518);
nand U1844 (N_1844,N_1562,N_1516);
or U1845 (N_1845,N_1494,N_1325);
nor U1846 (N_1846,N_1551,N_1678);
nor U1847 (N_1847,N_1383,N_1460);
nor U1848 (N_1848,N_1700,N_1437);
and U1849 (N_1849,N_1394,N_1616);
and U1850 (N_1850,N_1211,N_1454);
or U1851 (N_1851,N_1542,N_1556);
nand U1852 (N_1852,N_1771,N_1650);
nand U1853 (N_1853,N_1505,N_1408);
or U1854 (N_1854,N_1414,N_1474);
or U1855 (N_1855,N_1277,N_1498);
or U1856 (N_1856,N_1375,N_1315);
nor U1857 (N_1857,N_1795,N_1756);
nor U1858 (N_1858,N_1762,N_1218);
nand U1859 (N_1859,N_1775,N_1480);
or U1860 (N_1860,N_1264,N_1606);
or U1861 (N_1861,N_1417,N_1634);
nand U1862 (N_1862,N_1766,N_1400);
nor U1863 (N_1863,N_1343,N_1213);
nor U1864 (N_1864,N_1235,N_1413);
or U1865 (N_1865,N_1288,N_1492);
nor U1866 (N_1866,N_1366,N_1399);
xor U1867 (N_1867,N_1451,N_1258);
nor U1868 (N_1868,N_1614,N_1523);
nor U1869 (N_1869,N_1660,N_1450);
or U1870 (N_1870,N_1261,N_1714);
nand U1871 (N_1871,N_1351,N_1733);
and U1872 (N_1872,N_1726,N_1682);
nand U1873 (N_1873,N_1618,N_1545);
nor U1874 (N_1874,N_1722,N_1356);
or U1875 (N_1875,N_1689,N_1592);
and U1876 (N_1876,N_1217,N_1290);
and U1877 (N_1877,N_1384,N_1743);
nor U1878 (N_1878,N_1247,N_1742);
nand U1879 (N_1879,N_1554,N_1668);
or U1880 (N_1880,N_1308,N_1687);
or U1881 (N_1881,N_1254,N_1515);
or U1882 (N_1882,N_1433,N_1633);
nor U1883 (N_1883,N_1778,N_1701);
nand U1884 (N_1884,N_1575,N_1244);
nor U1885 (N_1885,N_1785,N_1528);
and U1886 (N_1886,N_1485,N_1436);
nand U1887 (N_1887,N_1200,N_1257);
or U1888 (N_1888,N_1458,N_1798);
and U1889 (N_1889,N_1744,N_1590);
nand U1890 (N_1890,N_1723,N_1468);
and U1891 (N_1891,N_1688,N_1794);
and U1892 (N_1892,N_1381,N_1768);
nor U1893 (N_1893,N_1405,N_1443);
and U1894 (N_1894,N_1656,N_1438);
nor U1895 (N_1895,N_1776,N_1728);
nor U1896 (N_1896,N_1521,N_1497);
and U1897 (N_1897,N_1206,N_1622);
xnor U1898 (N_1898,N_1341,N_1420);
or U1899 (N_1899,N_1564,N_1463);
nand U1900 (N_1900,N_1764,N_1725);
nand U1901 (N_1901,N_1663,N_1522);
nor U1902 (N_1902,N_1313,N_1234);
nor U1903 (N_1903,N_1285,N_1309);
or U1904 (N_1904,N_1537,N_1299);
xnor U1905 (N_1905,N_1560,N_1574);
nor U1906 (N_1906,N_1289,N_1621);
and U1907 (N_1907,N_1789,N_1423);
and U1908 (N_1908,N_1214,N_1333);
and U1909 (N_1909,N_1565,N_1535);
nand U1910 (N_1910,N_1750,N_1585);
nand U1911 (N_1911,N_1403,N_1401);
or U1912 (N_1912,N_1748,N_1291);
nand U1913 (N_1913,N_1259,N_1207);
and U1914 (N_1914,N_1388,N_1402);
nand U1915 (N_1915,N_1237,N_1638);
nand U1916 (N_1916,N_1486,N_1274);
xnor U1917 (N_1917,N_1550,N_1751);
nor U1918 (N_1918,N_1737,N_1712);
nand U1919 (N_1919,N_1339,N_1538);
nor U1920 (N_1920,N_1664,N_1662);
nor U1921 (N_1921,N_1377,N_1243);
or U1922 (N_1922,N_1788,N_1477);
or U1923 (N_1923,N_1434,N_1393);
nor U1924 (N_1924,N_1602,N_1484);
nor U1925 (N_1925,N_1284,N_1520);
nand U1926 (N_1926,N_1597,N_1746);
nand U1927 (N_1927,N_1478,N_1376);
nand U1928 (N_1928,N_1303,N_1628);
nand U1929 (N_1929,N_1559,N_1529);
xnor U1930 (N_1930,N_1435,N_1601);
or U1931 (N_1931,N_1525,N_1672);
nor U1932 (N_1932,N_1461,N_1357);
nand U1933 (N_1933,N_1763,N_1767);
nor U1934 (N_1934,N_1555,N_1530);
and U1935 (N_1935,N_1426,N_1304);
or U1936 (N_1936,N_1674,N_1365);
nand U1937 (N_1937,N_1705,N_1491);
nand U1938 (N_1938,N_1233,N_1387);
or U1939 (N_1939,N_1270,N_1342);
and U1940 (N_1940,N_1256,N_1398);
nor U1941 (N_1941,N_1587,N_1594);
nand U1942 (N_1942,N_1250,N_1588);
or U1943 (N_1943,N_1671,N_1418);
or U1944 (N_1944,N_1730,N_1268);
nand U1945 (N_1945,N_1310,N_1327);
xor U1946 (N_1946,N_1265,N_1360);
and U1947 (N_1947,N_1226,N_1368);
nor U1948 (N_1948,N_1769,N_1603);
nor U1949 (N_1949,N_1717,N_1513);
or U1950 (N_1950,N_1350,N_1488);
or U1951 (N_1951,N_1797,N_1536);
nor U1952 (N_1952,N_1716,N_1335);
and U1953 (N_1953,N_1249,N_1510);
nand U1954 (N_1954,N_1307,N_1262);
or U1955 (N_1955,N_1558,N_1472);
nor U1956 (N_1956,N_1389,N_1747);
nor U1957 (N_1957,N_1598,N_1727);
nand U1958 (N_1958,N_1758,N_1729);
nor U1959 (N_1959,N_1607,N_1577);
nor U1960 (N_1960,N_1487,N_1658);
or U1961 (N_1961,N_1665,N_1739);
and U1962 (N_1962,N_1425,N_1745);
xnor U1963 (N_1963,N_1362,N_1212);
and U1964 (N_1964,N_1275,N_1786);
nor U1965 (N_1965,N_1373,N_1509);
or U1966 (N_1966,N_1511,N_1791);
nand U1967 (N_1967,N_1306,N_1221);
and U1968 (N_1968,N_1352,N_1493);
or U1969 (N_1969,N_1567,N_1321);
or U1970 (N_1970,N_1452,N_1367);
and U1971 (N_1971,N_1605,N_1297);
and U1972 (N_1972,N_1267,N_1546);
and U1973 (N_1973,N_1316,N_1232);
nand U1974 (N_1974,N_1738,N_1260);
xor U1975 (N_1975,N_1449,N_1580);
or U1976 (N_1976,N_1427,N_1346);
nand U1977 (N_1977,N_1282,N_1675);
nor U1978 (N_1978,N_1629,N_1557);
or U1979 (N_1979,N_1749,N_1455);
or U1980 (N_1980,N_1442,N_1441);
and U1981 (N_1981,N_1228,N_1599);
nor U1982 (N_1982,N_1203,N_1709);
and U1983 (N_1983,N_1345,N_1385);
nand U1984 (N_1984,N_1371,N_1708);
nand U1985 (N_1985,N_1332,N_1540);
nor U1986 (N_1986,N_1240,N_1483);
and U1987 (N_1987,N_1252,N_1386);
or U1988 (N_1988,N_1777,N_1613);
nor U1989 (N_1989,N_1532,N_1390);
and U1990 (N_1990,N_1595,N_1457);
or U1991 (N_1991,N_1312,N_1430);
and U1992 (N_1992,N_1576,N_1784);
or U1993 (N_1993,N_1344,N_1755);
nor U1994 (N_1994,N_1759,N_1573);
nand U1995 (N_1995,N_1323,N_1246);
and U1996 (N_1996,N_1765,N_1692);
and U1997 (N_1997,N_1287,N_1783);
nand U1998 (N_1998,N_1683,N_1429);
nor U1999 (N_1999,N_1462,N_1732);
or U2000 (N_2000,N_1770,N_1761);
nand U2001 (N_2001,N_1412,N_1760);
or U2002 (N_2002,N_1652,N_1624);
nor U2003 (N_2003,N_1549,N_1253);
nor U2004 (N_2004,N_1501,N_1229);
nor U2005 (N_2005,N_1647,N_1544);
and U2006 (N_2006,N_1465,N_1502);
or U2007 (N_2007,N_1453,N_1547);
nor U2008 (N_2008,N_1799,N_1735);
or U2009 (N_2009,N_1507,N_1703);
or U2010 (N_2010,N_1481,N_1506);
nor U2011 (N_2011,N_1208,N_1395);
and U2012 (N_2012,N_1239,N_1619);
and U2013 (N_2013,N_1715,N_1329);
nand U2014 (N_2014,N_1415,N_1334);
and U2015 (N_2015,N_1657,N_1584);
nand U2016 (N_2016,N_1610,N_1406);
or U2017 (N_2017,N_1230,N_1231);
nor U2018 (N_2018,N_1279,N_1361);
and U2019 (N_2019,N_1503,N_1222);
nand U2020 (N_2020,N_1711,N_1531);
nand U2021 (N_2021,N_1470,N_1358);
or U2022 (N_2022,N_1654,N_1236);
and U2023 (N_2023,N_1796,N_1591);
nor U2024 (N_2024,N_1479,N_1741);
nand U2025 (N_2025,N_1640,N_1635);
nor U2026 (N_2026,N_1295,N_1227);
nor U2027 (N_2027,N_1719,N_1754);
nor U2028 (N_2028,N_1681,N_1278);
and U2029 (N_2029,N_1609,N_1611);
nand U2030 (N_2030,N_1482,N_1680);
nand U2031 (N_2031,N_1407,N_1469);
or U2032 (N_2032,N_1720,N_1685);
or U2033 (N_2033,N_1673,N_1263);
or U2034 (N_2034,N_1561,N_1517);
and U2035 (N_2035,N_1271,N_1238);
and U2036 (N_2036,N_1779,N_1615);
nor U2037 (N_2037,N_1363,N_1582);
nand U2038 (N_2038,N_1331,N_1773);
nand U2039 (N_2039,N_1500,N_1348);
or U2040 (N_2040,N_1215,N_1792);
nand U2041 (N_2041,N_1706,N_1641);
nand U2042 (N_2042,N_1704,N_1677);
nand U2043 (N_2043,N_1645,N_1242);
and U2044 (N_2044,N_1464,N_1428);
nor U2045 (N_2045,N_1353,N_1534);
nor U2046 (N_2046,N_1637,N_1790);
nor U2047 (N_2047,N_1370,N_1757);
and U2048 (N_2048,N_1539,N_1684);
xnor U2049 (N_2049,N_1676,N_1317);
and U2050 (N_2050,N_1495,N_1439);
nand U2051 (N_2051,N_1330,N_1432);
nor U2052 (N_2052,N_1409,N_1533);
nor U2053 (N_2053,N_1379,N_1691);
nand U2054 (N_2054,N_1568,N_1382);
nor U2055 (N_2055,N_1459,N_1422);
and U2056 (N_2056,N_1627,N_1300);
nor U2057 (N_2057,N_1661,N_1571);
and U2058 (N_2058,N_1445,N_1793);
xnor U2059 (N_2059,N_1311,N_1440);
nand U2060 (N_2060,N_1552,N_1608);
nor U2061 (N_2061,N_1416,N_1581);
or U2062 (N_2062,N_1219,N_1305);
nand U2063 (N_2063,N_1630,N_1697);
and U2064 (N_2064,N_1731,N_1651);
or U2065 (N_2065,N_1202,N_1296);
nand U2066 (N_2066,N_1636,N_1216);
and U2067 (N_2067,N_1293,N_1298);
or U2068 (N_2068,N_1780,N_1695);
nor U2069 (N_2069,N_1667,N_1721);
nor U2070 (N_2070,N_1679,N_1266);
nand U2071 (N_2071,N_1527,N_1543);
nor U2072 (N_2072,N_1421,N_1374);
nor U2073 (N_2073,N_1707,N_1419);
nand U2074 (N_2074,N_1476,N_1391);
nor U2075 (N_2075,N_1740,N_1466);
and U2076 (N_2076,N_1578,N_1626);
nor U2077 (N_2077,N_1693,N_1372);
nor U2078 (N_2078,N_1508,N_1248);
nor U2079 (N_2079,N_1220,N_1471);
nor U2080 (N_2080,N_1241,N_1586);
and U2081 (N_2081,N_1646,N_1686);
and U2082 (N_2082,N_1355,N_1649);
nor U2083 (N_2083,N_1302,N_1318);
nand U2084 (N_2084,N_1753,N_1690);
nand U2085 (N_2085,N_1600,N_1512);
nand U2086 (N_2086,N_1378,N_1347);
and U2087 (N_2087,N_1589,N_1380);
nand U2088 (N_2088,N_1774,N_1648);
nor U2089 (N_2089,N_1696,N_1286);
and U2090 (N_2090,N_1710,N_1713);
nand U2091 (N_2091,N_1772,N_1782);
nor U2092 (N_2092,N_1337,N_1694);
or U2093 (N_2093,N_1205,N_1570);
and U2094 (N_2094,N_1255,N_1734);
and U2095 (N_2095,N_1519,N_1336);
and U2096 (N_2096,N_1447,N_1572);
nor U2097 (N_2097,N_1340,N_1354);
and U2098 (N_2098,N_1702,N_1781);
and U2099 (N_2099,N_1269,N_1273);
nand U2100 (N_2100,N_1443,N_1577);
nor U2101 (N_2101,N_1527,N_1695);
nand U2102 (N_2102,N_1273,N_1221);
nor U2103 (N_2103,N_1444,N_1356);
xor U2104 (N_2104,N_1533,N_1711);
nor U2105 (N_2105,N_1738,N_1259);
and U2106 (N_2106,N_1488,N_1787);
or U2107 (N_2107,N_1353,N_1729);
or U2108 (N_2108,N_1787,N_1478);
nand U2109 (N_2109,N_1243,N_1276);
and U2110 (N_2110,N_1266,N_1484);
and U2111 (N_2111,N_1476,N_1725);
and U2112 (N_2112,N_1785,N_1555);
nand U2113 (N_2113,N_1230,N_1579);
nor U2114 (N_2114,N_1420,N_1755);
nand U2115 (N_2115,N_1436,N_1669);
nand U2116 (N_2116,N_1522,N_1397);
nor U2117 (N_2117,N_1296,N_1653);
and U2118 (N_2118,N_1752,N_1535);
nor U2119 (N_2119,N_1356,N_1323);
or U2120 (N_2120,N_1464,N_1621);
nand U2121 (N_2121,N_1333,N_1607);
and U2122 (N_2122,N_1636,N_1253);
nand U2123 (N_2123,N_1558,N_1276);
nand U2124 (N_2124,N_1318,N_1650);
xnor U2125 (N_2125,N_1720,N_1749);
nor U2126 (N_2126,N_1201,N_1396);
or U2127 (N_2127,N_1510,N_1417);
and U2128 (N_2128,N_1304,N_1274);
and U2129 (N_2129,N_1604,N_1537);
nor U2130 (N_2130,N_1709,N_1359);
nor U2131 (N_2131,N_1749,N_1625);
nand U2132 (N_2132,N_1415,N_1563);
nand U2133 (N_2133,N_1229,N_1226);
nor U2134 (N_2134,N_1683,N_1341);
nand U2135 (N_2135,N_1498,N_1436);
or U2136 (N_2136,N_1713,N_1592);
nor U2137 (N_2137,N_1321,N_1295);
or U2138 (N_2138,N_1605,N_1390);
nor U2139 (N_2139,N_1518,N_1410);
and U2140 (N_2140,N_1335,N_1351);
nand U2141 (N_2141,N_1372,N_1496);
nand U2142 (N_2142,N_1789,N_1626);
nor U2143 (N_2143,N_1282,N_1217);
xor U2144 (N_2144,N_1443,N_1351);
or U2145 (N_2145,N_1451,N_1261);
and U2146 (N_2146,N_1425,N_1771);
and U2147 (N_2147,N_1250,N_1317);
xor U2148 (N_2148,N_1482,N_1536);
or U2149 (N_2149,N_1440,N_1208);
and U2150 (N_2150,N_1502,N_1376);
nor U2151 (N_2151,N_1717,N_1712);
nand U2152 (N_2152,N_1351,N_1209);
and U2153 (N_2153,N_1274,N_1707);
or U2154 (N_2154,N_1591,N_1773);
xnor U2155 (N_2155,N_1656,N_1205);
or U2156 (N_2156,N_1475,N_1455);
nor U2157 (N_2157,N_1710,N_1530);
nor U2158 (N_2158,N_1533,N_1527);
and U2159 (N_2159,N_1634,N_1420);
or U2160 (N_2160,N_1539,N_1285);
or U2161 (N_2161,N_1337,N_1218);
nor U2162 (N_2162,N_1398,N_1267);
and U2163 (N_2163,N_1761,N_1576);
nor U2164 (N_2164,N_1798,N_1226);
nor U2165 (N_2165,N_1692,N_1444);
nand U2166 (N_2166,N_1322,N_1432);
and U2167 (N_2167,N_1463,N_1524);
nand U2168 (N_2168,N_1439,N_1335);
nor U2169 (N_2169,N_1371,N_1277);
nor U2170 (N_2170,N_1380,N_1244);
nor U2171 (N_2171,N_1385,N_1418);
and U2172 (N_2172,N_1325,N_1393);
or U2173 (N_2173,N_1347,N_1240);
or U2174 (N_2174,N_1598,N_1647);
nor U2175 (N_2175,N_1380,N_1781);
or U2176 (N_2176,N_1298,N_1241);
or U2177 (N_2177,N_1717,N_1215);
and U2178 (N_2178,N_1400,N_1735);
nor U2179 (N_2179,N_1404,N_1439);
and U2180 (N_2180,N_1747,N_1723);
or U2181 (N_2181,N_1516,N_1764);
nor U2182 (N_2182,N_1648,N_1591);
nand U2183 (N_2183,N_1369,N_1786);
nand U2184 (N_2184,N_1682,N_1286);
and U2185 (N_2185,N_1335,N_1223);
nand U2186 (N_2186,N_1514,N_1249);
or U2187 (N_2187,N_1320,N_1285);
nor U2188 (N_2188,N_1572,N_1732);
and U2189 (N_2189,N_1513,N_1451);
or U2190 (N_2190,N_1475,N_1535);
or U2191 (N_2191,N_1550,N_1319);
nand U2192 (N_2192,N_1291,N_1318);
and U2193 (N_2193,N_1618,N_1782);
and U2194 (N_2194,N_1481,N_1708);
and U2195 (N_2195,N_1254,N_1267);
nor U2196 (N_2196,N_1797,N_1216);
xnor U2197 (N_2197,N_1363,N_1612);
nand U2198 (N_2198,N_1466,N_1249);
and U2199 (N_2199,N_1601,N_1304);
or U2200 (N_2200,N_1554,N_1235);
or U2201 (N_2201,N_1760,N_1426);
nor U2202 (N_2202,N_1704,N_1523);
nand U2203 (N_2203,N_1387,N_1243);
nand U2204 (N_2204,N_1672,N_1479);
or U2205 (N_2205,N_1300,N_1455);
or U2206 (N_2206,N_1264,N_1238);
or U2207 (N_2207,N_1677,N_1758);
and U2208 (N_2208,N_1211,N_1312);
or U2209 (N_2209,N_1644,N_1458);
and U2210 (N_2210,N_1367,N_1469);
or U2211 (N_2211,N_1220,N_1592);
xnor U2212 (N_2212,N_1427,N_1552);
or U2213 (N_2213,N_1267,N_1462);
nor U2214 (N_2214,N_1618,N_1631);
and U2215 (N_2215,N_1687,N_1761);
nand U2216 (N_2216,N_1428,N_1243);
and U2217 (N_2217,N_1709,N_1396);
nor U2218 (N_2218,N_1744,N_1455);
and U2219 (N_2219,N_1767,N_1467);
and U2220 (N_2220,N_1245,N_1574);
nor U2221 (N_2221,N_1455,N_1684);
nand U2222 (N_2222,N_1206,N_1269);
or U2223 (N_2223,N_1750,N_1673);
nor U2224 (N_2224,N_1584,N_1581);
or U2225 (N_2225,N_1646,N_1699);
nand U2226 (N_2226,N_1278,N_1661);
or U2227 (N_2227,N_1759,N_1514);
and U2228 (N_2228,N_1513,N_1370);
and U2229 (N_2229,N_1343,N_1260);
and U2230 (N_2230,N_1790,N_1743);
nor U2231 (N_2231,N_1228,N_1701);
nor U2232 (N_2232,N_1511,N_1281);
and U2233 (N_2233,N_1695,N_1581);
and U2234 (N_2234,N_1683,N_1786);
and U2235 (N_2235,N_1293,N_1707);
and U2236 (N_2236,N_1210,N_1461);
nand U2237 (N_2237,N_1352,N_1758);
nor U2238 (N_2238,N_1332,N_1406);
nor U2239 (N_2239,N_1498,N_1388);
nand U2240 (N_2240,N_1326,N_1216);
nor U2241 (N_2241,N_1607,N_1683);
and U2242 (N_2242,N_1469,N_1632);
or U2243 (N_2243,N_1335,N_1307);
or U2244 (N_2244,N_1686,N_1244);
nand U2245 (N_2245,N_1576,N_1615);
or U2246 (N_2246,N_1227,N_1585);
and U2247 (N_2247,N_1560,N_1539);
nor U2248 (N_2248,N_1690,N_1444);
or U2249 (N_2249,N_1299,N_1555);
or U2250 (N_2250,N_1263,N_1235);
nor U2251 (N_2251,N_1334,N_1259);
nand U2252 (N_2252,N_1250,N_1648);
or U2253 (N_2253,N_1485,N_1480);
and U2254 (N_2254,N_1651,N_1624);
and U2255 (N_2255,N_1783,N_1756);
nor U2256 (N_2256,N_1335,N_1261);
and U2257 (N_2257,N_1544,N_1614);
nor U2258 (N_2258,N_1732,N_1309);
nand U2259 (N_2259,N_1725,N_1357);
nor U2260 (N_2260,N_1251,N_1658);
and U2261 (N_2261,N_1401,N_1235);
and U2262 (N_2262,N_1435,N_1395);
or U2263 (N_2263,N_1436,N_1235);
and U2264 (N_2264,N_1347,N_1245);
and U2265 (N_2265,N_1757,N_1538);
xor U2266 (N_2266,N_1328,N_1376);
or U2267 (N_2267,N_1717,N_1304);
nand U2268 (N_2268,N_1213,N_1639);
or U2269 (N_2269,N_1618,N_1789);
and U2270 (N_2270,N_1467,N_1540);
nand U2271 (N_2271,N_1313,N_1780);
nand U2272 (N_2272,N_1747,N_1683);
or U2273 (N_2273,N_1512,N_1362);
nand U2274 (N_2274,N_1426,N_1607);
and U2275 (N_2275,N_1313,N_1761);
nand U2276 (N_2276,N_1601,N_1401);
nor U2277 (N_2277,N_1294,N_1335);
nor U2278 (N_2278,N_1786,N_1624);
nor U2279 (N_2279,N_1612,N_1610);
and U2280 (N_2280,N_1282,N_1528);
or U2281 (N_2281,N_1636,N_1656);
and U2282 (N_2282,N_1341,N_1518);
nor U2283 (N_2283,N_1785,N_1499);
and U2284 (N_2284,N_1380,N_1462);
and U2285 (N_2285,N_1523,N_1346);
and U2286 (N_2286,N_1470,N_1622);
nand U2287 (N_2287,N_1493,N_1518);
and U2288 (N_2288,N_1710,N_1407);
or U2289 (N_2289,N_1465,N_1576);
nand U2290 (N_2290,N_1327,N_1457);
nor U2291 (N_2291,N_1779,N_1407);
and U2292 (N_2292,N_1586,N_1331);
and U2293 (N_2293,N_1385,N_1249);
nor U2294 (N_2294,N_1224,N_1709);
or U2295 (N_2295,N_1333,N_1798);
or U2296 (N_2296,N_1329,N_1757);
and U2297 (N_2297,N_1388,N_1240);
or U2298 (N_2298,N_1587,N_1531);
nand U2299 (N_2299,N_1357,N_1595);
or U2300 (N_2300,N_1713,N_1266);
or U2301 (N_2301,N_1523,N_1240);
nor U2302 (N_2302,N_1622,N_1606);
or U2303 (N_2303,N_1485,N_1479);
or U2304 (N_2304,N_1507,N_1631);
nand U2305 (N_2305,N_1692,N_1712);
nand U2306 (N_2306,N_1716,N_1775);
and U2307 (N_2307,N_1639,N_1378);
nand U2308 (N_2308,N_1402,N_1523);
nor U2309 (N_2309,N_1341,N_1467);
nor U2310 (N_2310,N_1707,N_1630);
or U2311 (N_2311,N_1751,N_1262);
and U2312 (N_2312,N_1395,N_1710);
nand U2313 (N_2313,N_1440,N_1732);
or U2314 (N_2314,N_1751,N_1316);
nor U2315 (N_2315,N_1209,N_1662);
and U2316 (N_2316,N_1262,N_1362);
and U2317 (N_2317,N_1651,N_1203);
or U2318 (N_2318,N_1406,N_1782);
nor U2319 (N_2319,N_1597,N_1283);
nand U2320 (N_2320,N_1274,N_1779);
and U2321 (N_2321,N_1370,N_1440);
nor U2322 (N_2322,N_1618,N_1411);
nand U2323 (N_2323,N_1311,N_1529);
or U2324 (N_2324,N_1539,N_1436);
nand U2325 (N_2325,N_1538,N_1289);
or U2326 (N_2326,N_1364,N_1460);
nor U2327 (N_2327,N_1396,N_1527);
and U2328 (N_2328,N_1468,N_1712);
or U2329 (N_2329,N_1753,N_1780);
xnor U2330 (N_2330,N_1578,N_1379);
nand U2331 (N_2331,N_1681,N_1569);
or U2332 (N_2332,N_1398,N_1726);
nor U2333 (N_2333,N_1424,N_1298);
nor U2334 (N_2334,N_1738,N_1217);
nand U2335 (N_2335,N_1290,N_1433);
nand U2336 (N_2336,N_1454,N_1339);
nand U2337 (N_2337,N_1319,N_1579);
nor U2338 (N_2338,N_1255,N_1494);
and U2339 (N_2339,N_1701,N_1674);
or U2340 (N_2340,N_1289,N_1384);
and U2341 (N_2341,N_1363,N_1488);
and U2342 (N_2342,N_1328,N_1637);
nor U2343 (N_2343,N_1485,N_1683);
and U2344 (N_2344,N_1337,N_1259);
or U2345 (N_2345,N_1297,N_1541);
nor U2346 (N_2346,N_1506,N_1256);
or U2347 (N_2347,N_1677,N_1294);
or U2348 (N_2348,N_1591,N_1231);
and U2349 (N_2349,N_1391,N_1561);
or U2350 (N_2350,N_1525,N_1540);
and U2351 (N_2351,N_1421,N_1501);
nand U2352 (N_2352,N_1791,N_1252);
or U2353 (N_2353,N_1670,N_1673);
and U2354 (N_2354,N_1371,N_1454);
or U2355 (N_2355,N_1479,N_1463);
nor U2356 (N_2356,N_1513,N_1488);
nor U2357 (N_2357,N_1774,N_1401);
and U2358 (N_2358,N_1642,N_1437);
nand U2359 (N_2359,N_1768,N_1408);
nand U2360 (N_2360,N_1359,N_1353);
nor U2361 (N_2361,N_1611,N_1354);
or U2362 (N_2362,N_1679,N_1793);
and U2363 (N_2363,N_1706,N_1207);
nand U2364 (N_2364,N_1244,N_1417);
and U2365 (N_2365,N_1406,N_1779);
or U2366 (N_2366,N_1745,N_1293);
nor U2367 (N_2367,N_1342,N_1580);
and U2368 (N_2368,N_1607,N_1680);
and U2369 (N_2369,N_1393,N_1436);
and U2370 (N_2370,N_1435,N_1436);
and U2371 (N_2371,N_1715,N_1687);
nor U2372 (N_2372,N_1773,N_1735);
and U2373 (N_2373,N_1380,N_1523);
nand U2374 (N_2374,N_1699,N_1768);
and U2375 (N_2375,N_1521,N_1458);
nand U2376 (N_2376,N_1419,N_1546);
or U2377 (N_2377,N_1584,N_1771);
nand U2378 (N_2378,N_1463,N_1354);
nor U2379 (N_2379,N_1707,N_1446);
and U2380 (N_2380,N_1391,N_1650);
nor U2381 (N_2381,N_1740,N_1651);
or U2382 (N_2382,N_1763,N_1362);
nand U2383 (N_2383,N_1332,N_1243);
nand U2384 (N_2384,N_1783,N_1429);
nor U2385 (N_2385,N_1344,N_1700);
and U2386 (N_2386,N_1477,N_1258);
nor U2387 (N_2387,N_1642,N_1555);
and U2388 (N_2388,N_1219,N_1792);
or U2389 (N_2389,N_1324,N_1680);
xnor U2390 (N_2390,N_1630,N_1281);
xnor U2391 (N_2391,N_1771,N_1264);
nand U2392 (N_2392,N_1218,N_1302);
nand U2393 (N_2393,N_1544,N_1221);
xnor U2394 (N_2394,N_1322,N_1377);
nor U2395 (N_2395,N_1311,N_1307);
or U2396 (N_2396,N_1560,N_1672);
nand U2397 (N_2397,N_1383,N_1340);
or U2398 (N_2398,N_1493,N_1221);
or U2399 (N_2399,N_1519,N_1458);
or U2400 (N_2400,N_2028,N_1817);
nand U2401 (N_2401,N_1821,N_2367);
nor U2402 (N_2402,N_2214,N_1888);
nand U2403 (N_2403,N_2198,N_2130);
and U2404 (N_2404,N_2396,N_2019);
nand U2405 (N_2405,N_2320,N_2277);
or U2406 (N_2406,N_2363,N_1879);
nand U2407 (N_2407,N_1987,N_1921);
nand U2408 (N_2408,N_2301,N_2240);
nand U2409 (N_2409,N_1918,N_1942);
nand U2410 (N_2410,N_2316,N_2163);
xnor U2411 (N_2411,N_2091,N_2058);
nand U2412 (N_2412,N_1800,N_2179);
nor U2413 (N_2413,N_2069,N_2232);
nand U2414 (N_2414,N_2144,N_1899);
and U2415 (N_2415,N_2123,N_1859);
or U2416 (N_2416,N_2215,N_1949);
nor U2417 (N_2417,N_2095,N_2221);
nor U2418 (N_2418,N_1841,N_2298);
nor U2419 (N_2419,N_2013,N_1816);
nand U2420 (N_2420,N_1901,N_1881);
and U2421 (N_2421,N_2390,N_1847);
nor U2422 (N_2422,N_1979,N_2098);
and U2423 (N_2423,N_2127,N_2300);
or U2424 (N_2424,N_1951,N_1889);
nor U2425 (N_2425,N_2336,N_2334);
nor U2426 (N_2426,N_1833,N_2016);
nor U2427 (N_2427,N_1999,N_2075);
or U2428 (N_2428,N_1933,N_2242);
or U2429 (N_2429,N_2158,N_1935);
xor U2430 (N_2430,N_2128,N_2213);
or U2431 (N_2431,N_1814,N_1818);
or U2432 (N_2432,N_2072,N_2211);
xor U2433 (N_2433,N_1971,N_2088);
nor U2434 (N_2434,N_2278,N_2041);
nand U2435 (N_2435,N_1939,N_1848);
or U2436 (N_2436,N_2011,N_2249);
nand U2437 (N_2437,N_2138,N_2023);
nand U2438 (N_2438,N_2205,N_2150);
nor U2439 (N_2439,N_2100,N_1916);
or U2440 (N_2440,N_2229,N_1801);
and U2441 (N_2441,N_2122,N_2006);
and U2442 (N_2442,N_2148,N_1895);
and U2443 (N_2443,N_2125,N_2385);
or U2444 (N_2444,N_2237,N_1956);
nand U2445 (N_2445,N_1910,N_2197);
xor U2446 (N_2446,N_2105,N_1970);
and U2447 (N_2447,N_2387,N_1966);
nor U2448 (N_2448,N_2145,N_2044);
nand U2449 (N_2449,N_1840,N_1946);
nor U2450 (N_2450,N_2021,N_2292);
and U2451 (N_2451,N_2296,N_1976);
nand U2452 (N_2452,N_2132,N_1823);
and U2453 (N_2453,N_2331,N_1986);
or U2454 (N_2454,N_2370,N_1827);
nor U2455 (N_2455,N_2110,N_2184);
nand U2456 (N_2456,N_1891,N_2384);
nor U2457 (N_2457,N_2012,N_1957);
nor U2458 (N_2458,N_2297,N_2046);
or U2459 (N_2459,N_2313,N_1968);
xnor U2460 (N_2460,N_1866,N_2325);
or U2461 (N_2461,N_2056,N_2020);
and U2462 (N_2462,N_2225,N_1998);
nor U2463 (N_2463,N_2305,N_1996);
nand U2464 (N_2464,N_1914,N_1884);
and U2465 (N_2465,N_1872,N_2053);
and U2466 (N_2466,N_2260,N_1948);
or U2467 (N_2467,N_2285,N_1836);
and U2468 (N_2468,N_2193,N_2171);
and U2469 (N_2469,N_2153,N_2040);
xnor U2470 (N_2470,N_2323,N_2361);
or U2471 (N_2471,N_1977,N_2365);
nor U2472 (N_2472,N_2084,N_1927);
and U2473 (N_2473,N_2154,N_2177);
nor U2474 (N_2474,N_2061,N_1932);
xnor U2475 (N_2475,N_2135,N_2005);
and U2476 (N_2476,N_2304,N_2085);
or U2477 (N_2477,N_2227,N_2126);
nand U2478 (N_2478,N_2342,N_2347);
and U2479 (N_2479,N_2322,N_2048);
nor U2480 (N_2480,N_2341,N_2386);
nor U2481 (N_2481,N_1940,N_2137);
or U2482 (N_2482,N_2271,N_2243);
nor U2483 (N_2483,N_2395,N_1911);
nand U2484 (N_2484,N_1943,N_1965);
nor U2485 (N_2485,N_1984,N_1964);
nor U2486 (N_2486,N_2355,N_1804);
and U2487 (N_2487,N_2199,N_2094);
and U2488 (N_2488,N_2168,N_2017);
nor U2489 (N_2489,N_1845,N_2228);
nand U2490 (N_2490,N_2121,N_1862);
nor U2491 (N_2491,N_1811,N_2287);
and U2492 (N_2492,N_1885,N_2022);
and U2493 (N_2493,N_2052,N_1808);
nor U2494 (N_2494,N_2303,N_2245);
nand U2495 (N_2495,N_1989,N_1991);
nor U2496 (N_2496,N_2230,N_1950);
nor U2497 (N_2497,N_2160,N_2062);
nor U2498 (N_2498,N_2195,N_2210);
nor U2499 (N_2499,N_2087,N_2073);
or U2500 (N_2500,N_2155,N_2343);
or U2501 (N_2501,N_2004,N_2328);
and U2502 (N_2502,N_2254,N_2136);
xor U2503 (N_2503,N_2166,N_2108);
nor U2504 (N_2504,N_2309,N_2369);
xnor U2505 (N_2505,N_2172,N_2295);
and U2506 (N_2506,N_1887,N_2180);
or U2507 (N_2507,N_2200,N_2247);
or U2508 (N_2508,N_1819,N_2008);
or U2509 (N_2509,N_2364,N_2324);
or U2510 (N_2510,N_2076,N_2266);
nand U2511 (N_2511,N_2031,N_1923);
and U2512 (N_2512,N_1997,N_1904);
or U2513 (N_2513,N_1825,N_2107);
or U2514 (N_2514,N_1969,N_2169);
nand U2515 (N_2515,N_2290,N_1805);
and U2516 (N_2516,N_1907,N_2000);
nor U2517 (N_2517,N_2173,N_2238);
nand U2518 (N_2518,N_2188,N_2143);
nand U2519 (N_2519,N_2042,N_2190);
nand U2520 (N_2520,N_1876,N_2033);
and U2521 (N_2521,N_1990,N_2070);
xnor U2522 (N_2522,N_2124,N_2244);
nor U2523 (N_2523,N_1936,N_2089);
or U2524 (N_2524,N_2256,N_2079);
nand U2525 (N_2525,N_2026,N_2083);
nor U2526 (N_2526,N_2257,N_2286);
nor U2527 (N_2527,N_1865,N_2362);
nand U2528 (N_2528,N_2332,N_2263);
and U2529 (N_2529,N_2111,N_2201);
or U2530 (N_2530,N_2183,N_1992);
xor U2531 (N_2531,N_2035,N_2146);
nand U2532 (N_2532,N_2038,N_1878);
or U2533 (N_2533,N_1812,N_2139);
nand U2534 (N_2534,N_1975,N_2078);
nand U2535 (N_2535,N_1851,N_2253);
or U2536 (N_2536,N_1852,N_2231);
nor U2537 (N_2537,N_2092,N_1826);
nand U2538 (N_2538,N_2330,N_2074);
xor U2539 (N_2539,N_1874,N_1974);
nor U2540 (N_2540,N_2233,N_2064);
nor U2541 (N_2541,N_2359,N_1839);
nand U2542 (N_2542,N_2009,N_2115);
nor U2543 (N_2543,N_2134,N_2170);
and U2544 (N_2544,N_2186,N_2161);
or U2545 (N_2545,N_2374,N_2120);
or U2546 (N_2546,N_2152,N_2372);
nand U2547 (N_2547,N_1810,N_1820);
nand U2548 (N_2548,N_2222,N_2279);
nor U2549 (N_2549,N_2175,N_1925);
or U2550 (N_2550,N_1880,N_2375);
and U2551 (N_2551,N_2234,N_1963);
nand U2552 (N_2552,N_2348,N_1838);
nor U2553 (N_2553,N_1831,N_2142);
nor U2554 (N_2554,N_2015,N_2340);
nor U2555 (N_2555,N_1843,N_2101);
nor U2556 (N_2556,N_2209,N_2051);
or U2557 (N_2557,N_1917,N_2093);
or U2558 (N_2558,N_2356,N_2252);
nor U2559 (N_2559,N_1875,N_2068);
or U2560 (N_2560,N_2259,N_2036);
or U2561 (N_2561,N_1985,N_2306);
nor U2562 (N_2562,N_2357,N_1908);
or U2563 (N_2563,N_2147,N_1815);
or U2564 (N_2564,N_2001,N_2241);
or U2565 (N_2565,N_2319,N_2333);
nand U2566 (N_2566,N_2294,N_2371);
and U2567 (N_2567,N_2315,N_2381);
or U2568 (N_2568,N_1824,N_1809);
and U2569 (N_2569,N_1941,N_1929);
and U2570 (N_2570,N_2077,N_2344);
or U2571 (N_2571,N_1954,N_2182);
nand U2572 (N_2572,N_2339,N_2276);
or U2573 (N_2573,N_1822,N_1897);
and U2574 (N_2574,N_1924,N_2030);
nor U2575 (N_2575,N_2149,N_2216);
nor U2576 (N_2576,N_1803,N_2226);
or U2577 (N_2577,N_2258,N_2174);
nand U2578 (N_2578,N_2368,N_1928);
nor U2579 (N_2579,N_2164,N_1861);
nand U2580 (N_2580,N_1994,N_2097);
and U2581 (N_2581,N_1903,N_2312);
nor U2582 (N_2582,N_2165,N_2099);
nor U2583 (N_2583,N_2102,N_1930);
nand U2584 (N_2584,N_1909,N_2047);
and U2585 (N_2585,N_1894,N_2194);
and U2586 (N_2586,N_2255,N_2321);
nor U2587 (N_2587,N_2103,N_1853);
or U2588 (N_2588,N_1871,N_2379);
and U2589 (N_2589,N_2350,N_2060);
nand U2590 (N_2590,N_2129,N_2086);
or U2591 (N_2591,N_1902,N_1867);
or U2592 (N_2592,N_2131,N_2096);
or U2593 (N_2593,N_1882,N_2159);
xnor U2594 (N_2594,N_1858,N_1958);
nand U2595 (N_2595,N_1883,N_1906);
or U2596 (N_2596,N_1868,N_2311);
or U2597 (N_2597,N_1886,N_1983);
and U2598 (N_2598,N_2349,N_1857);
or U2599 (N_2599,N_1869,N_2187);
nand U2600 (N_2600,N_1849,N_1898);
nand U2601 (N_2601,N_2081,N_2066);
nand U2602 (N_2602,N_2265,N_2289);
and U2603 (N_2603,N_1813,N_1850);
nand U2604 (N_2604,N_2029,N_1860);
or U2605 (N_2605,N_1828,N_2220);
nor U2606 (N_2606,N_2267,N_1972);
and U2607 (N_2607,N_2112,N_2351);
and U2608 (N_2608,N_2065,N_2394);
and U2609 (N_2609,N_2327,N_2273);
nand U2610 (N_2610,N_2104,N_2151);
nor U2611 (N_2611,N_1959,N_1900);
or U2612 (N_2612,N_2141,N_2235);
and U2613 (N_2613,N_1913,N_2007);
nand U2614 (N_2614,N_2025,N_2185);
or U2615 (N_2615,N_2397,N_2354);
and U2616 (N_2616,N_2281,N_2133);
and U2617 (N_2617,N_2119,N_2360);
or U2618 (N_2618,N_2251,N_2314);
nor U2619 (N_2619,N_1806,N_2291);
and U2620 (N_2620,N_1870,N_2157);
and U2621 (N_2621,N_2326,N_2398);
nor U2622 (N_2622,N_2204,N_2176);
and U2623 (N_2623,N_1944,N_1807);
or U2624 (N_2624,N_2318,N_2202);
nor U2625 (N_2625,N_2037,N_1835);
nand U2626 (N_2626,N_1905,N_1896);
or U2627 (N_2627,N_2071,N_2307);
and U2628 (N_2628,N_1982,N_2346);
nor U2629 (N_2629,N_1978,N_2399);
and U2630 (N_2630,N_2329,N_2140);
or U2631 (N_2631,N_1837,N_2208);
nand U2632 (N_2632,N_2181,N_2293);
and U2633 (N_2633,N_2014,N_2106);
nor U2634 (N_2634,N_2239,N_1973);
and U2635 (N_2635,N_1863,N_1953);
and U2636 (N_2636,N_2063,N_1892);
nand U2637 (N_2637,N_2270,N_2080);
nand U2638 (N_2638,N_2219,N_2049);
xnor U2639 (N_2639,N_1915,N_2217);
and U2640 (N_2640,N_2032,N_2027);
nand U2641 (N_2641,N_1829,N_2310);
and U2642 (N_2642,N_2280,N_1952);
nand U2643 (N_2643,N_2380,N_1912);
xnor U2644 (N_2644,N_1980,N_2335);
or U2645 (N_2645,N_2043,N_1955);
and U2646 (N_2646,N_2382,N_1830);
or U2647 (N_2647,N_2236,N_2116);
nor U2648 (N_2648,N_2352,N_2261);
or U2649 (N_2649,N_1802,N_1844);
or U2650 (N_2650,N_2248,N_2057);
and U2651 (N_2651,N_2250,N_2262);
or U2652 (N_2652,N_2189,N_2376);
xor U2653 (N_2653,N_2067,N_2109);
nor U2654 (N_2654,N_1890,N_2167);
nor U2655 (N_2655,N_1961,N_2393);
and U2656 (N_2656,N_2338,N_2118);
or U2657 (N_2657,N_2207,N_2272);
nor U2658 (N_2658,N_2358,N_1962);
or U2659 (N_2659,N_2090,N_2366);
nand U2660 (N_2660,N_2392,N_1993);
or U2661 (N_2661,N_2218,N_1945);
or U2662 (N_2662,N_1842,N_2224);
or U2663 (N_2663,N_2059,N_1873);
and U2664 (N_2664,N_2082,N_2018);
nor U2665 (N_2665,N_2383,N_1947);
nor U2666 (N_2666,N_2345,N_1995);
or U2667 (N_2667,N_2039,N_2113);
nor U2668 (N_2668,N_1864,N_2389);
or U2669 (N_2669,N_2388,N_1934);
or U2670 (N_2670,N_1931,N_2288);
or U2671 (N_2671,N_2283,N_2045);
and U2672 (N_2672,N_1893,N_2002);
nand U2673 (N_2673,N_2282,N_2246);
and U2674 (N_2674,N_2178,N_2050);
or U2675 (N_2675,N_1919,N_2117);
and U2676 (N_2676,N_2114,N_2308);
nor U2677 (N_2677,N_2391,N_2034);
nor U2678 (N_2678,N_2269,N_1981);
or U2679 (N_2679,N_2203,N_2192);
or U2680 (N_2680,N_1988,N_2055);
or U2681 (N_2681,N_1877,N_2302);
nor U2682 (N_2682,N_2284,N_1960);
nand U2683 (N_2683,N_2353,N_2162);
nand U2684 (N_2684,N_2206,N_1856);
and U2685 (N_2685,N_2373,N_1846);
nand U2686 (N_2686,N_2010,N_1920);
and U2687 (N_2687,N_1832,N_1926);
nor U2688 (N_2688,N_2377,N_2264);
or U2689 (N_2689,N_2024,N_1938);
nand U2690 (N_2690,N_1937,N_2275);
nand U2691 (N_2691,N_2378,N_1855);
nor U2692 (N_2692,N_2337,N_2156);
or U2693 (N_2693,N_2212,N_1854);
nor U2694 (N_2694,N_2191,N_2223);
nand U2695 (N_2695,N_1967,N_2268);
or U2696 (N_2696,N_1834,N_1922);
or U2697 (N_2697,N_2054,N_2003);
xnor U2698 (N_2698,N_2274,N_2299);
nor U2699 (N_2699,N_2196,N_2317);
or U2700 (N_2700,N_1976,N_1943);
nand U2701 (N_2701,N_1857,N_2043);
and U2702 (N_2702,N_2321,N_1886);
nor U2703 (N_2703,N_2161,N_1829);
nand U2704 (N_2704,N_2272,N_1986);
or U2705 (N_2705,N_2161,N_2125);
nor U2706 (N_2706,N_2313,N_2189);
or U2707 (N_2707,N_2266,N_2133);
or U2708 (N_2708,N_2313,N_2336);
and U2709 (N_2709,N_1818,N_1957);
and U2710 (N_2710,N_2139,N_2163);
and U2711 (N_2711,N_2376,N_2204);
nand U2712 (N_2712,N_1823,N_2030);
or U2713 (N_2713,N_2323,N_1803);
nor U2714 (N_2714,N_2303,N_1989);
or U2715 (N_2715,N_1827,N_2195);
and U2716 (N_2716,N_2374,N_1939);
nand U2717 (N_2717,N_2130,N_2176);
or U2718 (N_2718,N_1915,N_2307);
nor U2719 (N_2719,N_2229,N_2121);
or U2720 (N_2720,N_2089,N_2198);
nor U2721 (N_2721,N_2101,N_1824);
nand U2722 (N_2722,N_1974,N_1839);
nor U2723 (N_2723,N_2267,N_2285);
or U2724 (N_2724,N_2139,N_2207);
nor U2725 (N_2725,N_1810,N_2157);
or U2726 (N_2726,N_2267,N_1845);
nand U2727 (N_2727,N_2378,N_1853);
and U2728 (N_2728,N_2113,N_1997);
nand U2729 (N_2729,N_2313,N_2353);
or U2730 (N_2730,N_2262,N_1802);
or U2731 (N_2731,N_2336,N_1985);
and U2732 (N_2732,N_1804,N_1880);
or U2733 (N_2733,N_1838,N_2032);
nor U2734 (N_2734,N_2020,N_2100);
nor U2735 (N_2735,N_2004,N_2124);
nand U2736 (N_2736,N_2228,N_2079);
nor U2737 (N_2737,N_1811,N_2200);
and U2738 (N_2738,N_2133,N_2148);
nor U2739 (N_2739,N_2210,N_2111);
or U2740 (N_2740,N_1947,N_2045);
nand U2741 (N_2741,N_2376,N_1994);
or U2742 (N_2742,N_1848,N_2194);
and U2743 (N_2743,N_2344,N_1847);
nor U2744 (N_2744,N_2371,N_2210);
nand U2745 (N_2745,N_2372,N_1837);
nand U2746 (N_2746,N_2304,N_2121);
or U2747 (N_2747,N_2274,N_1844);
nand U2748 (N_2748,N_2136,N_2139);
nor U2749 (N_2749,N_1974,N_2011);
and U2750 (N_2750,N_2273,N_1833);
and U2751 (N_2751,N_1835,N_1957);
nand U2752 (N_2752,N_2384,N_2127);
and U2753 (N_2753,N_1932,N_2143);
nor U2754 (N_2754,N_2222,N_2359);
or U2755 (N_2755,N_2398,N_2311);
and U2756 (N_2756,N_2030,N_2358);
or U2757 (N_2757,N_2165,N_2239);
nor U2758 (N_2758,N_2091,N_2326);
and U2759 (N_2759,N_2170,N_1818);
or U2760 (N_2760,N_2077,N_1934);
or U2761 (N_2761,N_1839,N_1932);
and U2762 (N_2762,N_2020,N_1822);
nand U2763 (N_2763,N_2112,N_1818);
or U2764 (N_2764,N_2062,N_1816);
xor U2765 (N_2765,N_2036,N_1856);
nand U2766 (N_2766,N_2216,N_2119);
nand U2767 (N_2767,N_1908,N_2010);
nor U2768 (N_2768,N_2336,N_2342);
or U2769 (N_2769,N_2149,N_1843);
or U2770 (N_2770,N_2115,N_2266);
nand U2771 (N_2771,N_1991,N_2109);
or U2772 (N_2772,N_2013,N_2355);
or U2773 (N_2773,N_2385,N_2148);
nand U2774 (N_2774,N_2118,N_2172);
and U2775 (N_2775,N_2053,N_2080);
nand U2776 (N_2776,N_2012,N_1979);
and U2777 (N_2777,N_2288,N_2246);
or U2778 (N_2778,N_1998,N_2045);
or U2779 (N_2779,N_1836,N_2072);
or U2780 (N_2780,N_2240,N_1894);
and U2781 (N_2781,N_2281,N_2207);
nand U2782 (N_2782,N_1960,N_2005);
nor U2783 (N_2783,N_1964,N_2027);
nand U2784 (N_2784,N_2300,N_2056);
nor U2785 (N_2785,N_2396,N_1912);
and U2786 (N_2786,N_2369,N_2067);
nor U2787 (N_2787,N_2013,N_2255);
and U2788 (N_2788,N_1852,N_2238);
or U2789 (N_2789,N_1807,N_1916);
nand U2790 (N_2790,N_1916,N_2108);
nand U2791 (N_2791,N_1815,N_1990);
or U2792 (N_2792,N_2190,N_2003);
nor U2793 (N_2793,N_2278,N_2000);
nand U2794 (N_2794,N_2234,N_1952);
xnor U2795 (N_2795,N_1807,N_2287);
or U2796 (N_2796,N_1843,N_2315);
nor U2797 (N_2797,N_2182,N_2298);
nand U2798 (N_2798,N_1902,N_1864);
nor U2799 (N_2799,N_2169,N_2118);
or U2800 (N_2800,N_1832,N_2057);
nor U2801 (N_2801,N_1915,N_1839);
nor U2802 (N_2802,N_2382,N_2149);
nand U2803 (N_2803,N_2219,N_1862);
nand U2804 (N_2804,N_2203,N_2127);
or U2805 (N_2805,N_1944,N_2105);
or U2806 (N_2806,N_2030,N_2177);
or U2807 (N_2807,N_2241,N_1945);
and U2808 (N_2808,N_2095,N_2336);
or U2809 (N_2809,N_2085,N_2190);
or U2810 (N_2810,N_2393,N_1969);
and U2811 (N_2811,N_2105,N_2318);
nand U2812 (N_2812,N_2311,N_2258);
nor U2813 (N_2813,N_2370,N_1868);
or U2814 (N_2814,N_2242,N_2007);
nand U2815 (N_2815,N_1860,N_2330);
and U2816 (N_2816,N_1832,N_2049);
nand U2817 (N_2817,N_1810,N_1984);
or U2818 (N_2818,N_2167,N_2161);
and U2819 (N_2819,N_2287,N_2182);
and U2820 (N_2820,N_2173,N_1819);
nor U2821 (N_2821,N_2242,N_2352);
or U2822 (N_2822,N_2350,N_2130);
or U2823 (N_2823,N_1912,N_1859);
and U2824 (N_2824,N_2141,N_2148);
xor U2825 (N_2825,N_1915,N_2218);
and U2826 (N_2826,N_2077,N_2141);
nor U2827 (N_2827,N_1809,N_2338);
and U2828 (N_2828,N_1803,N_2329);
or U2829 (N_2829,N_2238,N_1985);
nand U2830 (N_2830,N_2113,N_1889);
nand U2831 (N_2831,N_2189,N_1851);
nand U2832 (N_2832,N_2393,N_2235);
nand U2833 (N_2833,N_1989,N_2117);
and U2834 (N_2834,N_2074,N_1867);
or U2835 (N_2835,N_1885,N_2118);
or U2836 (N_2836,N_2091,N_2210);
or U2837 (N_2837,N_2251,N_1906);
nand U2838 (N_2838,N_1892,N_1874);
and U2839 (N_2839,N_1919,N_2131);
and U2840 (N_2840,N_2188,N_2251);
or U2841 (N_2841,N_2116,N_2042);
and U2842 (N_2842,N_2284,N_1917);
or U2843 (N_2843,N_2222,N_2070);
and U2844 (N_2844,N_2121,N_2389);
or U2845 (N_2845,N_1885,N_2135);
or U2846 (N_2846,N_2169,N_2245);
nand U2847 (N_2847,N_1898,N_2334);
nor U2848 (N_2848,N_1843,N_2269);
xor U2849 (N_2849,N_1920,N_2340);
or U2850 (N_2850,N_2333,N_1877);
nand U2851 (N_2851,N_1833,N_2271);
nor U2852 (N_2852,N_1839,N_2159);
nor U2853 (N_2853,N_2375,N_2148);
and U2854 (N_2854,N_2250,N_2042);
nor U2855 (N_2855,N_2280,N_2128);
and U2856 (N_2856,N_1882,N_2084);
or U2857 (N_2857,N_2012,N_2392);
or U2858 (N_2858,N_2166,N_1990);
and U2859 (N_2859,N_2091,N_2152);
and U2860 (N_2860,N_1902,N_2220);
nor U2861 (N_2861,N_2284,N_2096);
nand U2862 (N_2862,N_2192,N_2169);
nor U2863 (N_2863,N_2194,N_2383);
nor U2864 (N_2864,N_1859,N_2012);
or U2865 (N_2865,N_1991,N_2099);
and U2866 (N_2866,N_1931,N_2295);
nand U2867 (N_2867,N_2073,N_1992);
or U2868 (N_2868,N_2201,N_1867);
and U2869 (N_2869,N_2221,N_2002);
nor U2870 (N_2870,N_2204,N_1896);
or U2871 (N_2871,N_2323,N_1957);
nand U2872 (N_2872,N_1808,N_1984);
nand U2873 (N_2873,N_2081,N_1800);
or U2874 (N_2874,N_2065,N_2103);
and U2875 (N_2875,N_2332,N_2087);
nand U2876 (N_2876,N_2274,N_2007);
nor U2877 (N_2877,N_2182,N_2297);
nand U2878 (N_2878,N_1915,N_2232);
nor U2879 (N_2879,N_1820,N_2245);
or U2880 (N_2880,N_2292,N_2118);
and U2881 (N_2881,N_1991,N_2229);
nor U2882 (N_2882,N_1849,N_2332);
nand U2883 (N_2883,N_2106,N_2047);
nand U2884 (N_2884,N_1860,N_1828);
xor U2885 (N_2885,N_2266,N_2003);
or U2886 (N_2886,N_1966,N_2334);
and U2887 (N_2887,N_1861,N_2123);
nor U2888 (N_2888,N_2100,N_2338);
nor U2889 (N_2889,N_2259,N_1968);
or U2890 (N_2890,N_1962,N_2179);
nand U2891 (N_2891,N_1900,N_1840);
and U2892 (N_2892,N_2031,N_2351);
nor U2893 (N_2893,N_1940,N_2146);
nand U2894 (N_2894,N_2024,N_1942);
nor U2895 (N_2895,N_2183,N_2150);
or U2896 (N_2896,N_1818,N_2103);
and U2897 (N_2897,N_1971,N_2151);
nand U2898 (N_2898,N_1936,N_1942);
or U2899 (N_2899,N_2046,N_1823);
or U2900 (N_2900,N_2262,N_2360);
and U2901 (N_2901,N_1946,N_2173);
nand U2902 (N_2902,N_1977,N_1810);
or U2903 (N_2903,N_1857,N_2326);
nor U2904 (N_2904,N_1867,N_2399);
nor U2905 (N_2905,N_2119,N_1942);
and U2906 (N_2906,N_2225,N_2346);
nor U2907 (N_2907,N_2183,N_2316);
nor U2908 (N_2908,N_2067,N_1848);
nor U2909 (N_2909,N_2177,N_1880);
or U2910 (N_2910,N_2330,N_2097);
nor U2911 (N_2911,N_2060,N_2278);
nor U2912 (N_2912,N_2167,N_2222);
or U2913 (N_2913,N_2396,N_1832);
nand U2914 (N_2914,N_1926,N_2295);
nand U2915 (N_2915,N_1893,N_2014);
nor U2916 (N_2916,N_2053,N_2170);
nand U2917 (N_2917,N_2247,N_1999);
nor U2918 (N_2918,N_2037,N_2214);
nand U2919 (N_2919,N_1906,N_1930);
nand U2920 (N_2920,N_2183,N_1939);
or U2921 (N_2921,N_2084,N_1957);
nor U2922 (N_2922,N_2393,N_2105);
nand U2923 (N_2923,N_2186,N_2210);
nor U2924 (N_2924,N_1898,N_2067);
nand U2925 (N_2925,N_2200,N_1955);
or U2926 (N_2926,N_2287,N_1848);
and U2927 (N_2927,N_1877,N_2246);
nand U2928 (N_2928,N_2146,N_1816);
or U2929 (N_2929,N_1856,N_2180);
xnor U2930 (N_2930,N_2223,N_1843);
nor U2931 (N_2931,N_1850,N_2020);
or U2932 (N_2932,N_2074,N_1917);
nor U2933 (N_2933,N_2381,N_2339);
nand U2934 (N_2934,N_2329,N_2009);
and U2935 (N_2935,N_1952,N_2371);
nor U2936 (N_2936,N_1967,N_2385);
and U2937 (N_2937,N_2234,N_2226);
and U2938 (N_2938,N_2062,N_1930);
or U2939 (N_2939,N_2309,N_1847);
nand U2940 (N_2940,N_2009,N_2074);
nor U2941 (N_2941,N_1996,N_2026);
or U2942 (N_2942,N_2248,N_2076);
and U2943 (N_2943,N_1988,N_2334);
nand U2944 (N_2944,N_1871,N_2211);
or U2945 (N_2945,N_2099,N_2387);
and U2946 (N_2946,N_1909,N_1991);
nand U2947 (N_2947,N_1996,N_2025);
nand U2948 (N_2948,N_1898,N_2299);
and U2949 (N_2949,N_2386,N_1936);
or U2950 (N_2950,N_2272,N_2146);
or U2951 (N_2951,N_2081,N_1883);
xor U2952 (N_2952,N_2005,N_2326);
and U2953 (N_2953,N_2131,N_2336);
nand U2954 (N_2954,N_2221,N_1930);
nand U2955 (N_2955,N_2118,N_2330);
or U2956 (N_2956,N_2362,N_1926);
and U2957 (N_2957,N_2399,N_2272);
nor U2958 (N_2958,N_2122,N_2146);
nor U2959 (N_2959,N_2322,N_1935);
or U2960 (N_2960,N_1873,N_1942);
or U2961 (N_2961,N_2081,N_1864);
or U2962 (N_2962,N_2114,N_1986);
and U2963 (N_2963,N_1939,N_1892);
or U2964 (N_2964,N_2211,N_2087);
nand U2965 (N_2965,N_1911,N_1884);
xnor U2966 (N_2966,N_2135,N_2028);
nand U2967 (N_2967,N_2159,N_1938);
nand U2968 (N_2968,N_2218,N_2322);
nor U2969 (N_2969,N_2290,N_2329);
nor U2970 (N_2970,N_1919,N_2158);
nor U2971 (N_2971,N_2017,N_2247);
or U2972 (N_2972,N_2247,N_2103);
and U2973 (N_2973,N_1916,N_2059);
and U2974 (N_2974,N_2196,N_2096);
and U2975 (N_2975,N_2270,N_2068);
xor U2976 (N_2976,N_1971,N_1973);
or U2977 (N_2977,N_2078,N_1810);
or U2978 (N_2978,N_1949,N_2196);
and U2979 (N_2979,N_2196,N_2282);
nand U2980 (N_2980,N_2193,N_1812);
nor U2981 (N_2981,N_1854,N_2015);
nor U2982 (N_2982,N_2283,N_2176);
and U2983 (N_2983,N_2224,N_1917);
xnor U2984 (N_2984,N_2029,N_1837);
and U2985 (N_2985,N_1854,N_2163);
and U2986 (N_2986,N_2353,N_2233);
nor U2987 (N_2987,N_2167,N_2344);
or U2988 (N_2988,N_2301,N_1858);
nand U2989 (N_2989,N_2138,N_1923);
nor U2990 (N_2990,N_1852,N_2135);
or U2991 (N_2991,N_2175,N_1870);
and U2992 (N_2992,N_1832,N_2151);
or U2993 (N_2993,N_1907,N_2171);
or U2994 (N_2994,N_2275,N_1849);
nor U2995 (N_2995,N_1993,N_2137);
nand U2996 (N_2996,N_1961,N_2050);
and U2997 (N_2997,N_2178,N_2068);
or U2998 (N_2998,N_2299,N_2259);
or U2999 (N_2999,N_2162,N_2120);
or UO_0 (O_0,N_2538,N_2460);
nor UO_1 (O_1,N_2976,N_2753);
nor UO_2 (O_2,N_2447,N_2959);
and UO_3 (O_3,N_2663,N_2672);
nand UO_4 (O_4,N_2895,N_2838);
or UO_5 (O_5,N_2806,N_2691);
nor UO_6 (O_6,N_2519,N_2665);
and UO_7 (O_7,N_2795,N_2891);
or UO_8 (O_8,N_2690,N_2751);
nor UO_9 (O_9,N_2905,N_2455);
and UO_10 (O_10,N_2513,N_2743);
nand UO_11 (O_11,N_2523,N_2558);
and UO_12 (O_12,N_2869,N_2479);
nor UO_13 (O_13,N_2956,N_2821);
xor UO_14 (O_14,N_2733,N_2585);
nand UO_15 (O_15,N_2598,N_2920);
nand UO_16 (O_16,N_2911,N_2488);
or UO_17 (O_17,N_2605,N_2704);
nand UO_18 (O_18,N_2910,N_2796);
or UO_19 (O_19,N_2638,N_2937);
nand UO_20 (O_20,N_2689,N_2909);
nor UO_21 (O_21,N_2531,N_2450);
nor UO_22 (O_22,N_2584,N_2773);
or UO_23 (O_23,N_2422,N_2565);
or UO_24 (O_24,N_2681,N_2483);
nand UO_25 (O_25,N_2501,N_2781);
and UO_26 (O_26,N_2514,N_2544);
and UO_27 (O_27,N_2946,N_2508);
xnor UO_28 (O_28,N_2750,N_2746);
or UO_29 (O_29,N_2504,N_2988);
nor UO_30 (O_30,N_2581,N_2683);
and UO_31 (O_31,N_2528,N_2768);
nor UO_32 (O_32,N_2694,N_2735);
or UO_33 (O_33,N_2809,N_2529);
nand UO_34 (O_34,N_2440,N_2530);
or UO_35 (O_35,N_2614,N_2702);
nand UO_36 (O_36,N_2679,N_2968);
xnor UO_37 (O_37,N_2548,N_2520);
and UO_38 (O_38,N_2729,N_2426);
nand UO_39 (O_39,N_2668,N_2960);
nor UO_40 (O_40,N_2433,N_2536);
or UO_41 (O_41,N_2493,N_2557);
or UO_42 (O_42,N_2606,N_2687);
nand UO_43 (O_43,N_2772,N_2967);
nand UO_44 (O_44,N_2963,N_2686);
nand UO_45 (O_45,N_2862,N_2715);
and UO_46 (O_46,N_2877,N_2471);
or UO_47 (O_47,N_2794,N_2615);
nor UO_48 (O_48,N_2873,N_2936);
or UO_49 (O_49,N_2607,N_2637);
or UO_50 (O_50,N_2599,N_2412);
xor UO_51 (O_51,N_2416,N_2660);
nor UO_52 (O_52,N_2926,N_2820);
and UO_53 (O_53,N_2575,N_2823);
nand UO_54 (O_54,N_2849,N_2828);
or UO_55 (O_55,N_2646,N_2600);
and UO_56 (O_56,N_2414,N_2723);
nand UO_57 (O_57,N_2495,N_2973);
and UO_58 (O_58,N_2579,N_2954);
nor UO_59 (O_59,N_2644,N_2512);
nand UO_60 (O_60,N_2618,N_2405);
nand UO_61 (O_61,N_2899,N_2788);
nor UO_62 (O_62,N_2448,N_2658);
and UO_63 (O_63,N_2627,N_2863);
xor UO_64 (O_64,N_2678,N_2650);
nor UO_65 (O_65,N_2943,N_2507);
or UO_66 (O_66,N_2780,N_2952);
nand UO_67 (O_67,N_2940,N_2592);
nor UO_68 (O_68,N_2880,N_2941);
and UO_69 (O_69,N_2874,N_2769);
nor UO_70 (O_70,N_2680,N_2883);
nand UO_71 (O_71,N_2748,N_2760);
or UO_72 (O_72,N_2784,N_2634);
nor UO_73 (O_73,N_2496,N_2609);
and UO_74 (O_74,N_2871,N_2583);
nor UO_75 (O_75,N_2975,N_2935);
or UO_76 (O_76,N_2697,N_2511);
nand UO_77 (O_77,N_2787,N_2930);
and UO_78 (O_78,N_2965,N_2827);
nand UO_79 (O_79,N_2987,N_2861);
nor UO_80 (O_80,N_2664,N_2497);
nand UO_81 (O_81,N_2904,N_2752);
and UO_82 (O_82,N_2986,N_2684);
and UO_83 (O_83,N_2424,N_2813);
nand UO_84 (O_84,N_2503,N_2620);
nor UO_85 (O_85,N_2624,N_2951);
and UO_86 (O_86,N_2983,N_2613);
nand UO_87 (O_87,N_2559,N_2626);
nor UO_88 (O_88,N_2594,N_2586);
and UO_89 (O_89,N_2841,N_2623);
or UO_90 (O_90,N_2535,N_2408);
or UO_91 (O_91,N_2695,N_2649);
nand UO_92 (O_92,N_2725,N_2582);
and UO_93 (O_93,N_2825,N_2742);
xnor UO_94 (O_94,N_2429,N_2853);
nor UO_95 (O_95,N_2984,N_2846);
nand UO_96 (O_96,N_2884,N_2700);
or UO_97 (O_97,N_2947,N_2670);
nor UO_98 (O_98,N_2801,N_2767);
xor UO_99 (O_99,N_2855,N_2716);
or UO_100 (O_100,N_2561,N_2674);
and UO_101 (O_101,N_2766,N_2553);
nand UO_102 (O_102,N_2587,N_2541);
nand UO_103 (O_103,N_2419,N_2761);
nor UO_104 (O_104,N_2992,N_2890);
or UO_105 (O_105,N_2934,N_2982);
nand UO_106 (O_106,N_2696,N_2907);
nand UO_107 (O_107,N_2754,N_2865);
or UO_108 (O_108,N_2518,N_2990);
and UO_109 (O_109,N_2692,N_2738);
nor UO_110 (O_110,N_2453,N_2659);
and UO_111 (O_111,N_2734,N_2791);
nor UO_112 (O_112,N_2554,N_2886);
nand UO_113 (O_113,N_2655,N_2682);
nor UO_114 (O_114,N_2740,N_2532);
nor UO_115 (O_115,N_2506,N_2651);
nand UO_116 (O_116,N_2807,N_2489);
nand UO_117 (O_117,N_2875,N_2601);
nor UO_118 (O_118,N_2434,N_2792);
or UO_119 (O_119,N_2621,N_2906);
nand UO_120 (O_120,N_2510,N_2472);
or UO_121 (O_121,N_2499,N_2549);
and UO_122 (O_122,N_2953,N_2629);
nand UO_123 (O_123,N_2747,N_2402);
nor UO_124 (O_124,N_2677,N_2662);
nand UO_125 (O_125,N_2521,N_2755);
and UO_126 (O_126,N_2491,N_2852);
nor UO_127 (O_127,N_2958,N_2826);
and UO_128 (O_128,N_2957,N_2411);
and UO_129 (O_129,N_2647,N_2654);
nor UO_130 (O_130,N_2915,N_2708);
and UO_131 (O_131,N_2400,N_2616);
and UO_132 (O_132,N_2407,N_2860);
and UO_133 (O_133,N_2591,N_2872);
nor UO_134 (O_134,N_2648,N_2657);
nor UO_135 (O_135,N_2524,N_2949);
nor UO_136 (O_136,N_2597,N_2927);
nor UO_137 (O_137,N_2469,N_2671);
nand UO_138 (O_138,N_2676,N_2573);
nand UO_139 (O_139,N_2569,N_2824);
nand UO_140 (O_140,N_2608,N_2745);
nand UO_141 (O_141,N_2756,N_2439);
nor UO_142 (O_142,N_2685,N_2441);
xnor UO_143 (O_143,N_2759,N_2458);
nor UO_144 (O_144,N_2919,N_2771);
or UO_145 (O_145,N_2570,N_2763);
and UO_146 (O_146,N_2912,N_2913);
xor UO_147 (O_147,N_2485,N_2551);
nand UO_148 (O_148,N_2705,N_2486);
or UO_149 (O_149,N_2580,N_2893);
nor UO_150 (O_150,N_2534,N_2552);
and UO_151 (O_151,N_2818,N_2509);
and UO_152 (O_152,N_2588,N_2526);
nand UO_153 (O_153,N_2466,N_2430);
nor UO_154 (O_154,N_2473,N_2435);
and UO_155 (O_155,N_2834,N_2706);
and UO_156 (O_156,N_2870,N_2892);
nor UO_157 (O_157,N_2989,N_2737);
and UO_158 (O_158,N_2778,N_2793);
or UO_159 (O_159,N_2475,N_2401);
and UO_160 (O_160,N_2639,N_2502);
nand UO_161 (O_161,N_2550,N_2903);
nand UO_162 (O_162,N_2921,N_2437);
or UO_163 (O_163,N_2652,N_2864);
xor UO_164 (O_164,N_2995,N_2720);
or UO_165 (O_165,N_2595,N_2908);
and UO_166 (O_166,N_2850,N_2974);
nand UO_167 (O_167,N_2979,N_2445);
and UO_168 (O_168,N_2642,N_2894);
nor UO_169 (O_169,N_2924,N_2925);
and UO_170 (O_170,N_2463,N_2977);
or UO_171 (O_171,N_2409,N_2836);
and UO_172 (O_172,N_2722,N_2922);
and UO_173 (O_173,N_2882,N_2931);
nand UO_174 (O_174,N_2476,N_2540);
nand UO_175 (O_175,N_2833,N_2785);
or UO_176 (O_176,N_2711,N_2994);
nor UO_177 (O_177,N_2462,N_2403);
or UO_178 (O_178,N_2630,N_2596);
and UO_179 (O_179,N_2449,N_2480);
nand UO_180 (O_180,N_2413,N_2612);
nor UO_181 (O_181,N_2611,N_2467);
or UO_182 (O_182,N_2576,N_2939);
nor UO_183 (O_183,N_2928,N_2802);
nor UO_184 (O_184,N_2633,N_2560);
nand UO_185 (O_185,N_2783,N_2436);
nor UO_186 (O_186,N_2803,N_2970);
nand UO_187 (O_187,N_2537,N_2847);
and UO_188 (O_188,N_2464,N_2428);
and UO_189 (O_189,N_2545,N_2427);
nor UO_190 (O_190,N_2896,N_2902);
nand UO_191 (O_191,N_2574,N_2492);
nand UO_192 (O_192,N_2443,N_2432);
or UO_193 (O_193,N_2942,N_2844);
nand UO_194 (O_194,N_2719,N_2468);
nand UO_195 (O_195,N_2804,N_2993);
nand UO_196 (O_196,N_2800,N_2945);
nand UO_197 (O_197,N_2856,N_2829);
and UO_198 (O_198,N_2969,N_2868);
nand UO_199 (O_199,N_2619,N_2789);
nor UO_200 (O_200,N_2563,N_2693);
nor UO_201 (O_201,N_2730,N_2415);
or UO_202 (O_202,N_2636,N_2516);
and UO_203 (O_203,N_2900,N_2808);
nor UO_204 (O_204,N_2901,N_2562);
nand UO_205 (O_205,N_2765,N_2525);
or UO_206 (O_206,N_2688,N_2840);
nor UO_207 (O_207,N_2878,N_2498);
or UO_208 (O_208,N_2461,N_2567);
nor UO_209 (O_209,N_2452,N_2406);
and UO_210 (O_210,N_2950,N_2811);
or UO_211 (O_211,N_2932,N_2917);
and UO_212 (O_212,N_2887,N_2707);
nor UO_213 (O_213,N_2459,N_2955);
nor UO_214 (O_214,N_2985,N_2972);
nor UO_215 (O_215,N_2490,N_2898);
or UO_216 (O_216,N_2779,N_2617);
nor UO_217 (O_217,N_2423,N_2465);
or UO_218 (O_218,N_2832,N_2799);
nand UO_219 (O_219,N_2656,N_2929);
and UO_220 (O_220,N_2602,N_2709);
xnor UO_221 (O_221,N_2876,N_2640);
nor UO_222 (O_222,N_2918,N_2718);
nand UO_223 (O_223,N_2797,N_2961);
and UO_224 (O_224,N_2845,N_2944);
nor UO_225 (O_225,N_2555,N_2885);
nor UO_226 (O_226,N_2717,N_2888);
and UO_227 (O_227,N_2749,N_2425);
nand UO_228 (O_228,N_2482,N_2522);
nand UO_229 (O_229,N_2736,N_2810);
nand UO_230 (O_230,N_2487,N_2431);
and UO_231 (O_231,N_2782,N_2835);
nor UO_232 (O_232,N_2542,N_2698);
or UO_233 (O_233,N_2744,N_2857);
nor UO_234 (O_234,N_2699,N_2661);
nand UO_235 (O_235,N_2966,N_2997);
and UO_236 (O_236,N_2572,N_2964);
and UO_237 (O_237,N_2631,N_2484);
and UO_238 (O_238,N_2675,N_2477);
and UO_239 (O_239,N_2446,N_2547);
nor UO_240 (O_240,N_2897,N_2478);
or UO_241 (O_241,N_2645,N_2666);
nor UO_242 (O_242,N_2669,N_2933);
nand UO_243 (O_243,N_2978,N_2643);
nor UO_244 (O_244,N_2991,N_2938);
nor UO_245 (O_245,N_2815,N_2577);
nor UO_246 (O_246,N_2632,N_2854);
or UO_247 (O_247,N_2420,N_2816);
or UO_248 (O_248,N_2590,N_2962);
and UO_249 (O_249,N_2971,N_2879);
nor UO_250 (O_250,N_2517,N_2775);
nor UO_251 (O_251,N_2859,N_2851);
nor UO_252 (O_252,N_2653,N_2527);
or UO_253 (O_253,N_2712,N_2474);
or UO_254 (O_254,N_2757,N_2604);
and UO_255 (O_255,N_2673,N_2889);
nand UO_256 (O_256,N_2814,N_2451);
and UO_257 (O_257,N_2457,N_2539);
or UO_258 (O_258,N_2830,N_2721);
and UO_259 (O_259,N_2500,N_2593);
or UO_260 (O_260,N_2566,N_2404);
and UO_261 (O_261,N_2843,N_2418);
or UO_262 (O_262,N_2635,N_2837);
and UO_263 (O_263,N_2777,N_2948);
nand UO_264 (O_264,N_2724,N_2831);
and UO_265 (O_265,N_2641,N_2494);
nand UO_266 (O_266,N_2710,N_2858);
nor UO_267 (O_267,N_2739,N_2438);
nand UO_268 (O_268,N_2442,N_2625);
and UO_269 (O_269,N_2764,N_2533);
and UO_270 (O_270,N_2564,N_2505);
nand UO_271 (O_271,N_2470,N_2667);
nor UO_272 (O_272,N_2568,N_2776);
or UO_273 (O_273,N_2543,N_2881);
nor UO_274 (O_274,N_2714,N_2822);
xnor UO_275 (O_275,N_2603,N_2812);
and UO_276 (O_276,N_2546,N_2410);
or UO_277 (O_277,N_2628,N_2914);
nor UO_278 (O_278,N_2713,N_2732);
nor UO_279 (O_279,N_2727,N_2578);
or UO_280 (O_280,N_2556,N_2798);
and UO_281 (O_281,N_2774,N_2421);
and UO_282 (O_282,N_2726,N_2703);
and UO_283 (O_283,N_2916,N_2999);
nor UO_284 (O_284,N_2867,N_2998);
nor UO_285 (O_285,N_2454,N_2786);
and UO_286 (O_286,N_2728,N_2701);
and UO_287 (O_287,N_2790,N_2923);
and UO_288 (O_288,N_2456,N_2762);
nand UO_289 (O_289,N_2770,N_2839);
nor UO_290 (O_290,N_2444,N_2980);
xor UO_291 (O_291,N_2622,N_2481);
nor UO_292 (O_292,N_2819,N_2589);
and UO_293 (O_293,N_2996,N_2866);
nor UO_294 (O_294,N_2571,N_2817);
nor UO_295 (O_295,N_2848,N_2731);
nand UO_296 (O_296,N_2417,N_2741);
nor UO_297 (O_297,N_2610,N_2758);
and UO_298 (O_298,N_2515,N_2805);
and UO_299 (O_299,N_2981,N_2842);
and UO_300 (O_300,N_2783,N_2428);
or UO_301 (O_301,N_2686,N_2856);
nor UO_302 (O_302,N_2896,N_2654);
and UO_303 (O_303,N_2484,N_2856);
and UO_304 (O_304,N_2599,N_2499);
and UO_305 (O_305,N_2644,N_2540);
or UO_306 (O_306,N_2677,N_2737);
nor UO_307 (O_307,N_2878,N_2681);
nor UO_308 (O_308,N_2451,N_2418);
nand UO_309 (O_309,N_2464,N_2921);
and UO_310 (O_310,N_2575,N_2984);
and UO_311 (O_311,N_2889,N_2916);
and UO_312 (O_312,N_2533,N_2900);
nand UO_313 (O_313,N_2449,N_2953);
nand UO_314 (O_314,N_2657,N_2425);
nor UO_315 (O_315,N_2585,N_2445);
nor UO_316 (O_316,N_2628,N_2581);
nor UO_317 (O_317,N_2586,N_2460);
and UO_318 (O_318,N_2591,N_2815);
and UO_319 (O_319,N_2974,N_2498);
or UO_320 (O_320,N_2644,N_2499);
and UO_321 (O_321,N_2434,N_2721);
or UO_322 (O_322,N_2415,N_2884);
and UO_323 (O_323,N_2795,N_2445);
nor UO_324 (O_324,N_2991,N_2541);
xor UO_325 (O_325,N_2759,N_2844);
or UO_326 (O_326,N_2807,N_2573);
nor UO_327 (O_327,N_2956,N_2610);
and UO_328 (O_328,N_2559,N_2547);
nand UO_329 (O_329,N_2426,N_2770);
and UO_330 (O_330,N_2478,N_2487);
nor UO_331 (O_331,N_2432,N_2541);
nand UO_332 (O_332,N_2787,N_2877);
nor UO_333 (O_333,N_2400,N_2540);
nor UO_334 (O_334,N_2587,N_2798);
nand UO_335 (O_335,N_2956,N_2552);
nor UO_336 (O_336,N_2742,N_2852);
nor UO_337 (O_337,N_2524,N_2798);
and UO_338 (O_338,N_2448,N_2843);
and UO_339 (O_339,N_2852,N_2629);
and UO_340 (O_340,N_2414,N_2687);
or UO_341 (O_341,N_2835,N_2418);
or UO_342 (O_342,N_2443,N_2723);
or UO_343 (O_343,N_2752,N_2981);
xnor UO_344 (O_344,N_2854,N_2654);
or UO_345 (O_345,N_2419,N_2718);
and UO_346 (O_346,N_2584,N_2460);
or UO_347 (O_347,N_2665,N_2926);
nand UO_348 (O_348,N_2673,N_2839);
or UO_349 (O_349,N_2780,N_2973);
nand UO_350 (O_350,N_2547,N_2576);
or UO_351 (O_351,N_2416,N_2592);
nand UO_352 (O_352,N_2476,N_2802);
nor UO_353 (O_353,N_2697,N_2571);
and UO_354 (O_354,N_2558,N_2470);
nor UO_355 (O_355,N_2638,N_2810);
xnor UO_356 (O_356,N_2515,N_2827);
nand UO_357 (O_357,N_2445,N_2937);
and UO_358 (O_358,N_2911,N_2993);
and UO_359 (O_359,N_2737,N_2963);
and UO_360 (O_360,N_2417,N_2534);
or UO_361 (O_361,N_2433,N_2799);
or UO_362 (O_362,N_2481,N_2557);
nand UO_363 (O_363,N_2840,N_2976);
and UO_364 (O_364,N_2901,N_2983);
and UO_365 (O_365,N_2654,N_2625);
nand UO_366 (O_366,N_2517,N_2753);
nand UO_367 (O_367,N_2644,N_2406);
nand UO_368 (O_368,N_2465,N_2637);
nand UO_369 (O_369,N_2644,N_2464);
nor UO_370 (O_370,N_2445,N_2820);
nand UO_371 (O_371,N_2848,N_2769);
nor UO_372 (O_372,N_2743,N_2763);
nor UO_373 (O_373,N_2909,N_2511);
or UO_374 (O_374,N_2595,N_2645);
nor UO_375 (O_375,N_2615,N_2503);
nor UO_376 (O_376,N_2481,N_2582);
nor UO_377 (O_377,N_2998,N_2805);
nand UO_378 (O_378,N_2817,N_2641);
nand UO_379 (O_379,N_2511,N_2404);
nor UO_380 (O_380,N_2908,N_2769);
nor UO_381 (O_381,N_2678,N_2952);
or UO_382 (O_382,N_2678,N_2665);
nand UO_383 (O_383,N_2517,N_2727);
or UO_384 (O_384,N_2573,N_2791);
nor UO_385 (O_385,N_2415,N_2854);
nand UO_386 (O_386,N_2603,N_2539);
xor UO_387 (O_387,N_2513,N_2432);
nand UO_388 (O_388,N_2717,N_2494);
and UO_389 (O_389,N_2444,N_2879);
nor UO_390 (O_390,N_2830,N_2564);
and UO_391 (O_391,N_2851,N_2767);
or UO_392 (O_392,N_2788,N_2662);
or UO_393 (O_393,N_2559,N_2940);
or UO_394 (O_394,N_2481,N_2606);
nor UO_395 (O_395,N_2605,N_2717);
nor UO_396 (O_396,N_2664,N_2511);
nor UO_397 (O_397,N_2850,N_2667);
and UO_398 (O_398,N_2448,N_2720);
nand UO_399 (O_399,N_2641,N_2978);
nand UO_400 (O_400,N_2913,N_2972);
or UO_401 (O_401,N_2863,N_2723);
or UO_402 (O_402,N_2767,N_2431);
nor UO_403 (O_403,N_2831,N_2799);
or UO_404 (O_404,N_2785,N_2497);
nand UO_405 (O_405,N_2913,N_2884);
and UO_406 (O_406,N_2749,N_2851);
or UO_407 (O_407,N_2745,N_2702);
nand UO_408 (O_408,N_2471,N_2726);
nand UO_409 (O_409,N_2970,N_2776);
xnor UO_410 (O_410,N_2772,N_2830);
nor UO_411 (O_411,N_2517,N_2574);
xnor UO_412 (O_412,N_2947,N_2601);
or UO_413 (O_413,N_2880,N_2437);
and UO_414 (O_414,N_2742,N_2724);
or UO_415 (O_415,N_2815,N_2475);
nand UO_416 (O_416,N_2591,N_2731);
or UO_417 (O_417,N_2812,N_2568);
nand UO_418 (O_418,N_2563,N_2603);
and UO_419 (O_419,N_2651,N_2504);
nor UO_420 (O_420,N_2985,N_2560);
nand UO_421 (O_421,N_2707,N_2877);
nand UO_422 (O_422,N_2996,N_2641);
and UO_423 (O_423,N_2492,N_2415);
and UO_424 (O_424,N_2808,N_2593);
or UO_425 (O_425,N_2463,N_2688);
and UO_426 (O_426,N_2637,N_2600);
or UO_427 (O_427,N_2982,N_2679);
nor UO_428 (O_428,N_2792,N_2584);
nor UO_429 (O_429,N_2956,N_2974);
nand UO_430 (O_430,N_2623,N_2913);
and UO_431 (O_431,N_2969,N_2695);
nand UO_432 (O_432,N_2750,N_2861);
nand UO_433 (O_433,N_2716,N_2453);
and UO_434 (O_434,N_2641,N_2519);
nand UO_435 (O_435,N_2813,N_2601);
xnor UO_436 (O_436,N_2923,N_2589);
nor UO_437 (O_437,N_2999,N_2712);
nand UO_438 (O_438,N_2879,N_2537);
nor UO_439 (O_439,N_2811,N_2962);
or UO_440 (O_440,N_2947,N_2985);
and UO_441 (O_441,N_2961,N_2457);
nor UO_442 (O_442,N_2923,N_2421);
and UO_443 (O_443,N_2930,N_2811);
nand UO_444 (O_444,N_2683,N_2633);
and UO_445 (O_445,N_2983,N_2576);
nor UO_446 (O_446,N_2665,N_2633);
or UO_447 (O_447,N_2786,N_2801);
or UO_448 (O_448,N_2796,N_2929);
and UO_449 (O_449,N_2763,N_2914);
nor UO_450 (O_450,N_2691,N_2409);
nand UO_451 (O_451,N_2407,N_2861);
nand UO_452 (O_452,N_2746,N_2918);
and UO_453 (O_453,N_2672,N_2738);
or UO_454 (O_454,N_2522,N_2542);
nand UO_455 (O_455,N_2976,N_2762);
nand UO_456 (O_456,N_2801,N_2566);
or UO_457 (O_457,N_2910,N_2746);
or UO_458 (O_458,N_2471,N_2643);
or UO_459 (O_459,N_2939,N_2465);
nand UO_460 (O_460,N_2960,N_2522);
nor UO_461 (O_461,N_2513,N_2589);
nor UO_462 (O_462,N_2860,N_2511);
and UO_463 (O_463,N_2510,N_2622);
nor UO_464 (O_464,N_2549,N_2770);
or UO_465 (O_465,N_2976,N_2643);
xnor UO_466 (O_466,N_2779,N_2666);
nand UO_467 (O_467,N_2575,N_2997);
or UO_468 (O_468,N_2984,N_2905);
nor UO_469 (O_469,N_2462,N_2488);
nand UO_470 (O_470,N_2741,N_2596);
or UO_471 (O_471,N_2712,N_2986);
and UO_472 (O_472,N_2466,N_2852);
and UO_473 (O_473,N_2531,N_2846);
nor UO_474 (O_474,N_2914,N_2799);
nand UO_475 (O_475,N_2831,N_2774);
nor UO_476 (O_476,N_2908,N_2487);
or UO_477 (O_477,N_2805,N_2555);
and UO_478 (O_478,N_2834,N_2951);
nand UO_479 (O_479,N_2823,N_2811);
or UO_480 (O_480,N_2670,N_2474);
or UO_481 (O_481,N_2960,N_2873);
nor UO_482 (O_482,N_2645,N_2550);
and UO_483 (O_483,N_2648,N_2565);
nand UO_484 (O_484,N_2852,N_2870);
xor UO_485 (O_485,N_2816,N_2582);
and UO_486 (O_486,N_2745,N_2513);
or UO_487 (O_487,N_2572,N_2710);
nand UO_488 (O_488,N_2631,N_2514);
nor UO_489 (O_489,N_2535,N_2915);
and UO_490 (O_490,N_2433,N_2515);
nor UO_491 (O_491,N_2871,N_2519);
and UO_492 (O_492,N_2697,N_2640);
or UO_493 (O_493,N_2848,N_2775);
or UO_494 (O_494,N_2526,N_2472);
and UO_495 (O_495,N_2522,N_2718);
and UO_496 (O_496,N_2762,N_2452);
nand UO_497 (O_497,N_2902,N_2839);
nand UO_498 (O_498,N_2752,N_2875);
or UO_499 (O_499,N_2912,N_2674);
endmodule